
module mult_N256_CC256 ( clk, rst, g_input, e_input, o );
  input [255:0] g_input;
  input [0:0] e_input;
  output [511:0] o;
  input clk, rst;
  wire   \add_42/carry[511] , \add_42/carry[510] , \add_42/carry[509] ,
         \add_42/carry[508] , \add_42/carry[507] , \add_42/carry[506] ,
         \add_42/carry[505] , \add_42/carry[504] , \add_42/carry[503] ,
         \add_42/carry[502] , \add_42/carry[501] , \add_42/carry[500] ,
         \add_42/carry[499] , \add_42/carry[498] , \add_42/carry[497] ,
         \add_42/carry[496] , \add_42/carry[495] , \add_42/carry[494] ,
         \add_42/carry[493] , \add_42/carry[492] , \add_42/carry[491] ,
         \add_42/carry[490] , \add_42/carry[489] , \add_42/carry[488] ,
         \add_42/carry[487] , \add_42/carry[486] , \add_42/carry[485] ,
         \add_42/carry[484] , \add_42/carry[483] , \add_42/carry[482] ,
         \add_42/carry[481] , \add_42/carry[480] , \add_42/carry[479] ,
         \add_42/carry[478] , \add_42/carry[477] , \add_42/carry[476] ,
         \add_42/carry[475] , \add_42/carry[474] , \add_42/carry[473] ,
         \add_42/carry[472] , \add_42/carry[471] , \add_42/carry[470] ,
         \add_42/carry[469] , \add_42/carry[468] , \add_42/carry[467] ,
         \add_42/carry[466] , \add_42/carry[465] , \add_42/carry[464] ,
         \add_42/carry[463] , \add_42/carry[462] , \add_42/carry[461] ,
         \add_42/carry[460] , \add_42/carry[459] , \add_42/carry[458] ,
         \add_42/carry[457] , \add_42/carry[456] , \add_42/carry[455] ,
         \add_42/carry[454] , \add_42/carry[453] , \add_42/carry[452] ,
         \add_42/carry[451] , \add_42/carry[450] , \add_42/carry[449] ,
         \add_42/carry[448] , \add_42/carry[447] , \add_42/carry[446] ,
         \add_42/carry[445] , \add_42/carry[444] , \add_42/carry[443] ,
         \add_42/carry[442] , \add_42/carry[441] , \add_42/carry[440] ,
         \add_42/carry[439] , \add_42/carry[438] , \add_42/carry[437] ,
         \add_42/carry[436] , \add_42/carry[435] , \add_42/carry[434] ,
         \add_42/carry[433] , \add_42/carry[432] , \add_42/carry[431] ,
         \add_42/carry[430] , \add_42/carry[429] , \add_42/carry[428] ,
         \add_42/carry[427] , \add_42/carry[426] , \add_42/carry[425] ,
         \add_42/carry[424] , \add_42/carry[423] , \add_42/carry[422] ,
         \add_42/carry[421] , \add_42/carry[420] , \add_42/carry[419] ,
         \add_42/carry[418] , \add_42/carry[417] , \add_42/carry[416] ,
         \add_42/carry[415] , \add_42/carry[414] , \add_42/carry[413] ,
         \add_42/carry[412] , \add_42/carry[411] , \add_42/carry[410] ,
         \add_42/carry[409] , \add_42/carry[408] , \add_42/carry[407] ,
         \add_42/carry[406] , \add_42/carry[405] , \add_42/carry[404] ,
         \add_42/carry[403] , \add_42/carry[402] , \add_42/carry[401] ,
         \add_42/carry[400] , \add_42/carry[399] , \add_42/carry[398] ,
         \add_42/carry[397] , \add_42/carry[396] , \add_42/carry[395] ,
         \add_42/carry[394] , \add_42/carry[393] , \add_42/carry[392] ,
         \add_42/carry[391] , \add_42/carry[390] , \add_42/carry[389] ,
         \add_42/carry[388] , \add_42/carry[387] , \add_42/carry[386] ,
         \add_42/carry[385] , \add_42/carry[384] , \add_42/carry[383] ,
         \add_42/carry[382] , \add_42/carry[381] , \add_42/carry[380] ,
         \add_42/carry[379] , \add_42/carry[378] , \add_42/carry[377] ,
         \add_42/carry[376] , \add_42/carry[375] , \add_42/carry[374] ,
         \add_42/carry[373] , \add_42/carry[372] , \add_42/carry[371] ,
         \add_42/carry[370] , \add_42/carry[369] , \add_42/carry[368] ,
         \add_42/carry[367] , \add_42/carry[366] , \add_42/carry[365] ,
         \add_42/carry[364] , \add_42/carry[363] , \add_42/carry[362] ,
         \add_42/carry[361] , \add_42/carry[360] , \add_42/carry[359] ,
         \add_42/carry[358] , \add_42/carry[357] , \add_42/carry[356] ,
         \add_42/carry[355] , \add_42/carry[354] , \add_42/carry[353] ,
         \add_42/carry[352] , \add_42/carry[351] , \add_42/carry[350] ,
         \add_42/carry[349] , \add_42/carry[348] , \add_42/carry[347] ,
         \add_42/carry[346] , \add_42/carry[345] , \add_42/carry[344] ,
         \add_42/carry[343] , \add_42/carry[342] , \add_42/carry[341] ,
         \add_42/carry[340] , \add_42/carry[339] , \add_42/carry[338] ,
         \add_42/carry[337] , \add_42/carry[336] , \add_42/carry[335] ,
         \add_42/carry[334] , \add_42/carry[333] , \add_42/carry[332] ,
         \add_42/carry[331] , \add_42/carry[330] , \add_42/carry[329] ,
         \add_42/carry[328] , \add_42/carry[327] , \add_42/carry[326] ,
         \add_42/carry[325] , \add_42/carry[324] , \add_42/carry[323] ,
         \add_42/carry[322] , \add_42/carry[321] , \add_42/carry[320] ,
         \add_42/carry[319] , \add_42/carry[318] , \add_42/carry[317] ,
         \add_42/carry[316] , \add_42/carry[315] , \add_42/carry[314] ,
         \add_42/carry[313] , \add_42/carry[312] , \add_42/carry[311] ,
         \add_42/carry[310] , \add_42/carry[309] , \add_42/carry[308] ,
         \add_42/carry[307] , \add_42/carry[306] , \add_42/carry[305] ,
         \add_42/carry[304] , \add_42/carry[303] , \add_42/carry[302] ,
         \add_42/carry[301] , \add_42/carry[300] , \add_42/carry[299] ,
         \add_42/carry[298] , \add_42/carry[297] , \add_42/carry[296] ,
         \add_42/carry[295] , \add_42/carry[294] , \add_42/carry[293] ,
         \add_42/carry[292] , \add_42/carry[291] , \add_42/carry[290] ,
         \add_42/carry[289] , \add_42/carry[288] , \add_42/carry[287] ,
         \add_42/carry[286] , \add_42/carry[285] , \add_42/carry[284] ,
         \add_42/carry[283] , \add_42/carry[282] , \add_42/carry[281] ,
         \add_42/carry[280] , \add_42/carry[279] , \add_42/carry[278] ,
         \add_42/carry[277] , \add_42/carry[276] , \add_42/carry[275] ,
         \add_42/carry[274] , \add_42/carry[273] , \add_42/carry[272] ,
         \add_42/carry[271] , \add_42/carry[270] , \add_42/carry[269] ,
         \add_42/carry[268] , \add_42/carry[267] , \add_42/carry[266] ,
         \add_42/carry[265] , \add_42/carry[264] , \add_42/carry[263] ,
         \add_42/carry[262] , \add_42/carry[261] , \add_42/carry[260] ,
         \add_42/carry[259] , \add_42/carry[258] , \add_42/carry[257] ,
         \add_42/carry[256] , n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769;
  wire   [511:0] sreg;
  assign o[254] = sreg[254];
  assign o[253] = sreg[253];
  assign o[252] = sreg[252];
  assign o[251] = sreg[251];
  assign o[250] = sreg[250];
  assign o[249] = sreg[249];
  assign o[248] = sreg[248];
  assign o[247] = sreg[247];
  assign o[246] = sreg[246];
  assign o[245] = sreg[245];
  assign o[244] = sreg[244];
  assign o[243] = sreg[243];
  assign o[242] = sreg[242];
  assign o[241] = sreg[241];
  assign o[240] = sreg[240];
  assign o[239] = sreg[239];
  assign o[238] = sreg[238];
  assign o[237] = sreg[237];
  assign o[236] = sreg[236];
  assign o[235] = sreg[235];
  assign o[234] = sreg[234];
  assign o[233] = sreg[233];
  assign o[232] = sreg[232];
  assign o[231] = sreg[231];
  assign o[230] = sreg[230];
  assign o[229] = sreg[229];
  assign o[228] = sreg[228];
  assign o[227] = sreg[227];
  assign o[226] = sreg[226];
  assign o[225] = sreg[225];
  assign o[224] = sreg[224];
  assign o[223] = sreg[223];
  assign o[222] = sreg[222];
  assign o[221] = sreg[221];
  assign o[220] = sreg[220];
  assign o[219] = sreg[219];
  assign o[218] = sreg[218];
  assign o[217] = sreg[217];
  assign o[216] = sreg[216];
  assign o[215] = sreg[215];
  assign o[214] = sreg[214];
  assign o[213] = sreg[213];
  assign o[212] = sreg[212];
  assign o[211] = sreg[211];
  assign o[210] = sreg[210];
  assign o[209] = sreg[209];
  assign o[208] = sreg[208];
  assign o[207] = sreg[207];
  assign o[206] = sreg[206];
  assign o[205] = sreg[205];
  assign o[204] = sreg[204];
  assign o[203] = sreg[203];
  assign o[202] = sreg[202];
  assign o[201] = sreg[201];
  assign o[200] = sreg[200];
  assign o[199] = sreg[199];
  assign o[198] = sreg[198];
  assign o[197] = sreg[197];
  assign o[196] = sreg[196];
  assign o[195] = sreg[195];
  assign o[194] = sreg[194];
  assign o[193] = sreg[193];
  assign o[192] = sreg[192];
  assign o[191] = sreg[191];
  assign o[190] = sreg[190];
  assign o[189] = sreg[189];
  assign o[188] = sreg[188];
  assign o[187] = sreg[187];
  assign o[186] = sreg[186];
  assign o[185] = sreg[185];
  assign o[184] = sreg[184];
  assign o[183] = sreg[183];
  assign o[182] = sreg[182];
  assign o[181] = sreg[181];
  assign o[180] = sreg[180];
  assign o[179] = sreg[179];
  assign o[178] = sreg[178];
  assign o[177] = sreg[177];
  assign o[176] = sreg[176];
  assign o[175] = sreg[175];
  assign o[174] = sreg[174];
  assign o[173] = sreg[173];
  assign o[172] = sreg[172];
  assign o[171] = sreg[171];
  assign o[170] = sreg[170];
  assign o[169] = sreg[169];
  assign o[168] = sreg[168];
  assign o[167] = sreg[167];
  assign o[166] = sreg[166];
  assign o[165] = sreg[165];
  assign o[164] = sreg[164];
  assign o[163] = sreg[163];
  assign o[162] = sreg[162];
  assign o[161] = sreg[161];
  assign o[160] = sreg[160];
  assign o[159] = sreg[159];
  assign o[158] = sreg[158];
  assign o[157] = sreg[157];
  assign o[156] = sreg[156];
  assign o[155] = sreg[155];
  assign o[154] = sreg[154];
  assign o[153] = sreg[153];
  assign o[152] = sreg[152];
  assign o[151] = sreg[151];
  assign o[150] = sreg[150];
  assign o[149] = sreg[149];
  assign o[148] = sreg[148];
  assign o[147] = sreg[147];
  assign o[146] = sreg[146];
  assign o[145] = sreg[145];
  assign o[144] = sreg[144];
  assign o[143] = sreg[143];
  assign o[142] = sreg[142];
  assign o[141] = sreg[141];
  assign o[140] = sreg[140];
  assign o[139] = sreg[139];
  assign o[138] = sreg[138];
  assign o[137] = sreg[137];
  assign o[136] = sreg[136];
  assign o[135] = sreg[135];
  assign o[134] = sreg[134];
  assign o[133] = sreg[133];
  assign o[132] = sreg[132];
  assign o[131] = sreg[131];
  assign o[130] = sreg[130];
  assign o[129] = sreg[129];
  assign o[128] = sreg[128];
  assign o[127] = sreg[127];
  assign o[126] = sreg[126];
  assign o[125] = sreg[125];
  assign o[124] = sreg[124];
  assign o[123] = sreg[123];
  assign o[122] = sreg[122];
  assign o[121] = sreg[121];
  assign o[120] = sreg[120];
  assign o[119] = sreg[119];
  assign o[118] = sreg[118];
  assign o[117] = sreg[117];
  assign o[116] = sreg[116];
  assign o[115] = sreg[115];
  assign o[114] = sreg[114];
  assign o[113] = sreg[113];
  assign o[112] = sreg[112];
  assign o[111] = sreg[111];
  assign o[110] = sreg[110];
  assign o[109] = sreg[109];
  assign o[108] = sreg[108];
  assign o[107] = sreg[107];
  assign o[106] = sreg[106];
  assign o[105] = sreg[105];
  assign o[104] = sreg[104];
  assign o[103] = sreg[103];
  assign o[102] = sreg[102];
  assign o[101] = sreg[101];
  assign o[100] = sreg[100];
  assign o[99] = sreg[99];
  assign o[98] = sreg[98];
  assign o[97] = sreg[97];
  assign o[96] = sreg[96];
  assign o[95] = sreg[95];
  assign o[94] = sreg[94];
  assign o[93] = sreg[93];
  assign o[92] = sreg[92];
  assign o[91] = sreg[91];
  assign o[90] = sreg[90];
  assign o[89] = sreg[89];
  assign o[88] = sreg[88];
  assign o[87] = sreg[87];
  assign o[86] = sreg[86];
  assign o[85] = sreg[85];
  assign o[84] = sreg[84];
  assign o[83] = sreg[83];
  assign o[82] = sreg[82];
  assign o[81] = sreg[81];
  assign o[80] = sreg[80];
  assign o[79] = sreg[79];
  assign o[78] = sreg[78];
  assign o[77] = sreg[77];
  assign o[76] = sreg[76];
  assign o[75] = sreg[75];
  assign o[74] = sreg[74];
  assign o[73] = sreg[73];
  assign o[72] = sreg[72];
  assign o[71] = sreg[71];
  assign o[70] = sreg[70];
  assign o[69] = sreg[69];
  assign o[68] = sreg[68];
  assign o[67] = sreg[67];
  assign o[66] = sreg[66];
  assign o[65] = sreg[65];
  assign o[64] = sreg[64];
  assign o[63] = sreg[63];
  assign o[62] = sreg[62];
  assign o[61] = sreg[61];
  assign o[60] = sreg[60];
  assign o[59] = sreg[59];
  assign o[58] = sreg[58];
  assign o[57] = sreg[57];
  assign o[56] = sreg[56];
  assign o[55] = sreg[55];
  assign o[54] = sreg[54];
  assign o[53] = sreg[53];
  assign o[52] = sreg[52];
  assign o[51] = sreg[51];
  assign o[50] = sreg[50];
  assign o[49] = sreg[49];
  assign o[48] = sreg[48];
  assign o[47] = sreg[47];
  assign o[46] = sreg[46];
  assign o[45] = sreg[45];
  assign o[44] = sreg[44];
  assign o[43] = sreg[43];
  assign o[42] = sreg[42];
  assign o[41] = sreg[41];
  assign o[40] = sreg[40];
  assign o[39] = sreg[39];
  assign o[38] = sreg[38];
  assign o[37] = sreg[37];
  assign o[36] = sreg[36];
  assign o[35] = sreg[35];
  assign o[34] = sreg[34];
  assign o[33] = sreg[33];
  assign o[32] = sreg[32];
  assign o[31] = sreg[31];
  assign o[30] = sreg[30];
  assign o[29] = sreg[29];
  assign o[28] = sreg[28];
  assign o[27] = sreg[27];
  assign o[26] = sreg[26];
  assign o[25] = sreg[25];
  assign o[24] = sreg[24];
  assign o[23] = sreg[23];
  assign o[22] = sreg[22];
  assign o[21] = sreg[21];
  assign o[20] = sreg[20];
  assign o[19] = sreg[19];
  assign o[18] = sreg[18];
  assign o[17] = sreg[17];
  assign o[16] = sreg[16];
  assign o[15] = sreg[15];
  assign o[14] = sreg[14];
  assign o[13] = sreg[13];
  assign o[12] = sreg[12];
  assign o[11] = sreg[11];
  assign o[10] = sreg[10];
  assign o[9] = sreg[9];
  assign o[8] = sreg[8];
  assign o[7] = sreg[7];
  assign o[6] = sreg[6];
  assign o[5] = sreg[5];
  assign o[4] = sreg[4];
  assign o[3] = sreg[3];
  assign o[2] = sreg[2];
  assign o[1] = sreg[1];
  assign o[511] = \add_42/carry[511] ;

  DFF \sreg_reg[0]  ( .D(sreg[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[0]) );
  DFF \sreg_reg[1]  ( .D(sreg[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[1])
         );
  DFF \sreg_reg[2]  ( .D(sreg[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[2])
         );
  DFF \sreg_reg[3]  ( .D(sreg[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[3])
         );
  DFF \sreg_reg[4]  ( .D(sreg[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[4])
         );
  DFF \sreg_reg[5]  ( .D(sreg[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[5])
         );
  DFF \sreg_reg[6]  ( .D(sreg[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[6])
         );
  DFF \sreg_reg[7]  ( .D(sreg[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[7])
         );
  DFF \sreg_reg[8]  ( .D(sreg[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[8])
         );
  DFF \sreg_reg[9]  ( .D(sreg[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[9]) );
  DFF \sreg_reg[10]  ( .D(sreg[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[10]) );
  DFF \sreg_reg[11]  ( .D(sreg[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[11]) );
  DFF \sreg_reg[12]  ( .D(sreg[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[12]) );
  DFF \sreg_reg[13]  ( .D(sreg[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[13]) );
  DFF \sreg_reg[14]  ( .D(sreg[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[14]) );
  DFF \sreg_reg[15]  ( .D(sreg[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[15]) );
  DFF \sreg_reg[16]  ( .D(sreg[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[16]) );
  DFF \sreg_reg[17]  ( .D(sreg[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[17]) );
  DFF \sreg_reg[18]  ( .D(sreg[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[18]) );
  DFF \sreg_reg[19]  ( .D(sreg[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[19]) );
  DFF \sreg_reg[20]  ( .D(sreg[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[20]) );
  DFF \sreg_reg[21]  ( .D(sreg[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[21]) );
  DFF \sreg_reg[22]  ( .D(sreg[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[22]) );
  DFF \sreg_reg[23]  ( .D(sreg[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[23]) );
  DFF \sreg_reg[24]  ( .D(sreg[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[24]) );
  DFF \sreg_reg[25]  ( .D(sreg[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[25]) );
  DFF \sreg_reg[26]  ( .D(sreg[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[26]) );
  DFF \sreg_reg[27]  ( .D(sreg[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[27]) );
  DFF \sreg_reg[28]  ( .D(sreg[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[28]) );
  DFF \sreg_reg[29]  ( .D(sreg[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[29]) );
  DFF \sreg_reg[30]  ( .D(sreg[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[30]) );
  DFF \sreg_reg[31]  ( .D(sreg[32]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[31]) );
  DFF \sreg_reg[32]  ( .D(sreg[33]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[32]) );
  DFF \sreg_reg[33]  ( .D(sreg[34]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[33]) );
  DFF \sreg_reg[34]  ( .D(sreg[35]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[34]) );
  DFF \sreg_reg[35]  ( .D(sreg[36]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[35]) );
  DFF \sreg_reg[36]  ( .D(sreg[37]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[36]) );
  DFF \sreg_reg[37]  ( .D(sreg[38]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[37]) );
  DFF \sreg_reg[38]  ( .D(sreg[39]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[38]) );
  DFF \sreg_reg[39]  ( .D(sreg[40]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[39]) );
  DFF \sreg_reg[40]  ( .D(sreg[41]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[40]) );
  DFF \sreg_reg[41]  ( .D(sreg[42]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[41]) );
  DFF \sreg_reg[42]  ( .D(sreg[43]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[42]) );
  DFF \sreg_reg[43]  ( .D(sreg[44]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[43]) );
  DFF \sreg_reg[44]  ( .D(sreg[45]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[44]) );
  DFF \sreg_reg[45]  ( .D(sreg[46]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[45]) );
  DFF \sreg_reg[46]  ( .D(sreg[47]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[46]) );
  DFF \sreg_reg[47]  ( .D(sreg[48]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[47]) );
  DFF \sreg_reg[48]  ( .D(sreg[49]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[48]) );
  DFF \sreg_reg[49]  ( .D(sreg[50]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[49]) );
  DFF \sreg_reg[50]  ( .D(sreg[51]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[50]) );
  DFF \sreg_reg[51]  ( .D(sreg[52]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[51]) );
  DFF \sreg_reg[52]  ( .D(sreg[53]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[52]) );
  DFF \sreg_reg[53]  ( .D(sreg[54]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[53]) );
  DFF \sreg_reg[54]  ( .D(sreg[55]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[54]) );
  DFF \sreg_reg[55]  ( .D(sreg[56]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[55]) );
  DFF \sreg_reg[56]  ( .D(sreg[57]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[56]) );
  DFF \sreg_reg[57]  ( .D(sreg[58]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[57]) );
  DFF \sreg_reg[58]  ( .D(sreg[59]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[58]) );
  DFF \sreg_reg[59]  ( .D(sreg[60]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[59]) );
  DFF \sreg_reg[60]  ( .D(sreg[61]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[60]) );
  DFF \sreg_reg[61]  ( .D(sreg[62]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[61]) );
  DFF \sreg_reg[62]  ( .D(sreg[63]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[62]) );
  DFF \sreg_reg[63]  ( .D(sreg[64]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[63]) );
  DFF \sreg_reg[64]  ( .D(sreg[65]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[64]) );
  DFF \sreg_reg[65]  ( .D(sreg[66]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[65]) );
  DFF \sreg_reg[66]  ( .D(sreg[67]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[66]) );
  DFF \sreg_reg[67]  ( .D(sreg[68]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[67]) );
  DFF \sreg_reg[68]  ( .D(sreg[69]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[68]) );
  DFF \sreg_reg[69]  ( .D(sreg[70]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[69]) );
  DFF \sreg_reg[70]  ( .D(sreg[71]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[70]) );
  DFF \sreg_reg[71]  ( .D(sreg[72]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[71]) );
  DFF \sreg_reg[72]  ( .D(sreg[73]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[72]) );
  DFF \sreg_reg[73]  ( .D(sreg[74]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[73]) );
  DFF \sreg_reg[74]  ( .D(sreg[75]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[74]) );
  DFF \sreg_reg[75]  ( .D(sreg[76]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[75]) );
  DFF \sreg_reg[76]  ( .D(sreg[77]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[76]) );
  DFF \sreg_reg[77]  ( .D(sreg[78]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[77]) );
  DFF \sreg_reg[78]  ( .D(sreg[79]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[78]) );
  DFF \sreg_reg[79]  ( .D(sreg[80]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[79]) );
  DFF \sreg_reg[80]  ( .D(sreg[81]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[80]) );
  DFF \sreg_reg[81]  ( .D(sreg[82]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[81]) );
  DFF \sreg_reg[82]  ( .D(sreg[83]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[82]) );
  DFF \sreg_reg[83]  ( .D(sreg[84]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[83]) );
  DFF \sreg_reg[84]  ( .D(sreg[85]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[84]) );
  DFF \sreg_reg[85]  ( .D(sreg[86]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[85]) );
  DFF \sreg_reg[86]  ( .D(sreg[87]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[86]) );
  DFF \sreg_reg[87]  ( .D(sreg[88]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[87]) );
  DFF \sreg_reg[88]  ( .D(sreg[89]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[88]) );
  DFF \sreg_reg[89]  ( .D(sreg[90]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[89]) );
  DFF \sreg_reg[90]  ( .D(sreg[91]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[90]) );
  DFF \sreg_reg[91]  ( .D(sreg[92]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[91]) );
  DFF \sreg_reg[92]  ( .D(sreg[93]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[92]) );
  DFF \sreg_reg[93]  ( .D(sreg[94]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[93]) );
  DFF \sreg_reg[94]  ( .D(sreg[95]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[94]) );
  DFF \sreg_reg[95]  ( .D(sreg[96]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[95]) );
  DFF \sreg_reg[96]  ( .D(sreg[97]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[96]) );
  DFF \sreg_reg[97]  ( .D(sreg[98]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[97]) );
  DFF \sreg_reg[98]  ( .D(sreg[99]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[98]) );
  DFF \sreg_reg[99]  ( .D(sreg[100]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[99]) );
  DFF \sreg_reg[100]  ( .D(sreg[101]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[100]) );
  DFF \sreg_reg[101]  ( .D(sreg[102]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[101]) );
  DFF \sreg_reg[102]  ( .D(sreg[103]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[102]) );
  DFF \sreg_reg[103]  ( .D(sreg[104]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[103]) );
  DFF \sreg_reg[104]  ( .D(sreg[105]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[104]) );
  DFF \sreg_reg[105]  ( .D(sreg[106]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[105]) );
  DFF \sreg_reg[106]  ( .D(sreg[107]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[106]) );
  DFF \sreg_reg[107]  ( .D(sreg[108]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[107]) );
  DFF \sreg_reg[108]  ( .D(sreg[109]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[108]) );
  DFF \sreg_reg[109]  ( .D(sreg[110]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[109]) );
  DFF \sreg_reg[110]  ( .D(sreg[111]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[110]) );
  DFF \sreg_reg[111]  ( .D(sreg[112]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[111]) );
  DFF \sreg_reg[112]  ( .D(sreg[113]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[112]) );
  DFF \sreg_reg[113]  ( .D(sreg[114]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[113]) );
  DFF \sreg_reg[114]  ( .D(sreg[115]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[114]) );
  DFF \sreg_reg[115]  ( .D(sreg[116]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[115]) );
  DFF \sreg_reg[116]  ( .D(sreg[117]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[116]) );
  DFF \sreg_reg[117]  ( .D(sreg[118]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[117]) );
  DFF \sreg_reg[118]  ( .D(sreg[119]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[118]) );
  DFF \sreg_reg[119]  ( .D(sreg[120]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[119]) );
  DFF \sreg_reg[120]  ( .D(sreg[121]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[120]) );
  DFF \sreg_reg[121]  ( .D(sreg[122]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[121]) );
  DFF \sreg_reg[122]  ( .D(sreg[123]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[122]) );
  DFF \sreg_reg[123]  ( .D(sreg[124]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[123]) );
  DFF \sreg_reg[124]  ( .D(sreg[125]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[124]) );
  DFF \sreg_reg[125]  ( .D(sreg[126]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[125]) );
  DFF \sreg_reg[126]  ( .D(sreg[127]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[126]) );
  DFF \sreg_reg[127]  ( .D(sreg[128]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[127]) );
  DFF \sreg_reg[128]  ( .D(sreg[129]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[128]) );
  DFF \sreg_reg[129]  ( .D(sreg[130]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[129]) );
  DFF \sreg_reg[130]  ( .D(sreg[131]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[130]) );
  DFF \sreg_reg[131]  ( .D(sreg[132]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[131]) );
  DFF \sreg_reg[132]  ( .D(sreg[133]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[132]) );
  DFF \sreg_reg[133]  ( .D(sreg[134]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[133]) );
  DFF \sreg_reg[134]  ( .D(sreg[135]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[134]) );
  DFF \sreg_reg[135]  ( .D(sreg[136]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[135]) );
  DFF \sreg_reg[136]  ( .D(sreg[137]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[136]) );
  DFF \sreg_reg[137]  ( .D(sreg[138]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[137]) );
  DFF \sreg_reg[138]  ( .D(sreg[139]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[138]) );
  DFF \sreg_reg[139]  ( .D(sreg[140]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[139]) );
  DFF \sreg_reg[140]  ( .D(sreg[141]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[140]) );
  DFF \sreg_reg[141]  ( .D(sreg[142]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[141]) );
  DFF \sreg_reg[142]  ( .D(sreg[143]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[142]) );
  DFF \sreg_reg[143]  ( .D(sreg[144]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[143]) );
  DFF \sreg_reg[144]  ( .D(sreg[145]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[144]) );
  DFF \sreg_reg[145]  ( .D(sreg[146]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[145]) );
  DFF \sreg_reg[146]  ( .D(sreg[147]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[146]) );
  DFF \sreg_reg[147]  ( .D(sreg[148]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[147]) );
  DFF \sreg_reg[148]  ( .D(sreg[149]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[148]) );
  DFF \sreg_reg[149]  ( .D(sreg[150]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[149]) );
  DFF \sreg_reg[150]  ( .D(sreg[151]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[150]) );
  DFF \sreg_reg[151]  ( .D(sreg[152]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[151]) );
  DFF \sreg_reg[152]  ( .D(sreg[153]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[152]) );
  DFF \sreg_reg[153]  ( .D(sreg[154]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[153]) );
  DFF \sreg_reg[154]  ( .D(sreg[155]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[154]) );
  DFF \sreg_reg[155]  ( .D(sreg[156]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[155]) );
  DFF \sreg_reg[156]  ( .D(sreg[157]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[156]) );
  DFF \sreg_reg[157]  ( .D(sreg[158]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[157]) );
  DFF \sreg_reg[158]  ( .D(sreg[159]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[158]) );
  DFF \sreg_reg[159]  ( .D(sreg[160]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[159]) );
  DFF \sreg_reg[160]  ( .D(sreg[161]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[160]) );
  DFF \sreg_reg[161]  ( .D(sreg[162]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[161]) );
  DFF \sreg_reg[162]  ( .D(sreg[163]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[162]) );
  DFF \sreg_reg[163]  ( .D(sreg[164]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[163]) );
  DFF \sreg_reg[164]  ( .D(sreg[165]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[164]) );
  DFF \sreg_reg[165]  ( .D(sreg[166]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[165]) );
  DFF \sreg_reg[166]  ( .D(sreg[167]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[166]) );
  DFF \sreg_reg[167]  ( .D(sreg[168]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[167]) );
  DFF \sreg_reg[168]  ( .D(sreg[169]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[168]) );
  DFF \sreg_reg[169]  ( .D(sreg[170]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[169]) );
  DFF \sreg_reg[170]  ( .D(sreg[171]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[170]) );
  DFF \sreg_reg[171]  ( .D(sreg[172]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[171]) );
  DFF \sreg_reg[172]  ( .D(sreg[173]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[172]) );
  DFF \sreg_reg[173]  ( .D(sreg[174]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[173]) );
  DFF \sreg_reg[174]  ( .D(sreg[175]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[174]) );
  DFF \sreg_reg[175]  ( .D(sreg[176]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[175]) );
  DFF \sreg_reg[176]  ( .D(sreg[177]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[176]) );
  DFF \sreg_reg[177]  ( .D(sreg[178]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[177]) );
  DFF \sreg_reg[178]  ( .D(sreg[179]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[178]) );
  DFF \sreg_reg[179]  ( .D(sreg[180]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[179]) );
  DFF \sreg_reg[180]  ( .D(sreg[181]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[180]) );
  DFF \sreg_reg[181]  ( .D(sreg[182]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[181]) );
  DFF \sreg_reg[182]  ( .D(sreg[183]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[182]) );
  DFF \sreg_reg[183]  ( .D(sreg[184]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[183]) );
  DFF \sreg_reg[184]  ( .D(sreg[185]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[184]) );
  DFF \sreg_reg[185]  ( .D(sreg[186]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[185]) );
  DFF \sreg_reg[186]  ( .D(sreg[187]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[186]) );
  DFF \sreg_reg[187]  ( .D(sreg[188]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[187]) );
  DFF \sreg_reg[188]  ( .D(sreg[189]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[188]) );
  DFF \sreg_reg[189]  ( .D(sreg[190]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[189]) );
  DFF \sreg_reg[190]  ( .D(sreg[191]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[190]) );
  DFF \sreg_reg[191]  ( .D(sreg[192]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[191]) );
  DFF \sreg_reg[192]  ( .D(sreg[193]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[192]) );
  DFF \sreg_reg[193]  ( .D(sreg[194]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[193]) );
  DFF \sreg_reg[194]  ( .D(sreg[195]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[194]) );
  DFF \sreg_reg[195]  ( .D(sreg[196]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[195]) );
  DFF \sreg_reg[196]  ( .D(sreg[197]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[196]) );
  DFF \sreg_reg[197]  ( .D(sreg[198]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[197]) );
  DFF \sreg_reg[198]  ( .D(sreg[199]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[198]) );
  DFF \sreg_reg[199]  ( .D(sreg[200]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[199]) );
  DFF \sreg_reg[200]  ( .D(sreg[201]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[200]) );
  DFF \sreg_reg[201]  ( .D(sreg[202]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[201]) );
  DFF \sreg_reg[202]  ( .D(sreg[203]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[202]) );
  DFF \sreg_reg[203]  ( .D(sreg[204]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[203]) );
  DFF \sreg_reg[204]  ( .D(sreg[205]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[204]) );
  DFF \sreg_reg[205]  ( .D(sreg[206]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[205]) );
  DFF \sreg_reg[206]  ( .D(sreg[207]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[206]) );
  DFF \sreg_reg[207]  ( .D(sreg[208]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[207]) );
  DFF \sreg_reg[208]  ( .D(sreg[209]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[208]) );
  DFF \sreg_reg[209]  ( .D(sreg[210]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[209]) );
  DFF \sreg_reg[210]  ( .D(sreg[211]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[210]) );
  DFF \sreg_reg[211]  ( .D(sreg[212]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[211]) );
  DFF \sreg_reg[212]  ( .D(sreg[213]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[212]) );
  DFF \sreg_reg[213]  ( .D(sreg[214]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[213]) );
  DFF \sreg_reg[214]  ( .D(sreg[215]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[214]) );
  DFF \sreg_reg[215]  ( .D(sreg[216]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[215]) );
  DFF \sreg_reg[216]  ( .D(sreg[217]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[216]) );
  DFF \sreg_reg[217]  ( .D(sreg[218]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[217]) );
  DFF \sreg_reg[218]  ( .D(sreg[219]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[218]) );
  DFF \sreg_reg[219]  ( .D(sreg[220]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[219]) );
  DFF \sreg_reg[220]  ( .D(sreg[221]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[220]) );
  DFF \sreg_reg[221]  ( .D(sreg[222]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[221]) );
  DFF \sreg_reg[222]  ( .D(sreg[223]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[222]) );
  DFF \sreg_reg[223]  ( .D(sreg[224]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[223]) );
  DFF \sreg_reg[224]  ( .D(sreg[225]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[224]) );
  DFF \sreg_reg[225]  ( .D(sreg[226]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[225]) );
  DFF \sreg_reg[226]  ( .D(sreg[227]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[226]) );
  DFF \sreg_reg[227]  ( .D(sreg[228]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[227]) );
  DFF \sreg_reg[228]  ( .D(sreg[229]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[228]) );
  DFF \sreg_reg[229]  ( .D(sreg[230]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[229]) );
  DFF \sreg_reg[230]  ( .D(sreg[231]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[230]) );
  DFF \sreg_reg[231]  ( .D(sreg[232]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[231]) );
  DFF \sreg_reg[232]  ( .D(sreg[233]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[232]) );
  DFF \sreg_reg[233]  ( .D(sreg[234]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[233]) );
  DFF \sreg_reg[234]  ( .D(sreg[235]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[234]) );
  DFF \sreg_reg[235]  ( .D(sreg[236]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[235]) );
  DFF \sreg_reg[236]  ( .D(sreg[237]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[236]) );
  DFF \sreg_reg[237]  ( .D(sreg[238]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[237]) );
  DFF \sreg_reg[238]  ( .D(sreg[239]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[238]) );
  DFF \sreg_reg[239]  ( .D(sreg[240]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[239]) );
  DFF \sreg_reg[240]  ( .D(sreg[241]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[240]) );
  DFF \sreg_reg[241]  ( .D(sreg[242]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[241]) );
  DFF \sreg_reg[242]  ( .D(sreg[243]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[242]) );
  DFF \sreg_reg[243]  ( .D(sreg[244]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[243]) );
  DFF \sreg_reg[244]  ( .D(sreg[245]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[244]) );
  DFF \sreg_reg[245]  ( .D(sreg[246]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[245]) );
  DFF \sreg_reg[246]  ( .D(sreg[247]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[246]) );
  DFF \sreg_reg[247]  ( .D(sreg[248]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[247]) );
  DFF \sreg_reg[248]  ( .D(sreg[249]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[248]) );
  DFF \sreg_reg[249]  ( .D(sreg[250]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[249]) );
  DFF \sreg_reg[250]  ( .D(sreg[251]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[250]) );
  DFF \sreg_reg[251]  ( .D(sreg[252]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[251]) );
  DFF \sreg_reg[252]  ( .D(sreg[253]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[252]) );
  DFF \sreg_reg[253]  ( .D(sreg[254]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[253]) );
  DFF \sreg_reg[254]  ( .D(o[255]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[254]) );
  DFF \sreg_reg[255]  ( .D(o[256]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[255]) );
  DFF \sreg_reg[256]  ( .D(o[257]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[256]) );
  DFF \sreg_reg[257]  ( .D(o[258]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[257]) );
  DFF \sreg_reg[258]  ( .D(o[259]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[258]) );
  DFF \sreg_reg[259]  ( .D(o[260]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[259]) );
  DFF \sreg_reg[260]  ( .D(o[261]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[260]) );
  DFF \sreg_reg[261]  ( .D(o[262]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[261]) );
  DFF \sreg_reg[262]  ( .D(o[263]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[262]) );
  DFF \sreg_reg[263]  ( .D(o[264]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[263]) );
  DFF \sreg_reg[264]  ( .D(o[265]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[264]) );
  DFF \sreg_reg[265]  ( .D(o[266]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[265]) );
  DFF \sreg_reg[266]  ( .D(o[267]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[266]) );
  DFF \sreg_reg[267]  ( .D(o[268]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[267]) );
  DFF \sreg_reg[268]  ( .D(o[269]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[268]) );
  DFF \sreg_reg[269]  ( .D(o[270]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[269]) );
  DFF \sreg_reg[270]  ( .D(o[271]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[270]) );
  DFF \sreg_reg[271]  ( .D(o[272]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[271]) );
  DFF \sreg_reg[272]  ( .D(o[273]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[272]) );
  DFF \sreg_reg[273]  ( .D(o[274]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[273]) );
  DFF \sreg_reg[274]  ( .D(o[275]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[274]) );
  DFF \sreg_reg[275]  ( .D(o[276]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[275]) );
  DFF \sreg_reg[276]  ( .D(o[277]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[276]) );
  DFF \sreg_reg[277]  ( .D(o[278]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[277]) );
  DFF \sreg_reg[278]  ( .D(o[279]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[278]) );
  DFF \sreg_reg[279]  ( .D(o[280]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[279]) );
  DFF \sreg_reg[280]  ( .D(o[281]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[280]) );
  DFF \sreg_reg[281]  ( .D(o[282]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[281]) );
  DFF \sreg_reg[282]  ( .D(o[283]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[282]) );
  DFF \sreg_reg[283]  ( .D(o[284]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[283]) );
  DFF \sreg_reg[284]  ( .D(o[285]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[284]) );
  DFF \sreg_reg[285]  ( .D(o[286]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[285]) );
  DFF \sreg_reg[286]  ( .D(o[287]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[286]) );
  DFF \sreg_reg[287]  ( .D(o[288]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[287]) );
  DFF \sreg_reg[288]  ( .D(o[289]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[288]) );
  DFF \sreg_reg[289]  ( .D(o[290]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[289]) );
  DFF \sreg_reg[290]  ( .D(o[291]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[290]) );
  DFF \sreg_reg[291]  ( .D(o[292]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[291]) );
  DFF \sreg_reg[292]  ( .D(o[293]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[292]) );
  DFF \sreg_reg[293]  ( .D(o[294]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[293]) );
  DFF \sreg_reg[294]  ( .D(o[295]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[294]) );
  DFF \sreg_reg[295]  ( .D(o[296]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[295]) );
  DFF \sreg_reg[296]  ( .D(o[297]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[296]) );
  DFF \sreg_reg[297]  ( .D(o[298]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[297]) );
  DFF \sreg_reg[298]  ( .D(o[299]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[298]) );
  DFF \sreg_reg[299]  ( .D(o[300]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[299]) );
  DFF \sreg_reg[300]  ( .D(o[301]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[300]) );
  DFF \sreg_reg[301]  ( .D(o[302]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[301]) );
  DFF \sreg_reg[302]  ( .D(o[303]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[302]) );
  DFF \sreg_reg[303]  ( .D(o[304]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[303]) );
  DFF \sreg_reg[304]  ( .D(o[305]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[304]) );
  DFF \sreg_reg[305]  ( .D(o[306]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[305]) );
  DFF \sreg_reg[306]  ( .D(o[307]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[306]) );
  DFF \sreg_reg[307]  ( .D(o[308]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[307]) );
  DFF \sreg_reg[308]  ( .D(o[309]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[308]) );
  DFF \sreg_reg[309]  ( .D(o[310]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[309]) );
  DFF \sreg_reg[310]  ( .D(o[311]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[310]) );
  DFF \sreg_reg[311]  ( .D(o[312]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[311]) );
  DFF \sreg_reg[312]  ( .D(o[313]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[312]) );
  DFF \sreg_reg[313]  ( .D(o[314]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[313]) );
  DFF \sreg_reg[314]  ( .D(o[315]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[314]) );
  DFF \sreg_reg[315]  ( .D(o[316]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[315]) );
  DFF \sreg_reg[316]  ( .D(o[317]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[316]) );
  DFF \sreg_reg[317]  ( .D(o[318]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[317]) );
  DFF \sreg_reg[318]  ( .D(o[319]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[318]) );
  DFF \sreg_reg[319]  ( .D(o[320]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[319]) );
  DFF \sreg_reg[320]  ( .D(o[321]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[320]) );
  DFF \sreg_reg[321]  ( .D(o[322]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[321]) );
  DFF \sreg_reg[322]  ( .D(o[323]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[322]) );
  DFF \sreg_reg[323]  ( .D(o[324]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[323]) );
  DFF \sreg_reg[324]  ( .D(o[325]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[324]) );
  DFF \sreg_reg[325]  ( .D(o[326]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[325]) );
  DFF \sreg_reg[326]  ( .D(o[327]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[326]) );
  DFF \sreg_reg[327]  ( .D(o[328]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[327]) );
  DFF \sreg_reg[328]  ( .D(o[329]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[328]) );
  DFF \sreg_reg[329]  ( .D(o[330]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[329]) );
  DFF \sreg_reg[330]  ( .D(o[331]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[330]) );
  DFF \sreg_reg[331]  ( .D(o[332]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[331]) );
  DFF \sreg_reg[332]  ( .D(o[333]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[332]) );
  DFF \sreg_reg[333]  ( .D(o[334]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[333]) );
  DFF \sreg_reg[334]  ( .D(o[335]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[334]) );
  DFF \sreg_reg[335]  ( .D(o[336]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[335]) );
  DFF \sreg_reg[336]  ( .D(o[337]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[336]) );
  DFF \sreg_reg[337]  ( .D(o[338]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[337]) );
  DFF \sreg_reg[338]  ( .D(o[339]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[338]) );
  DFF \sreg_reg[339]  ( .D(o[340]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[339]) );
  DFF \sreg_reg[340]  ( .D(o[341]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[340]) );
  DFF \sreg_reg[341]  ( .D(o[342]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[341]) );
  DFF \sreg_reg[342]  ( .D(o[343]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[342]) );
  DFF \sreg_reg[343]  ( .D(o[344]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[343]) );
  DFF \sreg_reg[344]  ( .D(o[345]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[344]) );
  DFF \sreg_reg[345]  ( .D(o[346]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[345]) );
  DFF \sreg_reg[346]  ( .D(o[347]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[346]) );
  DFF \sreg_reg[347]  ( .D(o[348]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[347]) );
  DFF \sreg_reg[348]  ( .D(o[349]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[348]) );
  DFF \sreg_reg[349]  ( .D(o[350]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[349]) );
  DFF \sreg_reg[350]  ( .D(o[351]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[350]) );
  DFF \sreg_reg[351]  ( .D(o[352]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[351]) );
  DFF \sreg_reg[352]  ( .D(o[353]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[352]) );
  DFF \sreg_reg[353]  ( .D(o[354]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[353]) );
  DFF \sreg_reg[354]  ( .D(o[355]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[354]) );
  DFF \sreg_reg[355]  ( .D(o[356]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[355]) );
  DFF \sreg_reg[356]  ( .D(o[357]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[356]) );
  DFF \sreg_reg[357]  ( .D(o[358]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[357]) );
  DFF \sreg_reg[358]  ( .D(o[359]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[358]) );
  DFF \sreg_reg[359]  ( .D(o[360]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[359]) );
  DFF \sreg_reg[360]  ( .D(o[361]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[360]) );
  DFF \sreg_reg[361]  ( .D(o[362]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[361]) );
  DFF \sreg_reg[362]  ( .D(o[363]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[362]) );
  DFF \sreg_reg[363]  ( .D(o[364]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[363]) );
  DFF \sreg_reg[364]  ( .D(o[365]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[364]) );
  DFF \sreg_reg[365]  ( .D(o[366]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[365]) );
  DFF \sreg_reg[366]  ( .D(o[367]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[366]) );
  DFF \sreg_reg[367]  ( .D(o[368]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[367]) );
  DFF \sreg_reg[368]  ( .D(o[369]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[368]) );
  DFF \sreg_reg[369]  ( .D(o[370]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[369]) );
  DFF \sreg_reg[370]  ( .D(o[371]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[370]) );
  DFF \sreg_reg[371]  ( .D(o[372]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[371]) );
  DFF \sreg_reg[372]  ( .D(o[373]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[372]) );
  DFF \sreg_reg[373]  ( .D(o[374]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[373]) );
  DFF \sreg_reg[374]  ( .D(o[375]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[374]) );
  DFF \sreg_reg[375]  ( .D(o[376]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[375]) );
  DFF \sreg_reg[376]  ( .D(o[377]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[376]) );
  DFF \sreg_reg[377]  ( .D(o[378]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[377]) );
  DFF \sreg_reg[378]  ( .D(o[379]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[378]) );
  DFF \sreg_reg[379]  ( .D(o[380]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[379]) );
  DFF \sreg_reg[380]  ( .D(o[381]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[380]) );
  DFF \sreg_reg[381]  ( .D(o[382]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[381]) );
  DFF \sreg_reg[382]  ( .D(o[383]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[382]) );
  DFF \sreg_reg[383]  ( .D(o[384]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[383]) );
  DFF \sreg_reg[384]  ( .D(o[385]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[384]) );
  DFF \sreg_reg[385]  ( .D(o[386]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[385]) );
  DFF \sreg_reg[386]  ( .D(o[387]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[386]) );
  DFF \sreg_reg[387]  ( .D(o[388]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[387]) );
  DFF \sreg_reg[388]  ( .D(o[389]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[388]) );
  DFF \sreg_reg[389]  ( .D(o[390]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[389]) );
  DFF \sreg_reg[390]  ( .D(o[391]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[390]) );
  DFF \sreg_reg[391]  ( .D(o[392]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[391]) );
  DFF \sreg_reg[392]  ( .D(o[393]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[392]) );
  DFF \sreg_reg[393]  ( .D(o[394]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[393]) );
  DFF \sreg_reg[394]  ( .D(o[395]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[394]) );
  DFF \sreg_reg[395]  ( .D(o[396]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[395]) );
  DFF \sreg_reg[396]  ( .D(o[397]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[396]) );
  DFF \sreg_reg[397]  ( .D(o[398]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[397]) );
  DFF \sreg_reg[398]  ( .D(o[399]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[398]) );
  DFF \sreg_reg[399]  ( .D(o[400]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[399]) );
  DFF \sreg_reg[400]  ( .D(o[401]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[400]) );
  DFF \sreg_reg[401]  ( .D(o[402]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[401]) );
  DFF \sreg_reg[402]  ( .D(o[403]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[402]) );
  DFF \sreg_reg[403]  ( .D(o[404]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[403]) );
  DFF \sreg_reg[404]  ( .D(o[405]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[404]) );
  DFF \sreg_reg[405]  ( .D(o[406]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[405]) );
  DFF \sreg_reg[406]  ( .D(o[407]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[406]) );
  DFF \sreg_reg[407]  ( .D(o[408]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[407]) );
  DFF \sreg_reg[408]  ( .D(o[409]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[408]) );
  DFF \sreg_reg[409]  ( .D(o[410]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[409]) );
  DFF \sreg_reg[410]  ( .D(o[411]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[410]) );
  DFF \sreg_reg[411]  ( .D(o[412]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[411]) );
  DFF \sreg_reg[412]  ( .D(o[413]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[412]) );
  DFF \sreg_reg[413]  ( .D(o[414]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[413]) );
  DFF \sreg_reg[414]  ( .D(o[415]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[414]) );
  DFF \sreg_reg[415]  ( .D(o[416]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[415]) );
  DFF \sreg_reg[416]  ( .D(o[417]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[416]) );
  DFF \sreg_reg[417]  ( .D(o[418]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[417]) );
  DFF \sreg_reg[418]  ( .D(o[419]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[418]) );
  DFF \sreg_reg[419]  ( .D(o[420]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[419]) );
  DFF \sreg_reg[420]  ( .D(o[421]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[420]) );
  DFF \sreg_reg[421]  ( .D(o[422]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[421]) );
  DFF \sreg_reg[422]  ( .D(o[423]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[422]) );
  DFF \sreg_reg[423]  ( .D(o[424]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[423]) );
  DFF \sreg_reg[424]  ( .D(o[425]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[424]) );
  DFF \sreg_reg[425]  ( .D(o[426]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[425]) );
  DFF \sreg_reg[426]  ( .D(o[427]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[426]) );
  DFF \sreg_reg[427]  ( .D(o[428]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[427]) );
  DFF \sreg_reg[428]  ( .D(o[429]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[428]) );
  DFF \sreg_reg[429]  ( .D(o[430]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[429]) );
  DFF \sreg_reg[430]  ( .D(o[431]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[430]) );
  DFF \sreg_reg[431]  ( .D(o[432]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[431]) );
  DFF \sreg_reg[432]  ( .D(o[433]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[432]) );
  DFF \sreg_reg[433]  ( .D(o[434]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[433]) );
  DFF \sreg_reg[434]  ( .D(o[435]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[434]) );
  DFF \sreg_reg[435]  ( .D(o[436]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[435]) );
  DFF \sreg_reg[436]  ( .D(o[437]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[436]) );
  DFF \sreg_reg[437]  ( .D(o[438]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[437]) );
  DFF \sreg_reg[438]  ( .D(o[439]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[438]) );
  DFF \sreg_reg[439]  ( .D(o[440]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[439]) );
  DFF \sreg_reg[440]  ( .D(o[441]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[440]) );
  DFF \sreg_reg[441]  ( .D(o[442]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[441]) );
  DFF \sreg_reg[442]  ( .D(o[443]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[442]) );
  DFF \sreg_reg[443]  ( .D(o[444]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[443]) );
  DFF \sreg_reg[444]  ( .D(o[445]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[444]) );
  DFF \sreg_reg[445]  ( .D(o[446]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[445]) );
  DFF \sreg_reg[446]  ( .D(o[447]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[446]) );
  DFF \sreg_reg[447]  ( .D(o[448]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[447]) );
  DFF \sreg_reg[448]  ( .D(o[449]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[448]) );
  DFF \sreg_reg[449]  ( .D(o[450]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[449]) );
  DFF \sreg_reg[450]  ( .D(o[451]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[450]) );
  DFF \sreg_reg[451]  ( .D(o[452]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[451]) );
  DFF \sreg_reg[452]  ( .D(o[453]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[452]) );
  DFF \sreg_reg[453]  ( .D(o[454]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[453]) );
  DFF \sreg_reg[454]  ( .D(o[455]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[454]) );
  DFF \sreg_reg[455]  ( .D(o[456]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[455]) );
  DFF \sreg_reg[456]  ( .D(o[457]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[456]) );
  DFF \sreg_reg[457]  ( .D(o[458]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[457]) );
  DFF \sreg_reg[458]  ( .D(o[459]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[458]) );
  DFF \sreg_reg[459]  ( .D(o[460]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[459]) );
  DFF \sreg_reg[460]  ( .D(o[461]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[460]) );
  DFF \sreg_reg[461]  ( .D(o[462]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[461]) );
  DFF \sreg_reg[462]  ( .D(o[463]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[462]) );
  DFF \sreg_reg[463]  ( .D(o[464]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[463]) );
  DFF \sreg_reg[464]  ( .D(o[465]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[464]) );
  DFF \sreg_reg[465]  ( .D(o[466]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[465]) );
  DFF \sreg_reg[466]  ( .D(o[467]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[466]) );
  DFF \sreg_reg[467]  ( .D(o[468]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[467]) );
  DFF \sreg_reg[468]  ( .D(o[469]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[468]) );
  DFF \sreg_reg[469]  ( .D(o[470]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[469]) );
  DFF \sreg_reg[470]  ( .D(o[471]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[470]) );
  DFF \sreg_reg[471]  ( .D(o[472]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[471]) );
  DFF \sreg_reg[472]  ( .D(o[473]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[472]) );
  DFF \sreg_reg[473]  ( .D(o[474]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[473]) );
  DFF \sreg_reg[474]  ( .D(o[475]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[474]) );
  DFF \sreg_reg[475]  ( .D(o[476]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[475]) );
  DFF \sreg_reg[476]  ( .D(o[477]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[476]) );
  DFF \sreg_reg[477]  ( .D(o[478]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[477]) );
  DFF \sreg_reg[478]  ( .D(o[479]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[478]) );
  DFF \sreg_reg[479]  ( .D(o[480]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[479]) );
  DFF \sreg_reg[480]  ( .D(o[481]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[480]) );
  DFF \sreg_reg[481]  ( .D(o[482]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[481]) );
  DFF \sreg_reg[482]  ( .D(o[483]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[482]) );
  DFF \sreg_reg[483]  ( .D(o[484]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[483]) );
  DFF \sreg_reg[484]  ( .D(o[485]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[484]) );
  DFF \sreg_reg[485]  ( .D(o[486]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[485]) );
  DFF \sreg_reg[486]  ( .D(o[487]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[486]) );
  DFF \sreg_reg[487]  ( .D(o[488]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[487]) );
  DFF \sreg_reg[488]  ( .D(o[489]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[488]) );
  DFF \sreg_reg[489]  ( .D(o[490]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[489]) );
  DFF \sreg_reg[490]  ( .D(o[491]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[490]) );
  DFF \sreg_reg[491]  ( .D(o[492]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[491]) );
  DFF \sreg_reg[492]  ( .D(o[493]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[492]) );
  DFF \sreg_reg[493]  ( .D(o[494]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[493]) );
  DFF \sreg_reg[494]  ( .D(o[495]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[494]) );
  DFF \sreg_reg[495]  ( .D(o[496]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[495]) );
  DFF \sreg_reg[496]  ( .D(o[497]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[496]) );
  DFF \sreg_reg[497]  ( .D(o[498]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[497]) );
  DFF \sreg_reg[498]  ( .D(o[499]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[498]) );
  DFF \sreg_reg[499]  ( .D(o[500]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[499]) );
  DFF \sreg_reg[500]  ( .D(o[501]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[500]) );
  DFF \sreg_reg[501]  ( .D(o[502]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[501]) );
  DFF \sreg_reg[502]  ( .D(o[503]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[502]) );
  DFF \sreg_reg[503]  ( .D(o[504]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[503]) );
  DFF \sreg_reg[504]  ( .D(o[505]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[504]) );
  DFF \sreg_reg[505]  ( .D(o[506]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[505]) );
  DFF \sreg_reg[506]  ( .D(o[507]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[506]) );
  DFF \sreg_reg[507]  ( .D(o[508]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[507]) );
  DFF \sreg_reg[508]  ( .D(o[509]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[508]) );
  DFF \sreg_reg[509]  ( .D(o[510]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[509]) );
  DFF \sreg_reg[510]  ( .D(\add_42/carry[511] ), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[510]) );
  FADDER \add_42/U1_256  ( .CIN(sreg[256]), .IN0(n768), .IN1(
        \add_42/carry[256] ), .COUT(\add_42/carry[257] ), .SUM(o[256]) );
  FADDER \add_42/U1_257  ( .CIN(sreg[257]), .IN0(n767), .IN1(
        \add_42/carry[257] ), .COUT(\add_42/carry[258] ), .SUM(o[257]) );
  FADDER \add_42/U1_258  ( .CIN(sreg[258]), .IN0(n766), .IN1(
        \add_42/carry[258] ), .COUT(\add_42/carry[259] ), .SUM(o[258]) );
  FADDER \add_42/U1_259  ( .CIN(sreg[259]), .IN0(n765), .IN1(
        \add_42/carry[259] ), .COUT(\add_42/carry[260] ), .SUM(o[259]) );
  FADDER \add_42/U1_260  ( .CIN(sreg[260]), .IN0(n764), .IN1(
        \add_42/carry[260] ), .COUT(\add_42/carry[261] ), .SUM(o[260]) );
  FADDER \add_42/U1_261  ( .CIN(sreg[261]), .IN0(n763), .IN1(
        \add_42/carry[261] ), .COUT(\add_42/carry[262] ), .SUM(o[261]) );
  FADDER \add_42/U1_262  ( .CIN(sreg[262]), .IN0(n762), .IN1(
        \add_42/carry[262] ), .COUT(\add_42/carry[263] ), .SUM(o[262]) );
  FADDER \add_42/U1_263  ( .CIN(sreg[263]), .IN0(n761), .IN1(
        \add_42/carry[263] ), .COUT(\add_42/carry[264] ), .SUM(o[263]) );
  FADDER \add_42/U1_264  ( .CIN(sreg[264]), .IN0(n760), .IN1(
        \add_42/carry[264] ), .COUT(\add_42/carry[265] ), .SUM(o[264]) );
  FADDER \add_42/U1_265  ( .CIN(sreg[265]), .IN0(n759), .IN1(
        \add_42/carry[265] ), .COUT(\add_42/carry[266] ), .SUM(o[265]) );
  FADDER \add_42/U1_266  ( .CIN(sreg[266]), .IN0(n758), .IN1(
        \add_42/carry[266] ), .COUT(\add_42/carry[267] ), .SUM(o[266]) );
  FADDER \add_42/U1_267  ( .CIN(sreg[267]), .IN0(n757), .IN1(
        \add_42/carry[267] ), .COUT(\add_42/carry[268] ), .SUM(o[267]) );
  FADDER \add_42/U1_268  ( .CIN(sreg[268]), .IN0(n756), .IN1(
        \add_42/carry[268] ), .COUT(\add_42/carry[269] ), .SUM(o[268]) );
  FADDER \add_42/U1_269  ( .CIN(sreg[269]), .IN0(n755), .IN1(
        \add_42/carry[269] ), .COUT(\add_42/carry[270] ), .SUM(o[269]) );
  FADDER \add_42/U1_270  ( .CIN(sreg[270]), .IN0(n754), .IN1(
        \add_42/carry[270] ), .COUT(\add_42/carry[271] ), .SUM(o[270]) );
  FADDER \add_42/U1_271  ( .CIN(sreg[271]), .IN0(n753), .IN1(
        \add_42/carry[271] ), .COUT(\add_42/carry[272] ), .SUM(o[271]) );
  FADDER \add_42/U1_272  ( .CIN(sreg[272]), .IN0(n752), .IN1(
        \add_42/carry[272] ), .COUT(\add_42/carry[273] ), .SUM(o[272]) );
  FADDER \add_42/U1_273  ( .CIN(sreg[273]), .IN0(n751), .IN1(
        \add_42/carry[273] ), .COUT(\add_42/carry[274] ), .SUM(o[273]) );
  FADDER \add_42/U1_274  ( .CIN(sreg[274]), .IN0(n750), .IN1(
        \add_42/carry[274] ), .COUT(\add_42/carry[275] ), .SUM(o[274]) );
  FADDER \add_42/U1_275  ( .CIN(sreg[275]), .IN0(n749), .IN1(
        \add_42/carry[275] ), .COUT(\add_42/carry[276] ), .SUM(o[275]) );
  FADDER \add_42/U1_276  ( .CIN(sreg[276]), .IN0(n748), .IN1(
        \add_42/carry[276] ), .COUT(\add_42/carry[277] ), .SUM(o[276]) );
  FADDER \add_42/U1_277  ( .CIN(sreg[277]), .IN0(n747), .IN1(
        \add_42/carry[277] ), .COUT(\add_42/carry[278] ), .SUM(o[277]) );
  FADDER \add_42/U1_278  ( .CIN(sreg[278]), .IN0(n746), .IN1(
        \add_42/carry[278] ), .COUT(\add_42/carry[279] ), .SUM(o[278]) );
  FADDER \add_42/U1_279  ( .CIN(sreg[279]), .IN0(n745), .IN1(
        \add_42/carry[279] ), .COUT(\add_42/carry[280] ), .SUM(o[279]) );
  FADDER \add_42/U1_280  ( .CIN(sreg[280]), .IN0(n744), .IN1(
        \add_42/carry[280] ), .COUT(\add_42/carry[281] ), .SUM(o[280]) );
  FADDER \add_42/U1_281  ( .CIN(sreg[281]), .IN0(n743), .IN1(
        \add_42/carry[281] ), .COUT(\add_42/carry[282] ), .SUM(o[281]) );
  FADDER \add_42/U1_282  ( .CIN(sreg[282]), .IN0(n742), .IN1(
        \add_42/carry[282] ), .COUT(\add_42/carry[283] ), .SUM(o[282]) );
  FADDER \add_42/U1_283  ( .CIN(sreg[283]), .IN0(n741), .IN1(
        \add_42/carry[283] ), .COUT(\add_42/carry[284] ), .SUM(o[283]) );
  FADDER \add_42/U1_284  ( .CIN(sreg[284]), .IN0(n740), .IN1(
        \add_42/carry[284] ), .COUT(\add_42/carry[285] ), .SUM(o[284]) );
  FADDER \add_42/U1_285  ( .CIN(sreg[285]), .IN0(n739), .IN1(
        \add_42/carry[285] ), .COUT(\add_42/carry[286] ), .SUM(o[285]) );
  FADDER \add_42/U1_286  ( .CIN(sreg[286]), .IN0(n738), .IN1(
        \add_42/carry[286] ), .COUT(\add_42/carry[287] ), .SUM(o[286]) );
  FADDER \add_42/U1_287  ( .CIN(sreg[287]), .IN0(n737), .IN1(
        \add_42/carry[287] ), .COUT(\add_42/carry[288] ), .SUM(o[287]) );
  FADDER \add_42/U1_288  ( .CIN(sreg[288]), .IN0(n736), .IN1(
        \add_42/carry[288] ), .COUT(\add_42/carry[289] ), .SUM(o[288]) );
  FADDER \add_42/U1_289  ( .CIN(sreg[289]), .IN0(n735), .IN1(
        \add_42/carry[289] ), .COUT(\add_42/carry[290] ), .SUM(o[289]) );
  FADDER \add_42/U1_290  ( .CIN(sreg[290]), .IN0(n734), .IN1(
        \add_42/carry[290] ), .COUT(\add_42/carry[291] ), .SUM(o[290]) );
  FADDER \add_42/U1_291  ( .CIN(sreg[291]), .IN0(n733), .IN1(
        \add_42/carry[291] ), .COUT(\add_42/carry[292] ), .SUM(o[291]) );
  FADDER \add_42/U1_292  ( .CIN(sreg[292]), .IN0(n732), .IN1(
        \add_42/carry[292] ), .COUT(\add_42/carry[293] ), .SUM(o[292]) );
  FADDER \add_42/U1_293  ( .CIN(sreg[293]), .IN0(n731), .IN1(
        \add_42/carry[293] ), .COUT(\add_42/carry[294] ), .SUM(o[293]) );
  FADDER \add_42/U1_294  ( .CIN(sreg[294]), .IN0(n730), .IN1(
        \add_42/carry[294] ), .COUT(\add_42/carry[295] ), .SUM(o[294]) );
  FADDER \add_42/U1_295  ( .CIN(sreg[295]), .IN0(n729), .IN1(
        \add_42/carry[295] ), .COUT(\add_42/carry[296] ), .SUM(o[295]) );
  FADDER \add_42/U1_296  ( .CIN(sreg[296]), .IN0(n728), .IN1(
        \add_42/carry[296] ), .COUT(\add_42/carry[297] ), .SUM(o[296]) );
  FADDER \add_42/U1_297  ( .CIN(sreg[297]), .IN0(n727), .IN1(
        \add_42/carry[297] ), .COUT(\add_42/carry[298] ), .SUM(o[297]) );
  FADDER \add_42/U1_298  ( .CIN(sreg[298]), .IN0(n726), .IN1(
        \add_42/carry[298] ), .COUT(\add_42/carry[299] ), .SUM(o[298]) );
  FADDER \add_42/U1_299  ( .CIN(sreg[299]), .IN0(n725), .IN1(
        \add_42/carry[299] ), .COUT(\add_42/carry[300] ), .SUM(o[299]) );
  FADDER \add_42/U1_300  ( .CIN(sreg[300]), .IN0(n724), .IN1(
        \add_42/carry[300] ), .COUT(\add_42/carry[301] ), .SUM(o[300]) );
  FADDER \add_42/U1_301  ( .CIN(sreg[301]), .IN0(n723), .IN1(
        \add_42/carry[301] ), .COUT(\add_42/carry[302] ), .SUM(o[301]) );
  FADDER \add_42/U1_302  ( .CIN(sreg[302]), .IN0(n722), .IN1(
        \add_42/carry[302] ), .COUT(\add_42/carry[303] ), .SUM(o[302]) );
  FADDER \add_42/U1_303  ( .CIN(sreg[303]), .IN0(n721), .IN1(
        \add_42/carry[303] ), .COUT(\add_42/carry[304] ), .SUM(o[303]) );
  FADDER \add_42/U1_304  ( .CIN(sreg[304]), .IN0(n720), .IN1(
        \add_42/carry[304] ), .COUT(\add_42/carry[305] ), .SUM(o[304]) );
  FADDER \add_42/U1_305  ( .CIN(sreg[305]), .IN0(n719), .IN1(
        \add_42/carry[305] ), .COUT(\add_42/carry[306] ), .SUM(o[305]) );
  FADDER \add_42/U1_306  ( .CIN(sreg[306]), .IN0(n718), .IN1(
        \add_42/carry[306] ), .COUT(\add_42/carry[307] ), .SUM(o[306]) );
  FADDER \add_42/U1_307  ( .CIN(sreg[307]), .IN0(n717), .IN1(
        \add_42/carry[307] ), .COUT(\add_42/carry[308] ), .SUM(o[307]) );
  FADDER \add_42/U1_308  ( .CIN(sreg[308]), .IN0(n716), .IN1(
        \add_42/carry[308] ), .COUT(\add_42/carry[309] ), .SUM(o[308]) );
  FADDER \add_42/U1_309  ( .CIN(sreg[309]), .IN0(n715), .IN1(
        \add_42/carry[309] ), .COUT(\add_42/carry[310] ), .SUM(o[309]) );
  FADDER \add_42/U1_310  ( .CIN(sreg[310]), .IN0(n714), .IN1(
        \add_42/carry[310] ), .COUT(\add_42/carry[311] ), .SUM(o[310]) );
  FADDER \add_42/U1_311  ( .CIN(sreg[311]), .IN0(n713), .IN1(
        \add_42/carry[311] ), .COUT(\add_42/carry[312] ), .SUM(o[311]) );
  FADDER \add_42/U1_312  ( .CIN(sreg[312]), .IN0(n712), .IN1(
        \add_42/carry[312] ), .COUT(\add_42/carry[313] ), .SUM(o[312]) );
  FADDER \add_42/U1_313  ( .CIN(sreg[313]), .IN0(n711), .IN1(
        \add_42/carry[313] ), .COUT(\add_42/carry[314] ), .SUM(o[313]) );
  FADDER \add_42/U1_314  ( .CIN(sreg[314]), .IN0(n710), .IN1(
        \add_42/carry[314] ), .COUT(\add_42/carry[315] ), .SUM(o[314]) );
  FADDER \add_42/U1_315  ( .CIN(sreg[315]), .IN0(n709), .IN1(
        \add_42/carry[315] ), .COUT(\add_42/carry[316] ), .SUM(o[315]) );
  FADDER \add_42/U1_316  ( .CIN(sreg[316]), .IN0(n708), .IN1(
        \add_42/carry[316] ), .COUT(\add_42/carry[317] ), .SUM(o[316]) );
  FADDER \add_42/U1_317  ( .CIN(sreg[317]), .IN0(n707), .IN1(
        \add_42/carry[317] ), .COUT(\add_42/carry[318] ), .SUM(o[317]) );
  FADDER \add_42/U1_318  ( .CIN(sreg[318]), .IN0(n706), .IN1(
        \add_42/carry[318] ), .COUT(\add_42/carry[319] ), .SUM(o[318]) );
  FADDER \add_42/U1_319  ( .CIN(sreg[319]), .IN0(n705), .IN1(
        \add_42/carry[319] ), .COUT(\add_42/carry[320] ), .SUM(o[319]) );
  FADDER \add_42/U1_320  ( .CIN(sreg[320]), .IN0(n704), .IN1(
        \add_42/carry[320] ), .COUT(\add_42/carry[321] ), .SUM(o[320]) );
  FADDER \add_42/U1_321  ( .CIN(sreg[321]), .IN0(n703), .IN1(
        \add_42/carry[321] ), .COUT(\add_42/carry[322] ), .SUM(o[321]) );
  FADDER \add_42/U1_322  ( .CIN(sreg[322]), .IN0(n702), .IN1(
        \add_42/carry[322] ), .COUT(\add_42/carry[323] ), .SUM(o[322]) );
  FADDER \add_42/U1_323  ( .CIN(sreg[323]), .IN0(n701), .IN1(
        \add_42/carry[323] ), .COUT(\add_42/carry[324] ), .SUM(o[323]) );
  FADDER \add_42/U1_324  ( .CIN(sreg[324]), .IN0(n700), .IN1(
        \add_42/carry[324] ), .COUT(\add_42/carry[325] ), .SUM(o[324]) );
  FADDER \add_42/U1_325  ( .CIN(sreg[325]), .IN0(n699), .IN1(
        \add_42/carry[325] ), .COUT(\add_42/carry[326] ), .SUM(o[325]) );
  FADDER \add_42/U1_326  ( .CIN(sreg[326]), .IN0(n698), .IN1(
        \add_42/carry[326] ), .COUT(\add_42/carry[327] ), .SUM(o[326]) );
  FADDER \add_42/U1_327  ( .CIN(sreg[327]), .IN0(n697), .IN1(
        \add_42/carry[327] ), .COUT(\add_42/carry[328] ), .SUM(o[327]) );
  FADDER \add_42/U1_328  ( .CIN(sreg[328]), .IN0(n696), .IN1(
        \add_42/carry[328] ), .COUT(\add_42/carry[329] ), .SUM(o[328]) );
  FADDER \add_42/U1_329  ( .CIN(sreg[329]), .IN0(n695), .IN1(
        \add_42/carry[329] ), .COUT(\add_42/carry[330] ), .SUM(o[329]) );
  FADDER \add_42/U1_330  ( .CIN(sreg[330]), .IN0(n694), .IN1(
        \add_42/carry[330] ), .COUT(\add_42/carry[331] ), .SUM(o[330]) );
  FADDER \add_42/U1_331  ( .CIN(sreg[331]), .IN0(n693), .IN1(
        \add_42/carry[331] ), .COUT(\add_42/carry[332] ), .SUM(o[331]) );
  FADDER \add_42/U1_332  ( .CIN(sreg[332]), .IN0(n692), .IN1(
        \add_42/carry[332] ), .COUT(\add_42/carry[333] ), .SUM(o[332]) );
  FADDER \add_42/U1_333  ( .CIN(sreg[333]), .IN0(n691), .IN1(
        \add_42/carry[333] ), .COUT(\add_42/carry[334] ), .SUM(o[333]) );
  FADDER \add_42/U1_334  ( .CIN(sreg[334]), .IN0(n690), .IN1(
        \add_42/carry[334] ), .COUT(\add_42/carry[335] ), .SUM(o[334]) );
  FADDER \add_42/U1_335  ( .CIN(sreg[335]), .IN0(n689), .IN1(
        \add_42/carry[335] ), .COUT(\add_42/carry[336] ), .SUM(o[335]) );
  FADDER \add_42/U1_336  ( .CIN(sreg[336]), .IN0(n688), .IN1(
        \add_42/carry[336] ), .COUT(\add_42/carry[337] ), .SUM(o[336]) );
  FADDER \add_42/U1_337  ( .CIN(sreg[337]), .IN0(n687), .IN1(
        \add_42/carry[337] ), .COUT(\add_42/carry[338] ), .SUM(o[337]) );
  FADDER \add_42/U1_338  ( .CIN(sreg[338]), .IN0(n686), .IN1(
        \add_42/carry[338] ), .COUT(\add_42/carry[339] ), .SUM(o[338]) );
  FADDER \add_42/U1_339  ( .CIN(sreg[339]), .IN0(n685), .IN1(
        \add_42/carry[339] ), .COUT(\add_42/carry[340] ), .SUM(o[339]) );
  FADDER \add_42/U1_340  ( .CIN(sreg[340]), .IN0(n684), .IN1(
        \add_42/carry[340] ), .COUT(\add_42/carry[341] ), .SUM(o[340]) );
  FADDER \add_42/U1_341  ( .CIN(sreg[341]), .IN0(n683), .IN1(
        \add_42/carry[341] ), .COUT(\add_42/carry[342] ), .SUM(o[341]) );
  FADDER \add_42/U1_342  ( .CIN(sreg[342]), .IN0(n682), .IN1(
        \add_42/carry[342] ), .COUT(\add_42/carry[343] ), .SUM(o[342]) );
  FADDER \add_42/U1_343  ( .CIN(sreg[343]), .IN0(n681), .IN1(
        \add_42/carry[343] ), .COUT(\add_42/carry[344] ), .SUM(o[343]) );
  FADDER \add_42/U1_344  ( .CIN(sreg[344]), .IN0(n680), .IN1(
        \add_42/carry[344] ), .COUT(\add_42/carry[345] ), .SUM(o[344]) );
  FADDER \add_42/U1_345  ( .CIN(sreg[345]), .IN0(n679), .IN1(
        \add_42/carry[345] ), .COUT(\add_42/carry[346] ), .SUM(o[345]) );
  FADDER \add_42/U1_346  ( .CIN(sreg[346]), .IN0(n678), .IN1(
        \add_42/carry[346] ), .COUT(\add_42/carry[347] ), .SUM(o[346]) );
  FADDER \add_42/U1_347  ( .CIN(sreg[347]), .IN0(n677), .IN1(
        \add_42/carry[347] ), .COUT(\add_42/carry[348] ), .SUM(o[347]) );
  FADDER \add_42/U1_348  ( .CIN(sreg[348]), .IN0(n676), .IN1(
        \add_42/carry[348] ), .COUT(\add_42/carry[349] ), .SUM(o[348]) );
  FADDER \add_42/U1_349  ( .CIN(sreg[349]), .IN0(n675), .IN1(
        \add_42/carry[349] ), .COUT(\add_42/carry[350] ), .SUM(o[349]) );
  FADDER \add_42/U1_350  ( .CIN(sreg[350]), .IN0(n674), .IN1(
        \add_42/carry[350] ), .COUT(\add_42/carry[351] ), .SUM(o[350]) );
  FADDER \add_42/U1_351  ( .CIN(sreg[351]), .IN0(n673), .IN1(
        \add_42/carry[351] ), .COUT(\add_42/carry[352] ), .SUM(o[351]) );
  FADDER \add_42/U1_352  ( .CIN(sreg[352]), .IN0(n672), .IN1(
        \add_42/carry[352] ), .COUT(\add_42/carry[353] ), .SUM(o[352]) );
  FADDER \add_42/U1_353  ( .CIN(sreg[353]), .IN0(n671), .IN1(
        \add_42/carry[353] ), .COUT(\add_42/carry[354] ), .SUM(o[353]) );
  FADDER \add_42/U1_354  ( .CIN(sreg[354]), .IN0(n670), .IN1(
        \add_42/carry[354] ), .COUT(\add_42/carry[355] ), .SUM(o[354]) );
  FADDER \add_42/U1_355  ( .CIN(sreg[355]), .IN0(n669), .IN1(
        \add_42/carry[355] ), .COUT(\add_42/carry[356] ), .SUM(o[355]) );
  FADDER \add_42/U1_356  ( .CIN(sreg[356]), .IN0(n668), .IN1(
        \add_42/carry[356] ), .COUT(\add_42/carry[357] ), .SUM(o[356]) );
  FADDER \add_42/U1_357  ( .CIN(sreg[357]), .IN0(n667), .IN1(
        \add_42/carry[357] ), .COUT(\add_42/carry[358] ), .SUM(o[357]) );
  FADDER \add_42/U1_358  ( .CIN(sreg[358]), .IN0(n666), .IN1(
        \add_42/carry[358] ), .COUT(\add_42/carry[359] ), .SUM(o[358]) );
  FADDER \add_42/U1_359  ( .CIN(sreg[359]), .IN0(n665), .IN1(
        \add_42/carry[359] ), .COUT(\add_42/carry[360] ), .SUM(o[359]) );
  FADDER \add_42/U1_360  ( .CIN(sreg[360]), .IN0(n664), .IN1(
        \add_42/carry[360] ), .COUT(\add_42/carry[361] ), .SUM(o[360]) );
  FADDER \add_42/U1_361  ( .CIN(sreg[361]), .IN0(n663), .IN1(
        \add_42/carry[361] ), .COUT(\add_42/carry[362] ), .SUM(o[361]) );
  FADDER \add_42/U1_362  ( .CIN(sreg[362]), .IN0(n662), .IN1(
        \add_42/carry[362] ), .COUT(\add_42/carry[363] ), .SUM(o[362]) );
  FADDER \add_42/U1_363  ( .CIN(sreg[363]), .IN0(n661), .IN1(
        \add_42/carry[363] ), .COUT(\add_42/carry[364] ), .SUM(o[363]) );
  FADDER \add_42/U1_364  ( .CIN(sreg[364]), .IN0(n660), .IN1(
        \add_42/carry[364] ), .COUT(\add_42/carry[365] ), .SUM(o[364]) );
  FADDER \add_42/U1_365  ( .CIN(sreg[365]), .IN0(n659), .IN1(
        \add_42/carry[365] ), .COUT(\add_42/carry[366] ), .SUM(o[365]) );
  FADDER \add_42/U1_366  ( .CIN(sreg[366]), .IN0(n658), .IN1(
        \add_42/carry[366] ), .COUT(\add_42/carry[367] ), .SUM(o[366]) );
  FADDER \add_42/U1_367  ( .CIN(sreg[367]), .IN0(n657), .IN1(
        \add_42/carry[367] ), .COUT(\add_42/carry[368] ), .SUM(o[367]) );
  FADDER \add_42/U1_368  ( .CIN(sreg[368]), .IN0(n656), .IN1(
        \add_42/carry[368] ), .COUT(\add_42/carry[369] ), .SUM(o[368]) );
  FADDER \add_42/U1_369  ( .CIN(sreg[369]), .IN0(n655), .IN1(
        \add_42/carry[369] ), .COUT(\add_42/carry[370] ), .SUM(o[369]) );
  FADDER \add_42/U1_370  ( .CIN(sreg[370]), .IN0(n654), .IN1(
        \add_42/carry[370] ), .COUT(\add_42/carry[371] ), .SUM(o[370]) );
  FADDER \add_42/U1_371  ( .CIN(sreg[371]), .IN0(n653), .IN1(
        \add_42/carry[371] ), .COUT(\add_42/carry[372] ), .SUM(o[371]) );
  FADDER \add_42/U1_372  ( .CIN(sreg[372]), .IN0(n652), .IN1(
        \add_42/carry[372] ), .COUT(\add_42/carry[373] ), .SUM(o[372]) );
  FADDER \add_42/U1_373  ( .CIN(sreg[373]), .IN0(n651), .IN1(
        \add_42/carry[373] ), .COUT(\add_42/carry[374] ), .SUM(o[373]) );
  FADDER \add_42/U1_374  ( .CIN(sreg[374]), .IN0(n650), .IN1(
        \add_42/carry[374] ), .COUT(\add_42/carry[375] ), .SUM(o[374]) );
  FADDER \add_42/U1_375  ( .CIN(sreg[375]), .IN0(n649), .IN1(
        \add_42/carry[375] ), .COUT(\add_42/carry[376] ), .SUM(o[375]) );
  FADDER \add_42/U1_376  ( .CIN(sreg[376]), .IN0(n648), .IN1(
        \add_42/carry[376] ), .COUT(\add_42/carry[377] ), .SUM(o[376]) );
  FADDER \add_42/U1_377  ( .CIN(sreg[377]), .IN0(n647), .IN1(
        \add_42/carry[377] ), .COUT(\add_42/carry[378] ), .SUM(o[377]) );
  FADDER \add_42/U1_378  ( .CIN(sreg[378]), .IN0(n646), .IN1(
        \add_42/carry[378] ), .COUT(\add_42/carry[379] ), .SUM(o[378]) );
  FADDER \add_42/U1_379  ( .CIN(sreg[379]), .IN0(n645), .IN1(
        \add_42/carry[379] ), .COUT(\add_42/carry[380] ), .SUM(o[379]) );
  FADDER \add_42/U1_380  ( .CIN(sreg[380]), .IN0(n644), .IN1(
        \add_42/carry[380] ), .COUT(\add_42/carry[381] ), .SUM(o[380]) );
  FADDER \add_42/U1_381  ( .CIN(sreg[381]), .IN0(n643), .IN1(
        \add_42/carry[381] ), .COUT(\add_42/carry[382] ), .SUM(o[381]) );
  FADDER \add_42/U1_382  ( .CIN(sreg[382]), .IN0(n642), .IN1(
        \add_42/carry[382] ), .COUT(\add_42/carry[383] ), .SUM(o[382]) );
  FADDER \add_42/U1_383  ( .CIN(sreg[383]), .IN0(n641), .IN1(
        \add_42/carry[383] ), .COUT(\add_42/carry[384] ), .SUM(o[383]) );
  FADDER \add_42/U1_384  ( .CIN(sreg[384]), .IN0(n640), .IN1(
        \add_42/carry[384] ), .COUT(\add_42/carry[385] ), .SUM(o[384]) );
  FADDER \add_42/U1_385  ( .CIN(sreg[385]), .IN0(n639), .IN1(
        \add_42/carry[385] ), .COUT(\add_42/carry[386] ), .SUM(o[385]) );
  FADDER \add_42/U1_386  ( .CIN(sreg[386]), .IN0(n638), .IN1(
        \add_42/carry[386] ), .COUT(\add_42/carry[387] ), .SUM(o[386]) );
  FADDER \add_42/U1_387  ( .CIN(sreg[387]), .IN0(n637), .IN1(
        \add_42/carry[387] ), .COUT(\add_42/carry[388] ), .SUM(o[387]) );
  FADDER \add_42/U1_388  ( .CIN(sreg[388]), .IN0(n636), .IN1(
        \add_42/carry[388] ), .COUT(\add_42/carry[389] ), .SUM(o[388]) );
  FADDER \add_42/U1_389  ( .CIN(sreg[389]), .IN0(n635), .IN1(
        \add_42/carry[389] ), .COUT(\add_42/carry[390] ), .SUM(o[389]) );
  FADDER \add_42/U1_390  ( .CIN(sreg[390]), .IN0(n634), .IN1(
        \add_42/carry[390] ), .COUT(\add_42/carry[391] ), .SUM(o[390]) );
  FADDER \add_42/U1_391  ( .CIN(sreg[391]), .IN0(n633), .IN1(
        \add_42/carry[391] ), .COUT(\add_42/carry[392] ), .SUM(o[391]) );
  FADDER \add_42/U1_392  ( .CIN(sreg[392]), .IN0(n632), .IN1(
        \add_42/carry[392] ), .COUT(\add_42/carry[393] ), .SUM(o[392]) );
  FADDER \add_42/U1_393  ( .CIN(sreg[393]), .IN0(n631), .IN1(
        \add_42/carry[393] ), .COUT(\add_42/carry[394] ), .SUM(o[393]) );
  FADDER \add_42/U1_394  ( .CIN(sreg[394]), .IN0(n630), .IN1(
        \add_42/carry[394] ), .COUT(\add_42/carry[395] ), .SUM(o[394]) );
  FADDER \add_42/U1_395  ( .CIN(sreg[395]), .IN0(n629), .IN1(
        \add_42/carry[395] ), .COUT(\add_42/carry[396] ), .SUM(o[395]) );
  FADDER \add_42/U1_396  ( .CIN(sreg[396]), .IN0(n628), .IN1(
        \add_42/carry[396] ), .COUT(\add_42/carry[397] ), .SUM(o[396]) );
  FADDER \add_42/U1_397  ( .CIN(sreg[397]), .IN0(n627), .IN1(
        \add_42/carry[397] ), .COUT(\add_42/carry[398] ), .SUM(o[397]) );
  FADDER \add_42/U1_398  ( .CIN(sreg[398]), .IN0(n626), .IN1(
        \add_42/carry[398] ), .COUT(\add_42/carry[399] ), .SUM(o[398]) );
  FADDER \add_42/U1_399  ( .CIN(sreg[399]), .IN0(n625), .IN1(
        \add_42/carry[399] ), .COUT(\add_42/carry[400] ), .SUM(o[399]) );
  FADDER \add_42/U1_400  ( .CIN(sreg[400]), .IN0(n624), .IN1(
        \add_42/carry[400] ), .COUT(\add_42/carry[401] ), .SUM(o[400]) );
  FADDER \add_42/U1_401  ( .CIN(sreg[401]), .IN0(n623), .IN1(
        \add_42/carry[401] ), .COUT(\add_42/carry[402] ), .SUM(o[401]) );
  FADDER \add_42/U1_402  ( .CIN(sreg[402]), .IN0(n622), .IN1(
        \add_42/carry[402] ), .COUT(\add_42/carry[403] ), .SUM(o[402]) );
  FADDER \add_42/U1_403  ( .CIN(sreg[403]), .IN0(n621), .IN1(
        \add_42/carry[403] ), .COUT(\add_42/carry[404] ), .SUM(o[403]) );
  FADDER \add_42/U1_404  ( .CIN(sreg[404]), .IN0(n620), .IN1(
        \add_42/carry[404] ), .COUT(\add_42/carry[405] ), .SUM(o[404]) );
  FADDER \add_42/U1_405  ( .CIN(sreg[405]), .IN0(n619), .IN1(
        \add_42/carry[405] ), .COUT(\add_42/carry[406] ), .SUM(o[405]) );
  FADDER \add_42/U1_406  ( .CIN(sreg[406]), .IN0(n618), .IN1(
        \add_42/carry[406] ), .COUT(\add_42/carry[407] ), .SUM(o[406]) );
  FADDER \add_42/U1_407  ( .CIN(sreg[407]), .IN0(n617), .IN1(
        \add_42/carry[407] ), .COUT(\add_42/carry[408] ), .SUM(o[407]) );
  FADDER \add_42/U1_408  ( .CIN(sreg[408]), .IN0(n616), .IN1(
        \add_42/carry[408] ), .COUT(\add_42/carry[409] ), .SUM(o[408]) );
  FADDER \add_42/U1_409  ( .CIN(sreg[409]), .IN0(n615), .IN1(
        \add_42/carry[409] ), .COUT(\add_42/carry[410] ), .SUM(o[409]) );
  FADDER \add_42/U1_410  ( .CIN(sreg[410]), .IN0(n614), .IN1(
        \add_42/carry[410] ), .COUT(\add_42/carry[411] ), .SUM(o[410]) );
  FADDER \add_42/U1_411  ( .CIN(sreg[411]), .IN0(n613), .IN1(
        \add_42/carry[411] ), .COUT(\add_42/carry[412] ), .SUM(o[411]) );
  FADDER \add_42/U1_412  ( .CIN(sreg[412]), .IN0(n612), .IN1(
        \add_42/carry[412] ), .COUT(\add_42/carry[413] ), .SUM(o[412]) );
  FADDER \add_42/U1_413  ( .CIN(sreg[413]), .IN0(n611), .IN1(
        \add_42/carry[413] ), .COUT(\add_42/carry[414] ), .SUM(o[413]) );
  FADDER \add_42/U1_414  ( .CIN(sreg[414]), .IN0(n610), .IN1(
        \add_42/carry[414] ), .COUT(\add_42/carry[415] ), .SUM(o[414]) );
  FADDER \add_42/U1_415  ( .CIN(sreg[415]), .IN0(n609), .IN1(
        \add_42/carry[415] ), .COUT(\add_42/carry[416] ), .SUM(o[415]) );
  FADDER \add_42/U1_416  ( .CIN(sreg[416]), .IN0(n608), .IN1(
        \add_42/carry[416] ), .COUT(\add_42/carry[417] ), .SUM(o[416]) );
  FADDER \add_42/U1_417  ( .CIN(sreg[417]), .IN0(n607), .IN1(
        \add_42/carry[417] ), .COUT(\add_42/carry[418] ), .SUM(o[417]) );
  FADDER \add_42/U1_418  ( .CIN(sreg[418]), .IN0(n606), .IN1(
        \add_42/carry[418] ), .COUT(\add_42/carry[419] ), .SUM(o[418]) );
  FADDER \add_42/U1_419  ( .CIN(sreg[419]), .IN0(n605), .IN1(
        \add_42/carry[419] ), .COUT(\add_42/carry[420] ), .SUM(o[419]) );
  FADDER \add_42/U1_420  ( .CIN(sreg[420]), .IN0(n604), .IN1(
        \add_42/carry[420] ), .COUT(\add_42/carry[421] ), .SUM(o[420]) );
  FADDER \add_42/U1_421  ( .CIN(sreg[421]), .IN0(n603), .IN1(
        \add_42/carry[421] ), .COUT(\add_42/carry[422] ), .SUM(o[421]) );
  FADDER \add_42/U1_422  ( .CIN(sreg[422]), .IN0(n602), .IN1(
        \add_42/carry[422] ), .COUT(\add_42/carry[423] ), .SUM(o[422]) );
  FADDER \add_42/U1_423  ( .CIN(sreg[423]), .IN0(n601), .IN1(
        \add_42/carry[423] ), .COUT(\add_42/carry[424] ), .SUM(o[423]) );
  FADDER \add_42/U1_424  ( .CIN(sreg[424]), .IN0(n600), .IN1(
        \add_42/carry[424] ), .COUT(\add_42/carry[425] ), .SUM(o[424]) );
  FADDER \add_42/U1_425  ( .CIN(sreg[425]), .IN0(n599), .IN1(
        \add_42/carry[425] ), .COUT(\add_42/carry[426] ), .SUM(o[425]) );
  FADDER \add_42/U1_426  ( .CIN(sreg[426]), .IN0(n598), .IN1(
        \add_42/carry[426] ), .COUT(\add_42/carry[427] ), .SUM(o[426]) );
  FADDER \add_42/U1_427  ( .CIN(sreg[427]), .IN0(n597), .IN1(
        \add_42/carry[427] ), .COUT(\add_42/carry[428] ), .SUM(o[427]) );
  FADDER \add_42/U1_428  ( .CIN(sreg[428]), .IN0(n596), .IN1(
        \add_42/carry[428] ), .COUT(\add_42/carry[429] ), .SUM(o[428]) );
  FADDER \add_42/U1_429  ( .CIN(sreg[429]), .IN0(n595), .IN1(
        \add_42/carry[429] ), .COUT(\add_42/carry[430] ), .SUM(o[429]) );
  FADDER \add_42/U1_430  ( .CIN(sreg[430]), .IN0(n594), .IN1(
        \add_42/carry[430] ), .COUT(\add_42/carry[431] ), .SUM(o[430]) );
  FADDER \add_42/U1_431  ( .CIN(sreg[431]), .IN0(n593), .IN1(
        \add_42/carry[431] ), .COUT(\add_42/carry[432] ), .SUM(o[431]) );
  FADDER \add_42/U1_432  ( .CIN(sreg[432]), .IN0(n592), .IN1(
        \add_42/carry[432] ), .COUT(\add_42/carry[433] ), .SUM(o[432]) );
  FADDER \add_42/U1_433  ( .CIN(sreg[433]), .IN0(n591), .IN1(
        \add_42/carry[433] ), .COUT(\add_42/carry[434] ), .SUM(o[433]) );
  FADDER \add_42/U1_434  ( .CIN(sreg[434]), .IN0(n590), .IN1(
        \add_42/carry[434] ), .COUT(\add_42/carry[435] ), .SUM(o[434]) );
  FADDER \add_42/U1_435  ( .CIN(sreg[435]), .IN0(n589), .IN1(
        \add_42/carry[435] ), .COUT(\add_42/carry[436] ), .SUM(o[435]) );
  FADDER \add_42/U1_436  ( .CIN(sreg[436]), .IN0(n588), .IN1(
        \add_42/carry[436] ), .COUT(\add_42/carry[437] ), .SUM(o[436]) );
  FADDER \add_42/U1_437  ( .CIN(sreg[437]), .IN0(n587), .IN1(
        \add_42/carry[437] ), .COUT(\add_42/carry[438] ), .SUM(o[437]) );
  FADDER \add_42/U1_438  ( .CIN(sreg[438]), .IN0(n586), .IN1(
        \add_42/carry[438] ), .COUT(\add_42/carry[439] ), .SUM(o[438]) );
  FADDER \add_42/U1_439  ( .CIN(sreg[439]), .IN0(n585), .IN1(
        \add_42/carry[439] ), .COUT(\add_42/carry[440] ), .SUM(o[439]) );
  FADDER \add_42/U1_440  ( .CIN(sreg[440]), .IN0(n584), .IN1(
        \add_42/carry[440] ), .COUT(\add_42/carry[441] ), .SUM(o[440]) );
  FADDER \add_42/U1_441  ( .CIN(sreg[441]), .IN0(n583), .IN1(
        \add_42/carry[441] ), .COUT(\add_42/carry[442] ), .SUM(o[441]) );
  FADDER \add_42/U1_442  ( .CIN(sreg[442]), .IN0(n582), .IN1(
        \add_42/carry[442] ), .COUT(\add_42/carry[443] ), .SUM(o[442]) );
  FADDER \add_42/U1_443  ( .CIN(sreg[443]), .IN0(n581), .IN1(
        \add_42/carry[443] ), .COUT(\add_42/carry[444] ), .SUM(o[443]) );
  FADDER \add_42/U1_444  ( .CIN(sreg[444]), .IN0(n580), .IN1(
        \add_42/carry[444] ), .COUT(\add_42/carry[445] ), .SUM(o[444]) );
  FADDER \add_42/U1_445  ( .CIN(sreg[445]), .IN0(n579), .IN1(
        \add_42/carry[445] ), .COUT(\add_42/carry[446] ), .SUM(o[445]) );
  FADDER \add_42/U1_446  ( .CIN(sreg[446]), .IN0(n578), .IN1(
        \add_42/carry[446] ), .COUT(\add_42/carry[447] ), .SUM(o[446]) );
  FADDER \add_42/U1_447  ( .CIN(sreg[447]), .IN0(n577), .IN1(
        \add_42/carry[447] ), .COUT(\add_42/carry[448] ), .SUM(o[447]) );
  FADDER \add_42/U1_448  ( .CIN(sreg[448]), .IN0(n576), .IN1(
        \add_42/carry[448] ), .COUT(\add_42/carry[449] ), .SUM(o[448]) );
  FADDER \add_42/U1_449  ( .CIN(sreg[449]), .IN0(n575), .IN1(
        \add_42/carry[449] ), .COUT(\add_42/carry[450] ), .SUM(o[449]) );
  FADDER \add_42/U1_450  ( .CIN(sreg[450]), .IN0(n574), .IN1(
        \add_42/carry[450] ), .COUT(\add_42/carry[451] ), .SUM(o[450]) );
  FADDER \add_42/U1_451  ( .CIN(sreg[451]), .IN0(n573), .IN1(
        \add_42/carry[451] ), .COUT(\add_42/carry[452] ), .SUM(o[451]) );
  FADDER \add_42/U1_452  ( .CIN(sreg[452]), .IN0(n572), .IN1(
        \add_42/carry[452] ), .COUT(\add_42/carry[453] ), .SUM(o[452]) );
  FADDER \add_42/U1_453  ( .CIN(sreg[453]), .IN0(n571), .IN1(
        \add_42/carry[453] ), .COUT(\add_42/carry[454] ), .SUM(o[453]) );
  FADDER \add_42/U1_454  ( .CIN(sreg[454]), .IN0(n570), .IN1(
        \add_42/carry[454] ), .COUT(\add_42/carry[455] ), .SUM(o[454]) );
  FADDER \add_42/U1_455  ( .CIN(sreg[455]), .IN0(n569), .IN1(
        \add_42/carry[455] ), .COUT(\add_42/carry[456] ), .SUM(o[455]) );
  FADDER \add_42/U1_456  ( .CIN(sreg[456]), .IN0(n568), .IN1(
        \add_42/carry[456] ), .COUT(\add_42/carry[457] ), .SUM(o[456]) );
  FADDER \add_42/U1_457  ( .CIN(sreg[457]), .IN0(n567), .IN1(
        \add_42/carry[457] ), .COUT(\add_42/carry[458] ), .SUM(o[457]) );
  FADDER \add_42/U1_458  ( .CIN(sreg[458]), .IN0(n566), .IN1(
        \add_42/carry[458] ), .COUT(\add_42/carry[459] ), .SUM(o[458]) );
  FADDER \add_42/U1_459  ( .CIN(sreg[459]), .IN0(n565), .IN1(
        \add_42/carry[459] ), .COUT(\add_42/carry[460] ), .SUM(o[459]) );
  FADDER \add_42/U1_460  ( .CIN(sreg[460]), .IN0(n564), .IN1(
        \add_42/carry[460] ), .COUT(\add_42/carry[461] ), .SUM(o[460]) );
  FADDER \add_42/U1_461  ( .CIN(sreg[461]), .IN0(n563), .IN1(
        \add_42/carry[461] ), .COUT(\add_42/carry[462] ), .SUM(o[461]) );
  FADDER \add_42/U1_462  ( .CIN(sreg[462]), .IN0(n562), .IN1(
        \add_42/carry[462] ), .COUT(\add_42/carry[463] ), .SUM(o[462]) );
  FADDER \add_42/U1_463  ( .CIN(sreg[463]), .IN0(n561), .IN1(
        \add_42/carry[463] ), .COUT(\add_42/carry[464] ), .SUM(o[463]) );
  FADDER \add_42/U1_464  ( .CIN(sreg[464]), .IN0(n560), .IN1(
        \add_42/carry[464] ), .COUT(\add_42/carry[465] ), .SUM(o[464]) );
  FADDER \add_42/U1_465  ( .CIN(sreg[465]), .IN0(n559), .IN1(
        \add_42/carry[465] ), .COUT(\add_42/carry[466] ), .SUM(o[465]) );
  FADDER \add_42/U1_466  ( .CIN(sreg[466]), .IN0(n558), .IN1(
        \add_42/carry[466] ), .COUT(\add_42/carry[467] ), .SUM(o[466]) );
  FADDER \add_42/U1_467  ( .CIN(sreg[467]), .IN0(n557), .IN1(
        \add_42/carry[467] ), .COUT(\add_42/carry[468] ), .SUM(o[467]) );
  FADDER \add_42/U1_468  ( .CIN(sreg[468]), .IN0(n556), .IN1(
        \add_42/carry[468] ), .COUT(\add_42/carry[469] ), .SUM(o[468]) );
  FADDER \add_42/U1_469  ( .CIN(sreg[469]), .IN0(n555), .IN1(
        \add_42/carry[469] ), .COUT(\add_42/carry[470] ), .SUM(o[469]) );
  FADDER \add_42/U1_470  ( .CIN(sreg[470]), .IN0(n554), .IN1(
        \add_42/carry[470] ), .COUT(\add_42/carry[471] ), .SUM(o[470]) );
  FADDER \add_42/U1_471  ( .CIN(sreg[471]), .IN0(n553), .IN1(
        \add_42/carry[471] ), .COUT(\add_42/carry[472] ), .SUM(o[471]) );
  FADDER \add_42/U1_472  ( .CIN(sreg[472]), .IN0(n552), .IN1(
        \add_42/carry[472] ), .COUT(\add_42/carry[473] ), .SUM(o[472]) );
  FADDER \add_42/U1_473  ( .CIN(sreg[473]), .IN0(n551), .IN1(
        \add_42/carry[473] ), .COUT(\add_42/carry[474] ), .SUM(o[473]) );
  FADDER \add_42/U1_474  ( .CIN(sreg[474]), .IN0(n550), .IN1(
        \add_42/carry[474] ), .COUT(\add_42/carry[475] ), .SUM(o[474]) );
  FADDER \add_42/U1_475  ( .CIN(sreg[475]), .IN0(n549), .IN1(
        \add_42/carry[475] ), .COUT(\add_42/carry[476] ), .SUM(o[475]) );
  FADDER \add_42/U1_476  ( .CIN(sreg[476]), .IN0(n548), .IN1(
        \add_42/carry[476] ), .COUT(\add_42/carry[477] ), .SUM(o[476]) );
  FADDER \add_42/U1_477  ( .CIN(sreg[477]), .IN0(n547), .IN1(
        \add_42/carry[477] ), .COUT(\add_42/carry[478] ), .SUM(o[477]) );
  FADDER \add_42/U1_478  ( .CIN(sreg[478]), .IN0(n546), .IN1(
        \add_42/carry[478] ), .COUT(\add_42/carry[479] ), .SUM(o[478]) );
  FADDER \add_42/U1_479  ( .CIN(sreg[479]), .IN0(n545), .IN1(
        \add_42/carry[479] ), .COUT(\add_42/carry[480] ), .SUM(o[479]) );
  FADDER \add_42/U1_480  ( .CIN(sreg[480]), .IN0(n544), .IN1(
        \add_42/carry[480] ), .COUT(\add_42/carry[481] ), .SUM(o[480]) );
  FADDER \add_42/U1_481  ( .CIN(sreg[481]), .IN0(n543), .IN1(
        \add_42/carry[481] ), .COUT(\add_42/carry[482] ), .SUM(o[481]) );
  FADDER \add_42/U1_482  ( .CIN(sreg[482]), .IN0(n542), .IN1(
        \add_42/carry[482] ), .COUT(\add_42/carry[483] ), .SUM(o[482]) );
  FADDER \add_42/U1_483  ( .CIN(sreg[483]), .IN0(n541), .IN1(
        \add_42/carry[483] ), .COUT(\add_42/carry[484] ), .SUM(o[483]) );
  FADDER \add_42/U1_484  ( .CIN(sreg[484]), .IN0(n540), .IN1(
        \add_42/carry[484] ), .COUT(\add_42/carry[485] ), .SUM(o[484]) );
  FADDER \add_42/U1_485  ( .CIN(sreg[485]), .IN0(n539), .IN1(
        \add_42/carry[485] ), .COUT(\add_42/carry[486] ), .SUM(o[485]) );
  FADDER \add_42/U1_486  ( .CIN(sreg[486]), .IN0(n538), .IN1(
        \add_42/carry[486] ), .COUT(\add_42/carry[487] ), .SUM(o[486]) );
  FADDER \add_42/U1_487  ( .CIN(sreg[487]), .IN0(n537), .IN1(
        \add_42/carry[487] ), .COUT(\add_42/carry[488] ), .SUM(o[487]) );
  FADDER \add_42/U1_488  ( .CIN(sreg[488]), .IN0(n536), .IN1(
        \add_42/carry[488] ), .COUT(\add_42/carry[489] ), .SUM(o[488]) );
  FADDER \add_42/U1_489  ( .CIN(sreg[489]), .IN0(n535), .IN1(
        \add_42/carry[489] ), .COUT(\add_42/carry[490] ), .SUM(o[489]) );
  FADDER \add_42/U1_490  ( .CIN(sreg[490]), .IN0(n534), .IN1(
        \add_42/carry[490] ), .COUT(\add_42/carry[491] ), .SUM(o[490]) );
  FADDER \add_42/U1_491  ( .CIN(sreg[491]), .IN0(n533), .IN1(
        \add_42/carry[491] ), .COUT(\add_42/carry[492] ), .SUM(o[491]) );
  FADDER \add_42/U1_492  ( .CIN(sreg[492]), .IN0(n532), .IN1(
        \add_42/carry[492] ), .COUT(\add_42/carry[493] ), .SUM(o[492]) );
  FADDER \add_42/U1_493  ( .CIN(sreg[493]), .IN0(n531), .IN1(
        \add_42/carry[493] ), .COUT(\add_42/carry[494] ), .SUM(o[493]) );
  FADDER \add_42/U1_494  ( .CIN(sreg[494]), .IN0(n530), .IN1(
        \add_42/carry[494] ), .COUT(\add_42/carry[495] ), .SUM(o[494]) );
  FADDER \add_42/U1_495  ( .CIN(sreg[495]), .IN0(n529), .IN1(
        \add_42/carry[495] ), .COUT(\add_42/carry[496] ), .SUM(o[495]) );
  FADDER \add_42/U1_496  ( .CIN(sreg[496]), .IN0(n528), .IN1(
        \add_42/carry[496] ), .COUT(\add_42/carry[497] ), .SUM(o[496]) );
  FADDER \add_42/U1_497  ( .CIN(sreg[497]), .IN0(n527), .IN1(
        \add_42/carry[497] ), .COUT(\add_42/carry[498] ), .SUM(o[497]) );
  FADDER \add_42/U1_498  ( .CIN(sreg[498]), .IN0(n526), .IN1(
        \add_42/carry[498] ), .COUT(\add_42/carry[499] ), .SUM(o[498]) );
  FADDER \add_42/U1_499  ( .CIN(sreg[499]), .IN0(n525), .IN1(
        \add_42/carry[499] ), .COUT(\add_42/carry[500] ), .SUM(o[499]) );
  FADDER \add_42/U1_500  ( .CIN(sreg[500]), .IN0(n524), .IN1(
        \add_42/carry[500] ), .COUT(\add_42/carry[501] ), .SUM(o[500]) );
  FADDER \add_42/U1_501  ( .CIN(sreg[501]), .IN0(n523), .IN1(
        \add_42/carry[501] ), .COUT(\add_42/carry[502] ), .SUM(o[501]) );
  FADDER \add_42/U1_502  ( .CIN(sreg[502]), .IN0(n522), .IN1(
        \add_42/carry[502] ), .COUT(\add_42/carry[503] ), .SUM(o[502]) );
  FADDER \add_42/U1_503  ( .CIN(sreg[503]), .IN0(n521), .IN1(
        \add_42/carry[503] ), .COUT(\add_42/carry[504] ), .SUM(o[503]) );
  FADDER \add_42/U1_504  ( .CIN(sreg[504]), .IN0(n520), .IN1(
        \add_42/carry[504] ), .COUT(\add_42/carry[505] ), .SUM(o[504]) );
  FADDER \add_42/U1_505  ( .CIN(sreg[505]), .IN0(n519), .IN1(
        \add_42/carry[505] ), .COUT(\add_42/carry[506] ), .SUM(o[505]) );
  FADDER \add_42/U1_506  ( .CIN(sreg[506]), .IN0(n518), .IN1(
        \add_42/carry[506] ), .COUT(\add_42/carry[507] ), .SUM(o[506]) );
  FADDER \add_42/U1_507  ( .CIN(sreg[507]), .IN0(n517), .IN1(
        \add_42/carry[507] ), .COUT(\add_42/carry[508] ), .SUM(o[507]) );
  FADDER \add_42/U1_508  ( .CIN(sreg[508]), .IN0(n516), .IN1(
        \add_42/carry[508] ), .COUT(\add_42/carry[509] ), .SUM(o[508]) );
  FADDER \add_42/U1_509  ( .CIN(sreg[509]), .IN0(n515), .IN1(
        \add_42/carry[509] ), .COUT(\add_42/carry[510] ), .SUM(o[509]) );
  FADDER \add_42/U1_510  ( .CIN(sreg[510]), .IN0(n514), .IN1(
        \add_42/carry[510] ), .COUT(\add_42/carry[511] ), .SUM(o[510]) );
  AND U517 ( .A(sreg[255]), .B(n769), .Z(\add_42/carry[256] ) );
  XOR U518 ( .A(n769), .B(sreg[255]), .Z(o[255]) );
  AND U519 ( .A(g_input[255]), .B(e_input[0]), .Z(n514) );
  AND U520 ( .A(g_input[254]), .B(e_input[0]), .Z(n515) );
  AND U521 ( .A(g_input[253]), .B(e_input[0]), .Z(n516) );
  AND U522 ( .A(g_input[252]), .B(e_input[0]), .Z(n517) );
  AND U523 ( .A(g_input[251]), .B(e_input[0]), .Z(n518) );
  AND U524 ( .A(g_input[250]), .B(e_input[0]), .Z(n519) );
  AND U525 ( .A(g_input[249]), .B(e_input[0]), .Z(n520) );
  AND U526 ( .A(g_input[248]), .B(e_input[0]), .Z(n521) );
  AND U527 ( .A(g_input[247]), .B(e_input[0]), .Z(n522) );
  AND U528 ( .A(g_input[246]), .B(e_input[0]), .Z(n523) );
  AND U529 ( .A(g_input[245]), .B(e_input[0]), .Z(n524) );
  AND U530 ( .A(g_input[244]), .B(e_input[0]), .Z(n525) );
  AND U531 ( .A(g_input[243]), .B(e_input[0]), .Z(n526) );
  AND U532 ( .A(g_input[242]), .B(e_input[0]), .Z(n527) );
  AND U533 ( .A(g_input[241]), .B(e_input[0]), .Z(n528) );
  AND U534 ( .A(g_input[240]), .B(e_input[0]), .Z(n529) );
  AND U535 ( .A(g_input[239]), .B(e_input[0]), .Z(n530) );
  AND U536 ( .A(g_input[238]), .B(e_input[0]), .Z(n531) );
  AND U537 ( .A(g_input[237]), .B(e_input[0]), .Z(n532) );
  AND U538 ( .A(g_input[236]), .B(e_input[0]), .Z(n533) );
  AND U539 ( .A(g_input[235]), .B(e_input[0]), .Z(n534) );
  AND U540 ( .A(g_input[234]), .B(e_input[0]), .Z(n535) );
  AND U541 ( .A(g_input[233]), .B(e_input[0]), .Z(n536) );
  AND U542 ( .A(g_input[232]), .B(e_input[0]), .Z(n537) );
  AND U543 ( .A(g_input[231]), .B(e_input[0]), .Z(n538) );
  AND U544 ( .A(g_input[230]), .B(e_input[0]), .Z(n539) );
  AND U545 ( .A(g_input[229]), .B(e_input[0]), .Z(n540) );
  AND U546 ( .A(g_input[228]), .B(e_input[0]), .Z(n541) );
  AND U547 ( .A(g_input[227]), .B(e_input[0]), .Z(n542) );
  AND U548 ( .A(g_input[226]), .B(e_input[0]), .Z(n543) );
  AND U549 ( .A(g_input[225]), .B(e_input[0]), .Z(n544) );
  AND U550 ( .A(g_input[224]), .B(e_input[0]), .Z(n545) );
  AND U551 ( .A(g_input[223]), .B(e_input[0]), .Z(n546) );
  AND U552 ( .A(g_input[222]), .B(e_input[0]), .Z(n547) );
  AND U553 ( .A(g_input[221]), .B(e_input[0]), .Z(n548) );
  AND U554 ( .A(g_input[220]), .B(e_input[0]), .Z(n549) );
  AND U555 ( .A(g_input[219]), .B(e_input[0]), .Z(n550) );
  AND U556 ( .A(g_input[218]), .B(e_input[0]), .Z(n551) );
  AND U557 ( .A(g_input[217]), .B(e_input[0]), .Z(n552) );
  AND U558 ( .A(g_input[216]), .B(e_input[0]), .Z(n553) );
  AND U559 ( .A(g_input[215]), .B(e_input[0]), .Z(n554) );
  AND U560 ( .A(g_input[214]), .B(e_input[0]), .Z(n555) );
  AND U561 ( .A(g_input[213]), .B(e_input[0]), .Z(n556) );
  AND U562 ( .A(g_input[212]), .B(e_input[0]), .Z(n557) );
  AND U563 ( .A(g_input[211]), .B(e_input[0]), .Z(n558) );
  AND U564 ( .A(g_input[210]), .B(e_input[0]), .Z(n559) );
  AND U565 ( .A(g_input[209]), .B(e_input[0]), .Z(n560) );
  AND U566 ( .A(g_input[208]), .B(e_input[0]), .Z(n561) );
  AND U567 ( .A(g_input[207]), .B(e_input[0]), .Z(n562) );
  AND U568 ( .A(g_input[206]), .B(e_input[0]), .Z(n563) );
  AND U569 ( .A(g_input[205]), .B(e_input[0]), .Z(n564) );
  AND U570 ( .A(g_input[204]), .B(e_input[0]), .Z(n565) );
  AND U571 ( .A(g_input[203]), .B(e_input[0]), .Z(n566) );
  AND U572 ( .A(g_input[202]), .B(e_input[0]), .Z(n567) );
  AND U573 ( .A(g_input[201]), .B(e_input[0]), .Z(n568) );
  AND U574 ( .A(g_input[200]), .B(e_input[0]), .Z(n569) );
  AND U575 ( .A(g_input[199]), .B(e_input[0]), .Z(n570) );
  AND U576 ( .A(g_input[198]), .B(e_input[0]), .Z(n571) );
  AND U577 ( .A(g_input[197]), .B(e_input[0]), .Z(n572) );
  AND U578 ( .A(g_input[196]), .B(e_input[0]), .Z(n573) );
  AND U579 ( .A(g_input[195]), .B(e_input[0]), .Z(n574) );
  AND U580 ( .A(g_input[194]), .B(e_input[0]), .Z(n575) );
  AND U581 ( .A(g_input[193]), .B(e_input[0]), .Z(n576) );
  AND U582 ( .A(g_input[192]), .B(e_input[0]), .Z(n577) );
  AND U583 ( .A(g_input[191]), .B(e_input[0]), .Z(n578) );
  AND U584 ( .A(g_input[190]), .B(e_input[0]), .Z(n579) );
  AND U585 ( .A(g_input[189]), .B(e_input[0]), .Z(n580) );
  AND U586 ( .A(g_input[188]), .B(e_input[0]), .Z(n581) );
  AND U587 ( .A(g_input[187]), .B(e_input[0]), .Z(n582) );
  AND U588 ( .A(g_input[186]), .B(e_input[0]), .Z(n583) );
  AND U589 ( .A(g_input[185]), .B(e_input[0]), .Z(n584) );
  AND U590 ( .A(g_input[184]), .B(e_input[0]), .Z(n585) );
  AND U591 ( .A(g_input[183]), .B(e_input[0]), .Z(n586) );
  AND U592 ( .A(g_input[182]), .B(e_input[0]), .Z(n587) );
  AND U593 ( .A(g_input[181]), .B(e_input[0]), .Z(n588) );
  AND U594 ( .A(g_input[180]), .B(e_input[0]), .Z(n589) );
  AND U595 ( .A(g_input[179]), .B(e_input[0]), .Z(n590) );
  AND U596 ( .A(g_input[178]), .B(e_input[0]), .Z(n591) );
  AND U597 ( .A(g_input[177]), .B(e_input[0]), .Z(n592) );
  AND U598 ( .A(g_input[176]), .B(e_input[0]), .Z(n593) );
  AND U599 ( .A(g_input[175]), .B(e_input[0]), .Z(n594) );
  AND U600 ( .A(g_input[174]), .B(e_input[0]), .Z(n595) );
  AND U601 ( .A(g_input[173]), .B(e_input[0]), .Z(n596) );
  AND U602 ( .A(g_input[172]), .B(e_input[0]), .Z(n597) );
  AND U603 ( .A(g_input[171]), .B(e_input[0]), .Z(n598) );
  AND U604 ( .A(g_input[170]), .B(e_input[0]), .Z(n599) );
  AND U605 ( .A(g_input[169]), .B(e_input[0]), .Z(n600) );
  AND U606 ( .A(g_input[168]), .B(e_input[0]), .Z(n601) );
  AND U607 ( .A(g_input[167]), .B(e_input[0]), .Z(n602) );
  AND U608 ( .A(g_input[166]), .B(e_input[0]), .Z(n603) );
  AND U609 ( .A(g_input[165]), .B(e_input[0]), .Z(n604) );
  AND U610 ( .A(g_input[164]), .B(e_input[0]), .Z(n605) );
  AND U611 ( .A(g_input[163]), .B(e_input[0]), .Z(n606) );
  AND U612 ( .A(g_input[162]), .B(e_input[0]), .Z(n607) );
  AND U613 ( .A(g_input[161]), .B(e_input[0]), .Z(n608) );
  AND U614 ( .A(g_input[160]), .B(e_input[0]), .Z(n609) );
  AND U615 ( .A(g_input[159]), .B(e_input[0]), .Z(n610) );
  AND U616 ( .A(g_input[158]), .B(e_input[0]), .Z(n611) );
  AND U617 ( .A(g_input[157]), .B(e_input[0]), .Z(n612) );
  AND U618 ( .A(g_input[156]), .B(e_input[0]), .Z(n613) );
  AND U619 ( .A(g_input[155]), .B(e_input[0]), .Z(n614) );
  AND U620 ( .A(g_input[154]), .B(e_input[0]), .Z(n615) );
  AND U621 ( .A(g_input[153]), .B(e_input[0]), .Z(n616) );
  AND U622 ( .A(g_input[152]), .B(e_input[0]), .Z(n617) );
  AND U623 ( .A(g_input[151]), .B(e_input[0]), .Z(n618) );
  AND U624 ( .A(g_input[150]), .B(e_input[0]), .Z(n619) );
  AND U625 ( .A(g_input[149]), .B(e_input[0]), .Z(n620) );
  AND U626 ( .A(g_input[148]), .B(e_input[0]), .Z(n621) );
  AND U627 ( .A(g_input[147]), .B(e_input[0]), .Z(n622) );
  AND U628 ( .A(g_input[146]), .B(e_input[0]), .Z(n623) );
  AND U629 ( .A(g_input[145]), .B(e_input[0]), .Z(n624) );
  AND U630 ( .A(g_input[144]), .B(e_input[0]), .Z(n625) );
  AND U631 ( .A(g_input[143]), .B(e_input[0]), .Z(n626) );
  AND U632 ( .A(g_input[142]), .B(e_input[0]), .Z(n627) );
  AND U633 ( .A(g_input[141]), .B(e_input[0]), .Z(n628) );
  AND U634 ( .A(g_input[140]), .B(e_input[0]), .Z(n629) );
  AND U635 ( .A(g_input[139]), .B(e_input[0]), .Z(n630) );
  AND U636 ( .A(g_input[138]), .B(e_input[0]), .Z(n631) );
  AND U637 ( .A(g_input[137]), .B(e_input[0]), .Z(n632) );
  AND U638 ( .A(g_input[136]), .B(e_input[0]), .Z(n633) );
  AND U639 ( .A(g_input[135]), .B(e_input[0]), .Z(n634) );
  AND U640 ( .A(g_input[134]), .B(e_input[0]), .Z(n635) );
  AND U641 ( .A(g_input[133]), .B(e_input[0]), .Z(n636) );
  AND U642 ( .A(g_input[132]), .B(e_input[0]), .Z(n637) );
  AND U643 ( .A(g_input[131]), .B(e_input[0]), .Z(n638) );
  AND U644 ( .A(g_input[130]), .B(e_input[0]), .Z(n639) );
  AND U645 ( .A(g_input[129]), .B(e_input[0]), .Z(n640) );
  AND U646 ( .A(g_input[128]), .B(e_input[0]), .Z(n641) );
  AND U647 ( .A(g_input[127]), .B(e_input[0]), .Z(n642) );
  AND U648 ( .A(g_input[126]), .B(e_input[0]), .Z(n643) );
  AND U649 ( .A(g_input[125]), .B(e_input[0]), .Z(n644) );
  AND U650 ( .A(g_input[124]), .B(e_input[0]), .Z(n645) );
  AND U651 ( .A(g_input[123]), .B(e_input[0]), .Z(n646) );
  AND U652 ( .A(g_input[122]), .B(e_input[0]), .Z(n647) );
  AND U653 ( .A(g_input[121]), .B(e_input[0]), .Z(n648) );
  AND U654 ( .A(g_input[120]), .B(e_input[0]), .Z(n649) );
  AND U655 ( .A(g_input[119]), .B(e_input[0]), .Z(n650) );
  AND U656 ( .A(g_input[118]), .B(e_input[0]), .Z(n651) );
  AND U657 ( .A(g_input[117]), .B(e_input[0]), .Z(n652) );
  AND U658 ( .A(g_input[116]), .B(e_input[0]), .Z(n653) );
  AND U659 ( .A(g_input[115]), .B(e_input[0]), .Z(n654) );
  AND U660 ( .A(g_input[114]), .B(e_input[0]), .Z(n655) );
  AND U661 ( .A(g_input[113]), .B(e_input[0]), .Z(n656) );
  AND U662 ( .A(g_input[112]), .B(e_input[0]), .Z(n657) );
  AND U663 ( .A(g_input[111]), .B(e_input[0]), .Z(n658) );
  AND U664 ( .A(g_input[110]), .B(e_input[0]), .Z(n659) );
  AND U665 ( .A(g_input[109]), .B(e_input[0]), .Z(n660) );
  AND U666 ( .A(g_input[108]), .B(e_input[0]), .Z(n661) );
  AND U667 ( .A(g_input[107]), .B(e_input[0]), .Z(n662) );
  AND U668 ( .A(g_input[106]), .B(e_input[0]), .Z(n663) );
  AND U669 ( .A(g_input[105]), .B(e_input[0]), .Z(n664) );
  AND U670 ( .A(g_input[104]), .B(e_input[0]), .Z(n665) );
  AND U671 ( .A(g_input[103]), .B(e_input[0]), .Z(n666) );
  AND U672 ( .A(g_input[102]), .B(e_input[0]), .Z(n667) );
  AND U673 ( .A(g_input[101]), .B(e_input[0]), .Z(n668) );
  AND U674 ( .A(g_input[100]), .B(e_input[0]), .Z(n669) );
  AND U675 ( .A(g_input[99]), .B(e_input[0]), .Z(n670) );
  AND U676 ( .A(g_input[98]), .B(e_input[0]), .Z(n671) );
  AND U677 ( .A(g_input[97]), .B(e_input[0]), .Z(n672) );
  AND U678 ( .A(g_input[96]), .B(e_input[0]), .Z(n673) );
  AND U679 ( .A(g_input[95]), .B(e_input[0]), .Z(n674) );
  AND U680 ( .A(g_input[94]), .B(e_input[0]), .Z(n675) );
  AND U681 ( .A(g_input[93]), .B(e_input[0]), .Z(n676) );
  AND U682 ( .A(g_input[92]), .B(e_input[0]), .Z(n677) );
  AND U683 ( .A(g_input[91]), .B(e_input[0]), .Z(n678) );
  AND U684 ( .A(g_input[90]), .B(e_input[0]), .Z(n679) );
  AND U685 ( .A(g_input[89]), .B(e_input[0]), .Z(n680) );
  AND U686 ( .A(g_input[88]), .B(e_input[0]), .Z(n681) );
  AND U687 ( .A(g_input[87]), .B(e_input[0]), .Z(n682) );
  AND U688 ( .A(g_input[86]), .B(e_input[0]), .Z(n683) );
  AND U689 ( .A(g_input[85]), .B(e_input[0]), .Z(n684) );
  AND U690 ( .A(g_input[84]), .B(e_input[0]), .Z(n685) );
  AND U691 ( .A(g_input[83]), .B(e_input[0]), .Z(n686) );
  AND U692 ( .A(g_input[82]), .B(e_input[0]), .Z(n687) );
  AND U693 ( .A(g_input[81]), .B(e_input[0]), .Z(n688) );
  AND U694 ( .A(g_input[80]), .B(e_input[0]), .Z(n689) );
  AND U695 ( .A(g_input[79]), .B(e_input[0]), .Z(n690) );
  AND U696 ( .A(g_input[78]), .B(e_input[0]), .Z(n691) );
  AND U697 ( .A(g_input[77]), .B(e_input[0]), .Z(n692) );
  AND U698 ( .A(g_input[76]), .B(e_input[0]), .Z(n693) );
  AND U699 ( .A(g_input[75]), .B(e_input[0]), .Z(n694) );
  AND U700 ( .A(g_input[74]), .B(e_input[0]), .Z(n695) );
  AND U701 ( .A(g_input[73]), .B(e_input[0]), .Z(n696) );
  AND U702 ( .A(g_input[72]), .B(e_input[0]), .Z(n697) );
  AND U703 ( .A(g_input[71]), .B(e_input[0]), .Z(n698) );
  AND U704 ( .A(g_input[70]), .B(e_input[0]), .Z(n699) );
  AND U705 ( .A(g_input[69]), .B(e_input[0]), .Z(n700) );
  AND U706 ( .A(g_input[68]), .B(e_input[0]), .Z(n701) );
  AND U707 ( .A(g_input[67]), .B(e_input[0]), .Z(n702) );
  AND U708 ( .A(g_input[66]), .B(e_input[0]), .Z(n703) );
  AND U709 ( .A(g_input[65]), .B(e_input[0]), .Z(n704) );
  AND U710 ( .A(g_input[64]), .B(e_input[0]), .Z(n705) );
  AND U711 ( .A(g_input[63]), .B(e_input[0]), .Z(n706) );
  AND U712 ( .A(g_input[62]), .B(e_input[0]), .Z(n707) );
  AND U713 ( .A(g_input[61]), .B(e_input[0]), .Z(n708) );
  AND U714 ( .A(g_input[60]), .B(e_input[0]), .Z(n709) );
  AND U715 ( .A(g_input[59]), .B(e_input[0]), .Z(n710) );
  AND U716 ( .A(g_input[58]), .B(e_input[0]), .Z(n711) );
  AND U717 ( .A(g_input[57]), .B(e_input[0]), .Z(n712) );
  AND U718 ( .A(g_input[56]), .B(e_input[0]), .Z(n713) );
  AND U719 ( .A(g_input[55]), .B(e_input[0]), .Z(n714) );
  AND U720 ( .A(g_input[54]), .B(e_input[0]), .Z(n715) );
  AND U721 ( .A(g_input[53]), .B(e_input[0]), .Z(n716) );
  AND U722 ( .A(g_input[52]), .B(e_input[0]), .Z(n717) );
  AND U723 ( .A(g_input[51]), .B(e_input[0]), .Z(n718) );
  AND U724 ( .A(g_input[50]), .B(e_input[0]), .Z(n719) );
  AND U725 ( .A(g_input[49]), .B(e_input[0]), .Z(n720) );
  AND U726 ( .A(g_input[48]), .B(e_input[0]), .Z(n721) );
  AND U727 ( .A(g_input[47]), .B(e_input[0]), .Z(n722) );
  AND U728 ( .A(g_input[46]), .B(e_input[0]), .Z(n723) );
  AND U729 ( .A(g_input[45]), .B(e_input[0]), .Z(n724) );
  AND U730 ( .A(g_input[44]), .B(e_input[0]), .Z(n725) );
  AND U731 ( .A(g_input[43]), .B(e_input[0]), .Z(n726) );
  AND U732 ( .A(g_input[42]), .B(e_input[0]), .Z(n727) );
  AND U733 ( .A(g_input[41]), .B(e_input[0]), .Z(n728) );
  AND U734 ( .A(g_input[40]), .B(e_input[0]), .Z(n729) );
  AND U735 ( .A(g_input[39]), .B(e_input[0]), .Z(n730) );
  AND U736 ( .A(g_input[38]), .B(e_input[0]), .Z(n731) );
  AND U737 ( .A(g_input[37]), .B(e_input[0]), .Z(n732) );
  AND U738 ( .A(g_input[36]), .B(e_input[0]), .Z(n733) );
  AND U739 ( .A(g_input[35]), .B(e_input[0]), .Z(n734) );
  AND U740 ( .A(g_input[34]), .B(e_input[0]), .Z(n735) );
  AND U741 ( .A(g_input[33]), .B(e_input[0]), .Z(n736) );
  AND U742 ( .A(g_input[32]), .B(e_input[0]), .Z(n737) );
  AND U743 ( .A(g_input[31]), .B(e_input[0]), .Z(n738) );
  AND U744 ( .A(g_input[30]), .B(e_input[0]), .Z(n739) );
  AND U745 ( .A(g_input[29]), .B(e_input[0]), .Z(n740) );
  AND U746 ( .A(g_input[28]), .B(e_input[0]), .Z(n741) );
  AND U747 ( .A(g_input[27]), .B(e_input[0]), .Z(n742) );
  AND U748 ( .A(g_input[26]), .B(e_input[0]), .Z(n743) );
  AND U749 ( .A(g_input[25]), .B(e_input[0]), .Z(n744) );
  AND U750 ( .A(g_input[24]), .B(e_input[0]), .Z(n745) );
  AND U751 ( .A(g_input[23]), .B(e_input[0]), .Z(n746) );
  AND U752 ( .A(g_input[22]), .B(e_input[0]), .Z(n747) );
  AND U753 ( .A(g_input[21]), .B(e_input[0]), .Z(n748) );
  AND U754 ( .A(g_input[20]), .B(e_input[0]), .Z(n749) );
  AND U755 ( .A(g_input[19]), .B(e_input[0]), .Z(n750) );
  AND U756 ( .A(g_input[18]), .B(e_input[0]), .Z(n751) );
  AND U757 ( .A(g_input[17]), .B(e_input[0]), .Z(n752) );
  AND U758 ( .A(g_input[16]), .B(e_input[0]), .Z(n753) );
  AND U759 ( .A(g_input[15]), .B(e_input[0]), .Z(n754) );
  AND U760 ( .A(g_input[14]), .B(e_input[0]), .Z(n755) );
  AND U761 ( .A(g_input[13]), .B(e_input[0]), .Z(n756) );
  AND U762 ( .A(g_input[12]), .B(e_input[0]), .Z(n757) );
  AND U763 ( .A(g_input[11]), .B(e_input[0]), .Z(n758) );
  AND U764 ( .A(g_input[10]), .B(e_input[0]), .Z(n759) );
  AND U765 ( .A(g_input[9]), .B(e_input[0]), .Z(n760) );
  AND U766 ( .A(g_input[8]), .B(e_input[0]), .Z(n761) );
  AND U767 ( .A(g_input[7]), .B(e_input[0]), .Z(n762) );
  AND U768 ( .A(g_input[6]), .B(e_input[0]), .Z(n763) );
  AND U769 ( .A(g_input[5]), .B(e_input[0]), .Z(n764) );
  AND U770 ( .A(g_input[4]), .B(e_input[0]), .Z(n765) );
  AND U771 ( .A(g_input[3]), .B(e_input[0]), .Z(n766) );
  AND U772 ( .A(g_input[2]), .B(e_input[0]), .Z(n767) );
  AND U773 ( .A(g_input[1]), .B(e_input[0]), .Z(n768) );
  AND U774 ( .A(g_input[0]), .B(e_input[0]), .Z(n769) );
endmodule

