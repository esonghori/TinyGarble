
module compare_N16384_CC16 ( clk, rst, x, y, g );
  input [1023:0] x;
  input [1023:0] y;
  input clk, rst;
  output g;
  wire   ci, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120;

  DFF ci_reg ( .D(g), .CLK(clk), .RST(rst), .I(1'b1), .Q(ci) );
  XOR U1028 ( .A(y[3]), .B(n5107), .Z(n5108) );
  XOR U1029 ( .A(y[7]), .B(n5091), .Z(n5092) );
  XOR U1030 ( .A(y[11]), .B(n5075), .Z(n5076) );
  XOR U1031 ( .A(y[15]), .B(n5059), .Z(n5060) );
  XOR U1032 ( .A(y[19]), .B(n5043), .Z(n5044) );
  XOR U1033 ( .A(y[23]), .B(n5027), .Z(n5028) );
  XOR U1034 ( .A(y[27]), .B(n5011), .Z(n5012) );
  XOR U1035 ( .A(y[31]), .B(n4995), .Z(n4996) );
  XOR U1036 ( .A(y[35]), .B(n4979), .Z(n4980) );
  XOR U1037 ( .A(y[39]), .B(n4963), .Z(n4964) );
  XOR U1038 ( .A(y[43]), .B(n4947), .Z(n4948) );
  XOR U1039 ( .A(y[47]), .B(n4931), .Z(n4932) );
  XOR U1040 ( .A(y[51]), .B(n4915), .Z(n4916) );
  XOR U1041 ( .A(y[55]), .B(n4899), .Z(n4900) );
  XOR U1042 ( .A(y[59]), .B(n4883), .Z(n4884) );
  XOR U1043 ( .A(y[63]), .B(n4867), .Z(n4868) );
  XOR U1044 ( .A(y[67]), .B(n4851), .Z(n4852) );
  XOR U1045 ( .A(y[71]), .B(n4835), .Z(n4836) );
  XOR U1046 ( .A(y[75]), .B(n4819), .Z(n4820) );
  XOR U1047 ( .A(y[79]), .B(n4803), .Z(n4804) );
  XOR U1048 ( .A(y[83]), .B(n4787), .Z(n4788) );
  XOR U1049 ( .A(y[87]), .B(n4771), .Z(n4772) );
  XOR U1050 ( .A(y[91]), .B(n4755), .Z(n4756) );
  XOR U1051 ( .A(y[95]), .B(n4739), .Z(n4740) );
  XOR U1052 ( .A(y[99]), .B(n4723), .Z(n4724) );
  XOR U1053 ( .A(y[103]), .B(n4707), .Z(n4708) );
  XOR U1054 ( .A(y[107]), .B(n4691), .Z(n4692) );
  XOR U1055 ( .A(y[111]), .B(n4675), .Z(n4676) );
  XOR U1056 ( .A(y[115]), .B(n4659), .Z(n4660) );
  XOR U1057 ( .A(y[119]), .B(n4643), .Z(n4644) );
  XOR U1058 ( .A(y[123]), .B(n4627), .Z(n4628) );
  XOR U1059 ( .A(y[127]), .B(n4611), .Z(n4612) );
  XOR U1060 ( .A(y[131]), .B(n4595), .Z(n4596) );
  XOR U1061 ( .A(y[135]), .B(n4579), .Z(n4580) );
  XOR U1062 ( .A(y[139]), .B(n4563), .Z(n4564) );
  XOR U1063 ( .A(y[143]), .B(n4547), .Z(n4548) );
  XOR U1064 ( .A(y[147]), .B(n4531), .Z(n4532) );
  XOR U1065 ( .A(y[151]), .B(n4515), .Z(n4516) );
  XOR U1066 ( .A(y[155]), .B(n4499), .Z(n4500) );
  XOR U1067 ( .A(y[159]), .B(n4483), .Z(n4484) );
  XOR U1068 ( .A(y[163]), .B(n4467), .Z(n4468) );
  XOR U1069 ( .A(y[167]), .B(n4451), .Z(n4452) );
  XOR U1070 ( .A(y[171]), .B(n4435), .Z(n4436) );
  XOR U1071 ( .A(y[175]), .B(n4419), .Z(n4420) );
  XOR U1072 ( .A(y[179]), .B(n4403), .Z(n4404) );
  XOR U1073 ( .A(y[183]), .B(n4387), .Z(n4388) );
  XOR U1074 ( .A(y[187]), .B(n4371), .Z(n4372) );
  XOR U1075 ( .A(y[191]), .B(n4355), .Z(n4356) );
  XOR U1076 ( .A(y[195]), .B(n4339), .Z(n4340) );
  XOR U1077 ( .A(y[199]), .B(n4323), .Z(n4324) );
  XOR U1078 ( .A(y[203]), .B(n4307), .Z(n4308) );
  XOR U1079 ( .A(y[207]), .B(n4291), .Z(n4292) );
  XOR U1080 ( .A(y[211]), .B(n4275), .Z(n4276) );
  XOR U1081 ( .A(y[215]), .B(n4259), .Z(n4260) );
  XOR U1082 ( .A(y[219]), .B(n4243), .Z(n4244) );
  XOR U1083 ( .A(y[223]), .B(n4227), .Z(n4228) );
  XOR U1084 ( .A(y[227]), .B(n4211), .Z(n4212) );
  XOR U1085 ( .A(y[231]), .B(n4195), .Z(n4196) );
  XOR U1086 ( .A(y[235]), .B(n4179), .Z(n4180) );
  XOR U1087 ( .A(y[239]), .B(n4163), .Z(n4164) );
  XOR U1088 ( .A(y[243]), .B(n4147), .Z(n4148) );
  XOR U1089 ( .A(y[247]), .B(n4131), .Z(n4132) );
  XOR U1090 ( .A(y[251]), .B(n4115), .Z(n4116) );
  XOR U1091 ( .A(y[255]), .B(n4099), .Z(n4100) );
  XOR U1092 ( .A(y[259]), .B(n4083), .Z(n4084) );
  XOR U1093 ( .A(y[263]), .B(n4067), .Z(n4068) );
  XOR U1094 ( .A(y[267]), .B(n4051), .Z(n4052) );
  XOR U1095 ( .A(y[271]), .B(n4035), .Z(n4036) );
  XOR U1096 ( .A(y[275]), .B(n4019), .Z(n4020) );
  XOR U1097 ( .A(y[279]), .B(n4003), .Z(n4004) );
  XOR U1098 ( .A(y[283]), .B(n3987), .Z(n3988) );
  XOR U1099 ( .A(y[287]), .B(n3971), .Z(n3972) );
  XOR U1100 ( .A(y[291]), .B(n3955), .Z(n3956) );
  XOR U1101 ( .A(y[295]), .B(n3939), .Z(n3940) );
  XOR U1102 ( .A(y[299]), .B(n3923), .Z(n3924) );
  XOR U1103 ( .A(y[303]), .B(n3907), .Z(n3908) );
  XOR U1104 ( .A(y[307]), .B(n3891), .Z(n3892) );
  XOR U1105 ( .A(y[311]), .B(n3875), .Z(n3876) );
  XOR U1106 ( .A(y[315]), .B(n3859), .Z(n3860) );
  XOR U1107 ( .A(y[319]), .B(n3843), .Z(n3844) );
  XOR U1108 ( .A(y[323]), .B(n3827), .Z(n3828) );
  XOR U1109 ( .A(y[327]), .B(n3811), .Z(n3812) );
  XOR U1110 ( .A(y[331]), .B(n3795), .Z(n3796) );
  XOR U1111 ( .A(y[335]), .B(n3779), .Z(n3780) );
  XOR U1112 ( .A(y[339]), .B(n3763), .Z(n3764) );
  XOR U1113 ( .A(y[343]), .B(n3747), .Z(n3748) );
  XOR U1114 ( .A(y[347]), .B(n3731), .Z(n3732) );
  XOR U1115 ( .A(y[351]), .B(n3715), .Z(n3716) );
  XOR U1116 ( .A(y[355]), .B(n3699), .Z(n3700) );
  XOR U1117 ( .A(y[359]), .B(n3683), .Z(n3684) );
  XOR U1118 ( .A(y[363]), .B(n3667), .Z(n3668) );
  XOR U1119 ( .A(y[367]), .B(n3651), .Z(n3652) );
  XOR U1120 ( .A(y[371]), .B(n3635), .Z(n3636) );
  XOR U1121 ( .A(y[375]), .B(n3619), .Z(n3620) );
  XOR U1122 ( .A(y[379]), .B(n3603), .Z(n3604) );
  XOR U1123 ( .A(y[383]), .B(n3587), .Z(n3588) );
  XOR U1124 ( .A(y[387]), .B(n3571), .Z(n3572) );
  XOR U1125 ( .A(y[391]), .B(n3555), .Z(n3556) );
  XOR U1126 ( .A(y[395]), .B(n3539), .Z(n3540) );
  XOR U1127 ( .A(y[399]), .B(n3523), .Z(n3524) );
  XOR U1128 ( .A(y[403]), .B(n3507), .Z(n3508) );
  XOR U1129 ( .A(y[407]), .B(n3491), .Z(n3492) );
  XOR U1130 ( .A(y[411]), .B(n3475), .Z(n3476) );
  XOR U1131 ( .A(y[415]), .B(n3459), .Z(n3460) );
  XOR U1132 ( .A(y[419]), .B(n3443), .Z(n3444) );
  XOR U1133 ( .A(y[423]), .B(n3427), .Z(n3428) );
  XOR U1134 ( .A(y[427]), .B(n3411), .Z(n3412) );
  XOR U1135 ( .A(y[431]), .B(n3395), .Z(n3396) );
  XOR U1136 ( .A(y[435]), .B(n3379), .Z(n3380) );
  XOR U1137 ( .A(y[439]), .B(n3363), .Z(n3364) );
  XOR U1138 ( .A(y[443]), .B(n3347), .Z(n3348) );
  XOR U1139 ( .A(y[447]), .B(n3331), .Z(n3332) );
  XOR U1140 ( .A(y[451]), .B(n3315), .Z(n3316) );
  XOR U1141 ( .A(y[455]), .B(n3299), .Z(n3300) );
  XOR U1142 ( .A(y[459]), .B(n3283), .Z(n3284) );
  XOR U1143 ( .A(y[463]), .B(n3267), .Z(n3268) );
  XOR U1144 ( .A(y[467]), .B(n3251), .Z(n3252) );
  XOR U1145 ( .A(y[471]), .B(n3235), .Z(n3236) );
  XOR U1146 ( .A(y[475]), .B(n3219), .Z(n3220) );
  XOR U1147 ( .A(y[479]), .B(n3203), .Z(n3204) );
  XOR U1148 ( .A(y[483]), .B(n3187), .Z(n3188) );
  XOR U1149 ( .A(y[487]), .B(n3171), .Z(n3172) );
  XOR U1150 ( .A(y[491]), .B(n3155), .Z(n3156) );
  XOR U1151 ( .A(y[495]), .B(n3139), .Z(n3140) );
  XOR U1152 ( .A(y[499]), .B(n3123), .Z(n3124) );
  XOR U1153 ( .A(y[503]), .B(n3107), .Z(n3108) );
  XOR U1154 ( .A(y[507]), .B(n3091), .Z(n3092) );
  XOR U1155 ( .A(y[511]), .B(n3075), .Z(n3076) );
  XOR U1156 ( .A(y[515]), .B(n3059), .Z(n3060) );
  XOR U1157 ( .A(y[519]), .B(n3043), .Z(n3044) );
  XOR U1158 ( .A(y[523]), .B(n3027), .Z(n3028) );
  XOR U1159 ( .A(y[527]), .B(n3011), .Z(n3012) );
  XOR U1160 ( .A(y[531]), .B(n2995), .Z(n2996) );
  XOR U1161 ( .A(y[535]), .B(n2979), .Z(n2980) );
  XOR U1162 ( .A(y[539]), .B(n2963), .Z(n2964) );
  XOR U1163 ( .A(y[543]), .B(n2947), .Z(n2948) );
  XOR U1164 ( .A(y[547]), .B(n2931), .Z(n2932) );
  XOR U1165 ( .A(y[551]), .B(n2915), .Z(n2916) );
  XOR U1166 ( .A(y[555]), .B(n2899), .Z(n2900) );
  XOR U1167 ( .A(y[559]), .B(n2883), .Z(n2884) );
  XOR U1168 ( .A(y[563]), .B(n2867), .Z(n2868) );
  XOR U1169 ( .A(y[567]), .B(n2851), .Z(n2852) );
  XOR U1170 ( .A(y[571]), .B(n2835), .Z(n2836) );
  XOR U1171 ( .A(y[575]), .B(n2819), .Z(n2820) );
  XOR U1172 ( .A(y[579]), .B(n2803), .Z(n2804) );
  XOR U1173 ( .A(y[583]), .B(n2787), .Z(n2788) );
  XOR U1174 ( .A(y[587]), .B(n2771), .Z(n2772) );
  XOR U1175 ( .A(y[591]), .B(n2755), .Z(n2756) );
  XOR U1176 ( .A(y[595]), .B(n2739), .Z(n2740) );
  XOR U1177 ( .A(y[599]), .B(n2723), .Z(n2724) );
  XOR U1178 ( .A(y[603]), .B(n2707), .Z(n2708) );
  XOR U1179 ( .A(y[607]), .B(n2691), .Z(n2692) );
  XOR U1180 ( .A(y[611]), .B(n2675), .Z(n2676) );
  XOR U1181 ( .A(y[615]), .B(n2659), .Z(n2660) );
  XOR U1182 ( .A(y[619]), .B(n2643), .Z(n2644) );
  XOR U1183 ( .A(y[623]), .B(n2627), .Z(n2628) );
  XOR U1184 ( .A(y[627]), .B(n2611), .Z(n2612) );
  XOR U1185 ( .A(y[631]), .B(n2595), .Z(n2596) );
  XOR U1186 ( .A(y[635]), .B(n2579), .Z(n2580) );
  XOR U1187 ( .A(y[639]), .B(n2563), .Z(n2564) );
  XOR U1188 ( .A(y[643]), .B(n2547), .Z(n2548) );
  XOR U1189 ( .A(y[647]), .B(n2531), .Z(n2532) );
  XOR U1190 ( .A(y[651]), .B(n2515), .Z(n2516) );
  XOR U1191 ( .A(y[655]), .B(n2499), .Z(n2500) );
  XOR U1192 ( .A(y[659]), .B(n2483), .Z(n2484) );
  XOR U1193 ( .A(y[663]), .B(n2467), .Z(n2468) );
  XOR U1194 ( .A(y[667]), .B(n2451), .Z(n2452) );
  XOR U1195 ( .A(y[671]), .B(n2435), .Z(n2436) );
  XOR U1196 ( .A(y[675]), .B(n2419), .Z(n2420) );
  XOR U1197 ( .A(y[679]), .B(n2403), .Z(n2404) );
  XOR U1198 ( .A(y[683]), .B(n2387), .Z(n2388) );
  XOR U1199 ( .A(y[687]), .B(n2371), .Z(n2372) );
  XOR U1200 ( .A(y[691]), .B(n2355), .Z(n2356) );
  XOR U1201 ( .A(y[695]), .B(n2339), .Z(n2340) );
  XOR U1202 ( .A(y[699]), .B(n2323), .Z(n2324) );
  XOR U1203 ( .A(y[703]), .B(n2307), .Z(n2308) );
  XOR U1204 ( .A(y[707]), .B(n2291), .Z(n2292) );
  XOR U1205 ( .A(y[711]), .B(n2275), .Z(n2276) );
  XOR U1206 ( .A(y[715]), .B(n2259), .Z(n2260) );
  XOR U1207 ( .A(y[719]), .B(n2243), .Z(n2244) );
  XOR U1208 ( .A(y[723]), .B(n2227), .Z(n2228) );
  XOR U1209 ( .A(y[727]), .B(n2211), .Z(n2212) );
  XOR U1210 ( .A(y[731]), .B(n2195), .Z(n2196) );
  XOR U1211 ( .A(y[735]), .B(n2179), .Z(n2180) );
  XOR U1212 ( .A(y[739]), .B(n2163), .Z(n2164) );
  XOR U1213 ( .A(y[743]), .B(n2147), .Z(n2148) );
  XOR U1214 ( .A(y[747]), .B(n2131), .Z(n2132) );
  XOR U1215 ( .A(y[751]), .B(n2115), .Z(n2116) );
  XOR U1216 ( .A(y[755]), .B(n2099), .Z(n2100) );
  XOR U1217 ( .A(y[759]), .B(n2083), .Z(n2084) );
  XOR U1218 ( .A(y[763]), .B(n2067), .Z(n2068) );
  XOR U1219 ( .A(y[767]), .B(n2051), .Z(n2052) );
  XOR U1220 ( .A(y[771]), .B(n2035), .Z(n2036) );
  XOR U1221 ( .A(y[775]), .B(n2019), .Z(n2020) );
  XOR U1222 ( .A(y[779]), .B(n2003), .Z(n2004) );
  XOR U1223 ( .A(y[783]), .B(n1987), .Z(n1988) );
  XOR U1224 ( .A(y[787]), .B(n1971), .Z(n1972) );
  XOR U1225 ( .A(y[791]), .B(n1955), .Z(n1956) );
  XOR U1226 ( .A(y[795]), .B(n1939), .Z(n1940) );
  XOR U1227 ( .A(y[799]), .B(n1923), .Z(n1924) );
  XOR U1228 ( .A(y[803]), .B(n1907), .Z(n1908) );
  XOR U1229 ( .A(y[807]), .B(n1891), .Z(n1892) );
  XOR U1230 ( .A(y[811]), .B(n1875), .Z(n1876) );
  XOR U1231 ( .A(y[815]), .B(n1859), .Z(n1860) );
  XOR U1232 ( .A(y[819]), .B(n1843), .Z(n1844) );
  XOR U1233 ( .A(y[823]), .B(n1827), .Z(n1828) );
  XOR U1234 ( .A(y[827]), .B(n1811), .Z(n1812) );
  XOR U1235 ( .A(y[831]), .B(n1795), .Z(n1796) );
  XOR U1236 ( .A(y[835]), .B(n1779), .Z(n1780) );
  XOR U1237 ( .A(y[839]), .B(n1763), .Z(n1764) );
  XOR U1238 ( .A(y[843]), .B(n1747), .Z(n1748) );
  XOR U1239 ( .A(y[847]), .B(n1731), .Z(n1732) );
  XOR U1240 ( .A(y[851]), .B(n1715), .Z(n1716) );
  XOR U1241 ( .A(y[855]), .B(n1699), .Z(n1700) );
  XOR U1242 ( .A(y[859]), .B(n1683), .Z(n1684) );
  XOR U1243 ( .A(y[863]), .B(n1667), .Z(n1668) );
  XOR U1244 ( .A(y[867]), .B(n1651), .Z(n1652) );
  XOR U1245 ( .A(y[871]), .B(n1635), .Z(n1636) );
  XOR U1246 ( .A(y[875]), .B(n1619), .Z(n1620) );
  XOR U1247 ( .A(y[879]), .B(n1603), .Z(n1604) );
  XOR U1248 ( .A(y[883]), .B(n1587), .Z(n1588) );
  XOR U1249 ( .A(y[887]), .B(n1571), .Z(n1572) );
  XOR U1250 ( .A(y[891]), .B(n1555), .Z(n1556) );
  XOR U1251 ( .A(y[895]), .B(n1539), .Z(n1540) );
  XOR U1252 ( .A(y[899]), .B(n1523), .Z(n1524) );
  XOR U1253 ( .A(y[903]), .B(n1507), .Z(n1508) );
  XOR U1254 ( .A(y[907]), .B(n1491), .Z(n1492) );
  XOR U1255 ( .A(y[911]), .B(n1475), .Z(n1476) );
  XOR U1256 ( .A(y[915]), .B(n1459), .Z(n1460) );
  XOR U1257 ( .A(y[919]), .B(n1443), .Z(n1444) );
  XOR U1258 ( .A(y[923]), .B(n1427), .Z(n1428) );
  XOR U1259 ( .A(y[927]), .B(n1411), .Z(n1412) );
  XOR U1260 ( .A(y[931]), .B(n1395), .Z(n1396) );
  XOR U1261 ( .A(y[935]), .B(n1379), .Z(n1380) );
  XOR U1262 ( .A(y[939]), .B(n1363), .Z(n1364) );
  XOR U1263 ( .A(y[943]), .B(n1347), .Z(n1348) );
  XOR U1264 ( .A(y[947]), .B(n1331), .Z(n1332) );
  XOR U1265 ( .A(y[951]), .B(n1315), .Z(n1316) );
  XOR U1266 ( .A(y[955]), .B(n1299), .Z(n1300) );
  XOR U1267 ( .A(y[959]), .B(n1283), .Z(n1284) );
  XOR U1268 ( .A(y[963]), .B(n1267), .Z(n1268) );
  XOR U1269 ( .A(y[967]), .B(n1251), .Z(n1252) );
  XOR U1270 ( .A(y[971]), .B(n1235), .Z(n1236) );
  XOR U1271 ( .A(y[975]), .B(n1219), .Z(n1220) );
  XOR U1272 ( .A(y[979]), .B(n1203), .Z(n1204) );
  XOR U1273 ( .A(y[983]), .B(n1187), .Z(n1188) );
  XOR U1274 ( .A(y[987]), .B(n1171), .Z(n1172) );
  XOR U1275 ( .A(y[991]), .B(n1155), .Z(n1156) );
  XOR U1276 ( .A(y[995]), .B(n1139), .Z(n1140) );
  XOR U1277 ( .A(y[999]), .B(n1123), .Z(n1124) );
  XOR U1278 ( .A(y[1003]), .B(n1107), .Z(n1108) );
  XOR U1279 ( .A(y[1007]), .B(n1091), .Z(n1092) );
  XOR U1280 ( .A(y[1011]), .B(n1075), .Z(n1076) );
  XOR U1281 ( .A(y[1015]), .B(n1059), .Z(n1060) );
  XOR U1282 ( .A(y[1019]), .B(n1043), .Z(n1044) );
  XOR U1283 ( .A(y[4]), .B(n5103), .Z(n5104) );
  XOR U1284 ( .A(y[8]), .B(n5087), .Z(n5088) );
  XOR U1285 ( .A(y[12]), .B(n5071), .Z(n5072) );
  XOR U1286 ( .A(y[16]), .B(n5055), .Z(n5056) );
  XOR U1287 ( .A(y[20]), .B(n5039), .Z(n5040) );
  XOR U1288 ( .A(y[24]), .B(n5023), .Z(n5024) );
  XOR U1289 ( .A(y[28]), .B(n5007), .Z(n5008) );
  XOR U1290 ( .A(y[32]), .B(n4991), .Z(n4992) );
  XOR U1291 ( .A(y[36]), .B(n4975), .Z(n4976) );
  XOR U1292 ( .A(y[40]), .B(n4959), .Z(n4960) );
  XOR U1293 ( .A(y[44]), .B(n4943), .Z(n4944) );
  XOR U1294 ( .A(y[48]), .B(n4927), .Z(n4928) );
  XOR U1295 ( .A(y[52]), .B(n4911), .Z(n4912) );
  XOR U1296 ( .A(y[56]), .B(n4895), .Z(n4896) );
  XOR U1297 ( .A(y[60]), .B(n4879), .Z(n4880) );
  XOR U1298 ( .A(y[64]), .B(n4863), .Z(n4864) );
  XOR U1299 ( .A(y[68]), .B(n4847), .Z(n4848) );
  XOR U1300 ( .A(y[72]), .B(n4831), .Z(n4832) );
  XOR U1301 ( .A(y[76]), .B(n4815), .Z(n4816) );
  XOR U1302 ( .A(y[80]), .B(n4799), .Z(n4800) );
  XOR U1303 ( .A(y[84]), .B(n4783), .Z(n4784) );
  XOR U1304 ( .A(y[88]), .B(n4767), .Z(n4768) );
  XOR U1305 ( .A(y[92]), .B(n4751), .Z(n4752) );
  XOR U1306 ( .A(y[96]), .B(n4735), .Z(n4736) );
  XOR U1307 ( .A(y[100]), .B(n4719), .Z(n4720) );
  XOR U1308 ( .A(y[104]), .B(n4703), .Z(n4704) );
  XOR U1309 ( .A(y[108]), .B(n4687), .Z(n4688) );
  XOR U1310 ( .A(y[112]), .B(n4671), .Z(n4672) );
  XOR U1311 ( .A(y[116]), .B(n4655), .Z(n4656) );
  XOR U1312 ( .A(y[120]), .B(n4639), .Z(n4640) );
  XOR U1313 ( .A(y[124]), .B(n4623), .Z(n4624) );
  XOR U1314 ( .A(y[128]), .B(n4607), .Z(n4608) );
  XOR U1315 ( .A(y[132]), .B(n4591), .Z(n4592) );
  XOR U1316 ( .A(y[136]), .B(n4575), .Z(n4576) );
  XOR U1317 ( .A(y[140]), .B(n4559), .Z(n4560) );
  XOR U1318 ( .A(y[144]), .B(n4543), .Z(n4544) );
  XOR U1319 ( .A(y[148]), .B(n4527), .Z(n4528) );
  XOR U1320 ( .A(y[152]), .B(n4511), .Z(n4512) );
  XOR U1321 ( .A(y[156]), .B(n4495), .Z(n4496) );
  XOR U1322 ( .A(y[160]), .B(n4479), .Z(n4480) );
  XOR U1323 ( .A(y[164]), .B(n4463), .Z(n4464) );
  XOR U1324 ( .A(y[168]), .B(n4447), .Z(n4448) );
  XOR U1325 ( .A(y[172]), .B(n4431), .Z(n4432) );
  XOR U1326 ( .A(y[176]), .B(n4415), .Z(n4416) );
  XOR U1327 ( .A(y[180]), .B(n4399), .Z(n4400) );
  XOR U1328 ( .A(y[184]), .B(n4383), .Z(n4384) );
  XOR U1329 ( .A(y[188]), .B(n4367), .Z(n4368) );
  XOR U1330 ( .A(y[192]), .B(n4351), .Z(n4352) );
  XOR U1331 ( .A(y[196]), .B(n4335), .Z(n4336) );
  XOR U1332 ( .A(y[200]), .B(n4319), .Z(n4320) );
  XOR U1333 ( .A(y[204]), .B(n4303), .Z(n4304) );
  XOR U1334 ( .A(y[208]), .B(n4287), .Z(n4288) );
  XOR U1335 ( .A(y[212]), .B(n4271), .Z(n4272) );
  XOR U1336 ( .A(y[216]), .B(n4255), .Z(n4256) );
  XOR U1337 ( .A(y[220]), .B(n4239), .Z(n4240) );
  XOR U1338 ( .A(y[224]), .B(n4223), .Z(n4224) );
  XOR U1339 ( .A(y[228]), .B(n4207), .Z(n4208) );
  XOR U1340 ( .A(y[232]), .B(n4191), .Z(n4192) );
  XOR U1341 ( .A(y[236]), .B(n4175), .Z(n4176) );
  XOR U1342 ( .A(y[240]), .B(n4159), .Z(n4160) );
  XOR U1343 ( .A(y[244]), .B(n4143), .Z(n4144) );
  XOR U1344 ( .A(y[248]), .B(n4127), .Z(n4128) );
  XOR U1345 ( .A(y[252]), .B(n4111), .Z(n4112) );
  XOR U1346 ( .A(y[256]), .B(n4095), .Z(n4096) );
  XOR U1347 ( .A(y[260]), .B(n4079), .Z(n4080) );
  XOR U1348 ( .A(y[264]), .B(n4063), .Z(n4064) );
  XOR U1349 ( .A(y[268]), .B(n4047), .Z(n4048) );
  XOR U1350 ( .A(y[272]), .B(n4031), .Z(n4032) );
  XOR U1351 ( .A(y[276]), .B(n4015), .Z(n4016) );
  XOR U1352 ( .A(y[280]), .B(n3999), .Z(n4000) );
  XOR U1353 ( .A(y[284]), .B(n3983), .Z(n3984) );
  XOR U1354 ( .A(y[288]), .B(n3967), .Z(n3968) );
  XOR U1355 ( .A(y[292]), .B(n3951), .Z(n3952) );
  XOR U1356 ( .A(y[296]), .B(n3935), .Z(n3936) );
  XOR U1357 ( .A(y[300]), .B(n3919), .Z(n3920) );
  XOR U1358 ( .A(y[304]), .B(n3903), .Z(n3904) );
  XOR U1359 ( .A(y[308]), .B(n3887), .Z(n3888) );
  XOR U1360 ( .A(y[312]), .B(n3871), .Z(n3872) );
  XOR U1361 ( .A(y[316]), .B(n3855), .Z(n3856) );
  XOR U1362 ( .A(y[320]), .B(n3839), .Z(n3840) );
  XOR U1363 ( .A(y[324]), .B(n3823), .Z(n3824) );
  XOR U1364 ( .A(y[328]), .B(n3807), .Z(n3808) );
  XOR U1365 ( .A(y[332]), .B(n3791), .Z(n3792) );
  XOR U1366 ( .A(y[336]), .B(n3775), .Z(n3776) );
  XOR U1367 ( .A(y[340]), .B(n3759), .Z(n3760) );
  XOR U1368 ( .A(y[344]), .B(n3743), .Z(n3744) );
  XOR U1369 ( .A(y[348]), .B(n3727), .Z(n3728) );
  XOR U1370 ( .A(y[352]), .B(n3711), .Z(n3712) );
  XOR U1371 ( .A(y[356]), .B(n3695), .Z(n3696) );
  XOR U1372 ( .A(y[360]), .B(n3679), .Z(n3680) );
  XOR U1373 ( .A(y[364]), .B(n3663), .Z(n3664) );
  XOR U1374 ( .A(y[368]), .B(n3647), .Z(n3648) );
  XOR U1375 ( .A(y[372]), .B(n3631), .Z(n3632) );
  XOR U1376 ( .A(y[376]), .B(n3615), .Z(n3616) );
  XOR U1377 ( .A(y[380]), .B(n3599), .Z(n3600) );
  XOR U1378 ( .A(y[384]), .B(n3583), .Z(n3584) );
  XOR U1379 ( .A(y[388]), .B(n3567), .Z(n3568) );
  XOR U1380 ( .A(y[392]), .B(n3551), .Z(n3552) );
  XOR U1381 ( .A(y[396]), .B(n3535), .Z(n3536) );
  XOR U1382 ( .A(y[400]), .B(n3519), .Z(n3520) );
  XOR U1383 ( .A(y[404]), .B(n3503), .Z(n3504) );
  XOR U1384 ( .A(y[408]), .B(n3487), .Z(n3488) );
  XOR U1385 ( .A(y[412]), .B(n3471), .Z(n3472) );
  XOR U1386 ( .A(y[416]), .B(n3455), .Z(n3456) );
  XOR U1387 ( .A(y[420]), .B(n3439), .Z(n3440) );
  XOR U1388 ( .A(y[424]), .B(n3423), .Z(n3424) );
  XOR U1389 ( .A(y[428]), .B(n3407), .Z(n3408) );
  XOR U1390 ( .A(y[432]), .B(n3391), .Z(n3392) );
  XOR U1391 ( .A(y[436]), .B(n3375), .Z(n3376) );
  XOR U1392 ( .A(y[440]), .B(n3359), .Z(n3360) );
  XOR U1393 ( .A(y[444]), .B(n3343), .Z(n3344) );
  XOR U1394 ( .A(y[448]), .B(n3327), .Z(n3328) );
  XOR U1395 ( .A(y[452]), .B(n3311), .Z(n3312) );
  XOR U1396 ( .A(y[456]), .B(n3295), .Z(n3296) );
  XOR U1397 ( .A(y[460]), .B(n3279), .Z(n3280) );
  XOR U1398 ( .A(y[464]), .B(n3263), .Z(n3264) );
  XOR U1399 ( .A(y[468]), .B(n3247), .Z(n3248) );
  XOR U1400 ( .A(y[472]), .B(n3231), .Z(n3232) );
  XOR U1401 ( .A(y[476]), .B(n3215), .Z(n3216) );
  XOR U1402 ( .A(y[480]), .B(n3199), .Z(n3200) );
  XOR U1403 ( .A(y[484]), .B(n3183), .Z(n3184) );
  XOR U1404 ( .A(y[488]), .B(n3167), .Z(n3168) );
  XOR U1405 ( .A(y[492]), .B(n3151), .Z(n3152) );
  XOR U1406 ( .A(y[496]), .B(n3135), .Z(n3136) );
  XOR U1407 ( .A(y[500]), .B(n3119), .Z(n3120) );
  XOR U1408 ( .A(y[504]), .B(n3103), .Z(n3104) );
  XOR U1409 ( .A(y[508]), .B(n3087), .Z(n3088) );
  XOR U1410 ( .A(y[512]), .B(n3071), .Z(n3072) );
  XOR U1411 ( .A(y[516]), .B(n3055), .Z(n3056) );
  XOR U1412 ( .A(y[520]), .B(n3039), .Z(n3040) );
  XOR U1413 ( .A(y[524]), .B(n3023), .Z(n3024) );
  XOR U1414 ( .A(y[528]), .B(n3007), .Z(n3008) );
  XOR U1415 ( .A(y[532]), .B(n2991), .Z(n2992) );
  XOR U1416 ( .A(y[536]), .B(n2975), .Z(n2976) );
  XOR U1417 ( .A(y[540]), .B(n2959), .Z(n2960) );
  XOR U1418 ( .A(y[544]), .B(n2943), .Z(n2944) );
  XOR U1419 ( .A(y[548]), .B(n2927), .Z(n2928) );
  XOR U1420 ( .A(y[552]), .B(n2911), .Z(n2912) );
  XOR U1421 ( .A(y[556]), .B(n2895), .Z(n2896) );
  XOR U1422 ( .A(y[560]), .B(n2879), .Z(n2880) );
  XOR U1423 ( .A(y[564]), .B(n2863), .Z(n2864) );
  XOR U1424 ( .A(y[568]), .B(n2847), .Z(n2848) );
  XOR U1425 ( .A(y[572]), .B(n2831), .Z(n2832) );
  XOR U1426 ( .A(y[576]), .B(n2815), .Z(n2816) );
  XOR U1427 ( .A(y[580]), .B(n2799), .Z(n2800) );
  XOR U1428 ( .A(y[584]), .B(n2783), .Z(n2784) );
  XOR U1429 ( .A(y[588]), .B(n2767), .Z(n2768) );
  XOR U1430 ( .A(y[592]), .B(n2751), .Z(n2752) );
  XOR U1431 ( .A(y[596]), .B(n2735), .Z(n2736) );
  XOR U1432 ( .A(y[600]), .B(n2719), .Z(n2720) );
  XOR U1433 ( .A(y[604]), .B(n2703), .Z(n2704) );
  XOR U1434 ( .A(y[608]), .B(n2687), .Z(n2688) );
  XOR U1435 ( .A(y[612]), .B(n2671), .Z(n2672) );
  XOR U1436 ( .A(y[616]), .B(n2655), .Z(n2656) );
  XOR U1437 ( .A(y[620]), .B(n2639), .Z(n2640) );
  XOR U1438 ( .A(y[624]), .B(n2623), .Z(n2624) );
  XOR U1439 ( .A(y[628]), .B(n2607), .Z(n2608) );
  XOR U1440 ( .A(y[632]), .B(n2591), .Z(n2592) );
  XOR U1441 ( .A(y[636]), .B(n2575), .Z(n2576) );
  XOR U1442 ( .A(y[640]), .B(n2559), .Z(n2560) );
  XOR U1443 ( .A(y[644]), .B(n2543), .Z(n2544) );
  XOR U1444 ( .A(y[648]), .B(n2527), .Z(n2528) );
  XOR U1445 ( .A(y[652]), .B(n2511), .Z(n2512) );
  XOR U1446 ( .A(y[656]), .B(n2495), .Z(n2496) );
  XOR U1447 ( .A(y[660]), .B(n2479), .Z(n2480) );
  XOR U1448 ( .A(y[664]), .B(n2463), .Z(n2464) );
  XOR U1449 ( .A(y[668]), .B(n2447), .Z(n2448) );
  XOR U1450 ( .A(y[672]), .B(n2431), .Z(n2432) );
  XOR U1451 ( .A(y[676]), .B(n2415), .Z(n2416) );
  XOR U1452 ( .A(y[680]), .B(n2399), .Z(n2400) );
  XOR U1453 ( .A(y[684]), .B(n2383), .Z(n2384) );
  XOR U1454 ( .A(y[688]), .B(n2367), .Z(n2368) );
  XOR U1455 ( .A(y[692]), .B(n2351), .Z(n2352) );
  XOR U1456 ( .A(y[696]), .B(n2335), .Z(n2336) );
  XOR U1457 ( .A(y[700]), .B(n2319), .Z(n2320) );
  XOR U1458 ( .A(y[704]), .B(n2303), .Z(n2304) );
  XOR U1459 ( .A(y[708]), .B(n2287), .Z(n2288) );
  XOR U1460 ( .A(y[712]), .B(n2271), .Z(n2272) );
  XOR U1461 ( .A(y[716]), .B(n2255), .Z(n2256) );
  XOR U1462 ( .A(y[720]), .B(n2239), .Z(n2240) );
  XOR U1463 ( .A(y[724]), .B(n2223), .Z(n2224) );
  XOR U1464 ( .A(y[728]), .B(n2207), .Z(n2208) );
  XOR U1465 ( .A(y[732]), .B(n2191), .Z(n2192) );
  XOR U1466 ( .A(y[736]), .B(n2175), .Z(n2176) );
  XOR U1467 ( .A(y[740]), .B(n2159), .Z(n2160) );
  XOR U1468 ( .A(y[744]), .B(n2143), .Z(n2144) );
  XOR U1469 ( .A(y[748]), .B(n2127), .Z(n2128) );
  XOR U1470 ( .A(y[752]), .B(n2111), .Z(n2112) );
  XOR U1471 ( .A(y[756]), .B(n2095), .Z(n2096) );
  XOR U1472 ( .A(y[760]), .B(n2079), .Z(n2080) );
  XOR U1473 ( .A(y[764]), .B(n2063), .Z(n2064) );
  XOR U1474 ( .A(y[768]), .B(n2047), .Z(n2048) );
  XOR U1475 ( .A(y[772]), .B(n2031), .Z(n2032) );
  XOR U1476 ( .A(y[776]), .B(n2015), .Z(n2016) );
  XOR U1477 ( .A(y[780]), .B(n1999), .Z(n2000) );
  XOR U1478 ( .A(y[784]), .B(n1983), .Z(n1984) );
  XOR U1479 ( .A(y[788]), .B(n1967), .Z(n1968) );
  XOR U1480 ( .A(y[792]), .B(n1951), .Z(n1952) );
  XOR U1481 ( .A(y[796]), .B(n1935), .Z(n1936) );
  XOR U1482 ( .A(y[800]), .B(n1919), .Z(n1920) );
  XOR U1483 ( .A(y[804]), .B(n1903), .Z(n1904) );
  XOR U1484 ( .A(y[808]), .B(n1887), .Z(n1888) );
  XOR U1485 ( .A(y[812]), .B(n1871), .Z(n1872) );
  XOR U1486 ( .A(y[816]), .B(n1855), .Z(n1856) );
  XOR U1487 ( .A(y[820]), .B(n1839), .Z(n1840) );
  XOR U1488 ( .A(y[824]), .B(n1823), .Z(n1824) );
  XOR U1489 ( .A(y[828]), .B(n1807), .Z(n1808) );
  XOR U1490 ( .A(y[832]), .B(n1791), .Z(n1792) );
  XOR U1491 ( .A(y[836]), .B(n1775), .Z(n1776) );
  XOR U1492 ( .A(y[840]), .B(n1759), .Z(n1760) );
  XOR U1493 ( .A(y[844]), .B(n1743), .Z(n1744) );
  XOR U1494 ( .A(y[848]), .B(n1727), .Z(n1728) );
  XOR U1495 ( .A(y[852]), .B(n1711), .Z(n1712) );
  XOR U1496 ( .A(y[856]), .B(n1695), .Z(n1696) );
  XOR U1497 ( .A(y[860]), .B(n1679), .Z(n1680) );
  XOR U1498 ( .A(y[864]), .B(n1663), .Z(n1664) );
  XOR U1499 ( .A(y[868]), .B(n1647), .Z(n1648) );
  XOR U1500 ( .A(y[872]), .B(n1631), .Z(n1632) );
  XOR U1501 ( .A(y[876]), .B(n1615), .Z(n1616) );
  XOR U1502 ( .A(y[880]), .B(n1599), .Z(n1600) );
  XOR U1503 ( .A(y[884]), .B(n1583), .Z(n1584) );
  XOR U1504 ( .A(y[888]), .B(n1567), .Z(n1568) );
  XOR U1505 ( .A(y[892]), .B(n1551), .Z(n1552) );
  XOR U1506 ( .A(y[896]), .B(n1535), .Z(n1536) );
  XOR U1507 ( .A(y[900]), .B(n1519), .Z(n1520) );
  XOR U1508 ( .A(y[904]), .B(n1503), .Z(n1504) );
  XOR U1509 ( .A(y[908]), .B(n1487), .Z(n1488) );
  XOR U1510 ( .A(y[912]), .B(n1471), .Z(n1472) );
  XOR U1511 ( .A(y[916]), .B(n1455), .Z(n1456) );
  XOR U1512 ( .A(y[920]), .B(n1439), .Z(n1440) );
  XOR U1513 ( .A(y[924]), .B(n1423), .Z(n1424) );
  XOR U1514 ( .A(y[928]), .B(n1407), .Z(n1408) );
  XOR U1515 ( .A(y[932]), .B(n1391), .Z(n1392) );
  XOR U1516 ( .A(y[936]), .B(n1375), .Z(n1376) );
  XOR U1517 ( .A(y[940]), .B(n1359), .Z(n1360) );
  XOR U1518 ( .A(y[944]), .B(n1343), .Z(n1344) );
  XOR U1519 ( .A(y[948]), .B(n1327), .Z(n1328) );
  XOR U1520 ( .A(y[952]), .B(n1311), .Z(n1312) );
  XOR U1521 ( .A(y[956]), .B(n1295), .Z(n1296) );
  XOR U1522 ( .A(y[960]), .B(n1279), .Z(n1280) );
  XOR U1523 ( .A(y[964]), .B(n1263), .Z(n1264) );
  XOR U1524 ( .A(y[968]), .B(n1247), .Z(n1248) );
  XOR U1525 ( .A(y[972]), .B(n1231), .Z(n1232) );
  XOR U1526 ( .A(y[976]), .B(n1215), .Z(n1216) );
  XOR U1527 ( .A(y[980]), .B(n1199), .Z(n1200) );
  XOR U1528 ( .A(y[984]), .B(n1183), .Z(n1184) );
  XOR U1529 ( .A(y[988]), .B(n1167), .Z(n1168) );
  XOR U1530 ( .A(y[992]), .B(n1151), .Z(n1152) );
  XOR U1531 ( .A(y[996]), .B(n1135), .Z(n1136) );
  XOR U1532 ( .A(y[1000]), .B(n1119), .Z(n1120) );
  XOR U1533 ( .A(y[1004]), .B(n1103), .Z(n1104) );
  XOR U1534 ( .A(y[1008]), .B(n1087), .Z(n1088) );
  XOR U1535 ( .A(y[1012]), .B(n1071), .Z(n1072) );
  XOR U1536 ( .A(y[1016]), .B(n1055), .Z(n1056) );
  XOR U1537 ( .A(y[1020]), .B(n1039), .Z(n1040) );
  XOR U1538 ( .A(y[5]), .B(n5099), .Z(n5100) );
  XOR U1539 ( .A(y[9]), .B(n5083), .Z(n5084) );
  XOR U1540 ( .A(y[13]), .B(n5067), .Z(n5068) );
  XOR U1541 ( .A(y[17]), .B(n5051), .Z(n5052) );
  XOR U1542 ( .A(y[21]), .B(n5035), .Z(n5036) );
  XOR U1543 ( .A(y[25]), .B(n5019), .Z(n5020) );
  XOR U1544 ( .A(y[29]), .B(n5003), .Z(n5004) );
  XOR U1545 ( .A(y[33]), .B(n4987), .Z(n4988) );
  XOR U1546 ( .A(y[37]), .B(n4971), .Z(n4972) );
  XOR U1547 ( .A(y[41]), .B(n4955), .Z(n4956) );
  XOR U1548 ( .A(y[45]), .B(n4939), .Z(n4940) );
  XOR U1549 ( .A(y[49]), .B(n4923), .Z(n4924) );
  XOR U1550 ( .A(y[53]), .B(n4907), .Z(n4908) );
  XOR U1551 ( .A(y[57]), .B(n4891), .Z(n4892) );
  XOR U1552 ( .A(y[61]), .B(n4875), .Z(n4876) );
  XOR U1553 ( .A(y[65]), .B(n4859), .Z(n4860) );
  XOR U1554 ( .A(y[69]), .B(n4843), .Z(n4844) );
  XOR U1555 ( .A(y[73]), .B(n4827), .Z(n4828) );
  XOR U1556 ( .A(y[77]), .B(n4811), .Z(n4812) );
  XOR U1557 ( .A(y[81]), .B(n4795), .Z(n4796) );
  XOR U1558 ( .A(y[85]), .B(n4779), .Z(n4780) );
  XOR U1559 ( .A(y[89]), .B(n4763), .Z(n4764) );
  XOR U1560 ( .A(y[93]), .B(n4747), .Z(n4748) );
  XOR U1561 ( .A(y[97]), .B(n4731), .Z(n4732) );
  XOR U1562 ( .A(y[101]), .B(n4715), .Z(n4716) );
  XOR U1563 ( .A(y[105]), .B(n4699), .Z(n4700) );
  XOR U1564 ( .A(y[109]), .B(n4683), .Z(n4684) );
  XOR U1565 ( .A(y[113]), .B(n4667), .Z(n4668) );
  XOR U1566 ( .A(y[117]), .B(n4651), .Z(n4652) );
  XOR U1567 ( .A(y[121]), .B(n4635), .Z(n4636) );
  XOR U1568 ( .A(y[125]), .B(n4619), .Z(n4620) );
  XOR U1569 ( .A(y[129]), .B(n4603), .Z(n4604) );
  XOR U1570 ( .A(y[133]), .B(n4587), .Z(n4588) );
  XOR U1571 ( .A(y[137]), .B(n4571), .Z(n4572) );
  XOR U1572 ( .A(y[141]), .B(n4555), .Z(n4556) );
  XOR U1573 ( .A(y[145]), .B(n4539), .Z(n4540) );
  XOR U1574 ( .A(y[149]), .B(n4523), .Z(n4524) );
  XOR U1575 ( .A(y[153]), .B(n4507), .Z(n4508) );
  XOR U1576 ( .A(y[157]), .B(n4491), .Z(n4492) );
  XOR U1577 ( .A(y[161]), .B(n4475), .Z(n4476) );
  XOR U1578 ( .A(y[165]), .B(n4459), .Z(n4460) );
  XOR U1579 ( .A(y[169]), .B(n4443), .Z(n4444) );
  XOR U1580 ( .A(y[173]), .B(n4427), .Z(n4428) );
  XOR U1581 ( .A(y[177]), .B(n4411), .Z(n4412) );
  XOR U1582 ( .A(y[181]), .B(n4395), .Z(n4396) );
  XOR U1583 ( .A(y[185]), .B(n4379), .Z(n4380) );
  XOR U1584 ( .A(y[189]), .B(n4363), .Z(n4364) );
  XOR U1585 ( .A(y[193]), .B(n4347), .Z(n4348) );
  XOR U1586 ( .A(y[197]), .B(n4331), .Z(n4332) );
  XOR U1587 ( .A(y[201]), .B(n4315), .Z(n4316) );
  XOR U1588 ( .A(y[205]), .B(n4299), .Z(n4300) );
  XOR U1589 ( .A(y[209]), .B(n4283), .Z(n4284) );
  XOR U1590 ( .A(y[213]), .B(n4267), .Z(n4268) );
  XOR U1591 ( .A(y[217]), .B(n4251), .Z(n4252) );
  XOR U1592 ( .A(y[221]), .B(n4235), .Z(n4236) );
  XOR U1593 ( .A(y[225]), .B(n4219), .Z(n4220) );
  XOR U1594 ( .A(y[229]), .B(n4203), .Z(n4204) );
  XOR U1595 ( .A(y[233]), .B(n4187), .Z(n4188) );
  XOR U1596 ( .A(y[237]), .B(n4171), .Z(n4172) );
  XOR U1597 ( .A(y[241]), .B(n4155), .Z(n4156) );
  XOR U1598 ( .A(y[245]), .B(n4139), .Z(n4140) );
  XOR U1599 ( .A(y[249]), .B(n4123), .Z(n4124) );
  XOR U1600 ( .A(y[253]), .B(n4107), .Z(n4108) );
  XOR U1601 ( .A(y[257]), .B(n4091), .Z(n4092) );
  XOR U1602 ( .A(y[261]), .B(n4075), .Z(n4076) );
  XOR U1603 ( .A(y[265]), .B(n4059), .Z(n4060) );
  XOR U1604 ( .A(y[269]), .B(n4043), .Z(n4044) );
  XOR U1605 ( .A(y[273]), .B(n4027), .Z(n4028) );
  XOR U1606 ( .A(y[277]), .B(n4011), .Z(n4012) );
  XOR U1607 ( .A(y[281]), .B(n3995), .Z(n3996) );
  XOR U1608 ( .A(y[285]), .B(n3979), .Z(n3980) );
  XOR U1609 ( .A(y[289]), .B(n3963), .Z(n3964) );
  XOR U1610 ( .A(y[293]), .B(n3947), .Z(n3948) );
  XOR U1611 ( .A(y[297]), .B(n3931), .Z(n3932) );
  XOR U1612 ( .A(y[301]), .B(n3915), .Z(n3916) );
  XOR U1613 ( .A(y[305]), .B(n3899), .Z(n3900) );
  XOR U1614 ( .A(y[309]), .B(n3883), .Z(n3884) );
  XOR U1615 ( .A(y[313]), .B(n3867), .Z(n3868) );
  XOR U1616 ( .A(y[317]), .B(n3851), .Z(n3852) );
  XOR U1617 ( .A(y[321]), .B(n3835), .Z(n3836) );
  XOR U1618 ( .A(y[325]), .B(n3819), .Z(n3820) );
  XOR U1619 ( .A(y[329]), .B(n3803), .Z(n3804) );
  XOR U1620 ( .A(y[333]), .B(n3787), .Z(n3788) );
  XOR U1621 ( .A(y[337]), .B(n3771), .Z(n3772) );
  XOR U1622 ( .A(y[341]), .B(n3755), .Z(n3756) );
  XOR U1623 ( .A(y[345]), .B(n3739), .Z(n3740) );
  XOR U1624 ( .A(y[349]), .B(n3723), .Z(n3724) );
  XOR U1625 ( .A(y[353]), .B(n3707), .Z(n3708) );
  XOR U1626 ( .A(y[357]), .B(n3691), .Z(n3692) );
  XOR U1627 ( .A(y[361]), .B(n3675), .Z(n3676) );
  XOR U1628 ( .A(y[365]), .B(n3659), .Z(n3660) );
  XOR U1629 ( .A(y[369]), .B(n3643), .Z(n3644) );
  XOR U1630 ( .A(y[373]), .B(n3627), .Z(n3628) );
  XOR U1631 ( .A(y[377]), .B(n3611), .Z(n3612) );
  XOR U1632 ( .A(y[381]), .B(n3595), .Z(n3596) );
  XOR U1633 ( .A(y[385]), .B(n3579), .Z(n3580) );
  XOR U1634 ( .A(y[389]), .B(n3563), .Z(n3564) );
  XOR U1635 ( .A(y[393]), .B(n3547), .Z(n3548) );
  XOR U1636 ( .A(y[397]), .B(n3531), .Z(n3532) );
  XOR U1637 ( .A(y[401]), .B(n3515), .Z(n3516) );
  XOR U1638 ( .A(y[405]), .B(n3499), .Z(n3500) );
  XOR U1639 ( .A(y[409]), .B(n3483), .Z(n3484) );
  XOR U1640 ( .A(y[413]), .B(n3467), .Z(n3468) );
  XOR U1641 ( .A(y[417]), .B(n3451), .Z(n3452) );
  XOR U1642 ( .A(y[421]), .B(n3435), .Z(n3436) );
  XOR U1643 ( .A(y[425]), .B(n3419), .Z(n3420) );
  XOR U1644 ( .A(y[429]), .B(n3403), .Z(n3404) );
  XOR U1645 ( .A(y[433]), .B(n3387), .Z(n3388) );
  XOR U1646 ( .A(y[437]), .B(n3371), .Z(n3372) );
  XOR U1647 ( .A(y[441]), .B(n3355), .Z(n3356) );
  XOR U1648 ( .A(y[445]), .B(n3339), .Z(n3340) );
  XOR U1649 ( .A(y[449]), .B(n3323), .Z(n3324) );
  XOR U1650 ( .A(y[453]), .B(n3307), .Z(n3308) );
  XOR U1651 ( .A(y[457]), .B(n3291), .Z(n3292) );
  XOR U1652 ( .A(y[461]), .B(n3275), .Z(n3276) );
  XOR U1653 ( .A(y[465]), .B(n3259), .Z(n3260) );
  XOR U1654 ( .A(y[469]), .B(n3243), .Z(n3244) );
  XOR U1655 ( .A(y[473]), .B(n3227), .Z(n3228) );
  XOR U1656 ( .A(y[477]), .B(n3211), .Z(n3212) );
  XOR U1657 ( .A(y[481]), .B(n3195), .Z(n3196) );
  XOR U1658 ( .A(y[485]), .B(n3179), .Z(n3180) );
  XOR U1659 ( .A(y[489]), .B(n3163), .Z(n3164) );
  XOR U1660 ( .A(y[493]), .B(n3147), .Z(n3148) );
  XOR U1661 ( .A(y[497]), .B(n3131), .Z(n3132) );
  XOR U1662 ( .A(y[501]), .B(n3115), .Z(n3116) );
  XOR U1663 ( .A(y[505]), .B(n3099), .Z(n3100) );
  XOR U1664 ( .A(y[509]), .B(n3083), .Z(n3084) );
  XOR U1665 ( .A(y[513]), .B(n3067), .Z(n3068) );
  XOR U1666 ( .A(y[517]), .B(n3051), .Z(n3052) );
  XOR U1667 ( .A(y[521]), .B(n3035), .Z(n3036) );
  XOR U1668 ( .A(y[525]), .B(n3019), .Z(n3020) );
  XOR U1669 ( .A(y[529]), .B(n3003), .Z(n3004) );
  XOR U1670 ( .A(y[533]), .B(n2987), .Z(n2988) );
  XOR U1671 ( .A(y[537]), .B(n2971), .Z(n2972) );
  XOR U1672 ( .A(y[541]), .B(n2955), .Z(n2956) );
  XOR U1673 ( .A(y[545]), .B(n2939), .Z(n2940) );
  XOR U1674 ( .A(y[549]), .B(n2923), .Z(n2924) );
  XOR U1675 ( .A(y[553]), .B(n2907), .Z(n2908) );
  XOR U1676 ( .A(y[557]), .B(n2891), .Z(n2892) );
  XOR U1677 ( .A(y[561]), .B(n2875), .Z(n2876) );
  XOR U1678 ( .A(y[565]), .B(n2859), .Z(n2860) );
  XOR U1679 ( .A(y[569]), .B(n2843), .Z(n2844) );
  XOR U1680 ( .A(y[573]), .B(n2827), .Z(n2828) );
  XOR U1681 ( .A(y[577]), .B(n2811), .Z(n2812) );
  XOR U1682 ( .A(y[581]), .B(n2795), .Z(n2796) );
  XOR U1683 ( .A(y[585]), .B(n2779), .Z(n2780) );
  XOR U1684 ( .A(y[589]), .B(n2763), .Z(n2764) );
  XOR U1685 ( .A(y[593]), .B(n2747), .Z(n2748) );
  XOR U1686 ( .A(y[597]), .B(n2731), .Z(n2732) );
  XOR U1687 ( .A(y[601]), .B(n2715), .Z(n2716) );
  XOR U1688 ( .A(y[605]), .B(n2699), .Z(n2700) );
  XOR U1689 ( .A(y[609]), .B(n2683), .Z(n2684) );
  XOR U1690 ( .A(y[613]), .B(n2667), .Z(n2668) );
  XOR U1691 ( .A(y[617]), .B(n2651), .Z(n2652) );
  XOR U1692 ( .A(y[621]), .B(n2635), .Z(n2636) );
  XOR U1693 ( .A(y[625]), .B(n2619), .Z(n2620) );
  XOR U1694 ( .A(y[629]), .B(n2603), .Z(n2604) );
  XOR U1695 ( .A(y[633]), .B(n2587), .Z(n2588) );
  XOR U1696 ( .A(y[637]), .B(n2571), .Z(n2572) );
  XOR U1697 ( .A(y[641]), .B(n2555), .Z(n2556) );
  XOR U1698 ( .A(y[645]), .B(n2539), .Z(n2540) );
  XOR U1699 ( .A(y[649]), .B(n2523), .Z(n2524) );
  XOR U1700 ( .A(y[653]), .B(n2507), .Z(n2508) );
  XOR U1701 ( .A(y[657]), .B(n2491), .Z(n2492) );
  XOR U1702 ( .A(y[661]), .B(n2475), .Z(n2476) );
  XOR U1703 ( .A(y[665]), .B(n2459), .Z(n2460) );
  XOR U1704 ( .A(y[669]), .B(n2443), .Z(n2444) );
  XOR U1705 ( .A(y[673]), .B(n2427), .Z(n2428) );
  XOR U1706 ( .A(y[677]), .B(n2411), .Z(n2412) );
  XOR U1707 ( .A(y[681]), .B(n2395), .Z(n2396) );
  XOR U1708 ( .A(y[685]), .B(n2379), .Z(n2380) );
  XOR U1709 ( .A(y[689]), .B(n2363), .Z(n2364) );
  XOR U1710 ( .A(y[693]), .B(n2347), .Z(n2348) );
  XOR U1711 ( .A(y[697]), .B(n2331), .Z(n2332) );
  XOR U1712 ( .A(y[701]), .B(n2315), .Z(n2316) );
  XOR U1713 ( .A(y[705]), .B(n2299), .Z(n2300) );
  XOR U1714 ( .A(y[709]), .B(n2283), .Z(n2284) );
  XOR U1715 ( .A(y[713]), .B(n2267), .Z(n2268) );
  XOR U1716 ( .A(y[717]), .B(n2251), .Z(n2252) );
  XOR U1717 ( .A(y[721]), .B(n2235), .Z(n2236) );
  XOR U1718 ( .A(y[725]), .B(n2219), .Z(n2220) );
  XOR U1719 ( .A(y[729]), .B(n2203), .Z(n2204) );
  XOR U1720 ( .A(y[733]), .B(n2187), .Z(n2188) );
  XOR U1721 ( .A(y[737]), .B(n2171), .Z(n2172) );
  XOR U1722 ( .A(y[741]), .B(n2155), .Z(n2156) );
  XOR U1723 ( .A(y[745]), .B(n2139), .Z(n2140) );
  XOR U1724 ( .A(y[749]), .B(n2123), .Z(n2124) );
  XOR U1725 ( .A(y[753]), .B(n2107), .Z(n2108) );
  XOR U1726 ( .A(y[757]), .B(n2091), .Z(n2092) );
  XOR U1727 ( .A(y[761]), .B(n2075), .Z(n2076) );
  XOR U1728 ( .A(y[765]), .B(n2059), .Z(n2060) );
  XOR U1729 ( .A(y[769]), .B(n2043), .Z(n2044) );
  XOR U1730 ( .A(y[773]), .B(n2027), .Z(n2028) );
  XOR U1731 ( .A(y[777]), .B(n2011), .Z(n2012) );
  XOR U1732 ( .A(y[781]), .B(n1995), .Z(n1996) );
  XOR U1733 ( .A(y[785]), .B(n1979), .Z(n1980) );
  XOR U1734 ( .A(y[789]), .B(n1963), .Z(n1964) );
  XOR U1735 ( .A(y[793]), .B(n1947), .Z(n1948) );
  XOR U1736 ( .A(y[797]), .B(n1931), .Z(n1932) );
  XOR U1737 ( .A(y[801]), .B(n1915), .Z(n1916) );
  XOR U1738 ( .A(y[805]), .B(n1899), .Z(n1900) );
  XOR U1739 ( .A(y[809]), .B(n1883), .Z(n1884) );
  XOR U1740 ( .A(y[813]), .B(n1867), .Z(n1868) );
  XOR U1741 ( .A(y[817]), .B(n1851), .Z(n1852) );
  XOR U1742 ( .A(y[821]), .B(n1835), .Z(n1836) );
  XOR U1743 ( .A(y[825]), .B(n1819), .Z(n1820) );
  XOR U1744 ( .A(y[829]), .B(n1803), .Z(n1804) );
  XOR U1745 ( .A(y[833]), .B(n1787), .Z(n1788) );
  XOR U1746 ( .A(y[837]), .B(n1771), .Z(n1772) );
  XOR U1747 ( .A(y[841]), .B(n1755), .Z(n1756) );
  XOR U1748 ( .A(y[845]), .B(n1739), .Z(n1740) );
  XOR U1749 ( .A(y[849]), .B(n1723), .Z(n1724) );
  XOR U1750 ( .A(y[853]), .B(n1707), .Z(n1708) );
  XOR U1751 ( .A(y[857]), .B(n1691), .Z(n1692) );
  XOR U1752 ( .A(y[861]), .B(n1675), .Z(n1676) );
  XOR U1753 ( .A(y[865]), .B(n1659), .Z(n1660) );
  XOR U1754 ( .A(y[869]), .B(n1643), .Z(n1644) );
  XOR U1755 ( .A(y[873]), .B(n1627), .Z(n1628) );
  XOR U1756 ( .A(y[877]), .B(n1611), .Z(n1612) );
  XOR U1757 ( .A(y[881]), .B(n1595), .Z(n1596) );
  XOR U1758 ( .A(y[885]), .B(n1579), .Z(n1580) );
  XOR U1759 ( .A(y[889]), .B(n1563), .Z(n1564) );
  XOR U1760 ( .A(y[893]), .B(n1547), .Z(n1548) );
  XOR U1761 ( .A(y[897]), .B(n1531), .Z(n1532) );
  XOR U1762 ( .A(y[901]), .B(n1515), .Z(n1516) );
  XOR U1763 ( .A(y[905]), .B(n1499), .Z(n1500) );
  XOR U1764 ( .A(y[909]), .B(n1483), .Z(n1484) );
  XOR U1765 ( .A(y[913]), .B(n1467), .Z(n1468) );
  XOR U1766 ( .A(y[917]), .B(n1451), .Z(n1452) );
  XOR U1767 ( .A(y[921]), .B(n1435), .Z(n1436) );
  XOR U1768 ( .A(y[925]), .B(n1419), .Z(n1420) );
  XOR U1769 ( .A(y[929]), .B(n1403), .Z(n1404) );
  XOR U1770 ( .A(y[933]), .B(n1387), .Z(n1388) );
  XOR U1771 ( .A(y[937]), .B(n1371), .Z(n1372) );
  XOR U1772 ( .A(y[941]), .B(n1355), .Z(n1356) );
  XOR U1773 ( .A(y[945]), .B(n1339), .Z(n1340) );
  XOR U1774 ( .A(y[949]), .B(n1323), .Z(n1324) );
  XOR U1775 ( .A(y[953]), .B(n1307), .Z(n1308) );
  XOR U1776 ( .A(y[957]), .B(n1291), .Z(n1292) );
  XOR U1777 ( .A(y[961]), .B(n1275), .Z(n1276) );
  XOR U1778 ( .A(y[965]), .B(n1259), .Z(n1260) );
  XOR U1779 ( .A(y[969]), .B(n1243), .Z(n1244) );
  XOR U1780 ( .A(y[973]), .B(n1227), .Z(n1228) );
  XOR U1781 ( .A(y[977]), .B(n1211), .Z(n1212) );
  XOR U1782 ( .A(y[981]), .B(n1195), .Z(n1196) );
  XOR U1783 ( .A(y[985]), .B(n1179), .Z(n1180) );
  XOR U1784 ( .A(y[989]), .B(n1163), .Z(n1164) );
  XOR U1785 ( .A(y[993]), .B(n1147), .Z(n1148) );
  XOR U1786 ( .A(y[997]), .B(n1131), .Z(n1132) );
  XOR U1787 ( .A(y[1001]), .B(n1115), .Z(n1116) );
  XOR U1788 ( .A(y[1005]), .B(n1099), .Z(n1100) );
  XOR U1789 ( .A(y[1009]), .B(n1083), .Z(n1084) );
  XOR U1790 ( .A(y[1013]), .B(n1067), .Z(n1068) );
  XOR U1791 ( .A(y[1017]), .B(n1051), .Z(n1052) );
  XOR U1792 ( .A(y[1021]), .B(n1035), .Z(n1036) );
  XOR U1793 ( .A(y[2]), .B(n5111), .Z(n5112) );
  XOR U1794 ( .A(y[6]), .B(n5095), .Z(n5096) );
  XOR U1795 ( .A(y[10]), .B(n5079), .Z(n5080) );
  XOR U1796 ( .A(y[14]), .B(n5063), .Z(n5064) );
  XOR U1797 ( .A(y[18]), .B(n5047), .Z(n5048) );
  XOR U1798 ( .A(y[22]), .B(n5031), .Z(n5032) );
  XOR U1799 ( .A(y[26]), .B(n5015), .Z(n5016) );
  XOR U1800 ( .A(y[30]), .B(n4999), .Z(n5000) );
  XOR U1801 ( .A(y[34]), .B(n4983), .Z(n4984) );
  XOR U1802 ( .A(y[38]), .B(n4967), .Z(n4968) );
  XOR U1803 ( .A(y[42]), .B(n4951), .Z(n4952) );
  XOR U1804 ( .A(y[46]), .B(n4935), .Z(n4936) );
  XOR U1805 ( .A(y[50]), .B(n4919), .Z(n4920) );
  XOR U1806 ( .A(y[54]), .B(n4903), .Z(n4904) );
  XOR U1807 ( .A(y[58]), .B(n4887), .Z(n4888) );
  XOR U1808 ( .A(y[62]), .B(n4871), .Z(n4872) );
  XOR U1809 ( .A(y[66]), .B(n4855), .Z(n4856) );
  XOR U1810 ( .A(y[70]), .B(n4839), .Z(n4840) );
  XOR U1811 ( .A(y[74]), .B(n4823), .Z(n4824) );
  XOR U1812 ( .A(y[78]), .B(n4807), .Z(n4808) );
  XOR U1813 ( .A(y[82]), .B(n4791), .Z(n4792) );
  XOR U1814 ( .A(y[86]), .B(n4775), .Z(n4776) );
  XOR U1815 ( .A(y[90]), .B(n4759), .Z(n4760) );
  XOR U1816 ( .A(y[94]), .B(n4743), .Z(n4744) );
  XOR U1817 ( .A(y[98]), .B(n4727), .Z(n4728) );
  XOR U1818 ( .A(y[102]), .B(n4711), .Z(n4712) );
  XOR U1819 ( .A(y[106]), .B(n4695), .Z(n4696) );
  XOR U1820 ( .A(y[110]), .B(n4679), .Z(n4680) );
  XOR U1821 ( .A(y[114]), .B(n4663), .Z(n4664) );
  XOR U1822 ( .A(y[118]), .B(n4647), .Z(n4648) );
  XOR U1823 ( .A(y[122]), .B(n4631), .Z(n4632) );
  XOR U1824 ( .A(y[126]), .B(n4615), .Z(n4616) );
  XOR U1825 ( .A(y[130]), .B(n4599), .Z(n4600) );
  XOR U1826 ( .A(y[134]), .B(n4583), .Z(n4584) );
  XOR U1827 ( .A(y[138]), .B(n4567), .Z(n4568) );
  XOR U1828 ( .A(y[142]), .B(n4551), .Z(n4552) );
  XOR U1829 ( .A(y[146]), .B(n4535), .Z(n4536) );
  XOR U1830 ( .A(y[150]), .B(n4519), .Z(n4520) );
  XOR U1831 ( .A(y[154]), .B(n4503), .Z(n4504) );
  XOR U1832 ( .A(y[158]), .B(n4487), .Z(n4488) );
  XOR U1833 ( .A(y[162]), .B(n4471), .Z(n4472) );
  XOR U1834 ( .A(y[166]), .B(n4455), .Z(n4456) );
  XOR U1835 ( .A(y[170]), .B(n4439), .Z(n4440) );
  XOR U1836 ( .A(y[174]), .B(n4423), .Z(n4424) );
  XOR U1837 ( .A(y[178]), .B(n4407), .Z(n4408) );
  XOR U1838 ( .A(y[182]), .B(n4391), .Z(n4392) );
  XOR U1839 ( .A(y[186]), .B(n4375), .Z(n4376) );
  XOR U1840 ( .A(y[190]), .B(n4359), .Z(n4360) );
  XOR U1841 ( .A(y[194]), .B(n4343), .Z(n4344) );
  XOR U1842 ( .A(y[198]), .B(n4327), .Z(n4328) );
  XOR U1843 ( .A(y[202]), .B(n4311), .Z(n4312) );
  XOR U1844 ( .A(y[206]), .B(n4295), .Z(n4296) );
  XOR U1845 ( .A(y[210]), .B(n4279), .Z(n4280) );
  XOR U1846 ( .A(y[214]), .B(n4263), .Z(n4264) );
  XOR U1847 ( .A(y[218]), .B(n4247), .Z(n4248) );
  XOR U1848 ( .A(y[222]), .B(n4231), .Z(n4232) );
  XOR U1849 ( .A(y[226]), .B(n4215), .Z(n4216) );
  XOR U1850 ( .A(y[230]), .B(n4199), .Z(n4200) );
  XOR U1851 ( .A(y[234]), .B(n4183), .Z(n4184) );
  XOR U1852 ( .A(y[238]), .B(n4167), .Z(n4168) );
  XOR U1853 ( .A(y[242]), .B(n4151), .Z(n4152) );
  XOR U1854 ( .A(y[246]), .B(n4135), .Z(n4136) );
  XOR U1855 ( .A(y[250]), .B(n4119), .Z(n4120) );
  XOR U1856 ( .A(y[254]), .B(n4103), .Z(n4104) );
  XOR U1857 ( .A(y[258]), .B(n4087), .Z(n4088) );
  XOR U1858 ( .A(y[262]), .B(n4071), .Z(n4072) );
  XOR U1859 ( .A(y[266]), .B(n4055), .Z(n4056) );
  XOR U1860 ( .A(y[270]), .B(n4039), .Z(n4040) );
  XOR U1861 ( .A(y[274]), .B(n4023), .Z(n4024) );
  XOR U1862 ( .A(y[278]), .B(n4007), .Z(n4008) );
  XOR U1863 ( .A(y[282]), .B(n3991), .Z(n3992) );
  XOR U1864 ( .A(y[286]), .B(n3975), .Z(n3976) );
  XOR U1865 ( .A(y[290]), .B(n3959), .Z(n3960) );
  XOR U1866 ( .A(y[294]), .B(n3943), .Z(n3944) );
  XOR U1867 ( .A(y[298]), .B(n3927), .Z(n3928) );
  XOR U1868 ( .A(y[302]), .B(n3911), .Z(n3912) );
  XOR U1869 ( .A(y[306]), .B(n3895), .Z(n3896) );
  XOR U1870 ( .A(y[310]), .B(n3879), .Z(n3880) );
  XOR U1871 ( .A(y[314]), .B(n3863), .Z(n3864) );
  XOR U1872 ( .A(y[318]), .B(n3847), .Z(n3848) );
  XOR U1873 ( .A(y[322]), .B(n3831), .Z(n3832) );
  XOR U1874 ( .A(y[326]), .B(n3815), .Z(n3816) );
  XOR U1875 ( .A(y[330]), .B(n3799), .Z(n3800) );
  XOR U1876 ( .A(y[334]), .B(n3783), .Z(n3784) );
  XOR U1877 ( .A(y[338]), .B(n3767), .Z(n3768) );
  XOR U1878 ( .A(y[342]), .B(n3751), .Z(n3752) );
  XOR U1879 ( .A(y[346]), .B(n3735), .Z(n3736) );
  XOR U1880 ( .A(y[350]), .B(n3719), .Z(n3720) );
  XOR U1881 ( .A(y[354]), .B(n3703), .Z(n3704) );
  XOR U1882 ( .A(y[358]), .B(n3687), .Z(n3688) );
  XOR U1883 ( .A(y[362]), .B(n3671), .Z(n3672) );
  XOR U1884 ( .A(y[366]), .B(n3655), .Z(n3656) );
  XOR U1885 ( .A(y[370]), .B(n3639), .Z(n3640) );
  XOR U1886 ( .A(y[374]), .B(n3623), .Z(n3624) );
  XOR U1887 ( .A(y[378]), .B(n3607), .Z(n3608) );
  XOR U1888 ( .A(y[382]), .B(n3591), .Z(n3592) );
  XOR U1889 ( .A(y[386]), .B(n3575), .Z(n3576) );
  XOR U1890 ( .A(y[390]), .B(n3559), .Z(n3560) );
  XOR U1891 ( .A(y[394]), .B(n3543), .Z(n3544) );
  XOR U1892 ( .A(y[398]), .B(n3527), .Z(n3528) );
  XOR U1893 ( .A(y[402]), .B(n3511), .Z(n3512) );
  XOR U1894 ( .A(y[406]), .B(n3495), .Z(n3496) );
  XOR U1895 ( .A(y[410]), .B(n3479), .Z(n3480) );
  XOR U1896 ( .A(y[414]), .B(n3463), .Z(n3464) );
  XOR U1897 ( .A(y[418]), .B(n3447), .Z(n3448) );
  XOR U1898 ( .A(y[422]), .B(n3431), .Z(n3432) );
  XOR U1899 ( .A(y[426]), .B(n3415), .Z(n3416) );
  XOR U1900 ( .A(y[430]), .B(n3399), .Z(n3400) );
  XOR U1901 ( .A(y[434]), .B(n3383), .Z(n3384) );
  XOR U1902 ( .A(y[438]), .B(n3367), .Z(n3368) );
  XOR U1903 ( .A(y[442]), .B(n3351), .Z(n3352) );
  XOR U1904 ( .A(y[446]), .B(n3335), .Z(n3336) );
  XOR U1905 ( .A(y[450]), .B(n3319), .Z(n3320) );
  XOR U1906 ( .A(y[454]), .B(n3303), .Z(n3304) );
  XOR U1907 ( .A(y[458]), .B(n3287), .Z(n3288) );
  XOR U1908 ( .A(y[462]), .B(n3271), .Z(n3272) );
  XOR U1909 ( .A(y[466]), .B(n3255), .Z(n3256) );
  XOR U1910 ( .A(y[470]), .B(n3239), .Z(n3240) );
  XOR U1911 ( .A(y[474]), .B(n3223), .Z(n3224) );
  XOR U1912 ( .A(y[478]), .B(n3207), .Z(n3208) );
  XOR U1913 ( .A(y[482]), .B(n3191), .Z(n3192) );
  XOR U1914 ( .A(y[486]), .B(n3175), .Z(n3176) );
  XOR U1915 ( .A(y[490]), .B(n3159), .Z(n3160) );
  XOR U1916 ( .A(y[494]), .B(n3143), .Z(n3144) );
  XOR U1917 ( .A(y[498]), .B(n3127), .Z(n3128) );
  XOR U1918 ( .A(y[502]), .B(n3111), .Z(n3112) );
  XOR U1919 ( .A(y[506]), .B(n3095), .Z(n3096) );
  XOR U1920 ( .A(y[510]), .B(n3079), .Z(n3080) );
  XOR U1921 ( .A(y[514]), .B(n3063), .Z(n3064) );
  XOR U1922 ( .A(y[518]), .B(n3047), .Z(n3048) );
  XOR U1923 ( .A(y[522]), .B(n3031), .Z(n3032) );
  XOR U1924 ( .A(y[526]), .B(n3015), .Z(n3016) );
  XOR U1925 ( .A(y[530]), .B(n2999), .Z(n3000) );
  XOR U1926 ( .A(y[534]), .B(n2983), .Z(n2984) );
  XOR U1927 ( .A(y[538]), .B(n2967), .Z(n2968) );
  XOR U1928 ( .A(y[542]), .B(n2951), .Z(n2952) );
  XOR U1929 ( .A(y[546]), .B(n2935), .Z(n2936) );
  XOR U1930 ( .A(y[550]), .B(n2919), .Z(n2920) );
  XOR U1931 ( .A(y[554]), .B(n2903), .Z(n2904) );
  XOR U1932 ( .A(y[558]), .B(n2887), .Z(n2888) );
  XOR U1933 ( .A(y[562]), .B(n2871), .Z(n2872) );
  XOR U1934 ( .A(y[566]), .B(n2855), .Z(n2856) );
  XOR U1935 ( .A(y[570]), .B(n2839), .Z(n2840) );
  XOR U1936 ( .A(y[574]), .B(n2823), .Z(n2824) );
  XOR U1937 ( .A(y[578]), .B(n2807), .Z(n2808) );
  XOR U1938 ( .A(y[582]), .B(n2791), .Z(n2792) );
  XOR U1939 ( .A(y[586]), .B(n2775), .Z(n2776) );
  XOR U1940 ( .A(y[590]), .B(n2759), .Z(n2760) );
  XOR U1941 ( .A(y[594]), .B(n2743), .Z(n2744) );
  XOR U1942 ( .A(y[598]), .B(n2727), .Z(n2728) );
  XOR U1943 ( .A(y[602]), .B(n2711), .Z(n2712) );
  XOR U1944 ( .A(y[606]), .B(n2695), .Z(n2696) );
  XOR U1945 ( .A(y[610]), .B(n2679), .Z(n2680) );
  XOR U1946 ( .A(y[614]), .B(n2663), .Z(n2664) );
  XOR U1947 ( .A(y[618]), .B(n2647), .Z(n2648) );
  XOR U1948 ( .A(y[622]), .B(n2631), .Z(n2632) );
  XOR U1949 ( .A(y[626]), .B(n2615), .Z(n2616) );
  XOR U1950 ( .A(y[630]), .B(n2599), .Z(n2600) );
  XOR U1951 ( .A(y[634]), .B(n2583), .Z(n2584) );
  XOR U1952 ( .A(y[638]), .B(n2567), .Z(n2568) );
  XOR U1953 ( .A(y[642]), .B(n2551), .Z(n2552) );
  XOR U1954 ( .A(y[646]), .B(n2535), .Z(n2536) );
  XOR U1955 ( .A(y[650]), .B(n2519), .Z(n2520) );
  XOR U1956 ( .A(y[654]), .B(n2503), .Z(n2504) );
  XOR U1957 ( .A(y[658]), .B(n2487), .Z(n2488) );
  XOR U1958 ( .A(y[662]), .B(n2471), .Z(n2472) );
  XOR U1959 ( .A(y[666]), .B(n2455), .Z(n2456) );
  XOR U1960 ( .A(y[670]), .B(n2439), .Z(n2440) );
  XOR U1961 ( .A(y[674]), .B(n2423), .Z(n2424) );
  XOR U1962 ( .A(y[678]), .B(n2407), .Z(n2408) );
  XOR U1963 ( .A(y[682]), .B(n2391), .Z(n2392) );
  XOR U1964 ( .A(y[686]), .B(n2375), .Z(n2376) );
  XOR U1965 ( .A(y[690]), .B(n2359), .Z(n2360) );
  XOR U1966 ( .A(y[694]), .B(n2343), .Z(n2344) );
  XOR U1967 ( .A(y[698]), .B(n2327), .Z(n2328) );
  XOR U1968 ( .A(y[702]), .B(n2311), .Z(n2312) );
  XOR U1969 ( .A(y[706]), .B(n2295), .Z(n2296) );
  XOR U1970 ( .A(y[710]), .B(n2279), .Z(n2280) );
  XOR U1971 ( .A(y[714]), .B(n2263), .Z(n2264) );
  XOR U1972 ( .A(y[718]), .B(n2247), .Z(n2248) );
  XOR U1973 ( .A(y[722]), .B(n2231), .Z(n2232) );
  XOR U1974 ( .A(y[726]), .B(n2215), .Z(n2216) );
  XOR U1975 ( .A(y[730]), .B(n2199), .Z(n2200) );
  XOR U1976 ( .A(y[734]), .B(n2183), .Z(n2184) );
  XOR U1977 ( .A(y[738]), .B(n2167), .Z(n2168) );
  XOR U1978 ( .A(y[742]), .B(n2151), .Z(n2152) );
  XOR U1979 ( .A(y[746]), .B(n2135), .Z(n2136) );
  XOR U1980 ( .A(y[750]), .B(n2119), .Z(n2120) );
  XOR U1981 ( .A(y[754]), .B(n2103), .Z(n2104) );
  XOR U1982 ( .A(y[758]), .B(n2087), .Z(n2088) );
  XOR U1983 ( .A(y[762]), .B(n2071), .Z(n2072) );
  XOR U1984 ( .A(y[766]), .B(n2055), .Z(n2056) );
  XOR U1985 ( .A(y[770]), .B(n2039), .Z(n2040) );
  XOR U1986 ( .A(y[774]), .B(n2023), .Z(n2024) );
  XOR U1987 ( .A(y[778]), .B(n2007), .Z(n2008) );
  XOR U1988 ( .A(y[782]), .B(n1991), .Z(n1992) );
  XOR U1989 ( .A(y[786]), .B(n1975), .Z(n1976) );
  XOR U1990 ( .A(y[790]), .B(n1959), .Z(n1960) );
  XOR U1991 ( .A(y[794]), .B(n1943), .Z(n1944) );
  XOR U1992 ( .A(y[798]), .B(n1927), .Z(n1928) );
  XOR U1993 ( .A(y[802]), .B(n1911), .Z(n1912) );
  XOR U1994 ( .A(y[806]), .B(n1895), .Z(n1896) );
  XOR U1995 ( .A(y[810]), .B(n1879), .Z(n1880) );
  XOR U1996 ( .A(y[814]), .B(n1863), .Z(n1864) );
  XOR U1997 ( .A(y[818]), .B(n1847), .Z(n1848) );
  XOR U1998 ( .A(y[822]), .B(n1831), .Z(n1832) );
  XOR U1999 ( .A(y[826]), .B(n1815), .Z(n1816) );
  XOR U2000 ( .A(y[830]), .B(n1799), .Z(n1800) );
  XOR U2001 ( .A(y[834]), .B(n1783), .Z(n1784) );
  XOR U2002 ( .A(y[838]), .B(n1767), .Z(n1768) );
  XOR U2003 ( .A(y[842]), .B(n1751), .Z(n1752) );
  XOR U2004 ( .A(y[846]), .B(n1735), .Z(n1736) );
  XOR U2005 ( .A(y[850]), .B(n1719), .Z(n1720) );
  XOR U2006 ( .A(y[854]), .B(n1703), .Z(n1704) );
  XOR U2007 ( .A(y[858]), .B(n1687), .Z(n1688) );
  XOR U2008 ( .A(y[862]), .B(n1671), .Z(n1672) );
  XOR U2009 ( .A(y[866]), .B(n1655), .Z(n1656) );
  XOR U2010 ( .A(y[870]), .B(n1639), .Z(n1640) );
  XOR U2011 ( .A(y[874]), .B(n1623), .Z(n1624) );
  XOR U2012 ( .A(y[878]), .B(n1607), .Z(n1608) );
  XOR U2013 ( .A(y[882]), .B(n1591), .Z(n1592) );
  XOR U2014 ( .A(y[886]), .B(n1575), .Z(n1576) );
  XOR U2015 ( .A(y[890]), .B(n1559), .Z(n1560) );
  XOR U2016 ( .A(y[894]), .B(n1543), .Z(n1544) );
  XOR U2017 ( .A(y[898]), .B(n1527), .Z(n1528) );
  XOR U2018 ( .A(y[902]), .B(n1511), .Z(n1512) );
  XOR U2019 ( .A(y[906]), .B(n1495), .Z(n1496) );
  XOR U2020 ( .A(y[910]), .B(n1479), .Z(n1480) );
  XOR U2021 ( .A(y[914]), .B(n1463), .Z(n1464) );
  XOR U2022 ( .A(y[918]), .B(n1447), .Z(n1448) );
  XOR U2023 ( .A(y[922]), .B(n1431), .Z(n1432) );
  XOR U2024 ( .A(y[926]), .B(n1415), .Z(n1416) );
  XOR U2025 ( .A(y[930]), .B(n1399), .Z(n1400) );
  XOR U2026 ( .A(y[934]), .B(n1383), .Z(n1384) );
  XOR U2027 ( .A(y[938]), .B(n1367), .Z(n1368) );
  XOR U2028 ( .A(y[942]), .B(n1351), .Z(n1352) );
  XOR U2029 ( .A(y[946]), .B(n1335), .Z(n1336) );
  XOR U2030 ( .A(y[950]), .B(n1319), .Z(n1320) );
  XOR U2031 ( .A(y[954]), .B(n1303), .Z(n1304) );
  XOR U2032 ( .A(y[958]), .B(n1287), .Z(n1288) );
  XOR U2033 ( .A(y[962]), .B(n1271), .Z(n1272) );
  XOR U2034 ( .A(y[966]), .B(n1255), .Z(n1256) );
  XOR U2035 ( .A(y[970]), .B(n1239), .Z(n1240) );
  XOR U2036 ( .A(y[974]), .B(n1223), .Z(n1224) );
  XOR U2037 ( .A(y[978]), .B(n1207), .Z(n1208) );
  XOR U2038 ( .A(y[982]), .B(n1191), .Z(n1192) );
  XOR U2039 ( .A(y[986]), .B(n1175), .Z(n1176) );
  XOR U2040 ( .A(y[990]), .B(n1159), .Z(n1160) );
  XOR U2041 ( .A(y[994]), .B(n1143), .Z(n1144) );
  XOR U2042 ( .A(y[998]), .B(n1127), .Z(n1128) );
  XOR U2043 ( .A(y[1002]), .B(n1111), .Z(n1112) );
  XOR U2044 ( .A(y[1006]), .B(n1095), .Z(n1096) );
  XOR U2045 ( .A(y[1010]), .B(n1079), .Z(n1080) );
  XOR U2046 ( .A(y[1014]), .B(n1063), .Z(n1064) );
  XOR U2047 ( .A(y[1018]), .B(n1047), .Z(n1048) );
  XOR U2048 ( .A(y[1022]), .B(n1031), .Z(n1032) );
  XOR U2049 ( .A(n1026), .B(n1027), .Z(g) );
  AND U2050 ( .A(n1028), .B(n1029), .Z(n1026) );
  XOR U2051 ( .A(x[1023]), .B(n1027), .Z(n1029) );
  XNOR U2052 ( .A(y[1023]), .B(n1027), .Z(n1028) );
  XNOR U2053 ( .A(n1030), .B(n1031), .Z(n1027) );
  AND U2054 ( .A(n1032), .B(n1033), .Z(n1030) );
  XNOR U2055 ( .A(x[1022]), .B(n1031), .Z(n1033) );
  XOR U2056 ( .A(n1034), .B(n1035), .Z(n1031) );
  AND U2057 ( .A(n1036), .B(n1037), .Z(n1034) );
  XNOR U2058 ( .A(x[1021]), .B(n1035), .Z(n1037) );
  XOR U2059 ( .A(n1038), .B(n1039), .Z(n1035) );
  AND U2060 ( .A(n1040), .B(n1041), .Z(n1038) );
  XNOR U2061 ( .A(x[1020]), .B(n1039), .Z(n1041) );
  XOR U2062 ( .A(n1042), .B(n1043), .Z(n1039) );
  AND U2063 ( .A(n1044), .B(n1045), .Z(n1042) );
  XNOR U2064 ( .A(x[1019]), .B(n1043), .Z(n1045) );
  XOR U2065 ( .A(n1046), .B(n1047), .Z(n1043) );
  AND U2066 ( .A(n1048), .B(n1049), .Z(n1046) );
  XNOR U2067 ( .A(x[1018]), .B(n1047), .Z(n1049) );
  XOR U2068 ( .A(n1050), .B(n1051), .Z(n1047) );
  AND U2069 ( .A(n1052), .B(n1053), .Z(n1050) );
  XNOR U2070 ( .A(x[1017]), .B(n1051), .Z(n1053) );
  XOR U2071 ( .A(n1054), .B(n1055), .Z(n1051) );
  AND U2072 ( .A(n1056), .B(n1057), .Z(n1054) );
  XNOR U2073 ( .A(x[1016]), .B(n1055), .Z(n1057) );
  XOR U2074 ( .A(n1058), .B(n1059), .Z(n1055) );
  AND U2075 ( .A(n1060), .B(n1061), .Z(n1058) );
  XNOR U2076 ( .A(x[1015]), .B(n1059), .Z(n1061) );
  XOR U2077 ( .A(n1062), .B(n1063), .Z(n1059) );
  AND U2078 ( .A(n1064), .B(n1065), .Z(n1062) );
  XNOR U2079 ( .A(x[1014]), .B(n1063), .Z(n1065) );
  XOR U2080 ( .A(n1066), .B(n1067), .Z(n1063) );
  AND U2081 ( .A(n1068), .B(n1069), .Z(n1066) );
  XNOR U2082 ( .A(x[1013]), .B(n1067), .Z(n1069) );
  XOR U2083 ( .A(n1070), .B(n1071), .Z(n1067) );
  AND U2084 ( .A(n1072), .B(n1073), .Z(n1070) );
  XNOR U2085 ( .A(x[1012]), .B(n1071), .Z(n1073) );
  XOR U2086 ( .A(n1074), .B(n1075), .Z(n1071) );
  AND U2087 ( .A(n1076), .B(n1077), .Z(n1074) );
  XNOR U2088 ( .A(x[1011]), .B(n1075), .Z(n1077) );
  XOR U2089 ( .A(n1078), .B(n1079), .Z(n1075) );
  AND U2090 ( .A(n1080), .B(n1081), .Z(n1078) );
  XNOR U2091 ( .A(x[1010]), .B(n1079), .Z(n1081) );
  XOR U2092 ( .A(n1082), .B(n1083), .Z(n1079) );
  AND U2093 ( .A(n1084), .B(n1085), .Z(n1082) );
  XNOR U2094 ( .A(x[1009]), .B(n1083), .Z(n1085) );
  XOR U2095 ( .A(n1086), .B(n1087), .Z(n1083) );
  AND U2096 ( .A(n1088), .B(n1089), .Z(n1086) );
  XNOR U2097 ( .A(x[1008]), .B(n1087), .Z(n1089) );
  XOR U2098 ( .A(n1090), .B(n1091), .Z(n1087) );
  AND U2099 ( .A(n1092), .B(n1093), .Z(n1090) );
  XNOR U2100 ( .A(x[1007]), .B(n1091), .Z(n1093) );
  XOR U2101 ( .A(n1094), .B(n1095), .Z(n1091) );
  AND U2102 ( .A(n1096), .B(n1097), .Z(n1094) );
  XNOR U2103 ( .A(x[1006]), .B(n1095), .Z(n1097) );
  XOR U2104 ( .A(n1098), .B(n1099), .Z(n1095) );
  AND U2105 ( .A(n1100), .B(n1101), .Z(n1098) );
  XNOR U2106 ( .A(x[1005]), .B(n1099), .Z(n1101) );
  XOR U2107 ( .A(n1102), .B(n1103), .Z(n1099) );
  AND U2108 ( .A(n1104), .B(n1105), .Z(n1102) );
  XNOR U2109 ( .A(x[1004]), .B(n1103), .Z(n1105) );
  XOR U2110 ( .A(n1106), .B(n1107), .Z(n1103) );
  AND U2111 ( .A(n1108), .B(n1109), .Z(n1106) );
  XNOR U2112 ( .A(x[1003]), .B(n1107), .Z(n1109) );
  XOR U2113 ( .A(n1110), .B(n1111), .Z(n1107) );
  AND U2114 ( .A(n1112), .B(n1113), .Z(n1110) );
  XNOR U2115 ( .A(x[1002]), .B(n1111), .Z(n1113) );
  XOR U2116 ( .A(n1114), .B(n1115), .Z(n1111) );
  AND U2117 ( .A(n1116), .B(n1117), .Z(n1114) );
  XNOR U2118 ( .A(x[1001]), .B(n1115), .Z(n1117) );
  XOR U2119 ( .A(n1118), .B(n1119), .Z(n1115) );
  AND U2120 ( .A(n1120), .B(n1121), .Z(n1118) );
  XNOR U2121 ( .A(x[1000]), .B(n1119), .Z(n1121) );
  XOR U2122 ( .A(n1122), .B(n1123), .Z(n1119) );
  AND U2123 ( .A(n1124), .B(n1125), .Z(n1122) );
  XNOR U2124 ( .A(x[999]), .B(n1123), .Z(n1125) );
  XOR U2125 ( .A(n1126), .B(n1127), .Z(n1123) );
  AND U2126 ( .A(n1128), .B(n1129), .Z(n1126) );
  XNOR U2127 ( .A(x[998]), .B(n1127), .Z(n1129) );
  XOR U2128 ( .A(n1130), .B(n1131), .Z(n1127) );
  AND U2129 ( .A(n1132), .B(n1133), .Z(n1130) );
  XNOR U2130 ( .A(x[997]), .B(n1131), .Z(n1133) );
  XOR U2131 ( .A(n1134), .B(n1135), .Z(n1131) );
  AND U2132 ( .A(n1136), .B(n1137), .Z(n1134) );
  XNOR U2133 ( .A(x[996]), .B(n1135), .Z(n1137) );
  XOR U2134 ( .A(n1138), .B(n1139), .Z(n1135) );
  AND U2135 ( .A(n1140), .B(n1141), .Z(n1138) );
  XNOR U2136 ( .A(x[995]), .B(n1139), .Z(n1141) );
  XOR U2137 ( .A(n1142), .B(n1143), .Z(n1139) );
  AND U2138 ( .A(n1144), .B(n1145), .Z(n1142) );
  XNOR U2139 ( .A(x[994]), .B(n1143), .Z(n1145) );
  XOR U2140 ( .A(n1146), .B(n1147), .Z(n1143) );
  AND U2141 ( .A(n1148), .B(n1149), .Z(n1146) );
  XNOR U2142 ( .A(x[993]), .B(n1147), .Z(n1149) );
  XOR U2143 ( .A(n1150), .B(n1151), .Z(n1147) );
  AND U2144 ( .A(n1152), .B(n1153), .Z(n1150) );
  XNOR U2145 ( .A(x[992]), .B(n1151), .Z(n1153) );
  XOR U2146 ( .A(n1154), .B(n1155), .Z(n1151) );
  AND U2147 ( .A(n1156), .B(n1157), .Z(n1154) );
  XNOR U2148 ( .A(x[991]), .B(n1155), .Z(n1157) );
  XOR U2149 ( .A(n1158), .B(n1159), .Z(n1155) );
  AND U2150 ( .A(n1160), .B(n1161), .Z(n1158) );
  XNOR U2151 ( .A(x[990]), .B(n1159), .Z(n1161) );
  XOR U2152 ( .A(n1162), .B(n1163), .Z(n1159) );
  AND U2153 ( .A(n1164), .B(n1165), .Z(n1162) );
  XNOR U2154 ( .A(x[989]), .B(n1163), .Z(n1165) );
  XOR U2155 ( .A(n1166), .B(n1167), .Z(n1163) );
  AND U2156 ( .A(n1168), .B(n1169), .Z(n1166) );
  XNOR U2157 ( .A(x[988]), .B(n1167), .Z(n1169) );
  XOR U2158 ( .A(n1170), .B(n1171), .Z(n1167) );
  AND U2159 ( .A(n1172), .B(n1173), .Z(n1170) );
  XNOR U2160 ( .A(x[987]), .B(n1171), .Z(n1173) );
  XOR U2161 ( .A(n1174), .B(n1175), .Z(n1171) );
  AND U2162 ( .A(n1176), .B(n1177), .Z(n1174) );
  XNOR U2163 ( .A(x[986]), .B(n1175), .Z(n1177) );
  XOR U2164 ( .A(n1178), .B(n1179), .Z(n1175) );
  AND U2165 ( .A(n1180), .B(n1181), .Z(n1178) );
  XNOR U2166 ( .A(x[985]), .B(n1179), .Z(n1181) );
  XOR U2167 ( .A(n1182), .B(n1183), .Z(n1179) );
  AND U2168 ( .A(n1184), .B(n1185), .Z(n1182) );
  XNOR U2169 ( .A(x[984]), .B(n1183), .Z(n1185) );
  XOR U2170 ( .A(n1186), .B(n1187), .Z(n1183) );
  AND U2171 ( .A(n1188), .B(n1189), .Z(n1186) );
  XNOR U2172 ( .A(x[983]), .B(n1187), .Z(n1189) );
  XOR U2173 ( .A(n1190), .B(n1191), .Z(n1187) );
  AND U2174 ( .A(n1192), .B(n1193), .Z(n1190) );
  XNOR U2175 ( .A(x[982]), .B(n1191), .Z(n1193) );
  XOR U2176 ( .A(n1194), .B(n1195), .Z(n1191) );
  AND U2177 ( .A(n1196), .B(n1197), .Z(n1194) );
  XNOR U2178 ( .A(x[981]), .B(n1195), .Z(n1197) );
  XOR U2179 ( .A(n1198), .B(n1199), .Z(n1195) );
  AND U2180 ( .A(n1200), .B(n1201), .Z(n1198) );
  XNOR U2181 ( .A(x[980]), .B(n1199), .Z(n1201) );
  XOR U2182 ( .A(n1202), .B(n1203), .Z(n1199) );
  AND U2183 ( .A(n1204), .B(n1205), .Z(n1202) );
  XNOR U2184 ( .A(x[979]), .B(n1203), .Z(n1205) );
  XOR U2185 ( .A(n1206), .B(n1207), .Z(n1203) );
  AND U2186 ( .A(n1208), .B(n1209), .Z(n1206) );
  XNOR U2187 ( .A(x[978]), .B(n1207), .Z(n1209) );
  XOR U2188 ( .A(n1210), .B(n1211), .Z(n1207) );
  AND U2189 ( .A(n1212), .B(n1213), .Z(n1210) );
  XNOR U2190 ( .A(x[977]), .B(n1211), .Z(n1213) );
  XOR U2191 ( .A(n1214), .B(n1215), .Z(n1211) );
  AND U2192 ( .A(n1216), .B(n1217), .Z(n1214) );
  XNOR U2193 ( .A(x[976]), .B(n1215), .Z(n1217) );
  XOR U2194 ( .A(n1218), .B(n1219), .Z(n1215) );
  AND U2195 ( .A(n1220), .B(n1221), .Z(n1218) );
  XNOR U2196 ( .A(x[975]), .B(n1219), .Z(n1221) );
  XOR U2197 ( .A(n1222), .B(n1223), .Z(n1219) );
  AND U2198 ( .A(n1224), .B(n1225), .Z(n1222) );
  XNOR U2199 ( .A(x[974]), .B(n1223), .Z(n1225) );
  XOR U2200 ( .A(n1226), .B(n1227), .Z(n1223) );
  AND U2201 ( .A(n1228), .B(n1229), .Z(n1226) );
  XNOR U2202 ( .A(x[973]), .B(n1227), .Z(n1229) );
  XOR U2203 ( .A(n1230), .B(n1231), .Z(n1227) );
  AND U2204 ( .A(n1232), .B(n1233), .Z(n1230) );
  XNOR U2205 ( .A(x[972]), .B(n1231), .Z(n1233) );
  XOR U2206 ( .A(n1234), .B(n1235), .Z(n1231) );
  AND U2207 ( .A(n1236), .B(n1237), .Z(n1234) );
  XNOR U2208 ( .A(x[971]), .B(n1235), .Z(n1237) );
  XOR U2209 ( .A(n1238), .B(n1239), .Z(n1235) );
  AND U2210 ( .A(n1240), .B(n1241), .Z(n1238) );
  XNOR U2211 ( .A(x[970]), .B(n1239), .Z(n1241) );
  XOR U2212 ( .A(n1242), .B(n1243), .Z(n1239) );
  AND U2213 ( .A(n1244), .B(n1245), .Z(n1242) );
  XNOR U2214 ( .A(x[969]), .B(n1243), .Z(n1245) );
  XOR U2215 ( .A(n1246), .B(n1247), .Z(n1243) );
  AND U2216 ( .A(n1248), .B(n1249), .Z(n1246) );
  XNOR U2217 ( .A(x[968]), .B(n1247), .Z(n1249) );
  XOR U2218 ( .A(n1250), .B(n1251), .Z(n1247) );
  AND U2219 ( .A(n1252), .B(n1253), .Z(n1250) );
  XNOR U2220 ( .A(x[967]), .B(n1251), .Z(n1253) );
  XOR U2221 ( .A(n1254), .B(n1255), .Z(n1251) );
  AND U2222 ( .A(n1256), .B(n1257), .Z(n1254) );
  XNOR U2223 ( .A(x[966]), .B(n1255), .Z(n1257) );
  XOR U2224 ( .A(n1258), .B(n1259), .Z(n1255) );
  AND U2225 ( .A(n1260), .B(n1261), .Z(n1258) );
  XNOR U2226 ( .A(x[965]), .B(n1259), .Z(n1261) );
  XOR U2227 ( .A(n1262), .B(n1263), .Z(n1259) );
  AND U2228 ( .A(n1264), .B(n1265), .Z(n1262) );
  XNOR U2229 ( .A(x[964]), .B(n1263), .Z(n1265) );
  XOR U2230 ( .A(n1266), .B(n1267), .Z(n1263) );
  AND U2231 ( .A(n1268), .B(n1269), .Z(n1266) );
  XNOR U2232 ( .A(x[963]), .B(n1267), .Z(n1269) );
  XOR U2233 ( .A(n1270), .B(n1271), .Z(n1267) );
  AND U2234 ( .A(n1272), .B(n1273), .Z(n1270) );
  XNOR U2235 ( .A(x[962]), .B(n1271), .Z(n1273) );
  XOR U2236 ( .A(n1274), .B(n1275), .Z(n1271) );
  AND U2237 ( .A(n1276), .B(n1277), .Z(n1274) );
  XNOR U2238 ( .A(x[961]), .B(n1275), .Z(n1277) );
  XOR U2239 ( .A(n1278), .B(n1279), .Z(n1275) );
  AND U2240 ( .A(n1280), .B(n1281), .Z(n1278) );
  XNOR U2241 ( .A(x[960]), .B(n1279), .Z(n1281) );
  XOR U2242 ( .A(n1282), .B(n1283), .Z(n1279) );
  AND U2243 ( .A(n1284), .B(n1285), .Z(n1282) );
  XNOR U2244 ( .A(x[959]), .B(n1283), .Z(n1285) );
  XOR U2245 ( .A(n1286), .B(n1287), .Z(n1283) );
  AND U2246 ( .A(n1288), .B(n1289), .Z(n1286) );
  XNOR U2247 ( .A(x[958]), .B(n1287), .Z(n1289) );
  XOR U2248 ( .A(n1290), .B(n1291), .Z(n1287) );
  AND U2249 ( .A(n1292), .B(n1293), .Z(n1290) );
  XNOR U2250 ( .A(x[957]), .B(n1291), .Z(n1293) );
  XOR U2251 ( .A(n1294), .B(n1295), .Z(n1291) );
  AND U2252 ( .A(n1296), .B(n1297), .Z(n1294) );
  XNOR U2253 ( .A(x[956]), .B(n1295), .Z(n1297) );
  XOR U2254 ( .A(n1298), .B(n1299), .Z(n1295) );
  AND U2255 ( .A(n1300), .B(n1301), .Z(n1298) );
  XNOR U2256 ( .A(x[955]), .B(n1299), .Z(n1301) );
  XOR U2257 ( .A(n1302), .B(n1303), .Z(n1299) );
  AND U2258 ( .A(n1304), .B(n1305), .Z(n1302) );
  XNOR U2259 ( .A(x[954]), .B(n1303), .Z(n1305) );
  XOR U2260 ( .A(n1306), .B(n1307), .Z(n1303) );
  AND U2261 ( .A(n1308), .B(n1309), .Z(n1306) );
  XNOR U2262 ( .A(x[953]), .B(n1307), .Z(n1309) );
  XOR U2263 ( .A(n1310), .B(n1311), .Z(n1307) );
  AND U2264 ( .A(n1312), .B(n1313), .Z(n1310) );
  XNOR U2265 ( .A(x[952]), .B(n1311), .Z(n1313) );
  XOR U2266 ( .A(n1314), .B(n1315), .Z(n1311) );
  AND U2267 ( .A(n1316), .B(n1317), .Z(n1314) );
  XNOR U2268 ( .A(x[951]), .B(n1315), .Z(n1317) );
  XOR U2269 ( .A(n1318), .B(n1319), .Z(n1315) );
  AND U2270 ( .A(n1320), .B(n1321), .Z(n1318) );
  XNOR U2271 ( .A(x[950]), .B(n1319), .Z(n1321) );
  XOR U2272 ( .A(n1322), .B(n1323), .Z(n1319) );
  AND U2273 ( .A(n1324), .B(n1325), .Z(n1322) );
  XNOR U2274 ( .A(x[949]), .B(n1323), .Z(n1325) );
  XOR U2275 ( .A(n1326), .B(n1327), .Z(n1323) );
  AND U2276 ( .A(n1328), .B(n1329), .Z(n1326) );
  XNOR U2277 ( .A(x[948]), .B(n1327), .Z(n1329) );
  XOR U2278 ( .A(n1330), .B(n1331), .Z(n1327) );
  AND U2279 ( .A(n1332), .B(n1333), .Z(n1330) );
  XNOR U2280 ( .A(x[947]), .B(n1331), .Z(n1333) );
  XOR U2281 ( .A(n1334), .B(n1335), .Z(n1331) );
  AND U2282 ( .A(n1336), .B(n1337), .Z(n1334) );
  XNOR U2283 ( .A(x[946]), .B(n1335), .Z(n1337) );
  XOR U2284 ( .A(n1338), .B(n1339), .Z(n1335) );
  AND U2285 ( .A(n1340), .B(n1341), .Z(n1338) );
  XNOR U2286 ( .A(x[945]), .B(n1339), .Z(n1341) );
  XOR U2287 ( .A(n1342), .B(n1343), .Z(n1339) );
  AND U2288 ( .A(n1344), .B(n1345), .Z(n1342) );
  XNOR U2289 ( .A(x[944]), .B(n1343), .Z(n1345) );
  XOR U2290 ( .A(n1346), .B(n1347), .Z(n1343) );
  AND U2291 ( .A(n1348), .B(n1349), .Z(n1346) );
  XNOR U2292 ( .A(x[943]), .B(n1347), .Z(n1349) );
  XOR U2293 ( .A(n1350), .B(n1351), .Z(n1347) );
  AND U2294 ( .A(n1352), .B(n1353), .Z(n1350) );
  XNOR U2295 ( .A(x[942]), .B(n1351), .Z(n1353) );
  XOR U2296 ( .A(n1354), .B(n1355), .Z(n1351) );
  AND U2297 ( .A(n1356), .B(n1357), .Z(n1354) );
  XNOR U2298 ( .A(x[941]), .B(n1355), .Z(n1357) );
  XOR U2299 ( .A(n1358), .B(n1359), .Z(n1355) );
  AND U2300 ( .A(n1360), .B(n1361), .Z(n1358) );
  XNOR U2301 ( .A(x[940]), .B(n1359), .Z(n1361) );
  XOR U2302 ( .A(n1362), .B(n1363), .Z(n1359) );
  AND U2303 ( .A(n1364), .B(n1365), .Z(n1362) );
  XNOR U2304 ( .A(x[939]), .B(n1363), .Z(n1365) );
  XOR U2305 ( .A(n1366), .B(n1367), .Z(n1363) );
  AND U2306 ( .A(n1368), .B(n1369), .Z(n1366) );
  XNOR U2307 ( .A(x[938]), .B(n1367), .Z(n1369) );
  XOR U2308 ( .A(n1370), .B(n1371), .Z(n1367) );
  AND U2309 ( .A(n1372), .B(n1373), .Z(n1370) );
  XNOR U2310 ( .A(x[937]), .B(n1371), .Z(n1373) );
  XOR U2311 ( .A(n1374), .B(n1375), .Z(n1371) );
  AND U2312 ( .A(n1376), .B(n1377), .Z(n1374) );
  XNOR U2313 ( .A(x[936]), .B(n1375), .Z(n1377) );
  XOR U2314 ( .A(n1378), .B(n1379), .Z(n1375) );
  AND U2315 ( .A(n1380), .B(n1381), .Z(n1378) );
  XNOR U2316 ( .A(x[935]), .B(n1379), .Z(n1381) );
  XOR U2317 ( .A(n1382), .B(n1383), .Z(n1379) );
  AND U2318 ( .A(n1384), .B(n1385), .Z(n1382) );
  XNOR U2319 ( .A(x[934]), .B(n1383), .Z(n1385) );
  XOR U2320 ( .A(n1386), .B(n1387), .Z(n1383) );
  AND U2321 ( .A(n1388), .B(n1389), .Z(n1386) );
  XNOR U2322 ( .A(x[933]), .B(n1387), .Z(n1389) );
  XOR U2323 ( .A(n1390), .B(n1391), .Z(n1387) );
  AND U2324 ( .A(n1392), .B(n1393), .Z(n1390) );
  XNOR U2325 ( .A(x[932]), .B(n1391), .Z(n1393) );
  XOR U2326 ( .A(n1394), .B(n1395), .Z(n1391) );
  AND U2327 ( .A(n1396), .B(n1397), .Z(n1394) );
  XNOR U2328 ( .A(x[931]), .B(n1395), .Z(n1397) );
  XOR U2329 ( .A(n1398), .B(n1399), .Z(n1395) );
  AND U2330 ( .A(n1400), .B(n1401), .Z(n1398) );
  XNOR U2331 ( .A(x[930]), .B(n1399), .Z(n1401) );
  XOR U2332 ( .A(n1402), .B(n1403), .Z(n1399) );
  AND U2333 ( .A(n1404), .B(n1405), .Z(n1402) );
  XNOR U2334 ( .A(x[929]), .B(n1403), .Z(n1405) );
  XOR U2335 ( .A(n1406), .B(n1407), .Z(n1403) );
  AND U2336 ( .A(n1408), .B(n1409), .Z(n1406) );
  XNOR U2337 ( .A(x[928]), .B(n1407), .Z(n1409) );
  XOR U2338 ( .A(n1410), .B(n1411), .Z(n1407) );
  AND U2339 ( .A(n1412), .B(n1413), .Z(n1410) );
  XNOR U2340 ( .A(x[927]), .B(n1411), .Z(n1413) );
  XOR U2341 ( .A(n1414), .B(n1415), .Z(n1411) );
  AND U2342 ( .A(n1416), .B(n1417), .Z(n1414) );
  XNOR U2343 ( .A(x[926]), .B(n1415), .Z(n1417) );
  XOR U2344 ( .A(n1418), .B(n1419), .Z(n1415) );
  AND U2345 ( .A(n1420), .B(n1421), .Z(n1418) );
  XNOR U2346 ( .A(x[925]), .B(n1419), .Z(n1421) );
  XOR U2347 ( .A(n1422), .B(n1423), .Z(n1419) );
  AND U2348 ( .A(n1424), .B(n1425), .Z(n1422) );
  XNOR U2349 ( .A(x[924]), .B(n1423), .Z(n1425) );
  XOR U2350 ( .A(n1426), .B(n1427), .Z(n1423) );
  AND U2351 ( .A(n1428), .B(n1429), .Z(n1426) );
  XNOR U2352 ( .A(x[923]), .B(n1427), .Z(n1429) );
  XOR U2353 ( .A(n1430), .B(n1431), .Z(n1427) );
  AND U2354 ( .A(n1432), .B(n1433), .Z(n1430) );
  XNOR U2355 ( .A(x[922]), .B(n1431), .Z(n1433) );
  XOR U2356 ( .A(n1434), .B(n1435), .Z(n1431) );
  AND U2357 ( .A(n1436), .B(n1437), .Z(n1434) );
  XNOR U2358 ( .A(x[921]), .B(n1435), .Z(n1437) );
  XOR U2359 ( .A(n1438), .B(n1439), .Z(n1435) );
  AND U2360 ( .A(n1440), .B(n1441), .Z(n1438) );
  XNOR U2361 ( .A(x[920]), .B(n1439), .Z(n1441) );
  XOR U2362 ( .A(n1442), .B(n1443), .Z(n1439) );
  AND U2363 ( .A(n1444), .B(n1445), .Z(n1442) );
  XNOR U2364 ( .A(x[919]), .B(n1443), .Z(n1445) );
  XOR U2365 ( .A(n1446), .B(n1447), .Z(n1443) );
  AND U2366 ( .A(n1448), .B(n1449), .Z(n1446) );
  XNOR U2367 ( .A(x[918]), .B(n1447), .Z(n1449) );
  XOR U2368 ( .A(n1450), .B(n1451), .Z(n1447) );
  AND U2369 ( .A(n1452), .B(n1453), .Z(n1450) );
  XNOR U2370 ( .A(x[917]), .B(n1451), .Z(n1453) );
  XOR U2371 ( .A(n1454), .B(n1455), .Z(n1451) );
  AND U2372 ( .A(n1456), .B(n1457), .Z(n1454) );
  XNOR U2373 ( .A(x[916]), .B(n1455), .Z(n1457) );
  XOR U2374 ( .A(n1458), .B(n1459), .Z(n1455) );
  AND U2375 ( .A(n1460), .B(n1461), .Z(n1458) );
  XNOR U2376 ( .A(x[915]), .B(n1459), .Z(n1461) );
  XOR U2377 ( .A(n1462), .B(n1463), .Z(n1459) );
  AND U2378 ( .A(n1464), .B(n1465), .Z(n1462) );
  XNOR U2379 ( .A(x[914]), .B(n1463), .Z(n1465) );
  XOR U2380 ( .A(n1466), .B(n1467), .Z(n1463) );
  AND U2381 ( .A(n1468), .B(n1469), .Z(n1466) );
  XNOR U2382 ( .A(x[913]), .B(n1467), .Z(n1469) );
  XOR U2383 ( .A(n1470), .B(n1471), .Z(n1467) );
  AND U2384 ( .A(n1472), .B(n1473), .Z(n1470) );
  XNOR U2385 ( .A(x[912]), .B(n1471), .Z(n1473) );
  XOR U2386 ( .A(n1474), .B(n1475), .Z(n1471) );
  AND U2387 ( .A(n1476), .B(n1477), .Z(n1474) );
  XNOR U2388 ( .A(x[911]), .B(n1475), .Z(n1477) );
  XOR U2389 ( .A(n1478), .B(n1479), .Z(n1475) );
  AND U2390 ( .A(n1480), .B(n1481), .Z(n1478) );
  XNOR U2391 ( .A(x[910]), .B(n1479), .Z(n1481) );
  XOR U2392 ( .A(n1482), .B(n1483), .Z(n1479) );
  AND U2393 ( .A(n1484), .B(n1485), .Z(n1482) );
  XNOR U2394 ( .A(x[909]), .B(n1483), .Z(n1485) );
  XOR U2395 ( .A(n1486), .B(n1487), .Z(n1483) );
  AND U2396 ( .A(n1488), .B(n1489), .Z(n1486) );
  XNOR U2397 ( .A(x[908]), .B(n1487), .Z(n1489) );
  XOR U2398 ( .A(n1490), .B(n1491), .Z(n1487) );
  AND U2399 ( .A(n1492), .B(n1493), .Z(n1490) );
  XNOR U2400 ( .A(x[907]), .B(n1491), .Z(n1493) );
  XOR U2401 ( .A(n1494), .B(n1495), .Z(n1491) );
  AND U2402 ( .A(n1496), .B(n1497), .Z(n1494) );
  XNOR U2403 ( .A(x[906]), .B(n1495), .Z(n1497) );
  XOR U2404 ( .A(n1498), .B(n1499), .Z(n1495) );
  AND U2405 ( .A(n1500), .B(n1501), .Z(n1498) );
  XNOR U2406 ( .A(x[905]), .B(n1499), .Z(n1501) );
  XOR U2407 ( .A(n1502), .B(n1503), .Z(n1499) );
  AND U2408 ( .A(n1504), .B(n1505), .Z(n1502) );
  XNOR U2409 ( .A(x[904]), .B(n1503), .Z(n1505) );
  XOR U2410 ( .A(n1506), .B(n1507), .Z(n1503) );
  AND U2411 ( .A(n1508), .B(n1509), .Z(n1506) );
  XNOR U2412 ( .A(x[903]), .B(n1507), .Z(n1509) );
  XOR U2413 ( .A(n1510), .B(n1511), .Z(n1507) );
  AND U2414 ( .A(n1512), .B(n1513), .Z(n1510) );
  XNOR U2415 ( .A(x[902]), .B(n1511), .Z(n1513) );
  XOR U2416 ( .A(n1514), .B(n1515), .Z(n1511) );
  AND U2417 ( .A(n1516), .B(n1517), .Z(n1514) );
  XNOR U2418 ( .A(x[901]), .B(n1515), .Z(n1517) );
  XOR U2419 ( .A(n1518), .B(n1519), .Z(n1515) );
  AND U2420 ( .A(n1520), .B(n1521), .Z(n1518) );
  XNOR U2421 ( .A(x[900]), .B(n1519), .Z(n1521) );
  XOR U2422 ( .A(n1522), .B(n1523), .Z(n1519) );
  AND U2423 ( .A(n1524), .B(n1525), .Z(n1522) );
  XNOR U2424 ( .A(x[899]), .B(n1523), .Z(n1525) );
  XOR U2425 ( .A(n1526), .B(n1527), .Z(n1523) );
  AND U2426 ( .A(n1528), .B(n1529), .Z(n1526) );
  XNOR U2427 ( .A(x[898]), .B(n1527), .Z(n1529) );
  XOR U2428 ( .A(n1530), .B(n1531), .Z(n1527) );
  AND U2429 ( .A(n1532), .B(n1533), .Z(n1530) );
  XNOR U2430 ( .A(x[897]), .B(n1531), .Z(n1533) );
  XOR U2431 ( .A(n1534), .B(n1535), .Z(n1531) );
  AND U2432 ( .A(n1536), .B(n1537), .Z(n1534) );
  XNOR U2433 ( .A(x[896]), .B(n1535), .Z(n1537) );
  XOR U2434 ( .A(n1538), .B(n1539), .Z(n1535) );
  AND U2435 ( .A(n1540), .B(n1541), .Z(n1538) );
  XNOR U2436 ( .A(x[895]), .B(n1539), .Z(n1541) );
  XOR U2437 ( .A(n1542), .B(n1543), .Z(n1539) );
  AND U2438 ( .A(n1544), .B(n1545), .Z(n1542) );
  XNOR U2439 ( .A(x[894]), .B(n1543), .Z(n1545) );
  XOR U2440 ( .A(n1546), .B(n1547), .Z(n1543) );
  AND U2441 ( .A(n1548), .B(n1549), .Z(n1546) );
  XNOR U2442 ( .A(x[893]), .B(n1547), .Z(n1549) );
  XOR U2443 ( .A(n1550), .B(n1551), .Z(n1547) );
  AND U2444 ( .A(n1552), .B(n1553), .Z(n1550) );
  XNOR U2445 ( .A(x[892]), .B(n1551), .Z(n1553) );
  XOR U2446 ( .A(n1554), .B(n1555), .Z(n1551) );
  AND U2447 ( .A(n1556), .B(n1557), .Z(n1554) );
  XNOR U2448 ( .A(x[891]), .B(n1555), .Z(n1557) );
  XOR U2449 ( .A(n1558), .B(n1559), .Z(n1555) );
  AND U2450 ( .A(n1560), .B(n1561), .Z(n1558) );
  XNOR U2451 ( .A(x[890]), .B(n1559), .Z(n1561) );
  XOR U2452 ( .A(n1562), .B(n1563), .Z(n1559) );
  AND U2453 ( .A(n1564), .B(n1565), .Z(n1562) );
  XNOR U2454 ( .A(x[889]), .B(n1563), .Z(n1565) );
  XOR U2455 ( .A(n1566), .B(n1567), .Z(n1563) );
  AND U2456 ( .A(n1568), .B(n1569), .Z(n1566) );
  XNOR U2457 ( .A(x[888]), .B(n1567), .Z(n1569) );
  XOR U2458 ( .A(n1570), .B(n1571), .Z(n1567) );
  AND U2459 ( .A(n1572), .B(n1573), .Z(n1570) );
  XNOR U2460 ( .A(x[887]), .B(n1571), .Z(n1573) );
  XOR U2461 ( .A(n1574), .B(n1575), .Z(n1571) );
  AND U2462 ( .A(n1576), .B(n1577), .Z(n1574) );
  XNOR U2463 ( .A(x[886]), .B(n1575), .Z(n1577) );
  XOR U2464 ( .A(n1578), .B(n1579), .Z(n1575) );
  AND U2465 ( .A(n1580), .B(n1581), .Z(n1578) );
  XNOR U2466 ( .A(x[885]), .B(n1579), .Z(n1581) );
  XOR U2467 ( .A(n1582), .B(n1583), .Z(n1579) );
  AND U2468 ( .A(n1584), .B(n1585), .Z(n1582) );
  XNOR U2469 ( .A(x[884]), .B(n1583), .Z(n1585) );
  XOR U2470 ( .A(n1586), .B(n1587), .Z(n1583) );
  AND U2471 ( .A(n1588), .B(n1589), .Z(n1586) );
  XNOR U2472 ( .A(x[883]), .B(n1587), .Z(n1589) );
  XOR U2473 ( .A(n1590), .B(n1591), .Z(n1587) );
  AND U2474 ( .A(n1592), .B(n1593), .Z(n1590) );
  XNOR U2475 ( .A(x[882]), .B(n1591), .Z(n1593) );
  XOR U2476 ( .A(n1594), .B(n1595), .Z(n1591) );
  AND U2477 ( .A(n1596), .B(n1597), .Z(n1594) );
  XNOR U2478 ( .A(x[881]), .B(n1595), .Z(n1597) );
  XOR U2479 ( .A(n1598), .B(n1599), .Z(n1595) );
  AND U2480 ( .A(n1600), .B(n1601), .Z(n1598) );
  XNOR U2481 ( .A(x[880]), .B(n1599), .Z(n1601) );
  XOR U2482 ( .A(n1602), .B(n1603), .Z(n1599) );
  AND U2483 ( .A(n1604), .B(n1605), .Z(n1602) );
  XNOR U2484 ( .A(x[879]), .B(n1603), .Z(n1605) );
  XOR U2485 ( .A(n1606), .B(n1607), .Z(n1603) );
  AND U2486 ( .A(n1608), .B(n1609), .Z(n1606) );
  XNOR U2487 ( .A(x[878]), .B(n1607), .Z(n1609) );
  XOR U2488 ( .A(n1610), .B(n1611), .Z(n1607) );
  AND U2489 ( .A(n1612), .B(n1613), .Z(n1610) );
  XNOR U2490 ( .A(x[877]), .B(n1611), .Z(n1613) );
  XOR U2491 ( .A(n1614), .B(n1615), .Z(n1611) );
  AND U2492 ( .A(n1616), .B(n1617), .Z(n1614) );
  XNOR U2493 ( .A(x[876]), .B(n1615), .Z(n1617) );
  XOR U2494 ( .A(n1618), .B(n1619), .Z(n1615) );
  AND U2495 ( .A(n1620), .B(n1621), .Z(n1618) );
  XNOR U2496 ( .A(x[875]), .B(n1619), .Z(n1621) );
  XOR U2497 ( .A(n1622), .B(n1623), .Z(n1619) );
  AND U2498 ( .A(n1624), .B(n1625), .Z(n1622) );
  XNOR U2499 ( .A(x[874]), .B(n1623), .Z(n1625) );
  XOR U2500 ( .A(n1626), .B(n1627), .Z(n1623) );
  AND U2501 ( .A(n1628), .B(n1629), .Z(n1626) );
  XNOR U2502 ( .A(x[873]), .B(n1627), .Z(n1629) );
  XOR U2503 ( .A(n1630), .B(n1631), .Z(n1627) );
  AND U2504 ( .A(n1632), .B(n1633), .Z(n1630) );
  XNOR U2505 ( .A(x[872]), .B(n1631), .Z(n1633) );
  XOR U2506 ( .A(n1634), .B(n1635), .Z(n1631) );
  AND U2507 ( .A(n1636), .B(n1637), .Z(n1634) );
  XNOR U2508 ( .A(x[871]), .B(n1635), .Z(n1637) );
  XOR U2509 ( .A(n1638), .B(n1639), .Z(n1635) );
  AND U2510 ( .A(n1640), .B(n1641), .Z(n1638) );
  XNOR U2511 ( .A(x[870]), .B(n1639), .Z(n1641) );
  XOR U2512 ( .A(n1642), .B(n1643), .Z(n1639) );
  AND U2513 ( .A(n1644), .B(n1645), .Z(n1642) );
  XNOR U2514 ( .A(x[869]), .B(n1643), .Z(n1645) );
  XOR U2515 ( .A(n1646), .B(n1647), .Z(n1643) );
  AND U2516 ( .A(n1648), .B(n1649), .Z(n1646) );
  XNOR U2517 ( .A(x[868]), .B(n1647), .Z(n1649) );
  XOR U2518 ( .A(n1650), .B(n1651), .Z(n1647) );
  AND U2519 ( .A(n1652), .B(n1653), .Z(n1650) );
  XNOR U2520 ( .A(x[867]), .B(n1651), .Z(n1653) );
  XOR U2521 ( .A(n1654), .B(n1655), .Z(n1651) );
  AND U2522 ( .A(n1656), .B(n1657), .Z(n1654) );
  XNOR U2523 ( .A(x[866]), .B(n1655), .Z(n1657) );
  XOR U2524 ( .A(n1658), .B(n1659), .Z(n1655) );
  AND U2525 ( .A(n1660), .B(n1661), .Z(n1658) );
  XNOR U2526 ( .A(x[865]), .B(n1659), .Z(n1661) );
  XOR U2527 ( .A(n1662), .B(n1663), .Z(n1659) );
  AND U2528 ( .A(n1664), .B(n1665), .Z(n1662) );
  XNOR U2529 ( .A(x[864]), .B(n1663), .Z(n1665) );
  XOR U2530 ( .A(n1666), .B(n1667), .Z(n1663) );
  AND U2531 ( .A(n1668), .B(n1669), .Z(n1666) );
  XNOR U2532 ( .A(x[863]), .B(n1667), .Z(n1669) );
  XOR U2533 ( .A(n1670), .B(n1671), .Z(n1667) );
  AND U2534 ( .A(n1672), .B(n1673), .Z(n1670) );
  XNOR U2535 ( .A(x[862]), .B(n1671), .Z(n1673) );
  XOR U2536 ( .A(n1674), .B(n1675), .Z(n1671) );
  AND U2537 ( .A(n1676), .B(n1677), .Z(n1674) );
  XNOR U2538 ( .A(x[861]), .B(n1675), .Z(n1677) );
  XOR U2539 ( .A(n1678), .B(n1679), .Z(n1675) );
  AND U2540 ( .A(n1680), .B(n1681), .Z(n1678) );
  XNOR U2541 ( .A(x[860]), .B(n1679), .Z(n1681) );
  XOR U2542 ( .A(n1682), .B(n1683), .Z(n1679) );
  AND U2543 ( .A(n1684), .B(n1685), .Z(n1682) );
  XNOR U2544 ( .A(x[859]), .B(n1683), .Z(n1685) );
  XOR U2545 ( .A(n1686), .B(n1687), .Z(n1683) );
  AND U2546 ( .A(n1688), .B(n1689), .Z(n1686) );
  XNOR U2547 ( .A(x[858]), .B(n1687), .Z(n1689) );
  XOR U2548 ( .A(n1690), .B(n1691), .Z(n1687) );
  AND U2549 ( .A(n1692), .B(n1693), .Z(n1690) );
  XNOR U2550 ( .A(x[857]), .B(n1691), .Z(n1693) );
  XOR U2551 ( .A(n1694), .B(n1695), .Z(n1691) );
  AND U2552 ( .A(n1696), .B(n1697), .Z(n1694) );
  XNOR U2553 ( .A(x[856]), .B(n1695), .Z(n1697) );
  XOR U2554 ( .A(n1698), .B(n1699), .Z(n1695) );
  AND U2555 ( .A(n1700), .B(n1701), .Z(n1698) );
  XNOR U2556 ( .A(x[855]), .B(n1699), .Z(n1701) );
  XOR U2557 ( .A(n1702), .B(n1703), .Z(n1699) );
  AND U2558 ( .A(n1704), .B(n1705), .Z(n1702) );
  XNOR U2559 ( .A(x[854]), .B(n1703), .Z(n1705) );
  XOR U2560 ( .A(n1706), .B(n1707), .Z(n1703) );
  AND U2561 ( .A(n1708), .B(n1709), .Z(n1706) );
  XNOR U2562 ( .A(x[853]), .B(n1707), .Z(n1709) );
  XOR U2563 ( .A(n1710), .B(n1711), .Z(n1707) );
  AND U2564 ( .A(n1712), .B(n1713), .Z(n1710) );
  XNOR U2565 ( .A(x[852]), .B(n1711), .Z(n1713) );
  XOR U2566 ( .A(n1714), .B(n1715), .Z(n1711) );
  AND U2567 ( .A(n1716), .B(n1717), .Z(n1714) );
  XNOR U2568 ( .A(x[851]), .B(n1715), .Z(n1717) );
  XOR U2569 ( .A(n1718), .B(n1719), .Z(n1715) );
  AND U2570 ( .A(n1720), .B(n1721), .Z(n1718) );
  XNOR U2571 ( .A(x[850]), .B(n1719), .Z(n1721) );
  XOR U2572 ( .A(n1722), .B(n1723), .Z(n1719) );
  AND U2573 ( .A(n1724), .B(n1725), .Z(n1722) );
  XNOR U2574 ( .A(x[849]), .B(n1723), .Z(n1725) );
  XOR U2575 ( .A(n1726), .B(n1727), .Z(n1723) );
  AND U2576 ( .A(n1728), .B(n1729), .Z(n1726) );
  XNOR U2577 ( .A(x[848]), .B(n1727), .Z(n1729) );
  XOR U2578 ( .A(n1730), .B(n1731), .Z(n1727) );
  AND U2579 ( .A(n1732), .B(n1733), .Z(n1730) );
  XNOR U2580 ( .A(x[847]), .B(n1731), .Z(n1733) );
  XOR U2581 ( .A(n1734), .B(n1735), .Z(n1731) );
  AND U2582 ( .A(n1736), .B(n1737), .Z(n1734) );
  XNOR U2583 ( .A(x[846]), .B(n1735), .Z(n1737) );
  XOR U2584 ( .A(n1738), .B(n1739), .Z(n1735) );
  AND U2585 ( .A(n1740), .B(n1741), .Z(n1738) );
  XNOR U2586 ( .A(x[845]), .B(n1739), .Z(n1741) );
  XOR U2587 ( .A(n1742), .B(n1743), .Z(n1739) );
  AND U2588 ( .A(n1744), .B(n1745), .Z(n1742) );
  XNOR U2589 ( .A(x[844]), .B(n1743), .Z(n1745) );
  XOR U2590 ( .A(n1746), .B(n1747), .Z(n1743) );
  AND U2591 ( .A(n1748), .B(n1749), .Z(n1746) );
  XNOR U2592 ( .A(x[843]), .B(n1747), .Z(n1749) );
  XOR U2593 ( .A(n1750), .B(n1751), .Z(n1747) );
  AND U2594 ( .A(n1752), .B(n1753), .Z(n1750) );
  XNOR U2595 ( .A(x[842]), .B(n1751), .Z(n1753) );
  XOR U2596 ( .A(n1754), .B(n1755), .Z(n1751) );
  AND U2597 ( .A(n1756), .B(n1757), .Z(n1754) );
  XNOR U2598 ( .A(x[841]), .B(n1755), .Z(n1757) );
  XOR U2599 ( .A(n1758), .B(n1759), .Z(n1755) );
  AND U2600 ( .A(n1760), .B(n1761), .Z(n1758) );
  XNOR U2601 ( .A(x[840]), .B(n1759), .Z(n1761) );
  XOR U2602 ( .A(n1762), .B(n1763), .Z(n1759) );
  AND U2603 ( .A(n1764), .B(n1765), .Z(n1762) );
  XNOR U2604 ( .A(x[839]), .B(n1763), .Z(n1765) );
  XOR U2605 ( .A(n1766), .B(n1767), .Z(n1763) );
  AND U2606 ( .A(n1768), .B(n1769), .Z(n1766) );
  XNOR U2607 ( .A(x[838]), .B(n1767), .Z(n1769) );
  XOR U2608 ( .A(n1770), .B(n1771), .Z(n1767) );
  AND U2609 ( .A(n1772), .B(n1773), .Z(n1770) );
  XNOR U2610 ( .A(x[837]), .B(n1771), .Z(n1773) );
  XOR U2611 ( .A(n1774), .B(n1775), .Z(n1771) );
  AND U2612 ( .A(n1776), .B(n1777), .Z(n1774) );
  XNOR U2613 ( .A(x[836]), .B(n1775), .Z(n1777) );
  XOR U2614 ( .A(n1778), .B(n1779), .Z(n1775) );
  AND U2615 ( .A(n1780), .B(n1781), .Z(n1778) );
  XNOR U2616 ( .A(x[835]), .B(n1779), .Z(n1781) );
  XOR U2617 ( .A(n1782), .B(n1783), .Z(n1779) );
  AND U2618 ( .A(n1784), .B(n1785), .Z(n1782) );
  XNOR U2619 ( .A(x[834]), .B(n1783), .Z(n1785) );
  XOR U2620 ( .A(n1786), .B(n1787), .Z(n1783) );
  AND U2621 ( .A(n1788), .B(n1789), .Z(n1786) );
  XNOR U2622 ( .A(x[833]), .B(n1787), .Z(n1789) );
  XOR U2623 ( .A(n1790), .B(n1791), .Z(n1787) );
  AND U2624 ( .A(n1792), .B(n1793), .Z(n1790) );
  XNOR U2625 ( .A(x[832]), .B(n1791), .Z(n1793) );
  XOR U2626 ( .A(n1794), .B(n1795), .Z(n1791) );
  AND U2627 ( .A(n1796), .B(n1797), .Z(n1794) );
  XNOR U2628 ( .A(x[831]), .B(n1795), .Z(n1797) );
  XOR U2629 ( .A(n1798), .B(n1799), .Z(n1795) );
  AND U2630 ( .A(n1800), .B(n1801), .Z(n1798) );
  XNOR U2631 ( .A(x[830]), .B(n1799), .Z(n1801) );
  XOR U2632 ( .A(n1802), .B(n1803), .Z(n1799) );
  AND U2633 ( .A(n1804), .B(n1805), .Z(n1802) );
  XNOR U2634 ( .A(x[829]), .B(n1803), .Z(n1805) );
  XOR U2635 ( .A(n1806), .B(n1807), .Z(n1803) );
  AND U2636 ( .A(n1808), .B(n1809), .Z(n1806) );
  XNOR U2637 ( .A(x[828]), .B(n1807), .Z(n1809) );
  XOR U2638 ( .A(n1810), .B(n1811), .Z(n1807) );
  AND U2639 ( .A(n1812), .B(n1813), .Z(n1810) );
  XNOR U2640 ( .A(x[827]), .B(n1811), .Z(n1813) );
  XOR U2641 ( .A(n1814), .B(n1815), .Z(n1811) );
  AND U2642 ( .A(n1816), .B(n1817), .Z(n1814) );
  XNOR U2643 ( .A(x[826]), .B(n1815), .Z(n1817) );
  XOR U2644 ( .A(n1818), .B(n1819), .Z(n1815) );
  AND U2645 ( .A(n1820), .B(n1821), .Z(n1818) );
  XNOR U2646 ( .A(x[825]), .B(n1819), .Z(n1821) );
  XOR U2647 ( .A(n1822), .B(n1823), .Z(n1819) );
  AND U2648 ( .A(n1824), .B(n1825), .Z(n1822) );
  XNOR U2649 ( .A(x[824]), .B(n1823), .Z(n1825) );
  XOR U2650 ( .A(n1826), .B(n1827), .Z(n1823) );
  AND U2651 ( .A(n1828), .B(n1829), .Z(n1826) );
  XNOR U2652 ( .A(x[823]), .B(n1827), .Z(n1829) );
  XOR U2653 ( .A(n1830), .B(n1831), .Z(n1827) );
  AND U2654 ( .A(n1832), .B(n1833), .Z(n1830) );
  XNOR U2655 ( .A(x[822]), .B(n1831), .Z(n1833) );
  XOR U2656 ( .A(n1834), .B(n1835), .Z(n1831) );
  AND U2657 ( .A(n1836), .B(n1837), .Z(n1834) );
  XNOR U2658 ( .A(x[821]), .B(n1835), .Z(n1837) );
  XOR U2659 ( .A(n1838), .B(n1839), .Z(n1835) );
  AND U2660 ( .A(n1840), .B(n1841), .Z(n1838) );
  XNOR U2661 ( .A(x[820]), .B(n1839), .Z(n1841) );
  XOR U2662 ( .A(n1842), .B(n1843), .Z(n1839) );
  AND U2663 ( .A(n1844), .B(n1845), .Z(n1842) );
  XNOR U2664 ( .A(x[819]), .B(n1843), .Z(n1845) );
  XOR U2665 ( .A(n1846), .B(n1847), .Z(n1843) );
  AND U2666 ( .A(n1848), .B(n1849), .Z(n1846) );
  XNOR U2667 ( .A(x[818]), .B(n1847), .Z(n1849) );
  XOR U2668 ( .A(n1850), .B(n1851), .Z(n1847) );
  AND U2669 ( .A(n1852), .B(n1853), .Z(n1850) );
  XNOR U2670 ( .A(x[817]), .B(n1851), .Z(n1853) );
  XOR U2671 ( .A(n1854), .B(n1855), .Z(n1851) );
  AND U2672 ( .A(n1856), .B(n1857), .Z(n1854) );
  XNOR U2673 ( .A(x[816]), .B(n1855), .Z(n1857) );
  XOR U2674 ( .A(n1858), .B(n1859), .Z(n1855) );
  AND U2675 ( .A(n1860), .B(n1861), .Z(n1858) );
  XNOR U2676 ( .A(x[815]), .B(n1859), .Z(n1861) );
  XOR U2677 ( .A(n1862), .B(n1863), .Z(n1859) );
  AND U2678 ( .A(n1864), .B(n1865), .Z(n1862) );
  XNOR U2679 ( .A(x[814]), .B(n1863), .Z(n1865) );
  XOR U2680 ( .A(n1866), .B(n1867), .Z(n1863) );
  AND U2681 ( .A(n1868), .B(n1869), .Z(n1866) );
  XNOR U2682 ( .A(x[813]), .B(n1867), .Z(n1869) );
  XOR U2683 ( .A(n1870), .B(n1871), .Z(n1867) );
  AND U2684 ( .A(n1872), .B(n1873), .Z(n1870) );
  XNOR U2685 ( .A(x[812]), .B(n1871), .Z(n1873) );
  XOR U2686 ( .A(n1874), .B(n1875), .Z(n1871) );
  AND U2687 ( .A(n1876), .B(n1877), .Z(n1874) );
  XNOR U2688 ( .A(x[811]), .B(n1875), .Z(n1877) );
  XOR U2689 ( .A(n1878), .B(n1879), .Z(n1875) );
  AND U2690 ( .A(n1880), .B(n1881), .Z(n1878) );
  XNOR U2691 ( .A(x[810]), .B(n1879), .Z(n1881) );
  XOR U2692 ( .A(n1882), .B(n1883), .Z(n1879) );
  AND U2693 ( .A(n1884), .B(n1885), .Z(n1882) );
  XNOR U2694 ( .A(x[809]), .B(n1883), .Z(n1885) );
  XOR U2695 ( .A(n1886), .B(n1887), .Z(n1883) );
  AND U2696 ( .A(n1888), .B(n1889), .Z(n1886) );
  XNOR U2697 ( .A(x[808]), .B(n1887), .Z(n1889) );
  XOR U2698 ( .A(n1890), .B(n1891), .Z(n1887) );
  AND U2699 ( .A(n1892), .B(n1893), .Z(n1890) );
  XNOR U2700 ( .A(x[807]), .B(n1891), .Z(n1893) );
  XOR U2701 ( .A(n1894), .B(n1895), .Z(n1891) );
  AND U2702 ( .A(n1896), .B(n1897), .Z(n1894) );
  XNOR U2703 ( .A(x[806]), .B(n1895), .Z(n1897) );
  XOR U2704 ( .A(n1898), .B(n1899), .Z(n1895) );
  AND U2705 ( .A(n1900), .B(n1901), .Z(n1898) );
  XNOR U2706 ( .A(x[805]), .B(n1899), .Z(n1901) );
  XOR U2707 ( .A(n1902), .B(n1903), .Z(n1899) );
  AND U2708 ( .A(n1904), .B(n1905), .Z(n1902) );
  XNOR U2709 ( .A(x[804]), .B(n1903), .Z(n1905) );
  XOR U2710 ( .A(n1906), .B(n1907), .Z(n1903) );
  AND U2711 ( .A(n1908), .B(n1909), .Z(n1906) );
  XNOR U2712 ( .A(x[803]), .B(n1907), .Z(n1909) );
  XOR U2713 ( .A(n1910), .B(n1911), .Z(n1907) );
  AND U2714 ( .A(n1912), .B(n1913), .Z(n1910) );
  XNOR U2715 ( .A(x[802]), .B(n1911), .Z(n1913) );
  XOR U2716 ( .A(n1914), .B(n1915), .Z(n1911) );
  AND U2717 ( .A(n1916), .B(n1917), .Z(n1914) );
  XNOR U2718 ( .A(x[801]), .B(n1915), .Z(n1917) );
  XOR U2719 ( .A(n1918), .B(n1919), .Z(n1915) );
  AND U2720 ( .A(n1920), .B(n1921), .Z(n1918) );
  XNOR U2721 ( .A(x[800]), .B(n1919), .Z(n1921) );
  XOR U2722 ( .A(n1922), .B(n1923), .Z(n1919) );
  AND U2723 ( .A(n1924), .B(n1925), .Z(n1922) );
  XNOR U2724 ( .A(x[799]), .B(n1923), .Z(n1925) );
  XOR U2725 ( .A(n1926), .B(n1927), .Z(n1923) );
  AND U2726 ( .A(n1928), .B(n1929), .Z(n1926) );
  XNOR U2727 ( .A(x[798]), .B(n1927), .Z(n1929) );
  XOR U2728 ( .A(n1930), .B(n1931), .Z(n1927) );
  AND U2729 ( .A(n1932), .B(n1933), .Z(n1930) );
  XNOR U2730 ( .A(x[797]), .B(n1931), .Z(n1933) );
  XOR U2731 ( .A(n1934), .B(n1935), .Z(n1931) );
  AND U2732 ( .A(n1936), .B(n1937), .Z(n1934) );
  XNOR U2733 ( .A(x[796]), .B(n1935), .Z(n1937) );
  XOR U2734 ( .A(n1938), .B(n1939), .Z(n1935) );
  AND U2735 ( .A(n1940), .B(n1941), .Z(n1938) );
  XNOR U2736 ( .A(x[795]), .B(n1939), .Z(n1941) );
  XOR U2737 ( .A(n1942), .B(n1943), .Z(n1939) );
  AND U2738 ( .A(n1944), .B(n1945), .Z(n1942) );
  XNOR U2739 ( .A(x[794]), .B(n1943), .Z(n1945) );
  XOR U2740 ( .A(n1946), .B(n1947), .Z(n1943) );
  AND U2741 ( .A(n1948), .B(n1949), .Z(n1946) );
  XNOR U2742 ( .A(x[793]), .B(n1947), .Z(n1949) );
  XOR U2743 ( .A(n1950), .B(n1951), .Z(n1947) );
  AND U2744 ( .A(n1952), .B(n1953), .Z(n1950) );
  XNOR U2745 ( .A(x[792]), .B(n1951), .Z(n1953) );
  XOR U2746 ( .A(n1954), .B(n1955), .Z(n1951) );
  AND U2747 ( .A(n1956), .B(n1957), .Z(n1954) );
  XNOR U2748 ( .A(x[791]), .B(n1955), .Z(n1957) );
  XOR U2749 ( .A(n1958), .B(n1959), .Z(n1955) );
  AND U2750 ( .A(n1960), .B(n1961), .Z(n1958) );
  XNOR U2751 ( .A(x[790]), .B(n1959), .Z(n1961) );
  XOR U2752 ( .A(n1962), .B(n1963), .Z(n1959) );
  AND U2753 ( .A(n1964), .B(n1965), .Z(n1962) );
  XNOR U2754 ( .A(x[789]), .B(n1963), .Z(n1965) );
  XOR U2755 ( .A(n1966), .B(n1967), .Z(n1963) );
  AND U2756 ( .A(n1968), .B(n1969), .Z(n1966) );
  XNOR U2757 ( .A(x[788]), .B(n1967), .Z(n1969) );
  XOR U2758 ( .A(n1970), .B(n1971), .Z(n1967) );
  AND U2759 ( .A(n1972), .B(n1973), .Z(n1970) );
  XNOR U2760 ( .A(x[787]), .B(n1971), .Z(n1973) );
  XOR U2761 ( .A(n1974), .B(n1975), .Z(n1971) );
  AND U2762 ( .A(n1976), .B(n1977), .Z(n1974) );
  XNOR U2763 ( .A(x[786]), .B(n1975), .Z(n1977) );
  XOR U2764 ( .A(n1978), .B(n1979), .Z(n1975) );
  AND U2765 ( .A(n1980), .B(n1981), .Z(n1978) );
  XNOR U2766 ( .A(x[785]), .B(n1979), .Z(n1981) );
  XOR U2767 ( .A(n1982), .B(n1983), .Z(n1979) );
  AND U2768 ( .A(n1984), .B(n1985), .Z(n1982) );
  XNOR U2769 ( .A(x[784]), .B(n1983), .Z(n1985) );
  XOR U2770 ( .A(n1986), .B(n1987), .Z(n1983) );
  AND U2771 ( .A(n1988), .B(n1989), .Z(n1986) );
  XNOR U2772 ( .A(x[783]), .B(n1987), .Z(n1989) );
  XOR U2773 ( .A(n1990), .B(n1991), .Z(n1987) );
  AND U2774 ( .A(n1992), .B(n1993), .Z(n1990) );
  XNOR U2775 ( .A(x[782]), .B(n1991), .Z(n1993) );
  XOR U2776 ( .A(n1994), .B(n1995), .Z(n1991) );
  AND U2777 ( .A(n1996), .B(n1997), .Z(n1994) );
  XNOR U2778 ( .A(x[781]), .B(n1995), .Z(n1997) );
  XOR U2779 ( .A(n1998), .B(n1999), .Z(n1995) );
  AND U2780 ( .A(n2000), .B(n2001), .Z(n1998) );
  XNOR U2781 ( .A(x[780]), .B(n1999), .Z(n2001) );
  XOR U2782 ( .A(n2002), .B(n2003), .Z(n1999) );
  AND U2783 ( .A(n2004), .B(n2005), .Z(n2002) );
  XNOR U2784 ( .A(x[779]), .B(n2003), .Z(n2005) );
  XOR U2785 ( .A(n2006), .B(n2007), .Z(n2003) );
  AND U2786 ( .A(n2008), .B(n2009), .Z(n2006) );
  XNOR U2787 ( .A(x[778]), .B(n2007), .Z(n2009) );
  XOR U2788 ( .A(n2010), .B(n2011), .Z(n2007) );
  AND U2789 ( .A(n2012), .B(n2013), .Z(n2010) );
  XNOR U2790 ( .A(x[777]), .B(n2011), .Z(n2013) );
  XOR U2791 ( .A(n2014), .B(n2015), .Z(n2011) );
  AND U2792 ( .A(n2016), .B(n2017), .Z(n2014) );
  XNOR U2793 ( .A(x[776]), .B(n2015), .Z(n2017) );
  XOR U2794 ( .A(n2018), .B(n2019), .Z(n2015) );
  AND U2795 ( .A(n2020), .B(n2021), .Z(n2018) );
  XNOR U2796 ( .A(x[775]), .B(n2019), .Z(n2021) );
  XOR U2797 ( .A(n2022), .B(n2023), .Z(n2019) );
  AND U2798 ( .A(n2024), .B(n2025), .Z(n2022) );
  XNOR U2799 ( .A(x[774]), .B(n2023), .Z(n2025) );
  XOR U2800 ( .A(n2026), .B(n2027), .Z(n2023) );
  AND U2801 ( .A(n2028), .B(n2029), .Z(n2026) );
  XNOR U2802 ( .A(x[773]), .B(n2027), .Z(n2029) );
  XOR U2803 ( .A(n2030), .B(n2031), .Z(n2027) );
  AND U2804 ( .A(n2032), .B(n2033), .Z(n2030) );
  XNOR U2805 ( .A(x[772]), .B(n2031), .Z(n2033) );
  XOR U2806 ( .A(n2034), .B(n2035), .Z(n2031) );
  AND U2807 ( .A(n2036), .B(n2037), .Z(n2034) );
  XNOR U2808 ( .A(x[771]), .B(n2035), .Z(n2037) );
  XOR U2809 ( .A(n2038), .B(n2039), .Z(n2035) );
  AND U2810 ( .A(n2040), .B(n2041), .Z(n2038) );
  XNOR U2811 ( .A(x[770]), .B(n2039), .Z(n2041) );
  XOR U2812 ( .A(n2042), .B(n2043), .Z(n2039) );
  AND U2813 ( .A(n2044), .B(n2045), .Z(n2042) );
  XNOR U2814 ( .A(x[769]), .B(n2043), .Z(n2045) );
  XOR U2815 ( .A(n2046), .B(n2047), .Z(n2043) );
  AND U2816 ( .A(n2048), .B(n2049), .Z(n2046) );
  XNOR U2817 ( .A(x[768]), .B(n2047), .Z(n2049) );
  XOR U2818 ( .A(n2050), .B(n2051), .Z(n2047) );
  AND U2819 ( .A(n2052), .B(n2053), .Z(n2050) );
  XNOR U2820 ( .A(x[767]), .B(n2051), .Z(n2053) );
  XOR U2821 ( .A(n2054), .B(n2055), .Z(n2051) );
  AND U2822 ( .A(n2056), .B(n2057), .Z(n2054) );
  XNOR U2823 ( .A(x[766]), .B(n2055), .Z(n2057) );
  XOR U2824 ( .A(n2058), .B(n2059), .Z(n2055) );
  AND U2825 ( .A(n2060), .B(n2061), .Z(n2058) );
  XNOR U2826 ( .A(x[765]), .B(n2059), .Z(n2061) );
  XOR U2827 ( .A(n2062), .B(n2063), .Z(n2059) );
  AND U2828 ( .A(n2064), .B(n2065), .Z(n2062) );
  XNOR U2829 ( .A(x[764]), .B(n2063), .Z(n2065) );
  XOR U2830 ( .A(n2066), .B(n2067), .Z(n2063) );
  AND U2831 ( .A(n2068), .B(n2069), .Z(n2066) );
  XNOR U2832 ( .A(x[763]), .B(n2067), .Z(n2069) );
  XOR U2833 ( .A(n2070), .B(n2071), .Z(n2067) );
  AND U2834 ( .A(n2072), .B(n2073), .Z(n2070) );
  XNOR U2835 ( .A(x[762]), .B(n2071), .Z(n2073) );
  XOR U2836 ( .A(n2074), .B(n2075), .Z(n2071) );
  AND U2837 ( .A(n2076), .B(n2077), .Z(n2074) );
  XNOR U2838 ( .A(x[761]), .B(n2075), .Z(n2077) );
  XOR U2839 ( .A(n2078), .B(n2079), .Z(n2075) );
  AND U2840 ( .A(n2080), .B(n2081), .Z(n2078) );
  XNOR U2841 ( .A(x[760]), .B(n2079), .Z(n2081) );
  XOR U2842 ( .A(n2082), .B(n2083), .Z(n2079) );
  AND U2843 ( .A(n2084), .B(n2085), .Z(n2082) );
  XNOR U2844 ( .A(x[759]), .B(n2083), .Z(n2085) );
  XOR U2845 ( .A(n2086), .B(n2087), .Z(n2083) );
  AND U2846 ( .A(n2088), .B(n2089), .Z(n2086) );
  XNOR U2847 ( .A(x[758]), .B(n2087), .Z(n2089) );
  XOR U2848 ( .A(n2090), .B(n2091), .Z(n2087) );
  AND U2849 ( .A(n2092), .B(n2093), .Z(n2090) );
  XNOR U2850 ( .A(x[757]), .B(n2091), .Z(n2093) );
  XOR U2851 ( .A(n2094), .B(n2095), .Z(n2091) );
  AND U2852 ( .A(n2096), .B(n2097), .Z(n2094) );
  XNOR U2853 ( .A(x[756]), .B(n2095), .Z(n2097) );
  XOR U2854 ( .A(n2098), .B(n2099), .Z(n2095) );
  AND U2855 ( .A(n2100), .B(n2101), .Z(n2098) );
  XNOR U2856 ( .A(x[755]), .B(n2099), .Z(n2101) );
  XOR U2857 ( .A(n2102), .B(n2103), .Z(n2099) );
  AND U2858 ( .A(n2104), .B(n2105), .Z(n2102) );
  XNOR U2859 ( .A(x[754]), .B(n2103), .Z(n2105) );
  XOR U2860 ( .A(n2106), .B(n2107), .Z(n2103) );
  AND U2861 ( .A(n2108), .B(n2109), .Z(n2106) );
  XNOR U2862 ( .A(x[753]), .B(n2107), .Z(n2109) );
  XOR U2863 ( .A(n2110), .B(n2111), .Z(n2107) );
  AND U2864 ( .A(n2112), .B(n2113), .Z(n2110) );
  XNOR U2865 ( .A(x[752]), .B(n2111), .Z(n2113) );
  XOR U2866 ( .A(n2114), .B(n2115), .Z(n2111) );
  AND U2867 ( .A(n2116), .B(n2117), .Z(n2114) );
  XNOR U2868 ( .A(x[751]), .B(n2115), .Z(n2117) );
  XOR U2869 ( .A(n2118), .B(n2119), .Z(n2115) );
  AND U2870 ( .A(n2120), .B(n2121), .Z(n2118) );
  XNOR U2871 ( .A(x[750]), .B(n2119), .Z(n2121) );
  XOR U2872 ( .A(n2122), .B(n2123), .Z(n2119) );
  AND U2873 ( .A(n2124), .B(n2125), .Z(n2122) );
  XNOR U2874 ( .A(x[749]), .B(n2123), .Z(n2125) );
  XOR U2875 ( .A(n2126), .B(n2127), .Z(n2123) );
  AND U2876 ( .A(n2128), .B(n2129), .Z(n2126) );
  XNOR U2877 ( .A(x[748]), .B(n2127), .Z(n2129) );
  XOR U2878 ( .A(n2130), .B(n2131), .Z(n2127) );
  AND U2879 ( .A(n2132), .B(n2133), .Z(n2130) );
  XNOR U2880 ( .A(x[747]), .B(n2131), .Z(n2133) );
  XOR U2881 ( .A(n2134), .B(n2135), .Z(n2131) );
  AND U2882 ( .A(n2136), .B(n2137), .Z(n2134) );
  XNOR U2883 ( .A(x[746]), .B(n2135), .Z(n2137) );
  XOR U2884 ( .A(n2138), .B(n2139), .Z(n2135) );
  AND U2885 ( .A(n2140), .B(n2141), .Z(n2138) );
  XNOR U2886 ( .A(x[745]), .B(n2139), .Z(n2141) );
  XOR U2887 ( .A(n2142), .B(n2143), .Z(n2139) );
  AND U2888 ( .A(n2144), .B(n2145), .Z(n2142) );
  XNOR U2889 ( .A(x[744]), .B(n2143), .Z(n2145) );
  XOR U2890 ( .A(n2146), .B(n2147), .Z(n2143) );
  AND U2891 ( .A(n2148), .B(n2149), .Z(n2146) );
  XNOR U2892 ( .A(x[743]), .B(n2147), .Z(n2149) );
  XOR U2893 ( .A(n2150), .B(n2151), .Z(n2147) );
  AND U2894 ( .A(n2152), .B(n2153), .Z(n2150) );
  XNOR U2895 ( .A(x[742]), .B(n2151), .Z(n2153) );
  XOR U2896 ( .A(n2154), .B(n2155), .Z(n2151) );
  AND U2897 ( .A(n2156), .B(n2157), .Z(n2154) );
  XNOR U2898 ( .A(x[741]), .B(n2155), .Z(n2157) );
  XOR U2899 ( .A(n2158), .B(n2159), .Z(n2155) );
  AND U2900 ( .A(n2160), .B(n2161), .Z(n2158) );
  XNOR U2901 ( .A(x[740]), .B(n2159), .Z(n2161) );
  XOR U2902 ( .A(n2162), .B(n2163), .Z(n2159) );
  AND U2903 ( .A(n2164), .B(n2165), .Z(n2162) );
  XNOR U2904 ( .A(x[739]), .B(n2163), .Z(n2165) );
  XOR U2905 ( .A(n2166), .B(n2167), .Z(n2163) );
  AND U2906 ( .A(n2168), .B(n2169), .Z(n2166) );
  XNOR U2907 ( .A(x[738]), .B(n2167), .Z(n2169) );
  XOR U2908 ( .A(n2170), .B(n2171), .Z(n2167) );
  AND U2909 ( .A(n2172), .B(n2173), .Z(n2170) );
  XNOR U2910 ( .A(x[737]), .B(n2171), .Z(n2173) );
  XOR U2911 ( .A(n2174), .B(n2175), .Z(n2171) );
  AND U2912 ( .A(n2176), .B(n2177), .Z(n2174) );
  XNOR U2913 ( .A(x[736]), .B(n2175), .Z(n2177) );
  XOR U2914 ( .A(n2178), .B(n2179), .Z(n2175) );
  AND U2915 ( .A(n2180), .B(n2181), .Z(n2178) );
  XNOR U2916 ( .A(x[735]), .B(n2179), .Z(n2181) );
  XOR U2917 ( .A(n2182), .B(n2183), .Z(n2179) );
  AND U2918 ( .A(n2184), .B(n2185), .Z(n2182) );
  XNOR U2919 ( .A(x[734]), .B(n2183), .Z(n2185) );
  XOR U2920 ( .A(n2186), .B(n2187), .Z(n2183) );
  AND U2921 ( .A(n2188), .B(n2189), .Z(n2186) );
  XNOR U2922 ( .A(x[733]), .B(n2187), .Z(n2189) );
  XOR U2923 ( .A(n2190), .B(n2191), .Z(n2187) );
  AND U2924 ( .A(n2192), .B(n2193), .Z(n2190) );
  XNOR U2925 ( .A(x[732]), .B(n2191), .Z(n2193) );
  XOR U2926 ( .A(n2194), .B(n2195), .Z(n2191) );
  AND U2927 ( .A(n2196), .B(n2197), .Z(n2194) );
  XNOR U2928 ( .A(x[731]), .B(n2195), .Z(n2197) );
  XOR U2929 ( .A(n2198), .B(n2199), .Z(n2195) );
  AND U2930 ( .A(n2200), .B(n2201), .Z(n2198) );
  XNOR U2931 ( .A(x[730]), .B(n2199), .Z(n2201) );
  XOR U2932 ( .A(n2202), .B(n2203), .Z(n2199) );
  AND U2933 ( .A(n2204), .B(n2205), .Z(n2202) );
  XNOR U2934 ( .A(x[729]), .B(n2203), .Z(n2205) );
  XOR U2935 ( .A(n2206), .B(n2207), .Z(n2203) );
  AND U2936 ( .A(n2208), .B(n2209), .Z(n2206) );
  XNOR U2937 ( .A(x[728]), .B(n2207), .Z(n2209) );
  XOR U2938 ( .A(n2210), .B(n2211), .Z(n2207) );
  AND U2939 ( .A(n2212), .B(n2213), .Z(n2210) );
  XNOR U2940 ( .A(x[727]), .B(n2211), .Z(n2213) );
  XOR U2941 ( .A(n2214), .B(n2215), .Z(n2211) );
  AND U2942 ( .A(n2216), .B(n2217), .Z(n2214) );
  XNOR U2943 ( .A(x[726]), .B(n2215), .Z(n2217) );
  XOR U2944 ( .A(n2218), .B(n2219), .Z(n2215) );
  AND U2945 ( .A(n2220), .B(n2221), .Z(n2218) );
  XNOR U2946 ( .A(x[725]), .B(n2219), .Z(n2221) );
  XOR U2947 ( .A(n2222), .B(n2223), .Z(n2219) );
  AND U2948 ( .A(n2224), .B(n2225), .Z(n2222) );
  XNOR U2949 ( .A(x[724]), .B(n2223), .Z(n2225) );
  XOR U2950 ( .A(n2226), .B(n2227), .Z(n2223) );
  AND U2951 ( .A(n2228), .B(n2229), .Z(n2226) );
  XNOR U2952 ( .A(x[723]), .B(n2227), .Z(n2229) );
  XOR U2953 ( .A(n2230), .B(n2231), .Z(n2227) );
  AND U2954 ( .A(n2232), .B(n2233), .Z(n2230) );
  XNOR U2955 ( .A(x[722]), .B(n2231), .Z(n2233) );
  XOR U2956 ( .A(n2234), .B(n2235), .Z(n2231) );
  AND U2957 ( .A(n2236), .B(n2237), .Z(n2234) );
  XNOR U2958 ( .A(x[721]), .B(n2235), .Z(n2237) );
  XOR U2959 ( .A(n2238), .B(n2239), .Z(n2235) );
  AND U2960 ( .A(n2240), .B(n2241), .Z(n2238) );
  XNOR U2961 ( .A(x[720]), .B(n2239), .Z(n2241) );
  XOR U2962 ( .A(n2242), .B(n2243), .Z(n2239) );
  AND U2963 ( .A(n2244), .B(n2245), .Z(n2242) );
  XNOR U2964 ( .A(x[719]), .B(n2243), .Z(n2245) );
  XOR U2965 ( .A(n2246), .B(n2247), .Z(n2243) );
  AND U2966 ( .A(n2248), .B(n2249), .Z(n2246) );
  XNOR U2967 ( .A(x[718]), .B(n2247), .Z(n2249) );
  XOR U2968 ( .A(n2250), .B(n2251), .Z(n2247) );
  AND U2969 ( .A(n2252), .B(n2253), .Z(n2250) );
  XNOR U2970 ( .A(x[717]), .B(n2251), .Z(n2253) );
  XOR U2971 ( .A(n2254), .B(n2255), .Z(n2251) );
  AND U2972 ( .A(n2256), .B(n2257), .Z(n2254) );
  XNOR U2973 ( .A(x[716]), .B(n2255), .Z(n2257) );
  XOR U2974 ( .A(n2258), .B(n2259), .Z(n2255) );
  AND U2975 ( .A(n2260), .B(n2261), .Z(n2258) );
  XNOR U2976 ( .A(x[715]), .B(n2259), .Z(n2261) );
  XOR U2977 ( .A(n2262), .B(n2263), .Z(n2259) );
  AND U2978 ( .A(n2264), .B(n2265), .Z(n2262) );
  XNOR U2979 ( .A(x[714]), .B(n2263), .Z(n2265) );
  XOR U2980 ( .A(n2266), .B(n2267), .Z(n2263) );
  AND U2981 ( .A(n2268), .B(n2269), .Z(n2266) );
  XNOR U2982 ( .A(x[713]), .B(n2267), .Z(n2269) );
  XOR U2983 ( .A(n2270), .B(n2271), .Z(n2267) );
  AND U2984 ( .A(n2272), .B(n2273), .Z(n2270) );
  XNOR U2985 ( .A(x[712]), .B(n2271), .Z(n2273) );
  XOR U2986 ( .A(n2274), .B(n2275), .Z(n2271) );
  AND U2987 ( .A(n2276), .B(n2277), .Z(n2274) );
  XNOR U2988 ( .A(x[711]), .B(n2275), .Z(n2277) );
  XOR U2989 ( .A(n2278), .B(n2279), .Z(n2275) );
  AND U2990 ( .A(n2280), .B(n2281), .Z(n2278) );
  XNOR U2991 ( .A(x[710]), .B(n2279), .Z(n2281) );
  XOR U2992 ( .A(n2282), .B(n2283), .Z(n2279) );
  AND U2993 ( .A(n2284), .B(n2285), .Z(n2282) );
  XNOR U2994 ( .A(x[709]), .B(n2283), .Z(n2285) );
  XOR U2995 ( .A(n2286), .B(n2287), .Z(n2283) );
  AND U2996 ( .A(n2288), .B(n2289), .Z(n2286) );
  XNOR U2997 ( .A(x[708]), .B(n2287), .Z(n2289) );
  XOR U2998 ( .A(n2290), .B(n2291), .Z(n2287) );
  AND U2999 ( .A(n2292), .B(n2293), .Z(n2290) );
  XNOR U3000 ( .A(x[707]), .B(n2291), .Z(n2293) );
  XOR U3001 ( .A(n2294), .B(n2295), .Z(n2291) );
  AND U3002 ( .A(n2296), .B(n2297), .Z(n2294) );
  XNOR U3003 ( .A(x[706]), .B(n2295), .Z(n2297) );
  XOR U3004 ( .A(n2298), .B(n2299), .Z(n2295) );
  AND U3005 ( .A(n2300), .B(n2301), .Z(n2298) );
  XNOR U3006 ( .A(x[705]), .B(n2299), .Z(n2301) );
  XOR U3007 ( .A(n2302), .B(n2303), .Z(n2299) );
  AND U3008 ( .A(n2304), .B(n2305), .Z(n2302) );
  XNOR U3009 ( .A(x[704]), .B(n2303), .Z(n2305) );
  XOR U3010 ( .A(n2306), .B(n2307), .Z(n2303) );
  AND U3011 ( .A(n2308), .B(n2309), .Z(n2306) );
  XNOR U3012 ( .A(x[703]), .B(n2307), .Z(n2309) );
  XOR U3013 ( .A(n2310), .B(n2311), .Z(n2307) );
  AND U3014 ( .A(n2312), .B(n2313), .Z(n2310) );
  XNOR U3015 ( .A(x[702]), .B(n2311), .Z(n2313) );
  XOR U3016 ( .A(n2314), .B(n2315), .Z(n2311) );
  AND U3017 ( .A(n2316), .B(n2317), .Z(n2314) );
  XNOR U3018 ( .A(x[701]), .B(n2315), .Z(n2317) );
  XOR U3019 ( .A(n2318), .B(n2319), .Z(n2315) );
  AND U3020 ( .A(n2320), .B(n2321), .Z(n2318) );
  XNOR U3021 ( .A(x[700]), .B(n2319), .Z(n2321) );
  XOR U3022 ( .A(n2322), .B(n2323), .Z(n2319) );
  AND U3023 ( .A(n2324), .B(n2325), .Z(n2322) );
  XNOR U3024 ( .A(x[699]), .B(n2323), .Z(n2325) );
  XOR U3025 ( .A(n2326), .B(n2327), .Z(n2323) );
  AND U3026 ( .A(n2328), .B(n2329), .Z(n2326) );
  XNOR U3027 ( .A(x[698]), .B(n2327), .Z(n2329) );
  XOR U3028 ( .A(n2330), .B(n2331), .Z(n2327) );
  AND U3029 ( .A(n2332), .B(n2333), .Z(n2330) );
  XNOR U3030 ( .A(x[697]), .B(n2331), .Z(n2333) );
  XOR U3031 ( .A(n2334), .B(n2335), .Z(n2331) );
  AND U3032 ( .A(n2336), .B(n2337), .Z(n2334) );
  XNOR U3033 ( .A(x[696]), .B(n2335), .Z(n2337) );
  XOR U3034 ( .A(n2338), .B(n2339), .Z(n2335) );
  AND U3035 ( .A(n2340), .B(n2341), .Z(n2338) );
  XNOR U3036 ( .A(x[695]), .B(n2339), .Z(n2341) );
  XOR U3037 ( .A(n2342), .B(n2343), .Z(n2339) );
  AND U3038 ( .A(n2344), .B(n2345), .Z(n2342) );
  XNOR U3039 ( .A(x[694]), .B(n2343), .Z(n2345) );
  XOR U3040 ( .A(n2346), .B(n2347), .Z(n2343) );
  AND U3041 ( .A(n2348), .B(n2349), .Z(n2346) );
  XNOR U3042 ( .A(x[693]), .B(n2347), .Z(n2349) );
  XOR U3043 ( .A(n2350), .B(n2351), .Z(n2347) );
  AND U3044 ( .A(n2352), .B(n2353), .Z(n2350) );
  XNOR U3045 ( .A(x[692]), .B(n2351), .Z(n2353) );
  XOR U3046 ( .A(n2354), .B(n2355), .Z(n2351) );
  AND U3047 ( .A(n2356), .B(n2357), .Z(n2354) );
  XNOR U3048 ( .A(x[691]), .B(n2355), .Z(n2357) );
  XOR U3049 ( .A(n2358), .B(n2359), .Z(n2355) );
  AND U3050 ( .A(n2360), .B(n2361), .Z(n2358) );
  XNOR U3051 ( .A(x[690]), .B(n2359), .Z(n2361) );
  XOR U3052 ( .A(n2362), .B(n2363), .Z(n2359) );
  AND U3053 ( .A(n2364), .B(n2365), .Z(n2362) );
  XNOR U3054 ( .A(x[689]), .B(n2363), .Z(n2365) );
  XOR U3055 ( .A(n2366), .B(n2367), .Z(n2363) );
  AND U3056 ( .A(n2368), .B(n2369), .Z(n2366) );
  XNOR U3057 ( .A(x[688]), .B(n2367), .Z(n2369) );
  XOR U3058 ( .A(n2370), .B(n2371), .Z(n2367) );
  AND U3059 ( .A(n2372), .B(n2373), .Z(n2370) );
  XNOR U3060 ( .A(x[687]), .B(n2371), .Z(n2373) );
  XOR U3061 ( .A(n2374), .B(n2375), .Z(n2371) );
  AND U3062 ( .A(n2376), .B(n2377), .Z(n2374) );
  XNOR U3063 ( .A(x[686]), .B(n2375), .Z(n2377) );
  XOR U3064 ( .A(n2378), .B(n2379), .Z(n2375) );
  AND U3065 ( .A(n2380), .B(n2381), .Z(n2378) );
  XNOR U3066 ( .A(x[685]), .B(n2379), .Z(n2381) );
  XOR U3067 ( .A(n2382), .B(n2383), .Z(n2379) );
  AND U3068 ( .A(n2384), .B(n2385), .Z(n2382) );
  XNOR U3069 ( .A(x[684]), .B(n2383), .Z(n2385) );
  XOR U3070 ( .A(n2386), .B(n2387), .Z(n2383) );
  AND U3071 ( .A(n2388), .B(n2389), .Z(n2386) );
  XNOR U3072 ( .A(x[683]), .B(n2387), .Z(n2389) );
  XOR U3073 ( .A(n2390), .B(n2391), .Z(n2387) );
  AND U3074 ( .A(n2392), .B(n2393), .Z(n2390) );
  XNOR U3075 ( .A(x[682]), .B(n2391), .Z(n2393) );
  XOR U3076 ( .A(n2394), .B(n2395), .Z(n2391) );
  AND U3077 ( .A(n2396), .B(n2397), .Z(n2394) );
  XNOR U3078 ( .A(x[681]), .B(n2395), .Z(n2397) );
  XOR U3079 ( .A(n2398), .B(n2399), .Z(n2395) );
  AND U3080 ( .A(n2400), .B(n2401), .Z(n2398) );
  XNOR U3081 ( .A(x[680]), .B(n2399), .Z(n2401) );
  XOR U3082 ( .A(n2402), .B(n2403), .Z(n2399) );
  AND U3083 ( .A(n2404), .B(n2405), .Z(n2402) );
  XNOR U3084 ( .A(x[679]), .B(n2403), .Z(n2405) );
  XOR U3085 ( .A(n2406), .B(n2407), .Z(n2403) );
  AND U3086 ( .A(n2408), .B(n2409), .Z(n2406) );
  XNOR U3087 ( .A(x[678]), .B(n2407), .Z(n2409) );
  XOR U3088 ( .A(n2410), .B(n2411), .Z(n2407) );
  AND U3089 ( .A(n2412), .B(n2413), .Z(n2410) );
  XNOR U3090 ( .A(x[677]), .B(n2411), .Z(n2413) );
  XOR U3091 ( .A(n2414), .B(n2415), .Z(n2411) );
  AND U3092 ( .A(n2416), .B(n2417), .Z(n2414) );
  XNOR U3093 ( .A(x[676]), .B(n2415), .Z(n2417) );
  XOR U3094 ( .A(n2418), .B(n2419), .Z(n2415) );
  AND U3095 ( .A(n2420), .B(n2421), .Z(n2418) );
  XNOR U3096 ( .A(x[675]), .B(n2419), .Z(n2421) );
  XOR U3097 ( .A(n2422), .B(n2423), .Z(n2419) );
  AND U3098 ( .A(n2424), .B(n2425), .Z(n2422) );
  XNOR U3099 ( .A(x[674]), .B(n2423), .Z(n2425) );
  XOR U3100 ( .A(n2426), .B(n2427), .Z(n2423) );
  AND U3101 ( .A(n2428), .B(n2429), .Z(n2426) );
  XNOR U3102 ( .A(x[673]), .B(n2427), .Z(n2429) );
  XOR U3103 ( .A(n2430), .B(n2431), .Z(n2427) );
  AND U3104 ( .A(n2432), .B(n2433), .Z(n2430) );
  XNOR U3105 ( .A(x[672]), .B(n2431), .Z(n2433) );
  XOR U3106 ( .A(n2434), .B(n2435), .Z(n2431) );
  AND U3107 ( .A(n2436), .B(n2437), .Z(n2434) );
  XNOR U3108 ( .A(x[671]), .B(n2435), .Z(n2437) );
  XOR U3109 ( .A(n2438), .B(n2439), .Z(n2435) );
  AND U3110 ( .A(n2440), .B(n2441), .Z(n2438) );
  XNOR U3111 ( .A(x[670]), .B(n2439), .Z(n2441) );
  XOR U3112 ( .A(n2442), .B(n2443), .Z(n2439) );
  AND U3113 ( .A(n2444), .B(n2445), .Z(n2442) );
  XNOR U3114 ( .A(x[669]), .B(n2443), .Z(n2445) );
  XOR U3115 ( .A(n2446), .B(n2447), .Z(n2443) );
  AND U3116 ( .A(n2448), .B(n2449), .Z(n2446) );
  XNOR U3117 ( .A(x[668]), .B(n2447), .Z(n2449) );
  XOR U3118 ( .A(n2450), .B(n2451), .Z(n2447) );
  AND U3119 ( .A(n2452), .B(n2453), .Z(n2450) );
  XNOR U3120 ( .A(x[667]), .B(n2451), .Z(n2453) );
  XOR U3121 ( .A(n2454), .B(n2455), .Z(n2451) );
  AND U3122 ( .A(n2456), .B(n2457), .Z(n2454) );
  XNOR U3123 ( .A(x[666]), .B(n2455), .Z(n2457) );
  XOR U3124 ( .A(n2458), .B(n2459), .Z(n2455) );
  AND U3125 ( .A(n2460), .B(n2461), .Z(n2458) );
  XNOR U3126 ( .A(x[665]), .B(n2459), .Z(n2461) );
  XOR U3127 ( .A(n2462), .B(n2463), .Z(n2459) );
  AND U3128 ( .A(n2464), .B(n2465), .Z(n2462) );
  XNOR U3129 ( .A(x[664]), .B(n2463), .Z(n2465) );
  XOR U3130 ( .A(n2466), .B(n2467), .Z(n2463) );
  AND U3131 ( .A(n2468), .B(n2469), .Z(n2466) );
  XNOR U3132 ( .A(x[663]), .B(n2467), .Z(n2469) );
  XOR U3133 ( .A(n2470), .B(n2471), .Z(n2467) );
  AND U3134 ( .A(n2472), .B(n2473), .Z(n2470) );
  XNOR U3135 ( .A(x[662]), .B(n2471), .Z(n2473) );
  XOR U3136 ( .A(n2474), .B(n2475), .Z(n2471) );
  AND U3137 ( .A(n2476), .B(n2477), .Z(n2474) );
  XNOR U3138 ( .A(x[661]), .B(n2475), .Z(n2477) );
  XOR U3139 ( .A(n2478), .B(n2479), .Z(n2475) );
  AND U3140 ( .A(n2480), .B(n2481), .Z(n2478) );
  XNOR U3141 ( .A(x[660]), .B(n2479), .Z(n2481) );
  XOR U3142 ( .A(n2482), .B(n2483), .Z(n2479) );
  AND U3143 ( .A(n2484), .B(n2485), .Z(n2482) );
  XNOR U3144 ( .A(x[659]), .B(n2483), .Z(n2485) );
  XOR U3145 ( .A(n2486), .B(n2487), .Z(n2483) );
  AND U3146 ( .A(n2488), .B(n2489), .Z(n2486) );
  XNOR U3147 ( .A(x[658]), .B(n2487), .Z(n2489) );
  XOR U3148 ( .A(n2490), .B(n2491), .Z(n2487) );
  AND U3149 ( .A(n2492), .B(n2493), .Z(n2490) );
  XNOR U3150 ( .A(x[657]), .B(n2491), .Z(n2493) );
  XOR U3151 ( .A(n2494), .B(n2495), .Z(n2491) );
  AND U3152 ( .A(n2496), .B(n2497), .Z(n2494) );
  XNOR U3153 ( .A(x[656]), .B(n2495), .Z(n2497) );
  XOR U3154 ( .A(n2498), .B(n2499), .Z(n2495) );
  AND U3155 ( .A(n2500), .B(n2501), .Z(n2498) );
  XNOR U3156 ( .A(x[655]), .B(n2499), .Z(n2501) );
  XOR U3157 ( .A(n2502), .B(n2503), .Z(n2499) );
  AND U3158 ( .A(n2504), .B(n2505), .Z(n2502) );
  XNOR U3159 ( .A(x[654]), .B(n2503), .Z(n2505) );
  XOR U3160 ( .A(n2506), .B(n2507), .Z(n2503) );
  AND U3161 ( .A(n2508), .B(n2509), .Z(n2506) );
  XNOR U3162 ( .A(x[653]), .B(n2507), .Z(n2509) );
  XOR U3163 ( .A(n2510), .B(n2511), .Z(n2507) );
  AND U3164 ( .A(n2512), .B(n2513), .Z(n2510) );
  XNOR U3165 ( .A(x[652]), .B(n2511), .Z(n2513) );
  XOR U3166 ( .A(n2514), .B(n2515), .Z(n2511) );
  AND U3167 ( .A(n2516), .B(n2517), .Z(n2514) );
  XNOR U3168 ( .A(x[651]), .B(n2515), .Z(n2517) );
  XOR U3169 ( .A(n2518), .B(n2519), .Z(n2515) );
  AND U3170 ( .A(n2520), .B(n2521), .Z(n2518) );
  XNOR U3171 ( .A(x[650]), .B(n2519), .Z(n2521) );
  XOR U3172 ( .A(n2522), .B(n2523), .Z(n2519) );
  AND U3173 ( .A(n2524), .B(n2525), .Z(n2522) );
  XNOR U3174 ( .A(x[649]), .B(n2523), .Z(n2525) );
  XOR U3175 ( .A(n2526), .B(n2527), .Z(n2523) );
  AND U3176 ( .A(n2528), .B(n2529), .Z(n2526) );
  XNOR U3177 ( .A(x[648]), .B(n2527), .Z(n2529) );
  XOR U3178 ( .A(n2530), .B(n2531), .Z(n2527) );
  AND U3179 ( .A(n2532), .B(n2533), .Z(n2530) );
  XNOR U3180 ( .A(x[647]), .B(n2531), .Z(n2533) );
  XOR U3181 ( .A(n2534), .B(n2535), .Z(n2531) );
  AND U3182 ( .A(n2536), .B(n2537), .Z(n2534) );
  XNOR U3183 ( .A(x[646]), .B(n2535), .Z(n2537) );
  XOR U3184 ( .A(n2538), .B(n2539), .Z(n2535) );
  AND U3185 ( .A(n2540), .B(n2541), .Z(n2538) );
  XNOR U3186 ( .A(x[645]), .B(n2539), .Z(n2541) );
  XOR U3187 ( .A(n2542), .B(n2543), .Z(n2539) );
  AND U3188 ( .A(n2544), .B(n2545), .Z(n2542) );
  XNOR U3189 ( .A(x[644]), .B(n2543), .Z(n2545) );
  XOR U3190 ( .A(n2546), .B(n2547), .Z(n2543) );
  AND U3191 ( .A(n2548), .B(n2549), .Z(n2546) );
  XNOR U3192 ( .A(x[643]), .B(n2547), .Z(n2549) );
  XOR U3193 ( .A(n2550), .B(n2551), .Z(n2547) );
  AND U3194 ( .A(n2552), .B(n2553), .Z(n2550) );
  XNOR U3195 ( .A(x[642]), .B(n2551), .Z(n2553) );
  XOR U3196 ( .A(n2554), .B(n2555), .Z(n2551) );
  AND U3197 ( .A(n2556), .B(n2557), .Z(n2554) );
  XNOR U3198 ( .A(x[641]), .B(n2555), .Z(n2557) );
  XOR U3199 ( .A(n2558), .B(n2559), .Z(n2555) );
  AND U3200 ( .A(n2560), .B(n2561), .Z(n2558) );
  XNOR U3201 ( .A(x[640]), .B(n2559), .Z(n2561) );
  XOR U3202 ( .A(n2562), .B(n2563), .Z(n2559) );
  AND U3203 ( .A(n2564), .B(n2565), .Z(n2562) );
  XNOR U3204 ( .A(x[639]), .B(n2563), .Z(n2565) );
  XOR U3205 ( .A(n2566), .B(n2567), .Z(n2563) );
  AND U3206 ( .A(n2568), .B(n2569), .Z(n2566) );
  XNOR U3207 ( .A(x[638]), .B(n2567), .Z(n2569) );
  XOR U3208 ( .A(n2570), .B(n2571), .Z(n2567) );
  AND U3209 ( .A(n2572), .B(n2573), .Z(n2570) );
  XNOR U3210 ( .A(x[637]), .B(n2571), .Z(n2573) );
  XOR U3211 ( .A(n2574), .B(n2575), .Z(n2571) );
  AND U3212 ( .A(n2576), .B(n2577), .Z(n2574) );
  XNOR U3213 ( .A(x[636]), .B(n2575), .Z(n2577) );
  XOR U3214 ( .A(n2578), .B(n2579), .Z(n2575) );
  AND U3215 ( .A(n2580), .B(n2581), .Z(n2578) );
  XNOR U3216 ( .A(x[635]), .B(n2579), .Z(n2581) );
  XOR U3217 ( .A(n2582), .B(n2583), .Z(n2579) );
  AND U3218 ( .A(n2584), .B(n2585), .Z(n2582) );
  XNOR U3219 ( .A(x[634]), .B(n2583), .Z(n2585) );
  XOR U3220 ( .A(n2586), .B(n2587), .Z(n2583) );
  AND U3221 ( .A(n2588), .B(n2589), .Z(n2586) );
  XNOR U3222 ( .A(x[633]), .B(n2587), .Z(n2589) );
  XOR U3223 ( .A(n2590), .B(n2591), .Z(n2587) );
  AND U3224 ( .A(n2592), .B(n2593), .Z(n2590) );
  XNOR U3225 ( .A(x[632]), .B(n2591), .Z(n2593) );
  XOR U3226 ( .A(n2594), .B(n2595), .Z(n2591) );
  AND U3227 ( .A(n2596), .B(n2597), .Z(n2594) );
  XNOR U3228 ( .A(x[631]), .B(n2595), .Z(n2597) );
  XOR U3229 ( .A(n2598), .B(n2599), .Z(n2595) );
  AND U3230 ( .A(n2600), .B(n2601), .Z(n2598) );
  XNOR U3231 ( .A(x[630]), .B(n2599), .Z(n2601) );
  XOR U3232 ( .A(n2602), .B(n2603), .Z(n2599) );
  AND U3233 ( .A(n2604), .B(n2605), .Z(n2602) );
  XNOR U3234 ( .A(x[629]), .B(n2603), .Z(n2605) );
  XOR U3235 ( .A(n2606), .B(n2607), .Z(n2603) );
  AND U3236 ( .A(n2608), .B(n2609), .Z(n2606) );
  XNOR U3237 ( .A(x[628]), .B(n2607), .Z(n2609) );
  XOR U3238 ( .A(n2610), .B(n2611), .Z(n2607) );
  AND U3239 ( .A(n2612), .B(n2613), .Z(n2610) );
  XNOR U3240 ( .A(x[627]), .B(n2611), .Z(n2613) );
  XOR U3241 ( .A(n2614), .B(n2615), .Z(n2611) );
  AND U3242 ( .A(n2616), .B(n2617), .Z(n2614) );
  XNOR U3243 ( .A(x[626]), .B(n2615), .Z(n2617) );
  XOR U3244 ( .A(n2618), .B(n2619), .Z(n2615) );
  AND U3245 ( .A(n2620), .B(n2621), .Z(n2618) );
  XNOR U3246 ( .A(x[625]), .B(n2619), .Z(n2621) );
  XOR U3247 ( .A(n2622), .B(n2623), .Z(n2619) );
  AND U3248 ( .A(n2624), .B(n2625), .Z(n2622) );
  XNOR U3249 ( .A(x[624]), .B(n2623), .Z(n2625) );
  XOR U3250 ( .A(n2626), .B(n2627), .Z(n2623) );
  AND U3251 ( .A(n2628), .B(n2629), .Z(n2626) );
  XNOR U3252 ( .A(x[623]), .B(n2627), .Z(n2629) );
  XOR U3253 ( .A(n2630), .B(n2631), .Z(n2627) );
  AND U3254 ( .A(n2632), .B(n2633), .Z(n2630) );
  XNOR U3255 ( .A(x[622]), .B(n2631), .Z(n2633) );
  XOR U3256 ( .A(n2634), .B(n2635), .Z(n2631) );
  AND U3257 ( .A(n2636), .B(n2637), .Z(n2634) );
  XNOR U3258 ( .A(x[621]), .B(n2635), .Z(n2637) );
  XOR U3259 ( .A(n2638), .B(n2639), .Z(n2635) );
  AND U3260 ( .A(n2640), .B(n2641), .Z(n2638) );
  XNOR U3261 ( .A(x[620]), .B(n2639), .Z(n2641) );
  XOR U3262 ( .A(n2642), .B(n2643), .Z(n2639) );
  AND U3263 ( .A(n2644), .B(n2645), .Z(n2642) );
  XNOR U3264 ( .A(x[619]), .B(n2643), .Z(n2645) );
  XOR U3265 ( .A(n2646), .B(n2647), .Z(n2643) );
  AND U3266 ( .A(n2648), .B(n2649), .Z(n2646) );
  XNOR U3267 ( .A(x[618]), .B(n2647), .Z(n2649) );
  XOR U3268 ( .A(n2650), .B(n2651), .Z(n2647) );
  AND U3269 ( .A(n2652), .B(n2653), .Z(n2650) );
  XNOR U3270 ( .A(x[617]), .B(n2651), .Z(n2653) );
  XOR U3271 ( .A(n2654), .B(n2655), .Z(n2651) );
  AND U3272 ( .A(n2656), .B(n2657), .Z(n2654) );
  XNOR U3273 ( .A(x[616]), .B(n2655), .Z(n2657) );
  XOR U3274 ( .A(n2658), .B(n2659), .Z(n2655) );
  AND U3275 ( .A(n2660), .B(n2661), .Z(n2658) );
  XNOR U3276 ( .A(x[615]), .B(n2659), .Z(n2661) );
  XOR U3277 ( .A(n2662), .B(n2663), .Z(n2659) );
  AND U3278 ( .A(n2664), .B(n2665), .Z(n2662) );
  XNOR U3279 ( .A(x[614]), .B(n2663), .Z(n2665) );
  XOR U3280 ( .A(n2666), .B(n2667), .Z(n2663) );
  AND U3281 ( .A(n2668), .B(n2669), .Z(n2666) );
  XNOR U3282 ( .A(x[613]), .B(n2667), .Z(n2669) );
  XOR U3283 ( .A(n2670), .B(n2671), .Z(n2667) );
  AND U3284 ( .A(n2672), .B(n2673), .Z(n2670) );
  XNOR U3285 ( .A(x[612]), .B(n2671), .Z(n2673) );
  XOR U3286 ( .A(n2674), .B(n2675), .Z(n2671) );
  AND U3287 ( .A(n2676), .B(n2677), .Z(n2674) );
  XNOR U3288 ( .A(x[611]), .B(n2675), .Z(n2677) );
  XOR U3289 ( .A(n2678), .B(n2679), .Z(n2675) );
  AND U3290 ( .A(n2680), .B(n2681), .Z(n2678) );
  XNOR U3291 ( .A(x[610]), .B(n2679), .Z(n2681) );
  XOR U3292 ( .A(n2682), .B(n2683), .Z(n2679) );
  AND U3293 ( .A(n2684), .B(n2685), .Z(n2682) );
  XNOR U3294 ( .A(x[609]), .B(n2683), .Z(n2685) );
  XOR U3295 ( .A(n2686), .B(n2687), .Z(n2683) );
  AND U3296 ( .A(n2688), .B(n2689), .Z(n2686) );
  XNOR U3297 ( .A(x[608]), .B(n2687), .Z(n2689) );
  XOR U3298 ( .A(n2690), .B(n2691), .Z(n2687) );
  AND U3299 ( .A(n2692), .B(n2693), .Z(n2690) );
  XNOR U3300 ( .A(x[607]), .B(n2691), .Z(n2693) );
  XOR U3301 ( .A(n2694), .B(n2695), .Z(n2691) );
  AND U3302 ( .A(n2696), .B(n2697), .Z(n2694) );
  XNOR U3303 ( .A(x[606]), .B(n2695), .Z(n2697) );
  XOR U3304 ( .A(n2698), .B(n2699), .Z(n2695) );
  AND U3305 ( .A(n2700), .B(n2701), .Z(n2698) );
  XNOR U3306 ( .A(x[605]), .B(n2699), .Z(n2701) );
  XOR U3307 ( .A(n2702), .B(n2703), .Z(n2699) );
  AND U3308 ( .A(n2704), .B(n2705), .Z(n2702) );
  XNOR U3309 ( .A(x[604]), .B(n2703), .Z(n2705) );
  XOR U3310 ( .A(n2706), .B(n2707), .Z(n2703) );
  AND U3311 ( .A(n2708), .B(n2709), .Z(n2706) );
  XNOR U3312 ( .A(x[603]), .B(n2707), .Z(n2709) );
  XOR U3313 ( .A(n2710), .B(n2711), .Z(n2707) );
  AND U3314 ( .A(n2712), .B(n2713), .Z(n2710) );
  XNOR U3315 ( .A(x[602]), .B(n2711), .Z(n2713) );
  XOR U3316 ( .A(n2714), .B(n2715), .Z(n2711) );
  AND U3317 ( .A(n2716), .B(n2717), .Z(n2714) );
  XNOR U3318 ( .A(x[601]), .B(n2715), .Z(n2717) );
  XOR U3319 ( .A(n2718), .B(n2719), .Z(n2715) );
  AND U3320 ( .A(n2720), .B(n2721), .Z(n2718) );
  XNOR U3321 ( .A(x[600]), .B(n2719), .Z(n2721) );
  XOR U3322 ( .A(n2722), .B(n2723), .Z(n2719) );
  AND U3323 ( .A(n2724), .B(n2725), .Z(n2722) );
  XNOR U3324 ( .A(x[599]), .B(n2723), .Z(n2725) );
  XOR U3325 ( .A(n2726), .B(n2727), .Z(n2723) );
  AND U3326 ( .A(n2728), .B(n2729), .Z(n2726) );
  XNOR U3327 ( .A(x[598]), .B(n2727), .Z(n2729) );
  XOR U3328 ( .A(n2730), .B(n2731), .Z(n2727) );
  AND U3329 ( .A(n2732), .B(n2733), .Z(n2730) );
  XNOR U3330 ( .A(x[597]), .B(n2731), .Z(n2733) );
  XOR U3331 ( .A(n2734), .B(n2735), .Z(n2731) );
  AND U3332 ( .A(n2736), .B(n2737), .Z(n2734) );
  XNOR U3333 ( .A(x[596]), .B(n2735), .Z(n2737) );
  XOR U3334 ( .A(n2738), .B(n2739), .Z(n2735) );
  AND U3335 ( .A(n2740), .B(n2741), .Z(n2738) );
  XNOR U3336 ( .A(x[595]), .B(n2739), .Z(n2741) );
  XOR U3337 ( .A(n2742), .B(n2743), .Z(n2739) );
  AND U3338 ( .A(n2744), .B(n2745), .Z(n2742) );
  XNOR U3339 ( .A(x[594]), .B(n2743), .Z(n2745) );
  XOR U3340 ( .A(n2746), .B(n2747), .Z(n2743) );
  AND U3341 ( .A(n2748), .B(n2749), .Z(n2746) );
  XNOR U3342 ( .A(x[593]), .B(n2747), .Z(n2749) );
  XOR U3343 ( .A(n2750), .B(n2751), .Z(n2747) );
  AND U3344 ( .A(n2752), .B(n2753), .Z(n2750) );
  XNOR U3345 ( .A(x[592]), .B(n2751), .Z(n2753) );
  XOR U3346 ( .A(n2754), .B(n2755), .Z(n2751) );
  AND U3347 ( .A(n2756), .B(n2757), .Z(n2754) );
  XNOR U3348 ( .A(x[591]), .B(n2755), .Z(n2757) );
  XOR U3349 ( .A(n2758), .B(n2759), .Z(n2755) );
  AND U3350 ( .A(n2760), .B(n2761), .Z(n2758) );
  XNOR U3351 ( .A(x[590]), .B(n2759), .Z(n2761) );
  XOR U3352 ( .A(n2762), .B(n2763), .Z(n2759) );
  AND U3353 ( .A(n2764), .B(n2765), .Z(n2762) );
  XNOR U3354 ( .A(x[589]), .B(n2763), .Z(n2765) );
  XOR U3355 ( .A(n2766), .B(n2767), .Z(n2763) );
  AND U3356 ( .A(n2768), .B(n2769), .Z(n2766) );
  XNOR U3357 ( .A(x[588]), .B(n2767), .Z(n2769) );
  XOR U3358 ( .A(n2770), .B(n2771), .Z(n2767) );
  AND U3359 ( .A(n2772), .B(n2773), .Z(n2770) );
  XNOR U3360 ( .A(x[587]), .B(n2771), .Z(n2773) );
  XOR U3361 ( .A(n2774), .B(n2775), .Z(n2771) );
  AND U3362 ( .A(n2776), .B(n2777), .Z(n2774) );
  XNOR U3363 ( .A(x[586]), .B(n2775), .Z(n2777) );
  XOR U3364 ( .A(n2778), .B(n2779), .Z(n2775) );
  AND U3365 ( .A(n2780), .B(n2781), .Z(n2778) );
  XNOR U3366 ( .A(x[585]), .B(n2779), .Z(n2781) );
  XOR U3367 ( .A(n2782), .B(n2783), .Z(n2779) );
  AND U3368 ( .A(n2784), .B(n2785), .Z(n2782) );
  XNOR U3369 ( .A(x[584]), .B(n2783), .Z(n2785) );
  XOR U3370 ( .A(n2786), .B(n2787), .Z(n2783) );
  AND U3371 ( .A(n2788), .B(n2789), .Z(n2786) );
  XNOR U3372 ( .A(x[583]), .B(n2787), .Z(n2789) );
  XOR U3373 ( .A(n2790), .B(n2791), .Z(n2787) );
  AND U3374 ( .A(n2792), .B(n2793), .Z(n2790) );
  XNOR U3375 ( .A(x[582]), .B(n2791), .Z(n2793) );
  XOR U3376 ( .A(n2794), .B(n2795), .Z(n2791) );
  AND U3377 ( .A(n2796), .B(n2797), .Z(n2794) );
  XNOR U3378 ( .A(x[581]), .B(n2795), .Z(n2797) );
  XOR U3379 ( .A(n2798), .B(n2799), .Z(n2795) );
  AND U3380 ( .A(n2800), .B(n2801), .Z(n2798) );
  XNOR U3381 ( .A(x[580]), .B(n2799), .Z(n2801) );
  XOR U3382 ( .A(n2802), .B(n2803), .Z(n2799) );
  AND U3383 ( .A(n2804), .B(n2805), .Z(n2802) );
  XNOR U3384 ( .A(x[579]), .B(n2803), .Z(n2805) );
  XOR U3385 ( .A(n2806), .B(n2807), .Z(n2803) );
  AND U3386 ( .A(n2808), .B(n2809), .Z(n2806) );
  XNOR U3387 ( .A(x[578]), .B(n2807), .Z(n2809) );
  XOR U3388 ( .A(n2810), .B(n2811), .Z(n2807) );
  AND U3389 ( .A(n2812), .B(n2813), .Z(n2810) );
  XNOR U3390 ( .A(x[577]), .B(n2811), .Z(n2813) );
  XOR U3391 ( .A(n2814), .B(n2815), .Z(n2811) );
  AND U3392 ( .A(n2816), .B(n2817), .Z(n2814) );
  XNOR U3393 ( .A(x[576]), .B(n2815), .Z(n2817) );
  XOR U3394 ( .A(n2818), .B(n2819), .Z(n2815) );
  AND U3395 ( .A(n2820), .B(n2821), .Z(n2818) );
  XNOR U3396 ( .A(x[575]), .B(n2819), .Z(n2821) );
  XOR U3397 ( .A(n2822), .B(n2823), .Z(n2819) );
  AND U3398 ( .A(n2824), .B(n2825), .Z(n2822) );
  XNOR U3399 ( .A(x[574]), .B(n2823), .Z(n2825) );
  XOR U3400 ( .A(n2826), .B(n2827), .Z(n2823) );
  AND U3401 ( .A(n2828), .B(n2829), .Z(n2826) );
  XNOR U3402 ( .A(x[573]), .B(n2827), .Z(n2829) );
  XOR U3403 ( .A(n2830), .B(n2831), .Z(n2827) );
  AND U3404 ( .A(n2832), .B(n2833), .Z(n2830) );
  XNOR U3405 ( .A(x[572]), .B(n2831), .Z(n2833) );
  XOR U3406 ( .A(n2834), .B(n2835), .Z(n2831) );
  AND U3407 ( .A(n2836), .B(n2837), .Z(n2834) );
  XNOR U3408 ( .A(x[571]), .B(n2835), .Z(n2837) );
  XOR U3409 ( .A(n2838), .B(n2839), .Z(n2835) );
  AND U3410 ( .A(n2840), .B(n2841), .Z(n2838) );
  XNOR U3411 ( .A(x[570]), .B(n2839), .Z(n2841) );
  XOR U3412 ( .A(n2842), .B(n2843), .Z(n2839) );
  AND U3413 ( .A(n2844), .B(n2845), .Z(n2842) );
  XNOR U3414 ( .A(x[569]), .B(n2843), .Z(n2845) );
  XOR U3415 ( .A(n2846), .B(n2847), .Z(n2843) );
  AND U3416 ( .A(n2848), .B(n2849), .Z(n2846) );
  XNOR U3417 ( .A(x[568]), .B(n2847), .Z(n2849) );
  XOR U3418 ( .A(n2850), .B(n2851), .Z(n2847) );
  AND U3419 ( .A(n2852), .B(n2853), .Z(n2850) );
  XNOR U3420 ( .A(x[567]), .B(n2851), .Z(n2853) );
  XOR U3421 ( .A(n2854), .B(n2855), .Z(n2851) );
  AND U3422 ( .A(n2856), .B(n2857), .Z(n2854) );
  XNOR U3423 ( .A(x[566]), .B(n2855), .Z(n2857) );
  XOR U3424 ( .A(n2858), .B(n2859), .Z(n2855) );
  AND U3425 ( .A(n2860), .B(n2861), .Z(n2858) );
  XNOR U3426 ( .A(x[565]), .B(n2859), .Z(n2861) );
  XOR U3427 ( .A(n2862), .B(n2863), .Z(n2859) );
  AND U3428 ( .A(n2864), .B(n2865), .Z(n2862) );
  XNOR U3429 ( .A(x[564]), .B(n2863), .Z(n2865) );
  XOR U3430 ( .A(n2866), .B(n2867), .Z(n2863) );
  AND U3431 ( .A(n2868), .B(n2869), .Z(n2866) );
  XNOR U3432 ( .A(x[563]), .B(n2867), .Z(n2869) );
  XOR U3433 ( .A(n2870), .B(n2871), .Z(n2867) );
  AND U3434 ( .A(n2872), .B(n2873), .Z(n2870) );
  XNOR U3435 ( .A(x[562]), .B(n2871), .Z(n2873) );
  XOR U3436 ( .A(n2874), .B(n2875), .Z(n2871) );
  AND U3437 ( .A(n2876), .B(n2877), .Z(n2874) );
  XNOR U3438 ( .A(x[561]), .B(n2875), .Z(n2877) );
  XOR U3439 ( .A(n2878), .B(n2879), .Z(n2875) );
  AND U3440 ( .A(n2880), .B(n2881), .Z(n2878) );
  XNOR U3441 ( .A(x[560]), .B(n2879), .Z(n2881) );
  XOR U3442 ( .A(n2882), .B(n2883), .Z(n2879) );
  AND U3443 ( .A(n2884), .B(n2885), .Z(n2882) );
  XNOR U3444 ( .A(x[559]), .B(n2883), .Z(n2885) );
  XOR U3445 ( .A(n2886), .B(n2887), .Z(n2883) );
  AND U3446 ( .A(n2888), .B(n2889), .Z(n2886) );
  XNOR U3447 ( .A(x[558]), .B(n2887), .Z(n2889) );
  XOR U3448 ( .A(n2890), .B(n2891), .Z(n2887) );
  AND U3449 ( .A(n2892), .B(n2893), .Z(n2890) );
  XNOR U3450 ( .A(x[557]), .B(n2891), .Z(n2893) );
  XOR U3451 ( .A(n2894), .B(n2895), .Z(n2891) );
  AND U3452 ( .A(n2896), .B(n2897), .Z(n2894) );
  XNOR U3453 ( .A(x[556]), .B(n2895), .Z(n2897) );
  XOR U3454 ( .A(n2898), .B(n2899), .Z(n2895) );
  AND U3455 ( .A(n2900), .B(n2901), .Z(n2898) );
  XNOR U3456 ( .A(x[555]), .B(n2899), .Z(n2901) );
  XOR U3457 ( .A(n2902), .B(n2903), .Z(n2899) );
  AND U3458 ( .A(n2904), .B(n2905), .Z(n2902) );
  XNOR U3459 ( .A(x[554]), .B(n2903), .Z(n2905) );
  XOR U3460 ( .A(n2906), .B(n2907), .Z(n2903) );
  AND U3461 ( .A(n2908), .B(n2909), .Z(n2906) );
  XNOR U3462 ( .A(x[553]), .B(n2907), .Z(n2909) );
  XOR U3463 ( .A(n2910), .B(n2911), .Z(n2907) );
  AND U3464 ( .A(n2912), .B(n2913), .Z(n2910) );
  XNOR U3465 ( .A(x[552]), .B(n2911), .Z(n2913) );
  XOR U3466 ( .A(n2914), .B(n2915), .Z(n2911) );
  AND U3467 ( .A(n2916), .B(n2917), .Z(n2914) );
  XNOR U3468 ( .A(x[551]), .B(n2915), .Z(n2917) );
  XOR U3469 ( .A(n2918), .B(n2919), .Z(n2915) );
  AND U3470 ( .A(n2920), .B(n2921), .Z(n2918) );
  XNOR U3471 ( .A(x[550]), .B(n2919), .Z(n2921) );
  XOR U3472 ( .A(n2922), .B(n2923), .Z(n2919) );
  AND U3473 ( .A(n2924), .B(n2925), .Z(n2922) );
  XNOR U3474 ( .A(x[549]), .B(n2923), .Z(n2925) );
  XOR U3475 ( .A(n2926), .B(n2927), .Z(n2923) );
  AND U3476 ( .A(n2928), .B(n2929), .Z(n2926) );
  XNOR U3477 ( .A(x[548]), .B(n2927), .Z(n2929) );
  XOR U3478 ( .A(n2930), .B(n2931), .Z(n2927) );
  AND U3479 ( .A(n2932), .B(n2933), .Z(n2930) );
  XNOR U3480 ( .A(x[547]), .B(n2931), .Z(n2933) );
  XOR U3481 ( .A(n2934), .B(n2935), .Z(n2931) );
  AND U3482 ( .A(n2936), .B(n2937), .Z(n2934) );
  XNOR U3483 ( .A(x[546]), .B(n2935), .Z(n2937) );
  XOR U3484 ( .A(n2938), .B(n2939), .Z(n2935) );
  AND U3485 ( .A(n2940), .B(n2941), .Z(n2938) );
  XNOR U3486 ( .A(x[545]), .B(n2939), .Z(n2941) );
  XOR U3487 ( .A(n2942), .B(n2943), .Z(n2939) );
  AND U3488 ( .A(n2944), .B(n2945), .Z(n2942) );
  XNOR U3489 ( .A(x[544]), .B(n2943), .Z(n2945) );
  XOR U3490 ( .A(n2946), .B(n2947), .Z(n2943) );
  AND U3491 ( .A(n2948), .B(n2949), .Z(n2946) );
  XNOR U3492 ( .A(x[543]), .B(n2947), .Z(n2949) );
  XOR U3493 ( .A(n2950), .B(n2951), .Z(n2947) );
  AND U3494 ( .A(n2952), .B(n2953), .Z(n2950) );
  XNOR U3495 ( .A(x[542]), .B(n2951), .Z(n2953) );
  XOR U3496 ( .A(n2954), .B(n2955), .Z(n2951) );
  AND U3497 ( .A(n2956), .B(n2957), .Z(n2954) );
  XNOR U3498 ( .A(x[541]), .B(n2955), .Z(n2957) );
  XOR U3499 ( .A(n2958), .B(n2959), .Z(n2955) );
  AND U3500 ( .A(n2960), .B(n2961), .Z(n2958) );
  XNOR U3501 ( .A(x[540]), .B(n2959), .Z(n2961) );
  XOR U3502 ( .A(n2962), .B(n2963), .Z(n2959) );
  AND U3503 ( .A(n2964), .B(n2965), .Z(n2962) );
  XNOR U3504 ( .A(x[539]), .B(n2963), .Z(n2965) );
  XOR U3505 ( .A(n2966), .B(n2967), .Z(n2963) );
  AND U3506 ( .A(n2968), .B(n2969), .Z(n2966) );
  XNOR U3507 ( .A(x[538]), .B(n2967), .Z(n2969) );
  XOR U3508 ( .A(n2970), .B(n2971), .Z(n2967) );
  AND U3509 ( .A(n2972), .B(n2973), .Z(n2970) );
  XNOR U3510 ( .A(x[537]), .B(n2971), .Z(n2973) );
  XOR U3511 ( .A(n2974), .B(n2975), .Z(n2971) );
  AND U3512 ( .A(n2976), .B(n2977), .Z(n2974) );
  XNOR U3513 ( .A(x[536]), .B(n2975), .Z(n2977) );
  XOR U3514 ( .A(n2978), .B(n2979), .Z(n2975) );
  AND U3515 ( .A(n2980), .B(n2981), .Z(n2978) );
  XNOR U3516 ( .A(x[535]), .B(n2979), .Z(n2981) );
  XOR U3517 ( .A(n2982), .B(n2983), .Z(n2979) );
  AND U3518 ( .A(n2984), .B(n2985), .Z(n2982) );
  XNOR U3519 ( .A(x[534]), .B(n2983), .Z(n2985) );
  XOR U3520 ( .A(n2986), .B(n2987), .Z(n2983) );
  AND U3521 ( .A(n2988), .B(n2989), .Z(n2986) );
  XNOR U3522 ( .A(x[533]), .B(n2987), .Z(n2989) );
  XOR U3523 ( .A(n2990), .B(n2991), .Z(n2987) );
  AND U3524 ( .A(n2992), .B(n2993), .Z(n2990) );
  XNOR U3525 ( .A(x[532]), .B(n2991), .Z(n2993) );
  XOR U3526 ( .A(n2994), .B(n2995), .Z(n2991) );
  AND U3527 ( .A(n2996), .B(n2997), .Z(n2994) );
  XNOR U3528 ( .A(x[531]), .B(n2995), .Z(n2997) );
  XOR U3529 ( .A(n2998), .B(n2999), .Z(n2995) );
  AND U3530 ( .A(n3000), .B(n3001), .Z(n2998) );
  XNOR U3531 ( .A(x[530]), .B(n2999), .Z(n3001) );
  XOR U3532 ( .A(n3002), .B(n3003), .Z(n2999) );
  AND U3533 ( .A(n3004), .B(n3005), .Z(n3002) );
  XNOR U3534 ( .A(x[529]), .B(n3003), .Z(n3005) );
  XOR U3535 ( .A(n3006), .B(n3007), .Z(n3003) );
  AND U3536 ( .A(n3008), .B(n3009), .Z(n3006) );
  XNOR U3537 ( .A(x[528]), .B(n3007), .Z(n3009) );
  XOR U3538 ( .A(n3010), .B(n3011), .Z(n3007) );
  AND U3539 ( .A(n3012), .B(n3013), .Z(n3010) );
  XNOR U3540 ( .A(x[527]), .B(n3011), .Z(n3013) );
  XOR U3541 ( .A(n3014), .B(n3015), .Z(n3011) );
  AND U3542 ( .A(n3016), .B(n3017), .Z(n3014) );
  XNOR U3543 ( .A(x[526]), .B(n3015), .Z(n3017) );
  XOR U3544 ( .A(n3018), .B(n3019), .Z(n3015) );
  AND U3545 ( .A(n3020), .B(n3021), .Z(n3018) );
  XNOR U3546 ( .A(x[525]), .B(n3019), .Z(n3021) );
  XOR U3547 ( .A(n3022), .B(n3023), .Z(n3019) );
  AND U3548 ( .A(n3024), .B(n3025), .Z(n3022) );
  XNOR U3549 ( .A(x[524]), .B(n3023), .Z(n3025) );
  XOR U3550 ( .A(n3026), .B(n3027), .Z(n3023) );
  AND U3551 ( .A(n3028), .B(n3029), .Z(n3026) );
  XNOR U3552 ( .A(x[523]), .B(n3027), .Z(n3029) );
  XOR U3553 ( .A(n3030), .B(n3031), .Z(n3027) );
  AND U3554 ( .A(n3032), .B(n3033), .Z(n3030) );
  XNOR U3555 ( .A(x[522]), .B(n3031), .Z(n3033) );
  XOR U3556 ( .A(n3034), .B(n3035), .Z(n3031) );
  AND U3557 ( .A(n3036), .B(n3037), .Z(n3034) );
  XNOR U3558 ( .A(x[521]), .B(n3035), .Z(n3037) );
  XOR U3559 ( .A(n3038), .B(n3039), .Z(n3035) );
  AND U3560 ( .A(n3040), .B(n3041), .Z(n3038) );
  XNOR U3561 ( .A(x[520]), .B(n3039), .Z(n3041) );
  XOR U3562 ( .A(n3042), .B(n3043), .Z(n3039) );
  AND U3563 ( .A(n3044), .B(n3045), .Z(n3042) );
  XNOR U3564 ( .A(x[519]), .B(n3043), .Z(n3045) );
  XOR U3565 ( .A(n3046), .B(n3047), .Z(n3043) );
  AND U3566 ( .A(n3048), .B(n3049), .Z(n3046) );
  XNOR U3567 ( .A(x[518]), .B(n3047), .Z(n3049) );
  XOR U3568 ( .A(n3050), .B(n3051), .Z(n3047) );
  AND U3569 ( .A(n3052), .B(n3053), .Z(n3050) );
  XNOR U3570 ( .A(x[517]), .B(n3051), .Z(n3053) );
  XOR U3571 ( .A(n3054), .B(n3055), .Z(n3051) );
  AND U3572 ( .A(n3056), .B(n3057), .Z(n3054) );
  XNOR U3573 ( .A(x[516]), .B(n3055), .Z(n3057) );
  XOR U3574 ( .A(n3058), .B(n3059), .Z(n3055) );
  AND U3575 ( .A(n3060), .B(n3061), .Z(n3058) );
  XNOR U3576 ( .A(x[515]), .B(n3059), .Z(n3061) );
  XOR U3577 ( .A(n3062), .B(n3063), .Z(n3059) );
  AND U3578 ( .A(n3064), .B(n3065), .Z(n3062) );
  XNOR U3579 ( .A(x[514]), .B(n3063), .Z(n3065) );
  XOR U3580 ( .A(n3066), .B(n3067), .Z(n3063) );
  AND U3581 ( .A(n3068), .B(n3069), .Z(n3066) );
  XNOR U3582 ( .A(x[513]), .B(n3067), .Z(n3069) );
  XOR U3583 ( .A(n3070), .B(n3071), .Z(n3067) );
  AND U3584 ( .A(n3072), .B(n3073), .Z(n3070) );
  XNOR U3585 ( .A(x[512]), .B(n3071), .Z(n3073) );
  XOR U3586 ( .A(n3074), .B(n3075), .Z(n3071) );
  AND U3587 ( .A(n3076), .B(n3077), .Z(n3074) );
  XNOR U3588 ( .A(x[511]), .B(n3075), .Z(n3077) );
  XOR U3589 ( .A(n3078), .B(n3079), .Z(n3075) );
  AND U3590 ( .A(n3080), .B(n3081), .Z(n3078) );
  XNOR U3591 ( .A(x[510]), .B(n3079), .Z(n3081) );
  XOR U3592 ( .A(n3082), .B(n3083), .Z(n3079) );
  AND U3593 ( .A(n3084), .B(n3085), .Z(n3082) );
  XNOR U3594 ( .A(x[509]), .B(n3083), .Z(n3085) );
  XOR U3595 ( .A(n3086), .B(n3087), .Z(n3083) );
  AND U3596 ( .A(n3088), .B(n3089), .Z(n3086) );
  XNOR U3597 ( .A(x[508]), .B(n3087), .Z(n3089) );
  XOR U3598 ( .A(n3090), .B(n3091), .Z(n3087) );
  AND U3599 ( .A(n3092), .B(n3093), .Z(n3090) );
  XNOR U3600 ( .A(x[507]), .B(n3091), .Z(n3093) );
  XOR U3601 ( .A(n3094), .B(n3095), .Z(n3091) );
  AND U3602 ( .A(n3096), .B(n3097), .Z(n3094) );
  XNOR U3603 ( .A(x[506]), .B(n3095), .Z(n3097) );
  XOR U3604 ( .A(n3098), .B(n3099), .Z(n3095) );
  AND U3605 ( .A(n3100), .B(n3101), .Z(n3098) );
  XNOR U3606 ( .A(x[505]), .B(n3099), .Z(n3101) );
  XOR U3607 ( .A(n3102), .B(n3103), .Z(n3099) );
  AND U3608 ( .A(n3104), .B(n3105), .Z(n3102) );
  XNOR U3609 ( .A(x[504]), .B(n3103), .Z(n3105) );
  XOR U3610 ( .A(n3106), .B(n3107), .Z(n3103) );
  AND U3611 ( .A(n3108), .B(n3109), .Z(n3106) );
  XNOR U3612 ( .A(x[503]), .B(n3107), .Z(n3109) );
  XOR U3613 ( .A(n3110), .B(n3111), .Z(n3107) );
  AND U3614 ( .A(n3112), .B(n3113), .Z(n3110) );
  XNOR U3615 ( .A(x[502]), .B(n3111), .Z(n3113) );
  XOR U3616 ( .A(n3114), .B(n3115), .Z(n3111) );
  AND U3617 ( .A(n3116), .B(n3117), .Z(n3114) );
  XNOR U3618 ( .A(x[501]), .B(n3115), .Z(n3117) );
  XOR U3619 ( .A(n3118), .B(n3119), .Z(n3115) );
  AND U3620 ( .A(n3120), .B(n3121), .Z(n3118) );
  XNOR U3621 ( .A(x[500]), .B(n3119), .Z(n3121) );
  XOR U3622 ( .A(n3122), .B(n3123), .Z(n3119) );
  AND U3623 ( .A(n3124), .B(n3125), .Z(n3122) );
  XNOR U3624 ( .A(x[499]), .B(n3123), .Z(n3125) );
  XOR U3625 ( .A(n3126), .B(n3127), .Z(n3123) );
  AND U3626 ( .A(n3128), .B(n3129), .Z(n3126) );
  XNOR U3627 ( .A(x[498]), .B(n3127), .Z(n3129) );
  XOR U3628 ( .A(n3130), .B(n3131), .Z(n3127) );
  AND U3629 ( .A(n3132), .B(n3133), .Z(n3130) );
  XNOR U3630 ( .A(x[497]), .B(n3131), .Z(n3133) );
  XOR U3631 ( .A(n3134), .B(n3135), .Z(n3131) );
  AND U3632 ( .A(n3136), .B(n3137), .Z(n3134) );
  XNOR U3633 ( .A(x[496]), .B(n3135), .Z(n3137) );
  XOR U3634 ( .A(n3138), .B(n3139), .Z(n3135) );
  AND U3635 ( .A(n3140), .B(n3141), .Z(n3138) );
  XNOR U3636 ( .A(x[495]), .B(n3139), .Z(n3141) );
  XOR U3637 ( .A(n3142), .B(n3143), .Z(n3139) );
  AND U3638 ( .A(n3144), .B(n3145), .Z(n3142) );
  XNOR U3639 ( .A(x[494]), .B(n3143), .Z(n3145) );
  XOR U3640 ( .A(n3146), .B(n3147), .Z(n3143) );
  AND U3641 ( .A(n3148), .B(n3149), .Z(n3146) );
  XNOR U3642 ( .A(x[493]), .B(n3147), .Z(n3149) );
  XOR U3643 ( .A(n3150), .B(n3151), .Z(n3147) );
  AND U3644 ( .A(n3152), .B(n3153), .Z(n3150) );
  XNOR U3645 ( .A(x[492]), .B(n3151), .Z(n3153) );
  XOR U3646 ( .A(n3154), .B(n3155), .Z(n3151) );
  AND U3647 ( .A(n3156), .B(n3157), .Z(n3154) );
  XNOR U3648 ( .A(x[491]), .B(n3155), .Z(n3157) );
  XOR U3649 ( .A(n3158), .B(n3159), .Z(n3155) );
  AND U3650 ( .A(n3160), .B(n3161), .Z(n3158) );
  XNOR U3651 ( .A(x[490]), .B(n3159), .Z(n3161) );
  XOR U3652 ( .A(n3162), .B(n3163), .Z(n3159) );
  AND U3653 ( .A(n3164), .B(n3165), .Z(n3162) );
  XNOR U3654 ( .A(x[489]), .B(n3163), .Z(n3165) );
  XOR U3655 ( .A(n3166), .B(n3167), .Z(n3163) );
  AND U3656 ( .A(n3168), .B(n3169), .Z(n3166) );
  XNOR U3657 ( .A(x[488]), .B(n3167), .Z(n3169) );
  XOR U3658 ( .A(n3170), .B(n3171), .Z(n3167) );
  AND U3659 ( .A(n3172), .B(n3173), .Z(n3170) );
  XNOR U3660 ( .A(x[487]), .B(n3171), .Z(n3173) );
  XOR U3661 ( .A(n3174), .B(n3175), .Z(n3171) );
  AND U3662 ( .A(n3176), .B(n3177), .Z(n3174) );
  XNOR U3663 ( .A(x[486]), .B(n3175), .Z(n3177) );
  XOR U3664 ( .A(n3178), .B(n3179), .Z(n3175) );
  AND U3665 ( .A(n3180), .B(n3181), .Z(n3178) );
  XNOR U3666 ( .A(x[485]), .B(n3179), .Z(n3181) );
  XOR U3667 ( .A(n3182), .B(n3183), .Z(n3179) );
  AND U3668 ( .A(n3184), .B(n3185), .Z(n3182) );
  XNOR U3669 ( .A(x[484]), .B(n3183), .Z(n3185) );
  XOR U3670 ( .A(n3186), .B(n3187), .Z(n3183) );
  AND U3671 ( .A(n3188), .B(n3189), .Z(n3186) );
  XNOR U3672 ( .A(x[483]), .B(n3187), .Z(n3189) );
  XOR U3673 ( .A(n3190), .B(n3191), .Z(n3187) );
  AND U3674 ( .A(n3192), .B(n3193), .Z(n3190) );
  XNOR U3675 ( .A(x[482]), .B(n3191), .Z(n3193) );
  XOR U3676 ( .A(n3194), .B(n3195), .Z(n3191) );
  AND U3677 ( .A(n3196), .B(n3197), .Z(n3194) );
  XNOR U3678 ( .A(x[481]), .B(n3195), .Z(n3197) );
  XOR U3679 ( .A(n3198), .B(n3199), .Z(n3195) );
  AND U3680 ( .A(n3200), .B(n3201), .Z(n3198) );
  XNOR U3681 ( .A(x[480]), .B(n3199), .Z(n3201) );
  XOR U3682 ( .A(n3202), .B(n3203), .Z(n3199) );
  AND U3683 ( .A(n3204), .B(n3205), .Z(n3202) );
  XNOR U3684 ( .A(x[479]), .B(n3203), .Z(n3205) );
  XOR U3685 ( .A(n3206), .B(n3207), .Z(n3203) );
  AND U3686 ( .A(n3208), .B(n3209), .Z(n3206) );
  XNOR U3687 ( .A(x[478]), .B(n3207), .Z(n3209) );
  XOR U3688 ( .A(n3210), .B(n3211), .Z(n3207) );
  AND U3689 ( .A(n3212), .B(n3213), .Z(n3210) );
  XNOR U3690 ( .A(x[477]), .B(n3211), .Z(n3213) );
  XOR U3691 ( .A(n3214), .B(n3215), .Z(n3211) );
  AND U3692 ( .A(n3216), .B(n3217), .Z(n3214) );
  XNOR U3693 ( .A(x[476]), .B(n3215), .Z(n3217) );
  XOR U3694 ( .A(n3218), .B(n3219), .Z(n3215) );
  AND U3695 ( .A(n3220), .B(n3221), .Z(n3218) );
  XNOR U3696 ( .A(x[475]), .B(n3219), .Z(n3221) );
  XOR U3697 ( .A(n3222), .B(n3223), .Z(n3219) );
  AND U3698 ( .A(n3224), .B(n3225), .Z(n3222) );
  XNOR U3699 ( .A(x[474]), .B(n3223), .Z(n3225) );
  XOR U3700 ( .A(n3226), .B(n3227), .Z(n3223) );
  AND U3701 ( .A(n3228), .B(n3229), .Z(n3226) );
  XNOR U3702 ( .A(x[473]), .B(n3227), .Z(n3229) );
  XOR U3703 ( .A(n3230), .B(n3231), .Z(n3227) );
  AND U3704 ( .A(n3232), .B(n3233), .Z(n3230) );
  XNOR U3705 ( .A(x[472]), .B(n3231), .Z(n3233) );
  XOR U3706 ( .A(n3234), .B(n3235), .Z(n3231) );
  AND U3707 ( .A(n3236), .B(n3237), .Z(n3234) );
  XNOR U3708 ( .A(x[471]), .B(n3235), .Z(n3237) );
  XOR U3709 ( .A(n3238), .B(n3239), .Z(n3235) );
  AND U3710 ( .A(n3240), .B(n3241), .Z(n3238) );
  XNOR U3711 ( .A(x[470]), .B(n3239), .Z(n3241) );
  XOR U3712 ( .A(n3242), .B(n3243), .Z(n3239) );
  AND U3713 ( .A(n3244), .B(n3245), .Z(n3242) );
  XNOR U3714 ( .A(x[469]), .B(n3243), .Z(n3245) );
  XOR U3715 ( .A(n3246), .B(n3247), .Z(n3243) );
  AND U3716 ( .A(n3248), .B(n3249), .Z(n3246) );
  XNOR U3717 ( .A(x[468]), .B(n3247), .Z(n3249) );
  XOR U3718 ( .A(n3250), .B(n3251), .Z(n3247) );
  AND U3719 ( .A(n3252), .B(n3253), .Z(n3250) );
  XNOR U3720 ( .A(x[467]), .B(n3251), .Z(n3253) );
  XOR U3721 ( .A(n3254), .B(n3255), .Z(n3251) );
  AND U3722 ( .A(n3256), .B(n3257), .Z(n3254) );
  XNOR U3723 ( .A(x[466]), .B(n3255), .Z(n3257) );
  XOR U3724 ( .A(n3258), .B(n3259), .Z(n3255) );
  AND U3725 ( .A(n3260), .B(n3261), .Z(n3258) );
  XNOR U3726 ( .A(x[465]), .B(n3259), .Z(n3261) );
  XOR U3727 ( .A(n3262), .B(n3263), .Z(n3259) );
  AND U3728 ( .A(n3264), .B(n3265), .Z(n3262) );
  XNOR U3729 ( .A(x[464]), .B(n3263), .Z(n3265) );
  XOR U3730 ( .A(n3266), .B(n3267), .Z(n3263) );
  AND U3731 ( .A(n3268), .B(n3269), .Z(n3266) );
  XNOR U3732 ( .A(x[463]), .B(n3267), .Z(n3269) );
  XOR U3733 ( .A(n3270), .B(n3271), .Z(n3267) );
  AND U3734 ( .A(n3272), .B(n3273), .Z(n3270) );
  XNOR U3735 ( .A(x[462]), .B(n3271), .Z(n3273) );
  XOR U3736 ( .A(n3274), .B(n3275), .Z(n3271) );
  AND U3737 ( .A(n3276), .B(n3277), .Z(n3274) );
  XNOR U3738 ( .A(x[461]), .B(n3275), .Z(n3277) );
  XOR U3739 ( .A(n3278), .B(n3279), .Z(n3275) );
  AND U3740 ( .A(n3280), .B(n3281), .Z(n3278) );
  XNOR U3741 ( .A(x[460]), .B(n3279), .Z(n3281) );
  XOR U3742 ( .A(n3282), .B(n3283), .Z(n3279) );
  AND U3743 ( .A(n3284), .B(n3285), .Z(n3282) );
  XNOR U3744 ( .A(x[459]), .B(n3283), .Z(n3285) );
  XOR U3745 ( .A(n3286), .B(n3287), .Z(n3283) );
  AND U3746 ( .A(n3288), .B(n3289), .Z(n3286) );
  XNOR U3747 ( .A(x[458]), .B(n3287), .Z(n3289) );
  XOR U3748 ( .A(n3290), .B(n3291), .Z(n3287) );
  AND U3749 ( .A(n3292), .B(n3293), .Z(n3290) );
  XNOR U3750 ( .A(x[457]), .B(n3291), .Z(n3293) );
  XOR U3751 ( .A(n3294), .B(n3295), .Z(n3291) );
  AND U3752 ( .A(n3296), .B(n3297), .Z(n3294) );
  XNOR U3753 ( .A(x[456]), .B(n3295), .Z(n3297) );
  XOR U3754 ( .A(n3298), .B(n3299), .Z(n3295) );
  AND U3755 ( .A(n3300), .B(n3301), .Z(n3298) );
  XNOR U3756 ( .A(x[455]), .B(n3299), .Z(n3301) );
  XOR U3757 ( .A(n3302), .B(n3303), .Z(n3299) );
  AND U3758 ( .A(n3304), .B(n3305), .Z(n3302) );
  XNOR U3759 ( .A(x[454]), .B(n3303), .Z(n3305) );
  XOR U3760 ( .A(n3306), .B(n3307), .Z(n3303) );
  AND U3761 ( .A(n3308), .B(n3309), .Z(n3306) );
  XNOR U3762 ( .A(x[453]), .B(n3307), .Z(n3309) );
  XOR U3763 ( .A(n3310), .B(n3311), .Z(n3307) );
  AND U3764 ( .A(n3312), .B(n3313), .Z(n3310) );
  XNOR U3765 ( .A(x[452]), .B(n3311), .Z(n3313) );
  XOR U3766 ( .A(n3314), .B(n3315), .Z(n3311) );
  AND U3767 ( .A(n3316), .B(n3317), .Z(n3314) );
  XNOR U3768 ( .A(x[451]), .B(n3315), .Z(n3317) );
  XOR U3769 ( .A(n3318), .B(n3319), .Z(n3315) );
  AND U3770 ( .A(n3320), .B(n3321), .Z(n3318) );
  XNOR U3771 ( .A(x[450]), .B(n3319), .Z(n3321) );
  XOR U3772 ( .A(n3322), .B(n3323), .Z(n3319) );
  AND U3773 ( .A(n3324), .B(n3325), .Z(n3322) );
  XNOR U3774 ( .A(x[449]), .B(n3323), .Z(n3325) );
  XOR U3775 ( .A(n3326), .B(n3327), .Z(n3323) );
  AND U3776 ( .A(n3328), .B(n3329), .Z(n3326) );
  XNOR U3777 ( .A(x[448]), .B(n3327), .Z(n3329) );
  XOR U3778 ( .A(n3330), .B(n3331), .Z(n3327) );
  AND U3779 ( .A(n3332), .B(n3333), .Z(n3330) );
  XNOR U3780 ( .A(x[447]), .B(n3331), .Z(n3333) );
  XOR U3781 ( .A(n3334), .B(n3335), .Z(n3331) );
  AND U3782 ( .A(n3336), .B(n3337), .Z(n3334) );
  XNOR U3783 ( .A(x[446]), .B(n3335), .Z(n3337) );
  XOR U3784 ( .A(n3338), .B(n3339), .Z(n3335) );
  AND U3785 ( .A(n3340), .B(n3341), .Z(n3338) );
  XNOR U3786 ( .A(x[445]), .B(n3339), .Z(n3341) );
  XOR U3787 ( .A(n3342), .B(n3343), .Z(n3339) );
  AND U3788 ( .A(n3344), .B(n3345), .Z(n3342) );
  XNOR U3789 ( .A(x[444]), .B(n3343), .Z(n3345) );
  XOR U3790 ( .A(n3346), .B(n3347), .Z(n3343) );
  AND U3791 ( .A(n3348), .B(n3349), .Z(n3346) );
  XNOR U3792 ( .A(x[443]), .B(n3347), .Z(n3349) );
  XOR U3793 ( .A(n3350), .B(n3351), .Z(n3347) );
  AND U3794 ( .A(n3352), .B(n3353), .Z(n3350) );
  XNOR U3795 ( .A(x[442]), .B(n3351), .Z(n3353) );
  XOR U3796 ( .A(n3354), .B(n3355), .Z(n3351) );
  AND U3797 ( .A(n3356), .B(n3357), .Z(n3354) );
  XNOR U3798 ( .A(x[441]), .B(n3355), .Z(n3357) );
  XOR U3799 ( .A(n3358), .B(n3359), .Z(n3355) );
  AND U3800 ( .A(n3360), .B(n3361), .Z(n3358) );
  XNOR U3801 ( .A(x[440]), .B(n3359), .Z(n3361) );
  XOR U3802 ( .A(n3362), .B(n3363), .Z(n3359) );
  AND U3803 ( .A(n3364), .B(n3365), .Z(n3362) );
  XNOR U3804 ( .A(x[439]), .B(n3363), .Z(n3365) );
  XOR U3805 ( .A(n3366), .B(n3367), .Z(n3363) );
  AND U3806 ( .A(n3368), .B(n3369), .Z(n3366) );
  XNOR U3807 ( .A(x[438]), .B(n3367), .Z(n3369) );
  XOR U3808 ( .A(n3370), .B(n3371), .Z(n3367) );
  AND U3809 ( .A(n3372), .B(n3373), .Z(n3370) );
  XNOR U3810 ( .A(x[437]), .B(n3371), .Z(n3373) );
  XOR U3811 ( .A(n3374), .B(n3375), .Z(n3371) );
  AND U3812 ( .A(n3376), .B(n3377), .Z(n3374) );
  XNOR U3813 ( .A(x[436]), .B(n3375), .Z(n3377) );
  XOR U3814 ( .A(n3378), .B(n3379), .Z(n3375) );
  AND U3815 ( .A(n3380), .B(n3381), .Z(n3378) );
  XNOR U3816 ( .A(x[435]), .B(n3379), .Z(n3381) );
  XOR U3817 ( .A(n3382), .B(n3383), .Z(n3379) );
  AND U3818 ( .A(n3384), .B(n3385), .Z(n3382) );
  XNOR U3819 ( .A(x[434]), .B(n3383), .Z(n3385) );
  XOR U3820 ( .A(n3386), .B(n3387), .Z(n3383) );
  AND U3821 ( .A(n3388), .B(n3389), .Z(n3386) );
  XNOR U3822 ( .A(x[433]), .B(n3387), .Z(n3389) );
  XOR U3823 ( .A(n3390), .B(n3391), .Z(n3387) );
  AND U3824 ( .A(n3392), .B(n3393), .Z(n3390) );
  XNOR U3825 ( .A(x[432]), .B(n3391), .Z(n3393) );
  XOR U3826 ( .A(n3394), .B(n3395), .Z(n3391) );
  AND U3827 ( .A(n3396), .B(n3397), .Z(n3394) );
  XNOR U3828 ( .A(x[431]), .B(n3395), .Z(n3397) );
  XOR U3829 ( .A(n3398), .B(n3399), .Z(n3395) );
  AND U3830 ( .A(n3400), .B(n3401), .Z(n3398) );
  XNOR U3831 ( .A(x[430]), .B(n3399), .Z(n3401) );
  XOR U3832 ( .A(n3402), .B(n3403), .Z(n3399) );
  AND U3833 ( .A(n3404), .B(n3405), .Z(n3402) );
  XNOR U3834 ( .A(x[429]), .B(n3403), .Z(n3405) );
  XOR U3835 ( .A(n3406), .B(n3407), .Z(n3403) );
  AND U3836 ( .A(n3408), .B(n3409), .Z(n3406) );
  XNOR U3837 ( .A(x[428]), .B(n3407), .Z(n3409) );
  XOR U3838 ( .A(n3410), .B(n3411), .Z(n3407) );
  AND U3839 ( .A(n3412), .B(n3413), .Z(n3410) );
  XNOR U3840 ( .A(x[427]), .B(n3411), .Z(n3413) );
  XOR U3841 ( .A(n3414), .B(n3415), .Z(n3411) );
  AND U3842 ( .A(n3416), .B(n3417), .Z(n3414) );
  XNOR U3843 ( .A(x[426]), .B(n3415), .Z(n3417) );
  XOR U3844 ( .A(n3418), .B(n3419), .Z(n3415) );
  AND U3845 ( .A(n3420), .B(n3421), .Z(n3418) );
  XNOR U3846 ( .A(x[425]), .B(n3419), .Z(n3421) );
  XOR U3847 ( .A(n3422), .B(n3423), .Z(n3419) );
  AND U3848 ( .A(n3424), .B(n3425), .Z(n3422) );
  XNOR U3849 ( .A(x[424]), .B(n3423), .Z(n3425) );
  XOR U3850 ( .A(n3426), .B(n3427), .Z(n3423) );
  AND U3851 ( .A(n3428), .B(n3429), .Z(n3426) );
  XNOR U3852 ( .A(x[423]), .B(n3427), .Z(n3429) );
  XOR U3853 ( .A(n3430), .B(n3431), .Z(n3427) );
  AND U3854 ( .A(n3432), .B(n3433), .Z(n3430) );
  XNOR U3855 ( .A(x[422]), .B(n3431), .Z(n3433) );
  XOR U3856 ( .A(n3434), .B(n3435), .Z(n3431) );
  AND U3857 ( .A(n3436), .B(n3437), .Z(n3434) );
  XNOR U3858 ( .A(x[421]), .B(n3435), .Z(n3437) );
  XOR U3859 ( .A(n3438), .B(n3439), .Z(n3435) );
  AND U3860 ( .A(n3440), .B(n3441), .Z(n3438) );
  XNOR U3861 ( .A(x[420]), .B(n3439), .Z(n3441) );
  XOR U3862 ( .A(n3442), .B(n3443), .Z(n3439) );
  AND U3863 ( .A(n3444), .B(n3445), .Z(n3442) );
  XNOR U3864 ( .A(x[419]), .B(n3443), .Z(n3445) );
  XOR U3865 ( .A(n3446), .B(n3447), .Z(n3443) );
  AND U3866 ( .A(n3448), .B(n3449), .Z(n3446) );
  XNOR U3867 ( .A(x[418]), .B(n3447), .Z(n3449) );
  XOR U3868 ( .A(n3450), .B(n3451), .Z(n3447) );
  AND U3869 ( .A(n3452), .B(n3453), .Z(n3450) );
  XNOR U3870 ( .A(x[417]), .B(n3451), .Z(n3453) );
  XOR U3871 ( .A(n3454), .B(n3455), .Z(n3451) );
  AND U3872 ( .A(n3456), .B(n3457), .Z(n3454) );
  XNOR U3873 ( .A(x[416]), .B(n3455), .Z(n3457) );
  XOR U3874 ( .A(n3458), .B(n3459), .Z(n3455) );
  AND U3875 ( .A(n3460), .B(n3461), .Z(n3458) );
  XNOR U3876 ( .A(x[415]), .B(n3459), .Z(n3461) );
  XOR U3877 ( .A(n3462), .B(n3463), .Z(n3459) );
  AND U3878 ( .A(n3464), .B(n3465), .Z(n3462) );
  XNOR U3879 ( .A(x[414]), .B(n3463), .Z(n3465) );
  XOR U3880 ( .A(n3466), .B(n3467), .Z(n3463) );
  AND U3881 ( .A(n3468), .B(n3469), .Z(n3466) );
  XNOR U3882 ( .A(x[413]), .B(n3467), .Z(n3469) );
  XOR U3883 ( .A(n3470), .B(n3471), .Z(n3467) );
  AND U3884 ( .A(n3472), .B(n3473), .Z(n3470) );
  XNOR U3885 ( .A(x[412]), .B(n3471), .Z(n3473) );
  XOR U3886 ( .A(n3474), .B(n3475), .Z(n3471) );
  AND U3887 ( .A(n3476), .B(n3477), .Z(n3474) );
  XNOR U3888 ( .A(x[411]), .B(n3475), .Z(n3477) );
  XOR U3889 ( .A(n3478), .B(n3479), .Z(n3475) );
  AND U3890 ( .A(n3480), .B(n3481), .Z(n3478) );
  XNOR U3891 ( .A(x[410]), .B(n3479), .Z(n3481) );
  XOR U3892 ( .A(n3482), .B(n3483), .Z(n3479) );
  AND U3893 ( .A(n3484), .B(n3485), .Z(n3482) );
  XNOR U3894 ( .A(x[409]), .B(n3483), .Z(n3485) );
  XOR U3895 ( .A(n3486), .B(n3487), .Z(n3483) );
  AND U3896 ( .A(n3488), .B(n3489), .Z(n3486) );
  XNOR U3897 ( .A(x[408]), .B(n3487), .Z(n3489) );
  XOR U3898 ( .A(n3490), .B(n3491), .Z(n3487) );
  AND U3899 ( .A(n3492), .B(n3493), .Z(n3490) );
  XNOR U3900 ( .A(x[407]), .B(n3491), .Z(n3493) );
  XOR U3901 ( .A(n3494), .B(n3495), .Z(n3491) );
  AND U3902 ( .A(n3496), .B(n3497), .Z(n3494) );
  XNOR U3903 ( .A(x[406]), .B(n3495), .Z(n3497) );
  XOR U3904 ( .A(n3498), .B(n3499), .Z(n3495) );
  AND U3905 ( .A(n3500), .B(n3501), .Z(n3498) );
  XNOR U3906 ( .A(x[405]), .B(n3499), .Z(n3501) );
  XOR U3907 ( .A(n3502), .B(n3503), .Z(n3499) );
  AND U3908 ( .A(n3504), .B(n3505), .Z(n3502) );
  XNOR U3909 ( .A(x[404]), .B(n3503), .Z(n3505) );
  XOR U3910 ( .A(n3506), .B(n3507), .Z(n3503) );
  AND U3911 ( .A(n3508), .B(n3509), .Z(n3506) );
  XNOR U3912 ( .A(x[403]), .B(n3507), .Z(n3509) );
  XOR U3913 ( .A(n3510), .B(n3511), .Z(n3507) );
  AND U3914 ( .A(n3512), .B(n3513), .Z(n3510) );
  XNOR U3915 ( .A(x[402]), .B(n3511), .Z(n3513) );
  XOR U3916 ( .A(n3514), .B(n3515), .Z(n3511) );
  AND U3917 ( .A(n3516), .B(n3517), .Z(n3514) );
  XNOR U3918 ( .A(x[401]), .B(n3515), .Z(n3517) );
  XOR U3919 ( .A(n3518), .B(n3519), .Z(n3515) );
  AND U3920 ( .A(n3520), .B(n3521), .Z(n3518) );
  XNOR U3921 ( .A(x[400]), .B(n3519), .Z(n3521) );
  XOR U3922 ( .A(n3522), .B(n3523), .Z(n3519) );
  AND U3923 ( .A(n3524), .B(n3525), .Z(n3522) );
  XNOR U3924 ( .A(x[399]), .B(n3523), .Z(n3525) );
  XOR U3925 ( .A(n3526), .B(n3527), .Z(n3523) );
  AND U3926 ( .A(n3528), .B(n3529), .Z(n3526) );
  XNOR U3927 ( .A(x[398]), .B(n3527), .Z(n3529) );
  XOR U3928 ( .A(n3530), .B(n3531), .Z(n3527) );
  AND U3929 ( .A(n3532), .B(n3533), .Z(n3530) );
  XNOR U3930 ( .A(x[397]), .B(n3531), .Z(n3533) );
  XOR U3931 ( .A(n3534), .B(n3535), .Z(n3531) );
  AND U3932 ( .A(n3536), .B(n3537), .Z(n3534) );
  XNOR U3933 ( .A(x[396]), .B(n3535), .Z(n3537) );
  XOR U3934 ( .A(n3538), .B(n3539), .Z(n3535) );
  AND U3935 ( .A(n3540), .B(n3541), .Z(n3538) );
  XNOR U3936 ( .A(x[395]), .B(n3539), .Z(n3541) );
  XOR U3937 ( .A(n3542), .B(n3543), .Z(n3539) );
  AND U3938 ( .A(n3544), .B(n3545), .Z(n3542) );
  XNOR U3939 ( .A(x[394]), .B(n3543), .Z(n3545) );
  XOR U3940 ( .A(n3546), .B(n3547), .Z(n3543) );
  AND U3941 ( .A(n3548), .B(n3549), .Z(n3546) );
  XNOR U3942 ( .A(x[393]), .B(n3547), .Z(n3549) );
  XOR U3943 ( .A(n3550), .B(n3551), .Z(n3547) );
  AND U3944 ( .A(n3552), .B(n3553), .Z(n3550) );
  XNOR U3945 ( .A(x[392]), .B(n3551), .Z(n3553) );
  XOR U3946 ( .A(n3554), .B(n3555), .Z(n3551) );
  AND U3947 ( .A(n3556), .B(n3557), .Z(n3554) );
  XNOR U3948 ( .A(x[391]), .B(n3555), .Z(n3557) );
  XOR U3949 ( .A(n3558), .B(n3559), .Z(n3555) );
  AND U3950 ( .A(n3560), .B(n3561), .Z(n3558) );
  XNOR U3951 ( .A(x[390]), .B(n3559), .Z(n3561) );
  XOR U3952 ( .A(n3562), .B(n3563), .Z(n3559) );
  AND U3953 ( .A(n3564), .B(n3565), .Z(n3562) );
  XNOR U3954 ( .A(x[389]), .B(n3563), .Z(n3565) );
  XOR U3955 ( .A(n3566), .B(n3567), .Z(n3563) );
  AND U3956 ( .A(n3568), .B(n3569), .Z(n3566) );
  XNOR U3957 ( .A(x[388]), .B(n3567), .Z(n3569) );
  XOR U3958 ( .A(n3570), .B(n3571), .Z(n3567) );
  AND U3959 ( .A(n3572), .B(n3573), .Z(n3570) );
  XNOR U3960 ( .A(x[387]), .B(n3571), .Z(n3573) );
  XOR U3961 ( .A(n3574), .B(n3575), .Z(n3571) );
  AND U3962 ( .A(n3576), .B(n3577), .Z(n3574) );
  XNOR U3963 ( .A(x[386]), .B(n3575), .Z(n3577) );
  XOR U3964 ( .A(n3578), .B(n3579), .Z(n3575) );
  AND U3965 ( .A(n3580), .B(n3581), .Z(n3578) );
  XNOR U3966 ( .A(x[385]), .B(n3579), .Z(n3581) );
  XOR U3967 ( .A(n3582), .B(n3583), .Z(n3579) );
  AND U3968 ( .A(n3584), .B(n3585), .Z(n3582) );
  XNOR U3969 ( .A(x[384]), .B(n3583), .Z(n3585) );
  XOR U3970 ( .A(n3586), .B(n3587), .Z(n3583) );
  AND U3971 ( .A(n3588), .B(n3589), .Z(n3586) );
  XNOR U3972 ( .A(x[383]), .B(n3587), .Z(n3589) );
  XOR U3973 ( .A(n3590), .B(n3591), .Z(n3587) );
  AND U3974 ( .A(n3592), .B(n3593), .Z(n3590) );
  XNOR U3975 ( .A(x[382]), .B(n3591), .Z(n3593) );
  XOR U3976 ( .A(n3594), .B(n3595), .Z(n3591) );
  AND U3977 ( .A(n3596), .B(n3597), .Z(n3594) );
  XNOR U3978 ( .A(x[381]), .B(n3595), .Z(n3597) );
  XOR U3979 ( .A(n3598), .B(n3599), .Z(n3595) );
  AND U3980 ( .A(n3600), .B(n3601), .Z(n3598) );
  XNOR U3981 ( .A(x[380]), .B(n3599), .Z(n3601) );
  XOR U3982 ( .A(n3602), .B(n3603), .Z(n3599) );
  AND U3983 ( .A(n3604), .B(n3605), .Z(n3602) );
  XNOR U3984 ( .A(x[379]), .B(n3603), .Z(n3605) );
  XOR U3985 ( .A(n3606), .B(n3607), .Z(n3603) );
  AND U3986 ( .A(n3608), .B(n3609), .Z(n3606) );
  XNOR U3987 ( .A(x[378]), .B(n3607), .Z(n3609) );
  XOR U3988 ( .A(n3610), .B(n3611), .Z(n3607) );
  AND U3989 ( .A(n3612), .B(n3613), .Z(n3610) );
  XNOR U3990 ( .A(x[377]), .B(n3611), .Z(n3613) );
  XOR U3991 ( .A(n3614), .B(n3615), .Z(n3611) );
  AND U3992 ( .A(n3616), .B(n3617), .Z(n3614) );
  XNOR U3993 ( .A(x[376]), .B(n3615), .Z(n3617) );
  XOR U3994 ( .A(n3618), .B(n3619), .Z(n3615) );
  AND U3995 ( .A(n3620), .B(n3621), .Z(n3618) );
  XNOR U3996 ( .A(x[375]), .B(n3619), .Z(n3621) );
  XOR U3997 ( .A(n3622), .B(n3623), .Z(n3619) );
  AND U3998 ( .A(n3624), .B(n3625), .Z(n3622) );
  XNOR U3999 ( .A(x[374]), .B(n3623), .Z(n3625) );
  XOR U4000 ( .A(n3626), .B(n3627), .Z(n3623) );
  AND U4001 ( .A(n3628), .B(n3629), .Z(n3626) );
  XNOR U4002 ( .A(x[373]), .B(n3627), .Z(n3629) );
  XOR U4003 ( .A(n3630), .B(n3631), .Z(n3627) );
  AND U4004 ( .A(n3632), .B(n3633), .Z(n3630) );
  XNOR U4005 ( .A(x[372]), .B(n3631), .Z(n3633) );
  XOR U4006 ( .A(n3634), .B(n3635), .Z(n3631) );
  AND U4007 ( .A(n3636), .B(n3637), .Z(n3634) );
  XNOR U4008 ( .A(x[371]), .B(n3635), .Z(n3637) );
  XOR U4009 ( .A(n3638), .B(n3639), .Z(n3635) );
  AND U4010 ( .A(n3640), .B(n3641), .Z(n3638) );
  XNOR U4011 ( .A(x[370]), .B(n3639), .Z(n3641) );
  XOR U4012 ( .A(n3642), .B(n3643), .Z(n3639) );
  AND U4013 ( .A(n3644), .B(n3645), .Z(n3642) );
  XNOR U4014 ( .A(x[369]), .B(n3643), .Z(n3645) );
  XOR U4015 ( .A(n3646), .B(n3647), .Z(n3643) );
  AND U4016 ( .A(n3648), .B(n3649), .Z(n3646) );
  XNOR U4017 ( .A(x[368]), .B(n3647), .Z(n3649) );
  XOR U4018 ( .A(n3650), .B(n3651), .Z(n3647) );
  AND U4019 ( .A(n3652), .B(n3653), .Z(n3650) );
  XNOR U4020 ( .A(x[367]), .B(n3651), .Z(n3653) );
  XOR U4021 ( .A(n3654), .B(n3655), .Z(n3651) );
  AND U4022 ( .A(n3656), .B(n3657), .Z(n3654) );
  XNOR U4023 ( .A(x[366]), .B(n3655), .Z(n3657) );
  XOR U4024 ( .A(n3658), .B(n3659), .Z(n3655) );
  AND U4025 ( .A(n3660), .B(n3661), .Z(n3658) );
  XNOR U4026 ( .A(x[365]), .B(n3659), .Z(n3661) );
  XOR U4027 ( .A(n3662), .B(n3663), .Z(n3659) );
  AND U4028 ( .A(n3664), .B(n3665), .Z(n3662) );
  XNOR U4029 ( .A(x[364]), .B(n3663), .Z(n3665) );
  XOR U4030 ( .A(n3666), .B(n3667), .Z(n3663) );
  AND U4031 ( .A(n3668), .B(n3669), .Z(n3666) );
  XNOR U4032 ( .A(x[363]), .B(n3667), .Z(n3669) );
  XOR U4033 ( .A(n3670), .B(n3671), .Z(n3667) );
  AND U4034 ( .A(n3672), .B(n3673), .Z(n3670) );
  XNOR U4035 ( .A(x[362]), .B(n3671), .Z(n3673) );
  XOR U4036 ( .A(n3674), .B(n3675), .Z(n3671) );
  AND U4037 ( .A(n3676), .B(n3677), .Z(n3674) );
  XNOR U4038 ( .A(x[361]), .B(n3675), .Z(n3677) );
  XOR U4039 ( .A(n3678), .B(n3679), .Z(n3675) );
  AND U4040 ( .A(n3680), .B(n3681), .Z(n3678) );
  XNOR U4041 ( .A(x[360]), .B(n3679), .Z(n3681) );
  XOR U4042 ( .A(n3682), .B(n3683), .Z(n3679) );
  AND U4043 ( .A(n3684), .B(n3685), .Z(n3682) );
  XNOR U4044 ( .A(x[359]), .B(n3683), .Z(n3685) );
  XOR U4045 ( .A(n3686), .B(n3687), .Z(n3683) );
  AND U4046 ( .A(n3688), .B(n3689), .Z(n3686) );
  XNOR U4047 ( .A(x[358]), .B(n3687), .Z(n3689) );
  XOR U4048 ( .A(n3690), .B(n3691), .Z(n3687) );
  AND U4049 ( .A(n3692), .B(n3693), .Z(n3690) );
  XNOR U4050 ( .A(x[357]), .B(n3691), .Z(n3693) );
  XOR U4051 ( .A(n3694), .B(n3695), .Z(n3691) );
  AND U4052 ( .A(n3696), .B(n3697), .Z(n3694) );
  XNOR U4053 ( .A(x[356]), .B(n3695), .Z(n3697) );
  XOR U4054 ( .A(n3698), .B(n3699), .Z(n3695) );
  AND U4055 ( .A(n3700), .B(n3701), .Z(n3698) );
  XNOR U4056 ( .A(x[355]), .B(n3699), .Z(n3701) );
  XOR U4057 ( .A(n3702), .B(n3703), .Z(n3699) );
  AND U4058 ( .A(n3704), .B(n3705), .Z(n3702) );
  XNOR U4059 ( .A(x[354]), .B(n3703), .Z(n3705) );
  XOR U4060 ( .A(n3706), .B(n3707), .Z(n3703) );
  AND U4061 ( .A(n3708), .B(n3709), .Z(n3706) );
  XNOR U4062 ( .A(x[353]), .B(n3707), .Z(n3709) );
  XOR U4063 ( .A(n3710), .B(n3711), .Z(n3707) );
  AND U4064 ( .A(n3712), .B(n3713), .Z(n3710) );
  XNOR U4065 ( .A(x[352]), .B(n3711), .Z(n3713) );
  XOR U4066 ( .A(n3714), .B(n3715), .Z(n3711) );
  AND U4067 ( .A(n3716), .B(n3717), .Z(n3714) );
  XNOR U4068 ( .A(x[351]), .B(n3715), .Z(n3717) );
  XOR U4069 ( .A(n3718), .B(n3719), .Z(n3715) );
  AND U4070 ( .A(n3720), .B(n3721), .Z(n3718) );
  XNOR U4071 ( .A(x[350]), .B(n3719), .Z(n3721) );
  XOR U4072 ( .A(n3722), .B(n3723), .Z(n3719) );
  AND U4073 ( .A(n3724), .B(n3725), .Z(n3722) );
  XNOR U4074 ( .A(x[349]), .B(n3723), .Z(n3725) );
  XOR U4075 ( .A(n3726), .B(n3727), .Z(n3723) );
  AND U4076 ( .A(n3728), .B(n3729), .Z(n3726) );
  XNOR U4077 ( .A(x[348]), .B(n3727), .Z(n3729) );
  XOR U4078 ( .A(n3730), .B(n3731), .Z(n3727) );
  AND U4079 ( .A(n3732), .B(n3733), .Z(n3730) );
  XNOR U4080 ( .A(x[347]), .B(n3731), .Z(n3733) );
  XOR U4081 ( .A(n3734), .B(n3735), .Z(n3731) );
  AND U4082 ( .A(n3736), .B(n3737), .Z(n3734) );
  XNOR U4083 ( .A(x[346]), .B(n3735), .Z(n3737) );
  XOR U4084 ( .A(n3738), .B(n3739), .Z(n3735) );
  AND U4085 ( .A(n3740), .B(n3741), .Z(n3738) );
  XNOR U4086 ( .A(x[345]), .B(n3739), .Z(n3741) );
  XOR U4087 ( .A(n3742), .B(n3743), .Z(n3739) );
  AND U4088 ( .A(n3744), .B(n3745), .Z(n3742) );
  XNOR U4089 ( .A(x[344]), .B(n3743), .Z(n3745) );
  XOR U4090 ( .A(n3746), .B(n3747), .Z(n3743) );
  AND U4091 ( .A(n3748), .B(n3749), .Z(n3746) );
  XNOR U4092 ( .A(x[343]), .B(n3747), .Z(n3749) );
  XOR U4093 ( .A(n3750), .B(n3751), .Z(n3747) );
  AND U4094 ( .A(n3752), .B(n3753), .Z(n3750) );
  XNOR U4095 ( .A(x[342]), .B(n3751), .Z(n3753) );
  XOR U4096 ( .A(n3754), .B(n3755), .Z(n3751) );
  AND U4097 ( .A(n3756), .B(n3757), .Z(n3754) );
  XNOR U4098 ( .A(x[341]), .B(n3755), .Z(n3757) );
  XOR U4099 ( .A(n3758), .B(n3759), .Z(n3755) );
  AND U4100 ( .A(n3760), .B(n3761), .Z(n3758) );
  XNOR U4101 ( .A(x[340]), .B(n3759), .Z(n3761) );
  XOR U4102 ( .A(n3762), .B(n3763), .Z(n3759) );
  AND U4103 ( .A(n3764), .B(n3765), .Z(n3762) );
  XNOR U4104 ( .A(x[339]), .B(n3763), .Z(n3765) );
  XOR U4105 ( .A(n3766), .B(n3767), .Z(n3763) );
  AND U4106 ( .A(n3768), .B(n3769), .Z(n3766) );
  XNOR U4107 ( .A(x[338]), .B(n3767), .Z(n3769) );
  XOR U4108 ( .A(n3770), .B(n3771), .Z(n3767) );
  AND U4109 ( .A(n3772), .B(n3773), .Z(n3770) );
  XNOR U4110 ( .A(x[337]), .B(n3771), .Z(n3773) );
  XOR U4111 ( .A(n3774), .B(n3775), .Z(n3771) );
  AND U4112 ( .A(n3776), .B(n3777), .Z(n3774) );
  XNOR U4113 ( .A(x[336]), .B(n3775), .Z(n3777) );
  XOR U4114 ( .A(n3778), .B(n3779), .Z(n3775) );
  AND U4115 ( .A(n3780), .B(n3781), .Z(n3778) );
  XNOR U4116 ( .A(x[335]), .B(n3779), .Z(n3781) );
  XOR U4117 ( .A(n3782), .B(n3783), .Z(n3779) );
  AND U4118 ( .A(n3784), .B(n3785), .Z(n3782) );
  XNOR U4119 ( .A(x[334]), .B(n3783), .Z(n3785) );
  XOR U4120 ( .A(n3786), .B(n3787), .Z(n3783) );
  AND U4121 ( .A(n3788), .B(n3789), .Z(n3786) );
  XNOR U4122 ( .A(x[333]), .B(n3787), .Z(n3789) );
  XOR U4123 ( .A(n3790), .B(n3791), .Z(n3787) );
  AND U4124 ( .A(n3792), .B(n3793), .Z(n3790) );
  XNOR U4125 ( .A(x[332]), .B(n3791), .Z(n3793) );
  XOR U4126 ( .A(n3794), .B(n3795), .Z(n3791) );
  AND U4127 ( .A(n3796), .B(n3797), .Z(n3794) );
  XNOR U4128 ( .A(x[331]), .B(n3795), .Z(n3797) );
  XOR U4129 ( .A(n3798), .B(n3799), .Z(n3795) );
  AND U4130 ( .A(n3800), .B(n3801), .Z(n3798) );
  XNOR U4131 ( .A(x[330]), .B(n3799), .Z(n3801) );
  XOR U4132 ( .A(n3802), .B(n3803), .Z(n3799) );
  AND U4133 ( .A(n3804), .B(n3805), .Z(n3802) );
  XNOR U4134 ( .A(x[329]), .B(n3803), .Z(n3805) );
  XOR U4135 ( .A(n3806), .B(n3807), .Z(n3803) );
  AND U4136 ( .A(n3808), .B(n3809), .Z(n3806) );
  XNOR U4137 ( .A(x[328]), .B(n3807), .Z(n3809) );
  XOR U4138 ( .A(n3810), .B(n3811), .Z(n3807) );
  AND U4139 ( .A(n3812), .B(n3813), .Z(n3810) );
  XNOR U4140 ( .A(x[327]), .B(n3811), .Z(n3813) );
  XOR U4141 ( .A(n3814), .B(n3815), .Z(n3811) );
  AND U4142 ( .A(n3816), .B(n3817), .Z(n3814) );
  XNOR U4143 ( .A(x[326]), .B(n3815), .Z(n3817) );
  XOR U4144 ( .A(n3818), .B(n3819), .Z(n3815) );
  AND U4145 ( .A(n3820), .B(n3821), .Z(n3818) );
  XNOR U4146 ( .A(x[325]), .B(n3819), .Z(n3821) );
  XOR U4147 ( .A(n3822), .B(n3823), .Z(n3819) );
  AND U4148 ( .A(n3824), .B(n3825), .Z(n3822) );
  XNOR U4149 ( .A(x[324]), .B(n3823), .Z(n3825) );
  XOR U4150 ( .A(n3826), .B(n3827), .Z(n3823) );
  AND U4151 ( .A(n3828), .B(n3829), .Z(n3826) );
  XNOR U4152 ( .A(x[323]), .B(n3827), .Z(n3829) );
  XOR U4153 ( .A(n3830), .B(n3831), .Z(n3827) );
  AND U4154 ( .A(n3832), .B(n3833), .Z(n3830) );
  XNOR U4155 ( .A(x[322]), .B(n3831), .Z(n3833) );
  XOR U4156 ( .A(n3834), .B(n3835), .Z(n3831) );
  AND U4157 ( .A(n3836), .B(n3837), .Z(n3834) );
  XNOR U4158 ( .A(x[321]), .B(n3835), .Z(n3837) );
  XOR U4159 ( .A(n3838), .B(n3839), .Z(n3835) );
  AND U4160 ( .A(n3840), .B(n3841), .Z(n3838) );
  XNOR U4161 ( .A(x[320]), .B(n3839), .Z(n3841) );
  XOR U4162 ( .A(n3842), .B(n3843), .Z(n3839) );
  AND U4163 ( .A(n3844), .B(n3845), .Z(n3842) );
  XNOR U4164 ( .A(x[319]), .B(n3843), .Z(n3845) );
  XOR U4165 ( .A(n3846), .B(n3847), .Z(n3843) );
  AND U4166 ( .A(n3848), .B(n3849), .Z(n3846) );
  XNOR U4167 ( .A(x[318]), .B(n3847), .Z(n3849) );
  XOR U4168 ( .A(n3850), .B(n3851), .Z(n3847) );
  AND U4169 ( .A(n3852), .B(n3853), .Z(n3850) );
  XNOR U4170 ( .A(x[317]), .B(n3851), .Z(n3853) );
  XOR U4171 ( .A(n3854), .B(n3855), .Z(n3851) );
  AND U4172 ( .A(n3856), .B(n3857), .Z(n3854) );
  XNOR U4173 ( .A(x[316]), .B(n3855), .Z(n3857) );
  XOR U4174 ( .A(n3858), .B(n3859), .Z(n3855) );
  AND U4175 ( .A(n3860), .B(n3861), .Z(n3858) );
  XNOR U4176 ( .A(x[315]), .B(n3859), .Z(n3861) );
  XOR U4177 ( .A(n3862), .B(n3863), .Z(n3859) );
  AND U4178 ( .A(n3864), .B(n3865), .Z(n3862) );
  XNOR U4179 ( .A(x[314]), .B(n3863), .Z(n3865) );
  XOR U4180 ( .A(n3866), .B(n3867), .Z(n3863) );
  AND U4181 ( .A(n3868), .B(n3869), .Z(n3866) );
  XNOR U4182 ( .A(x[313]), .B(n3867), .Z(n3869) );
  XOR U4183 ( .A(n3870), .B(n3871), .Z(n3867) );
  AND U4184 ( .A(n3872), .B(n3873), .Z(n3870) );
  XNOR U4185 ( .A(x[312]), .B(n3871), .Z(n3873) );
  XOR U4186 ( .A(n3874), .B(n3875), .Z(n3871) );
  AND U4187 ( .A(n3876), .B(n3877), .Z(n3874) );
  XNOR U4188 ( .A(x[311]), .B(n3875), .Z(n3877) );
  XOR U4189 ( .A(n3878), .B(n3879), .Z(n3875) );
  AND U4190 ( .A(n3880), .B(n3881), .Z(n3878) );
  XNOR U4191 ( .A(x[310]), .B(n3879), .Z(n3881) );
  XOR U4192 ( .A(n3882), .B(n3883), .Z(n3879) );
  AND U4193 ( .A(n3884), .B(n3885), .Z(n3882) );
  XNOR U4194 ( .A(x[309]), .B(n3883), .Z(n3885) );
  XOR U4195 ( .A(n3886), .B(n3887), .Z(n3883) );
  AND U4196 ( .A(n3888), .B(n3889), .Z(n3886) );
  XNOR U4197 ( .A(x[308]), .B(n3887), .Z(n3889) );
  XOR U4198 ( .A(n3890), .B(n3891), .Z(n3887) );
  AND U4199 ( .A(n3892), .B(n3893), .Z(n3890) );
  XNOR U4200 ( .A(x[307]), .B(n3891), .Z(n3893) );
  XOR U4201 ( .A(n3894), .B(n3895), .Z(n3891) );
  AND U4202 ( .A(n3896), .B(n3897), .Z(n3894) );
  XNOR U4203 ( .A(x[306]), .B(n3895), .Z(n3897) );
  XOR U4204 ( .A(n3898), .B(n3899), .Z(n3895) );
  AND U4205 ( .A(n3900), .B(n3901), .Z(n3898) );
  XNOR U4206 ( .A(x[305]), .B(n3899), .Z(n3901) );
  XOR U4207 ( .A(n3902), .B(n3903), .Z(n3899) );
  AND U4208 ( .A(n3904), .B(n3905), .Z(n3902) );
  XNOR U4209 ( .A(x[304]), .B(n3903), .Z(n3905) );
  XOR U4210 ( .A(n3906), .B(n3907), .Z(n3903) );
  AND U4211 ( .A(n3908), .B(n3909), .Z(n3906) );
  XNOR U4212 ( .A(x[303]), .B(n3907), .Z(n3909) );
  XOR U4213 ( .A(n3910), .B(n3911), .Z(n3907) );
  AND U4214 ( .A(n3912), .B(n3913), .Z(n3910) );
  XNOR U4215 ( .A(x[302]), .B(n3911), .Z(n3913) );
  XOR U4216 ( .A(n3914), .B(n3915), .Z(n3911) );
  AND U4217 ( .A(n3916), .B(n3917), .Z(n3914) );
  XNOR U4218 ( .A(x[301]), .B(n3915), .Z(n3917) );
  XOR U4219 ( .A(n3918), .B(n3919), .Z(n3915) );
  AND U4220 ( .A(n3920), .B(n3921), .Z(n3918) );
  XNOR U4221 ( .A(x[300]), .B(n3919), .Z(n3921) );
  XOR U4222 ( .A(n3922), .B(n3923), .Z(n3919) );
  AND U4223 ( .A(n3924), .B(n3925), .Z(n3922) );
  XNOR U4224 ( .A(x[299]), .B(n3923), .Z(n3925) );
  XOR U4225 ( .A(n3926), .B(n3927), .Z(n3923) );
  AND U4226 ( .A(n3928), .B(n3929), .Z(n3926) );
  XNOR U4227 ( .A(x[298]), .B(n3927), .Z(n3929) );
  XOR U4228 ( .A(n3930), .B(n3931), .Z(n3927) );
  AND U4229 ( .A(n3932), .B(n3933), .Z(n3930) );
  XNOR U4230 ( .A(x[297]), .B(n3931), .Z(n3933) );
  XOR U4231 ( .A(n3934), .B(n3935), .Z(n3931) );
  AND U4232 ( .A(n3936), .B(n3937), .Z(n3934) );
  XNOR U4233 ( .A(x[296]), .B(n3935), .Z(n3937) );
  XOR U4234 ( .A(n3938), .B(n3939), .Z(n3935) );
  AND U4235 ( .A(n3940), .B(n3941), .Z(n3938) );
  XNOR U4236 ( .A(x[295]), .B(n3939), .Z(n3941) );
  XOR U4237 ( .A(n3942), .B(n3943), .Z(n3939) );
  AND U4238 ( .A(n3944), .B(n3945), .Z(n3942) );
  XNOR U4239 ( .A(x[294]), .B(n3943), .Z(n3945) );
  XOR U4240 ( .A(n3946), .B(n3947), .Z(n3943) );
  AND U4241 ( .A(n3948), .B(n3949), .Z(n3946) );
  XNOR U4242 ( .A(x[293]), .B(n3947), .Z(n3949) );
  XOR U4243 ( .A(n3950), .B(n3951), .Z(n3947) );
  AND U4244 ( .A(n3952), .B(n3953), .Z(n3950) );
  XNOR U4245 ( .A(x[292]), .B(n3951), .Z(n3953) );
  XOR U4246 ( .A(n3954), .B(n3955), .Z(n3951) );
  AND U4247 ( .A(n3956), .B(n3957), .Z(n3954) );
  XNOR U4248 ( .A(x[291]), .B(n3955), .Z(n3957) );
  XOR U4249 ( .A(n3958), .B(n3959), .Z(n3955) );
  AND U4250 ( .A(n3960), .B(n3961), .Z(n3958) );
  XNOR U4251 ( .A(x[290]), .B(n3959), .Z(n3961) );
  XOR U4252 ( .A(n3962), .B(n3963), .Z(n3959) );
  AND U4253 ( .A(n3964), .B(n3965), .Z(n3962) );
  XNOR U4254 ( .A(x[289]), .B(n3963), .Z(n3965) );
  XOR U4255 ( .A(n3966), .B(n3967), .Z(n3963) );
  AND U4256 ( .A(n3968), .B(n3969), .Z(n3966) );
  XNOR U4257 ( .A(x[288]), .B(n3967), .Z(n3969) );
  XOR U4258 ( .A(n3970), .B(n3971), .Z(n3967) );
  AND U4259 ( .A(n3972), .B(n3973), .Z(n3970) );
  XNOR U4260 ( .A(x[287]), .B(n3971), .Z(n3973) );
  XOR U4261 ( .A(n3974), .B(n3975), .Z(n3971) );
  AND U4262 ( .A(n3976), .B(n3977), .Z(n3974) );
  XNOR U4263 ( .A(x[286]), .B(n3975), .Z(n3977) );
  XOR U4264 ( .A(n3978), .B(n3979), .Z(n3975) );
  AND U4265 ( .A(n3980), .B(n3981), .Z(n3978) );
  XNOR U4266 ( .A(x[285]), .B(n3979), .Z(n3981) );
  XOR U4267 ( .A(n3982), .B(n3983), .Z(n3979) );
  AND U4268 ( .A(n3984), .B(n3985), .Z(n3982) );
  XNOR U4269 ( .A(x[284]), .B(n3983), .Z(n3985) );
  XOR U4270 ( .A(n3986), .B(n3987), .Z(n3983) );
  AND U4271 ( .A(n3988), .B(n3989), .Z(n3986) );
  XNOR U4272 ( .A(x[283]), .B(n3987), .Z(n3989) );
  XOR U4273 ( .A(n3990), .B(n3991), .Z(n3987) );
  AND U4274 ( .A(n3992), .B(n3993), .Z(n3990) );
  XNOR U4275 ( .A(x[282]), .B(n3991), .Z(n3993) );
  XOR U4276 ( .A(n3994), .B(n3995), .Z(n3991) );
  AND U4277 ( .A(n3996), .B(n3997), .Z(n3994) );
  XNOR U4278 ( .A(x[281]), .B(n3995), .Z(n3997) );
  XOR U4279 ( .A(n3998), .B(n3999), .Z(n3995) );
  AND U4280 ( .A(n4000), .B(n4001), .Z(n3998) );
  XNOR U4281 ( .A(x[280]), .B(n3999), .Z(n4001) );
  XOR U4282 ( .A(n4002), .B(n4003), .Z(n3999) );
  AND U4283 ( .A(n4004), .B(n4005), .Z(n4002) );
  XNOR U4284 ( .A(x[279]), .B(n4003), .Z(n4005) );
  XOR U4285 ( .A(n4006), .B(n4007), .Z(n4003) );
  AND U4286 ( .A(n4008), .B(n4009), .Z(n4006) );
  XNOR U4287 ( .A(x[278]), .B(n4007), .Z(n4009) );
  XOR U4288 ( .A(n4010), .B(n4011), .Z(n4007) );
  AND U4289 ( .A(n4012), .B(n4013), .Z(n4010) );
  XNOR U4290 ( .A(x[277]), .B(n4011), .Z(n4013) );
  XOR U4291 ( .A(n4014), .B(n4015), .Z(n4011) );
  AND U4292 ( .A(n4016), .B(n4017), .Z(n4014) );
  XNOR U4293 ( .A(x[276]), .B(n4015), .Z(n4017) );
  XOR U4294 ( .A(n4018), .B(n4019), .Z(n4015) );
  AND U4295 ( .A(n4020), .B(n4021), .Z(n4018) );
  XNOR U4296 ( .A(x[275]), .B(n4019), .Z(n4021) );
  XOR U4297 ( .A(n4022), .B(n4023), .Z(n4019) );
  AND U4298 ( .A(n4024), .B(n4025), .Z(n4022) );
  XNOR U4299 ( .A(x[274]), .B(n4023), .Z(n4025) );
  XOR U4300 ( .A(n4026), .B(n4027), .Z(n4023) );
  AND U4301 ( .A(n4028), .B(n4029), .Z(n4026) );
  XNOR U4302 ( .A(x[273]), .B(n4027), .Z(n4029) );
  XOR U4303 ( .A(n4030), .B(n4031), .Z(n4027) );
  AND U4304 ( .A(n4032), .B(n4033), .Z(n4030) );
  XNOR U4305 ( .A(x[272]), .B(n4031), .Z(n4033) );
  XOR U4306 ( .A(n4034), .B(n4035), .Z(n4031) );
  AND U4307 ( .A(n4036), .B(n4037), .Z(n4034) );
  XNOR U4308 ( .A(x[271]), .B(n4035), .Z(n4037) );
  XOR U4309 ( .A(n4038), .B(n4039), .Z(n4035) );
  AND U4310 ( .A(n4040), .B(n4041), .Z(n4038) );
  XNOR U4311 ( .A(x[270]), .B(n4039), .Z(n4041) );
  XOR U4312 ( .A(n4042), .B(n4043), .Z(n4039) );
  AND U4313 ( .A(n4044), .B(n4045), .Z(n4042) );
  XNOR U4314 ( .A(x[269]), .B(n4043), .Z(n4045) );
  XOR U4315 ( .A(n4046), .B(n4047), .Z(n4043) );
  AND U4316 ( .A(n4048), .B(n4049), .Z(n4046) );
  XNOR U4317 ( .A(x[268]), .B(n4047), .Z(n4049) );
  XOR U4318 ( .A(n4050), .B(n4051), .Z(n4047) );
  AND U4319 ( .A(n4052), .B(n4053), .Z(n4050) );
  XNOR U4320 ( .A(x[267]), .B(n4051), .Z(n4053) );
  XOR U4321 ( .A(n4054), .B(n4055), .Z(n4051) );
  AND U4322 ( .A(n4056), .B(n4057), .Z(n4054) );
  XNOR U4323 ( .A(x[266]), .B(n4055), .Z(n4057) );
  XOR U4324 ( .A(n4058), .B(n4059), .Z(n4055) );
  AND U4325 ( .A(n4060), .B(n4061), .Z(n4058) );
  XNOR U4326 ( .A(x[265]), .B(n4059), .Z(n4061) );
  XOR U4327 ( .A(n4062), .B(n4063), .Z(n4059) );
  AND U4328 ( .A(n4064), .B(n4065), .Z(n4062) );
  XNOR U4329 ( .A(x[264]), .B(n4063), .Z(n4065) );
  XOR U4330 ( .A(n4066), .B(n4067), .Z(n4063) );
  AND U4331 ( .A(n4068), .B(n4069), .Z(n4066) );
  XNOR U4332 ( .A(x[263]), .B(n4067), .Z(n4069) );
  XOR U4333 ( .A(n4070), .B(n4071), .Z(n4067) );
  AND U4334 ( .A(n4072), .B(n4073), .Z(n4070) );
  XNOR U4335 ( .A(x[262]), .B(n4071), .Z(n4073) );
  XOR U4336 ( .A(n4074), .B(n4075), .Z(n4071) );
  AND U4337 ( .A(n4076), .B(n4077), .Z(n4074) );
  XNOR U4338 ( .A(x[261]), .B(n4075), .Z(n4077) );
  XOR U4339 ( .A(n4078), .B(n4079), .Z(n4075) );
  AND U4340 ( .A(n4080), .B(n4081), .Z(n4078) );
  XNOR U4341 ( .A(x[260]), .B(n4079), .Z(n4081) );
  XOR U4342 ( .A(n4082), .B(n4083), .Z(n4079) );
  AND U4343 ( .A(n4084), .B(n4085), .Z(n4082) );
  XNOR U4344 ( .A(x[259]), .B(n4083), .Z(n4085) );
  XOR U4345 ( .A(n4086), .B(n4087), .Z(n4083) );
  AND U4346 ( .A(n4088), .B(n4089), .Z(n4086) );
  XNOR U4347 ( .A(x[258]), .B(n4087), .Z(n4089) );
  XOR U4348 ( .A(n4090), .B(n4091), .Z(n4087) );
  AND U4349 ( .A(n4092), .B(n4093), .Z(n4090) );
  XNOR U4350 ( .A(x[257]), .B(n4091), .Z(n4093) );
  XOR U4351 ( .A(n4094), .B(n4095), .Z(n4091) );
  AND U4352 ( .A(n4096), .B(n4097), .Z(n4094) );
  XNOR U4353 ( .A(x[256]), .B(n4095), .Z(n4097) );
  XOR U4354 ( .A(n4098), .B(n4099), .Z(n4095) );
  AND U4355 ( .A(n4100), .B(n4101), .Z(n4098) );
  XNOR U4356 ( .A(x[255]), .B(n4099), .Z(n4101) );
  XOR U4357 ( .A(n4102), .B(n4103), .Z(n4099) );
  AND U4358 ( .A(n4104), .B(n4105), .Z(n4102) );
  XNOR U4359 ( .A(x[254]), .B(n4103), .Z(n4105) );
  XOR U4360 ( .A(n4106), .B(n4107), .Z(n4103) );
  AND U4361 ( .A(n4108), .B(n4109), .Z(n4106) );
  XNOR U4362 ( .A(x[253]), .B(n4107), .Z(n4109) );
  XOR U4363 ( .A(n4110), .B(n4111), .Z(n4107) );
  AND U4364 ( .A(n4112), .B(n4113), .Z(n4110) );
  XNOR U4365 ( .A(x[252]), .B(n4111), .Z(n4113) );
  XOR U4366 ( .A(n4114), .B(n4115), .Z(n4111) );
  AND U4367 ( .A(n4116), .B(n4117), .Z(n4114) );
  XNOR U4368 ( .A(x[251]), .B(n4115), .Z(n4117) );
  XOR U4369 ( .A(n4118), .B(n4119), .Z(n4115) );
  AND U4370 ( .A(n4120), .B(n4121), .Z(n4118) );
  XNOR U4371 ( .A(x[250]), .B(n4119), .Z(n4121) );
  XOR U4372 ( .A(n4122), .B(n4123), .Z(n4119) );
  AND U4373 ( .A(n4124), .B(n4125), .Z(n4122) );
  XNOR U4374 ( .A(x[249]), .B(n4123), .Z(n4125) );
  XOR U4375 ( .A(n4126), .B(n4127), .Z(n4123) );
  AND U4376 ( .A(n4128), .B(n4129), .Z(n4126) );
  XNOR U4377 ( .A(x[248]), .B(n4127), .Z(n4129) );
  XOR U4378 ( .A(n4130), .B(n4131), .Z(n4127) );
  AND U4379 ( .A(n4132), .B(n4133), .Z(n4130) );
  XNOR U4380 ( .A(x[247]), .B(n4131), .Z(n4133) );
  XOR U4381 ( .A(n4134), .B(n4135), .Z(n4131) );
  AND U4382 ( .A(n4136), .B(n4137), .Z(n4134) );
  XNOR U4383 ( .A(x[246]), .B(n4135), .Z(n4137) );
  XOR U4384 ( .A(n4138), .B(n4139), .Z(n4135) );
  AND U4385 ( .A(n4140), .B(n4141), .Z(n4138) );
  XNOR U4386 ( .A(x[245]), .B(n4139), .Z(n4141) );
  XOR U4387 ( .A(n4142), .B(n4143), .Z(n4139) );
  AND U4388 ( .A(n4144), .B(n4145), .Z(n4142) );
  XNOR U4389 ( .A(x[244]), .B(n4143), .Z(n4145) );
  XOR U4390 ( .A(n4146), .B(n4147), .Z(n4143) );
  AND U4391 ( .A(n4148), .B(n4149), .Z(n4146) );
  XNOR U4392 ( .A(x[243]), .B(n4147), .Z(n4149) );
  XOR U4393 ( .A(n4150), .B(n4151), .Z(n4147) );
  AND U4394 ( .A(n4152), .B(n4153), .Z(n4150) );
  XNOR U4395 ( .A(x[242]), .B(n4151), .Z(n4153) );
  XOR U4396 ( .A(n4154), .B(n4155), .Z(n4151) );
  AND U4397 ( .A(n4156), .B(n4157), .Z(n4154) );
  XNOR U4398 ( .A(x[241]), .B(n4155), .Z(n4157) );
  XOR U4399 ( .A(n4158), .B(n4159), .Z(n4155) );
  AND U4400 ( .A(n4160), .B(n4161), .Z(n4158) );
  XNOR U4401 ( .A(x[240]), .B(n4159), .Z(n4161) );
  XOR U4402 ( .A(n4162), .B(n4163), .Z(n4159) );
  AND U4403 ( .A(n4164), .B(n4165), .Z(n4162) );
  XNOR U4404 ( .A(x[239]), .B(n4163), .Z(n4165) );
  XOR U4405 ( .A(n4166), .B(n4167), .Z(n4163) );
  AND U4406 ( .A(n4168), .B(n4169), .Z(n4166) );
  XNOR U4407 ( .A(x[238]), .B(n4167), .Z(n4169) );
  XOR U4408 ( .A(n4170), .B(n4171), .Z(n4167) );
  AND U4409 ( .A(n4172), .B(n4173), .Z(n4170) );
  XNOR U4410 ( .A(x[237]), .B(n4171), .Z(n4173) );
  XOR U4411 ( .A(n4174), .B(n4175), .Z(n4171) );
  AND U4412 ( .A(n4176), .B(n4177), .Z(n4174) );
  XNOR U4413 ( .A(x[236]), .B(n4175), .Z(n4177) );
  XOR U4414 ( .A(n4178), .B(n4179), .Z(n4175) );
  AND U4415 ( .A(n4180), .B(n4181), .Z(n4178) );
  XNOR U4416 ( .A(x[235]), .B(n4179), .Z(n4181) );
  XOR U4417 ( .A(n4182), .B(n4183), .Z(n4179) );
  AND U4418 ( .A(n4184), .B(n4185), .Z(n4182) );
  XNOR U4419 ( .A(x[234]), .B(n4183), .Z(n4185) );
  XOR U4420 ( .A(n4186), .B(n4187), .Z(n4183) );
  AND U4421 ( .A(n4188), .B(n4189), .Z(n4186) );
  XNOR U4422 ( .A(x[233]), .B(n4187), .Z(n4189) );
  XOR U4423 ( .A(n4190), .B(n4191), .Z(n4187) );
  AND U4424 ( .A(n4192), .B(n4193), .Z(n4190) );
  XNOR U4425 ( .A(x[232]), .B(n4191), .Z(n4193) );
  XOR U4426 ( .A(n4194), .B(n4195), .Z(n4191) );
  AND U4427 ( .A(n4196), .B(n4197), .Z(n4194) );
  XNOR U4428 ( .A(x[231]), .B(n4195), .Z(n4197) );
  XOR U4429 ( .A(n4198), .B(n4199), .Z(n4195) );
  AND U4430 ( .A(n4200), .B(n4201), .Z(n4198) );
  XNOR U4431 ( .A(x[230]), .B(n4199), .Z(n4201) );
  XOR U4432 ( .A(n4202), .B(n4203), .Z(n4199) );
  AND U4433 ( .A(n4204), .B(n4205), .Z(n4202) );
  XNOR U4434 ( .A(x[229]), .B(n4203), .Z(n4205) );
  XOR U4435 ( .A(n4206), .B(n4207), .Z(n4203) );
  AND U4436 ( .A(n4208), .B(n4209), .Z(n4206) );
  XNOR U4437 ( .A(x[228]), .B(n4207), .Z(n4209) );
  XOR U4438 ( .A(n4210), .B(n4211), .Z(n4207) );
  AND U4439 ( .A(n4212), .B(n4213), .Z(n4210) );
  XNOR U4440 ( .A(x[227]), .B(n4211), .Z(n4213) );
  XOR U4441 ( .A(n4214), .B(n4215), .Z(n4211) );
  AND U4442 ( .A(n4216), .B(n4217), .Z(n4214) );
  XNOR U4443 ( .A(x[226]), .B(n4215), .Z(n4217) );
  XOR U4444 ( .A(n4218), .B(n4219), .Z(n4215) );
  AND U4445 ( .A(n4220), .B(n4221), .Z(n4218) );
  XNOR U4446 ( .A(x[225]), .B(n4219), .Z(n4221) );
  XOR U4447 ( .A(n4222), .B(n4223), .Z(n4219) );
  AND U4448 ( .A(n4224), .B(n4225), .Z(n4222) );
  XNOR U4449 ( .A(x[224]), .B(n4223), .Z(n4225) );
  XOR U4450 ( .A(n4226), .B(n4227), .Z(n4223) );
  AND U4451 ( .A(n4228), .B(n4229), .Z(n4226) );
  XNOR U4452 ( .A(x[223]), .B(n4227), .Z(n4229) );
  XOR U4453 ( .A(n4230), .B(n4231), .Z(n4227) );
  AND U4454 ( .A(n4232), .B(n4233), .Z(n4230) );
  XNOR U4455 ( .A(x[222]), .B(n4231), .Z(n4233) );
  XOR U4456 ( .A(n4234), .B(n4235), .Z(n4231) );
  AND U4457 ( .A(n4236), .B(n4237), .Z(n4234) );
  XNOR U4458 ( .A(x[221]), .B(n4235), .Z(n4237) );
  XOR U4459 ( .A(n4238), .B(n4239), .Z(n4235) );
  AND U4460 ( .A(n4240), .B(n4241), .Z(n4238) );
  XNOR U4461 ( .A(x[220]), .B(n4239), .Z(n4241) );
  XOR U4462 ( .A(n4242), .B(n4243), .Z(n4239) );
  AND U4463 ( .A(n4244), .B(n4245), .Z(n4242) );
  XNOR U4464 ( .A(x[219]), .B(n4243), .Z(n4245) );
  XOR U4465 ( .A(n4246), .B(n4247), .Z(n4243) );
  AND U4466 ( .A(n4248), .B(n4249), .Z(n4246) );
  XNOR U4467 ( .A(x[218]), .B(n4247), .Z(n4249) );
  XOR U4468 ( .A(n4250), .B(n4251), .Z(n4247) );
  AND U4469 ( .A(n4252), .B(n4253), .Z(n4250) );
  XNOR U4470 ( .A(x[217]), .B(n4251), .Z(n4253) );
  XOR U4471 ( .A(n4254), .B(n4255), .Z(n4251) );
  AND U4472 ( .A(n4256), .B(n4257), .Z(n4254) );
  XNOR U4473 ( .A(x[216]), .B(n4255), .Z(n4257) );
  XOR U4474 ( .A(n4258), .B(n4259), .Z(n4255) );
  AND U4475 ( .A(n4260), .B(n4261), .Z(n4258) );
  XNOR U4476 ( .A(x[215]), .B(n4259), .Z(n4261) );
  XOR U4477 ( .A(n4262), .B(n4263), .Z(n4259) );
  AND U4478 ( .A(n4264), .B(n4265), .Z(n4262) );
  XNOR U4479 ( .A(x[214]), .B(n4263), .Z(n4265) );
  XOR U4480 ( .A(n4266), .B(n4267), .Z(n4263) );
  AND U4481 ( .A(n4268), .B(n4269), .Z(n4266) );
  XNOR U4482 ( .A(x[213]), .B(n4267), .Z(n4269) );
  XOR U4483 ( .A(n4270), .B(n4271), .Z(n4267) );
  AND U4484 ( .A(n4272), .B(n4273), .Z(n4270) );
  XNOR U4485 ( .A(x[212]), .B(n4271), .Z(n4273) );
  XOR U4486 ( .A(n4274), .B(n4275), .Z(n4271) );
  AND U4487 ( .A(n4276), .B(n4277), .Z(n4274) );
  XNOR U4488 ( .A(x[211]), .B(n4275), .Z(n4277) );
  XOR U4489 ( .A(n4278), .B(n4279), .Z(n4275) );
  AND U4490 ( .A(n4280), .B(n4281), .Z(n4278) );
  XNOR U4491 ( .A(x[210]), .B(n4279), .Z(n4281) );
  XOR U4492 ( .A(n4282), .B(n4283), .Z(n4279) );
  AND U4493 ( .A(n4284), .B(n4285), .Z(n4282) );
  XNOR U4494 ( .A(x[209]), .B(n4283), .Z(n4285) );
  XOR U4495 ( .A(n4286), .B(n4287), .Z(n4283) );
  AND U4496 ( .A(n4288), .B(n4289), .Z(n4286) );
  XNOR U4497 ( .A(x[208]), .B(n4287), .Z(n4289) );
  XOR U4498 ( .A(n4290), .B(n4291), .Z(n4287) );
  AND U4499 ( .A(n4292), .B(n4293), .Z(n4290) );
  XNOR U4500 ( .A(x[207]), .B(n4291), .Z(n4293) );
  XOR U4501 ( .A(n4294), .B(n4295), .Z(n4291) );
  AND U4502 ( .A(n4296), .B(n4297), .Z(n4294) );
  XNOR U4503 ( .A(x[206]), .B(n4295), .Z(n4297) );
  XOR U4504 ( .A(n4298), .B(n4299), .Z(n4295) );
  AND U4505 ( .A(n4300), .B(n4301), .Z(n4298) );
  XNOR U4506 ( .A(x[205]), .B(n4299), .Z(n4301) );
  XOR U4507 ( .A(n4302), .B(n4303), .Z(n4299) );
  AND U4508 ( .A(n4304), .B(n4305), .Z(n4302) );
  XNOR U4509 ( .A(x[204]), .B(n4303), .Z(n4305) );
  XOR U4510 ( .A(n4306), .B(n4307), .Z(n4303) );
  AND U4511 ( .A(n4308), .B(n4309), .Z(n4306) );
  XNOR U4512 ( .A(x[203]), .B(n4307), .Z(n4309) );
  XOR U4513 ( .A(n4310), .B(n4311), .Z(n4307) );
  AND U4514 ( .A(n4312), .B(n4313), .Z(n4310) );
  XNOR U4515 ( .A(x[202]), .B(n4311), .Z(n4313) );
  XOR U4516 ( .A(n4314), .B(n4315), .Z(n4311) );
  AND U4517 ( .A(n4316), .B(n4317), .Z(n4314) );
  XNOR U4518 ( .A(x[201]), .B(n4315), .Z(n4317) );
  XOR U4519 ( .A(n4318), .B(n4319), .Z(n4315) );
  AND U4520 ( .A(n4320), .B(n4321), .Z(n4318) );
  XNOR U4521 ( .A(x[200]), .B(n4319), .Z(n4321) );
  XOR U4522 ( .A(n4322), .B(n4323), .Z(n4319) );
  AND U4523 ( .A(n4324), .B(n4325), .Z(n4322) );
  XNOR U4524 ( .A(x[199]), .B(n4323), .Z(n4325) );
  XOR U4525 ( .A(n4326), .B(n4327), .Z(n4323) );
  AND U4526 ( .A(n4328), .B(n4329), .Z(n4326) );
  XNOR U4527 ( .A(x[198]), .B(n4327), .Z(n4329) );
  XOR U4528 ( .A(n4330), .B(n4331), .Z(n4327) );
  AND U4529 ( .A(n4332), .B(n4333), .Z(n4330) );
  XNOR U4530 ( .A(x[197]), .B(n4331), .Z(n4333) );
  XOR U4531 ( .A(n4334), .B(n4335), .Z(n4331) );
  AND U4532 ( .A(n4336), .B(n4337), .Z(n4334) );
  XNOR U4533 ( .A(x[196]), .B(n4335), .Z(n4337) );
  XOR U4534 ( .A(n4338), .B(n4339), .Z(n4335) );
  AND U4535 ( .A(n4340), .B(n4341), .Z(n4338) );
  XNOR U4536 ( .A(x[195]), .B(n4339), .Z(n4341) );
  XOR U4537 ( .A(n4342), .B(n4343), .Z(n4339) );
  AND U4538 ( .A(n4344), .B(n4345), .Z(n4342) );
  XNOR U4539 ( .A(x[194]), .B(n4343), .Z(n4345) );
  XOR U4540 ( .A(n4346), .B(n4347), .Z(n4343) );
  AND U4541 ( .A(n4348), .B(n4349), .Z(n4346) );
  XNOR U4542 ( .A(x[193]), .B(n4347), .Z(n4349) );
  XOR U4543 ( .A(n4350), .B(n4351), .Z(n4347) );
  AND U4544 ( .A(n4352), .B(n4353), .Z(n4350) );
  XNOR U4545 ( .A(x[192]), .B(n4351), .Z(n4353) );
  XOR U4546 ( .A(n4354), .B(n4355), .Z(n4351) );
  AND U4547 ( .A(n4356), .B(n4357), .Z(n4354) );
  XNOR U4548 ( .A(x[191]), .B(n4355), .Z(n4357) );
  XOR U4549 ( .A(n4358), .B(n4359), .Z(n4355) );
  AND U4550 ( .A(n4360), .B(n4361), .Z(n4358) );
  XNOR U4551 ( .A(x[190]), .B(n4359), .Z(n4361) );
  XOR U4552 ( .A(n4362), .B(n4363), .Z(n4359) );
  AND U4553 ( .A(n4364), .B(n4365), .Z(n4362) );
  XNOR U4554 ( .A(x[189]), .B(n4363), .Z(n4365) );
  XOR U4555 ( .A(n4366), .B(n4367), .Z(n4363) );
  AND U4556 ( .A(n4368), .B(n4369), .Z(n4366) );
  XNOR U4557 ( .A(x[188]), .B(n4367), .Z(n4369) );
  XOR U4558 ( .A(n4370), .B(n4371), .Z(n4367) );
  AND U4559 ( .A(n4372), .B(n4373), .Z(n4370) );
  XNOR U4560 ( .A(x[187]), .B(n4371), .Z(n4373) );
  XOR U4561 ( .A(n4374), .B(n4375), .Z(n4371) );
  AND U4562 ( .A(n4376), .B(n4377), .Z(n4374) );
  XNOR U4563 ( .A(x[186]), .B(n4375), .Z(n4377) );
  XOR U4564 ( .A(n4378), .B(n4379), .Z(n4375) );
  AND U4565 ( .A(n4380), .B(n4381), .Z(n4378) );
  XNOR U4566 ( .A(x[185]), .B(n4379), .Z(n4381) );
  XOR U4567 ( .A(n4382), .B(n4383), .Z(n4379) );
  AND U4568 ( .A(n4384), .B(n4385), .Z(n4382) );
  XNOR U4569 ( .A(x[184]), .B(n4383), .Z(n4385) );
  XOR U4570 ( .A(n4386), .B(n4387), .Z(n4383) );
  AND U4571 ( .A(n4388), .B(n4389), .Z(n4386) );
  XNOR U4572 ( .A(x[183]), .B(n4387), .Z(n4389) );
  XOR U4573 ( .A(n4390), .B(n4391), .Z(n4387) );
  AND U4574 ( .A(n4392), .B(n4393), .Z(n4390) );
  XNOR U4575 ( .A(x[182]), .B(n4391), .Z(n4393) );
  XOR U4576 ( .A(n4394), .B(n4395), .Z(n4391) );
  AND U4577 ( .A(n4396), .B(n4397), .Z(n4394) );
  XNOR U4578 ( .A(x[181]), .B(n4395), .Z(n4397) );
  XOR U4579 ( .A(n4398), .B(n4399), .Z(n4395) );
  AND U4580 ( .A(n4400), .B(n4401), .Z(n4398) );
  XNOR U4581 ( .A(x[180]), .B(n4399), .Z(n4401) );
  XOR U4582 ( .A(n4402), .B(n4403), .Z(n4399) );
  AND U4583 ( .A(n4404), .B(n4405), .Z(n4402) );
  XNOR U4584 ( .A(x[179]), .B(n4403), .Z(n4405) );
  XOR U4585 ( .A(n4406), .B(n4407), .Z(n4403) );
  AND U4586 ( .A(n4408), .B(n4409), .Z(n4406) );
  XNOR U4587 ( .A(x[178]), .B(n4407), .Z(n4409) );
  XOR U4588 ( .A(n4410), .B(n4411), .Z(n4407) );
  AND U4589 ( .A(n4412), .B(n4413), .Z(n4410) );
  XNOR U4590 ( .A(x[177]), .B(n4411), .Z(n4413) );
  XOR U4591 ( .A(n4414), .B(n4415), .Z(n4411) );
  AND U4592 ( .A(n4416), .B(n4417), .Z(n4414) );
  XNOR U4593 ( .A(x[176]), .B(n4415), .Z(n4417) );
  XOR U4594 ( .A(n4418), .B(n4419), .Z(n4415) );
  AND U4595 ( .A(n4420), .B(n4421), .Z(n4418) );
  XNOR U4596 ( .A(x[175]), .B(n4419), .Z(n4421) );
  XOR U4597 ( .A(n4422), .B(n4423), .Z(n4419) );
  AND U4598 ( .A(n4424), .B(n4425), .Z(n4422) );
  XNOR U4599 ( .A(x[174]), .B(n4423), .Z(n4425) );
  XOR U4600 ( .A(n4426), .B(n4427), .Z(n4423) );
  AND U4601 ( .A(n4428), .B(n4429), .Z(n4426) );
  XNOR U4602 ( .A(x[173]), .B(n4427), .Z(n4429) );
  XOR U4603 ( .A(n4430), .B(n4431), .Z(n4427) );
  AND U4604 ( .A(n4432), .B(n4433), .Z(n4430) );
  XNOR U4605 ( .A(x[172]), .B(n4431), .Z(n4433) );
  XOR U4606 ( .A(n4434), .B(n4435), .Z(n4431) );
  AND U4607 ( .A(n4436), .B(n4437), .Z(n4434) );
  XNOR U4608 ( .A(x[171]), .B(n4435), .Z(n4437) );
  XOR U4609 ( .A(n4438), .B(n4439), .Z(n4435) );
  AND U4610 ( .A(n4440), .B(n4441), .Z(n4438) );
  XNOR U4611 ( .A(x[170]), .B(n4439), .Z(n4441) );
  XOR U4612 ( .A(n4442), .B(n4443), .Z(n4439) );
  AND U4613 ( .A(n4444), .B(n4445), .Z(n4442) );
  XNOR U4614 ( .A(x[169]), .B(n4443), .Z(n4445) );
  XOR U4615 ( .A(n4446), .B(n4447), .Z(n4443) );
  AND U4616 ( .A(n4448), .B(n4449), .Z(n4446) );
  XNOR U4617 ( .A(x[168]), .B(n4447), .Z(n4449) );
  XOR U4618 ( .A(n4450), .B(n4451), .Z(n4447) );
  AND U4619 ( .A(n4452), .B(n4453), .Z(n4450) );
  XNOR U4620 ( .A(x[167]), .B(n4451), .Z(n4453) );
  XOR U4621 ( .A(n4454), .B(n4455), .Z(n4451) );
  AND U4622 ( .A(n4456), .B(n4457), .Z(n4454) );
  XNOR U4623 ( .A(x[166]), .B(n4455), .Z(n4457) );
  XOR U4624 ( .A(n4458), .B(n4459), .Z(n4455) );
  AND U4625 ( .A(n4460), .B(n4461), .Z(n4458) );
  XNOR U4626 ( .A(x[165]), .B(n4459), .Z(n4461) );
  XOR U4627 ( .A(n4462), .B(n4463), .Z(n4459) );
  AND U4628 ( .A(n4464), .B(n4465), .Z(n4462) );
  XNOR U4629 ( .A(x[164]), .B(n4463), .Z(n4465) );
  XOR U4630 ( .A(n4466), .B(n4467), .Z(n4463) );
  AND U4631 ( .A(n4468), .B(n4469), .Z(n4466) );
  XNOR U4632 ( .A(x[163]), .B(n4467), .Z(n4469) );
  XOR U4633 ( .A(n4470), .B(n4471), .Z(n4467) );
  AND U4634 ( .A(n4472), .B(n4473), .Z(n4470) );
  XNOR U4635 ( .A(x[162]), .B(n4471), .Z(n4473) );
  XOR U4636 ( .A(n4474), .B(n4475), .Z(n4471) );
  AND U4637 ( .A(n4476), .B(n4477), .Z(n4474) );
  XNOR U4638 ( .A(x[161]), .B(n4475), .Z(n4477) );
  XOR U4639 ( .A(n4478), .B(n4479), .Z(n4475) );
  AND U4640 ( .A(n4480), .B(n4481), .Z(n4478) );
  XNOR U4641 ( .A(x[160]), .B(n4479), .Z(n4481) );
  XOR U4642 ( .A(n4482), .B(n4483), .Z(n4479) );
  AND U4643 ( .A(n4484), .B(n4485), .Z(n4482) );
  XNOR U4644 ( .A(x[159]), .B(n4483), .Z(n4485) );
  XOR U4645 ( .A(n4486), .B(n4487), .Z(n4483) );
  AND U4646 ( .A(n4488), .B(n4489), .Z(n4486) );
  XNOR U4647 ( .A(x[158]), .B(n4487), .Z(n4489) );
  XOR U4648 ( .A(n4490), .B(n4491), .Z(n4487) );
  AND U4649 ( .A(n4492), .B(n4493), .Z(n4490) );
  XNOR U4650 ( .A(x[157]), .B(n4491), .Z(n4493) );
  XOR U4651 ( .A(n4494), .B(n4495), .Z(n4491) );
  AND U4652 ( .A(n4496), .B(n4497), .Z(n4494) );
  XNOR U4653 ( .A(x[156]), .B(n4495), .Z(n4497) );
  XOR U4654 ( .A(n4498), .B(n4499), .Z(n4495) );
  AND U4655 ( .A(n4500), .B(n4501), .Z(n4498) );
  XNOR U4656 ( .A(x[155]), .B(n4499), .Z(n4501) );
  XOR U4657 ( .A(n4502), .B(n4503), .Z(n4499) );
  AND U4658 ( .A(n4504), .B(n4505), .Z(n4502) );
  XNOR U4659 ( .A(x[154]), .B(n4503), .Z(n4505) );
  XOR U4660 ( .A(n4506), .B(n4507), .Z(n4503) );
  AND U4661 ( .A(n4508), .B(n4509), .Z(n4506) );
  XNOR U4662 ( .A(x[153]), .B(n4507), .Z(n4509) );
  XOR U4663 ( .A(n4510), .B(n4511), .Z(n4507) );
  AND U4664 ( .A(n4512), .B(n4513), .Z(n4510) );
  XNOR U4665 ( .A(x[152]), .B(n4511), .Z(n4513) );
  XOR U4666 ( .A(n4514), .B(n4515), .Z(n4511) );
  AND U4667 ( .A(n4516), .B(n4517), .Z(n4514) );
  XNOR U4668 ( .A(x[151]), .B(n4515), .Z(n4517) );
  XOR U4669 ( .A(n4518), .B(n4519), .Z(n4515) );
  AND U4670 ( .A(n4520), .B(n4521), .Z(n4518) );
  XNOR U4671 ( .A(x[150]), .B(n4519), .Z(n4521) );
  XOR U4672 ( .A(n4522), .B(n4523), .Z(n4519) );
  AND U4673 ( .A(n4524), .B(n4525), .Z(n4522) );
  XNOR U4674 ( .A(x[149]), .B(n4523), .Z(n4525) );
  XOR U4675 ( .A(n4526), .B(n4527), .Z(n4523) );
  AND U4676 ( .A(n4528), .B(n4529), .Z(n4526) );
  XNOR U4677 ( .A(x[148]), .B(n4527), .Z(n4529) );
  XOR U4678 ( .A(n4530), .B(n4531), .Z(n4527) );
  AND U4679 ( .A(n4532), .B(n4533), .Z(n4530) );
  XNOR U4680 ( .A(x[147]), .B(n4531), .Z(n4533) );
  XOR U4681 ( .A(n4534), .B(n4535), .Z(n4531) );
  AND U4682 ( .A(n4536), .B(n4537), .Z(n4534) );
  XNOR U4683 ( .A(x[146]), .B(n4535), .Z(n4537) );
  XOR U4684 ( .A(n4538), .B(n4539), .Z(n4535) );
  AND U4685 ( .A(n4540), .B(n4541), .Z(n4538) );
  XNOR U4686 ( .A(x[145]), .B(n4539), .Z(n4541) );
  XOR U4687 ( .A(n4542), .B(n4543), .Z(n4539) );
  AND U4688 ( .A(n4544), .B(n4545), .Z(n4542) );
  XNOR U4689 ( .A(x[144]), .B(n4543), .Z(n4545) );
  XOR U4690 ( .A(n4546), .B(n4547), .Z(n4543) );
  AND U4691 ( .A(n4548), .B(n4549), .Z(n4546) );
  XNOR U4692 ( .A(x[143]), .B(n4547), .Z(n4549) );
  XOR U4693 ( .A(n4550), .B(n4551), .Z(n4547) );
  AND U4694 ( .A(n4552), .B(n4553), .Z(n4550) );
  XNOR U4695 ( .A(x[142]), .B(n4551), .Z(n4553) );
  XOR U4696 ( .A(n4554), .B(n4555), .Z(n4551) );
  AND U4697 ( .A(n4556), .B(n4557), .Z(n4554) );
  XNOR U4698 ( .A(x[141]), .B(n4555), .Z(n4557) );
  XOR U4699 ( .A(n4558), .B(n4559), .Z(n4555) );
  AND U4700 ( .A(n4560), .B(n4561), .Z(n4558) );
  XNOR U4701 ( .A(x[140]), .B(n4559), .Z(n4561) );
  XOR U4702 ( .A(n4562), .B(n4563), .Z(n4559) );
  AND U4703 ( .A(n4564), .B(n4565), .Z(n4562) );
  XNOR U4704 ( .A(x[139]), .B(n4563), .Z(n4565) );
  XOR U4705 ( .A(n4566), .B(n4567), .Z(n4563) );
  AND U4706 ( .A(n4568), .B(n4569), .Z(n4566) );
  XNOR U4707 ( .A(x[138]), .B(n4567), .Z(n4569) );
  XOR U4708 ( .A(n4570), .B(n4571), .Z(n4567) );
  AND U4709 ( .A(n4572), .B(n4573), .Z(n4570) );
  XNOR U4710 ( .A(x[137]), .B(n4571), .Z(n4573) );
  XOR U4711 ( .A(n4574), .B(n4575), .Z(n4571) );
  AND U4712 ( .A(n4576), .B(n4577), .Z(n4574) );
  XNOR U4713 ( .A(x[136]), .B(n4575), .Z(n4577) );
  XOR U4714 ( .A(n4578), .B(n4579), .Z(n4575) );
  AND U4715 ( .A(n4580), .B(n4581), .Z(n4578) );
  XNOR U4716 ( .A(x[135]), .B(n4579), .Z(n4581) );
  XOR U4717 ( .A(n4582), .B(n4583), .Z(n4579) );
  AND U4718 ( .A(n4584), .B(n4585), .Z(n4582) );
  XNOR U4719 ( .A(x[134]), .B(n4583), .Z(n4585) );
  XOR U4720 ( .A(n4586), .B(n4587), .Z(n4583) );
  AND U4721 ( .A(n4588), .B(n4589), .Z(n4586) );
  XNOR U4722 ( .A(x[133]), .B(n4587), .Z(n4589) );
  XOR U4723 ( .A(n4590), .B(n4591), .Z(n4587) );
  AND U4724 ( .A(n4592), .B(n4593), .Z(n4590) );
  XNOR U4725 ( .A(x[132]), .B(n4591), .Z(n4593) );
  XOR U4726 ( .A(n4594), .B(n4595), .Z(n4591) );
  AND U4727 ( .A(n4596), .B(n4597), .Z(n4594) );
  XNOR U4728 ( .A(x[131]), .B(n4595), .Z(n4597) );
  XOR U4729 ( .A(n4598), .B(n4599), .Z(n4595) );
  AND U4730 ( .A(n4600), .B(n4601), .Z(n4598) );
  XNOR U4731 ( .A(x[130]), .B(n4599), .Z(n4601) );
  XOR U4732 ( .A(n4602), .B(n4603), .Z(n4599) );
  AND U4733 ( .A(n4604), .B(n4605), .Z(n4602) );
  XNOR U4734 ( .A(x[129]), .B(n4603), .Z(n4605) );
  XOR U4735 ( .A(n4606), .B(n4607), .Z(n4603) );
  AND U4736 ( .A(n4608), .B(n4609), .Z(n4606) );
  XNOR U4737 ( .A(x[128]), .B(n4607), .Z(n4609) );
  XOR U4738 ( .A(n4610), .B(n4611), .Z(n4607) );
  AND U4739 ( .A(n4612), .B(n4613), .Z(n4610) );
  XNOR U4740 ( .A(x[127]), .B(n4611), .Z(n4613) );
  XOR U4741 ( .A(n4614), .B(n4615), .Z(n4611) );
  AND U4742 ( .A(n4616), .B(n4617), .Z(n4614) );
  XNOR U4743 ( .A(x[126]), .B(n4615), .Z(n4617) );
  XOR U4744 ( .A(n4618), .B(n4619), .Z(n4615) );
  AND U4745 ( .A(n4620), .B(n4621), .Z(n4618) );
  XNOR U4746 ( .A(x[125]), .B(n4619), .Z(n4621) );
  XOR U4747 ( .A(n4622), .B(n4623), .Z(n4619) );
  AND U4748 ( .A(n4624), .B(n4625), .Z(n4622) );
  XNOR U4749 ( .A(x[124]), .B(n4623), .Z(n4625) );
  XOR U4750 ( .A(n4626), .B(n4627), .Z(n4623) );
  AND U4751 ( .A(n4628), .B(n4629), .Z(n4626) );
  XNOR U4752 ( .A(x[123]), .B(n4627), .Z(n4629) );
  XOR U4753 ( .A(n4630), .B(n4631), .Z(n4627) );
  AND U4754 ( .A(n4632), .B(n4633), .Z(n4630) );
  XNOR U4755 ( .A(x[122]), .B(n4631), .Z(n4633) );
  XOR U4756 ( .A(n4634), .B(n4635), .Z(n4631) );
  AND U4757 ( .A(n4636), .B(n4637), .Z(n4634) );
  XNOR U4758 ( .A(x[121]), .B(n4635), .Z(n4637) );
  XOR U4759 ( .A(n4638), .B(n4639), .Z(n4635) );
  AND U4760 ( .A(n4640), .B(n4641), .Z(n4638) );
  XNOR U4761 ( .A(x[120]), .B(n4639), .Z(n4641) );
  XOR U4762 ( .A(n4642), .B(n4643), .Z(n4639) );
  AND U4763 ( .A(n4644), .B(n4645), .Z(n4642) );
  XNOR U4764 ( .A(x[119]), .B(n4643), .Z(n4645) );
  XOR U4765 ( .A(n4646), .B(n4647), .Z(n4643) );
  AND U4766 ( .A(n4648), .B(n4649), .Z(n4646) );
  XNOR U4767 ( .A(x[118]), .B(n4647), .Z(n4649) );
  XOR U4768 ( .A(n4650), .B(n4651), .Z(n4647) );
  AND U4769 ( .A(n4652), .B(n4653), .Z(n4650) );
  XNOR U4770 ( .A(x[117]), .B(n4651), .Z(n4653) );
  XOR U4771 ( .A(n4654), .B(n4655), .Z(n4651) );
  AND U4772 ( .A(n4656), .B(n4657), .Z(n4654) );
  XNOR U4773 ( .A(x[116]), .B(n4655), .Z(n4657) );
  XOR U4774 ( .A(n4658), .B(n4659), .Z(n4655) );
  AND U4775 ( .A(n4660), .B(n4661), .Z(n4658) );
  XNOR U4776 ( .A(x[115]), .B(n4659), .Z(n4661) );
  XOR U4777 ( .A(n4662), .B(n4663), .Z(n4659) );
  AND U4778 ( .A(n4664), .B(n4665), .Z(n4662) );
  XNOR U4779 ( .A(x[114]), .B(n4663), .Z(n4665) );
  XOR U4780 ( .A(n4666), .B(n4667), .Z(n4663) );
  AND U4781 ( .A(n4668), .B(n4669), .Z(n4666) );
  XNOR U4782 ( .A(x[113]), .B(n4667), .Z(n4669) );
  XOR U4783 ( .A(n4670), .B(n4671), .Z(n4667) );
  AND U4784 ( .A(n4672), .B(n4673), .Z(n4670) );
  XNOR U4785 ( .A(x[112]), .B(n4671), .Z(n4673) );
  XOR U4786 ( .A(n4674), .B(n4675), .Z(n4671) );
  AND U4787 ( .A(n4676), .B(n4677), .Z(n4674) );
  XNOR U4788 ( .A(x[111]), .B(n4675), .Z(n4677) );
  XOR U4789 ( .A(n4678), .B(n4679), .Z(n4675) );
  AND U4790 ( .A(n4680), .B(n4681), .Z(n4678) );
  XNOR U4791 ( .A(x[110]), .B(n4679), .Z(n4681) );
  XOR U4792 ( .A(n4682), .B(n4683), .Z(n4679) );
  AND U4793 ( .A(n4684), .B(n4685), .Z(n4682) );
  XNOR U4794 ( .A(x[109]), .B(n4683), .Z(n4685) );
  XOR U4795 ( .A(n4686), .B(n4687), .Z(n4683) );
  AND U4796 ( .A(n4688), .B(n4689), .Z(n4686) );
  XNOR U4797 ( .A(x[108]), .B(n4687), .Z(n4689) );
  XOR U4798 ( .A(n4690), .B(n4691), .Z(n4687) );
  AND U4799 ( .A(n4692), .B(n4693), .Z(n4690) );
  XNOR U4800 ( .A(x[107]), .B(n4691), .Z(n4693) );
  XOR U4801 ( .A(n4694), .B(n4695), .Z(n4691) );
  AND U4802 ( .A(n4696), .B(n4697), .Z(n4694) );
  XNOR U4803 ( .A(x[106]), .B(n4695), .Z(n4697) );
  XOR U4804 ( .A(n4698), .B(n4699), .Z(n4695) );
  AND U4805 ( .A(n4700), .B(n4701), .Z(n4698) );
  XNOR U4806 ( .A(x[105]), .B(n4699), .Z(n4701) );
  XOR U4807 ( .A(n4702), .B(n4703), .Z(n4699) );
  AND U4808 ( .A(n4704), .B(n4705), .Z(n4702) );
  XNOR U4809 ( .A(x[104]), .B(n4703), .Z(n4705) );
  XOR U4810 ( .A(n4706), .B(n4707), .Z(n4703) );
  AND U4811 ( .A(n4708), .B(n4709), .Z(n4706) );
  XNOR U4812 ( .A(x[103]), .B(n4707), .Z(n4709) );
  XOR U4813 ( .A(n4710), .B(n4711), .Z(n4707) );
  AND U4814 ( .A(n4712), .B(n4713), .Z(n4710) );
  XNOR U4815 ( .A(x[102]), .B(n4711), .Z(n4713) );
  XOR U4816 ( .A(n4714), .B(n4715), .Z(n4711) );
  AND U4817 ( .A(n4716), .B(n4717), .Z(n4714) );
  XNOR U4818 ( .A(x[101]), .B(n4715), .Z(n4717) );
  XOR U4819 ( .A(n4718), .B(n4719), .Z(n4715) );
  AND U4820 ( .A(n4720), .B(n4721), .Z(n4718) );
  XNOR U4821 ( .A(x[100]), .B(n4719), .Z(n4721) );
  XOR U4822 ( .A(n4722), .B(n4723), .Z(n4719) );
  AND U4823 ( .A(n4724), .B(n4725), .Z(n4722) );
  XNOR U4824 ( .A(x[99]), .B(n4723), .Z(n4725) );
  XOR U4825 ( .A(n4726), .B(n4727), .Z(n4723) );
  AND U4826 ( .A(n4728), .B(n4729), .Z(n4726) );
  XNOR U4827 ( .A(x[98]), .B(n4727), .Z(n4729) );
  XOR U4828 ( .A(n4730), .B(n4731), .Z(n4727) );
  AND U4829 ( .A(n4732), .B(n4733), .Z(n4730) );
  XNOR U4830 ( .A(x[97]), .B(n4731), .Z(n4733) );
  XOR U4831 ( .A(n4734), .B(n4735), .Z(n4731) );
  AND U4832 ( .A(n4736), .B(n4737), .Z(n4734) );
  XNOR U4833 ( .A(x[96]), .B(n4735), .Z(n4737) );
  XOR U4834 ( .A(n4738), .B(n4739), .Z(n4735) );
  AND U4835 ( .A(n4740), .B(n4741), .Z(n4738) );
  XNOR U4836 ( .A(x[95]), .B(n4739), .Z(n4741) );
  XOR U4837 ( .A(n4742), .B(n4743), .Z(n4739) );
  AND U4838 ( .A(n4744), .B(n4745), .Z(n4742) );
  XNOR U4839 ( .A(x[94]), .B(n4743), .Z(n4745) );
  XOR U4840 ( .A(n4746), .B(n4747), .Z(n4743) );
  AND U4841 ( .A(n4748), .B(n4749), .Z(n4746) );
  XNOR U4842 ( .A(x[93]), .B(n4747), .Z(n4749) );
  XOR U4843 ( .A(n4750), .B(n4751), .Z(n4747) );
  AND U4844 ( .A(n4752), .B(n4753), .Z(n4750) );
  XNOR U4845 ( .A(x[92]), .B(n4751), .Z(n4753) );
  XOR U4846 ( .A(n4754), .B(n4755), .Z(n4751) );
  AND U4847 ( .A(n4756), .B(n4757), .Z(n4754) );
  XNOR U4848 ( .A(x[91]), .B(n4755), .Z(n4757) );
  XOR U4849 ( .A(n4758), .B(n4759), .Z(n4755) );
  AND U4850 ( .A(n4760), .B(n4761), .Z(n4758) );
  XNOR U4851 ( .A(x[90]), .B(n4759), .Z(n4761) );
  XOR U4852 ( .A(n4762), .B(n4763), .Z(n4759) );
  AND U4853 ( .A(n4764), .B(n4765), .Z(n4762) );
  XNOR U4854 ( .A(x[89]), .B(n4763), .Z(n4765) );
  XOR U4855 ( .A(n4766), .B(n4767), .Z(n4763) );
  AND U4856 ( .A(n4768), .B(n4769), .Z(n4766) );
  XNOR U4857 ( .A(x[88]), .B(n4767), .Z(n4769) );
  XOR U4858 ( .A(n4770), .B(n4771), .Z(n4767) );
  AND U4859 ( .A(n4772), .B(n4773), .Z(n4770) );
  XNOR U4860 ( .A(x[87]), .B(n4771), .Z(n4773) );
  XOR U4861 ( .A(n4774), .B(n4775), .Z(n4771) );
  AND U4862 ( .A(n4776), .B(n4777), .Z(n4774) );
  XNOR U4863 ( .A(x[86]), .B(n4775), .Z(n4777) );
  XOR U4864 ( .A(n4778), .B(n4779), .Z(n4775) );
  AND U4865 ( .A(n4780), .B(n4781), .Z(n4778) );
  XNOR U4866 ( .A(x[85]), .B(n4779), .Z(n4781) );
  XOR U4867 ( .A(n4782), .B(n4783), .Z(n4779) );
  AND U4868 ( .A(n4784), .B(n4785), .Z(n4782) );
  XNOR U4869 ( .A(x[84]), .B(n4783), .Z(n4785) );
  XOR U4870 ( .A(n4786), .B(n4787), .Z(n4783) );
  AND U4871 ( .A(n4788), .B(n4789), .Z(n4786) );
  XNOR U4872 ( .A(x[83]), .B(n4787), .Z(n4789) );
  XOR U4873 ( .A(n4790), .B(n4791), .Z(n4787) );
  AND U4874 ( .A(n4792), .B(n4793), .Z(n4790) );
  XNOR U4875 ( .A(x[82]), .B(n4791), .Z(n4793) );
  XOR U4876 ( .A(n4794), .B(n4795), .Z(n4791) );
  AND U4877 ( .A(n4796), .B(n4797), .Z(n4794) );
  XNOR U4878 ( .A(x[81]), .B(n4795), .Z(n4797) );
  XOR U4879 ( .A(n4798), .B(n4799), .Z(n4795) );
  AND U4880 ( .A(n4800), .B(n4801), .Z(n4798) );
  XNOR U4881 ( .A(x[80]), .B(n4799), .Z(n4801) );
  XOR U4882 ( .A(n4802), .B(n4803), .Z(n4799) );
  AND U4883 ( .A(n4804), .B(n4805), .Z(n4802) );
  XNOR U4884 ( .A(x[79]), .B(n4803), .Z(n4805) );
  XOR U4885 ( .A(n4806), .B(n4807), .Z(n4803) );
  AND U4886 ( .A(n4808), .B(n4809), .Z(n4806) );
  XNOR U4887 ( .A(x[78]), .B(n4807), .Z(n4809) );
  XOR U4888 ( .A(n4810), .B(n4811), .Z(n4807) );
  AND U4889 ( .A(n4812), .B(n4813), .Z(n4810) );
  XNOR U4890 ( .A(x[77]), .B(n4811), .Z(n4813) );
  XOR U4891 ( .A(n4814), .B(n4815), .Z(n4811) );
  AND U4892 ( .A(n4816), .B(n4817), .Z(n4814) );
  XNOR U4893 ( .A(x[76]), .B(n4815), .Z(n4817) );
  XOR U4894 ( .A(n4818), .B(n4819), .Z(n4815) );
  AND U4895 ( .A(n4820), .B(n4821), .Z(n4818) );
  XNOR U4896 ( .A(x[75]), .B(n4819), .Z(n4821) );
  XOR U4897 ( .A(n4822), .B(n4823), .Z(n4819) );
  AND U4898 ( .A(n4824), .B(n4825), .Z(n4822) );
  XNOR U4899 ( .A(x[74]), .B(n4823), .Z(n4825) );
  XOR U4900 ( .A(n4826), .B(n4827), .Z(n4823) );
  AND U4901 ( .A(n4828), .B(n4829), .Z(n4826) );
  XNOR U4902 ( .A(x[73]), .B(n4827), .Z(n4829) );
  XOR U4903 ( .A(n4830), .B(n4831), .Z(n4827) );
  AND U4904 ( .A(n4832), .B(n4833), .Z(n4830) );
  XNOR U4905 ( .A(x[72]), .B(n4831), .Z(n4833) );
  XOR U4906 ( .A(n4834), .B(n4835), .Z(n4831) );
  AND U4907 ( .A(n4836), .B(n4837), .Z(n4834) );
  XNOR U4908 ( .A(x[71]), .B(n4835), .Z(n4837) );
  XOR U4909 ( .A(n4838), .B(n4839), .Z(n4835) );
  AND U4910 ( .A(n4840), .B(n4841), .Z(n4838) );
  XNOR U4911 ( .A(x[70]), .B(n4839), .Z(n4841) );
  XOR U4912 ( .A(n4842), .B(n4843), .Z(n4839) );
  AND U4913 ( .A(n4844), .B(n4845), .Z(n4842) );
  XNOR U4914 ( .A(x[69]), .B(n4843), .Z(n4845) );
  XOR U4915 ( .A(n4846), .B(n4847), .Z(n4843) );
  AND U4916 ( .A(n4848), .B(n4849), .Z(n4846) );
  XNOR U4917 ( .A(x[68]), .B(n4847), .Z(n4849) );
  XOR U4918 ( .A(n4850), .B(n4851), .Z(n4847) );
  AND U4919 ( .A(n4852), .B(n4853), .Z(n4850) );
  XNOR U4920 ( .A(x[67]), .B(n4851), .Z(n4853) );
  XOR U4921 ( .A(n4854), .B(n4855), .Z(n4851) );
  AND U4922 ( .A(n4856), .B(n4857), .Z(n4854) );
  XNOR U4923 ( .A(x[66]), .B(n4855), .Z(n4857) );
  XOR U4924 ( .A(n4858), .B(n4859), .Z(n4855) );
  AND U4925 ( .A(n4860), .B(n4861), .Z(n4858) );
  XNOR U4926 ( .A(x[65]), .B(n4859), .Z(n4861) );
  XOR U4927 ( .A(n4862), .B(n4863), .Z(n4859) );
  AND U4928 ( .A(n4864), .B(n4865), .Z(n4862) );
  XNOR U4929 ( .A(x[64]), .B(n4863), .Z(n4865) );
  XOR U4930 ( .A(n4866), .B(n4867), .Z(n4863) );
  AND U4931 ( .A(n4868), .B(n4869), .Z(n4866) );
  XNOR U4932 ( .A(x[63]), .B(n4867), .Z(n4869) );
  XOR U4933 ( .A(n4870), .B(n4871), .Z(n4867) );
  AND U4934 ( .A(n4872), .B(n4873), .Z(n4870) );
  XNOR U4935 ( .A(x[62]), .B(n4871), .Z(n4873) );
  XOR U4936 ( .A(n4874), .B(n4875), .Z(n4871) );
  AND U4937 ( .A(n4876), .B(n4877), .Z(n4874) );
  XNOR U4938 ( .A(x[61]), .B(n4875), .Z(n4877) );
  XOR U4939 ( .A(n4878), .B(n4879), .Z(n4875) );
  AND U4940 ( .A(n4880), .B(n4881), .Z(n4878) );
  XNOR U4941 ( .A(x[60]), .B(n4879), .Z(n4881) );
  XOR U4942 ( .A(n4882), .B(n4883), .Z(n4879) );
  AND U4943 ( .A(n4884), .B(n4885), .Z(n4882) );
  XNOR U4944 ( .A(x[59]), .B(n4883), .Z(n4885) );
  XOR U4945 ( .A(n4886), .B(n4887), .Z(n4883) );
  AND U4946 ( .A(n4888), .B(n4889), .Z(n4886) );
  XNOR U4947 ( .A(x[58]), .B(n4887), .Z(n4889) );
  XOR U4948 ( .A(n4890), .B(n4891), .Z(n4887) );
  AND U4949 ( .A(n4892), .B(n4893), .Z(n4890) );
  XNOR U4950 ( .A(x[57]), .B(n4891), .Z(n4893) );
  XOR U4951 ( .A(n4894), .B(n4895), .Z(n4891) );
  AND U4952 ( .A(n4896), .B(n4897), .Z(n4894) );
  XNOR U4953 ( .A(x[56]), .B(n4895), .Z(n4897) );
  XOR U4954 ( .A(n4898), .B(n4899), .Z(n4895) );
  AND U4955 ( .A(n4900), .B(n4901), .Z(n4898) );
  XNOR U4956 ( .A(x[55]), .B(n4899), .Z(n4901) );
  XOR U4957 ( .A(n4902), .B(n4903), .Z(n4899) );
  AND U4958 ( .A(n4904), .B(n4905), .Z(n4902) );
  XNOR U4959 ( .A(x[54]), .B(n4903), .Z(n4905) );
  XOR U4960 ( .A(n4906), .B(n4907), .Z(n4903) );
  AND U4961 ( .A(n4908), .B(n4909), .Z(n4906) );
  XNOR U4962 ( .A(x[53]), .B(n4907), .Z(n4909) );
  XOR U4963 ( .A(n4910), .B(n4911), .Z(n4907) );
  AND U4964 ( .A(n4912), .B(n4913), .Z(n4910) );
  XNOR U4965 ( .A(x[52]), .B(n4911), .Z(n4913) );
  XOR U4966 ( .A(n4914), .B(n4915), .Z(n4911) );
  AND U4967 ( .A(n4916), .B(n4917), .Z(n4914) );
  XNOR U4968 ( .A(x[51]), .B(n4915), .Z(n4917) );
  XOR U4969 ( .A(n4918), .B(n4919), .Z(n4915) );
  AND U4970 ( .A(n4920), .B(n4921), .Z(n4918) );
  XNOR U4971 ( .A(x[50]), .B(n4919), .Z(n4921) );
  XOR U4972 ( .A(n4922), .B(n4923), .Z(n4919) );
  AND U4973 ( .A(n4924), .B(n4925), .Z(n4922) );
  XNOR U4974 ( .A(x[49]), .B(n4923), .Z(n4925) );
  XOR U4975 ( .A(n4926), .B(n4927), .Z(n4923) );
  AND U4976 ( .A(n4928), .B(n4929), .Z(n4926) );
  XNOR U4977 ( .A(x[48]), .B(n4927), .Z(n4929) );
  XOR U4978 ( .A(n4930), .B(n4931), .Z(n4927) );
  AND U4979 ( .A(n4932), .B(n4933), .Z(n4930) );
  XNOR U4980 ( .A(x[47]), .B(n4931), .Z(n4933) );
  XOR U4981 ( .A(n4934), .B(n4935), .Z(n4931) );
  AND U4982 ( .A(n4936), .B(n4937), .Z(n4934) );
  XNOR U4983 ( .A(x[46]), .B(n4935), .Z(n4937) );
  XOR U4984 ( .A(n4938), .B(n4939), .Z(n4935) );
  AND U4985 ( .A(n4940), .B(n4941), .Z(n4938) );
  XNOR U4986 ( .A(x[45]), .B(n4939), .Z(n4941) );
  XOR U4987 ( .A(n4942), .B(n4943), .Z(n4939) );
  AND U4988 ( .A(n4944), .B(n4945), .Z(n4942) );
  XNOR U4989 ( .A(x[44]), .B(n4943), .Z(n4945) );
  XOR U4990 ( .A(n4946), .B(n4947), .Z(n4943) );
  AND U4991 ( .A(n4948), .B(n4949), .Z(n4946) );
  XNOR U4992 ( .A(x[43]), .B(n4947), .Z(n4949) );
  XOR U4993 ( .A(n4950), .B(n4951), .Z(n4947) );
  AND U4994 ( .A(n4952), .B(n4953), .Z(n4950) );
  XNOR U4995 ( .A(x[42]), .B(n4951), .Z(n4953) );
  XOR U4996 ( .A(n4954), .B(n4955), .Z(n4951) );
  AND U4997 ( .A(n4956), .B(n4957), .Z(n4954) );
  XNOR U4998 ( .A(x[41]), .B(n4955), .Z(n4957) );
  XOR U4999 ( .A(n4958), .B(n4959), .Z(n4955) );
  AND U5000 ( .A(n4960), .B(n4961), .Z(n4958) );
  XNOR U5001 ( .A(x[40]), .B(n4959), .Z(n4961) );
  XOR U5002 ( .A(n4962), .B(n4963), .Z(n4959) );
  AND U5003 ( .A(n4964), .B(n4965), .Z(n4962) );
  XNOR U5004 ( .A(x[39]), .B(n4963), .Z(n4965) );
  XOR U5005 ( .A(n4966), .B(n4967), .Z(n4963) );
  AND U5006 ( .A(n4968), .B(n4969), .Z(n4966) );
  XNOR U5007 ( .A(x[38]), .B(n4967), .Z(n4969) );
  XOR U5008 ( .A(n4970), .B(n4971), .Z(n4967) );
  AND U5009 ( .A(n4972), .B(n4973), .Z(n4970) );
  XNOR U5010 ( .A(x[37]), .B(n4971), .Z(n4973) );
  XOR U5011 ( .A(n4974), .B(n4975), .Z(n4971) );
  AND U5012 ( .A(n4976), .B(n4977), .Z(n4974) );
  XNOR U5013 ( .A(x[36]), .B(n4975), .Z(n4977) );
  XOR U5014 ( .A(n4978), .B(n4979), .Z(n4975) );
  AND U5015 ( .A(n4980), .B(n4981), .Z(n4978) );
  XNOR U5016 ( .A(x[35]), .B(n4979), .Z(n4981) );
  XOR U5017 ( .A(n4982), .B(n4983), .Z(n4979) );
  AND U5018 ( .A(n4984), .B(n4985), .Z(n4982) );
  XNOR U5019 ( .A(x[34]), .B(n4983), .Z(n4985) );
  XOR U5020 ( .A(n4986), .B(n4987), .Z(n4983) );
  AND U5021 ( .A(n4988), .B(n4989), .Z(n4986) );
  XNOR U5022 ( .A(x[33]), .B(n4987), .Z(n4989) );
  XOR U5023 ( .A(n4990), .B(n4991), .Z(n4987) );
  AND U5024 ( .A(n4992), .B(n4993), .Z(n4990) );
  XNOR U5025 ( .A(x[32]), .B(n4991), .Z(n4993) );
  XOR U5026 ( .A(n4994), .B(n4995), .Z(n4991) );
  AND U5027 ( .A(n4996), .B(n4997), .Z(n4994) );
  XNOR U5028 ( .A(x[31]), .B(n4995), .Z(n4997) );
  XOR U5029 ( .A(n4998), .B(n4999), .Z(n4995) );
  AND U5030 ( .A(n5000), .B(n5001), .Z(n4998) );
  XNOR U5031 ( .A(x[30]), .B(n4999), .Z(n5001) );
  XOR U5032 ( .A(n5002), .B(n5003), .Z(n4999) );
  AND U5033 ( .A(n5004), .B(n5005), .Z(n5002) );
  XNOR U5034 ( .A(x[29]), .B(n5003), .Z(n5005) );
  XOR U5035 ( .A(n5006), .B(n5007), .Z(n5003) );
  AND U5036 ( .A(n5008), .B(n5009), .Z(n5006) );
  XNOR U5037 ( .A(x[28]), .B(n5007), .Z(n5009) );
  XOR U5038 ( .A(n5010), .B(n5011), .Z(n5007) );
  AND U5039 ( .A(n5012), .B(n5013), .Z(n5010) );
  XNOR U5040 ( .A(x[27]), .B(n5011), .Z(n5013) );
  XOR U5041 ( .A(n5014), .B(n5015), .Z(n5011) );
  AND U5042 ( .A(n5016), .B(n5017), .Z(n5014) );
  XNOR U5043 ( .A(x[26]), .B(n5015), .Z(n5017) );
  XOR U5044 ( .A(n5018), .B(n5019), .Z(n5015) );
  AND U5045 ( .A(n5020), .B(n5021), .Z(n5018) );
  XNOR U5046 ( .A(x[25]), .B(n5019), .Z(n5021) );
  XOR U5047 ( .A(n5022), .B(n5023), .Z(n5019) );
  AND U5048 ( .A(n5024), .B(n5025), .Z(n5022) );
  XNOR U5049 ( .A(x[24]), .B(n5023), .Z(n5025) );
  XOR U5050 ( .A(n5026), .B(n5027), .Z(n5023) );
  AND U5051 ( .A(n5028), .B(n5029), .Z(n5026) );
  XNOR U5052 ( .A(x[23]), .B(n5027), .Z(n5029) );
  XOR U5053 ( .A(n5030), .B(n5031), .Z(n5027) );
  AND U5054 ( .A(n5032), .B(n5033), .Z(n5030) );
  XNOR U5055 ( .A(x[22]), .B(n5031), .Z(n5033) );
  XOR U5056 ( .A(n5034), .B(n5035), .Z(n5031) );
  AND U5057 ( .A(n5036), .B(n5037), .Z(n5034) );
  XNOR U5058 ( .A(x[21]), .B(n5035), .Z(n5037) );
  XOR U5059 ( .A(n5038), .B(n5039), .Z(n5035) );
  AND U5060 ( .A(n5040), .B(n5041), .Z(n5038) );
  XNOR U5061 ( .A(x[20]), .B(n5039), .Z(n5041) );
  XOR U5062 ( .A(n5042), .B(n5043), .Z(n5039) );
  AND U5063 ( .A(n5044), .B(n5045), .Z(n5042) );
  XNOR U5064 ( .A(x[19]), .B(n5043), .Z(n5045) );
  XOR U5065 ( .A(n5046), .B(n5047), .Z(n5043) );
  AND U5066 ( .A(n5048), .B(n5049), .Z(n5046) );
  XNOR U5067 ( .A(x[18]), .B(n5047), .Z(n5049) );
  XOR U5068 ( .A(n5050), .B(n5051), .Z(n5047) );
  AND U5069 ( .A(n5052), .B(n5053), .Z(n5050) );
  XNOR U5070 ( .A(x[17]), .B(n5051), .Z(n5053) );
  XOR U5071 ( .A(n5054), .B(n5055), .Z(n5051) );
  AND U5072 ( .A(n5056), .B(n5057), .Z(n5054) );
  XNOR U5073 ( .A(x[16]), .B(n5055), .Z(n5057) );
  XOR U5074 ( .A(n5058), .B(n5059), .Z(n5055) );
  AND U5075 ( .A(n5060), .B(n5061), .Z(n5058) );
  XNOR U5076 ( .A(x[15]), .B(n5059), .Z(n5061) );
  XOR U5077 ( .A(n5062), .B(n5063), .Z(n5059) );
  AND U5078 ( .A(n5064), .B(n5065), .Z(n5062) );
  XNOR U5079 ( .A(x[14]), .B(n5063), .Z(n5065) );
  XOR U5080 ( .A(n5066), .B(n5067), .Z(n5063) );
  AND U5081 ( .A(n5068), .B(n5069), .Z(n5066) );
  XNOR U5082 ( .A(x[13]), .B(n5067), .Z(n5069) );
  XOR U5083 ( .A(n5070), .B(n5071), .Z(n5067) );
  AND U5084 ( .A(n5072), .B(n5073), .Z(n5070) );
  XNOR U5085 ( .A(x[12]), .B(n5071), .Z(n5073) );
  XOR U5086 ( .A(n5074), .B(n5075), .Z(n5071) );
  AND U5087 ( .A(n5076), .B(n5077), .Z(n5074) );
  XNOR U5088 ( .A(x[11]), .B(n5075), .Z(n5077) );
  XOR U5089 ( .A(n5078), .B(n5079), .Z(n5075) );
  AND U5090 ( .A(n5080), .B(n5081), .Z(n5078) );
  XNOR U5091 ( .A(x[10]), .B(n5079), .Z(n5081) );
  XOR U5092 ( .A(n5082), .B(n5083), .Z(n5079) );
  AND U5093 ( .A(n5084), .B(n5085), .Z(n5082) );
  XNOR U5094 ( .A(x[9]), .B(n5083), .Z(n5085) );
  XOR U5095 ( .A(n5086), .B(n5087), .Z(n5083) );
  AND U5096 ( .A(n5088), .B(n5089), .Z(n5086) );
  XNOR U5097 ( .A(x[8]), .B(n5087), .Z(n5089) );
  XOR U5098 ( .A(n5090), .B(n5091), .Z(n5087) );
  AND U5099 ( .A(n5092), .B(n5093), .Z(n5090) );
  XNOR U5100 ( .A(x[7]), .B(n5091), .Z(n5093) );
  XOR U5101 ( .A(n5094), .B(n5095), .Z(n5091) );
  AND U5102 ( .A(n5096), .B(n5097), .Z(n5094) );
  XNOR U5103 ( .A(x[6]), .B(n5095), .Z(n5097) );
  XOR U5104 ( .A(n5098), .B(n5099), .Z(n5095) );
  AND U5105 ( .A(n5100), .B(n5101), .Z(n5098) );
  XNOR U5106 ( .A(x[5]), .B(n5099), .Z(n5101) );
  XOR U5107 ( .A(n5102), .B(n5103), .Z(n5099) );
  AND U5108 ( .A(n5104), .B(n5105), .Z(n5102) );
  XNOR U5109 ( .A(x[4]), .B(n5103), .Z(n5105) );
  XOR U5110 ( .A(n5106), .B(n5107), .Z(n5103) );
  AND U5111 ( .A(n5108), .B(n5109), .Z(n5106) );
  XNOR U5112 ( .A(x[3]), .B(n5107), .Z(n5109) );
  XOR U5113 ( .A(n5110), .B(n5111), .Z(n5107) );
  AND U5114 ( .A(n5112), .B(n5113), .Z(n5110) );
  XNOR U5115 ( .A(x[2]), .B(n5111), .Z(n5113) );
  XOR U5116 ( .A(n5114), .B(n5115), .Z(n5111) );
  AND U5117 ( .A(n5116), .B(n5117), .Z(n5114) );
  XNOR U5118 ( .A(x[1]), .B(n5115), .Z(n5117) );
  XOR U5119 ( .A(y[1]), .B(n5115), .Z(n5116) );
  XOR U5120 ( .A(ci), .B(n5118), .Z(n5115) );
  NANDN U5121 ( .A(n5119), .B(n5120), .Z(n5118) );
  XOR U5122 ( .A(x[0]), .B(ci), .Z(n5120) );
  XOR U5123 ( .A(y[0]), .B(ci), .Z(n5119) );
endmodule

