
module hamming_N1600_CC8 ( clk, rst, x, y, o );
  input [199:0] x;
  input [199:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NANDN U203 ( .A(n732), .B(n733), .Z(n1) );
  NANDN U204 ( .A(n730), .B(n731), .Z(n2) );
  AND U205 ( .A(n1), .B(n2), .Z(n1033) );
  NAND U206 ( .A(n739), .B(n738), .Z(n3) );
  NANDN U207 ( .A(n740), .B(n741), .Z(n4) );
  NAND U208 ( .A(n3), .B(n4), .Z(n959) );
  NAND U209 ( .A(n639), .B(n638), .Z(n5) );
  NANDN U210 ( .A(n640), .B(n641), .Z(n6) );
  AND U211 ( .A(n5), .B(n6), .Z(n919) );
  NAND U212 ( .A(n377), .B(oglobal[0]), .Z(n7) );
  NANDN U213 ( .A(n378), .B(n379), .Z(n8) );
  NAND U214 ( .A(n7), .B(n8), .Z(n915) );
  NAND U215 ( .A(n936), .B(n935), .Z(n9) );
  XOR U216 ( .A(n936), .B(n935), .Z(n10) );
  NANDN U217 ( .A(n934), .B(n10), .Z(n11) );
  NAND U218 ( .A(n9), .B(n11), .Z(n1111) );
  XOR U219 ( .A(n946), .B(n944), .Z(n12) );
  NANDN U220 ( .A(n945), .B(n12), .Z(n13) );
  NAND U221 ( .A(n946), .B(n944), .Z(n14) );
  AND U222 ( .A(n13), .B(n14), .Z(n1133) );
  XOR U223 ( .A(n1043), .B(n1041), .Z(n15) );
  NANDN U224 ( .A(n1042), .B(n15), .Z(n16) );
  NAND U225 ( .A(n1043), .B(n1041), .Z(n17) );
  AND U226 ( .A(n16), .B(n17), .Z(n1140) );
  NAND U227 ( .A(n992), .B(n993), .Z(n18) );
  XOR U228 ( .A(n992), .B(n993), .Z(n19) );
  NANDN U229 ( .A(n991), .B(n19), .Z(n20) );
  NAND U230 ( .A(n18), .B(n20), .Z(n1136) );
  NAND U231 ( .A(n954), .B(n953), .Z(n21) );
  XOR U232 ( .A(n954), .B(n953), .Z(n22) );
  NANDN U233 ( .A(n952), .B(n22), .Z(n23) );
  NAND U234 ( .A(n21), .B(n23), .Z(n1113) );
  NAND U235 ( .A(n912), .B(n913), .Z(n24) );
  XOR U236 ( .A(n912), .B(n913), .Z(n25) );
  NANDN U237 ( .A(n911), .B(n25), .Z(n26) );
  NAND U238 ( .A(n24), .B(n26), .Z(n1118) );
  NAND U239 ( .A(n964), .B(n962), .Z(n27) );
  XOR U240 ( .A(n964), .B(n962), .Z(n28) );
  NANDN U241 ( .A(n963), .B(n28), .Z(n29) );
  NAND U242 ( .A(n27), .B(n29), .Z(n1145) );
  XOR U243 ( .A(n973), .B(n971), .Z(n30) );
  NANDN U244 ( .A(n972), .B(n30), .Z(n31) );
  NAND U245 ( .A(n973), .B(n971), .Z(n32) );
  AND U246 ( .A(n31), .B(n32), .Z(n1143) );
  NAND U247 ( .A(n649), .B(n647), .Z(n33) );
  XOR U248 ( .A(n649), .B(n647), .Z(n34) );
  NANDN U249 ( .A(n648), .B(n34), .Z(n35) );
  NAND U250 ( .A(n33), .B(n35), .Z(n978) );
  NAND U251 ( .A(n698), .B(n699), .Z(n36) );
  XOR U252 ( .A(n698), .B(n699), .Z(n37) );
  NANDN U253 ( .A(n697), .B(n37), .Z(n38) );
  NAND U254 ( .A(n36), .B(n38), .Z(n896) );
  NAND U255 ( .A(n843), .B(n844), .Z(n39) );
  XOR U256 ( .A(n843), .B(n844), .Z(n40) );
  NANDN U257 ( .A(n842), .B(n40), .Z(n41) );
  NAND U258 ( .A(n39), .B(n41), .Z(n1045) );
  NAND U259 ( .A(n1089), .B(n1088), .Z(n42) );
  XOR U260 ( .A(n1089), .B(n1088), .Z(n43) );
  NANDN U261 ( .A(n1090), .B(n43), .Z(n44) );
  NAND U262 ( .A(n42), .B(n44), .Z(n1160) );
  NAND U263 ( .A(n1195), .B(n1194), .Z(n45) );
  XOR U264 ( .A(n1195), .B(n1194), .Z(n46) );
  NANDN U265 ( .A(n1196), .B(n46), .Z(n47) );
  NAND U266 ( .A(n45), .B(n47), .Z(n1249) );
  NAND U267 ( .A(n1085), .B(n1087), .Z(n48) );
  XOR U268 ( .A(n1085), .B(n1087), .Z(n49) );
  NAND U269 ( .A(n49), .B(n1086), .Z(n50) );
  NAND U270 ( .A(n48), .B(n50), .Z(n1204) );
  NAND U271 ( .A(n1301), .B(n1303), .Z(n51) );
  XOR U272 ( .A(n1301), .B(n1303), .Z(n52) );
  NAND U273 ( .A(n52), .B(n1302), .Z(n53) );
  NAND U274 ( .A(n51), .B(n53), .Z(n1311) );
  XOR U275 ( .A(n767), .B(n768), .Z(n54) );
  NANDN U276 ( .A(n769), .B(n54), .Z(n55) );
  NAND U277 ( .A(n767), .B(n768), .Z(n56) );
  AND U278 ( .A(n55), .B(n56), .Z(n1079) );
  XNOR U279 ( .A(n1211), .B(n1210), .Z(n57) );
  XNOR U280 ( .A(n1212), .B(n57), .Z(n1209) );
  NAND U281 ( .A(n1306), .B(n1305), .Z(n58) );
  XOR U282 ( .A(n1306), .B(n1305), .Z(n59) );
  NANDN U283 ( .A(n1307), .B(n59), .Z(n60) );
  NAND U284 ( .A(n58), .B(n60), .Z(n1316) );
  NAND U285 ( .A(n391), .B(n390), .Z(n61) );
  NANDN U286 ( .A(n392), .B(n393), .Z(n62) );
  NAND U287 ( .A(n61), .B(n62), .Z(n993) );
  NANDN U288 ( .A(n864), .B(n865), .Z(n63) );
  NANDN U289 ( .A(n862), .B(n863), .Z(n64) );
  AND U290 ( .A(n63), .B(n64), .Z(n971) );
  NAND U291 ( .A(n716), .B(n715), .Z(n65) );
  NANDN U292 ( .A(n717), .B(n718), .Z(n66) );
  AND U293 ( .A(n65), .B(n66), .Z(n928) );
  NAND U294 ( .A(n933), .B(n931), .Z(n67) );
  XOR U295 ( .A(n933), .B(n931), .Z(n68) );
  NANDN U296 ( .A(n932), .B(n68), .Z(n69) );
  NAND U297 ( .A(n67), .B(n69), .Z(n1112) );
  XOR U298 ( .A(n940), .B(n938), .Z(n70) );
  NANDN U299 ( .A(n939), .B(n70), .Z(n71) );
  NAND U300 ( .A(n940), .B(n938), .Z(n72) );
  AND U301 ( .A(n71), .B(n72), .Z(n1132) );
  XOR U302 ( .A(n970), .B(n968), .Z(n73) );
  NANDN U303 ( .A(n969), .B(n73), .Z(n74) );
  NAND U304 ( .A(n970), .B(n968), .Z(n75) );
  AND U305 ( .A(n74), .B(n75), .Z(n1144) );
  NAND U306 ( .A(n1065), .B(n1067), .Z(n76) );
  XOR U307 ( .A(n1065), .B(n1067), .Z(n77) );
  NAND U308 ( .A(n77), .B(n1066), .Z(n78) );
  NAND U309 ( .A(n76), .B(n78), .Z(n1194) );
  NAND U310 ( .A(n1139), .B(n1138), .Z(n79) );
  XOR U311 ( .A(n1139), .B(n1138), .Z(n80) );
  NANDN U312 ( .A(n1140), .B(n80), .Z(n81) );
  NAND U313 ( .A(n79), .B(n81), .Z(n1255) );
  NAND U314 ( .A(n1118), .B(n1120), .Z(n82) );
  XOR U315 ( .A(n1118), .B(n1120), .Z(n83) );
  NAND U316 ( .A(n83), .B(n1119), .Z(n84) );
  NAND U317 ( .A(n82), .B(n84), .Z(n1253) );
  OR U318 ( .A(n1147), .B(n1148), .Z(n85) );
  OR U319 ( .A(n1146), .B(n1145), .Z(n86) );
  NAND U320 ( .A(n85), .B(n86), .Z(n1245) );
  XOR U321 ( .A(n850), .B(n848), .Z(n87) );
  NANDN U322 ( .A(n849), .B(n87), .Z(n88) );
  NAND U323 ( .A(n850), .B(n848), .Z(n89) );
  AND U324 ( .A(n88), .B(n89), .Z(n1046) );
  XOR U325 ( .A(n494), .B(n492), .Z(n90) );
  NANDN U326 ( .A(n493), .B(n90), .Z(n91) );
  NAND U327 ( .A(n494), .B(n492), .Z(n92) );
  AND U328 ( .A(n91), .B(n92), .Z(n998) );
  NAND U329 ( .A(n1000), .B(n999), .Z(n93) );
  XOR U330 ( .A(n1000), .B(n999), .Z(n94) );
  NANDN U331 ( .A(n1001), .B(n94), .Z(n95) );
  NAND U332 ( .A(n93), .B(n95), .Z(n1165) );
  NAND U333 ( .A(n1191), .B(n1193), .Z(n96) );
  XOR U334 ( .A(n1191), .B(n1193), .Z(n97) );
  NAND U335 ( .A(n97), .B(n1192), .Z(n98) );
  NAND U336 ( .A(n96), .B(n98), .Z(n1250) );
  NAND U337 ( .A(n1004), .B(n1005), .Z(n99) );
  XOR U338 ( .A(n1004), .B(n1005), .Z(n100) );
  NANDN U339 ( .A(n1003), .B(n100), .Z(n101) );
  NAND U340 ( .A(n99), .B(n101), .Z(n1176) );
  NANDN U341 ( .A(n1170), .B(n1173), .Z(n102) );
  OR U342 ( .A(n1173), .B(n1171), .Z(n103) );
  NAND U343 ( .A(n1172), .B(n103), .Z(n104) );
  NAND U344 ( .A(n102), .B(n104), .Z(n1226) );
  XOR U345 ( .A(n1084), .B(n1082), .Z(n105) );
  NANDN U346 ( .A(n1083), .B(n105), .Z(n106) );
  NAND U347 ( .A(n1084), .B(n1082), .Z(n107) );
  AND U348 ( .A(n106), .B(n107), .Z(n1202) );
  NAND U349 ( .A(n1207), .B(n1209), .Z(n108) );
  XOR U350 ( .A(n1207), .B(n1209), .Z(n109) );
  NAND U351 ( .A(n109), .B(n1208), .Z(n110) );
  NAND U352 ( .A(n108), .B(n110), .Z(n1278) );
  NAND U353 ( .A(n1312), .B(n1313), .Z(n111) );
  XOR U354 ( .A(n1312), .B(n1313), .Z(n112) );
  NAND U355 ( .A(n112), .B(n1311), .Z(n113) );
  NAND U356 ( .A(n111), .B(n113), .Z(n1325) );
  NAND U357 ( .A(n1318), .B(n1319), .Z(n114) );
  XOR U358 ( .A(n1318), .B(n1319), .Z(n115) );
  NANDN U359 ( .A(n1317), .B(n115), .Z(n116) );
  NAND U360 ( .A(n114), .B(n116), .Z(n1321) );
  NAND U361 ( .A(n655), .B(n654), .Z(n117) );
  NANDN U362 ( .A(n656), .B(n657), .Z(n118) );
  NAND U363 ( .A(n117), .B(n118), .Z(n934) );
  NAND U364 ( .A(n399), .B(n398), .Z(n119) );
  NANDN U365 ( .A(n400), .B(n401), .Z(n120) );
  AND U366 ( .A(n119), .B(n120), .Z(n991) );
  NAND U367 ( .A(n883), .B(n882), .Z(n121) );
  NANDN U368 ( .A(n884), .B(n885), .Z(n122) );
  AND U369 ( .A(n121), .B(n122), .Z(n985) );
  NAND U370 ( .A(n643), .B(n642), .Z(n123) );
  NANDN U371 ( .A(n644), .B(n645), .Z(n124) );
  NAND U372 ( .A(n123), .B(n124), .Z(n918) );
  NAND U373 ( .A(n712), .B(n711), .Z(n125) );
  NANDN U374 ( .A(n713), .B(n714), .Z(n126) );
  NAND U375 ( .A(n125), .B(n126), .Z(n925) );
  NAND U376 ( .A(n586), .B(n585), .Z(n127) );
  NANDN U377 ( .A(n587), .B(n588), .Z(n128) );
  AND U378 ( .A(n127), .B(n128), .Z(n962) );
  XOR U379 ( .A(n990), .B(n988), .Z(n129) );
  NANDN U380 ( .A(n989), .B(n129), .Z(n130) );
  NAND U381 ( .A(n990), .B(n988), .Z(n131) );
  AND U382 ( .A(n130), .B(n131), .Z(n1137) );
  NAND U383 ( .A(n960), .B(n961), .Z(n132) );
  XOR U384 ( .A(n960), .B(n961), .Z(n133) );
  NANDN U385 ( .A(n959), .B(n133), .Z(n134) );
  NAND U386 ( .A(n132), .B(n134), .Z(n1146) );
  NAND U387 ( .A(n869), .B(n867), .Z(n135) );
  XOR U388 ( .A(n869), .B(n867), .Z(n136) );
  NANDN U389 ( .A(n868), .B(n136), .Z(n137) );
  NAND U390 ( .A(n135), .B(n137), .Z(n1026) );
  XOR U391 ( .A(n834), .B(n832), .Z(n138) );
  NANDN U392 ( .A(n833), .B(n138), .Z(n139) );
  NAND U393 ( .A(n834), .B(n832), .Z(n140) );
  AND U394 ( .A(n139), .B(n140), .Z(n1066) );
  XOR U395 ( .A(n841), .B(n839), .Z(n141) );
  NANDN U396 ( .A(n840), .B(n141), .Z(n142) );
  NAND U397 ( .A(n841), .B(n839), .Z(n143) );
  AND U398 ( .A(n142), .B(n143), .Z(n979) );
  NAND U399 ( .A(n388), .B(n389), .Z(n144) );
  XOR U400 ( .A(n388), .B(n389), .Z(n145) );
  NANDN U401 ( .A(n387), .B(n145), .Z(n146) );
  NAND U402 ( .A(n144), .B(n146), .Z(n1019) );
  NAND U403 ( .A(n1073), .B(n1074), .Z(n147) );
  XOR U404 ( .A(n1073), .B(n1074), .Z(n148) );
  NANDN U405 ( .A(n1072), .B(n148), .Z(n149) );
  NAND U406 ( .A(n147), .B(n149), .Z(n1122) );
  NAND U407 ( .A(n1132), .B(n1134), .Z(n150) );
  XOR U408 ( .A(n1132), .B(n1134), .Z(n151) );
  NAND U409 ( .A(n151), .B(n1133), .Z(n152) );
  NAND U410 ( .A(n150), .B(n152), .Z(n1256) );
  NAND U411 ( .A(n1142), .B(n1144), .Z(n153) );
  XOR U412 ( .A(n1142), .B(n1144), .Z(n154) );
  NAND U413 ( .A(n154), .B(n1143), .Z(n155) );
  NAND U414 ( .A(n153), .B(n155), .Z(n1246) );
  NAND U415 ( .A(n490), .B(n491), .Z(n156) );
  XOR U416 ( .A(n490), .B(n491), .Z(n157) );
  NANDN U417 ( .A(n489), .B(n157), .Z(n158) );
  NAND U418 ( .A(n156), .B(n158), .Z(n997) );
  NAND U419 ( .A(n1129), .B(n1130), .Z(n159) );
  XOR U420 ( .A(n1129), .B(n1130), .Z(n160) );
  NANDN U421 ( .A(n1128), .B(n160), .Z(n161) );
  NAND U422 ( .A(n159), .B(n161), .Z(n1223) );
  XOR U423 ( .A(n1254), .B(n1252), .Z(n162) );
  NANDN U424 ( .A(n1253), .B(n162), .Z(n163) );
  NAND U425 ( .A(n1254), .B(n1252), .Z(n164) );
  AND U426 ( .A(n163), .B(n164), .Z(n1302) );
  NAND U427 ( .A(n1250), .B(n1249), .Z(n165) );
  XOR U428 ( .A(n1250), .B(n1249), .Z(n166) );
  NANDN U429 ( .A(n1251), .B(n166), .Z(n167) );
  NAND U430 ( .A(n165), .B(n167), .Z(n1300) );
  NAND U431 ( .A(n815), .B(n814), .Z(n168) );
  XOR U432 ( .A(n815), .B(n814), .Z(n169) );
  NANDN U433 ( .A(n813), .B(n169), .Z(n170) );
  NAND U434 ( .A(n168), .B(n170), .Z(n1000) );
  NAND U435 ( .A(n1160), .B(n1162), .Z(n171) );
  XOR U436 ( .A(n1160), .B(n1162), .Z(n172) );
  NAND U437 ( .A(n172), .B(n1161), .Z(n173) );
  NAND U438 ( .A(n171), .B(n173), .Z(n1225) );
  NAND U439 ( .A(n1108), .B(n1107), .Z(n174) );
  XOR U440 ( .A(n1108), .B(n1107), .Z(n175) );
  NANDN U441 ( .A(n1109), .B(n175), .Z(n176) );
  NAND U442 ( .A(n174), .B(n176), .Z(n1240) );
  XOR U443 ( .A(n822), .B(n820), .Z(n177) );
  NANDN U444 ( .A(n821), .B(n177), .Z(n178) );
  NAND U445 ( .A(n822), .B(n820), .Z(n179) );
  AND U446 ( .A(n178), .B(n179), .Z(n1086) );
  NAND U447 ( .A(n1078), .B(n1080), .Z(n180) );
  XOR U448 ( .A(n1078), .B(n1080), .Z(n181) );
  NAND U449 ( .A(n181), .B(n1079), .Z(n182) );
  NAND U450 ( .A(n180), .B(n182), .Z(n1207) );
  XOR U451 ( .A(n1210), .B(n1211), .Z(n183) );
  NANDN U452 ( .A(n1212), .B(n183), .Z(n184) );
  NAND U453 ( .A(n1210), .B(n1211), .Z(n185) );
  AND U454 ( .A(n184), .B(n185), .Z(n1277) );
  XNOR U455 ( .A(n768), .B(n767), .Z(n186) );
  XNOR U456 ( .A(n769), .B(n186), .Z(n892) );
  XOR U457 ( .A(n1316), .B(n1314), .Z(n187) );
  NANDN U458 ( .A(n1315), .B(n187), .Z(n188) );
  NAND U459 ( .A(n1316), .B(n1314), .Z(n189) );
  AND U460 ( .A(n188), .B(n189), .Z(n1322) );
  NANDN U461 ( .A(n394), .B(n395), .Z(n190) );
  NANDN U462 ( .A(n396), .B(n397), .Z(n191) );
  NAND U463 ( .A(n190), .B(n191), .Z(n992) );
  NANDN U464 ( .A(n854), .B(n855), .Z(n192) );
  NANDN U465 ( .A(n852), .B(n853), .Z(n193) );
  AND U466 ( .A(n192), .B(n193), .Z(n973) );
  NANDN U467 ( .A(n577), .B(n578), .Z(n194) );
  NANDN U468 ( .A(n579), .B(n580), .Z(n195) );
  NAND U469 ( .A(n194), .B(n195), .Z(n963) );
  NAND U470 ( .A(n573), .B(n572), .Z(n196) );
  NANDN U471 ( .A(n574), .B(n575), .Z(n197) );
  AND U472 ( .A(n196), .B(n197), .Z(n956) );
  XOR U473 ( .A(oglobal[1]), .B(n1040), .Z(n198) );
  NANDN U474 ( .A(n1039), .B(n198), .Z(n199) );
  NAND U475 ( .A(oglobal[1]), .B(n1040), .Z(n200) );
  AND U476 ( .A(n199), .B(n200), .Z(n1139) );
  XOR U477 ( .A(n987), .B(n985), .Z(n201) );
  NANDN U478 ( .A(n986), .B(n201), .Z(n202) );
  NAND U479 ( .A(n987), .B(n985), .Z(n203) );
  AND U480 ( .A(n202), .B(n203), .Z(n1135) );
  NAND U481 ( .A(n950), .B(n951), .Z(n204) );
  XOR U482 ( .A(n950), .B(n951), .Z(n205) );
  NANDN U483 ( .A(n949), .B(n205), .Z(n206) );
  NAND U484 ( .A(n204), .B(n206), .Z(n1114) );
  NAND U485 ( .A(n823), .B(n825), .Z(n207) );
  XOR U486 ( .A(n823), .B(n825), .Z(n208) );
  NAND U487 ( .A(n208), .B(n824), .Z(n209) );
  NAND U488 ( .A(n207), .B(n209), .Z(n1065) );
  NAND U489 ( .A(n838), .B(n836), .Z(n210) );
  XOR U490 ( .A(n838), .B(n836), .Z(n211) );
  NANDN U491 ( .A(n837), .B(n211), .Z(n212) );
  NAND U492 ( .A(n210), .B(n212), .Z(n980) );
  NAND U493 ( .A(n652), .B(n650), .Z(n213) );
  XOR U494 ( .A(n652), .B(n650), .Z(n214) );
  NANDN U495 ( .A(n651), .B(n214), .Z(n215) );
  NAND U496 ( .A(n213), .B(n215), .Z(n977) );
  NAND U497 ( .A(n673), .B(n671), .Z(n216) );
  XOR U498 ( .A(n673), .B(n671), .Z(n217) );
  NANDN U499 ( .A(n672), .B(n217), .Z(n218) );
  NAND U500 ( .A(n216), .B(n218), .Z(n1055) );
  XOR U501 ( .A(n484), .B(n485), .Z(n219) );
  NANDN U502 ( .A(n486), .B(n219), .Z(n220) );
  NAND U503 ( .A(n484), .B(n485), .Z(n221) );
  AND U504 ( .A(n220), .B(n221), .Z(n1069) );
  NAND U505 ( .A(n729), .B(n727), .Z(n222) );
  XOR U506 ( .A(n729), .B(n727), .Z(n223) );
  NANDN U507 ( .A(n728), .B(n223), .Z(n224) );
  NAND U508 ( .A(n222), .B(n224), .Z(n905) );
  NAND U509 ( .A(n592), .B(n590), .Z(n225) );
  XOR U510 ( .A(n592), .B(n590), .Z(n226) );
  NANDN U511 ( .A(n591), .B(n226), .Z(n227) );
  NAND U512 ( .A(n225), .B(n227), .Z(n897) );
  NAND U513 ( .A(n702), .B(n700), .Z(n228) );
  XOR U514 ( .A(n702), .B(n700), .Z(n229) );
  NANDN U515 ( .A(n701), .B(n229), .Z(n230) );
  NAND U516 ( .A(n228), .B(n230), .Z(n895) );
  NAND U517 ( .A(n1060), .B(n1061), .Z(n231) );
  XOR U518 ( .A(n1060), .B(n1061), .Z(n232) );
  NANDN U519 ( .A(n1059), .B(n232), .Z(n233) );
  NAND U520 ( .A(n231), .B(n233), .Z(n1196) );
  NAND U521 ( .A(n846), .B(n847), .Z(n234) );
  XOR U522 ( .A(n846), .B(n847), .Z(n235) );
  NANDN U523 ( .A(n845), .B(n235), .Z(n236) );
  NAND U524 ( .A(n234), .B(n236), .Z(n1048) );
  NAND U525 ( .A(n997), .B(n998), .Z(n237) );
  XOR U526 ( .A(n997), .B(n998), .Z(n238) );
  NANDN U527 ( .A(n996), .B(n238), .Z(n239) );
  NAND U528 ( .A(n237), .B(n239), .Z(n1167) );
  NANDN U529 ( .A(n1187), .B(n1190), .Z(n240) );
  OR U530 ( .A(n1190), .B(n1188), .Z(n241) );
  NAND U531 ( .A(n1189), .B(n241), .Z(n242) );
  NAND U532 ( .A(n240), .B(n242), .Z(n1251) );
  NAND U533 ( .A(n1156), .B(n1157), .Z(n243) );
  XOR U534 ( .A(n1156), .B(n1157), .Z(n244) );
  NANDN U535 ( .A(n1155), .B(n244), .Z(n245) );
  NAND U536 ( .A(n243), .B(n245), .Z(n1233) );
  OR U537 ( .A(n1246), .B(n1245), .Z(n246) );
  NANDN U538 ( .A(n1248), .B(n1247), .Z(n247) );
  NAND U539 ( .A(n246), .B(n247), .Z(n1299) );
  XOR U540 ( .A(n443), .B(n442), .Z(n248) );
  XNOR U541 ( .A(n444), .B(n248), .Z(n757) );
  NAND U542 ( .A(n1222), .B(n1224), .Z(n249) );
  XOR U543 ( .A(n1222), .B(n1224), .Z(n250) );
  NAND U544 ( .A(n250), .B(n1223), .Z(n251) );
  NAND U545 ( .A(n249), .B(n251), .Z(n1296) );
  NAND U546 ( .A(n1273), .B(n1274), .Z(n252) );
  XOR U547 ( .A(n1273), .B(n1274), .Z(n253) );
  NANDN U548 ( .A(n1272), .B(n253), .Z(n254) );
  NAND U549 ( .A(n252), .B(n254), .Z(n1290) );
  NAND U550 ( .A(n1104), .B(n1105), .Z(n255) );
  XOR U551 ( .A(n1104), .B(n1105), .Z(n256) );
  NANDN U552 ( .A(n1103), .B(n256), .Z(n257) );
  NAND U553 ( .A(n255), .B(n257), .Z(n1215) );
  NAND U554 ( .A(n1276), .B(n1278), .Z(n258) );
  XOR U555 ( .A(n1276), .B(n1278), .Z(n259) );
  NAND U556 ( .A(n259), .B(n1277), .Z(n260) );
  NAND U557 ( .A(n258), .B(n260), .Z(n1287) );
  NAND U558 ( .A(n1321), .B(n1323), .Z(n261) );
  XOR U559 ( .A(n1321), .B(n1323), .Z(n262) );
  NAND U560 ( .A(n262), .B(n1322), .Z(n263) );
  NAND U561 ( .A(n261), .B(n263), .Z(n1331) );
  NANDN U562 ( .A(n734), .B(n735), .Z(n264) );
  NANDN U563 ( .A(n736), .B(n737), .Z(n265) );
  NAND U564 ( .A(n264), .B(n265), .Z(n1034) );
  NAND U565 ( .A(n750), .B(n749), .Z(n266) );
  NANDN U566 ( .A(n751), .B(n752), .Z(n267) );
  AND U567 ( .A(n266), .B(n267), .Z(n960) );
  NAND U568 ( .A(n582), .B(n581), .Z(n268) );
  NANDN U569 ( .A(n583), .B(n584), .Z(n269) );
  AND U570 ( .A(n268), .B(n269), .Z(n964) );
  NAND U571 ( .A(n627), .B(n628), .Z(n270) );
  XOR U572 ( .A(n627), .B(n628), .Z(n271) );
  NANDN U573 ( .A(n626), .B(n271), .Z(n272) );
  NAND U574 ( .A(n270), .B(n272), .Z(n1013) );
  XOR U575 ( .A(n943), .B(n941), .Z(n273) );
  NANDN U576 ( .A(n942), .B(n273), .Z(n274) );
  NAND U577 ( .A(n943), .B(n941), .Z(n275) );
  AND U578 ( .A(n274), .B(n275), .Z(n1134) );
  NAND U579 ( .A(n915), .B(n916), .Z(n276) );
  XOR U580 ( .A(n915), .B(n916), .Z(n277) );
  NANDN U581 ( .A(n914), .B(n277), .Z(n278) );
  NAND U582 ( .A(n276), .B(n278), .Z(n1120) );
  NAND U583 ( .A(n958), .B(n956), .Z(n279) );
  XOR U584 ( .A(n958), .B(n956), .Z(n280) );
  NANDN U585 ( .A(n957), .B(n280), .Z(n281) );
  NAND U586 ( .A(n279), .B(n281), .Z(n1148) );
  XOR U587 ( .A(n967), .B(n965), .Z(n282) );
  NANDN U588 ( .A(n966), .B(n282), .Z(n283) );
  NAND U589 ( .A(n967), .B(n965), .Z(n284) );
  AND U590 ( .A(n283), .B(n284), .Z(n1142) );
  NAND U591 ( .A(n676), .B(n674), .Z(n285) );
  XOR U592 ( .A(n676), .B(n674), .Z(n286) );
  NANDN U593 ( .A(n675), .B(n286), .Z(n287) );
  NAND U594 ( .A(n285), .B(n287), .Z(n1053) );
  XOR U595 ( .A(n442), .B(n443), .Z(n288) );
  NANDN U596 ( .A(n444), .B(n288), .Z(n289) );
  NAND U597 ( .A(n442), .B(n443), .Z(n290) );
  AND U598 ( .A(n289), .B(n290), .Z(n1072) );
  NAND U599 ( .A(n1063), .B(n1064), .Z(n291) );
  XOR U600 ( .A(n1063), .B(n1064), .Z(n292) );
  NANDN U601 ( .A(n1062), .B(n292), .Z(n293) );
  NAND U602 ( .A(n291), .B(n293), .Z(n1195) );
  NAND U603 ( .A(n976), .B(n978), .Z(n294) );
  XOR U604 ( .A(n976), .B(n978), .Z(n295) );
  NAND U605 ( .A(n295), .B(n977), .Z(n296) );
  NAND U606 ( .A(n294), .B(n296), .Z(n1192) );
  NAND U607 ( .A(n1070), .B(n1071), .Z(n297) );
  XOR U608 ( .A(n1070), .B(n1071), .Z(n298) );
  NANDN U609 ( .A(n1069), .B(n298), .Z(n299) );
  NAND U610 ( .A(n297), .B(n299), .Z(n1123) );
  NAND U611 ( .A(n1110), .B(n1112), .Z(n300) );
  XOR U612 ( .A(n1110), .B(n1112), .Z(n301) );
  NAND U613 ( .A(n301), .B(n1111), .Z(n302) );
  NAND U614 ( .A(n300), .B(n302), .Z(n1261) );
  NAND U615 ( .A(n1135), .B(n1137), .Z(n303) );
  XOR U616 ( .A(n1135), .B(n1137), .Z(n304) );
  NAND U617 ( .A(n304), .B(n1136), .Z(n305) );
  NAND U618 ( .A(n303), .B(n305), .Z(n1258) );
  NAND U619 ( .A(n809), .B(n811), .Z(n306) );
  XOR U620 ( .A(n809), .B(n811), .Z(n307) );
  NAND U621 ( .A(n307), .B(n810), .Z(n308) );
  NAND U622 ( .A(n306), .B(n308), .Z(n1059) );
  NAND U623 ( .A(n763), .B(n764), .Z(n309) );
  XOR U624 ( .A(n763), .B(n764), .Z(n310) );
  NANDN U625 ( .A(n762), .B(n310), .Z(n311) );
  NAND U626 ( .A(n309), .B(n311), .Z(n1090) );
  NAND U627 ( .A(n894), .B(n896), .Z(n312) );
  XOR U628 ( .A(n894), .B(n896), .Z(n313) );
  NAND U629 ( .A(n313), .B(n895), .Z(n314) );
  NAND U630 ( .A(n312), .B(n314), .Z(n1107) );
  NANDN U631 ( .A(n1097), .B(n1100), .Z(n315) );
  OR U632 ( .A(n1100), .B(n1098), .Z(n316) );
  NAND U633 ( .A(n1099), .B(n316), .Z(n317) );
  NAND U634 ( .A(n315), .B(n317), .Z(n1161) );
  XNOR U635 ( .A(n485), .B(n484), .Z(n318) );
  XNOR U636 ( .A(n486), .B(n318), .Z(n756) );
  NAND U637 ( .A(n817), .B(n818), .Z(n319) );
  XOR U638 ( .A(n817), .B(n818), .Z(n320) );
  NANDN U639 ( .A(n816), .B(n320), .Z(n321) );
  NAND U640 ( .A(n319), .B(n321), .Z(n1001) );
  NAND U641 ( .A(n1300), .B(n1298), .Z(n322) );
  XOR U642 ( .A(n1300), .B(n1298), .Z(n323) );
  NANDN U643 ( .A(n1299), .B(n323), .Z(n324) );
  NAND U644 ( .A(n322), .B(n324), .Z(n1313) );
  NAND U645 ( .A(n1075), .B(n1077), .Z(n325) );
  XOR U646 ( .A(n1075), .B(n1077), .Z(n326) );
  NAND U647 ( .A(n326), .B(n1076), .Z(n327) );
  NAND U648 ( .A(n325), .B(n327), .Z(n1208) );
  OR U649 ( .A(n1295), .B(n1296), .Z(n328) );
  OR U650 ( .A(n1294), .B(n1293), .Z(n329) );
  AND U651 ( .A(n328), .B(n329), .Z(n1314) );
  NAND U652 ( .A(n891), .B(n892), .Z(n330) );
  XOR U653 ( .A(n891), .B(n892), .Z(n331) );
  NANDN U654 ( .A(n890), .B(n331), .Z(n332) );
  NAND U655 ( .A(n330), .B(n332), .Z(n1104) );
  NAND U656 ( .A(n1280), .B(n1281), .Z(n333) );
  XOR U657 ( .A(n1280), .B(n1281), .Z(n334) );
  NANDN U658 ( .A(n1279), .B(n334), .Z(n335) );
  NAND U659 ( .A(n333), .B(n335), .Z(n1285) );
  NAND U660 ( .A(n1290), .B(n1292), .Z(n336) );
  XOR U661 ( .A(n1290), .B(n1292), .Z(n337) );
  NAND U662 ( .A(n337), .B(n1291), .Z(n338) );
  NAND U663 ( .A(n336), .B(n338), .Z(n1319) );
  NAND U664 ( .A(n1331), .B(n1330), .Z(n339) );
  XOR U665 ( .A(n1331), .B(n1330), .Z(n340) );
  NANDN U666 ( .A(oglobal[7]), .B(n340), .Z(n341) );
  NAND U667 ( .A(n339), .B(n341), .Z(n1332) );
  XOR U668 ( .A(x[46]), .B(y[46]), .Z(n692) );
  XOR U669 ( .A(x[50]), .B(y[50]), .Z(n690) );
  XNOR U670 ( .A(x[48]), .B(y[48]), .Z(n691) );
  XOR U671 ( .A(n690), .B(n691), .Z(n693) );
  XOR U672 ( .A(n692), .B(n693), .Z(n837) );
  XOR U673 ( .A(x[52]), .B(y[52]), .Z(n680) );
  XOR U674 ( .A(x[56]), .B(y[56]), .Z(n678) );
  XNOR U675 ( .A(x[54]), .B(y[54]), .Z(n679) );
  XOR U676 ( .A(n678), .B(n679), .Z(n681) );
  XNOR U677 ( .A(n680), .B(n681), .Z(n838) );
  XOR U678 ( .A(x[40]), .B(y[40]), .Z(n568) );
  XOR U679 ( .A(x[44]), .B(y[44]), .Z(n566) );
  XNOR U680 ( .A(x[42]), .B(y[42]), .Z(n567) );
  XOR U681 ( .A(n566), .B(n567), .Z(n569) );
  XNOR U682 ( .A(n568), .B(n569), .Z(n836) );
  XNOR U683 ( .A(n838), .B(n836), .Z(n342) );
  XOR U684 ( .A(n837), .B(n342), .Z(n708) );
  XOR U685 ( .A(x[16]), .B(y[16]), .Z(n548) );
  XOR U686 ( .A(x[20]), .B(y[20]), .Z(n546) );
  XNOR U687 ( .A(x[18]), .B(y[18]), .Z(n547) );
  XOR U688 ( .A(n546), .B(n547), .Z(n549) );
  XOR U689 ( .A(n548), .B(n549), .Z(n834) );
  XOR U690 ( .A(x[10]), .B(y[10]), .Z(n542) );
  XOR U691 ( .A(x[14]), .B(y[14]), .Z(n540) );
  XNOR U692 ( .A(x[12]), .B(y[12]), .Z(n541) );
  XOR U693 ( .A(n540), .B(n541), .Z(n543) );
  XNOR U694 ( .A(n542), .B(n543), .Z(n833) );
  XOR U695 ( .A(x[4]), .B(y[4]), .Z(n510) );
  XOR U696 ( .A(x[8]), .B(y[8]), .Z(n508) );
  XNOR U697 ( .A(x[6]), .B(y[6]), .Z(n509) );
  XOR U698 ( .A(n508), .B(n509), .Z(n511) );
  XOR U699 ( .A(n510), .B(n511), .Z(n832) );
  XOR U700 ( .A(n833), .B(n832), .Z(n343) );
  XOR U701 ( .A(n834), .B(n343), .Z(n706) );
  XOR U702 ( .A(x[34]), .B(y[34]), .Z(n575) );
  XOR U703 ( .A(x[38]), .B(y[38]), .Z(n573) );
  XOR U704 ( .A(x[36]), .B(y[36]), .Z(n572) );
  XNOR U705 ( .A(n573), .B(n572), .Z(n574) );
  XOR U706 ( .A(n575), .B(n574), .Z(n850) );
  XOR U707 ( .A(x[22]), .B(y[22]), .Z(n523) );
  XOR U708 ( .A(x[26]), .B(y[26]), .Z(n521) );
  XNOR U709 ( .A(x[24]), .B(y[24]), .Z(n522) );
  XOR U710 ( .A(n521), .B(n522), .Z(n524) );
  XNOR U711 ( .A(n523), .B(n524), .Z(n849) );
  XOR U712 ( .A(x[28]), .B(y[28]), .Z(n529) );
  XOR U713 ( .A(x[32]), .B(y[32]), .Z(n527) );
  XNOR U714 ( .A(x[30]), .B(y[30]), .Z(n528) );
  XOR U715 ( .A(n527), .B(n528), .Z(n530) );
  XOR U716 ( .A(n529), .B(n530), .Z(n848) );
  XOR U717 ( .A(n849), .B(n848), .Z(n344) );
  XNOR U718 ( .A(n850), .B(n344), .Z(n705) );
  XNOR U719 ( .A(n706), .B(n705), .Z(n707) );
  XNOR U720 ( .A(n708), .B(n707), .Z(n821) );
  XOR U721 ( .A(x[147]), .B(y[147]), .Z(n609) );
  XOR U722 ( .A(x[173]), .B(y[173]), .Z(n607) );
  XNOR U723 ( .A(x[145]), .B(y[145]), .Z(n608) );
  XOR U724 ( .A(n607), .B(n608), .Z(n610) );
  XOR U725 ( .A(n609), .B(n610), .Z(n868) );
  XOR U726 ( .A(x[143]), .B(y[143]), .Z(n792) );
  XOR U727 ( .A(x[175]), .B(y[175]), .Z(n790) );
  XNOR U728 ( .A(x[141]), .B(y[141]), .Z(n791) );
  XOR U729 ( .A(n790), .B(n791), .Z(n793) );
  XNOR U730 ( .A(n792), .B(n793), .Z(n869) );
  XOR U731 ( .A(x[163]), .B(y[163]), .Z(n621) );
  XOR U732 ( .A(x[161]), .B(y[161]), .Z(n619) );
  XNOR U733 ( .A(x[159]), .B(y[159]), .Z(n620) );
  XOR U734 ( .A(n619), .B(n620), .Z(n622) );
  XNOR U735 ( .A(n621), .B(n622), .Z(n867) );
  XNOR U736 ( .A(n869), .B(n867), .Z(n345) );
  XNOR U737 ( .A(n868), .B(n345), .Z(n818) );
  XOR U738 ( .A(x[135]), .B(y[135]), .Z(n798) );
  XOR U739 ( .A(x[179]), .B(y[179]), .Z(n796) );
  XNOR U740 ( .A(x[133]), .B(y[133]), .Z(n797) );
  XOR U741 ( .A(n796), .B(n797), .Z(n799) );
  XOR U742 ( .A(n798), .B(n799), .Z(n728) );
  XOR U743 ( .A(x[131]), .B(y[131]), .Z(n418) );
  XOR U744 ( .A(x[181]), .B(y[181]), .Z(n416) );
  XNOR U745 ( .A(x[129]), .B(y[129]), .Z(n417) );
  XOR U746 ( .A(n416), .B(n417), .Z(n419) );
  XNOR U747 ( .A(n418), .B(n419), .Z(n729) );
  XOR U748 ( .A(x[139]), .B(y[139]), .Z(n804) );
  XOR U749 ( .A(x[177]), .B(y[177]), .Z(n802) );
  XNOR U750 ( .A(x[137]), .B(y[137]), .Z(n803) );
  XOR U751 ( .A(n802), .B(n803), .Z(n805) );
  XNOR U752 ( .A(n804), .B(n805), .Z(n727) );
  XNOR U753 ( .A(n729), .B(n727), .Z(n346) );
  XNOR U754 ( .A(n728), .B(n346), .Z(n817) );
  XOR U755 ( .A(x[81]), .B(y[81]), .Z(n425) );
  XOR U756 ( .A(x[79]), .B(y[79]), .Z(n423) );
  XNOR U757 ( .A(x[77]), .B(y[77]), .Z(n424) );
  XOR U758 ( .A(n423), .B(n424), .Z(n426) );
  XOR U759 ( .A(n425), .B(n426), .Z(n675) );
  XOR U760 ( .A(x[75]), .B(y[75]), .Z(n460) );
  XOR U761 ( .A(x[73]), .B(y[73]), .Z(n458) );
  XNOR U762 ( .A(x[71]), .B(y[71]), .Z(n459) );
  XOR U763 ( .A(n458), .B(n459), .Z(n461) );
  XNOR U764 ( .A(n460), .B(n461), .Z(n676) );
  XOR U765 ( .A(x[87]), .B(y[87]), .Z(n431) );
  XOR U766 ( .A(x[85]), .B(y[85]), .Z(n429) );
  XNOR U767 ( .A(x[83]), .B(y[83]), .Z(n430) );
  XOR U768 ( .A(n429), .B(n430), .Z(n432) );
  XNOR U769 ( .A(n431), .B(n432), .Z(n674) );
  XNOR U770 ( .A(n676), .B(n674), .Z(n347) );
  XOR U771 ( .A(n675), .B(n347), .Z(n490) );
  XOR U772 ( .A(x[99]), .B(y[99]), .Z(n467) );
  XOR U773 ( .A(x[97]), .B(y[97]), .Z(n465) );
  XNOR U774 ( .A(x[95]), .B(y[95]), .Z(n466) );
  XOR U775 ( .A(n465), .B(n466), .Z(n468) );
  XOR U776 ( .A(n467), .B(n468), .Z(n648) );
  XOR U777 ( .A(x[93]), .B(y[93]), .Z(n437) );
  XOR U778 ( .A(x[91]), .B(y[91]), .Z(n435) );
  XNOR U779 ( .A(x[89]), .B(y[89]), .Z(n436) );
  XOR U780 ( .A(n435), .B(n436), .Z(n438) );
  XNOR U781 ( .A(n437), .B(n438), .Z(n649) );
  XOR U782 ( .A(x[103]), .B(y[103]), .Z(n473) );
  XOR U783 ( .A(x[195]), .B(y[195]), .Z(n471) );
  XNOR U784 ( .A(x[101]), .B(y[101]), .Z(n472) );
  XOR U785 ( .A(n471), .B(n472), .Z(n474) );
  XNOR U786 ( .A(n473), .B(n474), .Z(n647) );
  XNOR U787 ( .A(n649), .B(n647), .Z(n348) );
  XOR U788 ( .A(n648), .B(n348), .Z(n491) );
  XOR U789 ( .A(x[63]), .B(y[63]), .Z(n448) );
  XOR U790 ( .A(x[61]), .B(y[61]), .Z(n446) );
  XNOR U791 ( .A(x[59]), .B(y[59]), .Z(n447) );
  XOR U792 ( .A(n446), .B(n447), .Z(n449) );
  XOR U793 ( .A(n448), .B(n449), .Z(n672) );
  XOR U794 ( .A(x[57]), .B(y[57]), .Z(n785) );
  XOR U795 ( .A(x[55]), .B(y[55]), .Z(n783) );
  XNOR U796 ( .A(x[53]), .B(y[53]), .Z(n784) );
  XOR U797 ( .A(n783), .B(n784), .Z(n786) );
  XNOR U798 ( .A(n785), .B(n786), .Z(n673) );
  XOR U799 ( .A(x[69]), .B(y[69]), .Z(n454) );
  XOR U800 ( .A(x[67]), .B(y[67]), .Z(n452) );
  XNOR U801 ( .A(x[65]), .B(y[65]), .Z(n453) );
  XOR U802 ( .A(n452), .B(n453), .Z(n455) );
  XNOR U803 ( .A(n454), .B(n455), .Z(n671) );
  XNOR U804 ( .A(n673), .B(n671), .Z(n349) );
  XNOR U805 ( .A(n672), .B(n349), .Z(n489) );
  XOR U806 ( .A(n491), .B(n489), .Z(n350) );
  XNOR U807 ( .A(n490), .B(n350), .Z(n816) );
  XOR U808 ( .A(n817), .B(n816), .Z(n351) );
  XOR U809 ( .A(n818), .B(n351), .Z(n822) );
  XOR U810 ( .A(x[184]), .B(y[184]), .Z(n516) );
  XOR U811 ( .A(x[188]), .B(y[188]), .Z(n515) );
  XOR U812 ( .A(x[186]), .B(y[186]), .Z(n514) );
  XOR U813 ( .A(n515), .B(n514), .Z(n517) );
  XNOR U814 ( .A(n516), .B(n517), .Z(n442) );
  XOR U815 ( .A(x[154]), .B(y[154]), .Z(n657) );
  XOR U816 ( .A(x[158]), .B(y[158]), .Z(n655) );
  XOR U817 ( .A(x[156]), .B(y[156]), .Z(n654) );
  XNOR U818 ( .A(n655), .B(n654), .Z(n656) );
  XNOR U819 ( .A(n657), .B(n656), .Z(n444) );
  XOR U820 ( .A(x[148]), .B(y[148]), .Z(n645) );
  XOR U821 ( .A(x[152]), .B(y[152]), .Z(n643) );
  XOR U822 ( .A(x[150]), .B(y[150]), .Z(n642) );
  XNOR U823 ( .A(n643), .B(n642), .Z(n644) );
  XOR U824 ( .A(n645), .B(n644), .Z(n443) );
  XOR U825 ( .A(x[166]), .B(y[166]), .Z(n562) );
  XOR U826 ( .A(x[170]), .B(y[170]), .Z(n560) );
  XNOR U827 ( .A(x[168]), .B(y[168]), .Z(n561) );
  XOR U828 ( .A(n560), .B(n561), .Z(n563) );
  XOR U829 ( .A(n562), .B(n563), .Z(n755) );
  XOR U830 ( .A(x[190]), .B(y[190]), .Z(n858) );
  XOR U831 ( .A(x[194]), .B(y[194]), .Z(n857) );
  XOR U832 ( .A(x[192]), .B(y[192]), .Z(n856) );
  XOR U833 ( .A(n857), .B(n856), .Z(n859) );
  XNOR U834 ( .A(n858), .B(n859), .Z(n484) );
  XOR U835 ( .A(x[142]), .B(y[142]), .Z(n722) );
  XOR U836 ( .A(x[146]), .B(y[146]), .Z(n720) );
  XOR U837 ( .A(x[144]), .B(y[144]), .Z(n719) );
  XNOR U838 ( .A(n720), .B(n719), .Z(n721) );
  XNOR U839 ( .A(n722), .B(n721), .Z(n486) );
  XOR U840 ( .A(x[136]), .B(y[136]), .Z(n741) );
  XOR U841 ( .A(x[140]), .B(y[140]), .Z(n739) );
  XOR U842 ( .A(x[138]), .B(y[138]), .Z(n738) );
  XNOR U843 ( .A(n739), .B(n738), .Z(n740) );
  XOR U844 ( .A(n741), .B(n740), .Z(n485) );
  XOR U845 ( .A(n755), .B(n756), .Z(n352) );
  XOR U846 ( .A(n757), .B(n352), .Z(n820) );
  XNOR U847 ( .A(n822), .B(n820), .Z(n353) );
  XNOR U848 ( .A(n821), .B(n353), .Z(n891) );
  XOR U849 ( .A(x[178]), .B(y[178]), .Z(n554) );
  XOR U850 ( .A(x[182]), .B(y[182]), .Z(n552) );
  XNOR U851 ( .A(x[180]), .B(y[180]), .Z(n553) );
  XOR U852 ( .A(n552), .B(n553), .Z(n555) );
  XOR U853 ( .A(n554), .B(n555), .Z(n626) );
  XOR U854 ( .A(x[160]), .B(y[160]), .Z(n686) );
  XOR U855 ( .A(x[164]), .B(y[164]), .Z(n684) );
  XNOR U856 ( .A(x[162]), .B(y[162]), .Z(n685) );
  XOR U857 ( .A(n684), .B(n685), .Z(n687) );
  XNOR U858 ( .A(n686), .B(n687), .Z(n628) );
  XOR U859 ( .A(x[172]), .B(y[172]), .Z(n535) );
  XOR U860 ( .A(x[176]), .B(y[176]), .Z(n533) );
  XNOR U861 ( .A(x[174]), .B(y[174]), .Z(n534) );
  XOR U862 ( .A(n533), .B(n534), .Z(n536) );
  XNOR U863 ( .A(n535), .B(n536), .Z(n627) );
  XNOR U864 ( .A(n628), .B(n627), .Z(n354) );
  XNOR U865 ( .A(n626), .B(n354), .Z(n813) );
  XOR U866 ( .A(x[199]), .B(y[199]), .Z(n395) );
  XNOR U867 ( .A(x[2]), .B(y[2]), .Z(n394) );
  XNOR U868 ( .A(n395), .B(n394), .Z(n397) );
  XNOR U869 ( .A(x[197]), .B(y[197]), .Z(n396) );
  XNOR U870 ( .A(n397), .B(n396), .Z(n826) );
  XOR U871 ( .A(x[122]), .B(y[122]), .Z(n735) );
  XNOR U872 ( .A(x[120]), .B(y[120]), .Z(n734) );
  XNOR U873 ( .A(n735), .B(n734), .Z(n737) );
  XNOR U874 ( .A(x[118]), .B(y[118]), .Z(n736) );
  XNOR U875 ( .A(n737), .B(n736), .Z(n829) );
  XOR U876 ( .A(x[116]), .B(y[116]), .Z(n578) );
  XNOR U877 ( .A(x[114]), .B(y[114]), .Z(n577) );
  XNOR U878 ( .A(n578), .B(n577), .Z(n580) );
  XNOR U879 ( .A(x[112]), .B(y[112]), .Z(n579) );
  XNOR U880 ( .A(n580), .B(n579), .Z(n827) );
  XNOR U881 ( .A(n829), .B(n827), .Z(n355) );
  XNOR U882 ( .A(n826), .B(n355), .Z(n815) );
  XOR U883 ( .A(x[130]), .B(y[130]), .Z(n745) );
  XOR U884 ( .A(x[134]), .B(y[134]), .Z(n743) );
  XOR U885 ( .A(x[132]), .B(y[132]), .Z(n742) );
  XNOR U886 ( .A(n743), .B(n742), .Z(n744) );
  XNOR U887 ( .A(n745), .B(n744), .Z(n825) );
  XOR U888 ( .A(x[128]), .B(y[128]), .Z(n731) );
  XNOR U889 ( .A(x[126]), .B(y[126]), .Z(n730) );
  XNOR U890 ( .A(n731), .B(n730), .Z(n733) );
  XNOR U891 ( .A(x[124]), .B(y[124]), .Z(n732) );
  XNOR U892 ( .A(n733), .B(n732), .Z(n824) );
  XOR U893 ( .A(x[196]), .B(y[196]), .Z(n379) );
  XOR U894 ( .A(x[198]), .B(y[198]), .Z(n377) );
  XNOR U895 ( .A(n377), .B(oglobal[0]), .Z(n378) );
  XNOR U896 ( .A(n379), .B(n378), .Z(n823) );
  XNOR U897 ( .A(n824), .B(n823), .Z(n356) );
  XNOR U898 ( .A(n825), .B(n356), .Z(n814) );
  XNOR U899 ( .A(n815), .B(n814), .Z(n357) );
  XOR U900 ( .A(n813), .B(n357), .Z(n890) );
  XOR U901 ( .A(x[165]), .B(y[165]), .Z(n597) );
  XOR U902 ( .A(x[169]), .B(y[169]), .Z(n594) );
  XNOR U903 ( .A(x[167]), .B(y[167]), .Z(n595) );
  XNOR U904 ( .A(n594), .B(n595), .Z(n596) );
  XNOR U905 ( .A(n597), .B(n596), .Z(n389) );
  XOR U906 ( .A(x[151]), .B(y[151]), .Z(n616) );
  XOR U907 ( .A(x[171]), .B(y[171]), .Z(n613) );
  XNOR U908 ( .A(x[149]), .B(y[149]), .Z(n614) );
  XNOR U909 ( .A(n613), .B(n614), .Z(n615) );
  XNOR U910 ( .A(n616), .B(n615), .Z(n388) );
  XOR U911 ( .A(x[155]), .B(y[155]), .Z(n603) );
  XOR U912 ( .A(x[157]), .B(y[157]), .Z(n600) );
  XNOR U913 ( .A(x[153]), .B(y[153]), .Z(n601) );
  XNOR U914 ( .A(n600), .B(n601), .Z(n602) );
  XOR U915 ( .A(n603), .B(n602), .Z(n387) );
  XOR U916 ( .A(n388), .B(n387), .Z(n358) );
  XNOR U917 ( .A(n389), .B(n358), .Z(n764) );
  XOR U918 ( .A(x[127]), .B(y[127]), .Z(n406) );
  XOR U919 ( .A(x[183]), .B(y[183]), .Z(n404) );
  XNOR U920 ( .A(x[125]), .B(y[125]), .Z(n405) );
  XOR U921 ( .A(n404), .B(n405), .Z(n407) );
  XOR U922 ( .A(n406), .B(n407), .Z(n591) );
  XOR U923 ( .A(x[119]), .B(y[119]), .Z(n885) );
  XOR U924 ( .A(x[187]), .B(y[187]), .Z(n883) );
  XOR U925 ( .A(x[117]), .B(y[117]), .Z(n882) );
  XNOR U926 ( .A(n883), .B(n882), .Z(n884) );
  XNOR U927 ( .A(n885), .B(n884), .Z(n592) );
  XOR U928 ( .A(x[123]), .B(y[123]), .Z(n412) );
  XOR U929 ( .A(x[185]), .B(y[185]), .Z(n410) );
  XNOR U930 ( .A(x[121]), .B(y[121]), .Z(n411) );
  XOR U931 ( .A(n410), .B(n411), .Z(n413) );
  XNOR U932 ( .A(n412), .B(n413), .Z(n590) );
  XNOR U933 ( .A(n592), .B(n590), .Z(n359) );
  XNOR U934 ( .A(n591), .B(n359), .Z(n763) );
  XOR U935 ( .A(x[111]), .B(y[111]), .Z(n872) );
  XOR U936 ( .A(x[191]), .B(y[191]), .Z(n870) );
  XNOR U937 ( .A(x[109]), .B(y[109]), .Z(n871) );
  XOR U938 ( .A(n870), .B(n871), .Z(n873) );
  XOR U939 ( .A(n872), .B(n873), .Z(n651) );
  XOR U940 ( .A(x[107]), .B(y[107]), .Z(n479) );
  XOR U941 ( .A(x[193]), .B(y[193]), .Z(n477) );
  XNOR U942 ( .A(x[105]), .B(y[105]), .Z(n478) );
  XOR U943 ( .A(n477), .B(n478), .Z(n480) );
  XNOR U944 ( .A(n479), .B(n480), .Z(n652) );
  XOR U945 ( .A(x[115]), .B(y[115]), .Z(n878) );
  XOR U946 ( .A(x[189]), .B(y[189]), .Z(n876) );
  XNOR U947 ( .A(x[113]), .B(y[113]), .Z(n877) );
  XOR U948 ( .A(n876), .B(n877), .Z(n879) );
  XNOR U949 ( .A(n878), .B(n879), .Z(n650) );
  XNOR U950 ( .A(n652), .B(n650), .Z(n360) );
  XOR U951 ( .A(n651), .B(n360), .Z(n762) );
  XOR U952 ( .A(n763), .B(n762), .Z(n361) );
  XOR U953 ( .A(n764), .B(n361), .Z(n767) );
  XOR U954 ( .A(x[88]), .B(y[88]), .Z(n718) );
  XOR U955 ( .A(x[92]), .B(y[92]), .Z(n716) );
  XOR U956 ( .A(x[90]), .B(y[90]), .Z(n715) );
  XNOR U957 ( .A(n716), .B(n715), .Z(n717) );
  XOR U958 ( .A(n718), .B(n717), .Z(n845) );
  XOR U959 ( .A(x[82]), .B(y[82]), .Z(n714) );
  XOR U960 ( .A(x[86]), .B(y[86]), .Z(n712) );
  XOR U961 ( .A(x[84]), .B(y[84]), .Z(n711) );
  XNOR U962 ( .A(n712), .B(n711), .Z(n713) );
  XNOR U963 ( .A(n714), .B(n713), .Z(n847) );
  XOR U964 ( .A(x[76]), .B(y[76]), .Z(n641) );
  XOR U965 ( .A(x[80]), .B(y[80]), .Z(n639) );
  XOR U966 ( .A(x[78]), .B(y[78]), .Z(n638) );
  XNOR U967 ( .A(n639), .B(n638), .Z(n640) );
  XNOR U968 ( .A(n641), .B(n640), .Z(n846) );
  XNOR U969 ( .A(n847), .B(n846), .Z(n362) );
  XNOR U970 ( .A(n845), .B(n362), .Z(n497) );
  XOR U971 ( .A(x[100]), .B(y[100]), .Z(n588) );
  XOR U972 ( .A(x[104]), .B(y[104]), .Z(n586) );
  XOR U973 ( .A(x[102]), .B(y[102]), .Z(n585) );
  XNOR U974 ( .A(n586), .B(n585), .Z(n587) );
  XOR U975 ( .A(n588), .B(n587), .Z(n842) );
  XOR U976 ( .A(x[106]), .B(y[106]), .Z(n584) );
  XOR U977 ( .A(x[110]), .B(y[110]), .Z(n582) );
  XOR U978 ( .A(x[108]), .B(y[108]), .Z(n581) );
  XNOR U979 ( .A(n582), .B(n581), .Z(n583) );
  XNOR U980 ( .A(n584), .B(n583), .Z(n844) );
  XOR U981 ( .A(x[94]), .B(y[94]), .Z(n752) );
  XOR U982 ( .A(x[98]), .B(y[98]), .Z(n750) );
  XOR U983 ( .A(x[96]), .B(y[96]), .Z(n749) );
  XNOR U984 ( .A(n750), .B(n749), .Z(n751) );
  XNOR U985 ( .A(n752), .B(n751), .Z(n843) );
  XNOR U986 ( .A(n844), .B(n843), .Z(n363) );
  XNOR U987 ( .A(n842), .B(n363), .Z(n496) );
  XOR U988 ( .A(x[64]), .B(y[64]), .Z(n660) );
  XOR U989 ( .A(x[66]), .B(y[66]), .Z(n658) );
  XNOR U990 ( .A(x[68]), .B(y[68]), .Z(n659) );
  XOR U991 ( .A(n658), .B(n659), .Z(n661) );
  XOR U992 ( .A(n660), .B(n661), .Z(n841) );
  XOR U993 ( .A(x[70]), .B(y[70]), .Z(n634) );
  XOR U994 ( .A(x[74]), .B(y[74]), .Z(n632) );
  XNOR U995 ( .A(x[72]), .B(y[72]), .Z(n633) );
  XOR U996 ( .A(n632), .B(n633), .Z(n635) );
  XNOR U997 ( .A(n634), .B(n635), .Z(n840) );
  XOR U998 ( .A(x[58]), .B(y[58]), .Z(n666) );
  XOR U999 ( .A(x[62]), .B(y[62]), .Z(n664) );
  XNOR U1000 ( .A(x[60]), .B(y[60]), .Z(n665) );
  XOR U1001 ( .A(n664), .B(n665), .Z(n667) );
  XOR U1002 ( .A(n666), .B(n667), .Z(n839) );
  XOR U1003 ( .A(n840), .B(n839), .Z(n364) );
  XOR U1004 ( .A(n841), .B(n364), .Z(n495) );
  XOR U1005 ( .A(n496), .B(n495), .Z(n365) );
  XNOR U1006 ( .A(n497), .B(n365), .Z(n769) );
  XOR U1007 ( .A(x[27]), .B(y[27]), .Z(n382) );
  XOR U1008 ( .A(x[25]), .B(y[25]), .Z(n380) );
  XNOR U1009 ( .A(x[23]), .B(y[23]), .Z(n381) );
  XOR U1010 ( .A(n380), .B(n381), .Z(n383) );
  XOR U1011 ( .A(n382), .B(n383), .Z(n697) );
  XOR U1012 ( .A(x[21]), .B(y[21]), .Z(n373) );
  XOR U1013 ( .A(x[19]), .B(y[19]), .Z(n371) );
  XNOR U1014 ( .A(x[17]), .B(y[17]), .Z(n372) );
  XOR U1015 ( .A(n371), .B(n372), .Z(n374) );
  XNOR U1016 ( .A(n373), .B(n374), .Z(n699) );
  XOR U1017 ( .A(x[33]), .B(y[33]), .Z(n393) );
  XOR U1018 ( .A(x[31]), .B(y[31]), .Z(n391) );
  XOR U1019 ( .A(x[29]), .B(y[29]), .Z(n390) );
  XNOR U1020 ( .A(n391), .B(n390), .Z(n392) );
  XNOR U1021 ( .A(n393), .B(n392), .Z(n698) );
  XNOR U1022 ( .A(n699), .B(n698), .Z(n366) );
  XNOR U1023 ( .A(n697), .B(n366), .Z(n494) );
  XOR U1024 ( .A(x[45]), .B(y[45]), .Z(n773) );
  XOR U1025 ( .A(x[43]), .B(y[43]), .Z(n771) );
  XNOR U1026 ( .A(x[41]), .B(y[41]), .Z(n772) );
  XOR U1027 ( .A(n771), .B(n772), .Z(n774) );
  XOR U1028 ( .A(n773), .B(n774), .Z(n701) );
  XOR U1029 ( .A(x[39]), .B(y[39]), .Z(n401) );
  XOR U1030 ( .A(x[37]), .B(y[37]), .Z(n399) );
  XOR U1031 ( .A(x[35]), .B(y[35]), .Z(n398) );
  XNOR U1032 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U1033 ( .A(n401), .B(n400), .Z(n702) );
  XOR U1034 ( .A(x[51]), .B(y[51]), .Z(n779) );
  XOR U1035 ( .A(x[49]), .B(y[49]), .Z(n777) );
  XNOR U1036 ( .A(x[47]), .B(y[47]), .Z(n778) );
  XOR U1037 ( .A(n777), .B(n778), .Z(n780) );
  XNOR U1038 ( .A(n779), .B(n780), .Z(n700) );
  XNOR U1039 ( .A(n702), .B(n700), .Z(n367) );
  XOR U1040 ( .A(n701), .B(n367), .Z(n493) );
  XOR U1041 ( .A(x[3]), .B(y[3]), .Z(n504) );
  XOR U1042 ( .A(x[1]), .B(y[1]), .Z(n502) );
  XNOR U1043 ( .A(x[0]), .B(y[0]), .Z(n503) );
  XOR U1044 ( .A(n502), .B(n503), .Z(n505) );
  XNOR U1045 ( .A(n504), .B(n505), .Z(n811) );
  XOR U1046 ( .A(x[13]), .B(y[13]), .Z(n863) );
  XNOR U1047 ( .A(x[11]), .B(y[11]), .Z(n862) );
  XNOR U1048 ( .A(n863), .B(n862), .Z(n865) );
  XNOR U1049 ( .A(x[15]), .B(y[15]), .Z(n864) );
  XNOR U1050 ( .A(n865), .B(n864), .Z(n810) );
  XOR U1051 ( .A(x[7]), .B(y[7]), .Z(n853) );
  XNOR U1052 ( .A(x[5]), .B(y[5]), .Z(n852) );
  XNOR U1053 ( .A(n853), .B(n852), .Z(n855) );
  XNOR U1054 ( .A(x[9]), .B(y[9]), .Z(n854) );
  XNOR U1055 ( .A(n855), .B(n854), .Z(n809) );
  XNOR U1056 ( .A(n810), .B(n809), .Z(n368) );
  XOR U1057 ( .A(n811), .B(n368), .Z(n492) );
  XOR U1058 ( .A(n493), .B(n492), .Z(n369) );
  XOR U1059 ( .A(n494), .B(n369), .Z(n768) );
  XNOR U1060 ( .A(n890), .B(n892), .Z(n370) );
  XNOR U1061 ( .A(n891), .B(n370), .Z(o[0]) );
  NANDN U1062 ( .A(n372), .B(n371), .Z(n376) );
  NANDN U1063 ( .A(n374), .B(n373), .Z(n375) );
  NAND U1064 ( .A(n376), .B(n375), .Z(n916) );
  NANDN U1065 ( .A(n381), .B(n380), .Z(n385) );
  NANDN U1066 ( .A(n383), .B(n382), .Z(n384) );
  AND U1067 ( .A(n385), .B(n384), .Z(n914) );
  XOR U1068 ( .A(n915), .B(n914), .Z(n386) );
  XNOR U1069 ( .A(n916), .B(n386), .Z(n1021) );
  XOR U1070 ( .A(n992), .B(n991), .Z(n402) );
  XNOR U1071 ( .A(n993), .B(n402), .Z(n1020) );
  IV U1072 ( .A(n1020), .Z(n1018) );
  XNOR U1073 ( .A(n1019), .B(n1018), .Z(n403) );
  XOR U1074 ( .A(n1021), .B(n403), .Z(n1006) );
  NANDN U1075 ( .A(n405), .B(n404), .Z(n409) );
  NANDN U1076 ( .A(n407), .B(n406), .Z(n408) );
  NAND U1077 ( .A(n409), .B(n408), .Z(n932) );
  NANDN U1078 ( .A(n411), .B(n410), .Z(n415) );
  NANDN U1079 ( .A(n413), .B(n412), .Z(n414) );
  AND U1080 ( .A(n415), .B(n414), .Z(n933) );
  NANDN U1081 ( .A(n417), .B(n416), .Z(n421) );
  NANDN U1082 ( .A(n419), .B(n418), .Z(n420) );
  AND U1083 ( .A(n421), .B(n420), .Z(n931) );
  XNOR U1084 ( .A(n933), .B(n931), .Z(n422) );
  XOR U1085 ( .A(n932), .B(n422), .Z(n1074) );
  NANDN U1086 ( .A(n424), .B(n423), .Z(n428) );
  NANDN U1087 ( .A(n426), .B(n425), .Z(n427) );
  AND U1088 ( .A(n428), .B(n427), .Z(n943) );
  NANDN U1089 ( .A(n430), .B(n429), .Z(n434) );
  NANDN U1090 ( .A(n432), .B(n431), .Z(n433) );
  NAND U1091 ( .A(n434), .B(n433), .Z(n942) );
  NANDN U1092 ( .A(n436), .B(n435), .Z(n440) );
  NANDN U1093 ( .A(n438), .B(n437), .Z(n439) );
  AND U1094 ( .A(n440), .B(n439), .Z(n941) );
  XOR U1095 ( .A(n942), .B(n941), .Z(n441) );
  XNOR U1096 ( .A(n943), .B(n441), .Z(n1073) );
  XNOR U1097 ( .A(n1073), .B(n1072), .Z(n445) );
  XNOR U1098 ( .A(n1074), .B(n445), .Z(n1008) );
  NANDN U1099 ( .A(n447), .B(n446), .Z(n451) );
  NANDN U1100 ( .A(n449), .B(n448), .Z(n450) );
  AND U1101 ( .A(n451), .B(n450), .Z(n940) );
  NANDN U1102 ( .A(n453), .B(n452), .Z(n457) );
  NANDN U1103 ( .A(n455), .B(n454), .Z(n456) );
  NAND U1104 ( .A(n457), .B(n456), .Z(n939) );
  NANDN U1105 ( .A(n459), .B(n458), .Z(n463) );
  NANDN U1106 ( .A(n461), .B(n460), .Z(n462) );
  AND U1107 ( .A(n463), .B(n462), .Z(n938) );
  XOR U1108 ( .A(n939), .B(n938), .Z(n464) );
  XNOR U1109 ( .A(n940), .B(n464), .Z(n1071) );
  NANDN U1110 ( .A(n466), .B(n465), .Z(n470) );
  NANDN U1111 ( .A(n468), .B(n467), .Z(n469) );
  AND U1112 ( .A(n470), .B(n469), .Z(n946) );
  NANDN U1113 ( .A(n472), .B(n471), .Z(n476) );
  NANDN U1114 ( .A(n474), .B(n473), .Z(n475) );
  NAND U1115 ( .A(n476), .B(n475), .Z(n945) );
  NANDN U1116 ( .A(n478), .B(n477), .Z(n482) );
  NANDN U1117 ( .A(n480), .B(n479), .Z(n481) );
  AND U1118 ( .A(n482), .B(n481), .Z(n944) );
  XOR U1119 ( .A(n945), .B(n944), .Z(n483) );
  XNOR U1120 ( .A(n946), .B(n483), .Z(n1070) );
  XNOR U1121 ( .A(n1070), .B(n1069), .Z(n487) );
  XNOR U1122 ( .A(n1071), .B(n487), .Z(n1007) );
  XNOR U1123 ( .A(n1008), .B(n1007), .Z(n488) );
  XNOR U1124 ( .A(n1006), .B(n488), .Z(n1077) );
  NANDN U1125 ( .A(n496), .B(n495), .Z(n500) );
  ANDN U1126 ( .B(n496), .A(n495), .Z(n498) );
  OR U1127 ( .A(n498), .B(n497), .Z(n499) );
  AND U1128 ( .A(n500), .B(n499), .Z(n996) );
  XNOR U1129 ( .A(n998), .B(n996), .Z(n501) );
  XNOR U1130 ( .A(n997), .B(n501), .Z(n1075) );
  IV U1131 ( .A(n1075), .Z(n630) );
  NANDN U1132 ( .A(n503), .B(n502), .Z(n507) );
  NANDN U1133 ( .A(n505), .B(n504), .Z(n506) );
  NAND U1134 ( .A(n507), .B(n506), .Z(n952) );
  NANDN U1135 ( .A(n509), .B(n508), .Z(n513) );
  NANDN U1136 ( .A(n511), .B(n510), .Z(n512) );
  AND U1137 ( .A(n513), .B(n512), .Z(n954) );
  NAND U1138 ( .A(n515), .B(n514), .Z(n519) );
  NAND U1139 ( .A(n517), .B(n516), .Z(n518) );
  AND U1140 ( .A(n519), .B(n518), .Z(n953) );
  XNOR U1141 ( .A(n954), .B(n953), .Z(n520) );
  XNOR U1142 ( .A(n952), .B(n520), .Z(n1064) );
  NANDN U1143 ( .A(n522), .B(n521), .Z(n526) );
  NANDN U1144 ( .A(n524), .B(n523), .Z(n525) );
  AND U1145 ( .A(n526), .B(n525), .Z(n1041) );
  NANDN U1146 ( .A(n528), .B(n527), .Z(n532) );
  NANDN U1147 ( .A(n530), .B(n529), .Z(n531) );
  AND U1148 ( .A(n532), .B(n531), .Z(n1043) );
  NANDN U1149 ( .A(n534), .B(n533), .Z(n538) );
  NANDN U1150 ( .A(n536), .B(n535), .Z(n537) );
  NAND U1151 ( .A(n538), .B(n537), .Z(n1042) );
  XOR U1152 ( .A(n1043), .B(n1042), .Z(n539) );
  XOR U1153 ( .A(n1041), .B(n539), .Z(n1063) );
  NANDN U1154 ( .A(n541), .B(n540), .Z(n545) );
  NANDN U1155 ( .A(n543), .B(n542), .Z(n544) );
  AND U1156 ( .A(n545), .B(n544), .Z(n950) );
  NANDN U1157 ( .A(n547), .B(n546), .Z(n551) );
  NANDN U1158 ( .A(n549), .B(n548), .Z(n550) );
  AND U1159 ( .A(n551), .B(n550), .Z(n951) );
  NANDN U1160 ( .A(n553), .B(n552), .Z(n557) );
  NANDN U1161 ( .A(n555), .B(n554), .Z(n556) );
  NAND U1162 ( .A(n557), .B(n556), .Z(n949) );
  XOR U1163 ( .A(n951), .B(n949), .Z(n558) );
  XNOR U1164 ( .A(n950), .B(n558), .Z(n1062) );
  XOR U1165 ( .A(n1063), .B(n1062), .Z(n559) );
  XOR U1166 ( .A(n1064), .B(n559), .Z(n1003) );
  NANDN U1167 ( .A(n561), .B(n560), .Z(n565) );
  NANDN U1168 ( .A(n563), .B(n562), .Z(n564) );
  NAND U1169 ( .A(n565), .B(n564), .Z(n957) );
  NANDN U1170 ( .A(n567), .B(n566), .Z(n571) );
  NANDN U1171 ( .A(n569), .B(n568), .Z(n570) );
  AND U1172 ( .A(n571), .B(n570), .Z(n958) );
  XNOR U1173 ( .A(n958), .B(n956), .Z(n576) );
  XOR U1174 ( .A(n957), .B(n576), .Z(n899) );
  XNOR U1175 ( .A(n964), .B(n962), .Z(n589) );
  XOR U1176 ( .A(n963), .B(n589), .Z(n898) );
  XNOR U1177 ( .A(n898), .B(n897), .Z(n593) );
  XNOR U1178 ( .A(n899), .B(n593), .Z(n1005) );
  NANDN U1179 ( .A(n595), .B(n594), .Z(n599) );
  NAND U1180 ( .A(n597), .B(n596), .Z(n598) );
  NAND U1181 ( .A(n599), .B(n598), .Z(n1040) );
  NANDN U1182 ( .A(n601), .B(n600), .Z(n605) );
  NAND U1183 ( .A(n603), .B(n602), .Z(n604) );
  AND U1184 ( .A(n605), .B(n604), .Z(n1039) );
  XNOR U1185 ( .A(n1039), .B(oglobal[1]), .Z(n606) );
  XOR U1186 ( .A(n1040), .B(n606), .Z(n1014) );
  NANDN U1187 ( .A(n608), .B(n607), .Z(n612) );
  NANDN U1188 ( .A(n610), .B(n609), .Z(n611) );
  AND U1189 ( .A(n612), .B(n611), .Z(n967) );
  NANDN U1190 ( .A(n614), .B(n613), .Z(n618) );
  NAND U1191 ( .A(n616), .B(n615), .Z(n617) );
  NAND U1192 ( .A(n618), .B(n617), .Z(n966) );
  NANDN U1193 ( .A(n620), .B(n619), .Z(n624) );
  NANDN U1194 ( .A(n622), .B(n621), .Z(n623) );
  AND U1195 ( .A(n624), .B(n623), .Z(n965) );
  XOR U1196 ( .A(n966), .B(n965), .Z(n625) );
  XNOR U1197 ( .A(n967), .B(n625), .Z(n1012) );
  XOR U1198 ( .A(n1012), .B(n1013), .Z(n1015) );
  XNOR U1199 ( .A(n1014), .B(n1015), .Z(n1004) );
  XNOR U1200 ( .A(n1005), .B(n1004), .Z(n629) );
  XNOR U1201 ( .A(n1003), .B(n629), .Z(n1076) );
  XNOR U1202 ( .A(n630), .B(n1076), .Z(n631) );
  XOR U1203 ( .A(n1077), .B(n631), .Z(n1080) );
  NANDN U1204 ( .A(n633), .B(n632), .Z(n637) );
  NANDN U1205 ( .A(n635), .B(n634), .Z(n636) );
  AND U1206 ( .A(n637), .B(n636), .Z(n917) );
  XOR U1207 ( .A(n919), .B(n918), .Z(n646) );
  XOR U1208 ( .A(n917), .B(n646), .Z(n976) );
  XNOR U1209 ( .A(n978), .B(n977), .Z(n653) );
  XNOR U1210 ( .A(n976), .B(n653), .Z(n1093) );
  NANDN U1211 ( .A(n659), .B(n658), .Z(n663) );
  NANDN U1212 ( .A(n661), .B(n660), .Z(n662) );
  AND U1213 ( .A(n663), .B(n662), .Z(n936) );
  NANDN U1214 ( .A(n665), .B(n664), .Z(n669) );
  NANDN U1215 ( .A(n667), .B(n666), .Z(n668) );
  AND U1216 ( .A(n669), .B(n668), .Z(n935) );
  XNOR U1217 ( .A(n936), .B(n935), .Z(n670) );
  XOR U1218 ( .A(n934), .B(n670), .Z(n1051) );
  IV U1219 ( .A(n1051), .Z(n1052) );
  XNOR U1220 ( .A(n1055), .B(n1053), .Z(n677) );
  XNOR U1221 ( .A(n1052), .B(n677), .Z(n1092) );
  NANDN U1222 ( .A(n679), .B(n678), .Z(n683) );
  NANDN U1223 ( .A(n681), .B(n680), .Z(n682) );
  NAND U1224 ( .A(n683), .B(n682), .Z(n913) );
  NANDN U1225 ( .A(n685), .B(n684), .Z(n689) );
  NANDN U1226 ( .A(n687), .B(n686), .Z(n688) );
  NAND U1227 ( .A(n689), .B(n688), .Z(n912) );
  NANDN U1228 ( .A(n691), .B(n690), .Z(n695) );
  NANDN U1229 ( .A(n693), .B(n692), .Z(n694) );
  AND U1230 ( .A(n695), .B(n694), .Z(n911) );
  XOR U1231 ( .A(n912), .B(n911), .Z(n696) );
  XNOR U1232 ( .A(n913), .B(n696), .Z(n894) );
  XNOR U1233 ( .A(n896), .B(n895), .Z(n703) );
  XNOR U1234 ( .A(n894), .B(n703), .Z(n1091) );
  XNOR U1235 ( .A(n1092), .B(n1091), .Z(n704) );
  XNOR U1236 ( .A(n1093), .B(n704), .Z(n1084) );
  NANDN U1237 ( .A(n706), .B(n705), .Z(n710) );
  NANDN U1238 ( .A(n708), .B(n707), .Z(n709) );
  AND U1239 ( .A(n710), .B(n709), .Z(n1082) );
  NAND U1240 ( .A(n720), .B(n719), .Z(n725) );
  IV U1241 ( .A(n721), .Z(n723) );
  NAND U1242 ( .A(n723), .B(n722), .Z(n724) );
  AND U1243 ( .A(n725), .B(n724), .Z(n924) );
  XNOR U1244 ( .A(n928), .B(n924), .Z(n726) );
  XOR U1245 ( .A(n925), .B(n726), .Z(n906) );
  XNOR U1246 ( .A(n1033), .B(n1034), .Z(n1036) );
  NAND U1247 ( .A(n743), .B(n742), .Z(n748) );
  IV U1248 ( .A(n744), .Z(n746) );
  NAND U1249 ( .A(n746), .B(n745), .Z(n747) );
  AND U1250 ( .A(n748), .B(n747), .Z(n961) );
  XNOR U1251 ( .A(n961), .B(n960), .Z(n753) );
  XOR U1252 ( .A(n959), .B(n753), .Z(n1035) );
  XNOR U1253 ( .A(n1036), .B(n1035), .Z(n904) );
  IV U1254 ( .A(n904), .Z(n903) );
  XNOR U1255 ( .A(n905), .B(n903), .Z(n754) );
  XNOR U1256 ( .A(n906), .B(n754), .Z(n1088) );
  NANDN U1257 ( .A(n756), .B(n755), .Z(n761) );
  ANDN U1258 ( .B(n756), .A(n755), .Z(n759) );
  IV U1259 ( .A(n757), .Z(n758) );
  OR U1260 ( .A(n759), .B(n758), .Z(n760) );
  AND U1261 ( .A(n761), .B(n760), .Z(n1089) );
  XNOR U1262 ( .A(n1089), .B(n1090), .Z(n765) );
  XNOR U1263 ( .A(n1088), .B(n765), .Z(n1083) );
  XNOR U1264 ( .A(n1082), .B(n1083), .Z(n766) );
  XNOR U1265 ( .A(n1084), .B(n766), .Z(n1078) );
  XOR U1266 ( .A(n1078), .B(n1079), .Z(n770) );
  XNOR U1267 ( .A(n1080), .B(n770), .Z(n1103) );
  NANDN U1268 ( .A(n772), .B(n771), .Z(n776) );
  NANDN U1269 ( .A(n774), .B(n773), .Z(n775) );
  AND U1270 ( .A(n776), .B(n775), .Z(n990) );
  NANDN U1271 ( .A(n778), .B(n777), .Z(n782) );
  NANDN U1272 ( .A(n780), .B(n779), .Z(n781) );
  NAND U1273 ( .A(n782), .B(n781), .Z(n989) );
  NANDN U1274 ( .A(n784), .B(n783), .Z(n788) );
  NANDN U1275 ( .A(n786), .B(n785), .Z(n787) );
  AND U1276 ( .A(n788), .B(n787), .Z(n988) );
  XOR U1277 ( .A(n989), .B(n988), .Z(n789) );
  XNOR U1278 ( .A(n990), .B(n789), .Z(n1061) );
  NANDN U1279 ( .A(n791), .B(n790), .Z(n795) );
  NANDN U1280 ( .A(n793), .B(n792), .Z(n794) );
  AND U1281 ( .A(n795), .B(n794), .Z(n968) );
  NANDN U1282 ( .A(n797), .B(n796), .Z(n801) );
  NANDN U1283 ( .A(n799), .B(n798), .Z(n800) );
  AND U1284 ( .A(n801), .B(n800), .Z(n970) );
  NANDN U1285 ( .A(n803), .B(n802), .Z(n807) );
  NANDN U1286 ( .A(n805), .B(n804), .Z(n806) );
  NAND U1287 ( .A(n807), .B(n806), .Z(n969) );
  XOR U1288 ( .A(n970), .B(n969), .Z(n808) );
  XNOR U1289 ( .A(n968), .B(n808), .Z(n1060) );
  XNOR U1290 ( .A(n1060), .B(n1059), .Z(n812) );
  XNOR U1291 ( .A(n1061), .B(n812), .Z(n999) );
  XNOR U1292 ( .A(n1000), .B(n1001), .Z(n819) );
  XNOR U1293 ( .A(n999), .B(n819), .Z(n1087) );
  OR U1294 ( .A(n827), .B(n826), .Z(n831) );
  AND U1295 ( .A(n827), .B(n826), .Z(n828) );
  OR U1296 ( .A(n829), .B(n828), .Z(n830) );
  AND U1297 ( .A(n831), .B(n830), .Z(n1067) );
  XOR U1298 ( .A(n1067), .B(n1066), .Z(n835) );
  XOR U1299 ( .A(n1065), .B(n835), .Z(n981) );
  XNOR U1300 ( .A(n980), .B(n979), .Z(n982) );
  XNOR U1301 ( .A(n981), .B(n982), .Z(n1100) );
  XNOR U1302 ( .A(n1048), .B(n1046), .Z(n851) );
  XNOR U1303 ( .A(n1045), .B(n851), .Z(n1099) );
  NAND U1304 ( .A(n857), .B(n856), .Z(n861) );
  NAND U1305 ( .A(n859), .B(n858), .Z(n860) );
  NAND U1306 ( .A(n861), .B(n860), .Z(n972) );
  XOR U1307 ( .A(n972), .B(n971), .Z(n866) );
  XNOR U1308 ( .A(n973), .B(n866), .Z(n1028) );
  NANDN U1309 ( .A(n871), .B(n870), .Z(n875) );
  NANDN U1310 ( .A(n873), .B(n872), .Z(n874) );
  AND U1311 ( .A(n875), .B(n874), .Z(n987) );
  NANDN U1312 ( .A(n877), .B(n876), .Z(n881) );
  NANDN U1313 ( .A(n879), .B(n878), .Z(n880) );
  NAND U1314 ( .A(n881), .B(n880), .Z(n986) );
  XOR U1315 ( .A(n986), .B(n985), .Z(n886) );
  XOR U1316 ( .A(n987), .B(n886), .Z(n1025) );
  IV U1317 ( .A(n1025), .Z(n1027) );
  XNOR U1318 ( .A(n1026), .B(n1027), .Z(n887) );
  XNOR U1319 ( .A(n1028), .B(n887), .Z(n1098) );
  IV U1320 ( .A(n1098), .Z(n1097) );
  XNOR U1321 ( .A(n1099), .B(n1097), .Z(n888) );
  XNOR U1322 ( .A(n1100), .B(n888), .Z(n1085) );
  XNOR U1323 ( .A(n1086), .B(n1085), .Z(n889) );
  XNOR U1324 ( .A(n1087), .B(n889), .Z(n1105) );
  XNOR U1325 ( .A(n1105), .B(n1104), .Z(n893) );
  XNOR U1326 ( .A(n1103), .B(n893), .Z(o[1]) );
  NANDN U1327 ( .A(n898), .B(n897), .Z(n902) );
  ANDN U1328 ( .B(n898), .A(n897), .Z(n900) );
  OR U1329 ( .A(n900), .B(n899), .Z(n901) );
  AND U1330 ( .A(n902), .B(n901), .Z(n1109) );
  NANDN U1331 ( .A(n905), .B(n903), .Z(n909) );
  AND U1332 ( .A(n905), .B(n904), .Z(n907) );
  NANDN U1333 ( .A(n907), .B(n906), .Z(n908) );
  AND U1334 ( .A(n909), .B(n908), .Z(n1108) );
  XOR U1335 ( .A(n1109), .B(n1108), .Z(n910) );
  XNOR U1336 ( .A(n1107), .B(n910), .Z(n1173) );
  NANDN U1337 ( .A(n918), .B(n917), .Z(n922) );
  ANDN U1338 ( .B(n918), .A(n917), .Z(n920) );
  NANDN U1339 ( .A(n920), .B(n919), .Z(n921) );
  AND U1340 ( .A(n922), .B(n921), .Z(n1119) );
  XOR U1341 ( .A(n1120), .B(n1119), .Z(n923) );
  XNOR U1342 ( .A(n1118), .B(n923), .Z(n1190) );
  IV U1343 ( .A(n924), .Z(n926) );
  NAND U1344 ( .A(n926), .B(n925), .Z(n930) );
  NOR U1345 ( .A(n926), .B(n925), .Z(n927) );
  OR U1346 ( .A(n928), .B(n927), .Z(n929) );
  AND U1347 ( .A(n930), .B(n929), .Z(n1110) );
  XNOR U1348 ( .A(n1112), .B(n1111), .Z(n937) );
  XNOR U1349 ( .A(n1110), .B(n937), .Z(n1189) );
  XOR U1350 ( .A(n1134), .B(n1133), .Z(n947) );
  XNOR U1351 ( .A(n1132), .B(n947), .Z(n1188) );
  IV U1352 ( .A(n1188), .Z(n1187) );
  XNOR U1353 ( .A(n1189), .B(n1187), .Z(n948) );
  XNOR U1354 ( .A(n1190), .B(n948), .Z(n1172) );
  XOR U1355 ( .A(n1113), .B(oglobal[2]), .Z(n955) );
  XNOR U1356 ( .A(n1114), .B(n955), .Z(n1152) );
  XNOR U1357 ( .A(n1146), .B(n1145), .Z(n1147) );
  XNOR U1358 ( .A(n1148), .B(n1147), .Z(n1150) );
  XOR U1359 ( .A(n1144), .B(n1143), .Z(n974) );
  XNOR U1360 ( .A(n1142), .B(n974), .Z(n1149) );
  XOR U1361 ( .A(n1150), .B(n1149), .Z(n1151) );
  XNOR U1362 ( .A(n1152), .B(n1151), .Z(n1171) );
  IV U1363 ( .A(n1171), .Z(n1170) );
  XNOR U1364 ( .A(n1172), .B(n1170), .Z(n975) );
  XOR U1365 ( .A(n1173), .B(n975), .Z(n1210) );
  OR U1366 ( .A(n980), .B(n979), .Z(n984) );
  OR U1367 ( .A(n982), .B(n981), .Z(n983) );
  AND U1368 ( .A(n984), .B(n983), .Z(n1193) );
  XNOR U1369 ( .A(n1137), .B(n1136), .Z(n994) );
  XNOR U1370 ( .A(n1135), .B(n994), .Z(n1191) );
  XNOR U1371 ( .A(n1193), .B(n1191), .Z(n995) );
  XNOR U1372 ( .A(n1192), .B(n995), .Z(n1164) );
  IV U1373 ( .A(n1164), .Z(n1163) );
  XNOR U1374 ( .A(n1167), .B(n1165), .Z(n1002) );
  XNOR U1375 ( .A(n1163), .B(n1002), .Z(n1177) );
  NANDN U1376 ( .A(n1007), .B(n1006), .Z(n1011) );
  ANDN U1377 ( .B(n1007), .A(n1006), .Z(n1009) );
  OR U1378 ( .A(n1009), .B(n1008), .Z(n1010) );
  AND U1379 ( .A(n1011), .B(n1010), .Z(n1175) );
  XOR U1380 ( .A(n1176), .B(n1175), .Z(n1178) );
  XOR U1381 ( .A(n1177), .B(n1178), .Z(n1212) );
  NANDN U1382 ( .A(n1013), .B(n1012), .Z(n1017) );
  OR U1383 ( .A(n1015), .B(n1014), .Z(n1016) );
  AND U1384 ( .A(n1017), .B(n1016), .Z(n1156) );
  NAND U1385 ( .A(n1018), .B(n1019), .Z(n1024) );
  ANDN U1386 ( .B(n1020), .A(n1019), .Z(n1022) );
  OR U1387 ( .A(n1022), .B(n1021), .Z(n1023) );
  AND U1388 ( .A(n1024), .B(n1023), .Z(n1157) );
  NAND U1389 ( .A(n1025), .B(n1026), .Z(n1031) );
  ANDN U1390 ( .B(n1027), .A(n1026), .Z(n1029) );
  OR U1391 ( .A(n1029), .B(n1028), .Z(n1030) );
  AND U1392 ( .A(n1031), .B(n1030), .Z(n1155) );
  XNOR U1393 ( .A(n1157), .B(n1155), .Z(n1032) );
  XNOR U1394 ( .A(n1156), .B(n1032), .Z(n1183) );
  NANDN U1395 ( .A(n1034), .B(n1033), .Z(n1038) );
  NAND U1396 ( .A(n1036), .B(n1035), .Z(n1037) );
  NAND U1397 ( .A(n1038), .B(n1037), .Z(n1138) );
  XNOR U1398 ( .A(n1139), .B(n1140), .Z(n1044) );
  XOR U1399 ( .A(n1138), .B(n1044), .Z(n1128) );
  OR U1400 ( .A(n1046), .B(n1045), .Z(n1050) );
  AND U1401 ( .A(n1046), .B(n1045), .Z(n1047) );
  OR U1402 ( .A(n1048), .B(n1047), .Z(n1049) );
  AND U1403 ( .A(n1050), .B(n1049), .Z(n1130) );
  NANDN U1404 ( .A(n1053), .B(n1051), .Z(n1057) );
  AND U1405 ( .A(n1053), .B(n1052), .Z(n1054) );
  OR U1406 ( .A(n1055), .B(n1054), .Z(n1056) );
  AND U1407 ( .A(n1057), .B(n1056), .Z(n1129) );
  XNOR U1408 ( .A(n1130), .B(n1129), .Z(n1058) );
  XNOR U1409 ( .A(n1128), .B(n1058), .Z(n1181) );
  XNOR U1410 ( .A(n1195), .B(n1194), .Z(n1068) );
  XNOR U1411 ( .A(n1196), .B(n1068), .Z(n1124) );
  XNOR U1412 ( .A(n1123), .B(n1122), .Z(n1125) );
  XNOR U1413 ( .A(n1124), .B(n1125), .Z(n1182) );
  XOR U1414 ( .A(n1181), .B(n1182), .Z(n1184) );
  XNOR U1415 ( .A(n1183), .B(n1184), .Z(n1211) );
  XNOR U1416 ( .A(n1208), .B(n1207), .Z(n1081) );
  XOR U1417 ( .A(n1209), .B(n1081), .Z(n1217) );
  OR U1418 ( .A(n1092), .B(n1091), .Z(n1096) );
  AND U1419 ( .A(n1092), .B(n1091), .Z(n1094) );
  OR U1420 ( .A(n1094), .B(n1093), .Z(n1095) );
  AND U1421 ( .A(n1096), .B(n1095), .Z(n1162) );
  XOR U1422 ( .A(n1162), .B(n1161), .Z(n1101) );
  XNOR U1423 ( .A(n1160), .B(n1101), .Z(n1201) );
  IV U1424 ( .A(n1201), .Z(n1200) );
  XNOR U1425 ( .A(n1204), .B(n1200), .Z(n1102) );
  XNOR U1426 ( .A(n1202), .B(n1102), .Z(n1216) );
  IV U1427 ( .A(n1216), .Z(n1214) );
  XNOR U1428 ( .A(n1214), .B(n1215), .Z(n1106) );
  XNOR U1429 ( .A(n1217), .B(n1106), .Z(o[2]) );
  XOR U1430 ( .A(n1261), .B(oglobal[3]), .Z(n1254) );
  NANDN U1431 ( .A(n1113), .B(oglobal[2]), .Z(n1117) );
  ANDN U1432 ( .B(n1113), .A(oglobal[2]), .Z(n1115) );
  OR U1433 ( .A(n1115), .B(n1114), .Z(n1116) );
  AND U1434 ( .A(n1117), .B(n1116), .Z(n1252) );
  XNOR U1435 ( .A(n1252), .B(n1253), .Z(n1121) );
  XNOR U1436 ( .A(n1254), .B(n1121), .Z(n1222) );
  NAND U1437 ( .A(n1123), .B(n1122), .Z(n1127) );
  NANDN U1438 ( .A(n1125), .B(n1124), .Z(n1126) );
  AND U1439 ( .A(n1127), .B(n1126), .Z(n1224) );
  XNOR U1440 ( .A(n1224), .B(n1223), .Z(n1131) );
  XNOR U1441 ( .A(n1222), .B(n1131), .Z(n1242) );
  XOR U1442 ( .A(n1258), .B(n1255), .Z(n1141) );
  XOR U1443 ( .A(n1256), .B(n1141), .Z(n1247) );
  XNOR U1444 ( .A(n1246), .B(n1245), .Z(n1248) );
  XOR U1445 ( .A(n1247), .B(n1248), .Z(n1234) );
  NAND U1446 ( .A(n1150), .B(n1149), .Z(n1154) );
  NAND U1447 ( .A(n1152), .B(n1151), .Z(n1153) );
  AND U1448 ( .A(n1154), .B(n1153), .Z(n1232) );
  XNOR U1449 ( .A(n1232), .B(n1233), .Z(n1158) );
  XNOR U1450 ( .A(n1234), .B(n1158), .Z(n1239) );
  IV U1451 ( .A(n1239), .Z(n1238) );
  XNOR U1452 ( .A(n1242), .B(n1238), .Z(n1159) );
  XNOR U1453 ( .A(n1240), .B(n1159), .Z(n1274) );
  NANDN U1454 ( .A(n1165), .B(n1163), .Z(n1169) );
  AND U1455 ( .A(n1165), .B(n1164), .Z(n1166) );
  OR U1456 ( .A(n1167), .B(n1166), .Z(n1168) );
  AND U1457 ( .A(n1169), .B(n1168), .Z(n1228) );
  XOR U1458 ( .A(n1228), .B(n1226), .Z(n1174) );
  XNOR U1459 ( .A(n1225), .B(n1174), .Z(n1273) );
  OR U1460 ( .A(n1176), .B(n1175), .Z(n1180) );
  NAND U1461 ( .A(n1178), .B(n1177), .Z(n1179) );
  NAND U1462 ( .A(n1180), .B(n1179), .Z(n1268) );
  NAND U1463 ( .A(n1182), .B(n1181), .Z(n1186) );
  NAND U1464 ( .A(n1184), .B(n1183), .Z(n1185) );
  NAND U1465 ( .A(n1186), .B(n1185), .Z(n1266) );
  IV U1466 ( .A(n1266), .Z(n1265) );
  XNOR U1467 ( .A(n1250), .B(n1249), .Z(n1197) );
  XNOR U1468 ( .A(n1251), .B(n1197), .Z(n1267) );
  XNOR U1469 ( .A(n1265), .B(n1267), .Z(n1198) );
  XNOR U1470 ( .A(n1268), .B(n1198), .Z(n1272) );
  XOR U1471 ( .A(n1273), .B(n1272), .Z(n1199) );
  XNOR U1472 ( .A(n1274), .B(n1199), .Z(n1280) );
  NANDN U1473 ( .A(n1202), .B(n1200), .Z(n1206) );
  AND U1474 ( .A(n1202), .B(n1201), .Z(n1203) );
  OR U1475 ( .A(n1204), .B(n1203), .Z(n1205) );
  AND U1476 ( .A(n1206), .B(n1205), .Z(n1276) );
  XNOR U1477 ( .A(n1278), .B(n1277), .Z(n1213) );
  XNOR U1478 ( .A(n1276), .B(n1213), .Z(n1281) );
  NAND U1479 ( .A(n1214), .B(n1215), .Z(n1220) );
  ANDN U1480 ( .B(n1216), .A(n1215), .Z(n1218) );
  OR U1481 ( .A(n1218), .B(n1217), .Z(n1219) );
  AND U1482 ( .A(n1220), .B(n1219), .Z(n1279) );
  XNOR U1483 ( .A(n1281), .B(n1279), .Z(n1221) );
  XNOR U1484 ( .A(n1280), .B(n1221), .Z(o[3]) );
  OR U1485 ( .A(n1226), .B(n1225), .Z(n1230) );
  AND U1486 ( .A(n1226), .B(n1225), .Z(n1227) );
  OR U1487 ( .A(n1228), .B(n1227), .Z(n1229) );
  AND U1488 ( .A(n1230), .B(n1229), .Z(n1294) );
  IV U1489 ( .A(n1232), .Z(n1231) );
  NANDN U1490 ( .A(n1233), .B(n1231), .Z(n1237) );
  AND U1491 ( .A(n1233), .B(n1232), .Z(n1235) );
  OR U1492 ( .A(n1235), .B(n1234), .Z(n1236) );
  AND U1493 ( .A(n1237), .B(n1236), .Z(n1293) );
  XNOR U1494 ( .A(n1294), .B(n1293), .Z(n1295) );
  XOR U1495 ( .A(n1296), .B(n1295), .Z(n1307) );
  NANDN U1496 ( .A(n1240), .B(n1238), .Z(n1244) );
  AND U1497 ( .A(n1240), .B(n1239), .Z(n1241) );
  OR U1498 ( .A(n1242), .B(n1241), .Z(n1243) );
  AND U1499 ( .A(n1244), .B(n1243), .Z(n1306) );
  NANDN U1500 ( .A(n1256), .B(n1255), .Z(n1260) );
  ANDN U1501 ( .B(n1256), .A(n1255), .Z(n1257) );
  OR U1502 ( .A(n1258), .B(n1257), .Z(n1259) );
  AND U1503 ( .A(n1260), .B(n1259), .Z(n1303) );
  ANDN U1504 ( .B(oglobal[3]), .A(n1261), .Z(n1297) );
  XOR U1505 ( .A(n1297), .B(oglobal[4]), .Z(n1301) );
  XNOR U1506 ( .A(n1303), .B(n1301), .Z(n1262) );
  XNOR U1507 ( .A(n1302), .B(n1262), .Z(n1298) );
  XNOR U1508 ( .A(n1300), .B(n1298), .Z(n1263) );
  XOR U1509 ( .A(n1299), .B(n1263), .Z(n1305) );
  XNOR U1510 ( .A(n1306), .B(n1305), .Z(n1264) );
  XNOR U1511 ( .A(n1307), .B(n1264), .Z(n1292) );
  NANDN U1512 ( .A(n1267), .B(n1265), .Z(n1271) );
  AND U1513 ( .A(n1267), .B(n1266), .Z(n1269) );
  OR U1514 ( .A(n1269), .B(n1268), .Z(n1270) );
  AND U1515 ( .A(n1271), .B(n1270), .Z(n1291) );
  XNOR U1516 ( .A(n1291), .B(n1290), .Z(n1275) );
  XNOR U1517 ( .A(n1292), .B(n1275), .Z(n1284) );
  IV U1518 ( .A(n1284), .Z(n1283) );
  XNOR U1519 ( .A(n1287), .B(n1285), .Z(n1282) );
  XNOR U1520 ( .A(n1283), .B(n1282), .Z(o[4]) );
  NANDN U1521 ( .A(n1285), .B(n1283), .Z(n1289) );
  AND U1522 ( .A(n1285), .B(n1284), .Z(n1286) );
  OR U1523 ( .A(n1287), .B(n1286), .Z(n1288) );
  AND U1524 ( .A(n1289), .B(n1288), .Z(n1318) );
  AND U1525 ( .A(n1297), .B(oglobal[4]), .Z(n1310) );
  XOR U1526 ( .A(n1310), .B(oglobal[5]), .Z(n1312) );
  XNOR U1527 ( .A(n1313), .B(n1311), .Z(n1304) );
  XOR U1528 ( .A(n1312), .B(n1304), .Z(n1315) );
  XOR U1529 ( .A(n1315), .B(n1316), .Z(n1308) );
  XNOR U1530 ( .A(n1314), .B(n1308), .Z(n1317) );
  XNOR U1531 ( .A(n1319), .B(n1317), .Z(n1309) );
  XNOR U1532 ( .A(n1318), .B(n1309), .Z(o[5]) );
  AND U1533 ( .A(n1310), .B(oglobal[5]), .Z(n1324) );
  XOR U1534 ( .A(oglobal[6]), .B(n1324), .Z(n1326) );
  XNOR U1535 ( .A(n1326), .B(n1325), .Z(n1323) );
  XOR U1536 ( .A(n1322), .B(n1321), .Z(n1320) );
  XNOR U1537 ( .A(n1323), .B(n1320), .Z(o[6]) );
  NAND U1538 ( .A(n1324), .B(oglobal[6]), .Z(n1328) );
  NAND U1539 ( .A(n1326), .B(n1325), .Z(n1327) );
  AND U1540 ( .A(n1328), .B(n1327), .Z(n1330) );
  XNOR U1541 ( .A(n1331), .B(n1330), .Z(n1329) );
  XNOR U1542 ( .A(oglobal[7]), .B(n1329), .Z(o[7]) );
  XNOR U1543 ( .A(n1332), .B(oglobal[8]), .Z(o[8]) );
  NANDN U1544 ( .A(n1332), .B(oglobal[8]), .Z(n1333) );
  XNOR U1545 ( .A(oglobal[9]), .B(n1333), .Z(o[9]) );
  NANDN U1546 ( .A(n1333), .B(oglobal[9]), .Z(n1334) );
  XNOR U1547 ( .A(oglobal[10]), .B(n1334), .Z(o[10]) );
endmodule

