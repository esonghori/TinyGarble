
module hamming_N1600_CC8 ( clk, rst, x, y, o );
  input [199:0] x;
  input [199:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NANDN U203 ( .A(n516), .B(n515), .Z(n1) );
  NANDN U204 ( .A(n514), .B(n513), .Z(n2) );
  AND U205 ( .A(n1), .B(n2), .Z(n859) );
  NANDN U206 ( .A(n746), .B(n745), .Z(n3) );
  NANDN U207 ( .A(n744), .B(n743), .Z(n4) );
  AND U208 ( .A(n3), .B(n4), .Z(n880) );
  NANDN U209 ( .A(n723), .B(n722), .Z(n5) );
  NANDN U210 ( .A(n721), .B(n720), .Z(n6) );
  NAND U211 ( .A(n5), .B(n6), .Z(n875) );
  NANDN U212 ( .A(n372), .B(n371), .Z(n7) );
  NANDN U213 ( .A(n370), .B(n369), .Z(n8) );
  NAND U214 ( .A(n7), .B(n8), .Z(n907) );
  NANDN U215 ( .A(n619), .B(n618), .Z(n9) );
  NANDN U216 ( .A(n617), .B(n616), .Z(n10) );
  AND U217 ( .A(n9), .B(n10), .Z(n980) );
  XOR U218 ( .A(n292), .B(n291), .Z(n11) );
  NANDN U219 ( .A(n290), .B(n11), .Z(n12) );
  NAND U220 ( .A(n292), .B(n291), .Z(n13) );
  AND U221 ( .A(n12), .B(n13), .Z(n931) );
  XOR U222 ( .A(n857), .B(n856), .Z(n14) );
  NANDN U223 ( .A(n858), .B(n14), .Z(n15) );
  NAND U224 ( .A(n857), .B(n856), .Z(n16) );
  AND U225 ( .A(n15), .B(n16), .Z(n1046) );
  NANDN U226 ( .A(n659), .B(n658), .Z(n17) );
  NANDN U227 ( .A(n657), .B(n656), .Z(n18) );
  NAND U228 ( .A(n17), .B(n18), .Z(n870) );
  NANDN U229 ( .A(n491), .B(n490), .Z(n19) );
  NANDN U230 ( .A(n489), .B(n488), .Z(n20) );
  AND U231 ( .A(n19), .B(n20), .Z(n863) );
  NAND U232 ( .A(n590), .B(n589), .Z(n21) );
  NANDN U233 ( .A(n588), .B(n587), .Z(n22) );
  NAND U234 ( .A(n21), .B(n22), .Z(n829) );
  NANDN U235 ( .A(n687), .B(n686), .Z(n23) );
  NANDN U236 ( .A(n685), .B(n684), .Z(n24) );
  NAND U237 ( .A(n23), .B(n24), .Z(n858) );
  NANDN U238 ( .A(n672), .B(n671), .Z(n25) );
  NANDN U239 ( .A(n670), .B(n669), .Z(n26) );
  NAND U240 ( .A(n25), .B(n26), .Z(n883) );
  NANDN U241 ( .A(n738), .B(n737), .Z(n27) );
  NANDN U242 ( .A(n736), .B(n735), .Z(n28) );
  NAND U243 ( .A(n27), .B(n28), .Z(n881) );
  NANDN U244 ( .A(n731), .B(n730), .Z(n29) );
  NANDN U245 ( .A(n729), .B(n728), .Z(n30) );
  NAND U246 ( .A(n29), .B(n30), .Z(n876) );
  NANDN U247 ( .A(n376), .B(n375), .Z(n31) );
  NANDN U248 ( .A(n374), .B(n373), .Z(n32) );
  AND U249 ( .A(n31), .B(n32), .Z(n906) );
  NANDN U250 ( .A(n627), .B(n626), .Z(n33) );
  NANDN U251 ( .A(n625), .B(n624), .Z(n34) );
  NAND U252 ( .A(n33), .B(n34), .Z(n972) );
  NANDN U253 ( .A(n615), .B(n614), .Z(n35) );
  NANDN U254 ( .A(n613), .B(n612), .Z(n36) );
  NAND U255 ( .A(n35), .B(n36), .Z(n981) );
  NANDN U256 ( .A(n361), .B(n360), .Z(n37) );
  NANDN U257 ( .A(n359), .B(n358), .Z(n38) );
  AND U258 ( .A(n37), .B(n38), .Z(n819) );
  NANDN U259 ( .A(n646), .B(n645), .Z(n39) );
  NANDN U260 ( .A(n644), .B(n643), .Z(n40) );
  AND U261 ( .A(n39), .B(n40), .Z(n817) );
  XNOR U262 ( .A(n932), .B(n931), .Z(n933) );
  NAND U263 ( .A(n322), .B(n321), .Z(n41) );
  XOR U264 ( .A(n321), .B(n322), .Z(n42) );
  NANDN U265 ( .A(n320), .B(n42), .Z(n43) );
  NAND U266 ( .A(n41), .B(n43), .Z(n997) );
  NAND U267 ( .A(n912), .B(n911), .Z(n44) );
  XOR U268 ( .A(n911), .B(n912), .Z(n45) );
  NANDN U269 ( .A(n910), .B(n45), .Z(n46) );
  NAND U270 ( .A(n44), .B(n46), .Z(n1111) );
  NAND U271 ( .A(n873), .B(n872), .Z(n47) );
  XOR U272 ( .A(n872), .B(n873), .Z(n48) );
  NANDN U273 ( .A(n871), .B(n48), .Z(n49) );
  NAND U274 ( .A(n47), .B(n49), .Z(n1052) );
  NAND U275 ( .A(n861), .B(n860), .Z(n50) );
  XOR U276 ( .A(n860), .B(n861), .Z(n51) );
  NAND U277 ( .A(n51), .B(n859), .Z(n52) );
  NAND U278 ( .A(n50), .B(n52), .Z(n1045) );
  NAND U279 ( .A(n1109), .B(n1108), .Z(n53) );
  XOR U280 ( .A(n1108), .B(n1109), .Z(n54) );
  NAND U281 ( .A(n54), .B(n1107), .Z(n55) );
  NAND U282 ( .A(n53), .B(n55), .Z(n1168) );
  NAND U283 ( .A(n497), .B(n496), .Z(n56) );
  XOR U284 ( .A(n496), .B(n497), .Z(n57) );
  NANDN U285 ( .A(n495), .B(n57), .Z(n58) );
  NAND U286 ( .A(n56), .B(n58), .Z(n964) );
  NANDN U287 ( .A(n435), .B(n434), .Z(n59) );
  NANDN U288 ( .A(n433), .B(n432), .Z(n60) );
  AND U289 ( .A(n59), .B(n60), .Z(n871) );
  NANDN U290 ( .A(n487), .B(n486), .Z(n61) );
  NANDN U291 ( .A(n485), .B(n484), .Z(n62) );
  NAND U292 ( .A(n61), .B(n62), .Z(n862) );
  NANDN U293 ( .A(n471), .B(n470), .Z(n63) );
  NANDN U294 ( .A(n469), .B(n468), .Z(n64) );
  NAND U295 ( .A(n63), .B(n64), .Z(n853) );
  NANDN U296 ( .A(n623), .B(n622), .Z(n65) );
  NANDN U297 ( .A(n621), .B(n620), .Z(n66) );
  AND U298 ( .A(n65), .B(n66), .Z(n982) );
  NANDN U299 ( .A(n357), .B(n356), .Z(n67) );
  NANDN U300 ( .A(n355), .B(n354), .Z(n68) );
  NAND U301 ( .A(n67), .B(n68), .Z(n820) );
  NANDN U302 ( .A(n650), .B(n649), .Z(n69) );
  NANDN U303 ( .A(n648), .B(n647), .Z(n70) );
  AND U304 ( .A(n69), .B(n70), .Z(n816) );
  NANDN U305 ( .A(n557), .B(n556), .Z(n71) );
  NANDN U306 ( .A(n555), .B(n554), .Z(n72) );
  AND U307 ( .A(n71), .B(n72), .Z(n798) );
  NAND U308 ( .A(n352), .B(n351), .Z(n73) );
  XOR U309 ( .A(n351), .B(n352), .Z(n74) );
  NANDN U310 ( .A(n353), .B(n74), .Z(n75) );
  NAND U311 ( .A(n73), .B(n75), .Z(n985) );
  NAND U312 ( .A(n870), .B(n869), .Z(n76) );
  XOR U313 ( .A(n869), .B(n870), .Z(n77) );
  NANDN U314 ( .A(n868), .B(n77), .Z(n78) );
  NAND U315 ( .A(n76), .B(n78), .Z(n1051) );
  NAND U316 ( .A(n831), .B(n829), .Z(n79) );
  XOR U317 ( .A(n829), .B(n831), .Z(n80) );
  NAND U318 ( .A(n80), .B(n830), .Z(n81) );
  NAND U319 ( .A(n79), .B(n81), .Z(n1057) );
  XNOR U320 ( .A(n1046), .B(n1045), .Z(n1047) );
  NAND U321 ( .A(n909), .B(n908), .Z(n82) );
  NANDN U322 ( .A(n907), .B(n906), .Z(n83) );
  AND U323 ( .A(n82), .B(n83), .Z(n1086) );
  XOR U324 ( .A(oglobal[1]), .B(n972), .Z(n84) );
  NANDN U325 ( .A(n973), .B(n84), .Z(n85) );
  NAND U326 ( .A(oglobal[1]), .B(n972), .Z(n86) );
  AND U327 ( .A(n85), .B(n86), .Z(n1080) );
  OR U328 ( .A(n806), .B(n807), .Z(n87) );
  NANDN U329 ( .A(n809), .B(n808), .Z(n88) );
  AND U330 ( .A(n87), .B(n88), .Z(n1094) );
  NAND U331 ( .A(n894), .B(n893), .Z(n89) );
  NANDN U332 ( .A(n896), .B(n895), .Z(n90) );
  AND U333 ( .A(n89), .B(n90), .Z(n1023) );
  NAND U334 ( .A(n400), .B(n399), .Z(n91) );
  NAND U335 ( .A(n398), .B(n397), .Z(n92) );
  NAND U336 ( .A(n91), .B(n92), .Z(n785) );
  XOR U337 ( .A(n999), .B(n997), .Z(n93) );
  NANDN U338 ( .A(n998), .B(n93), .Z(n94) );
  NAND U339 ( .A(n999), .B(n997), .Z(n95) );
  AND U340 ( .A(n94), .B(n95), .Z(n1103) );
  NAND U341 ( .A(n1092), .B(n1091), .Z(n96) );
  NANDN U342 ( .A(n1090), .B(n1089), .Z(n97) );
  AND U343 ( .A(n96), .B(n97), .Z(n1149) );
  NAND U344 ( .A(n1033), .B(n1032), .Z(n98) );
  XOR U345 ( .A(n1032), .B(n1033), .Z(n99) );
  NANDN U346 ( .A(n1034), .B(n99), .Z(n100) );
  NAND U347 ( .A(n98), .B(n100), .Z(n1140) );
  NAND U348 ( .A(n1037), .B(n1036), .Z(n101) );
  XOR U349 ( .A(n1036), .B(n1037), .Z(n102) );
  NANDN U350 ( .A(n1038), .B(n102), .Z(n103) );
  NAND U351 ( .A(n101), .B(n103), .Z(n1185) );
  XOR U352 ( .A(n1134), .B(n1132), .Z(n104) );
  NAND U353 ( .A(n104), .B(n1133), .Z(n105) );
  NAND U354 ( .A(n1134), .B(n1132), .Z(n106) );
  AND U355 ( .A(n105), .B(n106), .Z(n1137) );
  XOR U356 ( .A(n734), .B(n732), .Z(n107) );
  NANDN U357 ( .A(n733), .B(n107), .Z(n108) );
  NAND U358 ( .A(n734), .B(n732), .Z(n109) );
  AND U359 ( .A(n108), .B(n109), .Z(n952) );
  NAND U360 ( .A(n402), .B(n401), .Z(n110) );
  XOR U361 ( .A(n401), .B(n402), .Z(n111) );
  NANDN U362 ( .A(n403), .B(n111), .Z(n112) );
  NAND U363 ( .A(n110), .B(n112), .Z(n833) );
  NANDN U364 ( .A(n439), .B(n438), .Z(n113) );
  NANDN U365 ( .A(n437), .B(n436), .Z(n114) );
  NAND U366 ( .A(n113), .B(n114), .Z(n873) );
  NANDN U367 ( .A(n663), .B(n662), .Z(n115) );
  NANDN U368 ( .A(n661), .B(n660), .Z(n116) );
  NAND U369 ( .A(n115), .B(n116), .Z(n869) );
  NANDN U370 ( .A(n508), .B(n507), .Z(n117) );
  NANDN U371 ( .A(n506), .B(n505), .Z(n118) );
  AND U372 ( .A(n117), .B(n118), .Z(n861) );
  NANDN U373 ( .A(n668), .B(n667), .Z(n119) );
  NANDN U374 ( .A(n666), .B(n665), .Z(n120) );
  NAND U375 ( .A(n119), .B(n120), .Z(n884) );
  NANDN U376 ( .A(n742), .B(n741), .Z(n121) );
  NANDN U377 ( .A(n740), .B(n739), .Z(n122) );
  AND U378 ( .A(n121), .B(n122), .Z(n882) );
  NANDN U379 ( .A(n380), .B(n379), .Z(n123) );
  NANDN U380 ( .A(n378), .B(n377), .Z(n124) );
  AND U381 ( .A(n123), .B(n124), .Z(n908) );
  NANDN U382 ( .A(n631), .B(n630), .Z(n125) );
  NANDN U383 ( .A(n629), .B(n628), .Z(n126) );
  AND U384 ( .A(n125), .B(n126), .Z(n973) );
  NANDN U385 ( .A(n642), .B(n641), .Z(n127) );
  NANDN U386 ( .A(n640), .B(n639), .Z(n128) );
  NAND U387 ( .A(n127), .B(n128), .Z(n818) );
  XOR U388 ( .A(n503), .B(n502), .Z(n129) );
  NANDN U389 ( .A(n504), .B(n129), .Z(n130) );
  NAND U390 ( .A(n503), .B(n502), .Z(n131) );
  AND U391 ( .A(n130), .B(n131), .Z(n894) );
  NAND U392 ( .A(n455), .B(n453), .Z(n132) );
  XOR U393 ( .A(n453), .B(n455), .Z(n133) );
  NANDN U394 ( .A(n454), .B(n133), .Z(n134) );
  NAND U395 ( .A(n132), .B(n134), .Z(n841) );
  NAND U396 ( .A(n904), .B(n903), .Z(n135) );
  XOR U397 ( .A(n903), .B(n904), .Z(n136) );
  NANDN U398 ( .A(n905), .B(n136), .Z(n137) );
  NAND U399 ( .A(n135), .B(n137), .Z(n1085) );
  NAND U400 ( .A(n822), .B(n821), .Z(n138) );
  NANDN U401 ( .A(n820), .B(n819), .Z(n139) );
  AND U402 ( .A(n138), .B(n139), .Z(n1098) );
  NANDN U403 ( .A(n892), .B(n891), .Z(n140) );
  NANDN U404 ( .A(n890), .B(n889), .Z(n141) );
  AND U405 ( .A(n140), .B(n141), .Z(n1022) );
  NAND U406 ( .A(n1062), .B(n1063), .Z(n142) );
  XOR U407 ( .A(n1063), .B(n1062), .Z(n143) );
  NANDN U408 ( .A(n1064), .B(n143), .Z(n144) );
  NAND U409 ( .A(n142), .B(n144), .Z(n1172) );
  XOR U410 ( .A(n1105), .B(n1103), .Z(n145) );
  NANDN U411 ( .A(n1104), .B(n145), .Z(n146) );
  NAND U412 ( .A(n1105), .B(n1103), .Z(n147) );
  AND U413 ( .A(n146), .B(n147), .Z(n1166) );
  NAND U414 ( .A(oglobal[2]), .B(n1057), .Z(n148) );
  XOR U415 ( .A(n1057), .B(oglobal[2]), .Z(n149) );
  NAND U416 ( .A(n149), .B(n1058), .Z(n150) );
  NAND U417 ( .A(n148), .B(n150), .Z(n1156) );
  NANDN U418 ( .A(n1094), .B(n1093), .Z(n151) );
  NANDN U419 ( .A(n1096), .B(n1095), .Z(n152) );
  NAND U420 ( .A(n151), .B(n152), .Z(n1143) );
  NAND U421 ( .A(n1031), .B(n1030), .Z(n153) );
  NAND U422 ( .A(n1028), .B(n1029), .Z(n154) );
  NAND U423 ( .A(n153), .B(n154), .Z(n1141) );
  NAND U424 ( .A(n395), .B(n396), .Z(n155) );
  NANDN U425 ( .A(n394), .B(n393), .Z(n156) );
  NAND U426 ( .A(n155), .B(n156), .Z(n765) );
  XOR U427 ( .A(n1168), .B(n1169), .Z(n157) );
  NANDN U428 ( .A(n1170), .B(n157), .Z(n158) );
  NAND U429 ( .A(n1168), .B(n1169), .Z(n159) );
  AND U430 ( .A(n158), .B(n159), .Z(n1223) );
  NAND U431 ( .A(n1009), .B(n1007), .Z(n160) );
  XOR U432 ( .A(n1007), .B(n1009), .Z(n161) );
  NAND U433 ( .A(n161), .B(n1008), .Z(n162) );
  NAND U434 ( .A(n160), .B(n162), .Z(n1122) );
  NAND U435 ( .A(n1129), .B(n1128), .Z(n163) );
  NANDN U436 ( .A(n1131), .B(n1130), .Z(n164) );
  AND U437 ( .A(n163), .B(n164), .Z(n1136) );
  NAND U438 ( .A(n560), .B(n559), .Z(n165) );
  XOR U439 ( .A(n559), .B(n560), .Z(n166) );
  NANDN U440 ( .A(n558), .B(n166), .Z(n167) );
  NAND U441 ( .A(n165), .B(n167), .Z(n844) );
  NANDN U442 ( .A(n443), .B(n442), .Z(n168) );
  NANDN U443 ( .A(n441), .B(n440), .Z(n169) );
  NAND U444 ( .A(n168), .B(n169), .Z(n872) );
  NANDN U445 ( .A(n655), .B(n654), .Z(n170) );
  NANDN U446 ( .A(n653), .B(n652), .Z(n171) );
  AND U447 ( .A(n170), .B(n171), .Z(n868) );
  NANDN U448 ( .A(n483), .B(n482), .Z(n172) );
  NANDN U449 ( .A(n481), .B(n480), .Z(n173) );
  NAND U450 ( .A(n172), .B(n173), .Z(n865) );
  NANDN U451 ( .A(n594), .B(n593), .Z(n174) );
  NANDN U452 ( .A(n592), .B(n591), .Z(n175) );
  NAND U453 ( .A(n174), .B(n175), .Z(n830) );
  NANDN U454 ( .A(n611), .B(n610), .Z(n176) );
  NANDN U455 ( .A(n609), .B(n608), .Z(n177) );
  AND U456 ( .A(n176), .B(n177), .Z(n826) );
  NANDN U457 ( .A(n696), .B(n695), .Z(n178) );
  NANDN U458 ( .A(n694), .B(n693), .Z(n179) );
  AND U459 ( .A(n178), .B(n179), .Z(n856) );
  NANDN U460 ( .A(n512), .B(n511), .Z(n180) );
  NANDN U461 ( .A(n510), .B(n509), .Z(n181) );
  AND U462 ( .A(n180), .B(n181), .Z(n860) );
  NANDN U463 ( .A(n676), .B(n675), .Z(n182) );
  NANDN U464 ( .A(n674), .B(n673), .Z(n183) );
  NAND U465 ( .A(n182), .B(n183), .Z(n885) );
  NANDN U466 ( .A(n727), .B(n726), .Z(n184) );
  NANDN U467 ( .A(n725), .B(n724), .Z(n185) );
  NAND U468 ( .A(n184), .B(n185), .Z(n874) );
  NANDN U469 ( .A(n365), .B(n364), .Z(n186) );
  NANDN U470 ( .A(n363), .B(n362), .Z(n187) );
  AND U471 ( .A(n186), .B(n187), .Z(n821) );
  NANDN U472 ( .A(n413), .B(n412), .Z(n188) );
  NANDN U473 ( .A(n411), .B(n410), .Z(n189) );
  AND U474 ( .A(n188), .B(n189), .Z(n806) );
  NANDN U475 ( .A(n547), .B(n546), .Z(n190) );
  NANDN U476 ( .A(n545), .B(n544), .Z(n191) );
  AND U477 ( .A(n190), .B(n191), .Z(n799) );
  XOR U478 ( .A(n501), .B(n500), .Z(n192) );
  NANDN U479 ( .A(n499), .B(n192), .Z(n193) );
  NAND U480 ( .A(n501), .B(n500), .Z(n194) );
  AND U481 ( .A(n193), .B(n194), .Z(n893) );
  NAND U482 ( .A(n294), .B(n293), .Z(n195) );
  XOR U483 ( .A(n293), .B(n294), .Z(n196) );
  NANDN U484 ( .A(n295), .B(n196), .Z(n197) );
  NAND U485 ( .A(n195), .B(n197), .Z(n889) );
  NAND U486 ( .A(n368), .B(n367), .Z(n198) );
  XOR U487 ( .A(n367), .B(n368), .Z(n199) );
  NAND U488 ( .A(n199), .B(n366), .Z(n200) );
  NAND U489 ( .A(n198), .B(n200), .Z(n937) );
  XOR U490 ( .A(n350), .B(n349), .Z(n201) );
  NANDN U491 ( .A(n348), .B(n201), .Z(n202) );
  NAND U492 ( .A(n350), .B(n349), .Z(n203) );
  AND U493 ( .A(n202), .B(n203), .Z(n984) );
  XOR U494 ( .A(n494), .B(n493), .Z(n204) );
  NANDN U495 ( .A(n492), .B(n204), .Z(n205) );
  NAND U496 ( .A(n494), .B(n493), .Z(n206) );
  AND U497 ( .A(n205), .B(n206), .Z(n968) );
  XOR U498 ( .A(n700), .B(n699), .Z(n207) );
  NANDN U499 ( .A(n698), .B(n207), .Z(n208) );
  NAND U500 ( .A(n700), .B(n699), .Z(n209) );
  AND U501 ( .A(n208), .B(n209), .Z(n992) );
  NAND U502 ( .A(n915), .B(n916), .Z(n210) );
  NANDN U503 ( .A(n914), .B(n913), .Z(n211) );
  NAND U504 ( .A(n210), .B(n211), .Z(n1110) );
  NAND U505 ( .A(n841), .B(n840), .Z(n212) );
  XOR U506 ( .A(n840), .B(n841), .Z(n213) );
  NANDN U507 ( .A(n839), .B(n213), .Z(n214) );
  NAND U508 ( .A(n212), .B(n214), .Z(n1068) );
  NAND U509 ( .A(n882), .B(n880), .Z(n215) );
  XOR U510 ( .A(n880), .B(n882), .Z(n216) );
  NANDN U511 ( .A(n881), .B(n216), .Z(n217) );
  NAND U512 ( .A(n215), .B(n217), .Z(n1089) );
  NAND U513 ( .A(n983), .B(n982), .Z(n218) );
  NANDN U514 ( .A(n981), .B(n980), .Z(n219) );
  NAND U515 ( .A(n218), .B(n219), .Z(n1081) );
  NAND U516 ( .A(n817), .B(n816), .Z(n220) );
  XOR U517 ( .A(n816), .B(n817), .Z(n221) );
  NANDN U518 ( .A(n818), .B(n221), .Z(n222) );
  NAND U519 ( .A(n220), .B(n222), .Z(n1097) );
  NAND U520 ( .A(n805), .B(n803), .Z(n223) );
  XOR U521 ( .A(n803), .B(n805), .Z(n224) );
  NANDN U522 ( .A(n804), .B(n224), .Z(n225) );
  NAND U523 ( .A(n223), .B(n225), .Z(n1093) );
  NAND U524 ( .A(n383), .B(n384), .Z(n226) );
  NANDN U525 ( .A(n382), .B(n381), .Z(n227) );
  NAND U526 ( .A(n226), .B(n227), .Z(n912) );
  XOR U527 ( .A(n1061), .B(n1060), .Z(n228) );
  NANDN U528 ( .A(n1059), .B(n228), .Z(n229) );
  NAND U529 ( .A(n1061), .B(n1060), .Z(n230) );
  AND U530 ( .A(n229), .B(n230), .Z(n1171) );
  NAND U531 ( .A(n1119), .B(n1118), .Z(n231) );
  NAND U532 ( .A(n1116), .B(n1117), .Z(n232) );
  AND U533 ( .A(n231), .B(n232), .Z(n1169) );
  NAND U534 ( .A(n1088), .B(n1087), .Z(n233) );
  NANDN U535 ( .A(n1086), .B(n1085), .Z(n234) );
  AND U536 ( .A(n233), .B(n234), .Z(n1150) );
  NAND U537 ( .A(n520), .B(n519), .Z(n235) );
  XOR U538 ( .A(n519), .B(n520), .Z(n236) );
  NANDN U539 ( .A(n518), .B(n236), .Z(n237) );
  NAND U540 ( .A(n235), .B(n237), .Z(n759) );
  XOR U541 ( .A(n1165), .B(n1166), .Z(n238) );
  NANDN U542 ( .A(n1167), .B(n238), .Z(n239) );
  NAND U543 ( .A(n1165), .B(n1166), .Z(n240) );
  AND U544 ( .A(n239), .B(n240), .Z(n1221) );
  NANDN U545 ( .A(n1158), .B(n1157), .Z(n241) );
  NANDN U546 ( .A(n1156), .B(n1155), .Z(n242) );
  AND U547 ( .A(n241), .B(n242), .Z(n1208) );
  XOR U548 ( .A(n1139), .B(n1140), .Z(n243) );
  NANDN U549 ( .A(n1141), .B(n243), .Z(n244) );
  NAND U550 ( .A(n1139), .B(n1140), .Z(n245) );
  AND U551 ( .A(n244), .B(n245), .Z(n1202) );
  NAND U552 ( .A(n523), .B(n522), .Z(n246) );
  XOR U553 ( .A(n522), .B(n523), .Z(n247) );
  NANDN U554 ( .A(n524), .B(n247), .Z(n248) );
  NAND U555 ( .A(n246), .B(n248), .Z(n1007) );
  NAND U556 ( .A(n1200), .B(n1198), .Z(n249) );
  XOR U557 ( .A(n1198), .B(n1200), .Z(n250) );
  NANDN U558 ( .A(n1199), .B(n250), .Z(n251) );
  NAND U559 ( .A(n249), .B(n251), .Z(n1241) );
  XOR U560 ( .A(n1138), .B(n1137), .Z(n252) );
  NAND U561 ( .A(n252), .B(n1136), .Z(n253) );
  NAND U562 ( .A(n1138), .B(n1137), .Z(n254) );
  AND U563 ( .A(n253), .B(n254), .Z(n1228) );
  XNOR U564 ( .A(x[118]), .B(y[118]), .Z(n423) );
  XNOR U565 ( .A(x[120]), .B(y[120]), .Z(n421) );
  XNOR U566 ( .A(x[122]), .B(y[122]), .Z(n420) );
  XNOR U567 ( .A(n421), .B(n420), .Z(n422) );
  XNOR U568 ( .A(n423), .B(n422), .Z(n286) );
  XNOR U569 ( .A(x[197]), .B(y[197]), .Z(n710) );
  XNOR U570 ( .A(x[2]), .B(y[2]), .Z(n708) );
  XNOR U571 ( .A(x[199]), .B(y[199]), .Z(n707) );
  XNOR U572 ( .A(n708), .B(n707), .Z(n709) );
  XNOR U573 ( .A(n710), .B(n709), .Z(n284) );
  XNOR U574 ( .A(x[112]), .B(y[112]), .Z(n576) );
  XNOR U575 ( .A(x[114]), .B(y[114]), .Z(n574) );
  XNOR U576 ( .A(x[116]), .B(y[116]), .Z(n573) );
  XNOR U577 ( .A(n574), .B(n573), .Z(n575) );
  XOR U578 ( .A(n576), .B(n575), .Z(n285) );
  XOR U579 ( .A(n284), .B(n285), .Z(n255) );
  XOR U580 ( .A(n286), .B(n255), .Z(n388) );
  XNOR U581 ( .A(x[172]), .B(y[172]), .Z(n623) );
  XNOR U582 ( .A(x[176]), .B(y[176]), .Z(n621) );
  XOR U583 ( .A(x[174]), .B(y[174]), .Z(n620) );
  XNOR U584 ( .A(n621), .B(n620), .Z(n622) );
  XOR U585 ( .A(n623), .B(n622), .Z(n636) );
  XNOR U586 ( .A(x[160]), .B(y[160]), .Z(n471) );
  XNOR U587 ( .A(x[164]), .B(y[164]), .Z(n469) );
  XOR U588 ( .A(x[162]), .B(y[162]), .Z(n468) );
  XNOR U589 ( .A(n469), .B(n468), .Z(n470) );
  XOR U590 ( .A(n471), .B(n470), .Z(n633) );
  XNOR U591 ( .A(x[178]), .B(y[178]), .Z(n611) );
  XNOR U592 ( .A(x[182]), .B(y[182]), .Z(n609) );
  XOR U593 ( .A(x[180]), .B(y[180]), .Z(n608) );
  XNOR U594 ( .A(n609), .B(n608), .Z(n610) );
  XNOR U595 ( .A(n611), .B(n610), .Z(n634) );
  XNOR U596 ( .A(n633), .B(n634), .Z(n635) );
  XOR U597 ( .A(n636), .B(n635), .Z(n387) );
  IV U598 ( .A(n387), .Z(n385) );
  XNOR U599 ( .A(x[196]), .B(y[196]), .Z(n690) );
  XNOR U600 ( .A(x[198]), .B(y[198]), .Z(n688) );
  XOR U601 ( .A(oglobal[0]), .B(n688), .Z(n689) );
  XOR U602 ( .A(n690), .B(n689), .Z(n292) );
  XNOR U603 ( .A(x[124]), .B(y[124]), .Z(n429) );
  XNOR U604 ( .A(x[128]), .B(y[128]), .Z(n427) );
  XNOR U605 ( .A(x[126]), .B(y[126]), .Z(n426) );
  XNOR U606 ( .A(n427), .B(n426), .Z(n428) );
  XNOR U607 ( .A(n429), .B(n428), .Z(n290) );
  XNOR U608 ( .A(x[130]), .B(y[130]), .Z(n417) );
  XNOR U609 ( .A(x[132]), .B(y[132]), .Z(n415) );
  XNOR U610 ( .A(x[134]), .B(y[134]), .Z(n414) );
  XNOR U611 ( .A(n415), .B(n414), .Z(n416) );
  XOR U612 ( .A(n417), .B(n416), .Z(n291) );
  XOR U613 ( .A(n290), .B(n291), .Z(n256) );
  XOR U614 ( .A(n292), .B(n256), .Z(n386) );
  XNOR U615 ( .A(n385), .B(n386), .Z(n257) );
  XNOR U616 ( .A(n388), .B(n257), .Z(n752) );
  XNOR U617 ( .A(x[40]), .B(y[40]), .Z(n557) );
  XNOR U618 ( .A(x[44]), .B(y[44]), .Z(n555) );
  XOR U619 ( .A(x[42]), .B(y[42]), .Z(n554) );
  XNOR U620 ( .A(n555), .B(n554), .Z(n556) );
  XOR U621 ( .A(n557), .B(n556), .Z(n299) );
  XNOR U622 ( .A(x[52]), .B(y[52]), .Z(n465) );
  XNOR U623 ( .A(x[56]), .B(y[56]), .Z(n462) );
  XNOR U624 ( .A(x[54]), .B(y[54]), .Z(n463) );
  XOR U625 ( .A(n462), .B(n463), .Z(n464) );
  XOR U626 ( .A(n465), .B(n464), .Z(n296) );
  XNOR U627 ( .A(x[46]), .B(y[46]), .Z(n459) );
  XNOR U628 ( .A(x[50]), .B(y[50]), .Z(n456) );
  XNOR U629 ( .A(x[48]), .B(y[48]), .Z(n457) );
  XOR U630 ( .A(n456), .B(n457), .Z(n458) );
  XNOR U631 ( .A(n459), .B(n458), .Z(n297) );
  XNOR U632 ( .A(n296), .B(n297), .Z(n298) );
  XNOR U633 ( .A(n299), .B(n298), .Z(n519) );
  XNOR U634 ( .A(x[4]), .B(y[4]), .Z(n584) );
  XNOR U635 ( .A(x[6]), .B(y[6]), .Z(n581) );
  XNOR U636 ( .A(x[8]), .B(y[8]), .Z(n582) );
  XOR U637 ( .A(n581), .B(n582), .Z(n583) );
  XOR U638 ( .A(n584), .B(n583), .Z(n281) );
  XNOR U639 ( .A(x[16]), .B(y[16]), .Z(n605) );
  XNOR U640 ( .A(x[18]), .B(y[18]), .Z(n602) );
  XNOR U641 ( .A(x[20]), .B(y[20]), .Z(n603) );
  XOR U642 ( .A(n602), .B(n603), .Z(n604) );
  XOR U643 ( .A(n605), .B(n604), .Z(n278) );
  XNOR U644 ( .A(x[10]), .B(y[10]), .Z(n599) );
  XNOR U645 ( .A(x[12]), .B(y[12]), .Z(n596) );
  XNOR U646 ( .A(x[14]), .B(y[14]), .Z(n597) );
  XOR U647 ( .A(n596), .B(n597), .Z(n598) );
  XNOR U648 ( .A(n599), .B(n598), .Z(n279) );
  XNOR U649 ( .A(n278), .B(n279), .Z(n280) );
  XNOR U650 ( .A(n281), .B(n280), .Z(n520) );
  XNOR U651 ( .A(x[22]), .B(y[22]), .Z(n619) );
  XNOR U652 ( .A(x[26]), .B(y[26]), .Z(n617) );
  XOR U653 ( .A(x[24]), .B(y[24]), .Z(n616) );
  XNOR U654 ( .A(n617), .B(n616), .Z(n618) );
  XOR U655 ( .A(n619), .B(n618), .Z(n345) );
  XNOR U656 ( .A(x[28]), .B(y[28]), .Z(n615) );
  XNOR U657 ( .A(x[32]), .B(y[32]), .Z(n613) );
  XOR U658 ( .A(x[30]), .B(y[30]), .Z(n612) );
  XNOR U659 ( .A(n613), .B(n612), .Z(n614) );
  XOR U660 ( .A(n615), .B(n614), .Z(n342) );
  XNOR U661 ( .A(x[34]), .B(y[34]), .Z(n551) );
  XNOR U662 ( .A(x[38]), .B(y[38]), .Z(n549) );
  XNOR U663 ( .A(x[36]), .B(y[36]), .Z(n548) );
  XNOR U664 ( .A(n549), .B(n548), .Z(n550) );
  XOR U665 ( .A(n551), .B(n550), .Z(n343) );
  XNOR U666 ( .A(n342), .B(n343), .Z(n344) );
  XOR U667 ( .A(n345), .B(n344), .Z(n518) );
  XOR U668 ( .A(n520), .B(n518), .Z(n258) );
  XNOR U669 ( .A(n519), .B(n258), .Z(n396) );
  XNOR U670 ( .A(x[166]), .B(y[166]), .Z(n547) );
  XNOR U671 ( .A(x[170]), .B(y[170]), .Z(n545) );
  XOR U672 ( .A(x[168]), .B(y[168]), .Z(n544) );
  XNOR U673 ( .A(n545), .B(n544), .Z(n546) );
  XOR U674 ( .A(n547), .B(n546), .Z(n449) );
  XNOR U675 ( .A(x[154]), .B(y[154]), .Z(n483) );
  XNOR U676 ( .A(x[156]), .B(y[156]), .Z(n481) );
  XOR U677 ( .A(x[158]), .B(y[158]), .Z(n480) );
  XNOR U678 ( .A(n481), .B(n480), .Z(n482) );
  XNOR U679 ( .A(n483), .B(n482), .Z(n680) );
  XNOR U680 ( .A(x[148]), .B(y[148]), .Z(n512) );
  XNOR U681 ( .A(x[150]), .B(y[150]), .Z(n510) );
  XOR U682 ( .A(x[152]), .B(y[152]), .Z(n509) );
  XNOR U683 ( .A(n510), .B(n509), .Z(n511) );
  XOR U684 ( .A(n512), .B(n511), .Z(n678) );
  XNOR U685 ( .A(x[184]), .B(y[184]), .Z(n594) );
  XNOR U686 ( .A(x[186]), .B(y[186]), .Z(n592) );
  XOR U687 ( .A(x[188]), .B(y[188]), .Z(n591) );
  XNOR U688 ( .A(n592), .B(n591), .Z(n593) );
  XNOR U689 ( .A(n594), .B(n593), .Z(n677) );
  IV U690 ( .A(n677), .Z(n679) );
  XNOR U691 ( .A(n678), .B(n679), .Z(n259) );
  XNOR U692 ( .A(n680), .B(n259), .Z(n446) );
  XNOR U693 ( .A(x[190]), .B(y[190]), .Z(n317) );
  XNOR U694 ( .A(x[192]), .B(y[192]), .Z(n315) );
  XNOR U695 ( .A(x[194]), .B(y[194]), .Z(n314) );
  XNOR U696 ( .A(n315), .B(n314), .Z(n316) );
  XOR U697 ( .A(n317), .B(n316), .Z(n734) );
  XNOR U698 ( .A(x[136]), .B(y[136]), .Z(n407) );
  XNOR U699 ( .A(x[138]), .B(y[138]), .Z(n405) );
  XNOR U700 ( .A(x[140]), .B(y[140]), .Z(n404) );
  XNOR U701 ( .A(n405), .B(n404), .Z(n406) );
  XNOR U702 ( .A(n407), .B(n406), .Z(n733) );
  XNOR U703 ( .A(x[142]), .B(y[142]), .Z(n443) );
  XNOR U704 ( .A(x[146]), .B(y[146]), .Z(n441) );
  XOR U705 ( .A(x[144]), .B(y[144]), .Z(n440) );
  XNOR U706 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U707 ( .A(n443), .B(n442), .Z(n732) );
  XOR U708 ( .A(n733), .B(n732), .Z(n260) );
  XNOR U709 ( .A(n734), .B(n260), .Z(n447) );
  IV U710 ( .A(n447), .Z(n445) );
  XOR U711 ( .A(n446), .B(n445), .Z(n261) );
  XNOR U712 ( .A(n449), .B(n261), .Z(n394) );
  XNOR U713 ( .A(x[103]), .B(y[103]), .Z(n746) );
  XNOR U714 ( .A(x[195]), .B(y[195]), .Z(n744) );
  XOR U715 ( .A(x[101]), .B(y[101]), .Z(n743) );
  XNOR U716 ( .A(n744), .B(n743), .Z(n745) );
  XNOR U717 ( .A(n746), .B(n745), .Z(n500) );
  XNOR U718 ( .A(x[93]), .B(y[93]), .Z(n668) );
  XNOR U719 ( .A(x[91]), .B(y[91]), .Z(n666) );
  XOR U720 ( .A(x[89]), .B(y[89]), .Z(n665) );
  XNOR U721 ( .A(n666), .B(n665), .Z(n667) );
  XNOR U722 ( .A(n668), .B(n667), .Z(n501) );
  XNOR U723 ( .A(x[99]), .B(y[99]), .Z(n742) );
  XNOR U724 ( .A(x[97]), .B(y[97]), .Z(n740) );
  XOR U725 ( .A(x[95]), .B(y[95]), .Z(n739) );
  XNOR U726 ( .A(n740), .B(n739), .Z(n741) );
  XOR U727 ( .A(n742), .B(n741), .Z(n499) );
  XOR U728 ( .A(n501), .B(n499), .Z(n262) );
  XNOR U729 ( .A(n500), .B(n262), .Z(n534) );
  XNOR U730 ( .A(x[57]), .B(y[57]), .Z(n376) );
  XNOR U731 ( .A(x[55]), .B(y[55]), .Z(n374) );
  XOR U732 ( .A(x[53]), .B(y[53]), .Z(n373) );
  XNOR U733 ( .A(n374), .B(n373), .Z(n375) );
  XNOR U734 ( .A(n376), .B(n375), .Z(n494) );
  XNOR U735 ( .A(x[69]), .B(y[69]), .Z(n731) );
  XNOR U736 ( .A(x[67]), .B(y[67]), .Z(n729) );
  XOR U737 ( .A(x[65]), .B(y[65]), .Z(n728) );
  XNOR U738 ( .A(n729), .B(n728), .Z(n730) );
  XOR U739 ( .A(n731), .B(n730), .Z(n492) );
  XNOR U740 ( .A(x[63]), .B(y[63]), .Z(n723) );
  XNOR U741 ( .A(x[61]), .B(y[61]), .Z(n721) );
  XOR U742 ( .A(x[59]), .B(y[59]), .Z(n720) );
  XNOR U743 ( .A(n721), .B(n720), .Z(n722) );
  XNOR U744 ( .A(n723), .B(n722), .Z(n493) );
  XOR U745 ( .A(n492), .B(n493), .Z(n263) );
  XOR U746 ( .A(n494), .B(n263), .Z(n532) );
  XNOR U747 ( .A(x[87]), .B(y[87]), .Z(n676) );
  XNOR U748 ( .A(x[85]), .B(y[85]), .Z(n674) );
  XOR U749 ( .A(x[83]), .B(y[83]), .Z(n673) );
  XNOR U750 ( .A(n674), .B(n673), .Z(n675) );
  XOR U751 ( .A(n676), .B(n675), .Z(n497) );
  XNOR U752 ( .A(x[81]), .B(y[81]), .Z(n672) );
  XNOR U753 ( .A(x[79]), .B(y[79]), .Z(n670) );
  XOR U754 ( .A(x[77]), .B(y[77]), .Z(n669) );
  XNOR U755 ( .A(n670), .B(n669), .Z(n671) );
  XNOR U756 ( .A(n672), .B(n671), .Z(n495) );
  XNOR U757 ( .A(x[75]), .B(y[75]), .Z(n727) );
  XNOR U758 ( .A(x[73]), .B(y[73]), .Z(n725) );
  XOR U759 ( .A(x[71]), .B(y[71]), .Z(n724) );
  XNOR U760 ( .A(n725), .B(n724), .Z(n726) );
  XOR U761 ( .A(n727), .B(n726), .Z(n496) );
  XOR U762 ( .A(n495), .B(n496), .Z(n264) );
  XOR U763 ( .A(n497), .B(n264), .Z(n531) );
  IV U764 ( .A(n531), .Z(n533) );
  XNOR U765 ( .A(n532), .B(n533), .Z(n265) );
  XOR U766 ( .A(n534), .B(n265), .Z(n384) );
  XNOR U767 ( .A(x[135]), .B(y[135]), .Z(n361) );
  XNOR U768 ( .A(x[179]), .B(y[179]), .Z(n359) );
  XOR U769 ( .A(x[133]), .B(y[133]), .Z(n358) );
  XNOR U770 ( .A(n359), .B(n358), .Z(n360) );
  XOR U771 ( .A(n361), .B(n360), .Z(n402) );
  XNOR U772 ( .A(x[131]), .B(y[131]), .Z(n655) );
  XNOR U773 ( .A(x[181]), .B(y[181]), .Z(n653) );
  XOR U774 ( .A(x[129]), .B(y[129]), .Z(n652) );
  XNOR U775 ( .A(n653), .B(n652), .Z(n654) );
  XNOR U776 ( .A(n655), .B(n654), .Z(n403) );
  XNOR U777 ( .A(x[139]), .B(y[139]), .Z(n365) );
  XNOR U778 ( .A(x[177]), .B(y[177]), .Z(n363) );
  XOR U779 ( .A(x[137]), .B(y[137]), .Z(n362) );
  XNOR U780 ( .A(n363), .B(n362), .Z(n364) );
  XOR U781 ( .A(n365), .B(n364), .Z(n401) );
  XOR U782 ( .A(n403), .B(n401), .Z(n266) );
  XNOR U783 ( .A(n402), .B(n266), .Z(n381) );
  XNOR U784 ( .A(x[143]), .B(y[143]), .Z(n357) );
  XNOR U785 ( .A(x[175]), .B(y[175]), .Z(n355) );
  XOR U786 ( .A(x[141]), .B(y[141]), .Z(n354) );
  XNOR U787 ( .A(n355), .B(n354), .Z(n356) );
  XNOR U788 ( .A(n357), .B(n356), .Z(n322) );
  XNOR U789 ( .A(x[147]), .B(y[147]), .Z(n642) );
  XNOR U790 ( .A(x[173]), .B(y[173]), .Z(n640) );
  XOR U791 ( .A(x[145]), .B(y[145]), .Z(n639) );
  XNOR U792 ( .A(n640), .B(n639), .Z(n641) );
  XOR U793 ( .A(n642), .B(n641), .Z(n320) );
  XNOR U794 ( .A(x[163]), .B(y[163]), .Z(n650) );
  XNOR U795 ( .A(x[161]), .B(y[161]), .Z(n648) );
  XOR U796 ( .A(x[159]), .B(y[159]), .Z(n647) );
  XNOR U797 ( .A(n648), .B(n647), .Z(n649) );
  XNOR U798 ( .A(n650), .B(n649), .Z(n321) );
  XOR U799 ( .A(n320), .B(n321), .Z(n267) );
  XNOR U800 ( .A(n322), .B(n267), .Z(n382) );
  XNOR U801 ( .A(n381), .B(n382), .Z(n383) );
  XNOR U802 ( .A(n384), .B(n383), .Z(n393) );
  XNOR U803 ( .A(n394), .B(n393), .Z(n395) );
  XOR U804 ( .A(n396), .B(n395), .Z(n751) );
  XNOR U805 ( .A(n752), .B(n751), .Z(n753) );
  XNOR U806 ( .A(x[9]), .B(y[9]), .Z(n311) );
  XNOR U807 ( .A(x[7]), .B(y[7]), .Z(n309) );
  XNOR U808 ( .A(x[5]), .B(y[5]), .Z(n308) );
  XNOR U809 ( .A(n309), .B(n308), .Z(n310) );
  XNOR U810 ( .A(n311), .B(n310), .Z(n367) );
  XNOR U811 ( .A(x[1]), .B(y[1]), .Z(n588) );
  XOR U812 ( .A(x[0]), .B(y[0]), .Z(n587) );
  XNOR U813 ( .A(n588), .B(n587), .Z(n590) );
  XOR U814 ( .A(x[3]), .B(y[3]), .Z(n589) );
  XNOR U815 ( .A(n590), .B(n589), .Z(n368) );
  XNOR U816 ( .A(x[15]), .B(y[15]), .Z(n305) );
  XNOR U817 ( .A(x[13]), .B(y[13]), .Z(n303) );
  XNOR U818 ( .A(x[11]), .B(y[11]), .Z(n302) );
  XNOR U819 ( .A(n303), .B(n302), .Z(n304) );
  XNOR U820 ( .A(n305), .B(n304), .Z(n366) );
  XNOR U821 ( .A(n368), .B(n366), .Z(n268) );
  XNOR U822 ( .A(n367), .B(n268), .Z(n541) );
  XNOR U823 ( .A(x[33]), .B(y[33]), .Z(n704) );
  XNOR U824 ( .A(x[31]), .B(y[31]), .Z(n702) );
  XNOR U825 ( .A(x[29]), .B(y[29]), .Z(n701) );
  XNOR U826 ( .A(n702), .B(n701), .Z(n703) );
  XOR U827 ( .A(n704), .B(n703), .Z(n455) );
  XNOR U828 ( .A(x[27]), .B(y[27]), .Z(n696) );
  XNOR U829 ( .A(x[25]), .B(y[25]), .Z(n694) );
  XOR U830 ( .A(x[23]), .B(y[23]), .Z(n693) );
  XNOR U831 ( .A(n694), .B(n693), .Z(n695) );
  XNOR U832 ( .A(n696), .B(n695), .Z(n453) );
  XNOR U833 ( .A(x[21]), .B(y[21]), .Z(n687) );
  XNOR U834 ( .A(x[19]), .B(y[19]), .Z(n685) );
  XOR U835 ( .A(x[17]), .B(y[17]), .Z(n684) );
  XNOR U836 ( .A(n685), .B(n684), .Z(n686) );
  XOR U837 ( .A(n687), .B(n686), .Z(n454) );
  XOR U838 ( .A(n453), .B(n454), .Z(n269) );
  XOR U839 ( .A(n455), .B(n269), .Z(n538) );
  XNOR U840 ( .A(x[45]), .B(y[45]), .Z(n372) );
  XNOR U841 ( .A(x[43]), .B(y[43]), .Z(n370) );
  XOR U842 ( .A(x[41]), .B(y[41]), .Z(n369) );
  XNOR U843 ( .A(n370), .B(n369), .Z(n371) );
  XOR U844 ( .A(n372), .B(n371), .Z(n476) );
  XNOR U845 ( .A(x[39]), .B(y[39]), .Z(n716) );
  XNOR U846 ( .A(x[37]), .B(y[37]), .Z(n714) );
  XNOR U847 ( .A(x[35]), .B(y[35]), .Z(n713) );
  XNOR U848 ( .A(n714), .B(n713), .Z(n715) );
  XOR U849 ( .A(n716), .B(n715), .Z(n474) );
  IV U850 ( .A(n474), .Z(n472) );
  XNOR U851 ( .A(x[51]), .B(y[51]), .Z(n380) );
  XNOR U852 ( .A(x[49]), .B(y[49]), .Z(n378) );
  XOR U853 ( .A(x[47]), .B(y[47]), .Z(n377) );
  XNOR U854 ( .A(n378), .B(n377), .Z(n379) );
  XNOR U855 ( .A(n380), .B(n379), .Z(n473) );
  XOR U856 ( .A(n472), .B(n473), .Z(n270) );
  XNOR U857 ( .A(n476), .B(n270), .Z(n539) );
  XOR U858 ( .A(n538), .B(n539), .Z(n540) );
  XNOR U859 ( .A(n541), .B(n540), .Z(n523) );
  XNOR U860 ( .A(x[94]), .B(y[94]), .Z(n413) );
  XNOR U861 ( .A(x[98]), .B(y[98]), .Z(n411) );
  XOR U862 ( .A(x[96]), .B(y[96]), .Z(n410) );
  XNOR U863 ( .A(n411), .B(n410), .Z(n412) );
  XOR U864 ( .A(n413), .B(n412), .Z(n353) );
  XNOR U865 ( .A(x[100]), .B(y[100]), .Z(n564) );
  XNOR U866 ( .A(x[104]), .B(y[104]), .Z(n562) );
  XNOR U867 ( .A(x[102]), .B(y[102]), .Z(n561) );
  XNOR U868 ( .A(n562), .B(n561), .Z(n563) );
  XOR U869 ( .A(n564), .B(n563), .Z(n352) );
  XNOR U870 ( .A(x[106]), .B(y[106]), .Z(n570) );
  XNOR U871 ( .A(x[108]), .B(y[108]), .Z(n568) );
  XNOR U872 ( .A(x[110]), .B(y[110]), .Z(n567) );
  XNOR U873 ( .A(n568), .B(n567), .Z(n569) );
  XOR U874 ( .A(n570), .B(n569), .Z(n351) );
  XNOR U875 ( .A(n352), .B(n351), .Z(n271) );
  XNOR U876 ( .A(n353), .B(n271), .Z(n528) );
  XNOR U877 ( .A(x[58]), .B(y[58]), .Z(n491) );
  XNOR U878 ( .A(x[62]), .B(y[62]), .Z(n489) );
  XOR U879 ( .A(x[60]), .B(y[60]), .Z(n488) );
  XNOR U880 ( .A(n489), .B(n488), .Z(n490) );
  XOR U881 ( .A(n491), .B(n490), .Z(n294) );
  XNOR U882 ( .A(x[70]), .B(y[70]), .Z(n516) );
  XNOR U883 ( .A(x[74]), .B(y[74]), .Z(n514) );
  XOR U884 ( .A(x[72]), .B(y[72]), .Z(n513) );
  XNOR U885 ( .A(n514), .B(n513), .Z(n515) );
  XNOR U886 ( .A(n516), .B(n515), .Z(n295) );
  XNOR U887 ( .A(x[64]), .B(y[64]), .Z(n487) );
  XNOR U888 ( .A(x[68]), .B(y[68]), .Z(n485) );
  XOR U889 ( .A(x[66]), .B(y[66]), .Z(n484) );
  XNOR U890 ( .A(n485), .B(n484), .Z(n486) );
  XOR U891 ( .A(n487), .B(n486), .Z(n293) );
  XOR U892 ( .A(n295), .B(n293), .Z(n272) );
  XNOR U893 ( .A(n294), .B(n272), .Z(n525) );
  XNOR U894 ( .A(x[82]), .B(y[82]), .Z(n435) );
  XNOR U895 ( .A(x[86]), .B(y[86]), .Z(n433) );
  XOR U896 ( .A(x[84]), .B(y[84]), .Z(n432) );
  XNOR U897 ( .A(n433), .B(n432), .Z(n434) );
  XNOR U898 ( .A(n435), .B(n434), .Z(n350) );
  XNOR U899 ( .A(x[88]), .B(y[88]), .Z(n439) );
  XNOR U900 ( .A(x[92]), .B(y[92]), .Z(n437) );
  XOR U901 ( .A(x[90]), .B(y[90]), .Z(n436) );
  XNOR U902 ( .A(n437), .B(n436), .Z(n438) );
  XOR U903 ( .A(n439), .B(n438), .Z(n348) );
  XNOR U904 ( .A(x[76]), .B(y[76]), .Z(n508) );
  XNOR U905 ( .A(x[80]), .B(y[80]), .Z(n506) );
  XOR U906 ( .A(x[78]), .B(y[78]), .Z(n505) );
  XNOR U907 ( .A(n506), .B(n505), .Z(n507) );
  XNOR U908 ( .A(n508), .B(n507), .Z(n349) );
  XOR U909 ( .A(n348), .B(n349), .Z(n273) );
  XNOR U910 ( .A(n350), .B(n273), .Z(n526) );
  XNOR U911 ( .A(n525), .B(n526), .Z(n527) );
  XOR U912 ( .A(n528), .B(n527), .Z(n524) );
  XNOR U913 ( .A(x[111]), .B(y[111]), .Z(n332) );
  XNOR U914 ( .A(x[191]), .B(y[191]), .Z(n330) );
  XNOR U915 ( .A(x[109]), .B(y[109]), .Z(n329) );
  XOR U916 ( .A(n330), .B(n329), .Z(n331) );
  XOR U917 ( .A(n332), .B(n331), .Z(n504) );
  XNOR U918 ( .A(x[107]), .B(y[107]), .Z(n738) );
  XNOR U919 ( .A(x[193]), .B(y[193]), .Z(n736) );
  XOR U920 ( .A(x[105]), .B(y[105]), .Z(n735) );
  XNOR U921 ( .A(n736), .B(n735), .Z(n737) );
  XNOR U922 ( .A(n738), .B(n737), .Z(n502) );
  XNOR U923 ( .A(x[115]), .B(y[115]), .Z(n338) );
  XNOR U924 ( .A(x[189]), .B(y[189]), .Z(n336) );
  XNOR U925 ( .A(x[113]), .B(y[113]), .Z(n335) );
  XOR U926 ( .A(n336), .B(n335), .Z(n337) );
  XNOR U927 ( .A(n338), .B(n337), .Z(n503) );
  XNOR U928 ( .A(n502), .B(n503), .Z(n274) );
  XNOR U929 ( .A(n504), .B(n274), .Z(n399) );
  XNOR U930 ( .A(x[165]), .B(y[165]), .Z(n627) );
  XNOR U931 ( .A(x[169]), .B(y[169]), .Z(n625) );
  XOR U932 ( .A(x[167]), .B(y[167]), .Z(n624) );
  XNOR U933 ( .A(n625), .B(n624), .Z(n626) );
  XOR U934 ( .A(n627), .B(n626), .Z(n700) );
  XNOR U935 ( .A(x[151]), .B(y[151]), .Z(n646) );
  XNOR U936 ( .A(x[171]), .B(y[171]), .Z(n644) );
  XOR U937 ( .A(x[149]), .B(y[149]), .Z(n643) );
  XNOR U938 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U939 ( .A(n646), .B(n645), .Z(n698) );
  XNOR U940 ( .A(x[155]), .B(y[155]), .Z(n631) );
  XNOR U941 ( .A(x[157]), .B(y[157]), .Z(n629) );
  XOR U942 ( .A(x[153]), .B(y[153]), .Z(n628) );
  XNOR U943 ( .A(n629), .B(n628), .Z(n630) );
  XOR U944 ( .A(n631), .B(n630), .Z(n699) );
  XOR U945 ( .A(n698), .B(n699), .Z(n275) );
  XNOR U946 ( .A(n700), .B(n275), .Z(n397) );
  XNOR U947 ( .A(x[123]), .B(y[123]), .Z(n659) );
  XNOR U948 ( .A(x[185]), .B(y[185]), .Z(n657) );
  XOR U949 ( .A(x[121]), .B(y[121]), .Z(n656) );
  XNOR U950 ( .A(n657), .B(n656), .Z(n658) );
  XOR U951 ( .A(n659), .B(n658), .Z(n560) );
  XNOR U952 ( .A(x[127]), .B(y[127]), .Z(n663) );
  XNOR U953 ( .A(x[183]), .B(y[183]), .Z(n661) );
  XOR U954 ( .A(x[125]), .B(y[125]), .Z(n660) );
  XNOR U955 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U956 ( .A(n663), .B(n662), .Z(n558) );
  XNOR U957 ( .A(x[119]), .B(y[119]), .Z(n326) );
  XNOR U958 ( .A(x[187]), .B(y[187]), .Z(n324) );
  XNOR U959 ( .A(x[117]), .B(y[117]), .Z(n323) );
  XNOR U960 ( .A(n324), .B(n323), .Z(n325) );
  XNOR U961 ( .A(n326), .B(n325), .Z(n559) );
  XOR U962 ( .A(n558), .B(n559), .Z(n276) );
  XNOR U963 ( .A(n560), .B(n276), .Z(n398) );
  XOR U964 ( .A(n397), .B(n398), .Z(n400) );
  XNOR U965 ( .A(n399), .B(n400), .Z(n522) );
  XOR U966 ( .A(n524), .B(n522), .Z(n277) );
  XNOR U967 ( .A(n523), .B(n277), .Z(n754) );
  XOR U968 ( .A(n753), .B(n754), .Z(o[0]) );
  NANDN U969 ( .A(n279), .B(n278), .Z(n283) );
  NAND U970 ( .A(n281), .B(n280), .Z(n282) );
  NAND U971 ( .A(n283), .B(n282), .Z(n934) );
  NANDN U972 ( .A(n285), .B(n284), .Z(n289) );
  ANDN U973 ( .B(n285), .A(n284), .Z(n287) );
  NANDN U974 ( .A(n287), .B(n286), .Z(n288) );
  AND U975 ( .A(n289), .B(n288), .Z(n932) );
  XNOR U976 ( .A(n934), .B(n933), .Z(n892) );
  NANDN U977 ( .A(n297), .B(n296), .Z(n301) );
  NAND U978 ( .A(n299), .B(n298), .Z(n300) );
  AND U979 ( .A(n301), .B(n300), .Z(n890) );
  XNOR U980 ( .A(n889), .B(n890), .Z(n891) );
  XNOR U981 ( .A(n892), .B(n891), .Z(n776) );
  OR U982 ( .A(n303), .B(n302), .Z(n307) );
  OR U983 ( .A(n305), .B(n304), .Z(n306) );
  NAND U984 ( .A(n307), .B(n306), .Z(n811) );
  OR U985 ( .A(n309), .B(n308), .Z(n313) );
  OR U986 ( .A(n311), .B(n310), .Z(n312) );
  AND U987 ( .A(n313), .B(n312), .Z(n810) );
  XNOR U988 ( .A(n811), .B(n810), .Z(n812) );
  OR U989 ( .A(n315), .B(n314), .Z(n319) );
  OR U990 ( .A(n317), .B(n316), .Z(n318) );
  AND U991 ( .A(n319), .B(n318), .Z(n813) );
  XNOR U992 ( .A(n812), .B(n813), .Z(n999) );
  OR U993 ( .A(n324), .B(n323), .Z(n328) );
  OR U994 ( .A(n326), .B(n325), .Z(n327) );
  NAND U995 ( .A(n328), .B(n327), .Z(n898) );
  OR U996 ( .A(n330), .B(n329), .Z(n334) );
  NANDN U997 ( .A(n332), .B(n331), .Z(n333) );
  AND U998 ( .A(n334), .B(n333), .Z(n897) );
  XNOR U999 ( .A(n898), .B(n897), .Z(n899) );
  OR U1000 ( .A(n336), .B(n335), .Z(n340) );
  NANDN U1001 ( .A(n338), .B(n337), .Z(n339) );
  AND U1002 ( .A(n340), .B(n339), .Z(n900) );
  XOR U1003 ( .A(n899), .B(n900), .Z(n998) );
  XOR U1004 ( .A(n997), .B(n998), .Z(n341) );
  XOR U1005 ( .A(n999), .B(n341), .Z(n777) );
  XOR U1006 ( .A(n776), .B(n777), .Z(n778) );
  NANDN U1007 ( .A(n343), .B(n342), .Z(n347) );
  NAND U1008 ( .A(n345), .B(n344), .Z(n346) );
  NAND U1009 ( .A(n347), .B(n346), .Z(n986) );
  XOR U1010 ( .A(n984), .B(n985), .Z(n987) );
  XOR U1011 ( .A(n986), .B(n987), .Z(n779) );
  XOR U1012 ( .A(n778), .B(n779), .Z(n766) );
  XNOR U1013 ( .A(n820), .B(n819), .Z(n822) );
  XNOR U1014 ( .A(n822), .B(n821), .Z(n938) );
  XNOR U1015 ( .A(n938), .B(n937), .Z(n939) );
  XNOR U1016 ( .A(n907), .B(n906), .Z(n909) );
  XNOR U1017 ( .A(n909), .B(n908), .Z(n940) );
  XOR U1018 ( .A(n939), .B(n940), .Z(n910) );
  NANDN U1019 ( .A(n385), .B(n386), .Z(n391) );
  NOR U1020 ( .A(n387), .B(n386), .Z(n389) );
  OR U1021 ( .A(n389), .B(n388), .Z(n390) );
  NAND U1022 ( .A(n391), .B(n390), .Z(n911) );
  XNOR U1023 ( .A(n912), .B(n911), .Z(n392) );
  XNOR U1024 ( .A(n910), .B(n392), .Z(n764) );
  XNOR U1025 ( .A(n764), .B(n765), .Z(n767) );
  XNOR U1026 ( .A(n766), .B(n767), .Z(n1010) );
  OR U1027 ( .A(n405), .B(n404), .Z(n409) );
  OR U1028 ( .A(n407), .B(n406), .Z(n408) );
  AND U1029 ( .A(n409), .B(n408), .Z(n809) );
  OR U1030 ( .A(n415), .B(n414), .Z(n419) );
  OR U1031 ( .A(n417), .B(n416), .Z(n418) );
  AND U1032 ( .A(n419), .B(n418), .Z(n807) );
  XOR U1033 ( .A(n806), .B(n807), .Z(n808) );
  XNOR U1034 ( .A(n809), .B(n808), .Z(n977) );
  OR U1035 ( .A(n421), .B(n420), .Z(n425) );
  OR U1036 ( .A(n423), .B(n422), .Z(n424) );
  NAND U1037 ( .A(n425), .B(n424), .Z(n975) );
  OR U1038 ( .A(n427), .B(n426), .Z(n431) );
  OR U1039 ( .A(n429), .B(n428), .Z(n430) );
  AND U1040 ( .A(n431), .B(n430), .Z(n974) );
  XNOR U1041 ( .A(n975), .B(n974), .Z(n976) );
  XNOR U1042 ( .A(n977), .B(n976), .Z(n834) );
  XOR U1043 ( .A(n833), .B(n834), .Z(n835) );
  XNOR U1044 ( .A(n873), .B(n872), .Z(n444) );
  XNOR U1045 ( .A(n871), .B(n444), .Z(n836) );
  XOR U1046 ( .A(n835), .B(n836), .Z(n783) );
  NANDN U1047 ( .A(n445), .B(n446), .Z(n451) );
  NOR U1048 ( .A(n447), .B(n446), .Z(n448) );
  OR U1049 ( .A(n449), .B(n448), .Z(n450) );
  AND U1050 ( .A(n451), .B(n450), .Z(n784) );
  IV U1051 ( .A(n784), .Z(n782) );
  XOR U1052 ( .A(n783), .B(n782), .Z(n452) );
  XOR U1053 ( .A(n785), .B(n452), .Z(n760) );
  OR U1054 ( .A(n457), .B(n456), .Z(n461) );
  NANDN U1055 ( .A(n459), .B(n458), .Z(n460) );
  NAND U1056 ( .A(n461), .B(n460), .Z(n851) );
  OR U1057 ( .A(n463), .B(n462), .Z(n467) );
  NANDN U1058 ( .A(n465), .B(n464), .Z(n466) );
  AND U1059 ( .A(n467), .B(n466), .Z(n850) );
  XNOR U1060 ( .A(n851), .B(n850), .Z(n852) );
  XNOR U1061 ( .A(n852), .B(n853), .Z(n839) );
  NANDN U1062 ( .A(n472), .B(n473), .Z(n478) );
  NOR U1063 ( .A(n474), .B(n473), .Z(n475) );
  OR U1064 ( .A(n476), .B(n475), .Z(n477) );
  NAND U1065 ( .A(n478), .B(n477), .Z(n840) );
  XOR U1066 ( .A(n839), .B(n840), .Z(n479) );
  XNOR U1067 ( .A(n841), .B(n479), .Z(n773) );
  XNOR U1068 ( .A(n862), .B(n863), .Z(n864) );
  XOR U1069 ( .A(n865), .B(n864), .Z(n965) );
  IV U1070 ( .A(n965), .Z(n966) );
  IV U1071 ( .A(n964), .Z(n967) );
  XNOR U1072 ( .A(n968), .B(n967), .Z(n498) );
  XNOR U1073 ( .A(n966), .B(n498), .Z(n771) );
  XNOR U1074 ( .A(n893), .B(n894), .Z(n896) );
  XNOR U1075 ( .A(n860), .B(n859), .Z(n517) );
  XNOR U1076 ( .A(n861), .B(n517), .Z(n895) );
  XNOR U1077 ( .A(n896), .B(n895), .Z(n770) );
  XNOR U1078 ( .A(n771), .B(n770), .Z(n772) );
  XOR U1079 ( .A(n773), .B(n772), .Z(n758) );
  IV U1080 ( .A(n759), .Z(n757) );
  XNOR U1081 ( .A(n758), .B(n757), .Z(n521) );
  XOR U1082 ( .A(n760), .B(n521), .Z(n1009) );
  NANDN U1083 ( .A(n526), .B(n525), .Z(n530) );
  NAND U1084 ( .A(n528), .B(n527), .Z(n529) );
  NAND U1085 ( .A(n530), .B(n529), .Z(n916) );
  NANDN U1086 ( .A(n531), .B(n532), .Z(n537) );
  NOR U1087 ( .A(n533), .B(n532), .Z(n535) );
  OR U1088 ( .A(n535), .B(n534), .Z(n536) );
  NAND U1089 ( .A(n537), .B(n536), .Z(n913) );
  NAND U1090 ( .A(n539), .B(n538), .Z(n543) );
  NAND U1091 ( .A(n541), .B(n540), .Z(n542) );
  AND U1092 ( .A(n543), .B(n542), .Z(n914) );
  XNOR U1093 ( .A(n913), .B(n914), .Z(n915) );
  XNOR U1094 ( .A(n916), .B(n915), .Z(n793) );
  OR U1095 ( .A(n549), .B(n548), .Z(n553) );
  OR U1096 ( .A(n551), .B(n550), .Z(n552) );
  AND U1097 ( .A(n553), .B(n552), .Z(n797) );
  XNOR U1098 ( .A(n797), .B(n798), .Z(n800) );
  XNOR U1099 ( .A(n799), .B(n800), .Z(n843) );
  IV U1100 ( .A(n844), .Z(n842) );
  OR U1101 ( .A(n562), .B(n561), .Z(n566) );
  OR U1102 ( .A(n564), .B(n563), .Z(n565) );
  NAND U1103 ( .A(n566), .B(n565), .Z(n803) );
  OR U1104 ( .A(n568), .B(n567), .Z(n572) );
  OR U1105 ( .A(n570), .B(n569), .Z(n571) );
  NAND U1106 ( .A(n572), .B(n571), .Z(n805) );
  OR U1107 ( .A(n574), .B(n573), .Z(n578) );
  OR U1108 ( .A(n576), .B(n575), .Z(n577) );
  AND U1109 ( .A(n578), .B(n577), .Z(n804) );
  XOR U1110 ( .A(n805), .B(n804), .Z(n579) );
  XNOR U1111 ( .A(n803), .B(n579), .Z(n845) );
  XNOR U1112 ( .A(n842), .B(n845), .Z(n580) );
  XNOR U1113 ( .A(n843), .B(n580), .Z(n917) );
  OR U1114 ( .A(n582), .B(n581), .Z(n586) );
  NANDN U1115 ( .A(n584), .B(n583), .Z(n585) );
  NAND U1116 ( .A(n586), .B(n585), .Z(n831) );
  XNOR U1117 ( .A(n829), .B(n830), .Z(n595) );
  XOR U1118 ( .A(n831), .B(n595), .Z(n943) );
  OR U1119 ( .A(n597), .B(n596), .Z(n601) );
  NANDN U1120 ( .A(n599), .B(n598), .Z(n600) );
  NAND U1121 ( .A(n601), .B(n600), .Z(n823) );
  OR U1122 ( .A(n603), .B(n602), .Z(n607) );
  NANDN U1123 ( .A(n605), .B(n604), .Z(n606) );
  AND U1124 ( .A(n607), .B(n606), .Z(n824) );
  XNOR U1125 ( .A(n823), .B(n824), .Z(n825) );
  XOR U1126 ( .A(n825), .B(n826), .Z(n944) );
  XNOR U1127 ( .A(n943), .B(n944), .Z(n945) );
  XNOR U1128 ( .A(n981), .B(n980), .Z(n983) );
  XNOR U1129 ( .A(n983), .B(n982), .Z(n946) );
  XOR U1130 ( .A(n945), .B(n946), .Z(n918) );
  XOR U1131 ( .A(n917), .B(n918), .Z(n919) );
  XNOR U1132 ( .A(n973), .B(oglobal[1]), .Z(n632) );
  XNOR U1133 ( .A(n972), .B(n632), .Z(n1003) );
  NANDN U1134 ( .A(n634), .B(n633), .Z(n638) );
  NAND U1135 ( .A(n636), .B(n635), .Z(n637) );
  NAND U1136 ( .A(n638), .B(n637), .Z(n1000) );
  XNOR U1137 ( .A(n817), .B(n816), .Z(n651) );
  XNOR U1138 ( .A(n818), .B(n651), .Z(n1001) );
  XNOR U1139 ( .A(n1000), .B(n1001), .Z(n1002) );
  XOR U1140 ( .A(n1003), .B(n1002), .Z(n920) );
  XOR U1141 ( .A(n919), .B(n920), .Z(n792) );
  XNOR U1142 ( .A(n870), .B(n869), .Z(n664) );
  XNOR U1143 ( .A(n868), .B(n664), .Z(n959) );
  XNOR U1144 ( .A(n884), .B(n883), .Z(n886) );
  XNOR U1145 ( .A(n886), .B(n885), .Z(n958) );
  NANDN U1146 ( .A(n677), .B(n678), .Z(n683) );
  NOR U1147 ( .A(n679), .B(n678), .Z(n681) );
  OR U1148 ( .A(n681), .B(n680), .Z(n682) );
  NAND U1149 ( .A(n683), .B(n682), .Z(n957) );
  XOR U1150 ( .A(n958), .B(n957), .Z(n960) );
  XOR U1151 ( .A(n959), .B(n960), .Z(n927) );
  NANDN U1152 ( .A(n688), .B(oglobal[0]), .Z(n692) );
  OR U1153 ( .A(n690), .B(n689), .Z(n691) );
  AND U1154 ( .A(n692), .B(n691), .Z(n857) );
  XNOR U1155 ( .A(n857), .B(n856), .Z(n697) );
  XNOR U1156 ( .A(n858), .B(n697), .Z(n993) );
  OR U1157 ( .A(n702), .B(n701), .Z(n706) );
  OR U1158 ( .A(n704), .B(n703), .Z(n705) );
  NAND U1159 ( .A(n706), .B(n705), .Z(n905) );
  OR U1160 ( .A(n708), .B(n707), .Z(n712) );
  OR U1161 ( .A(n710), .B(n709), .Z(n711) );
  AND U1162 ( .A(n712), .B(n711), .Z(n904) );
  OR U1163 ( .A(n714), .B(n713), .Z(n718) );
  OR U1164 ( .A(n716), .B(n715), .Z(n717) );
  AND U1165 ( .A(n718), .B(n717), .Z(n903) );
  XNOR U1166 ( .A(n904), .B(n903), .Z(n719) );
  XOR U1167 ( .A(n905), .B(n719), .Z(n991) );
  XOR U1168 ( .A(n992), .B(n991), .Z(n994) );
  XOR U1169 ( .A(n993), .B(n994), .Z(n924) );
  XNOR U1170 ( .A(n875), .B(n874), .Z(n877) );
  XOR U1171 ( .A(n877), .B(n876), .Z(n951) );
  IV U1172 ( .A(n952), .Z(n950) );
  XNOR U1173 ( .A(n882), .B(n880), .Z(n747) );
  XNOR U1174 ( .A(n881), .B(n747), .Z(n953) );
  XNOR U1175 ( .A(n950), .B(n953), .Z(n748) );
  XNOR U1176 ( .A(n951), .B(n748), .Z(n925) );
  IV U1177 ( .A(n925), .Z(n923) );
  XOR U1178 ( .A(n924), .B(n923), .Z(n749) );
  XNOR U1179 ( .A(n927), .B(n749), .Z(n791) );
  XOR U1180 ( .A(n792), .B(n791), .Z(n794) );
  XNOR U1181 ( .A(n793), .B(n794), .Z(n1008) );
  XOR U1182 ( .A(n1007), .B(n1008), .Z(n750) );
  XOR U1183 ( .A(n1009), .B(n750), .Z(n1011) );
  XOR U1184 ( .A(n1010), .B(n1011), .Z(n1012) );
  NANDN U1185 ( .A(n752), .B(n751), .Z(n756) );
  NAND U1186 ( .A(n754), .B(n753), .Z(n755) );
  AND U1187 ( .A(n756), .B(n755), .Z(n1013) );
  XNOR U1188 ( .A(n1012), .B(n1013), .Z(o[1]) );
  NANDN U1189 ( .A(n757), .B(n758), .Z(n763) );
  NOR U1190 ( .A(n759), .B(n758), .Z(n761) );
  NANDN U1191 ( .A(n761), .B(n760), .Z(n762) );
  NAND U1192 ( .A(n763), .B(n762), .Z(n1132) );
  NAND U1193 ( .A(n765), .B(n764), .Z(n769) );
  NANDN U1194 ( .A(n767), .B(n766), .Z(n768) );
  NAND U1195 ( .A(n769), .B(n768), .Z(n1134) );
  NANDN U1196 ( .A(n771), .B(n770), .Z(n775) );
  NANDN U1197 ( .A(n773), .B(n772), .Z(n774) );
  AND U1198 ( .A(n775), .B(n774), .Z(n1109) );
  NAND U1199 ( .A(n777), .B(n776), .Z(n781) );
  NANDN U1200 ( .A(n779), .B(n778), .Z(n780) );
  AND U1201 ( .A(n781), .B(n780), .Z(n1107) );
  NANDN U1202 ( .A(n782), .B(n783), .Z(n788) );
  NOR U1203 ( .A(n784), .B(n783), .Z(n786) );
  NANDN U1204 ( .A(n786), .B(n785), .Z(n787) );
  AND U1205 ( .A(n788), .B(n787), .Z(n1108) );
  XNOR U1206 ( .A(n1107), .B(n1108), .Z(n789) );
  XNOR U1207 ( .A(n1109), .B(n789), .Z(n1133) );
  XOR U1208 ( .A(n1134), .B(n1133), .Z(n790) );
  XOR U1209 ( .A(n1132), .B(n790), .Z(n1016) );
  NANDN U1210 ( .A(n792), .B(n791), .Z(n796) );
  NANDN U1211 ( .A(n794), .B(n793), .Z(n795) );
  NAND U1212 ( .A(n796), .B(n795), .Z(n1125) );
  OR U1213 ( .A(n798), .B(n797), .Z(n802) );
  OR U1214 ( .A(n800), .B(n799), .Z(n801) );
  AND U1215 ( .A(n802), .B(n801), .Z(n1096) );
  XNOR U1216 ( .A(n1093), .B(n1094), .Z(n1095) );
  XNOR U1217 ( .A(n1096), .B(n1095), .Z(n1074) );
  NANDN U1218 ( .A(n811), .B(n810), .Z(n815) );
  NAND U1219 ( .A(n813), .B(n812), .Z(n814) );
  AND U1220 ( .A(n815), .B(n814), .Z(n1099) );
  XOR U1221 ( .A(n1097), .B(n1098), .Z(n1100) );
  XNOR U1222 ( .A(n1099), .B(n1100), .Z(n1073) );
  XOR U1223 ( .A(n1074), .B(n1073), .Z(n1075) );
  NANDN U1224 ( .A(n824), .B(n823), .Z(n828) );
  NANDN U1225 ( .A(n826), .B(n825), .Z(n827) );
  NAND U1226 ( .A(n828), .B(n827), .Z(n1058) );
  XOR U1227 ( .A(n1057), .B(oglobal[2]), .Z(n832) );
  XNOR U1228 ( .A(n1058), .B(n832), .Z(n1076) );
  XOR U1229 ( .A(n1075), .B(n1076), .Z(n1118) );
  NAND U1230 ( .A(n834), .B(n833), .Z(n838) );
  NAND U1231 ( .A(n836), .B(n835), .Z(n837) );
  AND U1232 ( .A(n838), .B(n837), .Z(n1066) );
  IV U1233 ( .A(n1066), .Z(n1067) );
  IV U1234 ( .A(n1068), .Z(n1065) );
  NANDN U1235 ( .A(n842), .B(n843), .Z(n848) );
  NOR U1236 ( .A(n844), .B(n843), .Z(n846) );
  OR U1237 ( .A(n846), .B(n845), .Z(n847) );
  NAND U1238 ( .A(n848), .B(n847), .Z(n1069) );
  XNOR U1239 ( .A(n1065), .B(n1069), .Z(n849) );
  XNOR U1240 ( .A(n1067), .B(n849), .Z(n1117) );
  NANDN U1241 ( .A(n851), .B(n850), .Z(n855) );
  NANDN U1242 ( .A(n853), .B(n852), .Z(n854) );
  NAND U1243 ( .A(n855), .B(n854), .Z(n1048) );
  XOR U1244 ( .A(n1048), .B(n1047), .Z(n1029) );
  NANDN U1245 ( .A(n863), .B(n862), .Z(n867) );
  NAND U1246 ( .A(n865), .B(n864), .Z(n866) );
  NAND U1247 ( .A(n867), .B(n866), .Z(n1053) );
  XOR U1248 ( .A(n1051), .B(n1052), .Z(n1054) );
  XNOR U1249 ( .A(n1053), .B(n1054), .Z(n1028) );
  XOR U1250 ( .A(n1029), .B(n1028), .Z(n1030) );
  OR U1251 ( .A(n875), .B(n874), .Z(n879) );
  OR U1252 ( .A(n877), .B(n876), .Z(n878) );
  NAND U1253 ( .A(n879), .B(n878), .Z(n1092) );
  OR U1254 ( .A(n884), .B(n883), .Z(n888) );
  OR U1255 ( .A(n886), .B(n885), .Z(n887) );
  AND U1256 ( .A(n888), .B(n887), .Z(n1090) );
  XNOR U1257 ( .A(n1089), .B(n1090), .Z(n1091) );
  XOR U1258 ( .A(n1092), .B(n1091), .Z(n1031) );
  XOR U1259 ( .A(n1030), .B(n1031), .Z(n1116) );
  XOR U1260 ( .A(n1117), .B(n1116), .Z(n1119) );
  XNOR U1261 ( .A(n1118), .B(n1119), .Z(n1129) );
  XNOR U1262 ( .A(n1022), .B(n1023), .Z(n1025) );
  NANDN U1263 ( .A(n898), .B(n897), .Z(n902) );
  NAND U1264 ( .A(n900), .B(n899), .Z(n901) );
  NAND U1265 ( .A(n902), .B(n901), .Z(n1088) );
  XNOR U1266 ( .A(n1085), .B(n1086), .Z(n1087) );
  XOR U1267 ( .A(n1088), .B(n1087), .Z(n1024) );
  XNOR U1268 ( .A(n1025), .B(n1024), .Z(n1112) );
  XNOR U1269 ( .A(n1111), .B(n1110), .Z(n1113) );
  XOR U1270 ( .A(n1112), .B(n1113), .Z(n1036) );
  NAND U1271 ( .A(n918), .B(n917), .Z(n922) );
  NAND U1272 ( .A(n920), .B(n919), .Z(n921) );
  AND U1273 ( .A(n922), .B(n921), .Z(n1037) );
  NANDN U1274 ( .A(n923), .B(n924), .Z(n929) );
  NOR U1275 ( .A(n925), .B(n924), .Z(n926) );
  OR U1276 ( .A(n927), .B(n926), .Z(n928) );
  NAND U1277 ( .A(n929), .B(n928), .Z(n1038) );
  XOR U1278 ( .A(n1037), .B(n1038), .Z(n930) );
  XNOR U1279 ( .A(n1036), .B(n930), .Z(n1128) );
  XNOR U1280 ( .A(n1129), .B(n1128), .Z(n1131) );
  NANDN U1281 ( .A(n932), .B(n931), .Z(n936) );
  NAND U1282 ( .A(n934), .B(n933), .Z(n935) );
  AND U1283 ( .A(n936), .B(n935), .Z(n1032) );
  NANDN U1284 ( .A(n938), .B(n937), .Z(n942) );
  NANDN U1285 ( .A(n940), .B(n939), .Z(n941) );
  NAND U1286 ( .A(n942), .B(n941), .Z(n1034) );
  NAND U1287 ( .A(n944), .B(n943), .Z(n948) );
  OR U1288 ( .A(n946), .B(n945), .Z(n947) );
  AND U1289 ( .A(n948), .B(n947), .Z(n1033) );
  XOR U1290 ( .A(n1034), .B(n1033), .Z(n949) );
  XNOR U1291 ( .A(n1032), .B(n949), .Z(n1061) );
  NANDN U1292 ( .A(n950), .B(n951), .Z(n956) );
  NOR U1293 ( .A(n952), .B(n951), .Z(n954) );
  OR U1294 ( .A(n954), .B(n953), .Z(n955) );
  NAND U1295 ( .A(n956), .B(n955), .Z(n1059) );
  NANDN U1296 ( .A(n958), .B(n957), .Z(n962) );
  NANDN U1297 ( .A(n960), .B(n959), .Z(n961) );
  AND U1298 ( .A(n962), .B(n961), .Z(n1060) );
  XOR U1299 ( .A(n1059), .B(n1060), .Z(n963) );
  XOR U1300 ( .A(n1061), .B(n963), .Z(n1039) );
  NANDN U1301 ( .A(n965), .B(n964), .Z(n971) );
  ANDN U1302 ( .B(n967), .A(n966), .Z(n969) );
  NANDN U1303 ( .A(n969), .B(n968), .Z(n970) );
  NAND U1304 ( .A(n971), .B(n970), .Z(n1062) );
  NANDN U1305 ( .A(n975), .B(n974), .Z(n979) );
  NANDN U1306 ( .A(n977), .B(n976), .Z(n978) );
  NAND U1307 ( .A(n979), .B(n978), .Z(n1079) );
  XNOR U1308 ( .A(n1080), .B(n1079), .Z(n1082) );
  XNOR U1309 ( .A(n1082), .B(n1081), .Z(n1063) );
  NANDN U1310 ( .A(n985), .B(n984), .Z(n989) );
  NANDN U1311 ( .A(n987), .B(n986), .Z(n988) );
  AND U1312 ( .A(n989), .B(n988), .Z(n1064) );
  XNOR U1313 ( .A(n1063), .B(n1064), .Z(n990) );
  XNOR U1314 ( .A(n1062), .B(n990), .Z(n1040) );
  XNOR U1315 ( .A(n1039), .B(n1040), .Z(n1041) );
  NANDN U1316 ( .A(n992), .B(n991), .Z(n996) );
  OR U1317 ( .A(n994), .B(n993), .Z(n995) );
  NAND U1318 ( .A(n996), .B(n995), .Z(n1105) );
  NANDN U1319 ( .A(n1001), .B(n1000), .Z(n1005) );
  NAND U1320 ( .A(n1003), .B(n1002), .Z(n1004) );
  AND U1321 ( .A(n1005), .B(n1004), .Z(n1104) );
  XNOR U1322 ( .A(n1103), .B(n1104), .Z(n1006) );
  XOR U1323 ( .A(n1105), .B(n1006), .Z(n1042) );
  XNOR U1324 ( .A(n1041), .B(n1042), .Z(n1130) );
  XNOR U1325 ( .A(n1131), .B(n1130), .Z(n1123) );
  XOR U1326 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U1327 ( .A(n1125), .B(n1124), .Z(n1017) );
  XOR U1328 ( .A(n1016), .B(n1017), .Z(n1019) );
  NAND U1329 ( .A(n1011), .B(n1010), .Z(n1015) );
  NANDN U1330 ( .A(n1013), .B(n1012), .Z(n1014) );
  AND U1331 ( .A(n1015), .B(n1014), .Z(n1018) );
  XOR U1332 ( .A(n1019), .B(n1018), .Z(o[2]) );
  NANDN U1333 ( .A(n1017), .B(n1016), .Z(n1021) );
  OR U1334 ( .A(n1019), .B(n1018), .Z(n1020) );
  NAND U1335 ( .A(n1021), .B(n1020), .Z(n1192) );
  OR U1336 ( .A(n1023), .B(n1022), .Z(n1027) );
  NANDN U1337 ( .A(n1025), .B(n1024), .Z(n1026) );
  AND U1338 ( .A(n1027), .B(n1026), .Z(n1139) );
  XOR U1339 ( .A(n1141), .B(n1140), .Z(n1035) );
  XNOR U1340 ( .A(n1139), .B(n1035), .Z(n1188) );
  NANDN U1341 ( .A(n1040), .B(n1039), .Z(n1044) );
  NAND U1342 ( .A(n1042), .B(n1041), .Z(n1043) );
  NAND U1343 ( .A(n1044), .B(n1043), .Z(n1186) );
  XNOR U1344 ( .A(n1185), .B(n1186), .Z(n1187) );
  XOR U1345 ( .A(n1188), .B(n1187), .Z(n1182) );
  NANDN U1346 ( .A(n1046), .B(n1045), .Z(n1050) );
  NAND U1347 ( .A(n1048), .B(n1047), .Z(n1049) );
  AND U1348 ( .A(n1050), .B(n1049), .Z(n1158) );
  NAND U1349 ( .A(n1052), .B(n1051), .Z(n1056) );
  NAND U1350 ( .A(n1054), .B(n1053), .Z(n1055) );
  AND U1351 ( .A(n1056), .B(n1055), .Z(n1148) );
  XOR U1352 ( .A(oglobal[3]), .B(n1148), .Z(n1155) );
  XNOR U1353 ( .A(n1155), .B(n1156), .Z(n1157) );
  XOR U1354 ( .A(n1158), .B(n1157), .Z(n1174) );
  XNOR U1355 ( .A(n1171), .B(n1172), .Z(n1173) );
  XNOR U1356 ( .A(n1174), .B(n1173), .Z(n1160) );
  NANDN U1357 ( .A(n1066), .B(n1065), .Z(n1072) );
  ANDN U1358 ( .B(n1068), .A(n1067), .Z(n1070) );
  NANDN U1359 ( .A(n1070), .B(n1069), .Z(n1071) );
  NAND U1360 ( .A(n1072), .B(n1071), .Z(n1159) );
  XOR U1361 ( .A(n1160), .B(n1159), .Z(n1162) );
  OR U1362 ( .A(n1074), .B(n1073), .Z(n1078) );
  NAND U1363 ( .A(n1076), .B(n1075), .Z(n1077) );
  AND U1364 ( .A(n1078), .B(n1077), .Z(n1165) );
  OR U1365 ( .A(n1080), .B(n1079), .Z(n1084) );
  OR U1366 ( .A(n1082), .B(n1081), .Z(n1083) );
  NAND U1367 ( .A(n1084), .B(n1083), .Z(n1152) );
  XNOR U1368 ( .A(n1150), .B(n1149), .Z(n1151) );
  XOR U1369 ( .A(n1152), .B(n1151), .Z(n1144) );
  NANDN U1370 ( .A(n1098), .B(n1097), .Z(n1102) );
  OR U1371 ( .A(n1100), .B(n1099), .Z(n1101) );
  AND U1372 ( .A(n1102), .B(n1101), .Z(n1142) );
  XNOR U1373 ( .A(n1143), .B(n1142), .Z(n1145) );
  XNOR U1374 ( .A(n1144), .B(n1145), .Z(n1167) );
  XNOR U1375 ( .A(n1167), .B(n1166), .Z(n1106) );
  XNOR U1376 ( .A(n1165), .B(n1106), .Z(n1161) );
  XNOR U1377 ( .A(n1162), .B(n1161), .Z(n1179) );
  NAND U1378 ( .A(n1111), .B(n1110), .Z(n1115) );
  NANDN U1379 ( .A(n1113), .B(n1112), .Z(n1114) );
  NAND U1380 ( .A(n1115), .B(n1114), .Z(n1170) );
  XOR U1381 ( .A(n1170), .B(n1169), .Z(n1120) );
  XOR U1382 ( .A(n1168), .B(n1120), .Z(n1180) );
  IV U1383 ( .A(n1180), .Z(n1178) );
  XNOR U1384 ( .A(n1179), .B(n1178), .Z(n1121) );
  XNOR U1385 ( .A(n1182), .B(n1121), .Z(n1193) );
  XNOR U1386 ( .A(n1192), .B(n1193), .Z(n1194) );
  NAND U1387 ( .A(n1123), .B(n1122), .Z(n1127) );
  NAND U1388 ( .A(n1125), .B(n1124), .Z(n1126) );
  AND U1389 ( .A(n1127), .B(n1126), .Z(n1138) );
  XNOR U1390 ( .A(n1136), .B(n1137), .Z(n1135) );
  XNOR U1391 ( .A(n1138), .B(n1135), .Z(n1195) );
  XNOR U1392 ( .A(n1194), .B(n1195), .Z(o[3]) );
  OR U1393 ( .A(n1143), .B(n1142), .Z(n1147) );
  NANDN U1394 ( .A(n1145), .B(n1144), .Z(n1146) );
  AND U1395 ( .A(n1147), .B(n1146), .Z(n1203) );
  XOR U1396 ( .A(n1202), .B(n1203), .Z(n1205) );
  ANDN U1397 ( .B(oglobal[3]), .A(n1148), .Z(n1201) );
  XOR U1398 ( .A(oglobal[4]), .B(n1201), .Z(n1211) );
  OR U1399 ( .A(n1150), .B(n1149), .Z(n1154) );
  OR U1400 ( .A(n1152), .B(n1151), .Z(n1153) );
  AND U1401 ( .A(n1154), .B(n1153), .Z(n1209) );
  XNOR U1402 ( .A(n1209), .B(n1208), .Z(n1210) );
  XNOR U1403 ( .A(n1211), .B(n1210), .Z(n1204) );
  XNOR U1404 ( .A(n1205), .B(n1204), .Z(n1217) );
  NANDN U1405 ( .A(n1160), .B(n1159), .Z(n1164) );
  NANDN U1406 ( .A(n1162), .B(n1161), .Z(n1163) );
  NAND U1407 ( .A(n1164), .B(n1163), .Z(n1214) );
  NAND U1408 ( .A(n1172), .B(n1171), .Z(n1176) );
  OR U1409 ( .A(n1174), .B(n1173), .Z(n1175) );
  AND U1410 ( .A(n1176), .B(n1175), .Z(n1220) );
  IV U1411 ( .A(n1220), .Z(n1222) );
  XNOR U1412 ( .A(n1223), .B(n1222), .Z(n1177) );
  XOR U1413 ( .A(n1221), .B(n1177), .Z(n1215) );
  XOR U1414 ( .A(n1214), .B(n1215), .Z(n1216) );
  XNOR U1415 ( .A(n1217), .B(n1216), .Z(n1200) );
  NANDN U1416 ( .A(n1178), .B(n1179), .Z(n1184) );
  NOR U1417 ( .A(n1180), .B(n1179), .Z(n1181) );
  OR U1418 ( .A(n1182), .B(n1181), .Z(n1183) );
  AND U1419 ( .A(n1184), .B(n1183), .Z(n1198) );
  NANDN U1420 ( .A(n1186), .B(n1185), .Z(n1190) );
  NAND U1421 ( .A(n1188), .B(n1187), .Z(n1189) );
  AND U1422 ( .A(n1190), .B(n1189), .Z(n1199) );
  XNOR U1423 ( .A(n1198), .B(n1199), .Z(n1191) );
  XOR U1424 ( .A(n1200), .B(n1191), .Z(n1229) );
  XOR U1425 ( .A(n1228), .B(n1229), .Z(n1230) );
  NANDN U1426 ( .A(n1193), .B(n1192), .Z(n1197) );
  NANDN U1427 ( .A(n1195), .B(n1194), .Z(n1196) );
  AND U1428 ( .A(n1197), .B(n1196), .Z(n1231) );
  XNOR U1429 ( .A(n1230), .B(n1231), .Z(o[4]) );
  NAND U1430 ( .A(n1201), .B(oglobal[4]), .Z(n1234) );
  XOR U1431 ( .A(oglobal[5]), .B(n1234), .Z(n1237) );
  NANDN U1432 ( .A(n1203), .B(n1202), .Z(n1207) );
  OR U1433 ( .A(n1205), .B(n1204), .Z(n1206) );
  AND U1434 ( .A(n1207), .B(n1206), .Z(n1236) );
  OR U1435 ( .A(n1209), .B(n1208), .Z(n1213) );
  OR U1436 ( .A(n1211), .B(n1210), .Z(n1212) );
  AND U1437 ( .A(n1213), .B(n1212), .Z(n1235) );
  XNOR U1438 ( .A(n1236), .B(n1235), .Z(n1238) );
  XNOR U1439 ( .A(n1237), .B(n1238), .Z(n1249) );
  NANDN U1440 ( .A(n1215), .B(n1214), .Z(n1219) );
  OR U1441 ( .A(n1217), .B(n1216), .Z(n1218) );
  NAND U1442 ( .A(n1219), .B(n1218), .Z(n1251) );
  NANDN U1443 ( .A(n1220), .B(n1221), .Z(n1226) );
  NOR U1444 ( .A(n1222), .B(n1221), .Z(n1224) );
  NANDN U1445 ( .A(n1224), .B(n1223), .Z(n1225) );
  AND U1446 ( .A(n1226), .B(n1225), .Z(n1248) );
  IV U1447 ( .A(n1248), .Z(n1247) );
  XNOR U1448 ( .A(n1251), .B(n1247), .Z(n1227) );
  XOR U1449 ( .A(n1249), .B(n1227), .Z(n1242) );
  XOR U1450 ( .A(n1241), .B(n1242), .Z(n1243) );
  NAND U1451 ( .A(n1229), .B(n1228), .Z(n1233) );
  NANDN U1452 ( .A(n1231), .B(n1230), .Z(n1232) );
  AND U1453 ( .A(n1233), .B(n1232), .Z(n1244) );
  XNOR U1454 ( .A(n1243), .B(n1244), .Z(o[5]) );
  NANDN U1455 ( .A(n1234), .B(oglobal[5]), .Z(n1260) );
  XOR U1456 ( .A(oglobal[6]), .B(n1260), .Z(n1262) );
  OR U1457 ( .A(n1236), .B(n1235), .Z(n1240) );
  NANDN U1458 ( .A(n1238), .B(n1237), .Z(n1239) );
  NAND U1459 ( .A(n1240), .B(n1239), .Z(n1261) );
  XOR U1460 ( .A(n1262), .B(n1261), .Z(n1255) );
  NAND U1461 ( .A(n1242), .B(n1241), .Z(n1246) );
  NANDN U1462 ( .A(n1244), .B(n1243), .Z(n1245) );
  NAND U1463 ( .A(n1246), .B(n1245), .Z(n1257) );
  OR U1464 ( .A(n1249), .B(n1247), .Z(n1253) );
  ANDN U1465 ( .B(n1249), .A(n1248), .Z(n1250) );
  OR U1466 ( .A(n1251), .B(n1250), .Z(n1252) );
  NAND U1467 ( .A(n1253), .B(n1252), .Z(n1256) );
  XOR U1468 ( .A(n1257), .B(n1256), .Z(n1254) );
  XOR U1469 ( .A(n1255), .B(n1254), .Z(o[6]) );
  NANDN U1470 ( .A(n1255), .B(n1254), .Z(n1259) );
  OR U1471 ( .A(n1257), .B(n1256), .Z(n1258) );
  AND U1472 ( .A(n1259), .B(n1258), .Z(n1265) );
  XNOR U1473 ( .A(n1265), .B(oglobal[7]), .Z(n1267) );
  NANDN U1474 ( .A(n1260), .B(oglobal[6]), .Z(n1264) );
  OR U1475 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U1476 ( .A(n1264), .B(n1263), .Z(n1266) );
  XOR U1477 ( .A(n1267), .B(n1266), .Z(o[7]) );
  NAND U1478 ( .A(n1265), .B(oglobal[7]), .Z(n1269) );
  OR U1479 ( .A(n1267), .B(n1266), .Z(n1268) );
  AND U1480 ( .A(n1269), .B(n1268), .Z(n1270) );
  XNOR U1481 ( .A(oglobal[8]), .B(n1270), .Z(o[8]) );
  NANDN U1482 ( .A(n1270), .B(oglobal[8]), .Z(n1271) );
  XNOR U1483 ( .A(oglobal[9]), .B(n1271), .Z(o[9]) );
  NANDN U1484 ( .A(n1271), .B(oglobal[9]), .Z(n1272) );
  XNOR U1485 ( .A(oglobal[10]), .B(n1272), .Z(o[10]) );
endmodule

