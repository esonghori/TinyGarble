
module sum_N1024_CC2 ( clk, rst, a, b, c );
  input [511:0] a;
  input [511:0] b;
  output [511:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[1]), .B(n2043), .Z(n1341) );
  XOR U4 ( .A(a[4]), .B(n2034), .Z(n108) );
  XOR U5 ( .A(a[7]), .B(n2025), .Z(n27) );
  XOR U6 ( .A(a[10]), .B(n2016), .Z(n1711) );
  XOR U7 ( .A(a[13]), .B(n2007), .Z(n1588) );
  XOR U8 ( .A(a[16]), .B(n1998), .Z(n1465) );
  XOR U9 ( .A(a[19]), .B(n1989), .Z(n1342) );
  XOR U10 ( .A(a[22]), .B(n1980), .Z(n1218) );
  XOR U11 ( .A(a[25]), .B(n1971), .Z(n1095) );
  XOR U12 ( .A(a[28]), .B(n1962), .Z(n972) );
  XOR U13 ( .A(a[31]), .B(n1953), .Z(n848) );
  XOR U14 ( .A(a[34]), .B(n1944), .Z(n725) );
  XOR U15 ( .A(a[37]), .B(n1935), .Z(n602) );
  XOR U16 ( .A(a[40]), .B(n1926), .Z(n478) );
  XOR U17 ( .A(a[43]), .B(n1917), .Z(n355) );
  XOR U18 ( .A(a[46]), .B(n1908), .Z(n232) );
  XOR U19 ( .A(a[49]), .B(n1899), .Z(n109) );
  XOR U20 ( .A(a[52]), .B(n1890), .Z(n57) );
  XOR U21 ( .A(a[55]), .B(n1881), .Z(n54) );
  XOR U22 ( .A(a[58]), .B(n1872), .Z(n51) );
  XOR U23 ( .A(a[61]), .B(n1863), .Z(n47) );
  XOR U24 ( .A(a[64]), .B(n1854), .Z(n44) );
  XOR U25 ( .A(a[67]), .B(n1845), .Z(n41) );
  XOR U26 ( .A(a[70]), .B(n1836), .Z(n37) );
  XOR U27 ( .A(a[73]), .B(n1827), .Z(n34) );
  XOR U28 ( .A(a[76]), .B(n1818), .Z(n31) );
  XOR U29 ( .A(a[79]), .B(n1809), .Z(n28) );
  XOR U30 ( .A(a[82]), .B(n1800), .Z(n24) );
  XOR U31 ( .A(a[85]), .B(n1791), .Z(n21) );
  XOR U32 ( .A(a[88]), .B(n1782), .Z(n18) );
  XOR U33 ( .A(a[91]), .B(n1773), .Z(n14) );
  XOR U34 ( .A(a[94]), .B(n1764), .Z(n11) );
  XOR U35 ( .A(a[97]), .B(n1755), .Z(n8) );
  XOR U36 ( .A(a[100]), .B(n1745), .Z(n1747) );
  XOR U37 ( .A(a[103]), .B(n1733), .Z(n1735) );
  XOR U38 ( .A(a[106]), .B(n1721), .Z(n1723) );
  XOR U39 ( .A(a[109]), .B(n1708), .Z(n1710) );
  XOR U40 ( .A(a[112]), .B(n1696), .Z(n1698) );
  XOR U41 ( .A(a[115]), .B(n1684), .Z(n1686) );
  XOR U42 ( .A(a[118]), .B(n1672), .Z(n1674) );
  XOR U43 ( .A(a[121]), .B(n1659), .Z(n1661) );
  XOR U44 ( .A(a[124]), .B(n1647), .Z(n1649) );
  XOR U45 ( .A(a[127]), .B(n1635), .Z(n1637) );
  XOR U46 ( .A(a[130]), .B(n1622), .Z(n1624) );
  XOR U47 ( .A(a[133]), .B(n1610), .Z(n1612) );
  XOR U48 ( .A(a[136]), .B(n1598), .Z(n1600) );
  XOR U49 ( .A(a[139]), .B(n1585), .Z(n1587) );
  XOR U50 ( .A(a[142]), .B(n1573), .Z(n1575) );
  XOR U51 ( .A(a[145]), .B(n1561), .Z(n1563) );
  XOR U52 ( .A(a[148]), .B(n1549), .Z(n1551) );
  XOR U53 ( .A(a[151]), .B(n1536), .Z(n1538) );
  XOR U54 ( .A(a[154]), .B(n1524), .Z(n1526) );
  XOR U55 ( .A(a[157]), .B(n1512), .Z(n1514) );
  XOR U56 ( .A(a[160]), .B(n1499), .Z(n1501) );
  XOR U57 ( .A(a[163]), .B(n1487), .Z(n1489) );
  XOR U58 ( .A(a[166]), .B(n1475), .Z(n1477) );
  XOR U59 ( .A(a[169]), .B(n1462), .Z(n1464) );
  XOR U60 ( .A(a[172]), .B(n1450), .Z(n1452) );
  XOR U61 ( .A(a[175]), .B(n1438), .Z(n1440) );
  XOR U62 ( .A(a[178]), .B(n1426), .Z(n1428) );
  XOR U63 ( .A(a[181]), .B(n1413), .Z(n1415) );
  XOR U64 ( .A(a[184]), .B(n1401), .Z(n1403) );
  XOR U65 ( .A(a[187]), .B(n1389), .Z(n1391) );
  XOR U66 ( .A(a[190]), .B(n1376), .Z(n1378) );
  XOR U67 ( .A(a[193]), .B(n1364), .Z(n1366) );
  XOR U68 ( .A(a[196]), .B(n1352), .Z(n1354) );
  XOR U69 ( .A(a[199]), .B(n1338), .Z(n1340) );
  XOR U70 ( .A(a[202]), .B(n1326), .Z(n1328) );
  XOR U71 ( .A(a[205]), .B(n1314), .Z(n1316) );
  XOR U72 ( .A(a[208]), .B(n1302), .Z(n1304) );
  XOR U73 ( .A(a[211]), .B(n1289), .Z(n1291) );
  XOR U74 ( .A(a[214]), .B(n1277), .Z(n1279) );
  XOR U75 ( .A(a[217]), .B(n1265), .Z(n1267) );
  XOR U76 ( .A(a[220]), .B(n1252), .Z(n1254) );
  XOR U77 ( .A(a[223]), .B(n1240), .Z(n1242) );
  XOR U78 ( .A(a[226]), .B(n1228), .Z(n1230) );
  XOR U79 ( .A(a[229]), .B(n1215), .Z(n1217) );
  XOR U80 ( .A(a[232]), .B(n1203), .Z(n1205) );
  XOR U81 ( .A(a[235]), .B(n1191), .Z(n1193) );
  XOR U82 ( .A(a[238]), .B(n1179), .Z(n1181) );
  XOR U83 ( .A(a[241]), .B(n1166), .Z(n1168) );
  XOR U84 ( .A(a[244]), .B(n1154), .Z(n1156) );
  XOR U85 ( .A(a[247]), .B(n1142), .Z(n1144) );
  XOR U86 ( .A(a[250]), .B(n1129), .Z(n1131) );
  XOR U87 ( .A(a[253]), .B(n1117), .Z(n1119) );
  XOR U88 ( .A(a[256]), .B(n1105), .Z(n1107) );
  XOR U89 ( .A(a[259]), .B(n1092), .Z(n1094) );
  XOR U90 ( .A(a[262]), .B(n1080), .Z(n1082) );
  XOR U91 ( .A(a[265]), .B(n1068), .Z(n1070) );
  XOR U92 ( .A(a[268]), .B(n1056), .Z(n1058) );
  XOR U93 ( .A(a[271]), .B(n1043), .Z(n1045) );
  XOR U94 ( .A(a[274]), .B(n1031), .Z(n1033) );
  XOR U95 ( .A(a[277]), .B(n1019), .Z(n1021) );
  XOR U96 ( .A(a[280]), .B(n1006), .Z(n1008) );
  XOR U97 ( .A(a[283]), .B(n994), .Z(n996) );
  XOR U98 ( .A(a[286]), .B(n982), .Z(n984) );
  XOR U99 ( .A(a[289]), .B(n969), .Z(n971) );
  XOR U100 ( .A(a[292]), .B(n957), .Z(n959) );
  XOR U101 ( .A(a[295]), .B(n945), .Z(n947) );
  XOR U102 ( .A(a[298]), .B(n933), .Z(n935) );
  XOR U103 ( .A(a[301]), .B(n919), .Z(n921) );
  XOR U104 ( .A(a[304]), .B(n907), .Z(n909) );
  XOR U105 ( .A(a[307]), .B(n895), .Z(n897) );
  XOR U106 ( .A(a[310]), .B(n882), .Z(n884) );
  XOR U107 ( .A(a[313]), .B(n870), .Z(n872) );
  XOR U108 ( .A(a[316]), .B(n858), .Z(n860) );
  XOR U109 ( .A(a[319]), .B(n845), .Z(n847) );
  XOR U110 ( .A(a[322]), .B(n833), .Z(n835) );
  XOR U111 ( .A(a[325]), .B(n821), .Z(n823) );
  XOR U112 ( .A(a[328]), .B(n809), .Z(n811) );
  XOR U113 ( .A(a[331]), .B(n796), .Z(n798) );
  XOR U114 ( .A(a[334]), .B(n784), .Z(n786) );
  XOR U115 ( .A(a[337]), .B(n772), .Z(n774) );
  XOR U116 ( .A(a[340]), .B(n759), .Z(n761) );
  XOR U117 ( .A(a[343]), .B(n747), .Z(n749) );
  XOR U118 ( .A(a[346]), .B(n735), .Z(n737) );
  XOR U119 ( .A(a[349]), .B(n722), .Z(n724) );
  XOR U120 ( .A(a[352]), .B(n710), .Z(n712) );
  XOR U121 ( .A(a[355]), .B(n698), .Z(n700) );
  XOR U122 ( .A(a[358]), .B(n686), .Z(n688) );
  XOR U123 ( .A(a[361]), .B(n673), .Z(n675) );
  XOR U124 ( .A(a[364]), .B(n661), .Z(n663) );
  XOR U125 ( .A(a[367]), .B(n649), .Z(n651) );
  XOR U126 ( .A(a[370]), .B(n636), .Z(n638) );
  XOR U127 ( .A(a[373]), .B(n624), .Z(n626) );
  XOR U128 ( .A(a[376]), .B(n612), .Z(n614) );
  XOR U129 ( .A(a[379]), .B(n599), .Z(n601) );
  XOR U130 ( .A(a[382]), .B(n587), .Z(n589) );
  XOR U131 ( .A(a[385]), .B(n575), .Z(n577) );
  XOR U132 ( .A(a[388]), .B(n563), .Z(n565) );
  XOR U133 ( .A(a[391]), .B(n550), .Z(n552) );
  XOR U134 ( .A(a[394]), .B(n538), .Z(n540) );
  XOR U135 ( .A(a[397]), .B(n526), .Z(n528) );
  XOR U136 ( .A(a[400]), .B(n512), .Z(n514) );
  XOR U137 ( .A(a[403]), .B(n500), .Z(n502) );
  XOR U138 ( .A(a[406]), .B(n488), .Z(n490) );
  XOR U139 ( .A(a[409]), .B(n475), .Z(n477) );
  XOR U140 ( .A(a[412]), .B(n463), .Z(n465) );
  XOR U141 ( .A(a[415]), .B(n451), .Z(n453) );
  XOR U142 ( .A(a[418]), .B(n439), .Z(n441) );
  XOR U143 ( .A(a[421]), .B(n426), .Z(n428) );
  XOR U144 ( .A(a[424]), .B(n414), .Z(n416) );
  XOR U145 ( .A(a[427]), .B(n402), .Z(n404) );
  XOR U146 ( .A(a[430]), .B(n389), .Z(n391) );
  XOR U147 ( .A(a[433]), .B(n377), .Z(n379) );
  XOR U148 ( .A(a[436]), .B(n365), .Z(n367) );
  XOR U149 ( .A(a[439]), .B(n352), .Z(n354) );
  XOR U150 ( .A(a[442]), .B(n340), .Z(n342) );
  XOR U151 ( .A(a[445]), .B(n328), .Z(n330) );
  XOR U152 ( .A(a[448]), .B(n316), .Z(n318) );
  XOR U153 ( .A(a[451]), .B(n303), .Z(n305) );
  XOR U154 ( .A(a[454]), .B(n291), .Z(n293) );
  XOR U155 ( .A(a[457]), .B(n279), .Z(n281) );
  XOR U156 ( .A(a[460]), .B(n266), .Z(n268) );
  XOR U157 ( .A(a[463]), .B(n254), .Z(n256) );
  XOR U158 ( .A(a[466]), .B(n242), .Z(n244) );
  XOR U159 ( .A(a[469]), .B(n229), .Z(n231) );
  XOR U160 ( .A(a[472]), .B(n217), .Z(n219) );
  XOR U161 ( .A(a[475]), .B(n205), .Z(n207) );
  XOR U162 ( .A(a[478]), .B(n193), .Z(n195) );
  XOR U163 ( .A(a[481]), .B(n180), .Z(n182) );
  XOR U164 ( .A(a[484]), .B(n168), .Z(n170) );
  XOR U165 ( .A(a[487]), .B(n156), .Z(n158) );
  XOR U166 ( .A(a[490]), .B(n143), .Z(n145) );
  XOR U167 ( .A(a[493]), .B(n131), .Z(n133) );
  XOR U168 ( .A(a[496]), .B(n119), .Z(n121) );
  XOR U169 ( .A(a[499]), .B(n105), .Z(n107) );
  XOR U170 ( .A(a[502]), .B(n93), .Z(n95) );
  XOR U171 ( .A(a[505]), .B(n81), .Z(n83) );
  XOR U172 ( .A(a[508]), .B(n69), .Z(n71) );
  XOR U173 ( .A(a[2]), .B(n2040), .Z(n930) );
  XOR U174 ( .A(a[5]), .B(n2031), .Z(n49) );
  XOR U175 ( .A(a[8]), .B(n2022), .Z(n16) );
  XOR U176 ( .A(a[11]), .B(n2013), .Z(n1670) );
  XOR U177 ( .A(a[14]), .B(n2004), .Z(n1547) );
  XOR U178 ( .A(a[17]), .B(n1995), .Z(n1424) );
  XOR U179 ( .A(a[20]), .B(n1986), .Z(n1300) );
  XOR U180 ( .A(a[23]), .B(n1977), .Z(n1177) );
  XOR U181 ( .A(a[26]), .B(n1968), .Z(n1054) );
  XOR U182 ( .A(a[29]), .B(n1959), .Z(n931) );
  XOR U183 ( .A(a[32]), .B(n1950), .Z(n807) );
  XOR U184 ( .A(a[35]), .B(n1941), .Z(n684) );
  XOR U185 ( .A(a[38]), .B(n1932), .Z(n561) );
  XOR U186 ( .A(a[41]), .B(n1923), .Z(n437) );
  XOR U187 ( .A(a[44]), .B(n1914), .Z(n314) );
  XOR U188 ( .A(a[47]), .B(n1905), .Z(n191) );
  XOR U189 ( .A(a[50]), .B(n1896), .Z(n67) );
  XOR U190 ( .A(a[53]), .B(n1887), .Z(n56) );
  XOR U191 ( .A(a[56]), .B(n1878), .Z(n53) );
  XOR U192 ( .A(a[59]), .B(n1869), .Z(n50) );
  XOR U193 ( .A(a[62]), .B(n1860), .Z(n46) );
  XOR U194 ( .A(a[65]), .B(n1851), .Z(n43) );
  XOR U195 ( .A(a[68]), .B(n1842), .Z(n40) );
  XOR U196 ( .A(a[71]), .B(n1833), .Z(n36) );
  XOR U197 ( .A(a[74]), .B(n1824), .Z(n33) );
  XOR U198 ( .A(a[77]), .B(n1815), .Z(n30) );
  XOR U199 ( .A(a[80]), .B(n1806), .Z(n26) );
  XOR U200 ( .A(a[83]), .B(n1797), .Z(n23) );
  XOR U201 ( .A(a[86]), .B(n1788), .Z(n20) );
  XOR U202 ( .A(a[89]), .B(n1779), .Z(n17) );
  XOR U203 ( .A(a[92]), .B(n1770), .Z(n13) );
  XOR U204 ( .A(a[95]), .B(n1761), .Z(n10) );
  XOR U205 ( .A(a[98]), .B(n1752), .Z(n7) );
  XOR U206 ( .A(a[101]), .B(n1741), .Z(n1743) );
  XOR U207 ( .A(a[104]), .B(n1729), .Z(n1731) );
  XOR U208 ( .A(a[107]), .B(n1717), .Z(n1719) );
  XOR U209 ( .A(a[110]), .B(n1704), .Z(n1706) );
  XOR U210 ( .A(a[113]), .B(n1692), .Z(n1694) );
  XOR U211 ( .A(a[116]), .B(n1680), .Z(n1682) );
  XOR U212 ( .A(a[119]), .B(n1667), .Z(n1669) );
  XOR U213 ( .A(a[122]), .B(n1655), .Z(n1657) );
  XOR U214 ( .A(a[125]), .B(n1643), .Z(n1645) );
  XOR U215 ( .A(a[128]), .B(n1631), .Z(n1633) );
  XOR U216 ( .A(a[131]), .B(n1618), .Z(n1620) );
  XOR U217 ( .A(a[134]), .B(n1606), .Z(n1608) );
  XOR U218 ( .A(a[137]), .B(n1594), .Z(n1596) );
  XOR U219 ( .A(a[140]), .B(n1581), .Z(n1583) );
  XOR U220 ( .A(a[143]), .B(n1569), .Z(n1571) );
  XOR U221 ( .A(a[146]), .B(n1557), .Z(n1559) );
  XOR U222 ( .A(a[149]), .B(n1544), .Z(n1546) );
  XOR U223 ( .A(a[152]), .B(n1532), .Z(n1534) );
  XOR U224 ( .A(a[155]), .B(n1520), .Z(n1522) );
  XOR U225 ( .A(a[158]), .B(n1508), .Z(n1510) );
  XOR U226 ( .A(a[161]), .B(n1495), .Z(n1497) );
  XOR U227 ( .A(a[164]), .B(n1483), .Z(n1485) );
  XOR U228 ( .A(a[167]), .B(n1471), .Z(n1473) );
  XOR U229 ( .A(a[170]), .B(n1458), .Z(n1460) );
  XOR U230 ( .A(a[173]), .B(n1446), .Z(n1448) );
  XOR U231 ( .A(a[176]), .B(n1434), .Z(n1436) );
  XOR U232 ( .A(a[179]), .B(n1421), .Z(n1423) );
  XOR U233 ( .A(a[182]), .B(n1409), .Z(n1411) );
  XOR U234 ( .A(a[185]), .B(n1397), .Z(n1399) );
  XOR U235 ( .A(a[188]), .B(n1385), .Z(n1387) );
  XOR U236 ( .A(a[191]), .B(n1372), .Z(n1374) );
  XOR U237 ( .A(a[194]), .B(n1360), .Z(n1362) );
  XOR U238 ( .A(a[197]), .B(n1348), .Z(n1350) );
  XOR U239 ( .A(a[200]), .B(n1334), .Z(n1336) );
  XOR U240 ( .A(a[203]), .B(n1322), .Z(n1324) );
  XOR U241 ( .A(a[206]), .B(n1310), .Z(n1312) );
  XOR U242 ( .A(a[209]), .B(n1297), .Z(n1299) );
  XOR U243 ( .A(a[212]), .B(n1285), .Z(n1287) );
  XOR U244 ( .A(a[215]), .B(n1273), .Z(n1275) );
  XOR U245 ( .A(a[218]), .B(n1261), .Z(n1263) );
  XOR U246 ( .A(a[221]), .B(n1248), .Z(n1250) );
  XOR U247 ( .A(a[224]), .B(n1236), .Z(n1238) );
  XOR U248 ( .A(a[227]), .B(n1224), .Z(n1226) );
  XOR U249 ( .A(a[230]), .B(n1211), .Z(n1213) );
  XOR U250 ( .A(a[233]), .B(n1199), .Z(n1201) );
  XOR U251 ( .A(a[236]), .B(n1187), .Z(n1189) );
  XOR U252 ( .A(a[239]), .B(n1174), .Z(n1176) );
  XOR U253 ( .A(a[242]), .B(n1162), .Z(n1164) );
  XOR U254 ( .A(a[245]), .B(n1150), .Z(n1152) );
  XOR U255 ( .A(a[248]), .B(n1138), .Z(n1140) );
  XOR U256 ( .A(a[251]), .B(n1125), .Z(n1127) );
  XOR U257 ( .A(a[254]), .B(n1113), .Z(n1115) );
  XOR U258 ( .A(a[257]), .B(n1101), .Z(n1103) );
  XOR U259 ( .A(a[260]), .B(n1088), .Z(n1090) );
  XOR U260 ( .A(a[263]), .B(n1076), .Z(n1078) );
  XOR U261 ( .A(a[266]), .B(n1064), .Z(n1066) );
  XOR U262 ( .A(a[269]), .B(n1051), .Z(n1053) );
  XOR U263 ( .A(a[272]), .B(n1039), .Z(n1041) );
  XOR U264 ( .A(a[275]), .B(n1027), .Z(n1029) );
  XOR U265 ( .A(a[278]), .B(n1015), .Z(n1017) );
  XOR U266 ( .A(a[281]), .B(n1002), .Z(n1004) );
  XOR U267 ( .A(a[284]), .B(n990), .Z(n992) );
  XOR U268 ( .A(a[287]), .B(n978), .Z(n980) );
  XOR U269 ( .A(a[290]), .B(n965), .Z(n967) );
  XOR U270 ( .A(a[293]), .B(n953), .Z(n955) );
  XOR U271 ( .A(a[296]), .B(n941), .Z(n943) );
  XOR U272 ( .A(a[299]), .B(n927), .Z(n929) );
  XOR U273 ( .A(a[302]), .B(n915), .Z(n917) );
  XOR U274 ( .A(a[305]), .B(n903), .Z(n905) );
  XOR U275 ( .A(a[308]), .B(n891), .Z(n893) );
  XOR U276 ( .A(a[311]), .B(n878), .Z(n880) );
  XOR U277 ( .A(a[314]), .B(n866), .Z(n868) );
  XOR U278 ( .A(a[317]), .B(n854), .Z(n856) );
  XOR U279 ( .A(a[320]), .B(n841), .Z(n843) );
  XOR U280 ( .A(a[323]), .B(n829), .Z(n831) );
  XOR U281 ( .A(a[326]), .B(n817), .Z(n819) );
  XOR U282 ( .A(a[329]), .B(n804), .Z(n806) );
  XOR U283 ( .A(a[332]), .B(n792), .Z(n794) );
  XOR U284 ( .A(a[335]), .B(n780), .Z(n782) );
  XOR U285 ( .A(a[338]), .B(n768), .Z(n770) );
  XOR U286 ( .A(a[341]), .B(n755), .Z(n757) );
  XOR U287 ( .A(a[344]), .B(n743), .Z(n745) );
  XOR U288 ( .A(a[347]), .B(n731), .Z(n733) );
  XOR U289 ( .A(a[350]), .B(n718), .Z(n720) );
  XOR U290 ( .A(a[353]), .B(n706), .Z(n708) );
  XOR U291 ( .A(a[356]), .B(n694), .Z(n696) );
  XOR U292 ( .A(a[359]), .B(n681), .Z(n683) );
  XOR U293 ( .A(a[362]), .B(n669), .Z(n671) );
  XOR U294 ( .A(a[365]), .B(n657), .Z(n659) );
  XOR U295 ( .A(a[368]), .B(n645), .Z(n647) );
  XOR U296 ( .A(a[371]), .B(n632), .Z(n634) );
  XOR U297 ( .A(a[374]), .B(n620), .Z(n622) );
  XOR U298 ( .A(a[377]), .B(n608), .Z(n610) );
  XOR U299 ( .A(a[380]), .B(n595), .Z(n597) );
  XOR U300 ( .A(a[383]), .B(n583), .Z(n585) );
  XOR U301 ( .A(a[386]), .B(n571), .Z(n573) );
  XOR U302 ( .A(a[389]), .B(n558), .Z(n560) );
  XOR U303 ( .A(a[392]), .B(n546), .Z(n548) );
  XOR U304 ( .A(a[395]), .B(n534), .Z(n536) );
  XOR U305 ( .A(a[398]), .B(n522), .Z(n524) );
  XOR U306 ( .A(a[401]), .B(n508), .Z(n510) );
  XOR U307 ( .A(a[404]), .B(n496), .Z(n498) );
  XOR U308 ( .A(a[407]), .B(n484), .Z(n486) );
  XOR U309 ( .A(a[410]), .B(n471), .Z(n473) );
  XOR U310 ( .A(a[413]), .B(n459), .Z(n461) );
  XOR U311 ( .A(a[416]), .B(n447), .Z(n449) );
  XOR U312 ( .A(a[419]), .B(n434), .Z(n436) );
  XOR U313 ( .A(a[422]), .B(n422), .Z(n424) );
  XOR U314 ( .A(a[425]), .B(n410), .Z(n412) );
  XOR U315 ( .A(a[428]), .B(n398), .Z(n400) );
  XOR U316 ( .A(a[431]), .B(n385), .Z(n387) );
  XOR U317 ( .A(a[434]), .B(n373), .Z(n375) );
  XOR U318 ( .A(a[437]), .B(n361), .Z(n363) );
  XOR U319 ( .A(a[440]), .B(n348), .Z(n350) );
  XOR U320 ( .A(a[443]), .B(n336), .Z(n338) );
  XOR U321 ( .A(a[446]), .B(n324), .Z(n326) );
  XOR U322 ( .A(a[449]), .B(n311), .Z(n313) );
  XOR U323 ( .A(a[452]), .B(n299), .Z(n301) );
  XOR U324 ( .A(a[455]), .B(n287), .Z(n289) );
  XOR U325 ( .A(a[458]), .B(n275), .Z(n277) );
  XOR U326 ( .A(a[461]), .B(n262), .Z(n264) );
  XOR U327 ( .A(a[464]), .B(n250), .Z(n252) );
  XOR U328 ( .A(a[467]), .B(n238), .Z(n240) );
  XOR U329 ( .A(a[470]), .B(n225), .Z(n227) );
  XOR U330 ( .A(a[473]), .B(n213), .Z(n215) );
  XOR U331 ( .A(a[476]), .B(n201), .Z(n203) );
  XOR U332 ( .A(a[479]), .B(n188), .Z(n190) );
  XOR U333 ( .A(a[482]), .B(n176), .Z(n178) );
  XOR U334 ( .A(a[485]), .B(n164), .Z(n166) );
  XOR U335 ( .A(a[488]), .B(n152), .Z(n154) );
  XOR U336 ( .A(a[491]), .B(n139), .Z(n141) );
  XOR U337 ( .A(a[494]), .B(n127), .Z(n129) );
  XOR U338 ( .A(a[497]), .B(n115), .Z(n117) );
  XOR U339 ( .A(a[500]), .B(n101), .Z(n103) );
  XOR U340 ( .A(a[503]), .B(n89), .Z(n91) );
  XOR U341 ( .A(a[506]), .B(n77), .Z(n79) );
  XOR U342 ( .A(a[509]), .B(n64), .Z(n66) );
  XOR U343 ( .A(a[3]), .B(n2037), .Z(n519) );
  XOR U344 ( .A(a[6]), .B(n2028), .Z(n38) );
  XOR U345 ( .A(a[9]), .B(n2019), .Z(n5) );
  XOR U346 ( .A(a[12]), .B(n2010), .Z(n1629) );
  XOR U347 ( .A(a[15]), .B(n2001), .Z(n1506) );
  XOR U348 ( .A(a[18]), .B(n1992), .Z(n1383) );
  XOR U349 ( .A(a[21]), .B(n1983), .Z(n1259) );
  XOR U350 ( .A(a[24]), .B(n1974), .Z(n1136) );
  XOR U351 ( .A(a[27]), .B(n1965), .Z(n1013) );
  XOR U352 ( .A(a[30]), .B(n1956), .Z(n889) );
  XOR U353 ( .A(a[33]), .B(n1947), .Z(n766) );
  XOR U354 ( .A(a[36]), .B(n1938), .Z(n643) );
  XOR U355 ( .A(a[39]), .B(n1929), .Z(n520) );
  XOR U356 ( .A(a[42]), .B(n1920), .Z(n396) );
  XOR U357 ( .A(a[45]), .B(n1911), .Z(n273) );
  XOR U358 ( .A(a[48]), .B(n1902), .Z(n150) );
  XOR U359 ( .A(a[51]), .B(n1893), .Z(n58) );
  XOR U360 ( .A(a[54]), .B(n1884), .Z(n55) );
  XOR U361 ( .A(a[57]), .B(n1875), .Z(n52) );
  XOR U362 ( .A(a[60]), .B(n1866), .Z(n48) );
  XOR U363 ( .A(a[63]), .B(n1857), .Z(n45) );
  XOR U364 ( .A(a[66]), .B(n1848), .Z(n42) );
  XOR U365 ( .A(a[69]), .B(n1839), .Z(n39) );
  XOR U366 ( .A(a[72]), .B(n1830), .Z(n35) );
  XOR U367 ( .A(a[75]), .B(n1821), .Z(n32) );
  XOR U368 ( .A(a[78]), .B(n1812), .Z(n29) );
  XOR U369 ( .A(a[81]), .B(n1803), .Z(n25) );
  XOR U370 ( .A(a[84]), .B(n1794), .Z(n22) );
  XOR U371 ( .A(a[87]), .B(n1785), .Z(n19) );
  XOR U372 ( .A(a[90]), .B(n1776), .Z(n15) );
  XOR U373 ( .A(a[93]), .B(n1767), .Z(n12) );
  XOR U374 ( .A(a[96]), .B(n1758), .Z(n9) );
  XOR U375 ( .A(a[99]), .B(n1749), .Z(n6) );
  XOR U376 ( .A(a[102]), .B(n1737), .Z(n1739) );
  XOR U377 ( .A(a[105]), .B(n1725), .Z(n1727) );
  XOR U378 ( .A(a[108]), .B(n1713), .Z(n1715) );
  XOR U379 ( .A(a[111]), .B(n1700), .Z(n1702) );
  XOR U380 ( .A(a[114]), .B(n1688), .Z(n1690) );
  XOR U381 ( .A(a[117]), .B(n1676), .Z(n1678) );
  XOR U382 ( .A(a[120]), .B(n1663), .Z(n1665) );
  XOR U383 ( .A(a[123]), .B(n1651), .Z(n1653) );
  XOR U384 ( .A(a[126]), .B(n1639), .Z(n1641) );
  XOR U385 ( .A(a[129]), .B(n1626), .Z(n1628) );
  XOR U386 ( .A(a[132]), .B(n1614), .Z(n1616) );
  XOR U387 ( .A(a[135]), .B(n1602), .Z(n1604) );
  XOR U388 ( .A(a[138]), .B(n1590), .Z(n1592) );
  XOR U389 ( .A(a[141]), .B(n1577), .Z(n1579) );
  XOR U390 ( .A(a[144]), .B(n1565), .Z(n1567) );
  XOR U391 ( .A(a[147]), .B(n1553), .Z(n1555) );
  XOR U392 ( .A(a[150]), .B(n1540), .Z(n1542) );
  XOR U393 ( .A(a[153]), .B(n1528), .Z(n1530) );
  XOR U394 ( .A(a[156]), .B(n1516), .Z(n1518) );
  XOR U395 ( .A(a[159]), .B(n1503), .Z(n1505) );
  XOR U396 ( .A(a[162]), .B(n1491), .Z(n1493) );
  XOR U397 ( .A(a[165]), .B(n1479), .Z(n1481) );
  XOR U398 ( .A(a[168]), .B(n1467), .Z(n1469) );
  XOR U399 ( .A(a[171]), .B(n1454), .Z(n1456) );
  XOR U400 ( .A(a[174]), .B(n1442), .Z(n1444) );
  XOR U401 ( .A(a[177]), .B(n1430), .Z(n1432) );
  XOR U402 ( .A(a[180]), .B(n1417), .Z(n1419) );
  XOR U403 ( .A(a[183]), .B(n1405), .Z(n1407) );
  XOR U404 ( .A(a[186]), .B(n1393), .Z(n1395) );
  XOR U405 ( .A(a[189]), .B(n1380), .Z(n1382) );
  XOR U406 ( .A(a[192]), .B(n1368), .Z(n1370) );
  XOR U407 ( .A(a[195]), .B(n1356), .Z(n1358) );
  XOR U408 ( .A(a[198]), .B(n1344), .Z(n1346) );
  XOR U409 ( .A(a[201]), .B(n1330), .Z(n1332) );
  XOR U410 ( .A(a[204]), .B(n1318), .Z(n1320) );
  XOR U411 ( .A(a[207]), .B(n1306), .Z(n1308) );
  XOR U412 ( .A(a[210]), .B(n1293), .Z(n1295) );
  XOR U413 ( .A(a[213]), .B(n1281), .Z(n1283) );
  XOR U414 ( .A(a[216]), .B(n1269), .Z(n1271) );
  XOR U415 ( .A(a[219]), .B(n1256), .Z(n1258) );
  XOR U416 ( .A(a[222]), .B(n1244), .Z(n1246) );
  XOR U417 ( .A(a[225]), .B(n1232), .Z(n1234) );
  XOR U418 ( .A(a[228]), .B(n1220), .Z(n1222) );
  XOR U419 ( .A(a[231]), .B(n1207), .Z(n1209) );
  XOR U420 ( .A(a[234]), .B(n1195), .Z(n1197) );
  XOR U421 ( .A(a[237]), .B(n1183), .Z(n1185) );
  XOR U422 ( .A(a[240]), .B(n1170), .Z(n1172) );
  XOR U423 ( .A(a[243]), .B(n1158), .Z(n1160) );
  XOR U424 ( .A(a[246]), .B(n1146), .Z(n1148) );
  XOR U425 ( .A(a[249]), .B(n1133), .Z(n1135) );
  XOR U426 ( .A(a[252]), .B(n1121), .Z(n1123) );
  XOR U427 ( .A(a[255]), .B(n1109), .Z(n1111) );
  XOR U428 ( .A(a[258]), .B(n1097), .Z(n1099) );
  XOR U429 ( .A(a[261]), .B(n1084), .Z(n1086) );
  XOR U430 ( .A(a[264]), .B(n1072), .Z(n1074) );
  XOR U431 ( .A(a[267]), .B(n1060), .Z(n1062) );
  XOR U432 ( .A(a[270]), .B(n1047), .Z(n1049) );
  XOR U433 ( .A(a[273]), .B(n1035), .Z(n1037) );
  XOR U434 ( .A(a[276]), .B(n1023), .Z(n1025) );
  XOR U435 ( .A(a[279]), .B(n1010), .Z(n1012) );
  XOR U436 ( .A(a[282]), .B(n998), .Z(n1000) );
  XOR U437 ( .A(a[285]), .B(n986), .Z(n988) );
  XOR U438 ( .A(a[288]), .B(n974), .Z(n976) );
  XOR U439 ( .A(a[291]), .B(n961), .Z(n963) );
  XOR U440 ( .A(a[294]), .B(n949), .Z(n951) );
  XOR U441 ( .A(a[297]), .B(n937), .Z(n939) );
  XOR U442 ( .A(a[300]), .B(n923), .Z(n925) );
  XOR U443 ( .A(a[303]), .B(n911), .Z(n913) );
  XOR U444 ( .A(a[306]), .B(n899), .Z(n901) );
  XOR U445 ( .A(a[309]), .B(n886), .Z(n888) );
  XOR U446 ( .A(a[312]), .B(n874), .Z(n876) );
  XOR U447 ( .A(a[315]), .B(n862), .Z(n864) );
  XOR U448 ( .A(a[318]), .B(n850), .Z(n852) );
  XOR U449 ( .A(a[321]), .B(n837), .Z(n839) );
  XOR U450 ( .A(a[324]), .B(n825), .Z(n827) );
  XOR U451 ( .A(a[327]), .B(n813), .Z(n815) );
  XOR U452 ( .A(a[330]), .B(n800), .Z(n802) );
  XOR U453 ( .A(a[333]), .B(n788), .Z(n790) );
  XOR U454 ( .A(a[336]), .B(n776), .Z(n778) );
  XOR U455 ( .A(a[339]), .B(n763), .Z(n765) );
  XOR U456 ( .A(a[342]), .B(n751), .Z(n753) );
  XOR U457 ( .A(a[345]), .B(n739), .Z(n741) );
  XOR U458 ( .A(a[348]), .B(n727), .Z(n729) );
  XOR U459 ( .A(a[351]), .B(n714), .Z(n716) );
  XOR U460 ( .A(a[354]), .B(n702), .Z(n704) );
  XOR U461 ( .A(a[357]), .B(n690), .Z(n692) );
  XOR U462 ( .A(a[360]), .B(n677), .Z(n679) );
  XOR U463 ( .A(a[363]), .B(n665), .Z(n667) );
  XOR U464 ( .A(a[366]), .B(n653), .Z(n655) );
  XOR U465 ( .A(a[369]), .B(n640), .Z(n642) );
  XOR U466 ( .A(a[372]), .B(n628), .Z(n630) );
  XOR U467 ( .A(a[375]), .B(n616), .Z(n618) );
  XOR U468 ( .A(a[378]), .B(n604), .Z(n606) );
  XOR U469 ( .A(a[381]), .B(n591), .Z(n593) );
  XOR U470 ( .A(a[384]), .B(n579), .Z(n581) );
  XOR U471 ( .A(a[387]), .B(n567), .Z(n569) );
  XOR U472 ( .A(a[390]), .B(n554), .Z(n556) );
  XOR U473 ( .A(a[393]), .B(n542), .Z(n544) );
  XOR U474 ( .A(a[396]), .B(n530), .Z(n532) );
  XOR U475 ( .A(a[399]), .B(n516), .Z(n518) );
  XOR U476 ( .A(a[402]), .B(n504), .Z(n506) );
  XOR U477 ( .A(a[405]), .B(n492), .Z(n494) );
  XOR U478 ( .A(a[408]), .B(n480), .Z(n482) );
  XOR U479 ( .A(a[411]), .B(n467), .Z(n469) );
  XOR U480 ( .A(a[414]), .B(n455), .Z(n457) );
  XOR U481 ( .A(a[417]), .B(n443), .Z(n445) );
  XOR U482 ( .A(a[420]), .B(n430), .Z(n432) );
  XOR U483 ( .A(a[423]), .B(n418), .Z(n420) );
  XOR U484 ( .A(a[426]), .B(n406), .Z(n408) );
  XOR U485 ( .A(a[429]), .B(n393), .Z(n395) );
  XOR U486 ( .A(a[432]), .B(n381), .Z(n383) );
  XOR U487 ( .A(a[435]), .B(n369), .Z(n371) );
  XOR U488 ( .A(a[438]), .B(n357), .Z(n359) );
  XOR U489 ( .A(a[441]), .B(n344), .Z(n346) );
  XOR U490 ( .A(a[444]), .B(n332), .Z(n334) );
  XOR U491 ( .A(a[447]), .B(n320), .Z(n322) );
  XOR U492 ( .A(a[450]), .B(n307), .Z(n309) );
  XOR U493 ( .A(a[453]), .B(n295), .Z(n297) );
  XOR U494 ( .A(a[456]), .B(n283), .Z(n285) );
  XOR U495 ( .A(a[459]), .B(n270), .Z(n272) );
  XOR U496 ( .A(a[462]), .B(n258), .Z(n260) );
  XOR U497 ( .A(a[465]), .B(n246), .Z(n248) );
  XOR U498 ( .A(a[468]), .B(n234), .Z(n236) );
  XOR U499 ( .A(a[471]), .B(n221), .Z(n223) );
  XOR U500 ( .A(a[474]), .B(n209), .Z(n211) );
  XOR U501 ( .A(a[477]), .B(n197), .Z(n199) );
  XOR U502 ( .A(a[480]), .B(n184), .Z(n186) );
  XOR U503 ( .A(a[483]), .B(n172), .Z(n174) );
  XOR U504 ( .A(a[486]), .B(n160), .Z(n162) );
  XOR U505 ( .A(a[489]), .B(n147), .Z(n149) );
  XOR U506 ( .A(a[492]), .B(n135), .Z(n137) );
  XOR U507 ( .A(a[495]), .B(n123), .Z(n125) );
  XOR U508 ( .A(a[498]), .B(n111), .Z(n113) );
  XOR U509 ( .A(a[501]), .B(n97), .Z(n99) );
  XOR U510 ( .A(a[504]), .B(n85), .Z(n87) );
  XOR U511 ( .A(a[507]), .B(n73), .Z(n75) );
  XOR U512 ( .A(a[510]), .B(n60), .Z(n62) );
  XOR U513 ( .A(n1), .B(n2), .Z(carry_on_d) );
  ANDN U514 ( .B(n3), .A(n4), .Z(n1) );
  XOR U515 ( .A(b[511]), .B(n2), .Z(n3) );
  XNOR U516 ( .A(b[9]), .B(n5), .Z(c[9]) );
  XNOR U517 ( .A(b[99]), .B(n6), .Z(c[99]) );
  XNOR U518 ( .A(b[98]), .B(n7), .Z(c[98]) );
  XNOR U519 ( .A(b[97]), .B(n8), .Z(c[97]) );
  XNOR U520 ( .A(b[96]), .B(n9), .Z(c[96]) );
  XNOR U521 ( .A(b[95]), .B(n10), .Z(c[95]) );
  XNOR U522 ( .A(b[94]), .B(n11), .Z(c[94]) );
  XNOR U523 ( .A(b[93]), .B(n12), .Z(c[93]) );
  XNOR U524 ( .A(b[92]), .B(n13), .Z(c[92]) );
  XNOR U525 ( .A(b[91]), .B(n14), .Z(c[91]) );
  XNOR U526 ( .A(b[90]), .B(n15), .Z(c[90]) );
  XNOR U527 ( .A(b[8]), .B(n16), .Z(c[8]) );
  XNOR U528 ( .A(b[89]), .B(n17), .Z(c[89]) );
  XNOR U529 ( .A(b[88]), .B(n18), .Z(c[88]) );
  XNOR U530 ( .A(b[87]), .B(n19), .Z(c[87]) );
  XNOR U531 ( .A(b[86]), .B(n20), .Z(c[86]) );
  XNOR U532 ( .A(b[85]), .B(n21), .Z(c[85]) );
  XNOR U533 ( .A(b[84]), .B(n22), .Z(c[84]) );
  XNOR U534 ( .A(b[83]), .B(n23), .Z(c[83]) );
  XNOR U535 ( .A(b[82]), .B(n24), .Z(c[82]) );
  XNOR U536 ( .A(b[81]), .B(n25), .Z(c[81]) );
  XNOR U537 ( .A(b[80]), .B(n26), .Z(c[80]) );
  XNOR U538 ( .A(b[7]), .B(n27), .Z(c[7]) );
  XNOR U539 ( .A(b[79]), .B(n28), .Z(c[79]) );
  XNOR U540 ( .A(b[78]), .B(n29), .Z(c[78]) );
  XNOR U541 ( .A(b[77]), .B(n30), .Z(c[77]) );
  XNOR U542 ( .A(b[76]), .B(n31), .Z(c[76]) );
  XNOR U543 ( .A(b[75]), .B(n32), .Z(c[75]) );
  XNOR U544 ( .A(b[74]), .B(n33), .Z(c[74]) );
  XNOR U545 ( .A(b[73]), .B(n34), .Z(c[73]) );
  XNOR U546 ( .A(b[72]), .B(n35), .Z(c[72]) );
  XNOR U547 ( .A(b[71]), .B(n36), .Z(c[71]) );
  XNOR U548 ( .A(b[70]), .B(n37), .Z(c[70]) );
  XNOR U549 ( .A(b[6]), .B(n38), .Z(c[6]) );
  XNOR U550 ( .A(b[69]), .B(n39), .Z(c[69]) );
  XNOR U551 ( .A(b[68]), .B(n40), .Z(c[68]) );
  XNOR U552 ( .A(b[67]), .B(n41), .Z(c[67]) );
  XNOR U553 ( .A(b[66]), .B(n42), .Z(c[66]) );
  XNOR U554 ( .A(b[65]), .B(n43), .Z(c[65]) );
  XNOR U555 ( .A(b[64]), .B(n44), .Z(c[64]) );
  XNOR U556 ( .A(b[63]), .B(n45), .Z(c[63]) );
  XNOR U557 ( .A(b[62]), .B(n46), .Z(c[62]) );
  XNOR U558 ( .A(b[61]), .B(n47), .Z(c[61]) );
  XNOR U559 ( .A(b[60]), .B(n48), .Z(c[60]) );
  XNOR U560 ( .A(b[5]), .B(n49), .Z(c[5]) );
  XNOR U561 ( .A(b[59]), .B(n50), .Z(c[59]) );
  XNOR U562 ( .A(b[58]), .B(n51), .Z(c[58]) );
  XNOR U563 ( .A(b[57]), .B(n52), .Z(c[57]) );
  XNOR U564 ( .A(b[56]), .B(n53), .Z(c[56]) );
  XNOR U565 ( .A(b[55]), .B(n54), .Z(c[55]) );
  XNOR U566 ( .A(b[54]), .B(n55), .Z(c[54]) );
  XNOR U567 ( .A(b[53]), .B(n56), .Z(c[53]) );
  XNOR U568 ( .A(b[52]), .B(n57), .Z(c[52]) );
  XNOR U569 ( .A(b[51]), .B(n58), .Z(c[51]) );
  XNOR U570 ( .A(b[511]), .B(n4), .Z(c[511]) );
  XNOR U571 ( .A(a[511]), .B(n2), .Z(n4) );
  XNOR U572 ( .A(n59), .B(n60), .Z(n2) );
  ANDN U573 ( .B(n61), .A(n62), .Z(n59) );
  XNOR U574 ( .A(b[510]), .B(n60), .Z(n61) );
  XNOR U575 ( .A(b[510]), .B(n62), .Z(c[510]) );
  XOR U576 ( .A(n63), .B(n64), .Z(n60) );
  ANDN U577 ( .B(n65), .A(n66), .Z(n63) );
  XNOR U578 ( .A(b[509]), .B(n64), .Z(n65) );
  XNOR U579 ( .A(b[50]), .B(n67), .Z(c[50]) );
  XNOR U580 ( .A(b[509]), .B(n66), .Z(c[509]) );
  XOR U581 ( .A(n68), .B(n69), .Z(n64) );
  ANDN U582 ( .B(n70), .A(n71), .Z(n68) );
  XNOR U583 ( .A(b[508]), .B(n69), .Z(n70) );
  XNOR U584 ( .A(b[508]), .B(n71), .Z(c[508]) );
  XOR U585 ( .A(n72), .B(n73), .Z(n69) );
  ANDN U586 ( .B(n74), .A(n75), .Z(n72) );
  XNOR U587 ( .A(b[507]), .B(n73), .Z(n74) );
  XNOR U588 ( .A(b[507]), .B(n75), .Z(c[507]) );
  XOR U589 ( .A(n76), .B(n77), .Z(n73) );
  ANDN U590 ( .B(n78), .A(n79), .Z(n76) );
  XNOR U591 ( .A(b[506]), .B(n77), .Z(n78) );
  XNOR U592 ( .A(b[506]), .B(n79), .Z(c[506]) );
  XOR U593 ( .A(n80), .B(n81), .Z(n77) );
  ANDN U594 ( .B(n82), .A(n83), .Z(n80) );
  XNOR U595 ( .A(b[505]), .B(n81), .Z(n82) );
  XNOR U596 ( .A(b[505]), .B(n83), .Z(c[505]) );
  XOR U597 ( .A(n84), .B(n85), .Z(n81) );
  ANDN U598 ( .B(n86), .A(n87), .Z(n84) );
  XNOR U599 ( .A(b[504]), .B(n85), .Z(n86) );
  XNOR U600 ( .A(b[504]), .B(n87), .Z(c[504]) );
  XOR U601 ( .A(n88), .B(n89), .Z(n85) );
  ANDN U602 ( .B(n90), .A(n91), .Z(n88) );
  XNOR U603 ( .A(b[503]), .B(n89), .Z(n90) );
  XNOR U604 ( .A(b[503]), .B(n91), .Z(c[503]) );
  XOR U605 ( .A(n92), .B(n93), .Z(n89) );
  ANDN U606 ( .B(n94), .A(n95), .Z(n92) );
  XNOR U607 ( .A(b[502]), .B(n93), .Z(n94) );
  XNOR U608 ( .A(b[502]), .B(n95), .Z(c[502]) );
  XOR U609 ( .A(n96), .B(n97), .Z(n93) );
  ANDN U610 ( .B(n98), .A(n99), .Z(n96) );
  XNOR U611 ( .A(b[501]), .B(n97), .Z(n98) );
  XNOR U612 ( .A(b[501]), .B(n99), .Z(c[501]) );
  XOR U613 ( .A(n100), .B(n101), .Z(n97) );
  ANDN U614 ( .B(n102), .A(n103), .Z(n100) );
  XNOR U615 ( .A(b[500]), .B(n101), .Z(n102) );
  XNOR U616 ( .A(b[500]), .B(n103), .Z(c[500]) );
  XOR U617 ( .A(n104), .B(n105), .Z(n101) );
  ANDN U618 ( .B(n106), .A(n107), .Z(n104) );
  XNOR U619 ( .A(b[499]), .B(n105), .Z(n106) );
  XNOR U620 ( .A(b[4]), .B(n108), .Z(c[4]) );
  XNOR U621 ( .A(b[49]), .B(n109), .Z(c[49]) );
  XNOR U622 ( .A(b[499]), .B(n107), .Z(c[499]) );
  XOR U623 ( .A(n110), .B(n111), .Z(n105) );
  ANDN U624 ( .B(n112), .A(n113), .Z(n110) );
  XNOR U625 ( .A(b[498]), .B(n111), .Z(n112) );
  XNOR U626 ( .A(b[498]), .B(n113), .Z(c[498]) );
  XOR U627 ( .A(n114), .B(n115), .Z(n111) );
  ANDN U628 ( .B(n116), .A(n117), .Z(n114) );
  XNOR U629 ( .A(b[497]), .B(n115), .Z(n116) );
  XNOR U630 ( .A(b[497]), .B(n117), .Z(c[497]) );
  XOR U631 ( .A(n118), .B(n119), .Z(n115) );
  ANDN U632 ( .B(n120), .A(n121), .Z(n118) );
  XNOR U633 ( .A(b[496]), .B(n119), .Z(n120) );
  XNOR U634 ( .A(b[496]), .B(n121), .Z(c[496]) );
  XOR U635 ( .A(n122), .B(n123), .Z(n119) );
  ANDN U636 ( .B(n124), .A(n125), .Z(n122) );
  XNOR U637 ( .A(b[495]), .B(n123), .Z(n124) );
  XNOR U638 ( .A(b[495]), .B(n125), .Z(c[495]) );
  XOR U639 ( .A(n126), .B(n127), .Z(n123) );
  ANDN U640 ( .B(n128), .A(n129), .Z(n126) );
  XNOR U641 ( .A(b[494]), .B(n127), .Z(n128) );
  XNOR U642 ( .A(b[494]), .B(n129), .Z(c[494]) );
  XOR U643 ( .A(n130), .B(n131), .Z(n127) );
  ANDN U644 ( .B(n132), .A(n133), .Z(n130) );
  XNOR U645 ( .A(b[493]), .B(n131), .Z(n132) );
  XNOR U646 ( .A(b[493]), .B(n133), .Z(c[493]) );
  XOR U647 ( .A(n134), .B(n135), .Z(n131) );
  ANDN U648 ( .B(n136), .A(n137), .Z(n134) );
  XNOR U649 ( .A(b[492]), .B(n135), .Z(n136) );
  XNOR U650 ( .A(b[492]), .B(n137), .Z(c[492]) );
  XOR U651 ( .A(n138), .B(n139), .Z(n135) );
  ANDN U652 ( .B(n140), .A(n141), .Z(n138) );
  XNOR U653 ( .A(b[491]), .B(n139), .Z(n140) );
  XNOR U654 ( .A(b[491]), .B(n141), .Z(c[491]) );
  XOR U655 ( .A(n142), .B(n143), .Z(n139) );
  ANDN U656 ( .B(n144), .A(n145), .Z(n142) );
  XNOR U657 ( .A(b[490]), .B(n143), .Z(n144) );
  XNOR U658 ( .A(b[490]), .B(n145), .Z(c[490]) );
  XOR U659 ( .A(n146), .B(n147), .Z(n143) );
  ANDN U660 ( .B(n148), .A(n149), .Z(n146) );
  XNOR U661 ( .A(b[489]), .B(n147), .Z(n148) );
  XNOR U662 ( .A(b[48]), .B(n150), .Z(c[48]) );
  XNOR U663 ( .A(b[489]), .B(n149), .Z(c[489]) );
  XOR U664 ( .A(n151), .B(n152), .Z(n147) );
  ANDN U665 ( .B(n153), .A(n154), .Z(n151) );
  XNOR U666 ( .A(b[488]), .B(n152), .Z(n153) );
  XNOR U667 ( .A(b[488]), .B(n154), .Z(c[488]) );
  XOR U668 ( .A(n155), .B(n156), .Z(n152) );
  ANDN U669 ( .B(n157), .A(n158), .Z(n155) );
  XNOR U670 ( .A(b[487]), .B(n156), .Z(n157) );
  XNOR U671 ( .A(b[487]), .B(n158), .Z(c[487]) );
  XOR U672 ( .A(n159), .B(n160), .Z(n156) );
  ANDN U673 ( .B(n161), .A(n162), .Z(n159) );
  XNOR U674 ( .A(b[486]), .B(n160), .Z(n161) );
  XNOR U675 ( .A(b[486]), .B(n162), .Z(c[486]) );
  XOR U676 ( .A(n163), .B(n164), .Z(n160) );
  ANDN U677 ( .B(n165), .A(n166), .Z(n163) );
  XNOR U678 ( .A(b[485]), .B(n164), .Z(n165) );
  XNOR U679 ( .A(b[485]), .B(n166), .Z(c[485]) );
  XOR U680 ( .A(n167), .B(n168), .Z(n164) );
  ANDN U681 ( .B(n169), .A(n170), .Z(n167) );
  XNOR U682 ( .A(b[484]), .B(n168), .Z(n169) );
  XNOR U683 ( .A(b[484]), .B(n170), .Z(c[484]) );
  XOR U684 ( .A(n171), .B(n172), .Z(n168) );
  ANDN U685 ( .B(n173), .A(n174), .Z(n171) );
  XNOR U686 ( .A(b[483]), .B(n172), .Z(n173) );
  XNOR U687 ( .A(b[483]), .B(n174), .Z(c[483]) );
  XOR U688 ( .A(n175), .B(n176), .Z(n172) );
  ANDN U689 ( .B(n177), .A(n178), .Z(n175) );
  XNOR U690 ( .A(b[482]), .B(n176), .Z(n177) );
  XNOR U691 ( .A(b[482]), .B(n178), .Z(c[482]) );
  XOR U692 ( .A(n179), .B(n180), .Z(n176) );
  ANDN U693 ( .B(n181), .A(n182), .Z(n179) );
  XNOR U694 ( .A(b[481]), .B(n180), .Z(n181) );
  XNOR U695 ( .A(b[481]), .B(n182), .Z(c[481]) );
  XOR U696 ( .A(n183), .B(n184), .Z(n180) );
  ANDN U697 ( .B(n185), .A(n186), .Z(n183) );
  XNOR U698 ( .A(b[480]), .B(n184), .Z(n185) );
  XNOR U699 ( .A(b[480]), .B(n186), .Z(c[480]) );
  XOR U700 ( .A(n187), .B(n188), .Z(n184) );
  ANDN U701 ( .B(n189), .A(n190), .Z(n187) );
  XNOR U702 ( .A(b[479]), .B(n188), .Z(n189) );
  XNOR U703 ( .A(b[47]), .B(n191), .Z(c[47]) );
  XNOR U704 ( .A(b[479]), .B(n190), .Z(c[479]) );
  XOR U705 ( .A(n192), .B(n193), .Z(n188) );
  ANDN U706 ( .B(n194), .A(n195), .Z(n192) );
  XNOR U707 ( .A(b[478]), .B(n193), .Z(n194) );
  XNOR U708 ( .A(b[478]), .B(n195), .Z(c[478]) );
  XOR U709 ( .A(n196), .B(n197), .Z(n193) );
  ANDN U710 ( .B(n198), .A(n199), .Z(n196) );
  XNOR U711 ( .A(b[477]), .B(n197), .Z(n198) );
  XNOR U712 ( .A(b[477]), .B(n199), .Z(c[477]) );
  XOR U713 ( .A(n200), .B(n201), .Z(n197) );
  ANDN U714 ( .B(n202), .A(n203), .Z(n200) );
  XNOR U715 ( .A(b[476]), .B(n201), .Z(n202) );
  XNOR U716 ( .A(b[476]), .B(n203), .Z(c[476]) );
  XOR U717 ( .A(n204), .B(n205), .Z(n201) );
  ANDN U718 ( .B(n206), .A(n207), .Z(n204) );
  XNOR U719 ( .A(b[475]), .B(n205), .Z(n206) );
  XNOR U720 ( .A(b[475]), .B(n207), .Z(c[475]) );
  XOR U721 ( .A(n208), .B(n209), .Z(n205) );
  ANDN U722 ( .B(n210), .A(n211), .Z(n208) );
  XNOR U723 ( .A(b[474]), .B(n209), .Z(n210) );
  XNOR U724 ( .A(b[474]), .B(n211), .Z(c[474]) );
  XOR U725 ( .A(n212), .B(n213), .Z(n209) );
  ANDN U726 ( .B(n214), .A(n215), .Z(n212) );
  XNOR U727 ( .A(b[473]), .B(n213), .Z(n214) );
  XNOR U728 ( .A(b[473]), .B(n215), .Z(c[473]) );
  XOR U729 ( .A(n216), .B(n217), .Z(n213) );
  ANDN U730 ( .B(n218), .A(n219), .Z(n216) );
  XNOR U731 ( .A(b[472]), .B(n217), .Z(n218) );
  XNOR U732 ( .A(b[472]), .B(n219), .Z(c[472]) );
  XOR U733 ( .A(n220), .B(n221), .Z(n217) );
  ANDN U734 ( .B(n222), .A(n223), .Z(n220) );
  XNOR U735 ( .A(b[471]), .B(n221), .Z(n222) );
  XNOR U736 ( .A(b[471]), .B(n223), .Z(c[471]) );
  XOR U737 ( .A(n224), .B(n225), .Z(n221) );
  ANDN U738 ( .B(n226), .A(n227), .Z(n224) );
  XNOR U739 ( .A(b[470]), .B(n225), .Z(n226) );
  XNOR U740 ( .A(b[470]), .B(n227), .Z(c[470]) );
  XOR U741 ( .A(n228), .B(n229), .Z(n225) );
  ANDN U742 ( .B(n230), .A(n231), .Z(n228) );
  XNOR U743 ( .A(b[469]), .B(n229), .Z(n230) );
  XNOR U744 ( .A(b[46]), .B(n232), .Z(c[46]) );
  XNOR U745 ( .A(b[469]), .B(n231), .Z(c[469]) );
  XOR U746 ( .A(n233), .B(n234), .Z(n229) );
  ANDN U747 ( .B(n235), .A(n236), .Z(n233) );
  XNOR U748 ( .A(b[468]), .B(n234), .Z(n235) );
  XNOR U749 ( .A(b[468]), .B(n236), .Z(c[468]) );
  XOR U750 ( .A(n237), .B(n238), .Z(n234) );
  ANDN U751 ( .B(n239), .A(n240), .Z(n237) );
  XNOR U752 ( .A(b[467]), .B(n238), .Z(n239) );
  XNOR U753 ( .A(b[467]), .B(n240), .Z(c[467]) );
  XOR U754 ( .A(n241), .B(n242), .Z(n238) );
  ANDN U755 ( .B(n243), .A(n244), .Z(n241) );
  XNOR U756 ( .A(b[466]), .B(n242), .Z(n243) );
  XNOR U757 ( .A(b[466]), .B(n244), .Z(c[466]) );
  XOR U758 ( .A(n245), .B(n246), .Z(n242) );
  ANDN U759 ( .B(n247), .A(n248), .Z(n245) );
  XNOR U760 ( .A(b[465]), .B(n246), .Z(n247) );
  XNOR U761 ( .A(b[465]), .B(n248), .Z(c[465]) );
  XOR U762 ( .A(n249), .B(n250), .Z(n246) );
  ANDN U763 ( .B(n251), .A(n252), .Z(n249) );
  XNOR U764 ( .A(b[464]), .B(n250), .Z(n251) );
  XNOR U765 ( .A(b[464]), .B(n252), .Z(c[464]) );
  XOR U766 ( .A(n253), .B(n254), .Z(n250) );
  ANDN U767 ( .B(n255), .A(n256), .Z(n253) );
  XNOR U768 ( .A(b[463]), .B(n254), .Z(n255) );
  XNOR U769 ( .A(b[463]), .B(n256), .Z(c[463]) );
  XOR U770 ( .A(n257), .B(n258), .Z(n254) );
  ANDN U771 ( .B(n259), .A(n260), .Z(n257) );
  XNOR U772 ( .A(b[462]), .B(n258), .Z(n259) );
  XNOR U773 ( .A(b[462]), .B(n260), .Z(c[462]) );
  XOR U774 ( .A(n261), .B(n262), .Z(n258) );
  ANDN U775 ( .B(n263), .A(n264), .Z(n261) );
  XNOR U776 ( .A(b[461]), .B(n262), .Z(n263) );
  XNOR U777 ( .A(b[461]), .B(n264), .Z(c[461]) );
  XOR U778 ( .A(n265), .B(n266), .Z(n262) );
  ANDN U779 ( .B(n267), .A(n268), .Z(n265) );
  XNOR U780 ( .A(b[460]), .B(n266), .Z(n267) );
  XNOR U781 ( .A(b[460]), .B(n268), .Z(c[460]) );
  XOR U782 ( .A(n269), .B(n270), .Z(n266) );
  ANDN U783 ( .B(n271), .A(n272), .Z(n269) );
  XNOR U784 ( .A(b[459]), .B(n270), .Z(n271) );
  XNOR U785 ( .A(b[45]), .B(n273), .Z(c[45]) );
  XNOR U786 ( .A(b[459]), .B(n272), .Z(c[459]) );
  XOR U787 ( .A(n274), .B(n275), .Z(n270) );
  ANDN U788 ( .B(n276), .A(n277), .Z(n274) );
  XNOR U789 ( .A(b[458]), .B(n275), .Z(n276) );
  XNOR U790 ( .A(b[458]), .B(n277), .Z(c[458]) );
  XOR U791 ( .A(n278), .B(n279), .Z(n275) );
  ANDN U792 ( .B(n280), .A(n281), .Z(n278) );
  XNOR U793 ( .A(b[457]), .B(n279), .Z(n280) );
  XNOR U794 ( .A(b[457]), .B(n281), .Z(c[457]) );
  XOR U795 ( .A(n282), .B(n283), .Z(n279) );
  ANDN U796 ( .B(n284), .A(n285), .Z(n282) );
  XNOR U797 ( .A(b[456]), .B(n283), .Z(n284) );
  XNOR U798 ( .A(b[456]), .B(n285), .Z(c[456]) );
  XOR U799 ( .A(n286), .B(n287), .Z(n283) );
  ANDN U800 ( .B(n288), .A(n289), .Z(n286) );
  XNOR U801 ( .A(b[455]), .B(n287), .Z(n288) );
  XNOR U802 ( .A(b[455]), .B(n289), .Z(c[455]) );
  XOR U803 ( .A(n290), .B(n291), .Z(n287) );
  ANDN U804 ( .B(n292), .A(n293), .Z(n290) );
  XNOR U805 ( .A(b[454]), .B(n291), .Z(n292) );
  XNOR U806 ( .A(b[454]), .B(n293), .Z(c[454]) );
  XOR U807 ( .A(n294), .B(n295), .Z(n291) );
  ANDN U808 ( .B(n296), .A(n297), .Z(n294) );
  XNOR U809 ( .A(b[453]), .B(n295), .Z(n296) );
  XNOR U810 ( .A(b[453]), .B(n297), .Z(c[453]) );
  XOR U811 ( .A(n298), .B(n299), .Z(n295) );
  ANDN U812 ( .B(n300), .A(n301), .Z(n298) );
  XNOR U813 ( .A(b[452]), .B(n299), .Z(n300) );
  XNOR U814 ( .A(b[452]), .B(n301), .Z(c[452]) );
  XOR U815 ( .A(n302), .B(n303), .Z(n299) );
  ANDN U816 ( .B(n304), .A(n305), .Z(n302) );
  XNOR U817 ( .A(b[451]), .B(n303), .Z(n304) );
  XNOR U818 ( .A(b[451]), .B(n305), .Z(c[451]) );
  XOR U819 ( .A(n306), .B(n307), .Z(n303) );
  ANDN U820 ( .B(n308), .A(n309), .Z(n306) );
  XNOR U821 ( .A(b[450]), .B(n307), .Z(n308) );
  XNOR U822 ( .A(b[450]), .B(n309), .Z(c[450]) );
  XOR U823 ( .A(n310), .B(n311), .Z(n307) );
  ANDN U824 ( .B(n312), .A(n313), .Z(n310) );
  XNOR U825 ( .A(b[449]), .B(n311), .Z(n312) );
  XNOR U826 ( .A(b[44]), .B(n314), .Z(c[44]) );
  XNOR U827 ( .A(b[449]), .B(n313), .Z(c[449]) );
  XOR U828 ( .A(n315), .B(n316), .Z(n311) );
  ANDN U829 ( .B(n317), .A(n318), .Z(n315) );
  XNOR U830 ( .A(b[448]), .B(n316), .Z(n317) );
  XNOR U831 ( .A(b[448]), .B(n318), .Z(c[448]) );
  XOR U832 ( .A(n319), .B(n320), .Z(n316) );
  ANDN U833 ( .B(n321), .A(n322), .Z(n319) );
  XNOR U834 ( .A(b[447]), .B(n320), .Z(n321) );
  XNOR U835 ( .A(b[447]), .B(n322), .Z(c[447]) );
  XOR U836 ( .A(n323), .B(n324), .Z(n320) );
  ANDN U837 ( .B(n325), .A(n326), .Z(n323) );
  XNOR U838 ( .A(b[446]), .B(n324), .Z(n325) );
  XNOR U839 ( .A(b[446]), .B(n326), .Z(c[446]) );
  XOR U840 ( .A(n327), .B(n328), .Z(n324) );
  ANDN U841 ( .B(n329), .A(n330), .Z(n327) );
  XNOR U842 ( .A(b[445]), .B(n328), .Z(n329) );
  XNOR U843 ( .A(b[445]), .B(n330), .Z(c[445]) );
  XOR U844 ( .A(n331), .B(n332), .Z(n328) );
  ANDN U845 ( .B(n333), .A(n334), .Z(n331) );
  XNOR U846 ( .A(b[444]), .B(n332), .Z(n333) );
  XNOR U847 ( .A(b[444]), .B(n334), .Z(c[444]) );
  XOR U848 ( .A(n335), .B(n336), .Z(n332) );
  ANDN U849 ( .B(n337), .A(n338), .Z(n335) );
  XNOR U850 ( .A(b[443]), .B(n336), .Z(n337) );
  XNOR U851 ( .A(b[443]), .B(n338), .Z(c[443]) );
  XOR U852 ( .A(n339), .B(n340), .Z(n336) );
  ANDN U853 ( .B(n341), .A(n342), .Z(n339) );
  XNOR U854 ( .A(b[442]), .B(n340), .Z(n341) );
  XNOR U855 ( .A(b[442]), .B(n342), .Z(c[442]) );
  XOR U856 ( .A(n343), .B(n344), .Z(n340) );
  ANDN U857 ( .B(n345), .A(n346), .Z(n343) );
  XNOR U858 ( .A(b[441]), .B(n344), .Z(n345) );
  XNOR U859 ( .A(b[441]), .B(n346), .Z(c[441]) );
  XOR U860 ( .A(n347), .B(n348), .Z(n344) );
  ANDN U861 ( .B(n349), .A(n350), .Z(n347) );
  XNOR U862 ( .A(b[440]), .B(n348), .Z(n349) );
  XNOR U863 ( .A(b[440]), .B(n350), .Z(c[440]) );
  XOR U864 ( .A(n351), .B(n352), .Z(n348) );
  ANDN U865 ( .B(n353), .A(n354), .Z(n351) );
  XNOR U866 ( .A(b[439]), .B(n352), .Z(n353) );
  XNOR U867 ( .A(b[43]), .B(n355), .Z(c[43]) );
  XNOR U868 ( .A(b[439]), .B(n354), .Z(c[439]) );
  XOR U869 ( .A(n356), .B(n357), .Z(n352) );
  ANDN U870 ( .B(n358), .A(n359), .Z(n356) );
  XNOR U871 ( .A(b[438]), .B(n357), .Z(n358) );
  XNOR U872 ( .A(b[438]), .B(n359), .Z(c[438]) );
  XOR U873 ( .A(n360), .B(n361), .Z(n357) );
  ANDN U874 ( .B(n362), .A(n363), .Z(n360) );
  XNOR U875 ( .A(b[437]), .B(n361), .Z(n362) );
  XNOR U876 ( .A(b[437]), .B(n363), .Z(c[437]) );
  XOR U877 ( .A(n364), .B(n365), .Z(n361) );
  ANDN U878 ( .B(n366), .A(n367), .Z(n364) );
  XNOR U879 ( .A(b[436]), .B(n365), .Z(n366) );
  XNOR U880 ( .A(b[436]), .B(n367), .Z(c[436]) );
  XOR U881 ( .A(n368), .B(n369), .Z(n365) );
  ANDN U882 ( .B(n370), .A(n371), .Z(n368) );
  XNOR U883 ( .A(b[435]), .B(n369), .Z(n370) );
  XNOR U884 ( .A(b[435]), .B(n371), .Z(c[435]) );
  XOR U885 ( .A(n372), .B(n373), .Z(n369) );
  ANDN U886 ( .B(n374), .A(n375), .Z(n372) );
  XNOR U887 ( .A(b[434]), .B(n373), .Z(n374) );
  XNOR U888 ( .A(b[434]), .B(n375), .Z(c[434]) );
  XOR U889 ( .A(n376), .B(n377), .Z(n373) );
  ANDN U890 ( .B(n378), .A(n379), .Z(n376) );
  XNOR U891 ( .A(b[433]), .B(n377), .Z(n378) );
  XNOR U892 ( .A(b[433]), .B(n379), .Z(c[433]) );
  XOR U893 ( .A(n380), .B(n381), .Z(n377) );
  ANDN U894 ( .B(n382), .A(n383), .Z(n380) );
  XNOR U895 ( .A(b[432]), .B(n381), .Z(n382) );
  XNOR U896 ( .A(b[432]), .B(n383), .Z(c[432]) );
  XOR U897 ( .A(n384), .B(n385), .Z(n381) );
  ANDN U898 ( .B(n386), .A(n387), .Z(n384) );
  XNOR U899 ( .A(b[431]), .B(n385), .Z(n386) );
  XNOR U900 ( .A(b[431]), .B(n387), .Z(c[431]) );
  XOR U901 ( .A(n388), .B(n389), .Z(n385) );
  ANDN U902 ( .B(n390), .A(n391), .Z(n388) );
  XNOR U903 ( .A(b[430]), .B(n389), .Z(n390) );
  XNOR U904 ( .A(b[430]), .B(n391), .Z(c[430]) );
  XOR U905 ( .A(n392), .B(n393), .Z(n389) );
  ANDN U906 ( .B(n394), .A(n395), .Z(n392) );
  XNOR U907 ( .A(b[429]), .B(n393), .Z(n394) );
  XNOR U908 ( .A(b[42]), .B(n396), .Z(c[42]) );
  XNOR U909 ( .A(b[429]), .B(n395), .Z(c[429]) );
  XOR U910 ( .A(n397), .B(n398), .Z(n393) );
  ANDN U911 ( .B(n399), .A(n400), .Z(n397) );
  XNOR U912 ( .A(b[428]), .B(n398), .Z(n399) );
  XNOR U913 ( .A(b[428]), .B(n400), .Z(c[428]) );
  XOR U914 ( .A(n401), .B(n402), .Z(n398) );
  ANDN U915 ( .B(n403), .A(n404), .Z(n401) );
  XNOR U916 ( .A(b[427]), .B(n402), .Z(n403) );
  XNOR U917 ( .A(b[427]), .B(n404), .Z(c[427]) );
  XOR U918 ( .A(n405), .B(n406), .Z(n402) );
  ANDN U919 ( .B(n407), .A(n408), .Z(n405) );
  XNOR U920 ( .A(b[426]), .B(n406), .Z(n407) );
  XNOR U921 ( .A(b[426]), .B(n408), .Z(c[426]) );
  XOR U922 ( .A(n409), .B(n410), .Z(n406) );
  ANDN U923 ( .B(n411), .A(n412), .Z(n409) );
  XNOR U924 ( .A(b[425]), .B(n410), .Z(n411) );
  XNOR U925 ( .A(b[425]), .B(n412), .Z(c[425]) );
  XOR U926 ( .A(n413), .B(n414), .Z(n410) );
  ANDN U927 ( .B(n415), .A(n416), .Z(n413) );
  XNOR U928 ( .A(b[424]), .B(n414), .Z(n415) );
  XNOR U929 ( .A(b[424]), .B(n416), .Z(c[424]) );
  XOR U930 ( .A(n417), .B(n418), .Z(n414) );
  ANDN U931 ( .B(n419), .A(n420), .Z(n417) );
  XNOR U932 ( .A(b[423]), .B(n418), .Z(n419) );
  XNOR U933 ( .A(b[423]), .B(n420), .Z(c[423]) );
  XOR U934 ( .A(n421), .B(n422), .Z(n418) );
  ANDN U935 ( .B(n423), .A(n424), .Z(n421) );
  XNOR U936 ( .A(b[422]), .B(n422), .Z(n423) );
  XNOR U937 ( .A(b[422]), .B(n424), .Z(c[422]) );
  XOR U938 ( .A(n425), .B(n426), .Z(n422) );
  ANDN U939 ( .B(n427), .A(n428), .Z(n425) );
  XNOR U940 ( .A(b[421]), .B(n426), .Z(n427) );
  XNOR U941 ( .A(b[421]), .B(n428), .Z(c[421]) );
  XOR U942 ( .A(n429), .B(n430), .Z(n426) );
  ANDN U943 ( .B(n431), .A(n432), .Z(n429) );
  XNOR U944 ( .A(b[420]), .B(n430), .Z(n431) );
  XNOR U945 ( .A(b[420]), .B(n432), .Z(c[420]) );
  XOR U946 ( .A(n433), .B(n434), .Z(n430) );
  ANDN U947 ( .B(n435), .A(n436), .Z(n433) );
  XNOR U948 ( .A(b[419]), .B(n434), .Z(n435) );
  XNOR U949 ( .A(b[41]), .B(n437), .Z(c[41]) );
  XNOR U950 ( .A(b[419]), .B(n436), .Z(c[419]) );
  XOR U951 ( .A(n438), .B(n439), .Z(n434) );
  ANDN U952 ( .B(n440), .A(n441), .Z(n438) );
  XNOR U953 ( .A(b[418]), .B(n439), .Z(n440) );
  XNOR U954 ( .A(b[418]), .B(n441), .Z(c[418]) );
  XOR U955 ( .A(n442), .B(n443), .Z(n439) );
  ANDN U956 ( .B(n444), .A(n445), .Z(n442) );
  XNOR U957 ( .A(b[417]), .B(n443), .Z(n444) );
  XNOR U958 ( .A(b[417]), .B(n445), .Z(c[417]) );
  XOR U959 ( .A(n446), .B(n447), .Z(n443) );
  ANDN U960 ( .B(n448), .A(n449), .Z(n446) );
  XNOR U961 ( .A(b[416]), .B(n447), .Z(n448) );
  XNOR U962 ( .A(b[416]), .B(n449), .Z(c[416]) );
  XOR U963 ( .A(n450), .B(n451), .Z(n447) );
  ANDN U964 ( .B(n452), .A(n453), .Z(n450) );
  XNOR U965 ( .A(b[415]), .B(n451), .Z(n452) );
  XNOR U966 ( .A(b[415]), .B(n453), .Z(c[415]) );
  XOR U967 ( .A(n454), .B(n455), .Z(n451) );
  ANDN U968 ( .B(n456), .A(n457), .Z(n454) );
  XNOR U969 ( .A(b[414]), .B(n455), .Z(n456) );
  XNOR U970 ( .A(b[414]), .B(n457), .Z(c[414]) );
  XOR U971 ( .A(n458), .B(n459), .Z(n455) );
  ANDN U972 ( .B(n460), .A(n461), .Z(n458) );
  XNOR U973 ( .A(b[413]), .B(n459), .Z(n460) );
  XNOR U974 ( .A(b[413]), .B(n461), .Z(c[413]) );
  XOR U975 ( .A(n462), .B(n463), .Z(n459) );
  ANDN U976 ( .B(n464), .A(n465), .Z(n462) );
  XNOR U977 ( .A(b[412]), .B(n463), .Z(n464) );
  XNOR U978 ( .A(b[412]), .B(n465), .Z(c[412]) );
  XOR U979 ( .A(n466), .B(n467), .Z(n463) );
  ANDN U980 ( .B(n468), .A(n469), .Z(n466) );
  XNOR U981 ( .A(b[411]), .B(n467), .Z(n468) );
  XNOR U982 ( .A(b[411]), .B(n469), .Z(c[411]) );
  XOR U983 ( .A(n470), .B(n471), .Z(n467) );
  ANDN U984 ( .B(n472), .A(n473), .Z(n470) );
  XNOR U985 ( .A(b[410]), .B(n471), .Z(n472) );
  XNOR U986 ( .A(b[410]), .B(n473), .Z(c[410]) );
  XOR U987 ( .A(n474), .B(n475), .Z(n471) );
  ANDN U988 ( .B(n476), .A(n477), .Z(n474) );
  XNOR U989 ( .A(b[409]), .B(n475), .Z(n476) );
  XNOR U990 ( .A(b[40]), .B(n478), .Z(c[40]) );
  XNOR U991 ( .A(b[409]), .B(n477), .Z(c[409]) );
  XOR U992 ( .A(n479), .B(n480), .Z(n475) );
  ANDN U993 ( .B(n481), .A(n482), .Z(n479) );
  XNOR U994 ( .A(b[408]), .B(n480), .Z(n481) );
  XNOR U995 ( .A(b[408]), .B(n482), .Z(c[408]) );
  XOR U996 ( .A(n483), .B(n484), .Z(n480) );
  ANDN U997 ( .B(n485), .A(n486), .Z(n483) );
  XNOR U998 ( .A(b[407]), .B(n484), .Z(n485) );
  XNOR U999 ( .A(b[407]), .B(n486), .Z(c[407]) );
  XOR U1000 ( .A(n487), .B(n488), .Z(n484) );
  ANDN U1001 ( .B(n489), .A(n490), .Z(n487) );
  XNOR U1002 ( .A(b[406]), .B(n488), .Z(n489) );
  XNOR U1003 ( .A(b[406]), .B(n490), .Z(c[406]) );
  XOR U1004 ( .A(n491), .B(n492), .Z(n488) );
  ANDN U1005 ( .B(n493), .A(n494), .Z(n491) );
  XNOR U1006 ( .A(b[405]), .B(n492), .Z(n493) );
  XNOR U1007 ( .A(b[405]), .B(n494), .Z(c[405]) );
  XOR U1008 ( .A(n495), .B(n496), .Z(n492) );
  ANDN U1009 ( .B(n497), .A(n498), .Z(n495) );
  XNOR U1010 ( .A(b[404]), .B(n496), .Z(n497) );
  XNOR U1011 ( .A(b[404]), .B(n498), .Z(c[404]) );
  XOR U1012 ( .A(n499), .B(n500), .Z(n496) );
  ANDN U1013 ( .B(n501), .A(n502), .Z(n499) );
  XNOR U1014 ( .A(b[403]), .B(n500), .Z(n501) );
  XNOR U1015 ( .A(b[403]), .B(n502), .Z(c[403]) );
  XOR U1016 ( .A(n503), .B(n504), .Z(n500) );
  ANDN U1017 ( .B(n505), .A(n506), .Z(n503) );
  XNOR U1018 ( .A(b[402]), .B(n504), .Z(n505) );
  XNOR U1019 ( .A(b[402]), .B(n506), .Z(c[402]) );
  XOR U1020 ( .A(n507), .B(n508), .Z(n504) );
  ANDN U1021 ( .B(n509), .A(n510), .Z(n507) );
  XNOR U1022 ( .A(b[401]), .B(n508), .Z(n509) );
  XNOR U1023 ( .A(b[401]), .B(n510), .Z(c[401]) );
  XOR U1024 ( .A(n511), .B(n512), .Z(n508) );
  ANDN U1025 ( .B(n513), .A(n514), .Z(n511) );
  XNOR U1026 ( .A(b[400]), .B(n512), .Z(n513) );
  XNOR U1027 ( .A(b[400]), .B(n514), .Z(c[400]) );
  XOR U1028 ( .A(n515), .B(n516), .Z(n512) );
  ANDN U1029 ( .B(n517), .A(n518), .Z(n515) );
  XNOR U1030 ( .A(b[399]), .B(n516), .Z(n517) );
  XNOR U1031 ( .A(b[3]), .B(n519), .Z(c[3]) );
  XNOR U1032 ( .A(b[39]), .B(n520), .Z(c[39]) );
  XNOR U1033 ( .A(b[399]), .B(n518), .Z(c[399]) );
  XOR U1034 ( .A(n521), .B(n522), .Z(n516) );
  ANDN U1035 ( .B(n523), .A(n524), .Z(n521) );
  XNOR U1036 ( .A(b[398]), .B(n522), .Z(n523) );
  XNOR U1037 ( .A(b[398]), .B(n524), .Z(c[398]) );
  XOR U1038 ( .A(n525), .B(n526), .Z(n522) );
  ANDN U1039 ( .B(n527), .A(n528), .Z(n525) );
  XNOR U1040 ( .A(b[397]), .B(n526), .Z(n527) );
  XNOR U1041 ( .A(b[397]), .B(n528), .Z(c[397]) );
  XOR U1042 ( .A(n529), .B(n530), .Z(n526) );
  ANDN U1043 ( .B(n531), .A(n532), .Z(n529) );
  XNOR U1044 ( .A(b[396]), .B(n530), .Z(n531) );
  XNOR U1045 ( .A(b[396]), .B(n532), .Z(c[396]) );
  XOR U1046 ( .A(n533), .B(n534), .Z(n530) );
  ANDN U1047 ( .B(n535), .A(n536), .Z(n533) );
  XNOR U1048 ( .A(b[395]), .B(n534), .Z(n535) );
  XNOR U1049 ( .A(b[395]), .B(n536), .Z(c[395]) );
  XOR U1050 ( .A(n537), .B(n538), .Z(n534) );
  ANDN U1051 ( .B(n539), .A(n540), .Z(n537) );
  XNOR U1052 ( .A(b[394]), .B(n538), .Z(n539) );
  XNOR U1053 ( .A(b[394]), .B(n540), .Z(c[394]) );
  XOR U1054 ( .A(n541), .B(n542), .Z(n538) );
  ANDN U1055 ( .B(n543), .A(n544), .Z(n541) );
  XNOR U1056 ( .A(b[393]), .B(n542), .Z(n543) );
  XNOR U1057 ( .A(b[393]), .B(n544), .Z(c[393]) );
  XOR U1058 ( .A(n545), .B(n546), .Z(n542) );
  ANDN U1059 ( .B(n547), .A(n548), .Z(n545) );
  XNOR U1060 ( .A(b[392]), .B(n546), .Z(n547) );
  XNOR U1061 ( .A(b[392]), .B(n548), .Z(c[392]) );
  XOR U1062 ( .A(n549), .B(n550), .Z(n546) );
  ANDN U1063 ( .B(n551), .A(n552), .Z(n549) );
  XNOR U1064 ( .A(b[391]), .B(n550), .Z(n551) );
  XNOR U1065 ( .A(b[391]), .B(n552), .Z(c[391]) );
  XOR U1066 ( .A(n553), .B(n554), .Z(n550) );
  ANDN U1067 ( .B(n555), .A(n556), .Z(n553) );
  XNOR U1068 ( .A(b[390]), .B(n554), .Z(n555) );
  XNOR U1069 ( .A(b[390]), .B(n556), .Z(c[390]) );
  XOR U1070 ( .A(n557), .B(n558), .Z(n554) );
  ANDN U1071 ( .B(n559), .A(n560), .Z(n557) );
  XNOR U1072 ( .A(b[389]), .B(n558), .Z(n559) );
  XNOR U1073 ( .A(b[38]), .B(n561), .Z(c[38]) );
  XNOR U1074 ( .A(b[389]), .B(n560), .Z(c[389]) );
  XOR U1075 ( .A(n562), .B(n563), .Z(n558) );
  ANDN U1076 ( .B(n564), .A(n565), .Z(n562) );
  XNOR U1077 ( .A(b[388]), .B(n563), .Z(n564) );
  XNOR U1078 ( .A(b[388]), .B(n565), .Z(c[388]) );
  XOR U1079 ( .A(n566), .B(n567), .Z(n563) );
  ANDN U1080 ( .B(n568), .A(n569), .Z(n566) );
  XNOR U1081 ( .A(b[387]), .B(n567), .Z(n568) );
  XNOR U1082 ( .A(b[387]), .B(n569), .Z(c[387]) );
  XOR U1083 ( .A(n570), .B(n571), .Z(n567) );
  ANDN U1084 ( .B(n572), .A(n573), .Z(n570) );
  XNOR U1085 ( .A(b[386]), .B(n571), .Z(n572) );
  XNOR U1086 ( .A(b[386]), .B(n573), .Z(c[386]) );
  XOR U1087 ( .A(n574), .B(n575), .Z(n571) );
  ANDN U1088 ( .B(n576), .A(n577), .Z(n574) );
  XNOR U1089 ( .A(b[385]), .B(n575), .Z(n576) );
  XNOR U1090 ( .A(b[385]), .B(n577), .Z(c[385]) );
  XOR U1091 ( .A(n578), .B(n579), .Z(n575) );
  ANDN U1092 ( .B(n580), .A(n581), .Z(n578) );
  XNOR U1093 ( .A(b[384]), .B(n579), .Z(n580) );
  XNOR U1094 ( .A(b[384]), .B(n581), .Z(c[384]) );
  XOR U1095 ( .A(n582), .B(n583), .Z(n579) );
  ANDN U1096 ( .B(n584), .A(n585), .Z(n582) );
  XNOR U1097 ( .A(b[383]), .B(n583), .Z(n584) );
  XNOR U1098 ( .A(b[383]), .B(n585), .Z(c[383]) );
  XOR U1099 ( .A(n586), .B(n587), .Z(n583) );
  ANDN U1100 ( .B(n588), .A(n589), .Z(n586) );
  XNOR U1101 ( .A(b[382]), .B(n587), .Z(n588) );
  XNOR U1102 ( .A(b[382]), .B(n589), .Z(c[382]) );
  XOR U1103 ( .A(n590), .B(n591), .Z(n587) );
  ANDN U1104 ( .B(n592), .A(n593), .Z(n590) );
  XNOR U1105 ( .A(b[381]), .B(n591), .Z(n592) );
  XNOR U1106 ( .A(b[381]), .B(n593), .Z(c[381]) );
  XOR U1107 ( .A(n594), .B(n595), .Z(n591) );
  ANDN U1108 ( .B(n596), .A(n597), .Z(n594) );
  XNOR U1109 ( .A(b[380]), .B(n595), .Z(n596) );
  XNOR U1110 ( .A(b[380]), .B(n597), .Z(c[380]) );
  XOR U1111 ( .A(n598), .B(n599), .Z(n595) );
  ANDN U1112 ( .B(n600), .A(n601), .Z(n598) );
  XNOR U1113 ( .A(b[379]), .B(n599), .Z(n600) );
  XNOR U1114 ( .A(b[37]), .B(n602), .Z(c[37]) );
  XNOR U1115 ( .A(b[379]), .B(n601), .Z(c[379]) );
  XOR U1116 ( .A(n603), .B(n604), .Z(n599) );
  ANDN U1117 ( .B(n605), .A(n606), .Z(n603) );
  XNOR U1118 ( .A(b[378]), .B(n604), .Z(n605) );
  XNOR U1119 ( .A(b[378]), .B(n606), .Z(c[378]) );
  XOR U1120 ( .A(n607), .B(n608), .Z(n604) );
  ANDN U1121 ( .B(n609), .A(n610), .Z(n607) );
  XNOR U1122 ( .A(b[377]), .B(n608), .Z(n609) );
  XNOR U1123 ( .A(b[377]), .B(n610), .Z(c[377]) );
  XOR U1124 ( .A(n611), .B(n612), .Z(n608) );
  ANDN U1125 ( .B(n613), .A(n614), .Z(n611) );
  XNOR U1126 ( .A(b[376]), .B(n612), .Z(n613) );
  XNOR U1127 ( .A(b[376]), .B(n614), .Z(c[376]) );
  XOR U1128 ( .A(n615), .B(n616), .Z(n612) );
  ANDN U1129 ( .B(n617), .A(n618), .Z(n615) );
  XNOR U1130 ( .A(b[375]), .B(n616), .Z(n617) );
  XNOR U1131 ( .A(b[375]), .B(n618), .Z(c[375]) );
  XOR U1132 ( .A(n619), .B(n620), .Z(n616) );
  ANDN U1133 ( .B(n621), .A(n622), .Z(n619) );
  XNOR U1134 ( .A(b[374]), .B(n620), .Z(n621) );
  XNOR U1135 ( .A(b[374]), .B(n622), .Z(c[374]) );
  XOR U1136 ( .A(n623), .B(n624), .Z(n620) );
  ANDN U1137 ( .B(n625), .A(n626), .Z(n623) );
  XNOR U1138 ( .A(b[373]), .B(n624), .Z(n625) );
  XNOR U1139 ( .A(b[373]), .B(n626), .Z(c[373]) );
  XOR U1140 ( .A(n627), .B(n628), .Z(n624) );
  ANDN U1141 ( .B(n629), .A(n630), .Z(n627) );
  XNOR U1142 ( .A(b[372]), .B(n628), .Z(n629) );
  XNOR U1143 ( .A(b[372]), .B(n630), .Z(c[372]) );
  XOR U1144 ( .A(n631), .B(n632), .Z(n628) );
  ANDN U1145 ( .B(n633), .A(n634), .Z(n631) );
  XNOR U1146 ( .A(b[371]), .B(n632), .Z(n633) );
  XNOR U1147 ( .A(b[371]), .B(n634), .Z(c[371]) );
  XOR U1148 ( .A(n635), .B(n636), .Z(n632) );
  ANDN U1149 ( .B(n637), .A(n638), .Z(n635) );
  XNOR U1150 ( .A(b[370]), .B(n636), .Z(n637) );
  XNOR U1151 ( .A(b[370]), .B(n638), .Z(c[370]) );
  XOR U1152 ( .A(n639), .B(n640), .Z(n636) );
  ANDN U1153 ( .B(n641), .A(n642), .Z(n639) );
  XNOR U1154 ( .A(b[369]), .B(n640), .Z(n641) );
  XNOR U1155 ( .A(b[36]), .B(n643), .Z(c[36]) );
  XNOR U1156 ( .A(b[369]), .B(n642), .Z(c[369]) );
  XOR U1157 ( .A(n644), .B(n645), .Z(n640) );
  ANDN U1158 ( .B(n646), .A(n647), .Z(n644) );
  XNOR U1159 ( .A(b[368]), .B(n645), .Z(n646) );
  XNOR U1160 ( .A(b[368]), .B(n647), .Z(c[368]) );
  XOR U1161 ( .A(n648), .B(n649), .Z(n645) );
  ANDN U1162 ( .B(n650), .A(n651), .Z(n648) );
  XNOR U1163 ( .A(b[367]), .B(n649), .Z(n650) );
  XNOR U1164 ( .A(b[367]), .B(n651), .Z(c[367]) );
  XOR U1165 ( .A(n652), .B(n653), .Z(n649) );
  ANDN U1166 ( .B(n654), .A(n655), .Z(n652) );
  XNOR U1167 ( .A(b[366]), .B(n653), .Z(n654) );
  XNOR U1168 ( .A(b[366]), .B(n655), .Z(c[366]) );
  XOR U1169 ( .A(n656), .B(n657), .Z(n653) );
  ANDN U1170 ( .B(n658), .A(n659), .Z(n656) );
  XNOR U1171 ( .A(b[365]), .B(n657), .Z(n658) );
  XNOR U1172 ( .A(b[365]), .B(n659), .Z(c[365]) );
  XOR U1173 ( .A(n660), .B(n661), .Z(n657) );
  ANDN U1174 ( .B(n662), .A(n663), .Z(n660) );
  XNOR U1175 ( .A(b[364]), .B(n661), .Z(n662) );
  XNOR U1176 ( .A(b[364]), .B(n663), .Z(c[364]) );
  XOR U1177 ( .A(n664), .B(n665), .Z(n661) );
  ANDN U1178 ( .B(n666), .A(n667), .Z(n664) );
  XNOR U1179 ( .A(b[363]), .B(n665), .Z(n666) );
  XNOR U1180 ( .A(b[363]), .B(n667), .Z(c[363]) );
  XOR U1181 ( .A(n668), .B(n669), .Z(n665) );
  ANDN U1182 ( .B(n670), .A(n671), .Z(n668) );
  XNOR U1183 ( .A(b[362]), .B(n669), .Z(n670) );
  XNOR U1184 ( .A(b[362]), .B(n671), .Z(c[362]) );
  XOR U1185 ( .A(n672), .B(n673), .Z(n669) );
  ANDN U1186 ( .B(n674), .A(n675), .Z(n672) );
  XNOR U1187 ( .A(b[361]), .B(n673), .Z(n674) );
  XNOR U1188 ( .A(b[361]), .B(n675), .Z(c[361]) );
  XOR U1189 ( .A(n676), .B(n677), .Z(n673) );
  ANDN U1190 ( .B(n678), .A(n679), .Z(n676) );
  XNOR U1191 ( .A(b[360]), .B(n677), .Z(n678) );
  XNOR U1192 ( .A(b[360]), .B(n679), .Z(c[360]) );
  XOR U1193 ( .A(n680), .B(n681), .Z(n677) );
  ANDN U1194 ( .B(n682), .A(n683), .Z(n680) );
  XNOR U1195 ( .A(b[359]), .B(n681), .Z(n682) );
  XNOR U1196 ( .A(b[35]), .B(n684), .Z(c[35]) );
  XNOR U1197 ( .A(b[359]), .B(n683), .Z(c[359]) );
  XOR U1198 ( .A(n685), .B(n686), .Z(n681) );
  ANDN U1199 ( .B(n687), .A(n688), .Z(n685) );
  XNOR U1200 ( .A(b[358]), .B(n686), .Z(n687) );
  XNOR U1201 ( .A(b[358]), .B(n688), .Z(c[358]) );
  XOR U1202 ( .A(n689), .B(n690), .Z(n686) );
  ANDN U1203 ( .B(n691), .A(n692), .Z(n689) );
  XNOR U1204 ( .A(b[357]), .B(n690), .Z(n691) );
  XNOR U1205 ( .A(b[357]), .B(n692), .Z(c[357]) );
  XOR U1206 ( .A(n693), .B(n694), .Z(n690) );
  ANDN U1207 ( .B(n695), .A(n696), .Z(n693) );
  XNOR U1208 ( .A(b[356]), .B(n694), .Z(n695) );
  XNOR U1209 ( .A(b[356]), .B(n696), .Z(c[356]) );
  XOR U1210 ( .A(n697), .B(n698), .Z(n694) );
  ANDN U1211 ( .B(n699), .A(n700), .Z(n697) );
  XNOR U1212 ( .A(b[355]), .B(n698), .Z(n699) );
  XNOR U1213 ( .A(b[355]), .B(n700), .Z(c[355]) );
  XOR U1214 ( .A(n701), .B(n702), .Z(n698) );
  ANDN U1215 ( .B(n703), .A(n704), .Z(n701) );
  XNOR U1216 ( .A(b[354]), .B(n702), .Z(n703) );
  XNOR U1217 ( .A(b[354]), .B(n704), .Z(c[354]) );
  XOR U1218 ( .A(n705), .B(n706), .Z(n702) );
  ANDN U1219 ( .B(n707), .A(n708), .Z(n705) );
  XNOR U1220 ( .A(b[353]), .B(n706), .Z(n707) );
  XNOR U1221 ( .A(b[353]), .B(n708), .Z(c[353]) );
  XOR U1222 ( .A(n709), .B(n710), .Z(n706) );
  ANDN U1223 ( .B(n711), .A(n712), .Z(n709) );
  XNOR U1224 ( .A(b[352]), .B(n710), .Z(n711) );
  XNOR U1225 ( .A(b[352]), .B(n712), .Z(c[352]) );
  XOR U1226 ( .A(n713), .B(n714), .Z(n710) );
  ANDN U1227 ( .B(n715), .A(n716), .Z(n713) );
  XNOR U1228 ( .A(b[351]), .B(n714), .Z(n715) );
  XNOR U1229 ( .A(b[351]), .B(n716), .Z(c[351]) );
  XOR U1230 ( .A(n717), .B(n718), .Z(n714) );
  ANDN U1231 ( .B(n719), .A(n720), .Z(n717) );
  XNOR U1232 ( .A(b[350]), .B(n718), .Z(n719) );
  XNOR U1233 ( .A(b[350]), .B(n720), .Z(c[350]) );
  XOR U1234 ( .A(n721), .B(n722), .Z(n718) );
  ANDN U1235 ( .B(n723), .A(n724), .Z(n721) );
  XNOR U1236 ( .A(b[349]), .B(n722), .Z(n723) );
  XNOR U1237 ( .A(b[34]), .B(n725), .Z(c[34]) );
  XNOR U1238 ( .A(b[349]), .B(n724), .Z(c[349]) );
  XOR U1239 ( .A(n726), .B(n727), .Z(n722) );
  ANDN U1240 ( .B(n728), .A(n729), .Z(n726) );
  XNOR U1241 ( .A(b[348]), .B(n727), .Z(n728) );
  XNOR U1242 ( .A(b[348]), .B(n729), .Z(c[348]) );
  XOR U1243 ( .A(n730), .B(n731), .Z(n727) );
  ANDN U1244 ( .B(n732), .A(n733), .Z(n730) );
  XNOR U1245 ( .A(b[347]), .B(n731), .Z(n732) );
  XNOR U1246 ( .A(b[347]), .B(n733), .Z(c[347]) );
  XOR U1247 ( .A(n734), .B(n735), .Z(n731) );
  ANDN U1248 ( .B(n736), .A(n737), .Z(n734) );
  XNOR U1249 ( .A(b[346]), .B(n735), .Z(n736) );
  XNOR U1250 ( .A(b[346]), .B(n737), .Z(c[346]) );
  XOR U1251 ( .A(n738), .B(n739), .Z(n735) );
  ANDN U1252 ( .B(n740), .A(n741), .Z(n738) );
  XNOR U1253 ( .A(b[345]), .B(n739), .Z(n740) );
  XNOR U1254 ( .A(b[345]), .B(n741), .Z(c[345]) );
  XOR U1255 ( .A(n742), .B(n743), .Z(n739) );
  ANDN U1256 ( .B(n744), .A(n745), .Z(n742) );
  XNOR U1257 ( .A(b[344]), .B(n743), .Z(n744) );
  XNOR U1258 ( .A(b[344]), .B(n745), .Z(c[344]) );
  XOR U1259 ( .A(n746), .B(n747), .Z(n743) );
  ANDN U1260 ( .B(n748), .A(n749), .Z(n746) );
  XNOR U1261 ( .A(b[343]), .B(n747), .Z(n748) );
  XNOR U1262 ( .A(b[343]), .B(n749), .Z(c[343]) );
  XOR U1263 ( .A(n750), .B(n751), .Z(n747) );
  ANDN U1264 ( .B(n752), .A(n753), .Z(n750) );
  XNOR U1265 ( .A(b[342]), .B(n751), .Z(n752) );
  XNOR U1266 ( .A(b[342]), .B(n753), .Z(c[342]) );
  XOR U1267 ( .A(n754), .B(n755), .Z(n751) );
  ANDN U1268 ( .B(n756), .A(n757), .Z(n754) );
  XNOR U1269 ( .A(b[341]), .B(n755), .Z(n756) );
  XNOR U1270 ( .A(b[341]), .B(n757), .Z(c[341]) );
  XOR U1271 ( .A(n758), .B(n759), .Z(n755) );
  ANDN U1272 ( .B(n760), .A(n761), .Z(n758) );
  XNOR U1273 ( .A(b[340]), .B(n759), .Z(n760) );
  XNOR U1274 ( .A(b[340]), .B(n761), .Z(c[340]) );
  XOR U1275 ( .A(n762), .B(n763), .Z(n759) );
  ANDN U1276 ( .B(n764), .A(n765), .Z(n762) );
  XNOR U1277 ( .A(b[339]), .B(n763), .Z(n764) );
  XNOR U1278 ( .A(b[33]), .B(n766), .Z(c[33]) );
  XNOR U1279 ( .A(b[339]), .B(n765), .Z(c[339]) );
  XOR U1280 ( .A(n767), .B(n768), .Z(n763) );
  ANDN U1281 ( .B(n769), .A(n770), .Z(n767) );
  XNOR U1282 ( .A(b[338]), .B(n768), .Z(n769) );
  XNOR U1283 ( .A(b[338]), .B(n770), .Z(c[338]) );
  XOR U1284 ( .A(n771), .B(n772), .Z(n768) );
  ANDN U1285 ( .B(n773), .A(n774), .Z(n771) );
  XNOR U1286 ( .A(b[337]), .B(n772), .Z(n773) );
  XNOR U1287 ( .A(b[337]), .B(n774), .Z(c[337]) );
  XOR U1288 ( .A(n775), .B(n776), .Z(n772) );
  ANDN U1289 ( .B(n777), .A(n778), .Z(n775) );
  XNOR U1290 ( .A(b[336]), .B(n776), .Z(n777) );
  XNOR U1291 ( .A(b[336]), .B(n778), .Z(c[336]) );
  XOR U1292 ( .A(n779), .B(n780), .Z(n776) );
  ANDN U1293 ( .B(n781), .A(n782), .Z(n779) );
  XNOR U1294 ( .A(b[335]), .B(n780), .Z(n781) );
  XNOR U1295 ( .A(b[335]), .B(n782), .Z(c[335]) );
  XOR U1296 ( .A(n783), .B(n784), .Z(n780) );
  ANDN U1297 ( .B(n785), .A(n786), .Z(n783) );
  XNOR U1298 ( .A(b[334]), .B(n784), .Z(n785) );
  XNOR U1299 ( .A(b[334]), .B(n786), .Z(c[334]) );
  XOR U1300 ( .A(n787), .B(n788), .Z(n784) );
  ANDN U1301 ( .B(n789), .A(n790), .Z(n787) );
  XNOR U1302 ( .A(b[333]), .B(n788), .Z(n789) );
  XNOR U1303 ( .A(b[333]), .B(n790), .Z(c[333]) );
  XOR U1304 ( .A(n791), .B(n792), .Z(n788) );
  ANDN U1305 ( .B(n793), .A(n794), .Z(n791) );
  XNOR U1306 ( .A(b[332]), .B(n792), .Z(n793) );
  XNOR U1307 ( .A(b[332]), .B(n794), .Z(c[332]) );
  XOR U1308 ( .A(n795), .B(n796), .Z(n792) );
  ANDN U1309 ( .B(n797), .A(n798), .Z(n795) );
  XNOR U1310 ( .A(b[331]), .B(n796), .Z(n797) );
  XNOR U1311 ( .A(b[331]), .B(n798), .Z(c[331]) );
  XOR U1312 ( .A(n799), .B(n800), .Z(n796) );
  ANDN U1313 ( .B(n801), .A(n802), .Z(n799) );
  XNOR U1314 ( .A(b[330]), .B(n800), .Z(n801) );
  XNOR U1315 ( .A(b[330]), .B(n802), .Z(c[330]) );
  XOR U1316 ( .A(n803), .B(n804), .Z(n800) );
  ANDN U1317 ( .B(n805), .A(n806), .Z(n803) );
  XNOR U1318 ( .A(b[329]), .B(n804), .Z(n805) );
  XNOR U1319 ( .A(b[32]), .B(n807), .Z(c[32]) );
  XNOR U1320 ( .A(b[329]), .B(n806), .Z(c[329]) );
  XOR U1321 ( .A(n808), .B(n809), .Z(n804) );
  ANDN U1322 ( .B(n810), .A(n811), .Z(n808) );
  XNOR U1323 ( .A(b[328]), .B(n809), .Z(n810) );
  XNOR U1324 ( .A(b[328]), .B(n811), .Z(c[328]) );
  XOR U1325 ( .A(n812), .B(n813), .Z(n809) );
  ANDN U1326 ( .B(n814), .A(n815), .Z(n812) );
  XNOR U1327 ( .A(b[327]), .B(n813), .Z(n814) );
  XNOR U1328 ( .A(b[327]), .B(n815), .Z(c[327]) );
  XOR U1329 ( .A(n816), .B(n817), .Z(n813) );
  ANDN U1330 ( .B(n818), .A(n819), .Z(n816) );
  XNOR U1331 ( .A(b[326]), .B(n817), .Z(n818) );
  XNOR U1332 ( .A(b[326]), .B(n819), .Z(c[326]) );
  XOR U1333 ( .A(n820), .B(n821), .Z(n817) );
  ANDN U1334 ( .B(n822), .A(n823), .Z(n820) );
  XNOR U1335 ( .A(b[325]), .B(n821), .Z(n822) );
  XNOR U1336 ( .A(b[325]), .B(n823), .Z(c[325]) );
  XOR U1337 ( .A(n824), .B(n825), .Z(n821) );
  ANDN U1338 ( .B(n826), .A(n827), .Z(n824) );
  XNOR U1339 ( .A(b[324]), .B(n825), .Z(n826) );
  XNOR U1340 ( .A(b[324]), .B(n827), .Z(c[324]) );
  XOR U1341 ( .A(n828), .B(n829), .Z(n825) );
  ANDN U1342 ( .B(n830), .A(n831), .Z(n828) );
  XNOR U1343 ( .A(b[323]), .B(n829), .Z(n830) );
  XNOR U1344 ( .A(b[323]), .B(n831), .Z(c[323]) );
  XOR U1345 ( .A(n832), .B(n833), .Z(n829) );
  ANDN U1346 ( .B(n834), .A(n835), .Z(n832) );
  XNOR U1347 ( .A(b[322]), .B(n833), .Z(n834) );
  XNOR U1348 ( .A(b[322]), .B(n835), .Z(c[322]) );
  XOR U1349 ( .A(n836), .B(n837), .Z(n833) );
  ANDN U1350 ( .B(n838), .A(n839), .Z(n836) );
  XNOR U1351 ( .A(b[321]), .B(n837), .Z(n838) );
  XNOR U1352 ( .A(b[321]), .B(n839), .Z(c[321]) );
  XOR U1353 ( .A(n840), .B(n841), .Z(n837) );
  ANDN U1354 ( .B(n842), .A(n843), .Z(n840) );
  XNOR U1355 ( .A(b[320]), .B(n841), .Z(n842) );
  XNOR U1356 ( .A(b[320]), .B(n843), .Z(c[320]) );
  XOR U1357 ( .A(n844), .B(n845), .Z(n841) );
  ANDN U1358 ( .B(n846), .A(n847), .Z(n844) );
  XNOR U1359 ( .A(b[319]), .B(n845), .Z(n846) );
  XNOR U1360 ( .A(b[31]), .B(n848), .Z(c[31]) );
  XNOR U1361 ( .A(b[319]), .B(n847), .Z(c[319]) );
  XOR U1362 ( .A(n849), .B(n850), .Z(n845) );
  ANDN U1363 ( .B(n851), .A(n852), .Z(n849) );
  XNOR U1364 ( .A(b[318]), .B(n850), .Z(n851) );
  XNOR U1365 ( .A(b[318]), .B(n852), .Z(c[318]) );
  XOR U1366 ( .A(n853), .B(n854), .Z(n850) );
  ANDN U1367 ( .B(n855), .A(n856), .Z(n853) );
  XNOR U1368 ( .A(b[317]), .B(n854), .Z(n855) );
  XNOR U1369 ( .A(b[317]), .B(n856), .Z(c[317]) );
  XOR U1370 ( .A(n857), .B(n858), .Z(n854) );
  ANDN U1371 ( .B(n859), .A(n860), .Z(n857) );
  XNOR U1372 ( .A(b[316]), .B(n858), .Z(n859) );
  XNOR U1373 ( .A(b[316]), .B(n860), .Z(c[316]) );
  XOR U1374 ( .A(n861), .B(n862), .Z(n858) );
  ANDN U1375 ( .B(n863), .A(n864), .Z(n861) );
  XNOR U1376 ( .A(b[315]), .B(n862), .Z(n863) );
  XNOR U1377 ( .A(b[315]), .B(n864), .Z(c[315]) );
  XOR U1378 ( .A(n865), .B(n866), .Z(n862) );
  ANDN U1379 ( .B(n867), .A(n868), .Z(n865) );
  XNOR U1380 ( .A(b[314]), .B(n866), .Z(n867) );
  XNOR U1381 ( .A(b[314]), .B(n868), .Z(c[314]) );
  XOR U1382 ( .A(n869), .B(n870), .Z(n866) );
  ANDN U1383 ( .B(n871), .A(n872), .Z(n869) );
  XNOR U1384 ( .A(b[313]), .B(n870), .Z(n871) );
  XNOR U1385 ( .A(b[313]), .B(n872), .Z(c[313]) );
  XOR U1386 ( .A(n873), .B(n874), .Z(n870) );
  ANDN U1387 ( .B(n875), .A(n876), .Z(n873) );
  XNOR U1388 ( .A(b[312]), .B(n874), .Z(n875) );
  XNOR U1389 ( .A(b[312]), .B(n876), .Z(c[312]) );
  XOR U1390 ( .A(n877), .B(n878), .Z(n874) );
  ANDN U1391 ( .B(n879), .A(n880), .Z(n877) );
  XNOR U1392 ( .A(b[311]), .B(n878), .Z(n879) );
  XNOR U1393 ( .A(b[311]), .B(n880), .Z(c[311]) );
  XOR U1394 ( .A(n881), .B(n882), .Z(n878) );
  ANDN U1395 ( .B(n883), .A(n884), .Z(n881) );
  XNOR U1396 ( .A(b[310]), .B(n882), .Z(n883) );
  XNOR U1397 ( .A(b[310]), .B(n884), .Z(c[310]) );
  XOR U1398 ( .A(n885), .B(n886), .Z(n882) );
  ANDN U1399 ( .B(n887), .A(n888), .Z(n885) );
  XNOR U1400 ( .A(b[309]), .B(n886), .Z(n887) );
  XNOR U1401 ( .A(b[30]), .B(n889), .Z(c[30]) );
  XNOR U1402 ( .A(b[309]), .B(n888), .Z(c[309]) );
  XOR U1403 ( .A(n890), .B(n891), .Z(n886) );
  ANDN U1404 ( .B(n892), .A(n893), .Z(n890) );
  XNOR U1405 ( .A(b[308]), .B(n891), .Z(n892) );
  XNOR U1406 ( .A(b[308]), .B(n893), .Z(c[308]) );
  XOR U1407 ( .A(n894), .B(n895), .Z(n891) );
  ANDN U1408 ( .B(n896), .A(n897), .Z(n894) );
  XNOR U1409 ( .A(b[307]), .B(n895), .Z(n896) );
  XNOR U1410 ( .A(b[307]), .B(n897), .Z(c[307]) );
  XOR U1411 ( .A(n898), .B(n899), .Z(n895) );
  ANDN U1412 ( .B(n900), .A(n901), .Z(n898) );
  XNOR U1413 ( .A(b[306]), .B(n899), .Z(n900) );
  XNOR U1414 ( .A(b[306]), .B(n901), .Z(c[306]) );
  XOR U1415 ( .A(n902), .B(n903), .Z(n899) );
  ANDN U1416 ( .B(n904), .A(n905), .Z(n902) );
  XNOR U1417 ( .A(b[305]), .B(n903), .Z(n904) );
  XNOR U1418 ( .A(b[305]), .B(n905), .Z(c[305]) );
  XOR U1419 ( .A(n906), .B(n907), .Z(n903) );
  ANDN U1420 ( .B(n908), .A(n909), .Z(n906) );
  XNOR U1421 ( .A(b[304]), .B(n907), .Z(n908) );
  XNOR U1422 ( .A(b[304]), .B(n909), .Z(c[304]) );
  XOR U1423 ( .A(n910), .B(n911), .Z(n907) );
  ANDN U1424 ( .B(n912), .A(n913), .Z(n910) );
  XNOR U1425 ( .A(b[303]), .B(n911), .Z(n912) );
  XNOR U1426 ( .A(b[303]), .B(n913), .Z(c[303]) );
  XOR U1427 ( .A(n914), .B(n915), .Z(n911) );
  ANDN U1428 ( .B(n916), .A(n917), .Z(n914) );
  XNOR U1429 ( .A(b[302]), .B(n915), .Z(n916) );
  XNOR U1430 ( .A(b[302]), .B(n917), .Z(c[302]) );
  XOR U1431 ( .A(n918), .B(n919), .Z(n915) );
  ANDN U1432 ( .B(n920), .A(n921), .Z(n918) );
  XNOR U1433 ( .A(b[301]), .B(n919), .Z(n920) );
  XNOR U1434 ( .A(b[301]), .B(n921), .Z(c[301]) );
  XOR U1435 ( .A(n922), .B(n923), .Z(n919) );
  ANDN U1436 ( .B(n924), .A(n925), .Z(n922) );
  XNOR U1437 ( .A(b[300]), .B(n923), .Z(n924) );
  XNOR U1438 ( .A(b[300]), .B(n925), .Z(c[300]) );
  XOR U1439 ( .A(n926), .B(n927), .Z(n923) );
  ANDN U1440 ( .B(n928), .A(n929), .Z(n926) );
  XNOR U1441 ( .A(b[299]), .B(n927), .Z(n928) );
  XNOR U1442 ( .A(b[2]), .B(n930), .Z(c[2]) );
  XNOR U1443 ( .A(b[29]), .B(n931), .Z(c[29]) );
  XNOR U1444 ( .A(b[299]), .B(n929), .Z(c[299]) );
  XOR U1445 ( .A(n932), .B(n933), .Z(n927) );
  ANDN U1446 ( .B(n934), .A(n935), .Z(n932) );
  XNOR U1447 ( .A(b[298]), .B(n933), .Z(n934) );
  XNOR U1448 ( .A(b[298]), .B(n935), .Z(c[298]) );
  XOR U1449 ( .A(n936), .B(n937), .Z(n933) );
  ANDN U1450 ( .B(n938), .A(n939), .Z(n936) );
  XNOR U1451 ( .A(b[297]), .B(n937), .Z(n938) );
  XNOR U1452 ( .A(b[297]), .B(n939), .Z(c[297]) );
  XOR U1453 ( .A(n940), .B(n941), .Z(n937) );
  ANDN U1454 ( .B(n942), .A(n943), .Z(n940) );
  XNOR U1455 ( .A(b[296]), .B(n941), .Z(n942) );
  XNOR U1456 ( .A(b[296]), .B(n943), .Z(c[296]) );
  XOR U1457 ( .A(n944), .B(n945), .Z(n941) );
  ANDN U1458 ( .B(n946), .A(n947), .Z(n944) );
  XNOR U1459 ( .A(b[295]), .B(n945), .Z(n946) );
  XNOR U1460 ( .A(b[295]), .B(n947), .Z(c[295]) );
  XOR U1461 ( .A(n948), .B(n949), .Z(n945) );
  ANDN U1462 ( .B(n950), .A(n951), .Z(n948) );
  XNOR U1463 ( .A(b[294]), .B(n949), .Z(n950) );
  XNOR U1464 ( .A(b[294]), .B(n951), .Z(c[294]) );
  XOR U1465 ( .A(n952), .B(n953), .Z(n949) );
  ANDN U1466 ( .B(n954), .A(n955), .Z(n952) );
  XNOR U1467 ( .A(b[293]), .B(n953), .Z(n954) );
  XNOR U1468 ( .A(b[293]), .B(n955), .Z(c[293]) );
  XOR U1469 ( .A(n956), .B(n957), .Z(n953) );
  ANDN U1470 ( .B(n958), .A(n959), .Z(n956) );
  XNOR U1471 ( .A(b[292]), .B(n957), .Z(n958) );
  XNOR U1472 ( .A(b[292]), .B(n959), .Z(c[292]) );
  XOR U1473 ( .A(n960), .B(n961), .Z(n957) );
  ANDN U1474 ( .B(n962), .A(n963), .Z(n960) );
  XNOR U1475 ( .A(b[291]), .B(n961), .Z(n962) );
  XNOR U1476 ( .A(b[291]), .B(n963), .Z(c[291]) );
  XOR U1477 ( .A(n964), .B(n965), .Z(n961) );
  ANDN U1478 ( .B(n966), .A(n967), .Z(n964) );
  XNOR U1479 ( .A(b[290]), .B(n965), .Z(n966) );
  XNOR U1480 ( .A(b[290]), .B(n967), .Z(c[290]) );
  XOR U1481 ( .A(n968), .B(n969), .Z(n965) );
  ANDN U1482 ( .B(n970), .A(n971), .Z(n968) );
  XNOR U1483 ( .A(b[289]), .B(n969), .Z(n970) );
  XNOR U1484 ( .A(b[28]), .B(n972), .Z(c[28]) );
  XNOR U1485 ( .A(b[289]), .B(n971), .Z(c[289]) );
  XOR U1486 ( .A(n973), .B(n974), .Z(n969) );
  ANDN U1487 ( .B(n975), .A(n976), .Z(n973) );
  XNOR U1488 ( .A(b[288]), .B(n974), .Z(n975) );
  XNOR U1489 ( .A(b[288]), .B(n976), .Z(c[288]) );
  XOR U1490 ( .A(n977), .B(n978), .Z(n974) );
  ANDN U1491 ( .B(n979), .A(n980), .Z(n977) );
  XNOR U1492 ( .A(b[287]), .B(n978), .Z(n979) );
  XNOR U1493 ( .A(b[287]), .B(n980), .Z(c[287]) );
  XOR U1494 ( .A(n981), .B(n982), .Z(n978) );
  ANDN U1495 ( .B(n983), .A(n984), .Z(n981) );
  XNOR U1496 ( .A(b[286]), .B(n982), .Z(n983) );
  XNOR U1497 ( .A(b[286]), .B(n984), .Z(c[286]) );
  XOR U1498 ( .A(n985), .B(n986), .Z(n982) );
  ANDN U1499 ( .B(n987), .A(n988), .Z(n985) );
  XNOR U1500 ( .A(b[285]), .B(n986), .Z(n987) );
  XNOR U1501 ( .A(b[285]), .B(n988), .Z(c[285]) );
  XOR U1502 ( .A(n989), .B(n990), .Z(n986) );
  ANDN U1503 ( .B(n991), .A(n992), .Z(n989) );
  XNOR U1504 ( .A(b[284]), .B(n990), .Z(n991) );
  XNOR U1505 ( .A(b[284]), .B(n992), .Z(c[284]) );
  XOR U1506 ( .A(n993), .B(n994), .Z(n990) );
  ANDN U1507 ( .B(n995), .A(n996), .Z(n993) );
  XNOR U1508 ( .A(b[283]), .B(n994), .Z(n995) );
  XNOR U1509 ( .A(b[283]), .B(n996), .Z(c[283]) );
  XOR U1510 ( .A(n997), .B(n998), .Z(n994) );
  ANDN U1511 ( .B(n999), .A(n1000), .Z(n997) );
  XNOR U1512 ( .A(b[282]), .B(n998), .Z(n999) );
  XNOR U1513 ( .A(b[282]), .B(n1000), .Z(c[282]) );
  XOR U1514 ( .A(n1001), .B(n1002), .Z(n998) );
  ANDN U1515 ( .B(n1003), .A(n1004), .Z(n1001) );
  XNOR U1516 ( .A(b[281]), .B(n1002), .Z(n1003) );
  XNOR U1517 ( .A(b[281]), .B(n1004), .Z(c[281]) );
  XOR U1518 ( .A(n1005), .B(n1006), .Z(n1002) );
  ANDN U1519 ( .B(n1007), .A(n1008), .Z(n1005) );
  XNOR U1520 ( .A(b[280]), .B(n1006), .Z(n1007) );
  XNOR U1521 ( .A(b[280]), .B(n1008), .Z(c[280]) );
  XOR U1522 ( .A(n1009), .B(n1010), .Z(n1006) );
  ANDN U1523 ( .B(n1011), .A(n1012), .Z(n1009) );
  XNOR U1524 ( .A(b[279]), .B(n1010), .Z(n1011) );
  XNOR U1525 ( .A(b[27]), .B(n1013), .Z(c[27]) );
  XNOR U1526 ( .A(b[279]), .B(n1012), .Z(c[279]) );
  XOR U1527 ( .A(n1014), .B(n1015), .Z(n1010) );
  ANDN U1528 ( .B(n1016), .A(n1017), .Z(n1014) );
  XNOR U1529 ( .A(b[278]), .B(n1015), .Z(n1016) );
  XNOR U1530 ( .A(b[278]), .B(n1017), .Z(c[278]) );
  XOR U1531 ( .A(n1018), .B(n1019), .Z(n1015) );
  ANDN U1532 ( .B(n1020), .A(n1021), .Z(n1018) );
  XNOR U1533 ( .A(b[277]), .B(n1019), .Z(n1020) );
  XNOR U1534 ( .A(b[277]), .B(n1021), .Z(c[277]) );
  XOR U1535 ( .A(n1022), .B(n1023), .Z(n1019) );
  ANDN U1536 ( .B(n1024), .A(n1025), .Z(n1022) );
  XNOR U1537 ( .A(b[276]), .B(n1023), .Z(n1024) );
  XNOR U1538 ( .A(b[276]), .B(n1025), .Z(c[276]) );
  XOR U1539 ( .A(n1026), .B(n1027), .Z(n1023) );
  ANDN U1540 ( .B(n1028), .A(n1029), .Z(n1026) );
  XNOR U1541 ( .A(b[275]), .B(n1027), .Z(n1028) );
  XNOR U1542 ( .A(b[275]), .B(n1029), .Z(c[275]) );
  XOR U1543 ( .A(n1030), .B(n1031), .Z(n1027) );
  ANDN U1544 ( .B(n1032), .A(n1033), .Z(n1030) );
  XNOR U1545 ( .A(b[274]), .B(n1031), .Z(n1032) );
  XNOR U1546 ( .A(b[274]), .B(n1033), .Z(c[274]) );
  XOR U1547 ( .A(n1034), .B(n1035), .Z(n1031) );
  ANDN U1548 ( .B(n1036), .A(n1037), .Z(n1034) );
  XNOR U1549 ( .A(b[273]), .B(n1035), .Z(n1036) );
  XNOR U1550 ( .A(b[273]), .B(n1037), .Z(c[273]) );
  XOR U1551 ( .A(n1038), .B(n1039), .Z(n1035) );
  ANDN U1552 ( .B(n1040), .A(n1041), .Z(n1038) );
  XNOR U1553 ( .A(b[272]), .B(n1039), .Z(n1040) );
  XNOR U1554 ( .A(b[272]), .B(n1041), .Z(c[272]) );
  XOR U1555 ( .A(n1042), .B(n1043), .Z(n1039) );
  ANDN U1556 ( .B(n1044), .A(n1045), .Z(n1042) );
  XNOR U1557 ( .A(b[271]), .B(n1043), .Z(n1044) );
  XNOR U1558 ( .A(b[271]), .B(n1045), .Z(c[271]) );
  XOR U1559 ( .A(n1046), .B(n1047), .Z(n1043) );
  ANDN U1560 ( .B(n1048), .A(n1049), .Z(n1046) );
  XNOR U1561 ( .A(b[270]), .B(n1047), .Z(n1048) );
  XNOR U1562 ( .A(b[270]), .B(n1049), .Z(c[270]) );
  XOR U1563 ( .A(n1050), .B(n1051), .Z(n1047) );
  ANDN U1564 ( .B(n1052), .A(n1053), .Z(n1050) );
  XNOR U1565 ( .A(b[269]), .B(n1051), .Z(n1052) );
  XNOR U1566 ( .A(b[26]), .B(n1054), .Z(c[26]) );
  XNOR U1567 ( .A(b[269]), .B(n1053), .Z(c[269]) );
  XOR U1568 ( .A(n1055), .B(n1056), .Z(n1051) );
  ANDN U1569 ( .B(n1057), .A(n1058), .Z(n1055) );
  XNOR U1570 ( .A(b[268]), .B(n1056), .Z(n1057) );
  XNOR U1571 ( .A(b[268]), .B(n1058), .Z(c[268]) );
  XOR U1572 ( .A(n1059), .B(n1060), .Z(n1056) );
  ANDN U1573 ( .B(n1061), .A(n1062), .Z(n1059) );
  XNOR U1574 ( .A(b[267]), .B(n1060), .Z(n1061) );
  XNOR U1575 ( .A(b[267]), .B(n1062), .Z(c[267]) );
  XOR U1576 ( .A(n1063), .B(n1064), .Z(n1060) );
  ANDN U1577 ( .B(n1065), .A(n1066), .Z(n1063) );
  XNOR U1578 ( .A(b[266]), .B(n1064), .Z(n1065) );
  XNOR U1579 ( .A(b[266]), .B(n1066), .Z(c[266]) );
  XOR U1580 ( .A(n1067), .B(n1068), .Z(n1064) );
  ANDN U1581 ( .B(n1069), .A(n1070), .Z(n1067) );
  XNOR U1582 ( .A(b[265]), .B(n1068), .Z(n1069) );
  XNOR U1583 ( .A(b[265]), .B(n1070), .Z(c[265]) );
  XOR U1584 ( .A(n1071), .B(n1072), .Z(n1068) );
  ANDN U1585 ( .B(n1073), .A(n1074), .Z(n1071) );
  XNOR U1586 ( .A(b[264]), .B(n1072), .Z(n1073) );
  XNOR U1587 ( .A(b[264]), .B(n1074), .Z(c[264]) );
  XOR U1588 ( .A(n1075), .B(n1076), .Z(n1072) );
  ANDN U1589 ( .B(n1077), .A(n1078), .Z(n1075) );
  XNOR U1590 ( .A(b[263]), .B(n1076), .Z(n1077) );
  XNOR U1591 ( .A(b[263]), .B(n1078), .Z(c[263]) );
  XOR U1592 ( .A(n1079), .B(n1080), .Z(n1076) );
  ANDN U1593 ( .B(n1081), .A(n1082), .Z(n1079) );
  XNOR U1594 ( .A(b[262]), .B(n1080), .Z(n1081) );
  XNOR U1595 ( .A(b[262]), .B(n1082), .Z(c[262]) );
  XOR U1596 ( .A(n1083), .B(n1084), .Z(n1080) );
  ANDN U1597 ( .B(n1085), .A(n1086), .Z(n1083) );
  XNOR U1598 ( .A(b[261]), .B(n1084), .Z(n1085) );
  XNOR U1599 ( .A(b[261]), .B(n1086), .Z(c[261]) );
  XOR U1600 ( .A(n1087), .B(n1088), .Z(n1084) );
  ANDN U1601 ( .B(n1089), .A(n1090), .Z(n1087) );
  XNOR U1602 ( .A(b[260]), .B(n1088), .Z(n1089) );
  XNOR U1603 ( .A(b[260]), .B(n1090), .Z(c[260]) );
  XOR U1604 ( .A(n1091), .B(n1092), .Z(n1088) );
  ANDN U1605 ( .B(n1093), .A(n1094), .Z(n1091) );
  XNOR U1606 ( .A(b[259]), .B(n1092), .Z(n1093) );
  XNOR U1607 ( .A(b[25]), .B(n1095), .Z(c[25]) );
  XNOR U1608 ( .A(b[259]), .B(n1094), .Z(c[259]) );
  XOR U1609 ( .A(n1096), .B(n1097), .Z(n1092) );
  ANDN U1610 ( .B(n1098), .A(n1099), .Z(n1096) );
  XNOR U1611 ( .A(b[258]), .B(n1097), .Z(n1098) );
  XNOR U1612 ( .A(b[258]), .B(n1099), .Z(c[258]) );
  XOR U1613 ( .A(n1100), .B(n1101), .Z(n1097) );
  ANDN U1614 ( .B(n1102), .A(n1103), .Z(n1100) );
  XNOR U1615 ( .A(b[257]), .B(n1101), .Z(n1102) );
  XNOR U1616 ( .A(b[257]), .B(n1103), .Z(c[257]) );
  XOR U1617 ( .A(n1104), .B(n1105), .Z(n1101) );
  ANDN U1618 ( .B(n1106), .A(n1107), .Z(n1104) );
  XNOR U1619 ( .A(b[256]), .B(n1105), .Z(n1106) );
  XNOR U1620 ( .A(b[256]), .B(n1107), .Z(c[256]) );
  XOR U1621 ( .A(n1108), .B(n1109), .Z(n1105) );
  ANDN U1622 ( .B(n1110), .A(n1111), .Z(n1108) );
  XNOR U1623 ( .A(b[255]), .B(n1109), .Z(n1110) );
  XNOR U1624 ( .A(b[255]), .B(n1111), .Z(c[255]) );
  XOR U1625 ( .A(n1112), .B(n1113), .Z(n1109) );
  ANDN U1626 ( .B(n1114), .A(n1115), .Z(n1112) );
  XNOR U1627 ( .A(b[254]), .B(n1113), .Z(n1114) );
  XNOR U1628 ( .A(b[254]), .B(n1115), .Z(c[254]) );
  XOR U1629 ( .A(n1116), .B(n1117), .Z(n1113) );
  ANDN U1630 ( .B(n1118), .A(n1119), .Z(n1116) );
  XNOR U1631 ( .A(b[253]), .B(n1117), .Z(n1118) );
  XNOR U1632 ( .A(b[253]), .B(n1119), .Z(c[253]) );
  XOR U1633 ( .A(n1120), .B(n1121), .Z(n1117) );
  ANDN U1634 ( .B(n1122), .A(n1123), .Z(n1120) );
  XNOR U1635 ( .A(b[252]), .B(n1121), .Z(n1122) );
  XNOR U1636 ( .A(b[252]), .B(n1123), .Z(c[252]) );
  XOR U1637 ( .A(n1124), .B(n1125), .Z(n1121) );
  ANDN U1638 ( .B(n1126), .A(n1127), .Z(n1124) );
  XNOR U1639 ( .A(b[251]), .B(n1125), .Z(n1126) );
  XNOR U1640 ( .A(b[251]), .B(n1127), .Z(c[251]) );
  XOR U1641 ( .A(n1128), .B(n1129), .Z(n1125) );
  ANDN U1642 ( .B(n1130), .A(n1131), .Z(n1128) );
  XNOR U1643 ( .A(b[250]), .B(n1129), .Z(n1130) );
  XNOR U1644 ( .A(b[250]), .B(n1131), .Z(c[250]) );
  XOR U1645 ( .A(n1132), .B(n1133), .Z(n1129) );
  ANDN U1646 ( .B(n1134), .A(n1135), .Z(n1132) );
  XNOR U1647 ( .A(b[249]), .B(n1133), .Z(n1134) );
  XNOR U1648 ( .A(b[24]), .B(n1136), .Z(c[24]) );
  XNOR U1649 ( .A(b[249]), .B(n1135), .Z(c[249]) );
  XOR U1650 ( .A(n1137), .B(n1138), .Z(n1133) );
  ANDN U1651 ( .B(n1139), .A(n1140), .Z(n1137) );
  XNOR U1652 ( .A(b[248]), .B(n1138), .Z(n1139) );
  XNOR U1653 ( .A(b[248]), .B(n1140), .Z(c[248]) );
  XOR U1654 ( .A(n1141), .B(n1142), .Z(n1138) );
  ANDN U1655 ( .B(n1143), .A(n1144), .Z(n1141) );
  XNOR U1656 ( .A(b[247]), .B(n1142), .Z(n1143) );
  XNOR U1657 ( .A(b[247]), .B(n1144), .Z(c[247]) );
  XOR U1658 ( .A(n1145), .B(n1146), .Z(n1142) );
  ANDN U1659 ( .B(n1147), .A(n1148), .Z(n1145) );
  XNOR U1660 ( .A(b[246]), .B(n1146), .Z(n1147) );
  XNOR U1661 ( .A(b[246]), .B(n1148), .Z(c[246]) );
  XOR U1662 ( .A(n1149), .B(n1150), .Z(n1146) );
  ANDN U1663 ( .B(n1151), .A(n1152), .Z(n1149) );
  XNOR U1664 ( .A(b[245]), .B(n1150), .Z(n1151) );
  XNOR U1665 ( .A(b[245]), .B(n1152), .Z(c[245]) );
  XOR U1666 ( .A(n1153), .B(n1154), .Z(n1150) );
  ANDN U1667 ( .B(n1155), .A(n1156), .Z(n1153) );
  XNOR U1668 ( .A(b[244]), .B(n1154), .Z(n1155) );
  XNOR U1669 ( .A(b[244]), .B(n1156), .Z(c[244]) );
  XOR U1670 ( .A(n1157), .B(n1158), .Z(n1154) );
  ANDN U1671 ( .B(n1159), .A(n1160), .Z(n1157) );
  XNOR U1672 ( .A(b[243]), .B(n1158), .Z(n1159) );
  XNOR U1673 ( .A(b[243]), .B(n1160), .Z(c[243]) );
  XOR U1674 ( .A(n1161), .B(n1162), .Z(n1158) );
  ANDN U1675 ( .B(n1163), .A(n1164), .Z(n1161) );
  XNOR U1676 ( .A(b[242]), .B(n1162), .Z(n1163) );
  XNOR U1677 ( .A(b[242]), .B(n1164), .Z(c[242]) );
  XOR U1678 ( .A(n1165), .B(n1166), .Z(n1162) );
  ANDN U1679 ( .B(n1167), .A(n1168), .Z(n1165) );
  XNOR U1680 ( .A(b[241]), .B(n1166), .Z(n1167) );
  XNOR U1681 ( .A(b[241]), .B(n1168), .Z(c[241]) );
  XOR U1682 ( .A(n1169), .B(n1170), .Z(n1166) );
  ANDN U1683 ( .B(n1171), .A(n1172), .Z(n1169) );
  XNOR U1684 ( .A(b[240]), .B(n1170), .Z(n1171) );
  XNOR U1685 ( .A(b[240]), .B(n1172), .Z(c[240]) );
  XOR U1686 ( .A(n1173), .B(n1174), .Z(n1170) );
  ANDN U1687 ( .B(n1175), .A(n1176), .Z(n1173) );
  XNOR U1688 ( .A(b[239]), .B(n1174), .Z(n1175) );
  XNOR U1689 ( .A(b[23]), .B(n1177), .Z(c[23]) );
  XNOR U1690 ( .A(b[239]), .B(n1176), .Z(c[239]) );
  XOR U1691 ( .A(n1178), .B(n1179), .Z(n1174) );
  ANDN U1692 ( .B(n1180), .A(n1181), .Z(n1178) );
  XNOR U1693 ( .A(b[238]), .B(n1179), .Z(n1180) );
  XNOR U1694 ( .A(b[238]), .B(n1181), .Z(c[238]) );
  XOR U1695 ( .A(n1182), .B(n1183), .Z(n1179) );
  ANDN U1696 ( .B(n1184), .A(n1185), .Z(n1182) );
  XNOR U1697 ( .A(b[237]), .B(n1183), .Z(n1184) );
  XNOR U1698 ( .A(b[237]), .B(n1185), .Z(c[237]) );
  XOR U1699 ( .A(n1186), .B(n1187), .Z(n1183) );
  ANDN U1700 ( .B(n1188), .A(n1189), .Z(n1186) );
  XNOR U1701 ( .A(b[236]), .B(n1187), .Z(n1188) );
  XNOR U1702 ( .A(b[236]), .B(n1189), .Z(c[236]) );
  XOR U1703 ( .A(n1190), .B(n1191), .Z(n1187) );
  ANDN U1704 ( .B(n1192), .A(n1193), .Z(n1190) );
  XNOR U1705 ( .A(b[235]), .B(n1191), .Z(n1192) );
  XNOR U1706 ( .A(b[235]), .B(n1193), .Z(c[235]) );
  XOR U1707 ( .A(n1194), .B(n1195), .Z(n1191) );
  ANDN U1708 ( .B(n1196), .A(n1197), .Z(n1194) );
  XNOR U1709 ( .A(b[234]), .B(n1195), .Z(n1196) );
  XNOR U1710 ( .A(b[234]), .B(n1197), .Z(c[234]) );
  XOR U1711 ( .A(n1198), .B(n1199), .Z(n1195) );
  ANDN U1712 ( .B(n1200), .A(n1201), .Z(n1198) );
  XNOR U1713 ( .A(b[233]), .B(n1199), .Z(n1200) );
  XNOR U1714 ( .A(b[233]), .B(n1201), .Z(c[233]) );
  XOR U1715 ( .A(n1202), .B(n1203), .Z(n1199) );
  ANDN U1716 ( .B(n1204), .A(n1205), .Z(n1202) );
  XNOR U1717 ( .A(b[232]), .B(n1203), .Z(n1204) );
  XNOR U1718 ( .A(b[232]), .B(n1205), .Z(c[232]) );
  XOR U1719 ( .A(n1206), .B(n1207), .Z(n1203) );
  ANDN U1720 ( .B(n1208), .A(n1209), .Z(n1206) );
  XNOR U1721 ( .A(b[231]), .B(n1207), .Z(n1208) );
  XNOR U1722 ( .A(b[231]), .B(n1209), .Z(c[231]) );
  XOR U1723 ( .A(n1210), .B(n1211), .Z(n1207) );
  ANDN U1724 ( .B(n1212), .A(n1213), .Z(n1210) );
  XNOR U1725 ( .A(b[230]), .B(n1211), .Z(n1212) );
  XNOR U1726 ( .A(b[230]), .B(n1213), .Z(c[230]) );
  XOR U1727 ( .A(n1214), .B(n1215), .Z(n1211) );
  ANDN U1728 ( .B(n1216), .A(n1217), .Z(n1214) );
  XNOR U1729 ( .A(b[229]), .B(n1215), .Z(n1216) );
  XNOR U1730 ( .A(b[22]), .B(n1218), .Z(c[22]) );
  XNOR U1731 ( .A(b[229]), .B(n1217), .Z(c[229]) );
  XOR U1732 ( .A(n1219), .B(n1220), .Z(n1215) );
  ANDN U1733 ( .B(n1221), .A(n1222), .Z(n1219) );
  XNOR U1734 ( .A(b[228]), .B(n1220), .Z(n1221) );
  XNOR U1735 ( .A(b[228]), .B(n1222), .Z(c[228]) );
  XOR U1736 ( .A(n1223), .B(n1224), .Z(n1220) );
  ANDN U1737 ( .B(n1225), .A(n1226), .Z(n1223) );
  XNOR U1738 ( .A(b[227]), .B(n1224), .Z(n1225) );
  XNOR U1739 ( .A(b[227]), .B(n1226), .Z(c[227]) );
  XOR U1740 ( .A(n1227), .B(n1228), .Z(n1224) );
  ANDN U1741 ( .B(n1229), .A(n1230), .Z(n1227) );
  XNOR U1742 ( .A(b[226]), .B(n1228), .Z(n1229) );
  XNOR U1743 ( .A(b[226]), .B(n1230), .Z(c[226]) );
  XOR U1744 ( .A(n1231), .B(n1232), .Z(n1228) );
  ANDN U1745 ( .B(n1233), .A(n1234), .Z(n1231) );
  XNOR U1746 ( .A(b[225]), .B(n1232), .Z(n1233) );
  XNOR U1747 ( .A(b[225]), .B(n1234), .Z(c[225]) );
  XOR U1748 ( .A(n1235), .B(n1236), .Z(n1232) );
  ANDN U1749 ( .B(n1237), .A(n1238), .Z(n1235) );
  XNOR U1750 ( .A(b[224]), .B(n1236), .Z(n1237) );
  XNOR U1751 ( .A(b[224]), .B(n1238), .Z(c[224]) );
  XOR U1752 ( .A(n1239), .B(n1240), .Z(n1236) );
  ANDN U1753 ( .B(n1241), .A(n1242), .Z(n1239) );
  XNOR U1754 ( .A(b[223]), .B(n1240), .Z(n1241) );
  XNOR U1755 ( .A(b[223]), .B(n1242), .Z(c[223]) );
  XOR U1756 ( .A(n1243), .B(n1244), .Z(n1240) );
  ANDN U1757 ( .B(n1245), .A(n1246), .Z(n1243) );
  XNOR U1758 ( .A(b[222]), .B(n1244), .Z(n1245) );
  XNOR U1759 ( .A(b[222]), .B(n1246), .Z(c[222]) );
  XOR U1760 ( .A(n1247), .B(n1248), .Z(n1244) );
  ANDN U1761 ( .B(n1249), .A(n1250), .Z(n1247) );
  XNOR U1762 ( .A(b[221]), .B(n1248), .Z(n1249) );
  XNOR U1763 ( .A(b[221]), .B(n1250), .Z(c[221]) );
  XOR U1764 ( .A(n1251), .B(n1252), .Z(n1248) );
  ANDN U1765 ( .B(n1253), .A(n1254), .Z(n1251) );
  XNOR U1766 ( .A(b[220]), .B(n1252), .Z(n1253) );
  XNOR U1767 ( .A(b[220]), .B(n1254), .Z(c[220]) );
  XOR U1768 ( .A(n1255), .B(n1256), .Z(n1252) );
  ANDN U1769 ( .B(n1257), .A(n1258), .Z(n1255) );
  XNOR U1770 ( .A(b[219]), .B(n1256), .Z(n1257) );
  XNOR U1771 ( .A(b[21]), .B(n1259), .Z(c[21]) );
  XNOR U1772 ( .A(b[219]), .B(n1258), .Z(c[219]) );
  XOR U1773 ( .A(n1260), .B(n1261), .Z(n1256) );
  ANDN U1774 ( .B(n1262), .A(n1263), .Z(n1260) );
  XNOR U1775 ( .A(b[218]), .B(n1261), .Z(n1262) );
  XNOR U1776 ( .A(b[218]), .B(n1263), .Z(c[218]) );
  XOR U1777 ( .A(n1264), .B(n1265), .Z(n1261) );
  ANDN U1778 ( .B(n1266), .A(n1267), .Z(n1264) );
  XNOR U1779 ( .A(b[217]), .B(n1265), .Z(n1266) );
  XNOR U1780 ( .A(b[217]), .B(n1267), .Z(c[217]) );
  XOR U1781 ( .A(n1268), .B(n1269), .Z(n1265) );
  ANDN U1782 ( .B(n1270), .A(n1271), .Z(n1268) );
  XNOR U1783 ( .A(b[216]), .B(n1269), .Z(n1270) );
  XNOR U1784 ( .A(b[216]), .B(n1271), .Z(c[216]) );
  XOR U1785 ( .A(n1272), .B(n1273), .Z(n1269) );
  ANDN U1786 ( .B(n1274), .A(n1275), .Z(n1272) );
  XNOR U1787 ( .A(b[215]), .B(n1273), .Z(n1274) );
  XNOR U1788 ( .A(b[215]), .B(n1275), .Z(c[215]) );
  XOR U1789 ( .A(n1276), .B(n1277), .Z(n1273) );
  ANDN U1790 ( .B(n1278), .A(n1279), .Z(n1276) );
  XNOR U1791 ( .A(b[214]), .B(n1277), .Z(n1278) );
  XNOR U1792 ( .A(b[214]), .B(n1279), .Z(c[214]) );
  XOR U1793 ( .A(n1280), .B(n1281), .Z(n1277) );
  ANDN U1794 ( .B(n1282), .A(n1283), .Z(n1280) );
  XNOR U1795 ( .A(b[213]), .B(n1281), .Z(n1282) );
  XNOR U1796 ( .A(b[213]), .B(n1283), .Z(c[213]) );
  XOR U1797 ( .A(n1284), .B(n1285), .Z(n1281) );
  ANDN U1798 ( .B(n1286), .A(n1287), .Z(n1284) );
  XNOR U1799 ( .A(b[212]), .B(n1285), .Z(n1286) );
  XNOR U1800 ( .A(b[212]), .B(n1287), .Z(c[212]) );
  XOR U1801 ( .A(n1288), .B(n1289), .Z(n1285) );
  ANDN U1802 ( .B(n1290), .A(n1291), .Z(n1288) );
  XNOR U1803 ( .A(b[211]), .B(n1289), .Z(n1290) );
  XNOR U1804 ( .A(b[211]), .B(n1291), .Z(c[211]) );
  XOR U1805 ( .A(n1292), .B(n1293), .Z(n1289) );
  ANDN U1806 ( .B(n1294), .A(n1295), .Z(n1292) );
  XNOR U1807 ( .A(b[210]), .B(n1293), .Z(n1294) );
  XNOR U1808 ( .A(b[210]), .B(n1295), .Z(c[210]) );
  XOR U1809 ( .A(n1296), .B(n1297), .Z(n1293) );
  ANDN U1810 ( .B(n1298), .A(n1299), .Z(n1296) );
  XNOR U1811 ( .A(b[209]), .B(n1297), .Z(n1298) );
  XNOR U1812 ( .A(b[20]), .B(n1300), .Z(c[20]) );
  XNOR U1813 ( .A(b[209]), .B(n1299), .Z(c[209]) );
  XOR U1814 ( .A(n1301), .B(n1302), .Z(n1297) );
  ANDN U1815 ( .B(n1303), .A(n1304), .Z(n1301) );
  XNOR U1816 ( .A(b[208]), .B(n1302), .Z(n1303) );
  XNOR U1817 ( .A(b[208]), .B(n1304), .Z(c[208]) );
  XOR U1818 ( .A(n1305), .B(n1306), .Z(n1302) );
  ANDN U1819 ( .B(n1307), .A(n1308), .Z(n1305) );
  XNOR U1820 ( .A(b[207]), .B(n1306), .Z(n1307) );
  XNOR U1821 ( .A(b[207]), .B(n1308), .Z(c[207]) );
  XOR U1822 ( .A(n1309), .B(n1310), .Z(n1306) );
  ANDN U1823 ( .B(n1311), .A(n1312), .Z(n1309) );
  XNOR U1824 ( .A(b[206]), .B(n1310), .Z(n1311) );
  XNOR U1825 ( .A(b[206]), .B(n1312), .Z(c[206]) );
  XOR U1826 ( .A(n1313), .B(n1314), .Z(n1310) );
  ANDN U1827 ( .B(n1315), .A(n1316), .Z(n1313) );
  XNOR U1828 ( .A(b[205]), .B(n1314), .Z(n1315) );
  XNOR U1829 ( .A(b[205]), .B(n1316), .Z(c[205]) );
  XOR U1830 ( .A(n1317), .B(n1318), .Z(n1314) );
  ANDN U1831 ( .B(n1319), .A(n1320), .Z(n1317) );
  XNOR U1832 ( .A(b[204]), .B(n1318), .Z(n1319) );
  XNOR U1833 ( .A(b[204]), .B(n1320), .Z(c[204]) );
  XOR U1834 ( .A(n1321), .B(n1322), .Z(n1318) );
  ANDN U1835 ( .B(n1323), .A(n1324), .Z(n1321) );
  XNOR U1836 ( .A(b[203]), .B(n1322), .Z(n1323) );
  XNOR U1837 ( .A(b[203]), .B(n1324), .Z(c[203]) );
  XOR U1838 ( .A(n1325), .B(n1326), .Z(n1322) );
  ANDN U1839 ( .B(n1327), .A(n1328), .Z(n1325) );
  XNOR U1840 ( .A(b[202]), .B(n1326), .Z(n1327) );
  XNOR U1841 ( .A(b[202]), .B(n1328), .Z(c[202]) );
  XOR U1842 ( .A(n1329), .B(n1330), .Z(n1326) );
  ANDN U1843 ( .B(n1331), .A(n1332), .Z(n1329) );
  XNOR U1844 ( .A(b[201]), .B(n1330), .Z(n1331) );
  XNOR U1845 ( .A(b[201]), .B(n1332), .Z(c[201]) );
  XOR U1846 ( .A(n1333), .B(n1334), .Z(n1330) );
  ANDN U1847 ( .B(n1335), .A(n1336), .Z(n1333) );
  XNOR U1848 ( .A(b[200]), .B(n1334), .Z(n1335) );
  XNOR U1849 ( .A(b[200]), .B(n1336), .Z(c[200]) );
  XOR U1850 ( .A(n1337), .B(n1338), .Z(n1334) );
  ANDN U1851 ( .B(n1339), .A(n1340), .Z(n1337) );
  XNOR U1852 ( .A(b[199]), .B(n1338), .Z(n1339) );
  XNOR U1853 ( .A(b[1]), .B(n1341), .Z(c[1]) );
  XNOR U1854 ( .A(b[19]), .B(n1342), .Z(c[19]) );
  XNOR U1855 ( .A(b[199]), .B(n1340), .Z(c[199]) );
  XOR U1856 ( .A(n1343), .B(n1344), .Z(n1338) );
  ANDN U1857 ( .B(n1345), .A(n1346), .Z(n1343) );
  XNOR U1858 ( .A(b[198]), .B(n1344), .Z(n1345) );
  XNOR U1859 ( .A(b[198]), .B(n1346), .Z(c[198]) );
  XOR U1860 ( .A(n1347), .B(n1348), .Z(n1344) );
  ANDN U1861 ( .B(n1349), .A(n1350), .Z(n1347) );
  XNOR U1862 ( .A(b[197]), .B(n1348), .Z(n1349) );
  XNOR U1863 ( .A(b[197]), .B(n1350), .Z(c[197]) );
  XOR U1864 ( .A(n1351), .B(n1352), .Z(n1348) );
  ANDN U1865 ( .B(n1353), .A(n1354), .Z(n1351) );
  XNOR U1866 ( .A(b[196]), .B(n1352), .Z(n1353) );
  XNOR U1867 ( .A(b[196]), .B(n1354), .Z(c[196]) );
  XOR U1868 ( .A(n1355), .B(n1356), .Z(n1352) );
  ANDN U1869 ( .B(n1357), .A(n1358), .Z(n1355) );
  XNOR U1870 ( .A(b[195]), .B(n1356), .Z(n1357) );
  XNOR U1871 ( .A(b[195]), .B(n1358), .Z(c[195]) );
  XOR U1872 ( .A(n1359), .B(n1360), .Z(n1356) );
  ANDN U1873 ( .B(n1361), .A(n1362), .Z(n1359) );
  XNOR U1874 ( .A(b[194]), .B(n1360), .Z(n1361) );
  XNOR U1875 ( .A(b[194]), .B(n1362), .Z(c[194]) );
  XOR U1876 ( .A(n1363), .B(n1364), .Z(n1360) );
  ANDN U1877 ( .B(n1365), .A(n1366), .Z(n1363) );
  XNOR U1878 ( .A(b[193]), .B(n1364), .Z(n1365) );
  XNOR U1879 ( .A(b[193]), .B(n1366), .Z(c[193]) );
  XOR U1880 ( .A(n1367), .B(n1368), .Z(n1364) );
  ANDN U1881 ( .B(n1369), .A(n1370), .Z(n1367) );
  XNOR U1882 ( .A(b[192]), .B(n1368), .Z(n1369) );
  XNOR U1883 ( .A(b[192]), .B(n1370), .Z(c[192]) );
  XOR U1884 ( .A(n1371), .B(n1372), .Z(n1368) );
  ANDN U1885 ( .B(n1373), .A(n1374), .Z(n1371) );
  XNOR U1886 ( .A(b[191]), .B(n1372), .Z(n1373) );
  XNOR U1887 ( .A(b[191]), .B(n1374), .Z(c[191]) );
  XOR U1888 ( .A(n1375), .B(n1376), .Z(n1372) );
  ANDN U1889 ( .B(n1377), .A(n1378), .Z(n1375) );
  XNOR U1890 ( .A(b[190]), .B(n1376), .Z(n1377) );
  XNOR U1891 ( .A(b[190]), .B(n1378), .Z(c[190]) );
  XOR U1892 ( .A(n1379), .B(n1380), .Z(n1376) );
  ANDN U1893 ( .B(n1381), .A(n1382), .Z(n1379) );
  XNOR U1894 ( .A(b[189]), .B(n1380), .Z(n1381) );
  XNOR U1895 ( .A(b[18]), .B(n1383), .Z(c[18]) );
  XNOR U1896 ( .A(b[189]), .B(n1382), .Z(c[189]) );
  XOR U1897 ( .A(n1384), .B(n1385), .Z(n1380) );
  ANDN U1898 ( .B(n1386), .A(n1387), .Z(n1384) );
  XNOR U1899 ( .A(b[188]), .B(n1385), .Z(n1386) );
  XNOR U1900 ( .A(b[188]), .B(n1387), .Z(c[188]) );
  XOR U1901 ( .A(n1388), .B(n1389), .Z(n1385) );
  ANDN U1902 ( .B(n1390), .A(n1391), .Z(n1388) );
  XNOR U1903 ( .A(b[187]), .B(n1389), .Z(n1390) );
  XNOR U1904 ( .A(b[187]), .B(n1391), .Z(c[187]) );
  XOR U1905 ( .A(n1392), .B(n1393), .Z(n1389) );
  ANDN U1906 ( .B(n1394), .A(n1395), .Z(n1392) );
  XNOR U1907 ( .A(b[186]), .B(n1393), .Z(n1394) );
  XNOR U1908 ( .A(b[186]), .B(n1395), .Z(c[186]) );
  XOR U1909 ( .A(n1396), .B(n1397), .Z(n1393) );
  ANDN U1910 ( .B(n1398), .A(n1399), .Z(n1396) );
  XNOR U1911 ( .A(b[185]), .B(n1397), .Z(n1398) );
  XNOR U1912 ( .A(b[185]), .B(n1399), .Z(c[185]) );
  XOR U1913 ( .A(n1400), .B(n1401), .Z(n1397) );
  ANDN U1914 ( .B(n1402), .A(n1403), .Z(n1400) );
  XNOR U1915 ( .A(b[184]), .B(n1401), .Z(n1402) );
  XNOR U1916 ( .A(b[184]), .B(n1403), .Z(c[184]) );
  XOR U1917 ( .A(n1404), .B(n1405), .Z(n1401) );
  ANDN U1918 ( .B(n1406), .A(n1407), .Z(n1404) );
  XNOR U1919 ( .A(b[183]), .B(n1405), .Z(n1406) );
  XNOR U1920 ( .A(b[183]), .B(n1407), .Z(c[183]) );
  XOR U1921 ( .A(n1408), .B(n1409), .Z(n1405) );
  ANDN U1922 ( .B(n1410), .A(n1411), .Z(n1408) );
  XNOR U1923 ( .A(b[182]), .B(n1409), .Z(n1410) );
  XNOR U1924 ( .A(b[182]), .B(n1411), .Z(c[182]) );
  XOR U1925 ( .A(n1412), .B(n1413), .Z(n1409) );
  ANDN U1926 ( .B(n1414), .A(n1415), .Z(n1412) );
  XNOR U1927 ( .A(b[181]), .B(n1413), .Z(n1414) );
  XNOR U1928 ( .A(b[181]), .B(n1415), .Z(c[181]) );
  XOR U1929 ( .A(n1416), .B(n1417), .Z(n1413) );
  ANDN U1930 ( .B(n1418), .A(n1419), .Z(n1416) );
  XNOR U1931 ( .A(b[180]), .B(n1417), .Z(n1418) );
  XNOR U1932 ( .A(b[180]), .B(n1419), .Z(c[180]) );
  XOR U1933 ( .A(n1420), .B(n1421), .Z(n1417) );
  ANDN U1934 ( .B(n1422), .A(n1423), .Z(n1420) );
  XNOR U1935 ( .A(b[179]), .B(n1421), .Z(n1422) );
  XNOR U1936 ( .A(b[17]), .B(n1424), .Z(c[17]) );
  XNOR U1937 ( .A(b[179]), .B(n1423), .Z(c[179]) );
  XOR U1938 ( .A(n1425), .B(n1426), .Z(n1421) );
  ANDN U1939 ( .B(n1427), .A(n1428), .Z(n1425) );
  XNOR U1940 ( .A(b[178]), .B(n1426), .Z(n1427) );
  XNOR U1941 ( .A(b[178]), .B(n1428), .Z(c[178]) );
  XOR U1942 ( .A(n1429), .B(n1430), .Z(n1426) );
  ANDN U1943 ( .B(n1431), .A(n1432), .Z(n1429) );
  XNOR U1944 ( .A(b[177]), .B(n1430), .Z(n1431) );
  XNOR U1945 ( .A(b[177]), .B(n1432), .Z(c[177]) );
  XOR U1946 ( .A(n1433), .B(n1434), .Z(n1430) );
  ANDN U1947 ( .B(n1435), .A(n1436), .Z(n1433) );
  XNOR U1948 ( .A(b[176]), .B(n1434), .Z(n1435) );
  XNOR U1949 ( .A(b[176]), .B(n1436), .Z(c[176]) );
  XOR U1950 ( .A(n1437), .B(n1438), .Z(n1434) );
  ANDN U1951 ( .B(n1439), .A(n1440), .Z(n1437) );
  XNOR U1952 ( .A(b[175]), .B(n1438), .Z(n1439) );
  XNOR U1953 ( .A(b[175]), .B(n1440), .Z(c[175]) );
  XOR U1954 ( .A(n1441), .B(n1442), .Z(n1438) );
  ANDN U1955 ( .B(n1443), .A(n1444), .Z(n1441) );
  XNOR U1956 ( .A(b[174]), .B(n1442), .Z(n1443) );
  XNOR U1957 ( .A(b[174]), .B(n1444), .Z(c[174]) );
  XOR U1958 ( .A(n1445), .B(n1446), .Z(n1442) );
  ANDN U1959 ( .B(n1447), .A(n1448), .Z(n1445) );
  XNOR U1960 ( .A(b[173]), .B(n1446), .Z(n1447) );
  XNOR U1961 ( .A(b[173]), .B(n1448), .Z(c[173]) );
  XOR U1962 ( .A(n1449), .B(n1450), .Z(n1446) );
  ANDN U1963 ( .B(n1451), .A(n1452), .Z(n1449) );
  XNOR U1964 ( .A(b[172]), .B(n1450), .Z(n1451) );
  XNOR U1965 ( .A(b[172]), .B(n1452), .Z(c[172]) );
  XOR U1966 ( .A(n1453), .B(n1454), .Z(n1450) );
  ANDN U1967 ( .B(n1455), .A(n1456), .Z(n1453) );
  XNOR U1968 ( .A(b[171]), .B(n1454), .Z(n1455) );
  XNOR U1969 ( .A(b[171]), .B(n1456), .Z(c[171]) );
  XOR U1970 ( .A(n1457), .B(n1458), .Z(n1454) );
  ANDN U1971 ( .B(n1459), .A(n1460), .Z(n1457) );
  XNOR U1972 ( .A(b[170]), .B(n1458), .Z(n1459) );
  XNOR U1973 ( .A(b[170]), .B(n1460), .Z(c[170]) );
  XOR U1974 ( .A(n1461), .B(n1462), .Z(n1458) );
  ANDN U1975 ( .B(n1463), .A(n1464), .Z(n1461) );
  XNOR U1976 ( .A(b[169]), .B(n1462), .Z(n1463) );
  XNOR U1977 ( .A(b[16]), .B(n1465), .Z(c[16]) );
  XNOR U1978 ( .A(b[169]), .B(n1464), .Z(c[169]) );
  XOR U1979 ( .A(n1466), .B(n1467), .Z(n1462) );
  ANDN U1980 ( .B(n1468), .A(n1469), .Z(n1466) );
  XNOR U1981 ( .A(b[168]), .B(n1467), .Z(n1468) );
  XNOR U1982 ( .A(b[168]), .B(n1469), .Z(c[168]) );
  XOR U1983 ( .A(n1470), .B(n1471), .Z(n1467) );
  ANDN U1984 ( .B(n1472), .A(n1473), .Z(n1470) );
  XNOR U1985 ( .A(b[167]), .B(n1471), .Z(n1472) );
  XNOR U1986 ( .A(b[167]), .B(n1473), .Z(c[167]) );
  XOR U1987 ( .A(n1474), .B(n1475), .Z(n1471) );
  ANDN U1988 ( .B(n1476), .A(n1477), .Z(n1474) );
  XNOR U1989 ( .A(b[166]), .B(n1475), .Z(n1476) );
  XNOR U1990 ( .A(b[166]), .B(n1477), .Z(c[166]) );
  XOR U1991 ( .A(n1478), .B(n1479), .Z(n1475) );
  ANDN U1992 ( .B(n1480), .A(n1481), .Z(n1478) );
  XNOR U1993 ( .A(b[165]), .B(n1479), .Z(n1480) );
  XNOR U1994 ( .A(b[165]), .B(n1481), .Z(c[165]) );
  XOR U1995 ( .A(n1482), .B(n1483), .Z(n1479) );
  ANDN U1996 ( .B(n1484), .A(n1485), .Z(n1482) );
  XNOR U1997 ( .A(b[164]), .B(n1483), .Z(n1484) );
  XNOR U1998 ( .A(b[164]), .B(n1485), .Z(c[164]) );
  XOR U1999 ( .A(n1486), .B(n1487), .Z(n1483) );
  ANDN U2000 ( .B(n1488), .A(n1489), .Z(n1486) );
  XNOR U2001 ( .A(b[163]), .B(n1487), .Z(n1488) );
  XNOR U2002 ( .A(b[163]), .B(n1489), .Z(c[163]) );
  XOR U2003 ( .A(n1490), .B(n1491), .Z(n1487) );
  ANDN U2004 ( .B(n1492), .A(n1493), .Z(n1490) );
  XNOR U2005 ( .A(b[162]), .B(n1491), .Z(n1492) );
  XNOR U2006 ( .A(b[162]), .B(n1493), .Z(c[162]) );
  XOR U2007 ( .A(n1494), .B(n1495), .Z(n1491) );
  ANDN U2008 ( .B(n1496), .A(n1497), .Z(n1494) );
  XNOR U2009 ( .A(b[161]), .B(n1495), .Z(n1496) );
  XNOR U2010 ( .A(b[161]), .B(n1497), .Z(c[161]) );
  XOR U2011 ( .A(n1498), .B(n1499), .Z(n1495) );
  ANDN U2012 ( .B(n1500), .A(n1501), .Z(n1498) );
  XNOR U2013 ( .A(b[160]), .B(n1499), .Z(n1500) );
  XNOR U2014 ( .A(b[160]), .B(n1501), .Z(c[160]) );
  XOR U2015 ( .A(n1502), .B(n1503), .Z(n1499) );
  ANDN U2016 ( .B(n1504), .A(n1505), .Z(n1502) );
  XNOR U2017 ( .A(b[159]), .B(n1503), .Z(n1504) );
  XNOR U2018 ( .A(b[15]), .B(n1506), .Z(c[15]) );
  XNOR U2019 ( .A(b[159]), .B(n1505), .Z(c[159]) );
  XOR U2020 ( .A(n1507), .B(n1508), .Z(n1503) );
  ANDN U2021 ( .B(n1509), .A(n1510), .Z(n1507) );
  XNOR U2022 ( .A(b[158]), .B(n1508), .Z(n1509) );
  XNOR U2023 ( .A(b[158]), .B(n1510), .Z(c[158]) );
  XOR U2024 ( .A(n1511), .B(n1512), .Z(n1508) );
  ANDN U2025 ( .B(n1513), .A(n1514), .Z(n1511) );
  XNOR U2026 ( .A(b[157]), .B(n1512), .Z(n1513) );
  XNOR U2027 ( .A(b[157]), .B(n1514), .Z(c[157]) );
  XOR U2028 ( .A(n1515), .B(n1516), .Z(n1512) );
  ANDN U2029 ( .B(n1517), .A(n1518), .Z(n1515) );
  XNOR U2030 ( .A(b[156]), .B(n1516), .Z(n1517) );
  XNOR U2031 ( .A(b[156]), .B(n1518), .Z(c[156]) );
  XOR U2032 ( .A(n1519), .B(n1520), .Z(n1516) );
  ANDN U2033 ( .B(n1521), .A(n1522), .Z(n1519) );
  XNOR U2034 ( .A(b[155]), .B(n1520), .Z(n1521) );
  XNOR U2035 ( .A(b[155]), .B(n1522), .Z(c[155]) );
  XOR U2036 ( .A(n1523), .B(n1524), .Z(n1520) );
  ANDN U2037 ( .B(n1525), .A(n1526), .Z(n1523) );
  XNOR U2038 ( .A(b[154]), .B(n1524), .Z(n1525) );
  XNOR U2039 ( .A(b[154]), .B(n1526), .Z(c[154]) );
  XOR U2040 ( .A(n1527), .B(n1528), .Z(n1524) );
  ANDN U2041 ( .B(n1529), .A(n1530), .Z(n1527) );
  XNOR U2042 ( .A(b[153]), .B(n1528), .Z(n1529) );
  XNOR U2043 ( .A(b[153]), .B(n1530), .Z(c[153]) );
  XOR U2044 ( .A(n1531), .B(n1532), .Z(n1528) );
  ANDN U2045 ( .B(n1533), .A(n1534), .Z(n1531) );
  XNOR U2046 ( .A(b[152]), .B(n1532), .Z(n1533) );
  XNOR U2047 ( .A(b[152]), .B(n1534), .Z(c[152]) );
  XOR U2048 ( .A(n1535), .B(n1536), .Z(n1532) );
  ANDN U2049 ( .B(n1537), .A(n1538), .Z(n1535) );
  XNOR U2050 ( .A(b[151]), .B(n1536), .Z(n1537) );
  XNOR U2051 ( .A(b[151]), .B(n1538), .Z(c[151]) );
  XOR U2052 ( .A(n1539), .B(n1540), .Z(n1536) );
  ANDN U2053 ( .B(n1541), .A(n1542), .Z(n1539) );
  XNOR U2054 ( .A(b[150]), .B(n1540), .Z(n1541) );
  XNOR U2055 ( .A(b[150]), .B(n1542), .Z(c[150]) );
  XOR U2056 ( .A(n1543), .B(n1544), .Z(n1540) );
  ANDN U2057 ( .B(n1545), .A(n1546), .Z(n1543) );
  XNOR U2058 ( .A(b[149]), .B(n1544), .Z(n1545) );
  XNOR U2059 ( .A(b[14]), .B(n1547), .Z(c[14]) );
  XNOR U2060 ( .A(b[149]), .B(n1546), .Z(c[149]) );
  XOR U2061 ( .A(n1548), .B(n1549), .Z(n1544) );
  ANDN U2062 ( .B(n1550), .A(n1551), .Z(n1548) );
  XNOR U2063 ( .A(b[148]), .B(n1549), .Z(n1550) );
  XNOR U2064 ( .A(b[148]), .B(n1551), .Z(c[148]) );
  XOR U2065 ( .A(n1552), .B(n1553), .Z(n1549) );
  ANDN U2066 ( .B(n1554), .A(n1555), .Z(n1552) );
  XNOR U2067 ( .A(b[147]), .B(n1553), .Z(n1554) );
  XNOR U2068 ( .A(b[147]), .B(n1555), .Z(c[147]) );
  XOR U2069 ( .A(n1556), .B(n1557), .Z(n1553) );
  ANDN U2070 ( .B(n1558), .A(n1559), .Z(n1556) );
  XNOR U2071 ( .A(b[146]), .B(n1557), .Z(n1558) );
  XNOR U2072 ( .A(b[146]), .B(n1559), .Z(c[146]) );
  XOR U2073 ( .A(n1560), .B(n1561), .Z(n1557) );
  ANDN U2074 ( .B(n1562), .A(n1563), .Z(n1560) );
  XNOR U2075 ( .A(b[145]), .B(n1561), .Z(n1562) );
  XNOR U2076 ( .A(b[145]), .B(n1563), .Z(c[145]) );
  XOR U2077 ( .A(n1564), .B(n1565), .Z(n1561) );
  ANDN U2078 ( .B(n1566), .A(n1567), .Z(n1564) );
  XNOR U2079 ( .A(b[144]), .B(n1565), .Z(n1566) );
  XNOR U2080 ( .A(b[144]), .B(n1567), .Z(c[144]) );
  XOR U2081 ( .A(n1568), .B(n1569), .Z(n1565) );
  ANDN U2082 ( .B(n1570), .A(n1571), .Z(n1568) );
  XNOR U2083 ( .A(b[143]), .B(n1569), .Z(n1570) );
  XNOR U2084 ( .A(b[143]), .B(n1571), .Z(c[143]) );
  XOR U2085 ( .A(n1572), .B(n1573), .Z(n1569) );
  ANDN U2086 ( .B(n1574), .A(n1575), .Z(n1572) );
  XNOR U2087 ( .A(b[142]), .B(n1573), .Z(n1574) );
  XNOR U2088 ( .A(b[142]), .B(n1575), .Z(c[142]) );
  XOR U2089 ( .A(n1576), .B(n1577), .Z(n1573) );
  ANDN U2090 ( .B(n1578), .A(n1579), .Z(n1576) );
  XNOR U2091 ( .A(b[141]), .B(n1577), .Z(n1578) );
  XNOR U2092 ( .A(b[141]), .B(n1579), .Z(c[141]) );
  XOR U2093 ( .A(n1580), .B(n1581), .Z(n1577) );
  ANDN U2094 ( .B(n1582), .A(n1583), .Z(n1580) );
  XNOR U2095 ( .A(b[140]), .B(n1581), .Z(n1582) );
  XNOR U2096 ( .A(b[140]), .B(n1583), .Z(c[140]) );
  XOR U2097 ( .A(n1584), .B(n1585), .Z(n1581) );
  ANDN U2098 ( .B(n1586), .A(n1587), .Z(n1584) );
  XNOR U2099 ( .A(b[139]), .B(n1585), .Z(n1586) );
  XNOR U2100 ( .A(b[13]), .B(n1588), .Z(c[13]) );
  XNOR U2101 ( .A(b[139]), .B(n1587), .Z(c[139]) );
  XOR U2102 ( .A(n1589), .B(n1590), .Z(n1585) );
  ANDN U2103 ( .B(n1591), .A(n1592), .Z(n1589) );
  XNOR U2104 ( .A(b[138]), .B(n1590), .Z(n1591) );
  XNOR U2105 ( .A(b[138]), .B(n1592), .Z(c[138]) );
  XOR U2106 ( .A(n1593), .B(n1594), .Z(n1590) );
  ANDN U2107 ( .B(n1595), .A(n1596), .Z(n1593) );
  XNOR U2108 ( .A(b[137]), .B(n1594), .Z(n1595) );
  XNOR U2109 ( .A(b[137]), .B(n1596), .Z(c[137]) );
  XOR U2110 ( .A(n1597), .B(n1598), .Z(n1594) );
  ANDN U2111 ( .B(n1599), .A(n1600), .Z(n1597) );
  XNOR U2112 ( .A(b[136]), .B(n1598), .Z(n1599) );
  XNOR U2113 ( .A(b[136]), .B(n1600), .Z(c[136]) );
  XOR U2114 ( .A(n1601), .B(n1602), .Z(n1598) );
  ANDN U2115 ( .B(n1603), .A(n1604), .Z(n1601) );
  XNOR U2116 ( .A(b[135]), .B(n1602), .Z(n1603) );
  XNOR U2117 ( .A(b[135]), .B(n1604), .Z(c[135]) );
  XOR U2118 ( .A(n1605), .B(n1606), .Z(n1602) );
  ANDN U2119 ( .B(n1607), .A(n1608), .Z(n1605) );
  XNOR U2120 ( .A(b[134]), .B(n1606), .Z(n1607) );
  XNOR U2121 ( .A(b[134]), .B(n1608), .Z(c[134]) );
  XOR U2122 ( .A(n1609), .B(n1610), .Z(n1606) );
  ANDN U2123 ( .B(n1611), .A(n1612), .Z(n1609) );
  XNOR U2124 ( .A(b[133]), .B(n1610), .Z(n1611) );
  XNOR U2125 ( .A(b[133]), .B(n1612), .Z(c[133]) );
  XOR U2126 ( .A(n1613), .B(n1614), .Z(n1610) );
  ANDN U2127 ( .B(n1615), .A(n1616), .Z(n1613) );
  XNOR U2128 ( .A(b[132]), .B(n1614), .Z(n1615) );
  XNOR U2129 ( .A(b[132]), .B(n1616), .Z(c[132]) );
  XOR U2130 ( .A(n1617), .B(n1618), .Z(n1614) );
  ANDN U2131 ( .B(n1619), .A(n1620), .Z(n1617) );
  XNOR U2132 ( .A(b[131]), .B(n1618), .Z(n1619) );
  XNOR U2133 ( .A(b[131]), .B(n1620), .Z(c[131]) );
  XOR U2134 ( .A(n1621), .B(n1622), .Z(n1618) );
  ANDN U2135 ( .B(n1623), .A(n1624), .Z(n1621) );
  XNOR U2136 ( .A(b[130]), .B(n1622), .Z(n1623) );
  XNOR U2137 ( .A(b[130]), .B(n1624), .Z(c[130]) );
  XOR U2138 ( .A(n1625), .B(n1626), .Z(n1622) );
  ANDN U2139 ( .B(n1627), .A(n1628), .Z(n1625) );
  XNOR U2140 ( .A(b[129]), .B(n1626), .Z(n1627) );
  XNOR U2141 ( .A(b[12]), .B(n1629), .Z(c[12]) );
  XNOR U2142 ( .A(b[129]), .B(n1628), .Z(c[129]) );
  XOR U2143 ( .A(n1630), .B(n1631), .Z(n1626) );
  ANDN U2144 ( .B(n1632), .A(n1633), .Z(n1630) );
  XNOR U2145 ( .A(b[128]), .B(n1631), .Z(n1632) );
  XNOR U2146 ( .A(b[128]), .B(n1633), .Z(c[128]) );
  XOR U2147 ( .A(n1634), .B(n1635), .Z(n1631) );
  ANDN U2148 ( .B(n1636), .A(n1637), .Z(n1634) );
  XNOR U2149 ( .A(b[127]), .B(n1635), .Z(n1636) );
  XNOR U2150 ( .A(b[127]), .B(n1637), .Z(c[127]) );
  XOR U2151 ( .A(n1638), .B(n1639), .Z(n1635) );
  ANDN U2152 ( .B(n1640), .A(n1641), .Z(n1638) );
  XNOR U2153 ( .A(b[126]), .B(n1639), .Z(n1640) );
  XNOR U2154 ( .A(b[126]), .B(n1641), .Z(c[126]) );
  XOR U2155 ( .A(n1642), .B(n1643), .Z(n1639) );
  ANDN U2156 ( .B(n1644), .A(n1645), .Z(n1642) );
  XNOR U2157 ( .A(b[125]), .B(n1643), .Z(n1644) );
  XNOR U2158 ( .A(b[125]), .B(n1645), .Z(c[125]) );
  XOR U2159 ( .A(n1646), .B(n1647), .Z(n1643) );
  ANDN U2160 ( .B(n1648), .A(n1649), .Z(n1646) );
  XNOR U2161 ( .A(b[124]), .B(n1647), .Z(n1648) );
  XNOR U2162 ( .A(b[124]), .B(n1649), .Z(c[124]) );
  XOR U2163 ( .A(n1650), .B(n1651), .Z(n1647) );
  ANDN U2164 ( .B(n1652), .A(n1653), .Z(n1650) );
  XNOR U2165 ( .A(b[123]), .B(n1651), .Z(n1652) );
  XNOR U2166 ( .A(b[123]), .B(n1653), .Z(c[123]) );
  XOR U2167 ( .A(n1654), .B(n1655), .Z(n1651) );
  ANDN U2168 ( .B(n1656), .A(n1657), .Z(n1654) );
  XNOR U2169 ( .A(b[122]), .B(n1655), .Z(n1656) );
  XNOR U2170 ( .A(b[122]), .B(n1657), .Z(c[122]) );
  XOR U2171 ( .A(n1658), .B(n1659), .Z(n1655) );
  ANDN U2172 ( .B(n1660), .A(n1661), .Z(n1658) );
  XNOR U2173 ( .A(b[121]), .B(n1659), .Z(n1660) );
  XNOR U2174 ( .A(b[121]), .B(n1661), .Z(c[121]) );
  XOR U2175 ( .A(n1662), .B(n1663), .Z(n1659) );
  ANDN U2176 ( .B(n1664), .A(n1665), .Z(n1662) );
  XNOR U2177 ( .A(b[120]), .B(n1663), .Z(n1664) );
  XNOR U2178 ( .A(b[120]), .B(n1665), .Z(c[120]) );
  XOR U2179 ( .A(n1666), .B(n1667), .Z(n1663) );
  ANDN U2180 ( .B(n1668), .A(n1669), .Z(n1666) );
  XNOR U2181 ( .A(b[119]), .B(n1667), .Z(n1668) );
  XNOR U2182 ( .A(b[11]), .B(n1670), .Z(c[11]) );
  XNOR U2183 ( .A(b[119]), .B(n1669), .Z(c[119]) );
  XOR U2184 ( .A(n1671), .B(n1672), .Z(n1667) );
  ANDN U2185 ( .B(n1673), .A(n1674), .Z(n1671) );
  XNOR U2186 ( .A(b[118]), .B(n1672), .Z(n1673) );
  XNOR U2187 ( .A(b[118]), .B(n1674), .Z(c[118]) );
  XOR U2188 ( .A(n1675), .B(n1676), .Z(n1672) );
  ANDN U2189 ( .B(n1677), .A(n1678), .Z(n1675) );
  XNOR U2190 ( .A(b[117]), .B(n1676), .Z(n1677) );
  XNOR U2191 ( .A(b[117]), .B(n1678), .Z(c[117]) );
  XOR U2192 ( .A(n1679), .B(n1680), .Z(n1676) );
  ANDN U2193 ( .B(n1681), .A(n1682), .Z(n1679) );
  XNOR U2194 ( .A(b[116]), .B(n1680), .Z(n1681) );
  XNOR U2195 ( .A(b[116]), .B(n1682), .Z(c[116]) );
  XOR U2196 ( .A(n1683), .B(n1684), .Z(n1680) );
  ANDN U2197 ( .B(n1685), .A(n1686), .Z(n1683) );
  XNOR U2198 ( .A(b[115]), .B(n1684), .Z(n1685) );
  XNOR U2199 ( .A(b[115]), .B(n1686), .Z(c[115]) );
  XOR U2200 ( .A(n1687), .B(n1688), .Z(n1684) );
  ANDN U2201 ( .B(n1689), .A(n1690), .Z(n1687) );
  XNOR U2202 ( .A(b[114]), .B(n1688), .Z(n1689) );
  XNOR U2203 ( .A(b[114]), .B(n1690), .Z(c[114]) );
  XOR U2204 ( .A(n1691), .B(n1692), .Z(n1688) );
  ANDN U2205 ( .B(n1693), .A(n1694), .Z(n1691) );
  XNOR U2206 ( .A(b[113]), .B(n1692), .Z(n1693) );
  XNOR U2207 ( .A(b[113]), .B(n1694), .Z(c[113]) );
  XOR U2208 ( .A(n1695), .B(n1696), .Z(n1692) );
  ANDN U2209 ( .B(n1697), .A(n1698), .Z(n1695) );
  XNOR U2210 ( .A(b[112]), .B(n1696), .Z(n1697) );
  XNOR U2211 ( .A(b[112]), .B(n1698), .Z(c[112]) );
  XOR U2212 ( .A(n1699), .B(n1700), .Z(n1696) );
  ANDN U2213 ( .B(n1701), .A(n1702), .Z(n1699) );
  XNOR U2214 ( .A(b[111]), .B(n1700), .Z(n1701) );
  XNOR U2215 ( .A(b[111]), .B(n1702), .Z(c[111]) );
  XOR U2216 ( .A(n1703), .B(n1704), .Z(n1700) );
  ANDN U2217 ( .B(n1705), .A(n1706), .Z(n1703) );
  XNOR U2218 ( .A(b[110]), .B(n1704), .Z(n1705) );
  XNOR U2219 ( .A(b[110]), .B(n1706), .Z(c[110]) );
  XOR U2220 ( .A(n1707), .B(n1708), .Z(n1704) );
  ANDN U2221 ( .B(n1709), .A(n1710), .Z(n1707) );
  XNOR U2222 ( .A(b[109]), .B(n1708), .Z(n1709) );
  XNOR U2223 ( .A(b[10]), .B(n1711), .Z(c[10]) );
  XNOR U2224 ( .A(b[109]), .B(n1710), .Z(c[109]) );
  XOR U2225 ( .A(n1712), .B(n1713), .Z(n1708) );
  ANDN U2226 ( .B(n1714), .A(n1715), .Z(n1712) );
  XNOR U2227 ( .A(b[108]), .B(n1713), .Z(n1714) );
  XNOR U2228 ( .A(b[108]), .B(n1715), .Z(c[108]) );
  XOR U2229 ( .A(n1716), .B(n1717), .Z(n1713) );
  ANDN U2230 ( .B(n1718), .A(n1719), .Z(n1716) );
  XNOR U2231 ( .A(b[107]), .B(n1717), .Z(n1718) );
  XNOR U2232 ( .A(b[107]), .B(n1719), .Z(c[107]) );
  XOR U2233 ( .A(n1720), .B(n1721), .Z(n1717) );
  ANDN U2234 ( .B(n1722), .A(n1723), .Z(n1720) );
  XNOR U2235 ( .A(b[106]), .B(n1721), .Z(n1722) );
  XNOR U2236 ( .A(b[106]), .B(n1723), .Z(c[106]) );
  XOR U2237 ( .A(n1724), .B(n1725), .Z(n1721) );
  ANDN U2238 ( .B(n1726), .A(n1727), .Z(n1724) );
  XNOR U2239 ( .A(b[105]), .B(n1725), .Z(n1726) );
  XNOR U2240 ( .A(b[105]), .B(n1727), .Z(c[105]) );
  XOR U2241 ( .A(n1728), .B(n1729), .Z(n1725) );
  ANDN U2242 ( .B(n1730), .A(n1731), .Z(n1728) );
  XNOR U2243 ( .A(b[104]), .B(n1729), .Z(n1730) );
  XNOR U2244 ( .A(b[104]), .B(n1731), .Z(c[104]) );
  XOR U2245 ( .A(n1732), .B(n1733), .Z(n1729) );
  ANDN U2246 ( .B(n1734), .A(n1735), .Z(n1732) );
  XNOR U2247 ( .A(b[103]), .B(n1733), .Z(n1734) );
  XNOR U2248 ( .A(b[103]), .B(n1735), .Z(c[103]) );
  XOR U2249 ( .A(n1736), .B(n1737), .Z(n1733) );
  ANDN U2250 ( .B(n1738), .A(n1739), .Z(n1736) );
  XNOR U2251 ( .A(b[102]), .B(n1737), .Z(n1738) );
  XNOR U2252 ( .A(b[102]), .B(n1739), .Z(c[102]) );
  XOR U2253 ( .A(n1740), .B(n1741), .Z(n1737) );
  ANDN U2254 ( .B(n1742), .A(n1743), .Z(n1740) );
  XNOR U2255 ( .A(b[101]), .B(n1741), .Z(n1742) );
  XNOR U2256 ( .A(b[101]), .B(n1743), .Z(c[101]) );
  XOR U2257 ( .A(n1744), .B(n1745), .Z(n1741) );
  ANDN U2258 ( .B(n1746), .A(n1747), .Z(n1744) );
  XNOR U2259 ( .A(b[100]), .B(n1745), .Z(n1746) );
  XNOR U2260 ( .A(b[100]), .B(n1747), .Z(c[100]) );
  XOR U2261 ( .A(n1748), .B(n1749), .Z(n1745) );
  ANDN U2262 ( .B(n1750), .A(n6), .Z(n1748) );
  XNOR U2263 ( .A(b[99]), .B(n1749), .Z(n1750) );
  XOR U2264 ( .A(n1751), .B(n1752), .Z(n1749) );
  ANDN U2265 ( .B(n1753), .A(n7), .Z(n1751) );
  XNOR U2266 ( .A(b[98]), .B(n1752), .Z(n1753) );
  XOR U2267 ( .A(n1754), .B(n1755), .Z(n1752) );
  ANDN U2268 ( .B(n1756), .A(n8), .Z(n1754) );
  XNOR U2269 ( .A(b[97]), .B(n1755), .Z(n1756) );
  XOR U2270 ( .A(n1757), .B(n1758), .Z(n1755) );
  ANDN U2271 ( .B(n1759), .A(n9), .Z(n1757) );
  XNOR U2272 ( .A(b[96]), .B(n1758), .Z(n1759) );
  XOR U2273 ( .A(n1760), .B(n1761), .Z(n1758) );
  ANDN U2274 ( .B(n1762), .A(n10), .Z(n1760) );
  XNOR U2275 ( .A(b[95]), .B(n1761), .Z(n1762) );
  XOR U2276 ( .A(n1763), .B(n1764), .Z(n1761) );
  ANDN U2277 ( .B(n1765), .A(n11), .Z(n1763) );
  XNOR U2278 ( .A(b[94]), .B(n1764), .Z(n1765) );
  XOR U2279 ( .A(n1766), .B(n1767), .Z(n1764) );
  ANDN U2280 ( .B(n1768), .A(n12), .Z(n1766) );
  XNOR U2281 ( .A(b[93]), .B(n1767), .Z(n1768) );
  XOR U2282 ( .A(n1769), .B(n1770), .Z(n1767) );
  ANDN U2283 ( .B(n1771), .A(n13), .Z(n1769) );
  XNOR U2284 ( .A(b[92]), .B(n1770), .Z(n1771) );
  XOR U2285 ( .A(n1772), .B(n1773), .Z(n1770) );
  ANDN U2286 ( .B(n1774), .A(n14), .Z(n1772) );
  XNOR U2287 ( .A(b[91]), .B(n1773), .Z(n1774) );
  XOR U2288 ( .A(n1775), .B(n1776), .Z(n1773) );
  ANDN U2289 ( .B(n1777), .A(n15), .Z(n1775) );
  XNOR U2290 ( .A(b[90]), .B(n1776), .Z(n1777) );
  XOR U2291 ( .A(n1778), .B(n1779), .Z(n1776) );
  ANDN U2292 ( .B(n1780), .A(n17), .Z(n1778) );
  XNOR U2293 ( .A(b[89]), .B(n1779), .Z(n1780) );
  XOR U2294 ( .A(n1781), .B(n1782), .Z(n1779) );
  ANDN U2295 ( .B(n1783), .A(n18), .Z(n1781) );
  XNOR U2296 ( .A(b[88]), .B(n1782), .Z(n1783) );
  XOR U2297 ( .A(n1784), .B(n1785), .Z(n1782) );
  ANDN U2298 ( .B(n1786), .A(n19), .Z(n1784) );
  XNOR U2299 ( .A(b[87]), .B(n1785), .Z(n1786) );
  XOR U2300 ( .A(n1787), .B(n1788), .Z(n1785) );
  ANDN U2301 ( .B(n1789), .A(n20), .Z(n1787) );
  XNOR U2302 ( .A(b[86]), .B(n1788), .Z(n1789) );
  XOR U2303 ( .A(n1790), .B(n1791), .Z(n1788) );
  ANDN U2304 ( .B(n1792), .A(n21), .Z(n1790) );
  XNOR U2305 ( .A(b[85]), .B(n1791), .Z(n1792) );
  XOR U2306 ( .A(n1793), .B(n1794), .Z(n1791) );
  ANDN U2307 ( .B(n1795), .A(n22), .Z(n1793) );
  XNOR U2308 ( .A(b[84]), .B(n1794), .Z(n1795) );
  XOR U2309 ( .A(n1796), .B(n1797), .Z(n1794) );
  ANDN U2310 ( .B(n1798), .A(n23), .Z(n1796) );
  XNOR U2311 ( .A(b[83]), .B(n1797), .Z(n1798) );
  XOR U2312 ( .A(n1799), .B(n1800), .Z(n1797) );
  ANDN U2313 ( .B(n1801), .A(n24), .Z(n1799) );
  XNOR U2314 ( .A(b[82]), .B(n1800), .Z(n1801) );
  XOR U2315 ( .A(n1802), .B(n1803), .Z(n1800) );
  ANDN U2316 ( .B(n1804), .A(n25), .Z(n1802) );
  XNOR U2317 ( .A(b[81]), .B(n1803), .Z(n1804) );
  XOR U2318 ( .A(n1805), .B(n1806), .Z(n1803) );
  ANDN U2319 ( .B(n1807), .A(n26), .Z(n1805) );
  XNOR U2320 ( .A(b[80]), .B(n1806), .Z(n1807) );
  XOR U2321 ( .A(n1808), .B(n1809), .Z(n1806) );
  ANDN U2322 ( .B(n1810), .A(n28), .Z(n1808) );
  XNOR U2323 ( .A(b[79]), .B(n1809), .Z(n1810) );
  XOR U2324 ( .A(n1811), .B(n1812), .Z(n1809) );
  ANDN U2325 ( .B(n1813), .A(n29), .Z(n1811) );
  XNOR U2326 ( .A(b[78]), .B(n1812), .Z(n1813) );
  XOR U2327 ( .A(n1814), .B(n1815), .Z(n1812) );
  ANDN U2328 ( .B(n1816), .A(n30), .Z(n1814) );
  XNOR U2329 ( .A(b[77]), .B(n1815), .Z(n1816) );
  XOR U2330 ( .A(n1817), .B(n1818), .Z(n1815) );
  ANDN U2331 ( .B(n1819), .A(n31), .Z(n1817) );
  XNOR U2332 ( .A(b[76]), .B(n1818), .Z(n1819) );
  XOR U2333 ( .A(n1820), .B(n1821), .Z(n1818) );
  ANDN U2334 ( .B(n1822), .A(n32), .Z(n1820) );
  XNOR U2335 ( .A(b[75]), .B(n1821), .Z(n1822) );
  XOR U2336 ( .A(n1823), .B(n1824), .Z(n1821) );
  ANDN U2337 ( .B(n1825), .A(n33), .Z(n1823) );
  XNOR U2338 ( .A(b[74]), .B(n1824), .Z(n1825) );
  XOR U2339 ( .A(n1826), .B(n1827), .Z(n1824) );
  ANDN U2340 ( .B(n1828), .A(n34), .Z(n1826) );
  XNOR U2341 ( .A(b[73]), .B(n1827), .Z(n1828) );
  XOR U2342 ( .A(n1829), .B(n1830), .Z(n1827) );
  ANDN U2343 ( .B(n1831), .A(n35), .Z(n1829) );
  XNOR U2344 ( .A(b[72]), .B(n1830), .Z(n1831) );
  XOR U2345 ( .A(n1832), .B(n1833), .Z(n1830) );
  ANDN U2346 ( .B(n1834), .A(n36), .Z(n1832) );
  XNOR U2347 ( .A(b[71]), .B(n1833), .Z(n1834) );
  XOR U2348 ( .A(n1835), .B(n1836), .Z(n1833) );
  ANDN U2349 ( .B(n1837), .A(n37), .Z(n1835) );
  XNOR U2350 ( .A(b[70]), .B(n1836), .Z(n1837) );
  XOR U2351 ( .A(n1838), .B(n1839), .Z(n1836) );
  ANDN U2352 ( .B(n1840), .A(n39), .Z(n1838) );
  XNOR U2353 ( .A(b[69]), .B(n1839), .Z(n1840) );
  XOR U2354 ( .A(n1841), .B(n1842), .Z(n1839) );
  ANDN U2355 ( .B(n1843), .A(n40), .Z(n1841) );
  XNOR U2356 ( .A(b[68]), .B(n1842), .Z(n1843) );
  XOR U2357 ( .A(n1844), .B(n1845), .Z(n1842) );
  ANDN U2358 ( .B(n1846), .A(n41), .Z(n1844) );
  XNOR U2359 ( .A(b[67]), .B(n1845), .Z(n1846) );
  XOR U2360 ( .A(n1847), .B(n1848), .Z(n1845) );
  ANDN U2361 ( .B(n1849), .A(n42), .Z(n1847) );
  XNOR U2362 ( .A(b[66]), .B(n1848), .Z(n1849) );
  XOR U2363 ( .A(n1850), .B(n1851), .Z(n1848) );
  ANDN U2364 ( .B(n1852), .A(n43), .Z(n1850) );
  XNOR U2365 ( .A(b[65]), .B(n1851), .Z(n1852) );
  XOR U2366 ( .A(n1853), .B(n1854), .Z(n1851) );
  ANDN U2367 ( .B(n1855), .A(n44), .Z(n1853) );
  XNOR U2368 ( .A(b[64]), .B(n1854), .Z(n1855) );
  XOR U2369 ( .A(n1856), .B(n1857), .Z(n1854) );
  ANDN U2370 ( .B(n1858), .A(n45), .Z(n1856) );
  XNOR U2371 ( .A(b[63]), .B(n1857), .Z(n1858) );
  XOR U2372 ( .A(n1859), .B(n1860), .Z(n1857) );
  ANDN U2373 ( .B(n1861), .A(n46), .Z(n1859) );
  XNOR U2374 ( .A(b[62]), .B(n1860), .Z(n1861) );
  XOR U2375 ( .A(n1862), .B(n1863), .Z(n1860) );
  ANDN U2376 ( .B(n1864), .A(n47), .Z(n1862) );
  XNOR U2377 ( .A(b[61]), .B(n1863), .Z(n1864) );
  XOR U2378 ( .A(n1865), .B(n1866), .Z(n1863) );
  ANDN U2379 ( .B(n1867), .A(n48), .Z(n1865) );
  XNOR U2380 ( .A(b[60]), .B(n1866), .Z(n1867) );
  XOR U2381 ( .A(n1868), .B(n1869), .Z(n1866) );
  ANDN U2382 ( .B(n1870), .A(n50), .Z(n1868) );
  XNOR U2383 ( .A(b[59]), .B(n1869), .Z(n1870) );
  XOR U2384 ( .A(n1871), .B(n1872), .Z(n1869) );
  ANDN U2385 ( .B(n1873), .A(n51), .Z(n1871) );
  XNOR U2386 ( .A(b[58]), .B(n1872), .Z(n1873) );
  XOR U2387 ( .A(n1874), .B(n1875), .Z(n1872) );
  ANDN U2388 ( .B(n1876), .A(n52), .Z(n1874) );
  XNOR U2389 ( .A(b[57]), .B(n1875), .Z(n1876) );
  XOR U2390 ( .A(n1877), .B(n1878), .Z(n1875) );
  ANDN U2391 ( .B(n1879), .A(n53), .Z(n1877) );
  XNOR U2392 ( .A(b[56]), .B(n1878), .Z(n1879) );
  XOR U2393 ( .A(n1880), .B(n1881), .Z(n1878) );
  ANDN U2394 ( .B(n1882), .A(n54), .Z(n1880) );
  XNOR U2395 ( .A(b[55]), .B(n1881), .Z(n1882) );
  XOR U2396 ( .A(n1883), .B(n1884), .Z(n1881) );
  ANDN U2397 ( .B(n1885), .A(n55), .Z(n1883) );
  XNOR U2398 ( .A(b[54]), .B(n1884), .Z(n1885) );
  XOR U2399 ( .A(n1886), .B(n1887), .Z(n1884) );
  ANDN U2400 ( .B(n1888), .A(n56), .Z(n1886) );
  XNOR U2401 ( .A(b[53]), .B(n1887), .Z(n1888) );
  XOR U2402 ( .A(n1889), .B(n1890), .Z(n1887) );
  ANDN U2403 ( .B(n1891), .A(n57), .Z(n1889) );
  XNOR U2404 ( .A(b[52]), .B(n1890), .Z(n1891) );
  XOR U2405 ( .A(n1892), .B(n1893), .Z(n1890) );
  ANDN U2406 ( .B(n1894), .A(n58), .Z(n1892) );
  XNOR U2407 ( .A(b[51]), .B(n1893), .Z(n1894) );
  XOR U2408 ( .A(n1895), .B(n1896), .Z(n1893) );
  ANDN U2409 ( .B(n1897), .A(n67), .Z(n1895) );
  XNOR U2410 ( .A(b[50]), .B(n1896), .Z(n1897) );
  XOR U2411 ( .A(n1898), .B(n1899), .Z(n1896) );
  ANDN U2412 ( .B(n1900), .A(n109), .Z(n1898) );
  XNOR U2413 ( .A(b[49]), .B(n1899), .Z(n1900) );
  XOR U2414 ( .A(n1901), .B(n1902), .Z(n1899) );
  ANDN U2415 ( .B(n1903), .A(n150), .Z(n1901) );
  XNOR U2416 ( .A(b[48]), .B(n1902), .Z(n1903) );
  XOR U2417 ( .A(n1904), .B(n1905), .Z(n1902) );
  ANDN U2418 ( .B(n1906), .A(n191), .Z(n1904) );
  XNOR U2419 ( .A(b[47]), .B(n1905), .Z(n1906) );
  XOR U2420 ( .A(n1907), .B(n1908), .Z(n1905) );
  ANDN U2421 ( .B(n1909), .A(n232), .Z(n1907) );
  XNOR U2422 ( .A(b[46]), .B(n1908), .Z(n1909) );
  XOR U2423 ( .A(n1910), .B(n1911), .Z(n1908) );
  ANDN U2424 ( .B(n1912), .A(n273), .Z(n1910) );
  XNOR U2425 ( .A(b[45]), .B(n1911), .Z(n1912) );
  XOR U2426 ( .A(n1913), .B(n1914), .Z(n1911) );
  ANDN U2427 ( .B(n1915), .A(n314), .Z(n1913) );
  XNOR U2428 ( .A(b[44]), .B(n1914), .Z(n1915) );
  XOR U2429 ( .A(n1916), .B(n1917), .Z(n1914) );
  ANDN U2430 ( .B(n1918), .A(n355), .Z(n1916) );
  XNOR U2431 ( .A(b[43]), .B(n1917), .Z(n1918) );
  XOR U2432 ( .A(n1919), .B(n1920), .Z(n1917) );
  ANDN U2433 ( .B(n1921), .A(n396), .Z(n1919) );
  XNOR U2434 ( .A(b[42]), .B(n1920), .Z(n1921) );
  XOR U2435 ( .A(n1922), .B(n1923), .Z(n1920) );
  ANDN U2436 ( .B(n1924), .A(n437), .Z(n1922) );
  XNOR U2437 ( .A(b[41]), .B(n1923), .Z(n1924) );
  XOR U2438 ( .A(n1925), .B(n1926), .Z(n1923) );
  ANDN U2439 ( .B(n1927), .A(n478), .Z(n1925) );
  XNOR U2440 ( .A(b[40]), .B(n1926), .Z(n1927) );
  XOR U2441 ( .A(n1928), .B(n1929), .Z(n1926) );
  ANDN U2442 ( .B(n1930), .A(n520), .Z(n1928) );
  XNOR U2443 ( .A(b[39]), .B(n1929), .Z(n1930) );
  XOR U2444 ( .A(n1931), .B(n1932), .Z(n1929) );
  ANDN U2445 ( .B(n1933), .A(n561), .Z(n1931) );
  XNOR U2446 ( .A(b[38]), .B(n1932), .Z(n1933) );
  XOR U2447 ( .A(n1934), .B(n1935), .Z(n1932) );
  ANDN U2448 ( .B(n1936), .A(n602), .Z(n1934) );
  XNOR U2449 ( .A(b[37]), .B(n1935), .Z(n1936) );
  XOR U2450 ( .A(n1937), .B(n1938), .Z(n1935) );
  ANDN U2451 ( .B(n1939), .A(n643), .Z(n1937) );
  XNOR U2452 ( .A(b[36]), .B(n1938), .Z(n1939) );
  XOR U2453 ( .A(n1940), .B(n1941), .Z(n1938) );
  ANDN U2454 ( .B(n1942), .A(n684), .Z(n1940) );
  XNOR U2455 ( .A(b[35]), .B(n1941), .Z(n1942) );
  XOR U2456 ( .A(n1943), .B(n1944), .Z(n1941) );
  ANDN U2457 ( .B(n1945), .A(n725), .Z(n1943) );
  XNOR U2458 ( .A(b[34]), .B(n1944), .Z(n1945) );
  XOR U2459 ( .A(n1946), .B(n1947), .Z(n1944) );
  ANDN U2460 ( .B(n1948), .A(n766), .Z(n1946) );
  XNOR U2461 ( .A(b[33]), .B(n1947), .Z(n1948) );
  XOR U2462 ( .A(n1949), .B(n1950), .Z(n1947) );
  ANDN U2463 ( .B(n1951), .A(n807), .Z(n1949) );
  XNOR U2464 ( .A(b[32]), .B(n1950), .Z(n1951) );
  XOR U2465 ( .A(n1952), .B(n1953), .Z(n1950) );
  ANDN U2466 ( .B(n1954), .A(n848), .Z(n1952) );
  XNOR U2467 ( .A(b[31]), .B(n1953), .Z(n1954) );
  XOR U2468 ( .A(n1955), .B(n1956), .Z(n1953) );
  ANDN U2469 ( .B(n1957), .A(n889), .Z(n1955) );
  XNOR U2470 ( .A(b[30]), .B(n1956), .Z(n1957) );
  XOR U2471 ( .A(n1958), .B(n1959), .Z(n1956) );
  ANDN U2472 ( .B(n1960), .A(n931), .Z(n1958) );
  XNOR U2473 ( .A(b[29]), .B(n1959), .Z(n1960) );
  XOR U2474 ( .A(n1961), .B(n1962), .Z(n1959) );
  ANDN U2475 ( .B(n1963), .A(n972), .Z(n1961) );
  XNOR U2476 ( .A(b[28]), .B(n1962), .Z(n1963) );
  XOR U2477 ( .A(n1964), .B(n1965), .Z(n1962) );
  ANDN U2478 ( .B(n1966), .A(n1013), .Z(n1964) );
  XNOR U2479 ( .A(b[27]), .B(n1965), .Z(n1966) );
  XOR U2480 ( .A(n1967), .B(n1968), .Z(n1965) );
  ANDN U2481 ( .B(n1969), .A(n1054), .Z(n1967) );
  XNOR U2482 ( .A(b[26]), .B(n1968), .Z(n1969) );
  XOR U2483 ( .A(n1970), .B(n1971), .Z(n1968) );
  ANDN U2484 ( .B(n1972), .A(n1095), .Z(n1970) );
  XNOR U2485 ( .A(b[25]), .B(n1971), .Z(n1972) );
  XOR U2486 ( .A(n1973), .B(n1974), .Z(n1971) );
  ANDN U2487 ( .B(n1975), .A(n1136), .Z(n1973) );
  XNOR U2488 ( .A(b[24]), .B(n1974), .Z(n1975) );
  XOR U2489 ( .A(n1976), .B(n1977), .Z(n1974) );
  ANDN U2490 ( .B(n1978), .A(n1177), .Z(n1976) );
  XNOR U2491 ( .A(b[23]), .B(n1977), .Z(n1978) );
  XOR U2492 ( .A(n1979), .B(n1980), .Z(n1977) );
  ANDN U2493 ( .B(n1981), .A(n1218), .Z(n1979) );
  XNOR U2494 ( .A(b[22]), .B(n1980), .Z(n1981) );
  XOR U2495 ( .A(n1982), .B(n1983), .Z(n1980) );
  ANDN U2496 ( .B(n1984), .A(n1259), .Z(n1982) );
  XNOR U2497 ( .A(b[21]), .B(n1983), .Z(n1984) );
  XOR U2498 ( .A(n1985), .B(n1986), .Z(n1983) );
  ANDN U2499 ( .B(n1987), .A(n1300), .Z(n1985) );
  XNOR U2500 ( .A(b[20]), .B(n1986), .Z(n1987) );
  XOR U2501 ( .A(n1988), .B(n1989), .Z(n1986) );
  ANDN U2502 ( .B(n1990), .A(n1342), .Z(n1988) );
  XNOR U2503 ( .A(b[19]), .B(n1989), .Z(n1990) );
  XOR U2504 ( .A(n1991), .B(n1992), .Z(n1989) );
  ANDN U2505 ( .B(n1993), .A(n1383), .Z(n1991) );
  XNOR U2506 ( .A(b[18]), .B(n1992), .Z(n1993) );
  XOR U2507 ( .A(n1994), .B(n1995), .Z(n1992) );
  ANDN U2508 ( .B(n1996), .A(n1424), .Z(n1994) );
  XNOR U2509 ( .A(b[17]), .B(n1995), .Z(n1996) );
  XOR U2510 ( .A(n1997), .B(n1998), .Z(n1995) );
  ANDN U2511 ( .B(n1999), .A(n1465), .Z(n1997) );
  XNOR U2512 ( .A(b[16]), .B(n1998), .Z(n1999) );
  XOR U2513 ( .A(n2000), .B(n2001), .Z(n1998) );
  ANDN U2514 ( .B(n2002), .A(n1506), .Z(n2000) );
  XNOR U2515 ( .A(b[15]), .B(n2001), .Z(n2002) );
  XOR U2516 ( .A(n2003), .B(n2004), .Z(n2001) );
  ANDN U2517 ( .B(n2005), .A(n1547), .Z(n2003) );
  XNOR U2518 ( .A(b[14]), .B(n2004), .Z(n2005) );
  XOR U2519 ( .A(n2006), .B(n2007), .Z(n2004) );
  ANDN U2520 ( .B(n2008), .A(n1588), .Z(n2006) );
  XNOR U2521 ( .A(b[13]), .B(n2007), .Z(n2008) );
  XOR U2522 ( .A(n2009), .B(n2010), .Z(n2007) );
  ANDN U2523 ( .B(n2011), .A(n1629), .Z(n2009) );
  XNOR U2524 ( .A(b[12]), .B(n2010), .Z(n2011) );
  XOR U2525 ( .A(n2012), .B(n2013), .Z(n2010) );
  ANDN U2526 ( .B(n2014), .A(n1670), .Z(n2012) );
  XNOR U2527 ( .A(b[11]), .B(n2013), .Z(n2014) );
  XOR U2528 ( .A(n2015), .B(n2016), .Z(n2013) );
  ANDN U2529 ( .B(n2017), .A(n1711), .Z(n2015) );
  XNOR U2530 ( .A(b[10]), .B(n2016), .Z(n2017) );
  XOR U2531 ( .A(n2018), .B(n2019), .Z(n2016) );
  ANDN U2532 ( .B(n2020), .A(n5), .Z(n2018) );
  XNOR U2533 ( .A(b[9]), .B(n2019), .Z(n2020) );
  XOR U2534 ( .A(n2021), .B(n2022), .Z(n2019) );
  ANDN U2535 ( .B(n2023), .A(n16), .Z(n2021) );
  XNOR U2536 ( .A(b[8]), .B(n2022), .Z(n2023) );
  XOR U2537 ( .A(n2024), .B(n2025), .Z(n2022) );
  ANDN U2538 ( .B(n2026), .A(n27), .Z(n2024) );
  XNOR U2539 ( .A(b[7]), .B(n2025), .Z(n2026) );
  XOR U2540 ( .A(n2027), .B(n2028), .Z(n2025) );
  ANDN U2541 ( .B(n2029), .A(n38), .Z(n2027) );
  XNOR U2542 ( .A(b[6]), .B(n2028), .Z(n2029) );
  XOR U2543 ( .A(n2030), .B(n2031), .Z(n2028) );
  ANDN U2544 ( .B(n2032), .A(n49), .Z(n2030) );
  XNOR U2545 ( .A(b[5]), .B(n2031), .Z(n2032) );
  XOR U2546 ( .A(n2033), .B(n2034), .Z(n2031) );
  ANDN U2547 ( .B(n2035), .A(n108), .Z(n2033) );
  XNOR U2548 ( .A(b[4]), .B(n2034), .Z(n2035) );
  XOR U2549 ( .A(n2036), .B(n2037), .Z(n2034) );
  ANDN U2550 ( .B(n2038), .A(n519), .Z(n2036) );
  XNOR U2551 ( .A(b[3]), .B(n2037), .Z(n2038) );
  XOR U2552 ( .A(n2039), .B(n2040), .Z(n2037) );
  ANDN U2553 ( .B(n2041), .A(n930), .Z(n2039) );
  XNOR U2554 ( .A(b[2]), .B(n2040), .Z(n2041) );
  XOR U2555 ( .A(n2042), .B(n2043), .Z(n2040) );
  ANDN U2556 ( .B(n2044), .A(n1341), .Z(n2042) );
  XNOR U2557 ( .A(b[1]), .B(n2043), .Z(n2044) );
  XOR U2558 ( .A(carry_on), .B(n2045), .Z(n2043) );
  NANDN U2559 ( .A(n2046), .B(n2047), .Z(n2045) );
  XOR U2560 ( .A(carry_on), .B(b[0]), .Z(n2047) );
  XNOR U2561 ( .A(b[0]), .B(n2046), .Z(c[0]) );
  XNOR U2562 ( .A(a[0]), .B(carry_on), .Z(n2046) );
endmodule

