
module hamming_N1600_CC16 ( clk, rst, x, y, o );
  input [99:0] x;
  input [99:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[10]) );
  XOR U114 ( .A(n401), .B(n400), .Z(n398) );
  XOR U115 ( .A(n447), .B(n446), .Z(n444) );
  XOR U116 ( .A(n359), .B(n358), .Z(n356) );
  XOR U117 ( .A(n315), .B(n314), .Z(n312) );
  XOR U118 ( .A(n243), .B(n245), .Z(n251) );
  XOR U119 ( .A(n73), .B(n77), .Z(n113) );
  XNOR U120 ( .A(oglobal[4]), .B(n50), .Z(n16) );
  XOR U121 ( .A(n335), .B(n334), .Z(n355) );
  XNOR U122 ( .A(n277), .B(n412), .Z(n249) );
  XOR U123 ( .A(n312), .B(n311), .Z(n344) );
  XNOR U124 ( .A(n145), .B(n212), .Z(n116) );
  XNOR U125 ( .A(oglobal[3]), .B(n82), .Z(n18) );
  XOR U126 ( .A(n156), .B(n158), .Z(n177) );
  XOR U127 ( .A(n379), .B(n378), .Z(n397) );
  XOR U128 ( .A(n423), .B(n422), .Z(n443) );
  XOR U129 ( .A(n91), .B(n93), .Z(n112) );
  XNOR U130 ( .A(n209), .B(n324), .Z(n182) );
  XNOR U131 ( .A(n249), .B(n368), .Z(n216) );
  XNOR U132 ( .A(oglobal[5]), .B(n35), .Z(n14) );
  XNOR U133 ( .A(oglobal[2]), .B(n148), .Z(n20) );
  XOR U134 ( .A(n12), .B(n13), .Z(o[6]) );
  XNOR U135 ( .A(n14), .B(n15), .Z(o[5]) );
  XNOR U136 ( .A(n16), .B(n17), .Z(o[4]) );
  XOR U137 ( .A(n18), .B(n19), .Z(o[3]) );
  XOR U138 ( .A(n20), .B(n21), .Z(o[2]) );
  XOR U139 ( .A(n22), .B(n23), .Z(o[1]) );
  XOR U140 ( .A(n24), .B(n25), .Z(o[10]) );
  XOR U141 ( .A(oglobal[10]), .B(n26), .Z(n25) );
  AND U142 ( .A(n24), .B(o[9]), .Z(n26) );
  XOR U143 ( .A(oglobal[9]), .B(n24), .Z(o[9]) );
  NOR U144 ( .A(o[8]), .B(n27), .Z(n24) );
  XNOR U145 ( .A(oglobal[8]), .B(n27), .Z(o[8]) );
  OR U146 ( .A(o[7]), .B(n28), .Z(n27) );
  XNOR U147 ( .A(oglobal[7]), .B(n28), .Z(o[7]) );
  XNOR U148 ( .A(n29), .B(n30), .Z(n28) );
  ANDN U149 ( .B(n31), .A(n13), .Z(n29) );
  XNOR U150 ( .A(oglobal[6]), .B(n30), .Z(n13) );
  NANDN U151 ( .A(n30), .B(n12), .Z(n31) );
  OR U152 ( .A(n32), .B(n33), .Z(n12) );
  XOR U153 ( .A(n34), .B(n35), .Z(n30) );
  ANDN U154 ( .B(n36), .A(n14), .Z(n34) );
  XOR U155 ( .A(n35), .B(n15), .Z(n36) );
  XOR U156 ( .A(n32), .B(n33), .Z(n15) );
  AND U157 ( .A(n37), .B(n38), .Z(n33) );
  OR U158 ( .A(n39), .B(n40), .Z(n38) );
  XOR U159 ( .A(n41), .B(n42), .Z(n37) );
  ANDN U160 ( .B(n43), .A(n44), .Z(n41) );
  XOR U161 ( .A(n45), .B(n46), .Z(n43) );
  OR U162 ( .A(n47), .B(n48), .Z(n32) );
  XOR U163 ( .A(n49), .B(n50), .Z(n35) );
  ANDN U164 ( .B(n51), .A(n16), .Z(n49) );
  XOR U165 ( .A(n50), .B(n17), .Z(n51) );
  XNOR U166 ( .A(n44), .B(n46), .Z(n17) );
  XOR U167 ( .A(n47), .B(n48), .Z(n46) );
  AND U168 ( .A(n52), .B(n53), .Z(n48) );
  OR U169 ( .A(n54), .B(n55), .Z(n53) );
  XOR U170 ( .A(n56), .B(n57), .Z(n52) );
  ANDN U171 ( .B(n58), .A(n59), .Z(n56) );
  XOR U172 ( .A(n60), .B(n61), .Z(n58) );
  OR U173 ( .A(n62), .B(n63), .Z(n47) );
  XOR U174 ( .A(n42), .B(n64), .Z(n44) );
  XOR U175 ( .A(n39), .B(n40), .Z(n64) );
  AND U176 ( .A(n65), .B(n66), .Z(n40) );
  OR U177 ( .A(n67), .B(n68), .Z(n66) );
  XOR U178 ( .A(n69), .B(n70), .Z(n65) );
  AND U179 ( .A(n71), .B(n72), .Z(n69) );
  XNOR U180 ( .A(n73), .B(n70), .Z(n72) );
  OR U181 ( .A(n74), .B(n75), .Z(n39) );
  IV U182 ( .A(n45), .Z(n42) );
  XOR U183 ( .A(n76), .B(n77), .Z(n45) );
  AND U184 ( .A(n78), .B(n79), .Z(n76) );
  XOR U185 ( .A(n77), .B(n80), .Z(n79) );
  XOR U186 ( .A(n81), .B(n82), .Z(n50) );
  ANDN U187 ( .B(n83), .A(n18), .Z(n81) );
  XNOR U188 ( .A(n82), .B(n19), .Z(n83) );
  XNOR U189 ( .A(n78), .B(n80), .Z(n19) );
  XNOR U190 ( .A(n59), .B(n61), .Z(n80) );
  XOR U191 ( .A(n62), .B(n63), .Z(n61) );
  AND U192 ( .A(n84), .B(n85), .Z(n63) );
  OR U193 ( .A(n86), .B(n87), .Z(n85) );
  XOR U194 ( .A(n88), .B(n89), .Z(n84) );
  AND U195 ( .A(n90), .B(n91), .Z(n88) );
  XOR U196 ( .A(n92), .B(n93), .Z(n90) );
  OR U197 ( .A(n94), .B(n95), .Z(n62) );
  XOR U198 ( .A(n57), .B(n96), .Z(n59) );
  XOR U199 ( .A(n54), .B(n55), .Z(n96) );
  AND U200 ( .A(n97), .B(n98), .Z(n55) );
  OR U201 ( .A(n99), .B(n100), .Z(n98) );
  XOR U202 ( .A(n101), .B(n102), .Z(n97) );
  AND U203 ( .A(n103), .B(n104), .Z(n101) );
  XNOR U204 ( .A(n105), .B(n102), .Z(n104) );
  OR U205 ( .A(n106), .B(n107), .Z(n54) );
  IV U206 ( .A(n60), .Z(n57) );
  XNOR U207 ( .A(n108), .B(n109), .Z(n60) );
  AND U208 ( .A(n110), .B(n111), .Z(n108) );
  XNOR U209 ( .A(n109), .B(n112), .Z(n111) );
  XOR U210 ( .A(n71), .B(n113), .Z(n78) );
  XNOR U211 ( .A(n114), .B(n115), .Z(n77) );
  AND U212 ( .A(n116), .B(n117), .Z(n114) );
  XNOR U213 ( .A(n115), .B(n118), .Z(n117) );
  XOR U214 ( .A(n74), .B(n75), .Z(n73) );
  AND U215 ( .A(n119), .B(n120), .Z(n75) );
  OR U216 ( .A(n121), .B(n122), .Z(n120) );
  XOR U217 ( .A(n123), .B(n124), .Z(n119) );
  ANDN U218 ( .B(n125), .A(n126), .Z(n123) );
  XOR U219 ( .A(n124), .B(n127), .Z(n125) );
  OR U220 ( .A(n128), .B(n129), .Z(n74) );
  XNOR U221 ( .A(n70), .B(n130), .Z(n71) );
  XOR U222 ( .A(n67), .B(n68), .Z(n130) );
  AND U223 ( .A(n131), .B(n132), .Z(n68) );
  OR U224 ( .A(n133), .B(n134), .Z(n132) );
  XOR U225 ( .A(n135), .B(n136), .Z(n131) );
  AND U226 ( .A(n137), .B(n138), .Z(n135) );
  XNOR U227 ( .A(n139), .B(n136), .Z(n138) );
  OR U228 ( .A(n140), .B(n141), .Z(n67) );
  XOR U229 ( .A(n142), .B(n143), .Z(n70) );
  AND U230 ( .A(n144), .B(n145), .Z(n142) );
  XOR U231 ( .A(n146), .B(n143), .Z(n144) );
  XOR U232 ( .A(n147), .B(n148), .Z(n82) );
  ANDN U233 ( .B(n149), .A(n20), .Z(n147) );
  XNOR U234 ( .A(n148), .B(n21), .Z(n149) );
  XNOR U235 ( .A(n116), .B(n118), .Z(n21) );
  XOR U236 ( .A(n110), .B(n112), .Z(n118) );
  XOR U237 ( .A(n94), .B(n95), .Z(n93) );
  AND U238 ( .A(n150), .B(n151), .Z(n95) );
  OR U239 ( .A(n152), .B(n153), .Z(n151) );
  XOR U240 ( .A(n154), .B(n155), .Z(n150) );
  NAND U241 ( .A(n156), .B(n157), .Z(n155) );
  XOR U242 ( .A(n154), .B(n158), .Z(n157) );
  OR U243 ( .A(n159), .B(n160), .Z(n94) );
  XOR U244 ( .A(n92), .B(n161), .Z(n91) );
  XOR U245 ( .A(n86), .B(n87), .Z(n161) );
  AND U246 ( .A(n162), .B(n163), .Z(n87) );
  OR U247 ( .A(n164), .B(n165), .Z(n163) );
  XOR U248 ( .A(n166), .B(n167), .Z(n162) );
  NAND U249 ( .A(n168), .B(n169), .Z(n167) );
  XNOR U250 ( .A(n166), .B(n170), .Z(n168) );
  OR U251 ( .A(n171), .B(n172), .Z(n86) );
  IV U252 ( .A(n89), .Z(n92) );
  XOR U253 ( .A(n173), .B(n174), .Z(n89) );
  NAND U254 ( .A(n175), .B(n176), .Z(n174) );
  XOR U255 ( .A(n173), .B(n177), .Z(n175) );
  XOR U256 ( .A(n103), .B(n178), .Z(n110) );
  XNOR U257 ( .A(n105), .B(n109), .Z(n178) );
  XNOR U258 ( .A(n179), .B(n180), .Z(n109) );
  NAND U259 ( .A(n181), .B(n182), .Z(n180) );
  XNOR U260 ( .A(n179), .B(n183), .Z(n181) );
  XOR U261 ( .A(n106), .B(n107), .Z(n105) );
  AND U262 ( .A(n184), .B(n185), .Z(n107) );
  OR U263 ( .A(n186), .B(n187), .Z(n185) );
  XOR U264 ( .A(n188), .B(n189), .Z(n184) );
  NAND U265 ( .A(n190), .B(n191), .Z(n189) );
  XNOR U266 ( .A(n188), .B(n192), .Z(n190) );
  OR U267 ( .A(n193), .B(n194), .Z(n106) );
  XNOR U268 ( .A(n102), .B(n195), .Z(n103) );
  XOR U269 ( .A(n99), .B(n100), .Z(n195) );
  AND U270 ( .A(n196), .B(n197), .Z(n100) );
  OR U271 ( .A(n198), .B(n199), .Z(n197) );
  XOR U272 ( .A(n200), .B(n201), .Z(n196) );
  NAND U273 ( .A(n202), .B(n203), .Z(n201) );
  XNOR U274 ( .A(n200), .B(n204), .Z(n202) );
  OR U275 ( .A(n205), .B(n206), .Z(n99) );
  XNOR U276 ( .A(n207), .B(n208), .Z(n102) );
  NAND U277 ( .A(n209), .B(n210), .Z(n208) );
  XOR U278 ( .A(n207), .B(n211), .Z(n210) );
  XNOR U279 ( .A(n146), .B(n115), .Z(n212) );
  XNOR U280 ( .A(n213), .B(n214), .Z(n115) );
  NAND U281 ( .A(n215), .B(n216), .Z(n214) );
  XNOR U282 ( .A(n213), .B(n217), .Z(n215) );
  XNOR U283 ( .A(n126), .B(n127), .Z(n146) );
  XNOR U284 ( .A(n128), .B(n129), .Z(n127) );
  AND U285 ( .A(n218), .B(n219), .Z(n129) );
  OR U286 ( .A(n220), .B(n221), .Z(n219) );
  XOR U287 ( .A(n222), .B(n223), .Z(n218) );
  NAND U288 ( .A(n224), .B(n225), .Z(n223) );
  XNOR U289 ( .A(n222), .B(n226), .Z(n224) );
  OR U290 ( .A(n227), .B(n228), .Z(n128) );
  XOR U291 ( .A(n124), .B(n229), .Z(n126) );
  XOR U292 ( .A(n121), .B(n122), .Z(n229) );
  AND U293 ( .A(n230), .B(n231), .Z(n122) );
  OR U294 ( .A(n232), .B(n233), .Z(n231) );
  XOR U295 ( .A(n234), .B(n235), .Z(n230) );
  NAND U296 ( .A(n236), .B(n237), .Z(n235) );
  XNOR U297 ( .A(n234), .B(n238), .Z(n236) );
  OR U298 ( .A(n239), .B(n240), .Z(n121) );
  XNOR U299 ( .A(n241), .B(n242), .Z(n124) );
  NAND U300 ( .A(n243), .B(n244), .Z(n242) );
  XOR U301 ( .A(n241), .B(n245), .Z(n244) );
  XOR U302 ( .A(n137), .B(n246), .Z(n145) );
  XNOR U303 ( .A(n139), .B(n143), .Z(n246) );
  XNOR U304 ( .A(n247), .B(n248), .Z(n143) );
  NAND U305 ( .A(n249), .B(n250), .Z(n248) );
  XOR U306 ( .A(n247), .B(n251), .Z(n250) );
  XOR U307 ( .A(n140), .B(n141), .Z(n139) );
  AND U308 ( .A(n252), .B(n253), .Z(n141) );
  OR U309 ( .A(n254), .B(n255), .Z(n253) );
  XOR U310 ( .A(n256), .B(n257), .Z(n252) );
  NAND U311 ( .A(n258), .B(n259), .Z(n257) );
  XNOR U312 ( .A(n256), .B(n260), .Z(n258) );
  OR U313 ( .A(n261), .B(n262), .Z(n140) );
  XNOR U314 ( .A(n136), .B(n263), .Z(n137) );
  XOR U315 ( .A(n133), .B(n134), .Z(n263) );
  AND U316 ( .A(n264), .B(n265), .Z(n134) );
  OR U317 ( .A(n266), .B(n267), .Z(n265) );
  XOR U318 ( .A(n268), .B(n269), .Z(n264) );
  NAND U319 ( .A(n270), .B(n271), .Z(n269) );
  XNOR U320 ( .A(n268), .B(n272), .Z(n270) );
  OR U321 ( .A(n273), .B(n274), .Z(n133) );
  XNOR U322 ( .A(n275), .B(n276), .Z(n136) );
  NAND U323 ( .A(n277), .B(n278), .Z(n276) );
  XOR U324 ( .A(n275), .B(n279), .Z(n278) );
  XNOR U325 ( .A(n280), .B(n281), .Z(n148) );
  NANDN U326 ( .A(n22), .B(n282), .Z(n281) );
  XNOR U327 ( .A(n280), .B(n23), .Z(n282) );
  XNOR U328 ( .A(n216), .B(n217), .Z(n23) );
  XOR U329 ( .A(n182), .B(n183), .Z(n217) );
  XOR U330 ( .A(n176), .B(n177), .Z(n183) );
  XOR U331 ( .A(n159), .B(n160), .Z(n158) );
  AND U332 ( .A(n283), .B(n284), .Z(n160) );
  OR U333 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U334 ( .A(n287), .B(n288), .Z(n283) );
  OR U335 ( .A(n289), .B(n290), .Z(n159) );
  XOR U336 ( .A(n153), .B(n291), .Z(n156) );
  XOR U337 ( .A(n152), .B(n154), .Z(n291) );
  ANDN U338 ( .B(n292), .A(n293), .Z(n154) );
  OR U339 ( .A(n294), .B(n295), .Z(n152) );
  AND U340 ( .A(n296), .B(n297), .Z(n153) );
  OR U341 ( .A(n298), .B(n299), .Z(n297) );
  OR U342 ( .A(n300), .B(n301), .Z(n296) );
  XOR U343 ( .A(n169), .B(n302), .Z(n176) );
  XNOR U344 ( .A(n173), .B(n170), .Z(n302) );
  XNOR U345 ( .A(n171), .B(n172), .Z(n170) );
  AND U346 ( .A(n303), .B(n304), .Z(n172) );
  OR U347 ( .A(n305), .B(n306), .Z(n304) );
  OR U348 ( .A(n307), .B(n308), .Z(n303) );
  OR U349 ( .A(n309), .B(n310), .Z(n171) );
  ANDN U350 ( .B(n311), .A(n312), .Z(n173) );
  XOR U351 ( .A(n165), .B(n313), .Z(n169) );
  XOR U352 ( .A(n164), .B(n166), .Z(n313) );
  ANDN U353 ( .B(n314), .A(n315), .Z(n166) );
  OR U354 ( .A(n316), .B(n317), .Z(n164) );
  AND U355 ( .A(n318), .B(n319), .Z(n165) );
  OR U356 ( .A(n320), .B(n321), .Z(n319) );
  OR U357 ( .A(n322), .B(n323), .Z(n318) );
  XNOR U358 ( .A(n179), .B(n211), .Z(n324) );
  XOR U359 ( .A(n191), .B(n192), .Z(n211) );
  XNOR U360 ( .A(n193), .B(n194), .Z(n192) );
  AND U361 ( .A(n325), .B(n326), .Z(n194) );
  OR U362 ( .A(n327), .B(n328), .Z(n326) );
  OR U363 ( .A(n329), .B(n330), .Z(n325) );
  OR U364 ( .A(n331), .B(n332), .Z(n193) );
  XOR U365 ( .A(n187), .B(n333), .Z(n191) );
  XOR U366 ( .A(n186), .B(n188), .Z(n333) );
  ANDN U367 ( .B(n334), .A(n335), .Z(n188) );
  OR U368 ( .A(n336), .B(n337), .Z(n186) );
  AND U369 ( .A(n338), .B(n339), .Z(n187) );
  OR U370 ( .A(n340), .B(n341), .Z(n339) );
  OR U371 ( .A(n342), .B(n343), .Z(n338) );
  OR U372 ( .A(n344), .B(n345), .Z(n179) );
  XOR U373 ( .A(n203), .B(n346), .Z(n209) );
  XOR U374 ( .A(n207), .B(n204), .Z(n346) );
  XNOR U375 ( .A(n205), .B(n206), .Z(n204) );
  AND U376 ( .A(n347), .B(n348), .Z(n206) );
  OR U377 ( .A(n349), .B(n350), .Z(n348) );
  OR U378 ( .A(n351), .B(n352), .Z(n347) );
  OR U379 ( .A(n353), .B(n354), .Z(n205) );
  OR U380 ( .A(n355), .B(n356), .Z(n207) );
  XOR U381 ( .A(n199), .B(n357), .Z(n203) );
  XOR U382 ( .A(n198), .B(n200), .Z(n357) );
  ANDN U383 ( .B(n358), .A(n359), .Z(n200) );
  OR U384 ( .A(n360), .B(n361), .Z(n198) );
  AND U385 ( .A(n362), .B(n363), .Z(n199) );
  OR U386 ( .A(n364), .B(n365), .Z(n363) );
  OR U387 ( .A(n366), .B(n367), .Z(n362) );
  XNOR U388 ( .A(n213), .B(n251), .Z(n368) );
  XOR U389 ( .A(n225), .B(n226), .Z(n245) );
  XNOR U390 ( .A(n227), .B(n228), .Z(n226) );
  AND U391 ( .A(n369), .B(n370), .Z(n228) );
  OR U392 ( .A(n371), .B(n372), .Z(n370) );
  OR U393 ( .A(n373), .B(n374), .Z(n369) );
  OR U394 ( .A(n375), .B(n376), .Z(n227) );
  XOR U395 ( .A(n221), .B(n377), .Z(n225) );
  XOR U396 ( .A(n220), .B(n222), .Z(n377) );
  ANDN U397 ( .B(n378), .A(n379), .Z(n222) );
  OR U398 ( .A(n380), .B(n381), .Z(n220) );
  AND U399 ( .A(n382), .B(n383), .Z(n221) );
  OR U400 ( .A(n384), .B(n385), .Z(n383) );
  OR U401 ( .A(n386), .B(n387), .Z(n382) );
  XOR U402 ( .A(n237), .B(n388), .Z(n243) );
  XOR U403 ( .A(n241), .B(n238), .Z(n388) );
  XNOR U404 ( .A(n239), .B(n240), .Z(n238) );
  AND U405 ( .A(n389), .B(n390), .Z(n240) );
  OR U406 ( .A(n391), .B(n392), .Z(n390) );
  OR U407 ( .A(n393), .B(n394), .Z(n389) );
  OR U408 ( .A(n395), .B(n396), .Z(n239) );
  OR U409 ( .A(n397), .B(n398), .Z(n241) );
  XOR U410 ( .A(n233), .B(n399), .Z(n237) );
  XOR U411 ( .A(n232), .B(n234), .Z(n399) );
  ANDN U412 ( .B(n400), .A(n401), .Z(n234) );
  OR U413 ( .A(n402), .B(n403), .Z(n232) );
  AND U414 ( .A(n404), .B(n405), .Z(n233) );
  OR U415 ( .A(n406), .B(n407), .Z(n405) );
  OR U416 ( .A(n408), .B(n409), .Z(n404) );
  OR U417 ( .A(n410), .B(n411), .Z(n213) );
  XNOR U418 ( .A(n247), .B(n279), .Z(n412) );
  XOR U419 ( .A(n259), .B(n260), .Z(n279) );
  XNOR U420 ( .A(n261), .B(n262), .Z(n260) );
  AND U421 ( .A(n413), .B(n414), .Z(n262) );
  OR U422 ( .A(n415), .B(n416), .Z(n414) );
  OR U423 ( .A(n417), .B(n418), .Z(n413) );
  OR U424 ( .A(n419), .B(n420), .Z(n261) );
  XOR U425 ( .A(n255), .B(n421), .Z(n259) );
  XOR U426 ( .A(n254), .B(n256), .Z(n421) );
  ANDN U427 ( .B(n422), .A(n423), .Z(n256) );
  OR U428 ( .A(n424), .B(n425), .Z(n254) );
  AND U429 ( .A(n426), .B(n427), .Z(n255) );
  OR U430 ( .A(n428), .B(n429), .Z(n427) );
  OR U431 ( .A(n430), .B(n431), .Z(n426) );
  OR U432 ( .A(n432), .B(n433), .Z(n247) );
  XOR U433 ( .A(n271), .B(n434), .Z(n277) );
  XOR U434 ( .A(n275), .B(n272), .Z(n434) );
  XNOR U435 ( .A(n273), .B(n274), .Z(n272) );
  AND U436 ( .A(n435), .B(n436), .Z(n274) );
  OR U437 ( .A(n437), .B(n438), .Z(n436) );
  OR U438 ( .A(n439), .B(n440), .Z(n435) );
  OR U439 ( .A(n441), .B(n442), .Z(n273) );
  OR U440 ( .A(n443), .B(n444), .Z(n275) );
  XOR U441 ( .A(n267), .B(n445), .Z(n271) );
  XOR U442 ( .A(n266), .B(n268), .Z(n445) );
  ANDN U443 ( .B(n446), .A(n447), .Z(n268) );
  OR U444 ( .A(n448), .B(n449), .Z(n266) );
  AND U445 ( .A(n450), .B(n451), .Z(n267) );
  OR U446 ( .A(n452), .B(n453), .Z(n451) );
  OR U447 ( .A(n454), .B(n455), .Z(n450) );
  XNOR U448 ( .A(oglobal[1]), .B(n280), .Z(n22) );
  ANDN U449 ( .B(oglobal[0]), .A(n456), .Z(n280) );
  XNOR U450 ( .A(oglobal[0]), .B(n456), .Z(o[0]) );
  XNOR U451 ( .A(n411), .B(n410), .Z(n456) );
  XNOR U452 ( .A(n345), .B(n344), .Z(n410) );
  XNOR U453 ( .A(n292), .B(n293), .Z(n311) );
  XOR U454 ( .A(n287), .B(n288), .Z(n293) );
  XOR U455 ( .A(n289), .B(n290), .Z(n288) );
  XNOR U456 ( .A(y[63]), .B(x[63]), .Z(n290) );
  XNOR U457 ( .A(y[62]), .B(x[62]), .Z(n289) );
  XNOR U458 ( .A(n285), .B(n286), .Z(n287) );
  XNOR U459 ( .A(y[61]), .B(x[61]), .Z(n286) );
  XNOR U460 ( .A(y[60]), .B(x[60]), .Z(n285) );
  XOR U461 ( .A(n300), .B(n301), .Z(n292) );
  XNOR U462 ( .A(n295), .B(n294), .Z(n301) );
  XNOR U463 ( .A(y[59]), .B(x[59]), .Z(n294) );
  XNOR U464 ( .A(y[58]), .B(x[58]), .Z(n295) );
  XNOR U465 ( .A(n298), .B(n299), .Z(n300) );
  XNOR U466 ( .A(y[57]), .B(x[57]), .Z(n299) );
  XNOR U467 ( .A(y[56]), .B(x[56]), .Z(n298) );
  XOR U468 ( .A(n307), .B(n308), .Z(n314) );
  XNOR U469 ( .A(n310), .B(n309), .Z(n308) );
  XNOR U470 ( .A(y[55]), .B(x[55]), .Z(n309) );
  XNOR U471 ( .A(y[54]), .B(x[54]), .Z(n310) );
  XNOR U472 ( .A(n305), .B(n306), .Z(n307) );
  XNOR U473 ( .A(y[53]), .B(x[53]), .Z(n306) );
  XNOR U474 ( .A(y[52]), .B(x[52]), .Z(n305) );
  XNOR U475 ( .A(n322), .B(n323), .Z(n315) );
  XNOR U476 ( .A(n317), .B(n316), .Z(n323) );
  XNOR U477 ( .A(y[51]), .B(x[51]), .Z(n316) );
  XNOR U478 ( .A(y[50]), .B(x[50]), .Z(n317) );
  XNOR U479 ( .A(n320), .B(n321), .Z(n322) );
  XNOR U480 ( .A(y[49]), .B(x[49]), .Z(n321) );
  XNOR U481 ( .A(y[48]), .B(x[48]), .Z(n320) );
  XNOR U482 ( .A(n356), .B(n355), .Z(n345) );
  XOR U483 ( .A(n329), .B(n330), .Z(n334) );
  XNOR U484 ( .A(n332), .B(n331), .Z(n330) );
  XNOR U485 ( .A(y[47]), .B(x[47]), .Z(n331) );
  XNOR U486 ( .A(y[46]), .B(x[46]), .Z(n332) );
  XNOR U487 ( .A(n327), .B(n328), .Z(n329) );
  XNOR U488 ( .A(y[45]), .B(x[45]), .Z(n328) );
  XNOR U489 ( .A(y[44]), .B(x[44]), .Z(n327) );
  XNOR U490 ( .A(n342), .B(n343), .Z(n335) );
  XNOR U491 ( .A(n337), .B(n336), .Z(n343) );
  XNOR U492 ( .A(y[43]), .B(x[43]), .Z(n336) );
  XNOR U493 ( .A(y[42]), .B(x[42]), .Z(n337) );
  XNOR U494 ( .A(n340), .B(n341), .Z(n342) );
  XNOR U495 ( .A(y[41]), .B(x[41]), .Z(n341) );
  XNOR U496 ( .A(y[40]), .B(x[40]), .Z(n340) );
  XOR U497 ( .A(n351), .B(n352), .Z(n358) );
  XNOR U498 ( .A(n354), .B(n353), .Z(n352) );
  XNOR U499 ( .A(y[39]), .B(x[39]), .Z(n353) );
  XNOR U500 ( .A(y[38]), .B(x[38]), .Z(n354) );
  XNOR U501 ( .A(n349), .B(n350), .Z(n351) );
  XNOR U502 ( .A(y[37]), .B(x[37]), .Z(n350) );
  XNOR U503 ( .A(y[36]), .B(x[36]), .Z(n349) );
  XNOR U504 ( .A(n366), .B(n367), .Z(n359) );
  XNOR U505 ( .A(n361), .B(n360), .Z(n367) );
  XNOR U506 ( .A(y[35]), .B(x[35]), .Z(n360) );
  XNOR U507 ( .A(y[34]), .B(x[34]), .Z(n361) );
  XNOR U508 ( .A(n364), .B(n365), .Z(n366) );
  XNOR U509 ( .A(y[33]), .B(x[33]), .Z(n365) );
  XNOR U510 ( .A(y[32]), .B(x[32]), .Z(n364) );
  XNOR U511 ( .A(n433), .B(n432), .Z(n411) );
  XNOR U512 ( .A(n398), .B(n397), .Z(n432) );
  XOR U513 ( .A(n373), .B(n374), .Z(n378) );
  XNOR U514 ( .A(n376), .B(n375), .Z(n374) );
  XNOR U515 ( .A(y[31]), .B(x[31]), .Z(n375) );
  XNOR U516 ( .A(y[30]), .B(x[30]), .Z(n376) );
  XNOR U517 ( .A(n371), .B(n372), .Z(n373) );
  XNOR U518 ( .A(y[29]), .B(x[29]), .Z(n372) );
  XNOR U519 ( .A(y[28]), .B(x[28]), .Z(n371) );
  XNOR U520 ( .A(n386), .B(n387), .Z(n379) );
  XNOR U521 ( .A(n381), .B(n380), .Z(n387) );
  XNOR U522 ( .A(y[27]), .B(x[27]), .Z(n380) );
  XNOR U523 ( .A(y[26]), .B(x[26]), .Z(n381) );
  XNOR U524 ( .A(n384), .B(n385), .Z(n386) );
  XNOR U525 ( .A(y[25]), .B(x[25]), .Z(n385) );
  XNOR U526 ( .A(y[24]), .B(x[24]), .Z(n384) );
  XOR U527 ( .A(n393), .B(n394), .Z(n400) );
  XNOR U528 ( .A(n396), .B(n395), .Z(n394) );
  XNOR U529 ( .A(y[23]), .B(x[23]), .Z(n395) );
  XNOR U530 ( .A(y[22]), .B(x[22]), .Z(n396) );
  XNOR U531 ( .A(n391), .B(n392), .Z(n393) );
  XNOR U532 ( .A(y[21]), .B(x[21]), .Z(n392) );
  XNOR U533 ( .A(y[20]), .B(x[20]), .Z(n391) );
  XNOR U534 ( .A(n408), .B(n409), .Z(n401) );
  XNOR U535 ( .A(n403), .B(n402), .Z(n409) );
  XNOR U536 ( .A(y[19]), .B(x[19]), .Z(n402) );
  XNOR U537 ( .A(y[18]), .B(x[18]), .Z(n403) );
  XNOR U538 ( .A(n406), .B(n407), .Z(n408) );
  XNOR U539 ( .A(y[17]), .B(x[17]), .Z(n407) );
  XNOR U540 ( .A(y[16]), .B(x[16]), .Z(n406) );
  XNOR U541 ( .A(n444), .B(n443), .Z(n433) );
  XOR U542 ( .A(n417), .B(n418), .Z(n422) );
  XNOR U543 ( .A(n420), .B(n419), .Z(n418) );
  XNOR U544 ( .A(y[15]), .B(x[15]), .Z(n419) );
  XNOR U545 ( .A(y[14]), .B(x[14]), .Z(n420) );
  XNOR U546 ( .A(n415), .B(n416), .Z(n417) );
  XNOR U547 ( .A(y[13]), .B(x[13]), .Z(n416) );
  XNOR U548 ( .A(y[12]), .B(x[12]), .Z(n415) );
  XNOR U549 ( .A(n430), .B(n431), .Z(n423) );
  XNOR U550 ( .A(n425), .B(n424), .Z(n431) );
  XNOR U551 ( .A(y[11]), .B(x[11]), .Z(n424) );
  XNOR U552 ( .A(y[10]), .B(x[10]), .Z(n425) );
  XNOR U553 ( .A(n428), .B(n429), .Z(n430) );
  XNOR U554 ( .A(y[9]), .B(x[9]), .Z(n429) );
  XNOR U555 ( .A(y[8]), .B(x[8]), .Z(n428) );
  XOR U556 ( .A(n439), .B(n440), .Z(n446) );
  XNOR U557 ( .A(n442), .B(n441), .Z(n440) );
  XNOR U558 ( .A(y[7]), .B(x[7]), .Z(n441) );
  XNOR U559 ( .A(y[6]), .B(x[6]), .Z(n442) );
  XNOR U560 ( .A(n437), .B(n438), .Z(n439) );
  XNOR U561 ( .A(y[5]), .B(x[5]), .Z(n438) );
  XNOR U562 ( .A(y[4]), .B(x[4]), .Z(n437) );
  XNOR U563 ( .A(n454), .B(n455), .Z(n447) );
  XNOR U564 ( .A(n449), .B(n448), .Z(n455) );
  XNOR U565 ( .A(y[3]), .B(x[3]), .Z(n448) );
  XNOR U566 ( .A(y[2]), .B(x[2]), .Z(n449) );
  XNOR U567 ( .A(n452), .B(n453), .Z(n454) );
  XNOR U568 ( .A(y[1]), .B(x[1]), .Z(n453) );
  XNOR U569 ( .A(y[0]), .B(x[0]), .Z(n452) );
endmodule

