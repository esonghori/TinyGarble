
module hamming_N16000_CC2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U18 ( .A(B[1]), .B(A[1]), .Z(n18) );
  XOR U19 ( .A(A[13]), .B(n19), .Z(SUM[13]) );
  NAND U20 ( .A(n20), .B(n21), .Z(n19) );
  NAND U21 ( .A(n22), .B(B[12]), .Z(n21) );
  NANDN U22 ( .A(A[12]), .B(n23), .Z(n22) );
  NANDN U23 ( .A(n23), .B(A[12]), .Z(n20) );
  XOR U24 ( .A(n23), .B(n24), .Z(SUM[12]) );
  XNOR U25 ( .A(B[12]), .B(A[12]), .Z(n24) );
  AND U26 ( .A(n25), .B(n26), .Z(n23) );
  NAND U27 ( .A(n27), .B(B[11]), .Z(n26) );
  NANDN U28 ( .A(A[11]), .B(n28), .Z(n27) );
  NANDN U29 ( .A(n28), .B(A[11]), .Z(n25) );
  XOR U30 ( .A(n28), .B(n29), .Z(SUM[11]) );
  XNOR U31 ( .A(B[11]), .B(A[11]), .Z(n29) );
  AND U32 ( .A(n30), .B(n31), .Z(n28) );
  NAND U33 ( .A(n32), .B(B[10]), .Z(n31) );
  NANDN U34 ( .A(A[10]), .B(n33), .Z(n32) );
  NANDN U35 ( .A(n33), .B(A[10]), .Z(n30) );
  XOR U36 ( .A(n33), .B(n34), .Z(SUM[10]) );
  XNOR U37 ( .A(B[10]), .B(A[10]), .Z(n34) );
  AND U38 ( .A(n35), .B(n36), .Z(n33) );
  NAND U39 ( .A(n37), .B(B[9]), .Z(n36) );
  NANDN U40 ( .A(A[9]), .B(n1), .Z(n37) );
  NANDN U41 ( .A(n1), .B(A[9]), .Z(n35) );
  AND U42 ( .A(n38), .B(n39), .Z(n1) );
  NAND U43 ( .A(n40), .B(B[8]), .Z(n39) );
  NANDN U44 ( .A(A[8]), .B(n3), .Z(n40) );
  NANDN U45 ( .A(n3), .B(A[8]), .Z(n38) );
  AND U46 ( .A(n41), .B(n42), .Z(n3) );
  NAND U47 ( .A(n43), .B(B[7]), .Z(n42) );
  NANDN U48 ( .A(A[7]), .B(n5), .Z(n43) );
  NANDN U49 ( .A(n5), .B(A[7]), .Z(n41) );
  AND U50 ( .A(n44), .B(n45), .Z(n5) );
  NAND U51 ( .A(n46), .B(B[6]), .Z(n45) );
  NANDN U52 ( .A(A[6]), .B(n7), .Z(n46) );
  NANDN U53 ( .A(n7), .B(A[6]), .Z(n44) );
  AND U54 ( .A(n47), .B(n48), .Z(n7) );
  NAND U55 ( .A(n49), .B(B[5]), .Z(n48) );
  NANDN U56 ( .A(A[5]), .B(n9), .Z(n49) );
  NANDN U57 ( .A(n9), .B(A[5]), .Z(n47) );
  AND U58 ( .A(n50), .B(n51), .Z(n9) );
  NAND U59 ( .A(n52), .B(B[4]), .Z(n51) );
  NANDN U60 ( .A(A[4]), .B(n11), .Z(n52) );
  NANDN U61 ( .A(n11), .B(A[4]), .Z(n50) );
  AND U62 ( .A(n53), .B(n54), .Z(n11) );
  NAND U63 ( .A(n55), .B(B[3]), .Z(n54) );
  NANDN U64 ( .A(A[3]), .B(n13), .Z(n55) );
  NANDN U65 ( .A(n13), .B(A[3]), .Z(n53) );
  AND U66 ( .A(n56), .B(n57), .Z(n13) );
  NAND U67 ( .A(n58), .B(B[2]), .Z(n57) );
  NANDN U68 ( .A(A[2]), .B(n15), .Z(n58) );
  NANDN U69 ( .A(n15), .B(A[2]), .Z(n56) );
  AND U70 ( .A(n59), .B(n60), .Z(n15) );
  NAND U71 ( .A(n61), .B(B[1]), .Z(n60) );
  OR U72 ( .A(n17), .B(A[1]), .Z(n61) );
  NAND U73 ( .A(n17), .B(A[1]), .Z(n59) );
  AND U74 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U75 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;

  IV U1 ( .A(B[12]), .Z(n1) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  XOR U20 ( .A(n20), .B(n1), .Z(SUM[12]) );
  AND U21 ( .A(n21), .B(n22), .Z(n20) );
  NAND U22 ( .A(n23), .B(B[11]), .Z(n22) );
  NANDN U23 ( .A(A[11]), .B(n24), .Z(n23) );
  NANDN U24 ( .A(n24), .B(A[11]), .Z(n21) );
  XOR U25 ( .A(n24), .B(n25), .Z(SUM[11]) );
  XNOR U26 ( .A(B[11]), .B(A[11]), .Z(n25) );
  AND U27 ( .A(n26), .B(n27), .Z(n24) );
  NAND U28 ( .A(n28), .B(B[10]), .Z(n27) );
  NANDN U29 ( .A(A[10]), .B(n29), .Z(n28) );
  NANDN U30 ( .A(n29), .B(A[10]), .Z(n26) );
  XOR U31 ( .A(n29), .B(n30), .Z(SUM[10]) );
  XNOR U32 ( .A(B[10]), .B(A[10]), .Z(n30) );
  AND U33 ( .A(n31), .B(n32), .Z(n29) );
  NAND U34 ( .A(n33), .B(B[9]), .Z(n32) );
  NANDN U35 ( .A(A[9]), .B(n2), .Z(n33) );
  NANDN U36 ( .A(n2), .B(A[9]), .Z(n31) );
  AND U37 ( .A(n34), .B(n35), .Z(n2) );
  NAND U38 ( .A(n36), .B(B[8]), .Z(n35) );
  NANDN U39 ( .A(A[8]), .B(n4), .Z(n36) );
  NANDN U40 ( .A(n4), .B(A[8]), .Z(n34) );
  AND U41 ( .A(n37), .B(n38), .Z(n4) );
  NAND U42 ( .A(n39), .B(B[7]), .Z(n38) );
  NANDN U43 ( .A(A[7]), .B(n6), .Z(n39) );
  NANDN U44 ( .A(n6), .B(A[7]), .Z(n37) );
  AND U45 ( .A(n40), .B(n41), .Z(n6) );
  NAND U46 ( .A(n42), .B(B[6]), .Z(n41) );
  NANDN U47 ( .A(A[6]), .B(n8), .Z(n42) );
  NANDN U48 ( .A(n8), .B(A[6]), .Z(n40) );
  AND U49 ( .A(n43), .B(n44), .Z(n8) );
  NAND U50 ( .A(n45), .B(B[5]), .Z(n44) );
  NANDN U51 ( .A(A[5]), .B(n10), .Z(n45) );
  NANDN U52 ( .A(n10), .B(A[5]), .Z(n43) );
  AND U53 ( .A(n46), .B(n47), .Z(n10) );
  NAND U54 ( .A(n48), .B(B[4]), .Z(n47) );
  NANDN U55 ( .A(A[4]), .B(n12), .Z(n48) );
  NANDN U56 ( .A(n12), .B(A[4]), .Z(n46) );
  AND U57 ( .A(n49), .B(n50), .Z(n12) );
  NAND U58 ( .A(n51), .B(B[3]), .Z(n50) );
  NANDN U59 ( .A(A[3]), .B(n14), .Z(n51) );
  NANDN U60 ( .A(n14), .B(A[3]), .Z(n49) );
  AND U61 ( .A(n52), .B(n53), .Z(n14) );
  NAND U62 ( .A(n54), .B(B[2]), .Z(n53) );
  NANDN U63 ( .A(A[2]), .B(n16), .Z(n54) );
  NANDN U64 ( .A(n16), .B(A[2]), .Z(n52) );
  AND U65 ( .A(n55), .B(n56), .Z(n16) );
  NAND U66 ( .A(n57), .B(B[1]), .Z(n56) );
  OR U67 ( .A(n18), .B(A[1]), .Z(n57) );
  NAND U68 ( .A(n18), .B(A[1]), .Z(n55) );
  AND U69 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U70 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_2 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[12]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[11]), .Z(n21) );
  NANDN U21 ( .A(A[11]), .B(n23), .Z(n22) );
  NANDN U22 ( .A(n23), .B(A[11]), .Z(n20) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[11]) );
  XNOR U24 ( .A(B[11]), .B(A[11]), .Z(n24) );
  AND U25 ( .A(n25), .B(n26), .Z(n23) );
  NAND U26 ( .A(n27), .B(B[10]), .Z(n26) );
  NANDN U27 ( .A(A[10]), .B(n28), .Z(n27) );
  NANDN U28 ( .A(n28), .B(A[10]), .Z(n25) );
  XOR U29 ( .A(n28), .B(n29), .Z(SUM[10]) );
  XNOR U30 ( .A(B[10]), .B(A[10]), .Z(n29) );
  AND U31 ( .A(n30), .B(n31), .Z(n28) );
  NAND U32 ( .A(n32), .B(B[9]), .Z(n31) );
  NANDN U33 ( .A(A[9]), .B(n2), .Z(n32) );
  NANDN U34 ( .A(n2), .B(A[9]), .Z(n30) );
  AND U35 ( .A(n33), .B(n34), .Z(n2) );
  NAND U36 ( .A(n35), .B(B[8]), .Z(n34) );
  NANDN U37 ( .A(A[8]), .B(n4), .Z(n35) );
  NANDN U38 ( .A(n4), .B(A[8]), .Z(n33) );
  AND U39 ( .A(n36), .B(n37), .Z(n4) );
  NAND U40 ( .A(n38), .B(B[7]), .Z(n37) );
  NANDN U41 ( .A(A[7]), .B(n6), .Z(n38) );
  NANDN U42 ( .A(n6), .B(A[7]), .Z(n36) );
  AND U43 ( .A(n39), .B(n40), .Z(n6) );
  NAND U44 ( .A(n41), .B(B[6]), .Z(n40) );
  NANDN U45 ( .A(A[6]), .B(n8), .Z(n41) );
  NANDN U46 ( .A(n8), .B(A[6]), .Z(n39) );
  AND U47 ( .A(n42), .B(n43), .Z(n8) );
  NAND U48 ( .A(n44), .B(B[5]), .Z(n43) );
  NANDN U49 ( .A(A[5]), .B(n10), .Z(n44) );
  NANDN U50 ( .A(n10), .B(A[5]), .Z(n42) );
  AND U51 ( .A(n45), .B(n46), .Z(n10) );
  NAND U52 ( .A(n47), .B(B[4]), .Z(n46) );
  NANDN U53 ( .A(A[4]), .B(n12), .Z(n47) );
  NANDN U54 ( .A(n12), .B(A[4]), .Z(n45) );
  AND U55 ( .A(n48), .B(n49), .Z(n12) );
  NAND U56 ( .A(n50), .B(B[3]), .Z(n49) );
  NANDN U57 ( .A(A[3]), .B(n14), .Z(n50) );
  NANDN U58 ( .A(n14), .B(A[3]), .Z(n48) );
  AND U59 ( .A(n51), .B(n52), .Z(n14) );
  NAND U60 ( .A(n53), .B(B[2]), .Z(n52) );
  NANDN U61 ( .A(A[2]), .B(n16), .Z(n53) );
  NANDN U62 ( .A(n16), .B(A[2]), .Z(n51) );
  AND U63 ( .A(n54), .B(n55), .Z(n16) );
  NAND U64 ( .A(n56), .B(B[1]), .Z(n55) );
  OR U65 ( .A(n18), .B(A[1]), .Z(n56) );
  NAND U66 ( .A(n18), .B(A[1]), .Z(n54) );
  AND U67 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U68 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_3 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[11]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[10]), .Z(n21) );
  NANDN U21 ( .A(A[10]), .B(n23), .Z(n22) );
  NANDN U22 ( .A(n23), .B(A[10]), .Z(n20) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[10]) );
  XNOR U24 ( .A(B[10]), .B(A[10]), .Z(n24) );
  AND U25 ( .A(n25), .B(n26), .Z(n23) );
  NAND U26 ( .A(n27), .B(B[9]), .Z(n26) );
  NANDN U27 ( .A(A[9]), .B(n2), .Z(n27) );
  NANDN U28 ( .A(n2), .B(A[9]), .Z(n25) );
  AND U29 ( .A(n28), .B(n29), .Z(n2) );
  NAND U30 ( .A(n30), .B(B[8]), .Z(n29) );
  NANDN U31 ( .A(A[8]), .B(n4), .Z(n30) );
  NANDN U32 ( .A(n4), .B(A[8]), .Z(n28) );
  AND U33 ( .A(n31), .B(n32), .Z(n4) );
  NAND U34 ( .A(n33), .B(B[7]), .Z(n32) );
  NANDN U35 ( .A(A[7]), .B(n6), .Z(n33) );
  NANDN U36 ( .A(n6), .B(A[7]), .Z(n31) );
  AND U37 ( .A(n34), .B(n35), .Z(n6) );
  NAND U38 ( .A(n36), .B(B[6]), .Z(n35) );
  NANDN U39 ( .A(A[6]), .B(n8), .Z(n36) );
  NANDN U40 ( .A(n8), .B(A[6]), .Z(n34) );
  AND U41 ( .A(n37), .B(n38), .Z(n8) );
  NAND U42 ( .A(n39), .B(B[5]), .Z(n38) );
  NANDN U43 ( .A(A[5]), .B(n10), .Z(n39) );
  NANDN U44 ( .A(n10), .B(A[5]), .Z(n37) );
  AND U45 ( .A(n40), .B(n41), .Z(n10) );
  NAND U46 ( .A(n42), .B(B[4]), .Z(n41) );
  NANDN U47 ( .A(A[4]), .B(n12), .Z(n42) );
  NANDN U48 ( .A(n12), .B(A[4]), .Z(n40) );
  AND U49 ( .A(n43), .B(n44), .Z(n12) );
  NAND U50 ( .A(n45), .B(B[3]), .Z(n44) );
  NANDN U51 ( .A(A[3]), .B(n14), .Z(n45) );
  NANDN U52 ( .A(n14), .B(A[3]), .Z(n43) );
  AND U53 ( .A(n46), .B(n47), .Z(n14) );
  NAND U54 ( .A(n48), .B(B[2]), .Z(n47) );
  NANDN U55 ( .A(A[2]), .B(n16), .Z(n48) );
  NANDN U56 ( .A(n16), .B(A[2]), .Z(n46) );
  AND U57 ( .A(n49), .B(n50), .Z(n16) );
  NAND U58 ( .A(n51), .B(B[1]), .Z(n50) );
  OR U59 ( .A(n18), .B(A[1]), .Z(n51) );
  NAND U60 ( .A(n18), .B(A[1]), .Z(n49) );
  AND U61 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U62 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_4 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[11]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[10]), .Z(n21) );
  NANDN U21 ( .A(A[10]), .B(n23), .Z(n22) );
  NANDN U22 ( .A(n23), .B(A[10]), .Z(n20) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[10]) );
  XNOR U24 ( .A(B[10]), .B(A[10]), .Z(n24) );
  AND U25 ( .A(n25), .B(n26), .Z(n23) );
  NAND U26 ( .A(n27), .B(B[9]), .Z(n26) );
  NANDN U27 ( .A(A[9]), .B(n2), .Z(n27) );
  NANDN U28 ( .A(n2), .B(A[9]), .Z(n25) );
  AND U29 ( .A(n28), .B(n29), .Z(n2) );
  NAND U30 ( .A(n30), .B(B[8]), .Z(n29) );
  NANDN U31 ( .A(A[8]), .B(n4), .Z(n30) );
  NANDN U32 ( .A(n4), .B(A[8]), .Z(n28) );
  AND U33 ( .A(n31), .B(n32), .Z(n4) );
  NAND U34 ( .A(n33), .B(B[7]), .Z(n32) );
  NANDN U35 ( .A(A[7]), .B(n6), .Z(n33) );
  NANDN U36 ( .A(n6), .B(A[7]), .Z(n31) );
  AND U37 ( .A(n34), .B(n35), .Z(n6) );
  NAND U38 ( .A(n36), .B(B[6]), .Z(n35) );
  NANDN U39 ( .A(A[6]), .B(n8), .Z(n36) );
  NANDN U40 ( .A(n8), .B(A[6]), .Z(n34) );
  AND U41 ( .A(n37), .B(n38), .Z(n8) );
  NAND U42 ( .A(n39), .B(B[5]), .Z(n38) );
  NANDN U43 ( .A(A[5]), .B(n10), .Z(n39) );
  NANDN U44 ( .A(n10), .B(A[5]), .Z(n37) );
  AND U45 ( .A(n40), .B(n41), .Z(n10) );
  NAND U46 ( .A(n42), .B(B[4]), .Z(n41) );
  NANDN U47 ( .A(A[4]), .B(n12), .Z(n42) );
  NANDN U48 ( .A(n12), .B(A[4]), .Z(n40) );
  AND U49 ( .A(n43), .B(n44), .Z(n12) );
  NAND U50 ( .A(n45), .B(B[3]), .Z(n44) );
  NANDN U51 ( .A(A[3]), .B(n14), .Z(n45) );
  NANDN U52 ( .A(n14), .B(A[3]), .Z(n43) );
  AND U53 ( .A(n46), .B(n47), .Z(n14) );
  NAND U54 ( .A(n48), .B(B[2]), .Z(n47) );
  NANDN U55 ( .A(A[2]), .B(n16), .Z(n48) );
  NANDN U56 ( .A(n16), .B(A[2]), .Z(n46) );
  AND U57 ( .A(n49), .B(n50), .Z(n16) );
  NAND U58 ( .A(n51), .B(B[1]), .Z(n50) );
  OR U59 ( .A(n18), .B(A[1]), .Z(n51) );
  NAND U60 ( .A(n18), .B(A[1]), .Z(n49) );
  AND U61 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U62 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_5 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49;

  AND U1 ( .A(n2), .B(B[10]), .Z(SUM[11]) );
  IV U2 ( .A(n22), .Z(n2) );
  IV U3 ( .A(B[10]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[9]) );
  XNOR U5 ( .A(B[9]), .B(A[9]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[8]) );
  XNOR U7 ( .A(B[8]), .B(A[8]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[7]) );
  XNOR U9 ( .A(B[7]), .B(A[7]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[6]) );
  XNOR U11 ( .A(B[6]), .B(A[6]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[5]) );
  XNOR U13 ( .A(B[5]), .B(A[5]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[4]) );
  XNOR U15 ( .A(B[4]), .B(A[4]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[3]) );
  XNOR U17 ( .A(B[3]), .B(A[3]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[2]) );
  XNOR U19 ( .A(B[2]), .B(A[2]), .Z(n19) );
  XOR U20 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U21 ( .A(B[1]), .B(A[1]), .Z(n21) );
  XOR U22 ( .A(n22), .B(n3), .Z(SUM[10]) );
  AND U23 ( .A(n23), .B(n24), .Z(n22) );
  NAND U24 ( .A(n25), .B(B[9]), .Z(n24) );
  NANDN U25 ( .A(A[9]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[9]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(n28), .B(B[8]), .Z(n27) );
  NANDN U29 ( .A(A[8]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[8]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(n31), .B(B[7]), .Z(n30) );
  NANDN U33 ( .A(A[7]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[7]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(n34), .B(B[6]), .Z(n33) );
  NANDN U37 ( .A(A[6]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[6]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(n37), .B(B[5]), .Z(n36) );
  NANDN U41 ( .A(A[5]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[5]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(n40), .B(B[4]), .Z(n39) );
  NANDN U45 ( .A(A[4]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[4]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(n43), .B(B[3]), .Z(n42) );
  NANDN U49 ( .A(A[3]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[3]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(n46), .B(B[2]), .Z(n45) );
  NANDN U53 ( .A(A[2]), .B(n18), .Z(n46) );
  NANDN U54 ( .A(n18), .B(A[2]), .Z(n44) );
  AND U55 ( .A(n47), .B(n48), .Z(n18) );
  NAND U56 ( .A(n49), .B(B[1]), .Z(n48) );
  OR U57 ( .A(n20), .B(A[1]), .Z(n49) );
  NAND U58 ( .A(n20), .B(A[1]), .Z(n47) );
  AND U59 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U60 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_6 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[9]), .Z(n21) );
  NANDN U21 ( .A(A[9]), .B(n2), .Z(n22) );
  NANDN U22 ( .A(n2), .B(A[9]), .Z(n20) );
  AND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(n25), .B(B[8]), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(n28), .B(B[7]), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(n31), .B(B[6]), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(n34), .B(B[5]), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(n37), .B(B[4]), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(n40), .B(B[3]), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(n43), .B(B[2]), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(n46), .B(B[1]), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(n18), .B(A[1]), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_7 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[9]), .Z(n21) );
  NANDN U21 ( .A(A[9]), .B(n2), .Z(n22) );
  NANDN U22 ( .A(n2), .B(A[9]), .Z(n20) );
  AND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(n25), .B(B[8]), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(n28), .B(B[7]), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(n31), .B(B[6]), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(n34), .B(B[5]), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(n37), .B(B[4]), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(n40), .B(B[3]), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(n43), .B(B[2]), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(n46), .B(B[1]), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(n18), .B(A[1]), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_8 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[9]), .Z(n21) );
  NANDN U21 ( .A(A[9]), .B(n2), .Z(n22) );
  NANDN U22 ( .A(n2), .B(A[9]), .Z(n20) );
  AND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(n25), .B(B[8]), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(n28), .B(B[7]), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(n31), .B(B[6]), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(n34), .B(B[5]), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(n37), .B(B[4]), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(n40), .B(B[3]), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(n43), .B(B[2]), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(n46), .B(B[1]), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(n18), .B(A[1]), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_9 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[9]), .Z(n21) );
  NANDN U21 ( .A(A[9]), .B(n2), .Z(n22) );
  NANDN U22 ( .A(n2), .B(A[9]), .Z(n20) );
  AND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(n25), .B(B[8]), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(n28), .B(B[7]), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(n31), .B(B[6]), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(n34), .B(B[5]), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(n37), .B(B[4]), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(n40), .B(B[3]), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(n43), .B(B[2]), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(n46), .B(B[1]), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(n18), .B(A[1]), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_10 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  AND U1 ( .A(n2), .B(B[9]), .Z(SUM[10]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[9]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[8]) );
  XNOR U6 ( .A(B[8]), .B(A[8]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[7]) );
  XNOR U8 ( .A(B[7]), .B(A[7]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[6]) );
  XNOR U10 ( .A(B[6]), .B(A[6]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[5]) );
  XNOR U12 ( .A(B[5]), .B(A[5]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[4]) );
  XNOR U14 ( .A(B[4]), .B(A[4]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U16 ( .A(B[3]), .B(A[3]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(SUM[1]) );
  XOR U20 ( .A(B[1]), .B(A[1]), .Z(n20) );
  AND U21 ( .A(n21), .B(n22), .Z(n4) );
  NAND U22 ( .A(n23), .B(B[8]), .Z(n22) );
  NANDN U23 ( .A(A[8]), .B(n5), .Z(n23) );
  NANDN U24 ( .A(n5), .B(A[8]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n5) );
  NAND U26 ( .A(n26), .B(B[7]), .Z(n25) );
  NANDN U27 ( .A(A[7]), .B(n7), .Z(n26) );
  NANDN U28 ( .A(n7), .B(A[7]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n7) );
  NAND U30 ( .A(n29), .B(B[6]), .Z(n28) );
  NANDN U31 ( .A(A[6]), .B(n9), .Z(n29) );
  NANDN U32 ( .A(n9), .B(A[6]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n9) );
  NAND U34 ( .A(n32), .B(B[5]), .Z(n31) );
  NANDN U35 ( .A(A[5]), .B(n11), .Z(n32) );
  NANDN U36 ( .A(n11), .B(A[5]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n11) );
  NAND U38 ( .A(n35), .B(B[4]), .Z(n34) );
  NANDN U39 ( .A(A[4]), .B(n13), .Z(n35) );
  NANDN U40 ( .A(n13), .B(A[4]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n13) );
  NAND U42 ( .A(n38), .B(B[3]), .Z(n37) );
  NANDN U43 ( .A(A[3]), .B(n15), .Z(n38) );
  NANDN U44 ( .A(n15), .B(A[3]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n15) );
  NAND U46 ( .A(n41), .B(B[2]), .Z(n40) );
  NANDN U47 ( .A(A[2]), .B(n17), .Z(n41) );
  NANDN U48 ( .A(n17), .B(A[2]), .Z(n39) );
  AND U49 ( .A(n42), .B(n43), .Z(n17) );
  NAND U50 ( .A(n44), .B(B[1]), .Z(n43) );
  OR U51 ( .A(n19), .B(A[1]), .Z(n44) );
  NAND U52 ( .A(n19), .B(A[1]), .Z(n42) );
  AND U53 ( .A(B[0]), .B(A[0]), .Z(n19) );
  XOR U54 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_11 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_12 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_13 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_14 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_15 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_16 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_17 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_18 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_19 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_20 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_21 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_22 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_23 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_24 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_25 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_26 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_27 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_28 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_29 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_30 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_31 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_32 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_33 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_34 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_35 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_36 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_37 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_38 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_39 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_40 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_41 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_42 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_43 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_44 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_45 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_46 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_47 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_48 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_49 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_50 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_51 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_52 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_53 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_54 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_55 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_56 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_57 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_58 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_59 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_60 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_61 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_62 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_63 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_64 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_65 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_66 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_67 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_68 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_69 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_70 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_71 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_72 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_73 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_74 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_75 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_76 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_77 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_78 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_79 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_80 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_81 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_82 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_83 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  AND U1 ( .A(n2), .B(B[6]), .Z(SUM[7]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[6]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[4]) );
  XNOR U8 ( .A(B[4]), .B(A[4]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[3]) );
  XNOR U10 ( .A(B[3]), .B(A[3]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[2]) );
  XNOR U12 ( .A(B[2]), .B(A[2]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[1]) );
  XOR U14 ( .A(B[1]), .B(A[1]), .Z(n14) );
  AND U15 ( .A(n15), .B(n16), .Z(n4) );
  NAND U16 ( .A(n17), .B(B[5]), .Z(n16) );
  NANDN U17 ( .A(A[5]), .B(n5), .Z(n17) );
  NANDN U18 ( .A(n5), .B(A[5]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n5) );
  NAND U20 ( .A(n20), .B(B[4]), .Z(n19) );
  NANDN U21 ( .A(A[4]), .B(n7), .Z(n20) );
  NANDN U22 ( .A(n7), .B(A[4]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n7) );
  NAND U24 ( .A(n23), .B(B[3]), .Z(n22) );
  NANDN U25 ( .A(A[3]), .B(n9), .Z(n23) );
  NANDN U26 ( .A(n9), .B(A[3]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n9) );
  NAND U28 ( .A(n26), .B(B[2]), .Z(n25) );
  NANDN U29 ( .A(A[2]), .B(n11), .Z(n26) );
  NANDN U30 ( .A(n11), .B(A[2]), .Z(n24) );
  AND U31 ( .A(n27), .B(n28), .Z(n11) );
  NAND U32 ( .A(n29), .B(B[1]), .Z(n28) );
  OR U33 ( .A(n13), .B(A[1]), .Z(n29) );
  NAND U34 ( .A(n13), .B(A[1]), .Z(n27) );
  AND U35 ( .A(B[0]), .B(A[0]), .Z(n13) );
  XOR U36 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_84 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_85 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_86 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_87 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_88 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_89 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_90 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_91 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_92 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_93 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_94 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_95 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_96 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_97 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_98 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_99 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_100 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_101 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_102 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_103 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_104 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_105 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_106 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_107 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_108 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_109 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_110 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_111 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_112 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_113 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_114 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_115 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_116 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_117 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_118 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_119 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_120 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_121 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_122 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_123 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_124 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_125 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_126 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_127 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_128 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_129 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_130 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_131 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_132 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_133 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_134 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_135 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_136 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_137 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_138 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_139 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_140 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_141 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_142 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_143 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_144 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_145 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_146 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_147 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_148 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_149 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_150 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_151 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_152 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_153 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_154 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_155 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_156 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_157 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_158 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_159 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_160 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_161 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_162 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_163 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_164 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_165 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_166 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_167 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_168 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_169 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_170 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_171 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_172 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_173 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_174 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_175 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_176 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_177 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_178 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_179 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_180 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_181 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_182 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_183 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_184 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_185 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_186 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_187 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_188 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_189 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_190 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_191 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_192 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_193 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_194 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_195 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_196 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_197 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_198 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_199 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_200 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_201 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_202 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_203 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_204 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_205 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_206 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_207 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_208 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_209 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_210 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_211 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_212 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_213 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_214 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_215 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_216 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_217 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_218 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_219 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_220 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_221 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_222 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_223 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_224 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_225 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_226 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_227 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_228 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_229 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_230 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_231 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_232 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_233 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_234 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_235 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_236 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_237 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_238 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_239 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_240 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_241 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_242 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_243 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_244 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_245 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_246 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_247 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_248 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_249 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_250 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_251 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_252 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_253 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_254 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_255 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_256 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_257 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_258 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_259 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_260 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_261 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_262 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_263 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_264 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_265 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_266 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_267 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_268 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_269 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_270 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_271 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_272 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_273 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_274 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_275 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_276 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_277 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_278 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_279 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_280 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_281 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_282 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_283 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_284 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_285 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_286 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_287 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_288 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_289 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_290 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_291 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_292 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_293 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_294 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_295 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_296 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_297 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_298 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_299 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_300 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_301 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_302 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_303 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_304 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_305 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_306 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_307 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_308 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_309 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_310 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_311 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_312 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_313 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_314 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_315 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_316 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_317 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_318 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_319 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_320 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_321 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_322 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_323 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_324 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_325 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_326 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_327 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_328 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_329 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_330 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_331 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_332 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_333 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;

  AND U1 ( .A(n2), .B(B[4]), .Z(SUM[5]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[4]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[3]) );
  XNOR U6 ( .A(B[3]), .B(A[3]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[2]) );
  XNOR U8 ( .A(B[2]), .B(A[2]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[1]) );
  XOR U10 ( .A(B[1]), .B(A[1]), .Z(n10) );
  AND U11 ( .A(n11), .B(n12), .Z(n4) );
  NAND U12 ( .A(n13), .B(B[3]), .Z(n12) );
  NANDN U13 ( .A(A[3]), .B(n5), .Z(n13) );
  NANDN U14 ( .A(n5), .B(A[3]), .Z(n11) );
  AND U15 ( .A(n14), .B(n15), .Z(n5) );
  NAND U16 ( .A(n16), .B(B[2]), .Z(n15) );
  NANDN U17 ( .A(A[2]), .B(n7), .Z(n16) );
  NANDN U18 ( .A(n7), .B(A[2]), .Z(n14) );
  AND U19 ( .A(n17), .B(n18), .Z(n7) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n9), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n9), .B(A[1]), .Z(n17) );
  AND U23 ( .A(B[0]), .B(A[0]), .Z(n9) );
  XOR U24 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2 ( clk, rst, x, y, o );
  input [7999:0] x;
  input [7999:0] y;
  output [13:0] o;
  input clk, rst;
  wire   N60579, N60580, N60581, N60582, N60592, N60593, N60594, N60595,
         N60596, N60605, N60606, N60607, N60608, N60609, N60618, N60619,
         N60620, N60621, N60622, N60631, N60632, N60633, N60634, N60635,
         N60644, N60645, N60646, N60647, N60648, N60657, N60658, N60659,
         N60660, N60661, N60670, N60671, N60672, N60673, N60674, N60683,
         N60684, N60685, N60686, N60687, N60696, N60697, N60698, N60699,
         N60700, N60709, N60710, N60711, N60712, N60713, N60722, N60723,
         N60724, N60725, N60726, N60735, N60736, N60737, N60738, N60739,
         N60748, N60749, N60750, N60751, N60752, N60761, N60762, N60763,
         N60764, N60765, N60774, N60775, N60776, N60777, N60778, N60787,
         N60788, N60789, N60790, N60791, N60800, N60801, N60802, N60803,
         N60804, N60813, N60814, N60815, N60816, N60817, N60826, N60827,
         N60828, N60829, N60830, N60839, N60840, N60841, N60842, N60843,
         N60852, N60853, N60854, N60855, N60856, N60865, N60866, N60867,
         N60868, N60869, N60878, N60879, N60880, N60881, N60882, N60891,
         N60892, N60893, N60894, N60895, N60904, N60905, N60906, N60907,
         N60908, N60917, N60918, N60919, N60920, N60921, N60930, N60931,
         N60932, N60933, N60934, N60943, N60944, N60945, N60946, N60947,
         N60956, N60957, N60958, N60959, N60960, N60969, N60970, N60971,
         N60972, N60973, N60982, N60983, N60984, N60985, N60986, N60995,
         N60996, N60997, N60998, N60999, N61008, N61009, N61010, N61011,
         N61012, N61021, N61022, N61023, N61024, N61025, N61034, N61035,
         N61036, N61037, N61038, N61047, N61048, N61049, N61050, N61051,
         N61060, N61061, N61062, N61063, N61064, N61073, N61074, N61075,
         N61076, N61077, N61086, N61087, N61088, N61089, N61090, N61099,
         N61100, N61101, N61102, N61103, N61112, N61113, N61114, N61115,
         N61116, N61125, N61126, N61127, N61128, N61129, N61138, N61139,
         N61140, N61141, N61142, N61151, N61152, N61153, N61154, N61155,
         N61164, N61165, N61166, N61167, N61168, N61177, N61178, N61179,
         N61180, N61181, N61190, N61191, N61192, N61193, N61194, N61203,
         N61204, N61205, N61206, N61207, N61216, N61217, N61218, N61219,
         N61220, N61229, N61230, N61231, N61232, N61233, N61242, N61243,
         N61244, N61245, N61246, N61255, N61256, N61257, N61258, N61259,
         N61268, N61269, N61270, N61271, N61272, N61281, N61282, N61283,
         N61284, N61285, N61294, N61295, N61296, N61297, N61298, N61307,
         N61308, N61309, N61310, N61311, N61320, N61321, N61322, N61323,
         N61324, N61333, N61334, N61335, N61336, N61337, N61346, N61347,
         N61348, N61349, N61350, N61359, N61360, N61361, N61362, N61363,
         N61372, N61373, N61374, N61375, N61376, N61385, N61386, N61387,
         N61388, N61389, N61398, N61399, N61400, N61401, N61402, N61411,
         N61412, N61413, N61414, N61415, N61424, N61425, N61426, N61427,
         N61428, N61437, N61438, N61439, N61440, N61441, N61450, N61451,
         N61452, N61453, N61454, N61463, N61464, N61465, N61466, N61467,
         N61476, N61477, N61478, N61479, N61480, N61489, N61490, N61491,
         N61492, N61493, N61502, N61503, N61504, N61505, N61506, N61515,
         N61516, N61517, N61518, N61519, N61528, N61529, N61530, N61531,
         N61532, N61541, N61542, N61543, N61544, N61545, N61554, N61555,
         N61556, N61557, N61558, N61567, N61568, N61569, N61570, N61571,
         N61580, N61581, N61582, N61583, N61584, N61593, N61594, N61595,
         N61596, N61597, N61606, N61607, N61608, N61609, N61610, N61619,
         N61620, N61621, N61622, N61623, N61632, N61633, N61634, N61635,
         N61636, N61645, N61646, N61647, N61648, N61649, N61658, N61659,
         N61660, N61661, N61662, N61671, N61672, N61673, N61674, N61675,
         N61684, N61685, N61686, N61687, N61688, N61697, N61698, N61699,
         N61700, N61701, N61710, N61711, N61712, N61713, N61714, N61723,
         N61724, N61725, N61726, N61727, N61736, N61737, N61738, N61739,
         N61740, N61749, N61750, N61751, N61752, N61753, N61762, N61763,
         N61764, N61765, N61766, N61775, N61776, N61777, N61778, N61779,
         N61788, N61789, N61790, N61791, N61792, N61801, N61802, N61803,
         N61804, N61805, N61814, N61815, N61816, N61817, N61818, N61827,
         N61828, N61829, N61830, N61831, N61840, N61841, N61842, N61843,
         N61844, N61853, N61854, N61855, N61856, N61857, N61866, N61867,
         N61868, N61869, N61870, N61879, N61880, N61881, N61882, N61883,
         N61892, N61893, N61894, N61895, N61896, N61905, N61906, N61907,
         N61908, N61909, N61918, N61919, N61920, N61921, N61922, N61931,
         N61932, N61933, N61934, N61935, N61944, N61945, N61946, N61947,
         N61948, N61957, N61958, N61959, N61960, N61961, N61970, N61971,
         N61972, N61973, N61974, N61983, N61984, N61985, N61986, N61987,
         N61996, N61997, N61998, N61999, N62000, N62009, N62010, N62011,
         N62012, N62013, N62022, N62023, N62024, N62025, N62026, N62035,
         N62036, N62037, N62038, N62039, N62048, N62049, N62050, N62051,
         N62052, N62061, N62062, N62063, N62064, N62065, N62074, N62075,
         N62076, N62077, N62078, N62087, N62088, N62089, N62090, N62091,
         N62100, N62101, N62102, N62103, N62104, N62113, N62114, N62115,
         N62116, N62117, N62126, N62127, N62128, N62129, N62130, N62139,
         N62140, N62141, N62142, N62143, N62152, N62153, N62154, N62155,
         N62156, N62165, N62166, N62167, N62168, N62169, N62178, N62179,
         N62180, N62181, N62182, N62191, N62192, N62193, N62194, N62195,
         N62204, N62205, N62206, N62207, N62208, N62217, N62218, N62219,
         N62220, N62221, N62230, N62231, N62232, N62233, N62234, N62243,
         N62244, N62245, N62246, N62247, N62256, N62257, N62258, N62259,
         N62260, N62269, N62270, N62271, N62272, N62273, N62282, N62283,
         N62284, N62285, N62286, N62295, N62296, N62297, N62298, N62299,
         N62308, N62309, N62310, N62311, N62312, N62321, N62322, N62323,
         N62324, N62325, N62334, N62335, N62336, N62337, N62338, N62347,
         N62348, N62349, N62350, N62351, N62360, N62361, N62362, N62363,
         N62364, N62373, N62374, N62375, N62376, N62377, N62386, N62387,
         N62388, N62389, N62390, N62399, N62400, N62401, N62402, N62403,
         N62412, N62413, N62414, N62415, N62416, N62425, N62426, N62427,
         N62428, N62429, N62438, N62439, N62440, N62441, N62442, N62451,
         N62452, N62453, N62454, N62455, N62464, N62465, N62466, N62467,
         N62468, N62477, N62478, N62479, N62480, N62481, N62490, N62491,
         N62492, N62493, N62494, N62503, N62504, N62505, N62506, N62507,
         N62516, N62517, N62518, N62519, N62520, N62529, N62530, N62531,
         N62532, N62533, N62542, N62543, N62544, N62545, N62546, N62555,
         N62556, N62557, N62558, N62559, N62568, N62569, N62570, N62571,
         N62572, N62581, N62582, N62583, N62584, N62585, N62594, N62595,
         N62596, N62597, N62598, N62607, N62608, N62609, N62610, N62611,
         N62620, N62621, N62622, N62623, N62624, N62633, N62634, N62635,
         N62636, N62637, N62646, N62647, N62648, N62649, N62650, N62659,
         N62660, N62661, N62662, N62663, N62672, N62673, N62674, N62675,
         N62676, N62685, N62686, N62687, N62688, N62689, N62698, N62699,
         N62700, N62701, N62702, N62711, N62712, N62713, N62714, N62715,
         N62724, N62725, N62726, N62727, N62728, N62737, N62738, N62739,
         N62740, N62741, N62750, N62751, N62752, N62753, N62754, N62763,
         N62764, N62765, N62766, N62767, N62776, N62777, N62778, N62779,
         N62780, N62789, N62790, N62791, N62792, N62793, N62802, N62803,
         N62804, N62805, N62806, N62815, N62816, N62817, N62818, N62819,
         N62828, N62829, N62830, N62831, N62832, N62841, N62842, N62843,
         N62844, N62845, N62854, N62855, N62856, N62857, N62858, N62867,
         N62868, N62869, N62870, N62871, N62880, N62881, N62882, N62883,
         N62884, N62893, N62894, N62895, N62896, N62897, N62906, N62907,
         N62908, N62909, N62910, N62919, N62920, N62921, N62922, N62923,
         N62932, N62933, N62934, N62935, N62936, N62945, N62946, N62947,
         N62948, N62949, N62958, N62959, N62960, N62961, N62962, N62971,
         N62972, N62973, N62974, N62975, N62984, N62985, N62986, N62987,
         N62988, N62997, N62998, N62999, N63000, N63001, N63010, N63011,
         N63012, N63013, N63014, N63023, N63024, N63025, N63026, N63027,
         N63036, N63037, N63038, N63039, N63040, N63049, N63050, N63051,
         N63052, N63053, N63062, N63063, N63064, N63065, N63066, N63075,
         N63076, N63077, N63078, N63079, N63088, N63089, N63090, N63091,
         N63092, N63101, N63102, N63103, N63104, N63105, N63114, N63115,
         N63116, N63117, N63118, N63127, N63128, N63129, N63130, N63131,
         N63140, N63141, N63142, N63143, N63144, N63153, N63154, N63155,
         N63156, N63157, N63166, N63167, N63168, N63169, N63170, N63179,
         N63180, N63181, N63182, N63183, N63192, N63193, N63194, N63195,
         N63196, N63205, N63206, N63207, N63208, N63209, N63218, N63219,
         N63220, N63221, N63222, N63231, N63232, N63233, N63234, N63235,
         N63244, N63245, N63246, N63247, N63248, N63257, N63258, N63259,
         N63260, N63261, N63270, N63271, N63272, N63273, N63274, N63283,
         N63284, N63285, N63286, N63287, N63296, N63297, N63298, N63299,
         N63300, N63309, N63310, N63311, N63312, N63313, N63322, N63323,
         N63324, N63325, N63326, N63335, N63336, N63337, N63338, N63339,
         N63348, N63349, N63350, N63351, N63352, N63361, N63362, N63363,
         N63364, N63365, N63374, N63375, N63376, N63377, N63378, N63387,
         N63388, N63389, N63390, N63391, N63400, N63401, N63402, N63403,
         N63404, N63413, N63414, N63415, N63416, N63417, N63426, N63427,
         N63428, N63429, N63430, N63439, N63440, N63441, N63442, N63443,
         N63452, N63453, N63454, N63455, N63456, N63465, N63466, N63467,
         N63468, N63469, N63478, N63479, N63480, N63481, N63482, N63491,
         N63492, N63493, N63494, N63495, N63504, N63505, N63506, N63507,
         N63508, N63517, N63518, N63519, N63520, N63521, N63530, N63531,
         N63532, N63533, N63534, N63543, N63544, N63545, N63546, N63547,
         N63556, N63557, N63558, N63559, N63560, N63569, N63570, N63571,
         N63572, N63573, N63582, N63583, N63584, N63585, N63586, N63595,
         N63596, N63597, N63598, N63599, N63608, N63609, N63610, N63611,
         N63612, N63621, N63622, N63623, N63624, N63625, N63634, N63635,
         N63636, N63637, N63638, N63647, N63648, N63649, N63650, N63651,
         N63660, N63661, N63662, N63663, N63664, N63673, N63674, N63675,
         N63676, N63677, N63686, N63687, N63688, N63689, N63690, N63699,
         N63700, N63701, N63702, N63703, N63712, N63713, N63714, N63715,
         N63716, N63725, N63726, N63727, N63728, N63729, N63738, N63739,
         N63740, N63741, N63742, N63751, N63752, N63753, N63754, N63755,
         N63764, N63765, N63766, N63767, N63768, N63777, N63778, N63779,
         N63780, N63781, N63790, N63791, N63792, N63793, N63794, N63803,
         N63804, N63805, N63806, N63807, N63816, N63817, N63818, N63819,
         N63820, N63829, N63830, N63831, N63832, N63833, N63842, N63843,
         N63844, N63845, N63846, N63855, N63856, N63857, N63858, N63859,
         N63868, N63869, N63870, N63871, N63872, N63881, N63882, N63883,
         N63884, N63885, N63894, N63895, N63896, N63897, N63898, N63907,
         N63908, N63909, N63910, N63911, N63920, N63921, N63922, N63923,
         N63924, N63933, N63934, N63935, N63936, N63937, N63946, N63947,
         N63948, N63949, N63950, N63959, N63960, N63961, N63962, N63963,
         N63972, N63973, N63974, N63975, N63976, N63985, N63986, N63987,
         N63988, N63989, N63998, N63999, N64000, N64001, N64002, N64011,
         N64012, N64013, N64014, N64015, N64024, N64025, N64026, N64027,
         N64028, N64037, N64038, N64039, N64040, N64041, N64050, N64051,
         N64052, N64053, N64054, N64063, N64064, N64065, N64066, N64067,
         N64076, N64077, N64078, N64079, N64080, N64089, N64090, N64091,
         N64092, N64093, N64102, N64103, N64104, N64105, N64106, N64115,
         N64116, N64117, N64118, N64119, N64128, N64129, N64130, N64131,
         N64132, N64141, N64142, N64143, N64144, N64145, N64154, N64155,
         N64156, N64157, N64158, N64167, N64168, N64169, N64170, N64171,
         N64180, N64181, N64182, N64183, N64184, N64193, N64194, N64195,
         N64196, N64197, N64206, N64207, N64208, N64209, N64210, N64219,
         N64220, N64221, N64222, N64223, N64232, N64233, N64234, N64235,
         N64236, N64245, N64246, N64247, N64248, N64249, N64258, N64259,
         N64260, N64261, N64262, N64271, N64272, N64273, N64274, N64275,
         N64284, N64285, N64286, N64287, N64288, N64297, N64298, N64299,
         N64300, N64301, N64310, N64311, N64312, N64313, N64314, N64323,
         N64324, N64325, N64326, N64327, N64336, N64337, N64338, N64339,
         N64340, N64349, N64350, N64351, N64352, N64353, N64362, N64363,
         N64364, N64365, N64366, N64375, N64376, N64377, N64378, N64379,
         N64388, N64389, N64390, N64391, N64392, N64401, N64402, N64403,
         N64404, N64405, N64414, N64415, N64416, N64417, N64418, N64427,
         N64428, N64429, N64430, N64431, N64440, N64441, N64442, N64443,
         N64444, N64453, N64454, N64455, N64456, N64457, N64466, N64467,
         N64468, N64469, N64470, N64479, N64480, N64481, N64482, N64483,
         N64492, N64493, N64494, N64495, N64496, N64505, N64506, N64507,
         N64508, N64509, N64518, N64519, N64520, N64521, N64522, N64531,
         N64532, N64533, N64534, N64535, N64544, N64545, N64546, N64547,
         N64548, N64557, N64558, N64559, N64560, N64561, N64570, N64571,
         N64572, N64573, N64574, N64583, N64584, N64585, N64586, N64587,
         N64596, N64597, N64598, N64599, N64600, N64609, N64610, N64611,
         N64612, N64613, N64622, N64623, N64624, N64625, N64626, N64635,
         N64636, N64637, N64638, N64639, N64648, N64649, N64650, N64651,
         N64652, N64661, N64662, N64663, N64664, N64665, N64674, N64675,
         N64676, N64677, N64678, N64687, N64688, N64689, N64690, N64691,
         N64700, N64701, N64702, N64703, N64704, N64713, N64714, N64715,
         N64716, N64717, N64726, N64727, N64728, N64729, N64730, N64739,
         N64740, N64741, N64742, N64743, N64752, N64753, N64754, N64755,
         N64756, N64765, N64766, N64767, N64768, N64769, N64778, N64779,
         N64780, N64781, N64782, N64791, N64792, N64793, N64794, N64795,
         N64804, N64805, N64806, N64807, N64808, N64817, N64818, N64819,
         N64820, N64821, N64830, N64831, N64832, N64833, N64834, N64843,
         N64844, N64845, N64846, N64847, N64856, N64857, N64858, N64859,
         N64860, N64869, N64870, N64871, N64872, N64873, N64882, N64883,
         N64884, N64885, N64886, N64895, N64896, N64897, N64898, N64899,
         N64908, N64909, N64910, N64911, N64912, N64921, N64922, N64923,
         N64924, N64925, N64926, N64934, N64935, N64936, N64937, N64938,
         N64939, N64947, N64948, N64949, N64950, N64951, N64952, N64960,
         N64961, N64962, N64963, N64964, N64965, N64973, N64974, N64975,
         N64976, N64977, N64978, N64986, N64987, N64988, N64989, N64990,
         N64991, N64999, N65000, N65001, N65002, N65003, N65004, N65012,
         N65013, N65014, N65015, N65016, N65017, N65025, N65026, N65027,
         N65028, N65029, N65030, N65038, N65039, N65040, N65041, N65042,
         N65043, N65051, N65052, N65053, N65054, N65055, N65056, N65064,
         N65065, N65066, N65067, N65068, N65069, N65077, N65078, N65079,
         N65080, N65081, N65082, N65090, N65091, N65092, N65093, N65094,
         N65095, N65103, N65104, N65105, N65106, N65107, N65108, N65116,
         N65117, N65118, N65119, N65120, N65121, N65129, N65130, N65131,
         N65132, N65133, N65134, N65142, N65143, N65144, N65145, N65146,
         N65147, N65155, N65156, N65157, N65158, N65159, N65160, N65168,
         N65169, N65170, N65171, N65172, N65173, N65181, N65182, N65183,
         N65184, N65185, N65186, N65194, N65195, N65196, N65197, N65198,
         N65199, N65207, N65208, N65209, N65210, N65211, N65212, N65220,
         N65221, N65222, N65223, N65224, N65225, N65233, N65234, N65235,
         N65236, N65237, N65238, N65246, N65247, N65248, N65249, N65250,
         N65251, N65259, N65260, N65261, N65262, N65263, N65264, N65272,
         N65273, N65274, N65275, N65276, N65277, N65285, N65286, N65287,
         N65288, N65289, N65290, N65298, N65299, N65300, N65301, N65302,
         N65303, N65311, N65312, N65313, N65314, N65315, N65316, N65324,
         N65325, N65326, N65327, N65328, N65329, N65337, N65338, N65339,
         N65340, N65341, N65342, N65350, N65351, N65352, N65353, N65354,
         N65355, N65363, N65364, N65365, N65366, N65367, N65368, N65376,
         N65377, N65378, N65379, N65380, N65381, N65389, N65390, N65391,
         N65392, N65393, N65394, N65402, N65403, N65404, N65405, N65406,
         N65407, N65415, N65416, N65417, N65418, N65419, N65420, N65428,
         N65429, N65430, N65431, N65432, N65433, N65441, N65442, N65443,
         N65444, N65445, N65446, N65454, N65455, N65456, N65457, N65458,
         N65459, N65467, N65468, N65469, N65470, N65471, N65472, N65480,
         N65481, N65482, N65483, N65484, N65485, N65493, N65494, N65495,
         N65496, N65497, N65498, N65506, N65507, N65508, N65509, N65510,
         N65511, N65519, N65520, N65521, N65522, N65523, N65524, N65532,
         N65533, N65534, N65535, N65536, N65537, N65545, N65546, N65547,
         N65548, N65549, N65550, N65558, N65559, N65560, N65561, N65562,
         N65563, N65571, N65572, N65573, N65574, N65575, N65576, N65584,
         N65585, N65586, N65587, N65588, N65589, N65597, N65598, N65599,
         N65600, N65601, N65602, N65610, N65611, N65612, N65613, N65614,
         N65615, N65623, N65624, N65625, N65626, N65627, N65628, N65636,
         N65637, N65638, N65639, N65640, N65641, N65649, N65650, N65651,
         N65652, N65653, N65654, N65662, N65663, N65664, N65665, N65666,
         N65667, N65675, N65676, N65677, N65678, N65679, N65680, N65688,
         N65689, N65690, N65691, N65692, N65693, N65701, N65702, N65703,
         N65704, N65705, N65706, N65714, N65715, N65716, N65717, N65718,
         N65719, N65727, N65728, N65729, N65730, N65731, N65732, N65740,
         N65741, N65742, N65743, N65744, N65745, N65753, N65754, N65755,
         N65756, N65757, N65758, N65766, N65767, N65768, N65769, N65770,
         N65771, N65779, N65780, N65781, N65782, N65783, N65784, N65792,
         N65793, N65794, N65795, N65796, N65797, N65805, N65806, N65807,
         N65808, N65809, N65810, N65818, N65819, N65820, N65821, N65822,
         N65823, N65831, N65832, N65833, N65834, N65835, N65836, N65844,
         N65845, N65846, N65847, N65848, N65849, N65857, N65858, N65859,
         N65860, N65861, N65862, N65870, N65871, N65872, N65873, N65874,
         N65875, N65883, N65884, N65885, N65886, N65887, N65888, N65896,
         N65897, N65898, N65899, N65900, N65901, N65909, N65910, N65911,
         N65912, N65913, N65914, N65922, N65923, N65924, N65925, N65926,
         N65927, N65935, N65936, N65937, N65938, N65939, N65940, N65948,
         N65949, N65950, N65951, N65952, N65953, N65961, N65962, N65963,
         N65964, N65965, N65966, N65974, N65975, N65976, N65977, N65978,
         N65979, N65987, N65988, N65989, N65990, N65991, N65992, N66000,
         N66001, N66002, N66003, N66004, N66005, N66013, N66014, N66015,
         N66016, N66017, N66018, N66026, N66027, N66028, N66029, N66030,
         N66031, N66039, N66040, N66041, N66042, N66043, N66044, N66052,
         N66053, N66054, N66055, N66056, N66057, N66065, N66066, N66067,
         N66068, N66069, N66070, N66078, N66079, N66080, N66081, N66082,
         N66083, N66091, N66092, N66093, N66094, N66095, N66096, N66104,
         N66105, N66106, N66107, N66108, N66109, N66117, N66118, N66119,
         N66120, N66121, N66122, N66130, N66131, N66132, N66133, N66134,
         N66135, N66143, N66144, N66145, N66146, N66147, N66148, N66156,
         N66157, N66158, N66159, N66160, N66161, N66169, N66170, N66171,
         N66172, N66173, N66174, N66182, N66183, N66184, N66185, N66186,
         N66187, N66195, N66196, N66197, N66198, N66199, N66200, N66208,
         N66209, N66210, N66211, N66212, N66213, N66221, N66222, N66223,
         N66224, N66225, N66226, N66234, N66235, N66236, N66237, N66238,
         N66239, N66247, N66248, N66249, N66250, N66251, N66252, N66260,
         N66261, N66262, N66263, N66264, N66265, N66273, N66274, N66275,
         N66276, N66277, N66278, N66286, N66287, N66288, N66289, N66290,
         N66291, N66299, N66300, N66301, N66302, N66303, N66304, N66312,
         N66313, N66314, N66315, N66316, N66317, N66325, N66326, N66327,
         N66328, N66329, N66330, N66338, N66339, N66340, N66341, N66342,
         N66343, N66351, N66352, N66353, N66354, N66355, N66356, N66364,
         N66365, N66366, N66367, N66368, N66369, N66377, N66378, N66379,
         N66380, N66381, N66382, N66390, N66391, N66392, N66393, N66394,
         N66395, N66403, N66404, N66405, N66406, N66407, N66408, N66416,
         N66417, N66418, N66419, N66420, N66421, N66429, N66430, N66431,
         N66432, N66433, N66434, N66442, N66443, N66444, N66445, N66446,
         N66447, N66455, N66456, N66457, N66458, N66459, N66460, N66468,
         N66469, N66470, N66471, N66472, N66473, N66481, N66482, N66483,
         N66484, N66485, N66486, N66494, N66495, N66496, N66497, N66498,
         N66499, N66507, N66508, N66509, N66510, N66511, N66512, N66520,
         N66521, N66522, N66523, N66524, N66525, N66533, N66534, N66535,
         N66536, N66537, N66538, N66546, N66547, N66548, N66549, N66550,
         N66551, N66559, N66560, N66561, N66562, N66563, N66564, N66572,
         N66573, N66574, N66575, N66576, N66577, N66585, N66586, N66587,
         N66588, N66589, N66590, N66598, N66599, N66600, N66601, N66602,
         N66603, N66611, N66612, N66613, N66614, N66615, N66616, N66624,
         N66625, N66626, N66627, N66628, N66629, N66637, N66638, N66639,
         N66640, N66641, N66642, N66650, N66651, N66652, N66653, N66654,
         N66655, N66663, N66664, N66665, N66666, N66667, N66668, N66676,
         N66677, N66678, N66679, N66680, N66681, N66689, N66690, N66691,
         N66692, N66693, N66694, N66702, N66703, N66704, N66705, N66706,
         N66707, N66715, N66716, N66717, N66718, N66719, N66720, N66728,
         N66729, N66730, N66731, N66732, N66733, N66741, N66742, N66743,
         N66744, N66745, N66746, N66754, N66755, N66756, N66757, N66758,
         N66759, N66767, N66768, N66769, N66770, N66771, N66772, N66780,
         N66781, N66782, N66783, N66784, N66785, N66793, N66794, N66795,
         N66796, N66797, N66798, N66806, N66807, N66808, N66809, N66810,
         N66811, N66819, N66820, N66821, N66822, N66823, N66824, N66832,
         N66833, N66834, N66835, N66836, N66837, N66845, N66846, N66847,
         N66848, N66849, N66850, N66858, N66859, N66860, N66861, N66862,
         N66863, N66871, N66872, N66873, N66874, N66875, N66876, N66884,
         N66885, N66886, N66887, N66888, N66889, N66897, N66898, N66899,
         N66900, N66901, N66902, N66910, N66911, N66912, N66913, N66914,
         N66915, N66923, N66924, N66925, N66926, N66927, N66928, N66936,
         N66937, N66938, N66939, N66940, N66941, N66949, N66950, N66951,
         N66952, N66953, N66954, N66962, N66963, N66964, N66965, N66966,
         N66967, N66975, N66976, N66977, N66978, N66979, N66980, N66988,
         N66989, N66990, N66991, N66992, N66993, N67001, N67002, N67003,
         N67004, N67005, N67006, N67014, N67015, N67016, N67017, N67018,
         N67019, N67027, N67028, N67029, N67030, N67031, N67032, N67040,
         N67041, N67042, N67043, N67044, N67045, N67053, N67054, N67055,
         N67056, N67057, N67058, N67066, N67067, N67068, N67069, N67070,
         N67071, N67079, N67080, N67081, N67082, N67083, N67084, N67092,
         N67093, N67094, N67095, N67096, N67097, N67098, N67105, N67106,
         N67107, N67108, N67109, N67110, N67111, N67118, N67119, N67120,
         N67121, N67122, N67123, N67124, N67131, N67132, N67133, N67134,
         N67135, N67136, N67137, N67144, N67145, N67146, N67147, N67148,
         N67149, N67150, N67157, N67158, N67159, N67160, N67161, N67162,
         N67163, N67170, N67171, N67172, N67173, N67174, N67175, N67176,
         N67183, N67184, N67185, N67186, N67187, N67188, N67189, N67196,
         N67197, N67198, N67199, N67200, N67201, N67202, N67209, N67210,
         N67211, N67212, N67213, N67214, N67215, N67222, N67223, N67224,
         N67225, N67226, N67227, N67228, N67235, N67236, N67237, N67238,
         N67239, N67240, N67241, N67248, N67249, N67250, N67251, N67252,
         N67253, N67254, N67261, N67262, N67263, N67264, N67265, N67266,
         N67267, N67274, N67275, N67276, N67277, N67278, N67279, N67280,
         N67287, N67288, N67289, N67290, N67291, N67292, N67293, N67300,
         N67301, N67302, N67303, N67304, N67305, N67306, N67313, N67314,
         N67315, N67316, N67317, N67318, N67319, N67326, N67327, N67328,
         N67329, N67330, N67331, N67332, N67339, N67340, N67341, N67342,
         N67343, N67344, N67345, N67352, N67353, N67354, N67355, N67356,
         N67357, N67358, N67365, N67366, N67367, N67368, N67369, N67370,
         N67371, N67378, N67379, N67380, N67381, N67382, N67383, N67384,
         N67391, N67392, N67393, N67394, N67395, N67396, N67397, N67404,
         N67405, N67406, N67407, N67408, N67409, N67410, N67417, N67418,
         N67419, N67420, N67421, N67422, N67423, N67430, N67431, N67432,
         N67433, N67434, N67435, N67436, N67443, N67444, N67445, N67446,
         N67447, N67448, N67449, N67456, N67457, N67458, N67459, N67460,
         N67461, N67462, N67469, N67470, N67471, N67472, N67473, N67474,
         N67475, N67482, N67483, N67484, N67485, N67486, N67487, N67488,
         N67495, N67496, N67497, N67498, N67499, N67500, N67501, N67508,
         N67509, N67510, N67511, N67512, N67513, N67514, N67521, N67522,
         N67523, N67524, N67525, N67526, N67527, N67534, N67535, N67536,
         N67537, N67538, N67539, N67540, N67547, N67548, N67549, N67550,
         N67551, N67552, N67553, N67560, N67561, N67562, N67563, N67564,
         N67565, N67566, N67573, N67574, N67575, N67576, N67577, N67578,
         N67579, N67586, N67587, N67588, N67589, N67590, N67591, N67592,
         N67599, N67600, N67601, N67602, N67603, N67604, N67605, N67612,
         N67613, N67614, N67615, N67616, N67617, N67618, N67625, N67626,
         N67627, N67628, N67629, N67630, N67631, N67638, N67639, N67640,
         N67641, N67642, N67643, N67644, N67651, N67652, N67653, N67654,
         N67655, N67656, N67657, N67664, N67665, N67666, N67667, N67668,
         N67669, N67670, N67677, N67678, N67679, N67680, N67681, N67682,
         N67683, N67690, N67691, N67692, N67693, N67694, N67695, N67696,
         N67703, N67704, N67705, N67706, N67707, N67708, N67709, N67716,
         N67717, N67718, N67719, N67720, N67721, N67722, N67729, N67730,
         N67731, N67732, N67733, N67734, N67735, N67742, N67743, N67744,
         N67745, N67746, N67747, N67748, N67755, N67756, N67757, N67758,
         N67759, N67760, N67761, N67768, N67769, N67770, N67771, N67772,
         N67773, N67774, N67781, N67782, N67783, N67784, N67785, N67786,
         N67787, N67794, N67795, N67796, N67797, N67798, N67799, N67800,
         N67807, N67808, N67809, N67810, N67811, N67812, N67813, N67820,
         N67821, N67822, N67823, N67824, N67825, N67826, N67833, N67834,
         N67835, N67836, N67837, N67838, N67839, N67846, N67847, N67848,
         N67849, N67850, N67851, N67852, N67859, N67860, N67861, N67862,
         N67863, N67864, N67865, N67872, N67873, N67874, N67875, N67876,
         N67877, N67878, N67885, N67886, N67887, N67888, N67889, N67890,
         N67891, N67898, N67899, N67900, N67901, N67902, N67903, N67904,
         N67911, N67912, N67913, N67914, N67915, N67916, N67917, N67924,
         N67925, N67926, N67927, N67928, N67929, N67930, N67937, N67938,
         N67939, N67940, N67941, N67942, N67943, N67950, N67951, N67952,
         N67953, N67954, N67955, N67956, N67963, N67964, N67965, N67966,
         N67967, N67968, N67969, N67976, N67977, N67978, N67979, N67980,
         N67981, N67982, N67989, N67990, N67991, N67992, N67993, N67994,
         N67995, N68002, N68003, N68004, N68005, N68006, N68007, N68008,
         N68015, N68016, N68017, N68018, N68019, N68020, N68021, N68028,
         N68029, N68030, N68031, N68032, N68033, N68034, N68041, N68042,
         N68043, N68044, N68045, N68046, N68047, N68054, N68055, N68056,
         N68057, N68058, N68059, N68060, N68067, N68068, N68069, N68070,
         N68071, N68072, N68073, N68080, N68081, N68082, N68083, N68084,
         N68085, N68086, N68093, N68094, N68095, N68096, N68097, N68098,
         N68099, N68106, N68107, N68108, N68109, N68110, N68111, N68112,
         N68119, N68120, N68121, N68122, N68123, N68124, N68125, N68132,
         N68133, N68134, N68135, N68136, N68137, N68138, N68145, N68146,
         N68147, N68148, N68149, N68150, N68151, N68158, N68159, N68160,
         N68161, N68162, N68163, N68164, N68171, N68172, N68173, N68174,
         N68175, N68176, N68177, N68178, N68184, N68185, N68186, N68187,
         N68188, N68189, N68190, N68191, N68197, N68198, N68199, N68200,
         N68201, N68202, N68203, N68204, N68210, N68211, N68212, N68213,
         N68214, N68215, N68216, N68217, N68223, N68224, N68225, N68226,
         N68227, N68228, N68229, N68230, N68236, N68237, N68238, N68239,
         N68240, N68241, N68242, N68243, N68249, N68250, N68251, N68252,
         N68253, N68254, N68255, N68256, N68262, N68263, N68264, N68265,
         N68266, N68267, N68268, N68269, N68275, N68276, N68277, N68278,
         N68279, N68280, N68281, N68282, N68288, N68289, N68290, N68291,
         N68292, N68293, N68294, N68295, N68301, N68302, N68303, N68304,
         N68305, N68306, N68307, N68308, N68314, N68315, N68316, N68317,
         N68318, N68319, N68320, N68321, N68327, N68328, N68329, N68330,
         N68331, N68332, N68333, N68334, N68340, N68341, N68342, N68343,
         N68344, N68345, N68346, N68347, N68353, N68354, N68355, N68356,
         N68357, N68358, N68359, N68360, N68366, N68367, N68368, N68369,
         N68370, N68371, N68372, N68373, N68379, N68380, N68381, N68382,
         N68383, N68384, N68385, N68386, N68392, N68393, N68394, N68395,
         N68396, N68397, N68398, N68399, N68405, N68406, N68407, N68408,
         N68409, N68410, N68411, N68412, N68418, N68419, N68420, N68421,
         N68422, N68423, N68424, N68425, N68431, N68432, N68433, N68434,
         N68435, N68436, N68437, N68438, N68444, N68445, N68446, N68447,
         N68448, N68449, N68450, N68451, N68457, N68458, N68459, N68460,
         N68461, N68462, N68463, N68464, N68470, N68471, N68472, N68473,
         N68474, N68475, N68476, N68477, N68483, N68484, N68485, N68486,
         N68487, N68488, N68489, N68490, N68496, N68497, N68498, N68499,
         N68500, N68501, N68502, N68503, N68509, N68510, N68511, N68512,
         N68513, N68514, N68515, N68516, N68522, N68523, N68524, N68525,
         N68526, N68527, N68528, N68529, N68535, N68536, N68537, N68538,
         N68539, N68540, N68541, N68542, N68548, N68549, N68550, N68551,
         N68552, N68553, N68554, N68555, N68561, N68562, N68563, N68564,
         N68565, N68566, N68567, N68568, N68574, N68575, N68576, N68577,
         N68578, N68579, N68580, N68581, N68587, N68588, N68589, N68590,
         N68591, N68592, N68593, N68594, N68600, N68601, N68602, N68603,
         N68604, N68605, N68606, N68607, N68613, N68614, N68615, N68616,
         N68617, N68618, N68619, N68620, N68626, N68627, N68628, N68629,
         N68630, N68631, N68632, N68633, N68639, N68640, N68641, N68642,
         N68643, N68644, N68645, N68646, N68652, N68653, N68654, N68655,
         N68656, N68657, N68658, N68659, N68665, N68666, N68667, N68668,
         N68669, N68670, N68671, N68672, N68678, N68679, N68680, N68681,
         N68682, N68683, N68684, N68685, N68691, N68692, N68693, N68694,
         N68695, N68696, N68697, N68698, N68704, N68705, N68706, N68707,
         N68708, N68709, N68710, N68711, N68717, N68718, N68719, N68720,
         N68721, N68722, N68723, N68724, N68725, N68730, N68731, N68732,
         N68733, N68734, N68735, N68736, N68737, N68738, N68743, N68744,
         N68745, N68746, N68747, N68748, N68749, N68750, N68751, N68756,
         N68757, N68758, N68759, N68760, N68761, N68762, N68763, N68764,
         N68769, N68770, N68771, N68772, N68773, N68774, N68775, N68776,
         N68777, N68782, N68783, N68784, N68785, N68786, N68787, N68788,
         N68789, N68790, N68795, N68796, N68797, N68798, N68799, N68800,
         N68801, N68802, N68803, N68808, N68809, N68810, N68811, N68812,
         N68813, N68814, N68815, N68816, N68821, N68822, N68823, N68824,
         N68825, N68826, N68827, N68828, N68829, N68834, N68835, N68836,
         N68837, N68838, N68839, N68840, N68841, N68842, N68847, N68848,
         N68849, N68850, N68851, N68852, N68853, N68854, N68855, N68860,
         N68861, N68862, N68863, N68864, N68865, N68866, N68867, N68868,
         N68873, N68874, N68875, N68876, N68877, N68878, N68879, N68880,
         N68881, N68886, N68887, N68888, N68889, N68890, N68891, N68892,
         N68893, N68894, N68899, N68900, N68901, N68902, N68903, N68904,
         N68905, N68906, N68907, N68912, N68913, N68914, N68915, N68916,
         N68917, N68918, N68919, N68920, N68925, N68926, N68927, N68928,
         N68929, N68930, N68931, N68932, N68933, N68938, N68939, N68940,
         N68941, N68942, N68943, N68944, N68945, N68946, N68951, N68952,
         N68953, N68954, N68955, N68956, N68957, N68958, N68959, N68964,
         N68965, N68966, N68967, N68968, N68969, N68970, N68971, N68972,
         N68977, N68978, N68979, N68980, N68981, N68982, N68983, N68984,
         N68985, N68990, N68991, N68992, N68993, N68994, N68995, N68996,
         N68997, N68998, N68999, N69003, N69004, N69005, N69006, N69007,
         N69008, N69009, N69010, N69011, N69012, N69016, N69017, N69018,
         N69019, N69020, N69021, N69022, N69023, N69024, N69025, N69029,
         N69030, N69031, N69032, N69033, N69034, N69035, N69036, N69037,
         N69038, N69042, N69043, N69044, N69045, N69046, N69047, N69048,
         N69049, N69050, N69051, N69055, N69056, N69057, N69058, N69059,
         N69060, N69061, N69062, N69063, N69064, N69068, N69069, N69070,
         N69071, N69072, N69073, N69074, N69075, N69076, N69077, N69081,
         N69082, N69083, N69084, N69085, N69086, N69087, N69088, N69089,
         N69090, N69094, N69095, N69096, N69097, N69098, N69099, N69100,
         N69101, N69102, N69103, N69107, N69108, N69109, N69110, N69111,
         N69112, N69113, N69114, N69115, N69116, N69120, N69121, N69122,
         N69123, N69124, N69125, N69126, N69127, N69128, N69129, N69130,
         N69133, N69134, N69135, N69136, N69137, N69138, N69139, N69140,
         N69141, N69142, N69143, N69146, N69147, N69148, N69149, N69150,
         N69151, N69152, N69153, N69154, N69155, N69156, N69159, N69160,
         N69161, N69162, N69163, N69164, N69165, N69166, N69167, N69168,
         N69169, N69172, N69173, N69174, N69175, N69176, N69177, N69178,
         N69179, N69180, N69181, N69182, N69185, N69186, N69187, N69188,
         N69189, N69190, N69191, N69192, N69193, N69194, N69195, N69196,
         N69198, N69199, N69200, N69201, N69202, N69203, N69204, N69205,
         N69206, N69207, N69208, N69209, N69211, N69212, N69213, N69214,
         N69215, N69216, N69217, N69218, N69219, N69220, N69221, N69222,
         N69224, N69225, N69226, N69227, N69228, N69229, N69230, N69231,
         N69232, N69233, N69234, N69235, N69236, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
         n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390,
         n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
         n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
         n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414,
         n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
         n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
         n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
         n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446,
         n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
         n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462,
         n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470,
         n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
         n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486,
         n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494,
         n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
         n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510,
         n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
         n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
         n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534,
         n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
         n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
         n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558,
         n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566,
         n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574,
         n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582,
         n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
         n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598,
         n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606,
         n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614,
         n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
         n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630,
         n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638,
         n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646,
         n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654,
         n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662,
         n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670,
         n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678,
         n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
         n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
         n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702,
         n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710,
         n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718,
         n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726,
         n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734,
         n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
         n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750,
         n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
         n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766,
         n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774,
         n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782,
         n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790,
         n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798,
         n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806,
         n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814,
         n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822,
         n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830,
         n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838,
         n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846,
         n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854,
         n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862,
         n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870,
         n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
         n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886,
         n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894,
         n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902,
         n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
         n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918,
         n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926,
         n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934,
         n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942,
         n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950,
         n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958,
         n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966,
         n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974,
         n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982,
         n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990,
         n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998,
         n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
         n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014,
         n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022,
         n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030,
         n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038,
         n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046,
         n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054,
         n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062,
         n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070,
         n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
         n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086,
         n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094,
         n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102,
         n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110,
         n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118,
         n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
         n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134,
         n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142,
         n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
         n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158,
         n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166,
         n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174,
         n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182,
         n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
         n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
         n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206,
         n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214,
         n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
         n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230,
         n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238,
         n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
         n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
         n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262,
         n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
         n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278,
         n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286,
         n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294,
         n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302,
         n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310,
         n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318,
         n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326,
         n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334,
         n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342,
         n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350,
         n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358,
         n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366,
         n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374,
         n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382,
         n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390,
         n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398,
         n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406,
         n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414,
         n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422,
         n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430,
         n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438,
         n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446,
         n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454,
         n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462,
         n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470,
         n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478,
         n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486,
         n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494,
         n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502,
         n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510,
         n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518,
         n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526,
         n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534,
         n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542,
         n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550,
         n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558,
         n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566,
         n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574,
         n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582,
         n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590,
         n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598,
         n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606,
         n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614,
         n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622,
         n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630,
         n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638,
         n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646,
         n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654,
         n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662,
         n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670,
         n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678,
         n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686,
         n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694,
         n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702,
         n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710,
         n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718,
         n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726,
         n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734,
         n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742,
         n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750,
         n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758,
         n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766,
         n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774,
         n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782,
         n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790,
         n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798,
         n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806,
         n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814,
         n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822,
         n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830,
         n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838,
         n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846,
         n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854,
         n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862,
         n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870,
         n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878,
         n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886,
         n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894,
         n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902,
         n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910,
         n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918,
         n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926,
         n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934,
         n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942,
         n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950,
         n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958,
         n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966,
         n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974,
         n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982,
         n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990,
         n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998,
         n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006,
         n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014,
         n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022,
         n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030,
         n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038,
         n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046,
         n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054,
         n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062,
         n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070,
         n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078,
         n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086,
         n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094,
         n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102,
         n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110,
         n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118,
         n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126,
         n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134,
         n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142,
         n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150,
         n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158,
         n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166,
         n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174,
         n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182,
         n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190,
         n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198,
         n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206,
         n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214,
         n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222,
         n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230,
         n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238,
         n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246,
         n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254,
         n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262,
         n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270,
         n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278,
         n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286,
         n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294,
         n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302,
         n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310,
         n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318,
         n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326,
         n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334,
         n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342,
         n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350,
         n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358,
         n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366,
         n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374,
         n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382,
         n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390,
         n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398,
         n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406,
         n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414,
         n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422,
         n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430,
         n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438,
         n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446,
         n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454,
         n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462,
         n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470,
         n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478,
         n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486,
         n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494,
         n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502,
         n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510,
         n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518,
         n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526,
         n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534,
         n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542,
         n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550,
         n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558,
         n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566,
         n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574,
         n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582,
         n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590,
         n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598,
         n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606,
         n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614,
         n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622,
         n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630,
         n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638,
         n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646,
         n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654,
         n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662,
         n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670,
         n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678,
         n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686,
         n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694,
         n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702,
         n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710,
         n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718,
         n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726,
         n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734,
         n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742,
         n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750,
         n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758,
         n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766,
         n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774,
         n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782,
         n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790,
         n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798,
         n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806,
         n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814,
         n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822,
         n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830,
         n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838,
         n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846,
         n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854,
         n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862,
         n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870,
         n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878,
         n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886,
         n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894,
         n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902,
         n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910,
         n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918,
         n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926,
         n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934,
         n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942,
         n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950,
         n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958,
         n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966,
         n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974,
         n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982,
         n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990,
         n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998,
         n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006,
         n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014,
         n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022,
         n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030,
         n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038,
         n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046,
         n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054,
         n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062,
         n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070,
         n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078,
         n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086,
         n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094,
         n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102,
         n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110,
         n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118,
         n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126,
         n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134,
         n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142,
         n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150,
         n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158,
         n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166,
         n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174,
         n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182,
         n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190,
         n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198,
         n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206,
         n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214,
         n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222,
         n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230,
         n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238,
         n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246,
         n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254,
         n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262,
         n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270,
         n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278,
         n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286,
         n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294,
         n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302,
         n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310,
         n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318,
         n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326,
         n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334,
         n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342,
         n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350,
         n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358,
         n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366,
         n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374,
         n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382,
         n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390,
         n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398,
         n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406,
         n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414,
         n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422,
         n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430,
         n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438,
         n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446,
         n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454,
         n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462,
         n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470,
         n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478,
         n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486,
         n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494,
         n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502,
         n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510,
         n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518,
         n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526,
         n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534,
         n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542,
         n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550,
         n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558,
         n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566,
         n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574,
         n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582,
         n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590,
         n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598,
         n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606,
         n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614,
         n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622,
         n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630,
         n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638,
         n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646,
         n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654,
         n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662,
         n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670,
         n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678,
         n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686,
         n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694,
         n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702,
         n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710,
         n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718,
         n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726,
         n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734,
         n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742,
         n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750,
         n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758,
         n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766,
         n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774,
         n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782,
         n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790,
         n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798,
         n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806,
         n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814,
         n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822,
         n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830,
         n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838,
         n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846,
         n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854,
         n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862,
         n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870,
         n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878,
         n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886,
         n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894,
         n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902,
         n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910,
         n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918,
         n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926,
         n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934,
         n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942,
         n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950,
         n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958,
         n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966,
         n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974,
         n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982,
         n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990,
         n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998,
         n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006,
         n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014,
         n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022,
         n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030,
         n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038,
         n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046,
         n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054,
         n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062,
         n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070,
         n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078,
         n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086,
         n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094,
         n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102,
         n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110,
         n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118,
         n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126,
         n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134,
         n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142,
         n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150,
         n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158,
         n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166,
         n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174,
         n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182,
         n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190,
         n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198,
         n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206,
         n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214,
         n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222,
         n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230,
         n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238,
         n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246,
         n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254,
         n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262,
         n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270,
         n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278,
         n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286,
         n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294,
         n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302,
         n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310,
         n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318,
         n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326,
         n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334,
         n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342,
         n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350,
         n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358,
         n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366,
         n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374,
         n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382,
         n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390,
         n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398,
         n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406,
         n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414,
         n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422,
         n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430,
         n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438,
         n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446,
         n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454,
         n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462,
         n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470,
         n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478,
         n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486,
         n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494,
         n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502,
         n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510,
         n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518,
         n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526,
         n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534,
         n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542,
         n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550,
         n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558,
         n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566,
         n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574,
         n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582,
         n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590,
         n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598,
         n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606,
         n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614,
         n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622,
         n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630,
         n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638,
         n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646,
         n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654,
         n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662,
         n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670,
         n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678,
         n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686,
         n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694,
         n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702,
         n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710,
         n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718,
         n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726,
         n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734,
         n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742,
         n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750,
         n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758,
         n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766,
         n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774,
         n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782,
         n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790,
         n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798,
         n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806,
         n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814,
         n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822,
         n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830,
         n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838,
         n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846,
         n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854,
         n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862,
         n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870,
         n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878,
         n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886,
         n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894,
         n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902,
         n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910,
         n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918,
         n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926,
         n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934,
         n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942,
         n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950,
         n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958,
         n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966,
         n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974,
         n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982,
         n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990,
         n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998,
         n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006,
         n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014,
         n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022,
         n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030,
         n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038,
         n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046,
         n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054,
         n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062,
         n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070,
         n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078,
         n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086,
         n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094,
         n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102,
         n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110,
         n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118,
         n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126,
         n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134,
         n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142,
         n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150,
         n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158,
         n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166,
         n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174,
         n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182,
         n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190,
         n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
         n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206,
         n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214,
         n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222,
         n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230,
         n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238,
         n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246,
         n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254,
         n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262,
         n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
         n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278,
         n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286,
         n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294,
         n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302,
         n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310,
         n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318,
         n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326,
         n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334,
         n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342,
         n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350,
         n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358,
         n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366,
         n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374,
         n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382,
         n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390,
         n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398,
         n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406,
         n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414,
         n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422,
         n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430,
         n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438,
         n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446,
         n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454,
         n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462,
         n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470,
         n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478,
         n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486,
         n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494,
         n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502,
         n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510,
         n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518,
         n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526,
         n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534,
         n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542,
         n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550,
         n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558,
         n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566,
         n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574,
         n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582,
         n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590,
         n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598,
         n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606,
         n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614,
         n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622,
         n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630,
         n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638,
         n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646,
         n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654,
         n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662,
         n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670,
         n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678,
         n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686,
         n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694,
         n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702,
         n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710,
         n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718,
         n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726,
         n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734,
         n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742,
         n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750,
         n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758,
         n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766,
         n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774,
         n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782,
         n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790,
         n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798,
         n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806,
         n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814,
         n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822,
         n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830,
         n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838,
         n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846,
         n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854,
         n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862,
         n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870,
         n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878,
         n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886,
         n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894,
         n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902,
         n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910,
         n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918,
         n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926,
         n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934,
         n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942,
         n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950,
         n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958,
         n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966,
         n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974,
         n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982,
         n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990,
         n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998,
         n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006,
         n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014,
         n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022,
         n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030,
         n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038,
         n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046,
         n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054,
         n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062,
         n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070,
         n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078,
         n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086,
         n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094,
         n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102,
         n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110,
         n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118,
         n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126,
         n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134,
         n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142,
         n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150,
         n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158,
         n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166,
         n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174,
         n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182,
         n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190,
         n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198,
         n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206,
         n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214,
         n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222,
         n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230,
         n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238,
         n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246,
         n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254,
         n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262,
         n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270,
         n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278,
         n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286,
         n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294,
         n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302,
         n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310,
         n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318,
         n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326,
         n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334,
         n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342,
         n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350,
         n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358,
         n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366,
         n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374,
         n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382,
         n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390,
         n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398,
         n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406,
         n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414,
         n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422,
         n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430,
         n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438,
         n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446,
         n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454,
         n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462,
         n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470,
         n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478,
         n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486,
         n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494,
         n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502,
         n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510,
         n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518,
         n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526,
         n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534,
         n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542,
         n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550,
         n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558,
         n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566,
         n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574,
         n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582,
         n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590,
         n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598,
         n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606,
         n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614,
         n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622,
         n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630,
         n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638,
         n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646,
         n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654,
         n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662,
         n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670,
         n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678,
         n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686,
         n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694,
         n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702,
         n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710,
         n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718,
         n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726,
         n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734,
         n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742,
         n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750,
         n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758,
         n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766,
         n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774,
         n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782,
         n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790,
         n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798,
         n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806,
         n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814,
         n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822,
         n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830,
         n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838,
         n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846,
         n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854,
         n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862,
         n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870,
         n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878,
         n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886,
         n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894,
         n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902,
         n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910,
         n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918,
         n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926,
         n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934,
         n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942,
         n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950,
         n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958,
         n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966,
         n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974,
         n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982,
         n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990,
         n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998,
         n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006,
         n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014,
         n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022,
         n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030,
         n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038,
         n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046,
         n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054,
         n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062,
         n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070,
         n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078,
         n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086,
         n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094,
         n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102,
         n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110,
         n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118,
         n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126,
         n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134,
         n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142,
         n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150,
         n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158,
         n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166,
         n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174,
         n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182,
         n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190,
         n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198,
         n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206,
         n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214,
         n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222,
         n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230,
         n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238,
         n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246,
         n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254,
         n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262,
         n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270,
         n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278,
         n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286,
         n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294,
         n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302,
         n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310,
         n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318,
         n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326,
         n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334,
         n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342,
         n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350,
         n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358,
         n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366,
         n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374,
         n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382,
         n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390,
         n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398,
         n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406,
         n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414,
         n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422,
         n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430,
         n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
         n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446,
         n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454,
         n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462,
         n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470,
         n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478,
         n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486,
         n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494,
         n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502,
         n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510,
         n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518,
         n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526,
         n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534,
         n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542,
         n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550,
         n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558,
         n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566,
         n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574,
         n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582,
         n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590,
         n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598,
         n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606,
         n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614,
         n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622,
         n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630,
         n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638,
         n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646,
         n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654,
         n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662,
         n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670,
         n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678,
         n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686,
         n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694,
         n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702,
         n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710,
         n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718,
         n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726,
         n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734,
         n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742,
         n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750,
         n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758,
         n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766,
         n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774,
         n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782,
         n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790,
         n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798,
         n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806,
         n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814,
         n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822,
         n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830,
         n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838,
         n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846,
         n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854,
         n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862,
         n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870,
         n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878,
         n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886,
         n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894,
         n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902,
         n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910,
         n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918,
         n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926,
         n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934,
         n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942,
         n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950,
         n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958,
         n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966,
         n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974,
         n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982,
         n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990,
         n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998,
         n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006,
         n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014,
         n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022,
         n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030,
         n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038,
         n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046,
         n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054,
         n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062,
         n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070,
         n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078,
         n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086,
         n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094,
         n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102,
         n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110,
         n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118,
         n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126,
         n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134,
         n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142,
         n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150,
         n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158,
         n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166,
         n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174,
         n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182,
         n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190,
         n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198,
         n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206,
         n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214,
         n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222,
         n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230,
         n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238,
         n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246,
         n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254,
         n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262,
         n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270,
         n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278,
         n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286,
         n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294,
         n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302,
         n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310,
         n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318,
         n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326,
         n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334,
         n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342,
         n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350,
         n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358,
         n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366,
         n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374,
         n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382,
         n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390,
         n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398,
         n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406,
         n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414,
         n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
         n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430,
         n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438,
         n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446,
         n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454,
         n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462,
         n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470,
         n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478,
         n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486,
         n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494,
         n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502,
         n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510,
         n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518,
         n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526,
         n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534,
         n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542,
         n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550,
         n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558,
         n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566,
         n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574,
         n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582,
         n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590,
         n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598,
         n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606,
         n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614,
         n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622,
         n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630,
         n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638,
         n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646,
         n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654,
         n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662,
         n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670,
         n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678,
         n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686,
         n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694,
         n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702,
         n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
         n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718,
         n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726,
         n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734,
         n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742,
         n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750,
         n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758,
         n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766,
         n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774,
         n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782,
         n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790,
         n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798,
         n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806,
         n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814,
         n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822,
         n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830,
         n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838,
         n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846,
         n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
         n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862,
         n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870,
         n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878,
         n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886,
         n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894,
         n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902,
         n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910,
         n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918,
         n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926,
         n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934,
         n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942,
         n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950,
         n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958,
         n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966,
         n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974,
         n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982,
         n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990,
         n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998,
         n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006,
         n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014,
         n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022,
         n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030,
         n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038,
         n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046,
         n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054,
         n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062,
         n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070,
         n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078,
         n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086,
         n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094,
         n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102,
         n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110,
         n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118,
         n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126,
         n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134,
         n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
         n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150,
         n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158,
         n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166,
         n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174,
         n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182,
         n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190,
         n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198,
         n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206,
         n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214,
         n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222,
         n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230,
         n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238,
         n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246,
         n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254,
         n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262,
         n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270,
         n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278,
         n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286,
         n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294,
         n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302,
         n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310,
         n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318,
         n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326,
         n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334,
         n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342,
         n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350,
         n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358,
         n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366,
         n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374,
         n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382,
         n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390,
         n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398,
         n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406,
         n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414,
         n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422,
         n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430,
         n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438,
         n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446,
         n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454,
         n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462,
         n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470,
         n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478,
         n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486,
         n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494,
         n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
         n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510,
         n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518,
         n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526,
         n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534,
         n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542,
         n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550,
         n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558,
         n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566,
         n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574,
         n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582,
         n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590,
         n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598,
         n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606,
         n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614,
         n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622,
         n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630,
         n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638,
         n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646,
         n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654,
         n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662,
         n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670,
         n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678,
         n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686,
         n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694,
         n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702,
         n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710,
         n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718,
         n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726,
         n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734,
         n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742,
         n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750,
         n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758,
         n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766,
         n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774,
         n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782,
         n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790,
         n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798,
         n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806,
         n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814,
         n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822,
         n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830,
         n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838,
         n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846,
         n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854,
         n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862,
         n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870,
         n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878,
         n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886,
         n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894,
         n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902,
         n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910,
         n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918,
         n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926,
         n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934,
         n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942,
         n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950,
         n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958,
         n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966,
         n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974,
         n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982,
         n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990,
         n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998,
         n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006,
         n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014,
         n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022,
         n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030,
         n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038,
         n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046,
         n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054,
         n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062,
         n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070,
         n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078,
         n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086,
         n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094,
         n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102,
         n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110,
         n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118,
         n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126,
         n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134,
         n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142,
         n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150,
         n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158,
         n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166,
         n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174,
         n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182,
         n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190,
         n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198,
         n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206,
         n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214,
         n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222,
         n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230,
         n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238,
         n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246,
         n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254,
         n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262,
         n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270,
         n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278,
         n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286,
         n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294,
         n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302,
         n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310,
         n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318,
         n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326,
         n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334,
         n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342,
         n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350,
         n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358,
         n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366,
         n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374,
         n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382,
         n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390,
         n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398,
         n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406,
         n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414,
         n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422,
         n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430,
         n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438,
         n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446,
         n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454,
         n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462,
         n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470,
         n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478,
         n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
         n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494,
         n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502,
         n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510,
         n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518,
         n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526,
         n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534,
         n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542,
         n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550,
         n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558,
         n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566,
         n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574,
         n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582,
         n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590,
         n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598,
         n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606,
         n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614,
         n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622,
         n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630,
         n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638,
         n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646,
         n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654,
         n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662,
         n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670,
         n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678,
         n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686,
         n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694,
         n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702,
         n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710,
         n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718,
         n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726,
         n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734,
         n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742,
         n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750,
         n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758,
         n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766,
         n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774,
         n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782,
         n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790,
         n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798,
         n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806,
         n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814,
         n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822,
         n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830,
         n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838,
         n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846,
         n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854,
         n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862,
         n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870,
         n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878,
         n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886,
         n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894,
         n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902,
         n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910,
         n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918,
         n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926,
         n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934,
         n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942,
         n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950,
         n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958,
         n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966,
         n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974,
         n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982,
         n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990,
         n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998,
         n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006,
         n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014,
         n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022,
         n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030,
         n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038,
         n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046,
         n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054,
         n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062,
         n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070,
         n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078,
         n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086,
         n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094,
         n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102,
         n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110,
         n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118,
         n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126,
         n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134,
         n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142,
         n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150,
         n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158,
         n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166,
         n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174,
         n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182,
         n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190,
         n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198,
         n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206,
         n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214,
         n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222,
         n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230,
         n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238,
         n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246,
         n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254,
         n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262,
         n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270,
         n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278,
         n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286,
         n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294,
         n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302,
         n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310,
         n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318,
         n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326,
         n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334,
         n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342,
         n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350,
         n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358,
         n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366,
         n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374,
         n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382,
         n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390,
         n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398,
         n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406,
         n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414,
         n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422,
         n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430,
         n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438,
         n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446,
         n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454,
         n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462,
         n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470,
         n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478,
         n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486,
         n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494,
         n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502,
         n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510,
         n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518,
         n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526,
         n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534,
         n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542,
         n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550,
         n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558,
         n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566,
         n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574,
         n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582,
         n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590,
         n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598,
         n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606,
         n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614,
         n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622,
         n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630,
         n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638,
         n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646,
         n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654,
         n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662,
         n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670,
         n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678,
         n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686,
         n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694,
         n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702,
         n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710,
         n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718,
         n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726,
         n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734,
         n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742,
         n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750,
         n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758,
         n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766,
         n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774,
         n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782,
         n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790,
         n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798,
         n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806,
         n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814,
         n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822,
         n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830,
         n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838,
         n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846,
         n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854,
         n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862,
         n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870,
         n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878,
         n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886,
         n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
         n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902,
         n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910,
         n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918,
         n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926,
         n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934,
         n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942,
         n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
         n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958,
         n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
         n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974,
         n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982,
         n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990,
         n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998,
         n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006,
         n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014,
         n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022,
         n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030,
         n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038,
         n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046,
         n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054,
         n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062,
         n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070,
         n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078,
         n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086,
         n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094,
         n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102,
         n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110,
         n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118,
         n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126,
         n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134,
         n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142,
         n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150,
         n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158,
         n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166,
         n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174,
         n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
         n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190,
         n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198,
         n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206,
         n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214,
         n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222,
         n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230,
         n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238,
         n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246,
         n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254,
         n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262,
         n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270,
         n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278,
         n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286,
         n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294,
         n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302,
         n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310,
         n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318,
         n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326,
         n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334,
         n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342,
         n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350,
         n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
         n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366,
         n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374,
         n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382,
         n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390,
         n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398,
         n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406,
         n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414,
         n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422,
         n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430,
         n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438,
         n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446,
         n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454,
         n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462,
         n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470,
         n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478,
         n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486,
         n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494,
         n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502,
         n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510,
         n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518,
         n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526,
         n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534,
         n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542,
         n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550,
         n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558,
         n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566,
         n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574,
         n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582,
         n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590,
         n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598,
         n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606,
         n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614,
         n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622,
         n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630,
         n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
         n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646,
         n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654,
         n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662,
         n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670,
         n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678,
         n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
         n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
         n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702,
         n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
         n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718,
         n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726,
         n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734,
         n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
         n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750,
         n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
         n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766,
         n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
         n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782,
         n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790,
         n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798,
         n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806,
         n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
         n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822,
         n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
         n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838,
         n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846,
         n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
         n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862,
         n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870,
         n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878,
         n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886,
         n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894,
         n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902,
         n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910,
         n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918,
         n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
         n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934,
         n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942,
         n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950,
         n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
         n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966,
         n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974,
         n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982,
         n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990,
         n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998,
         n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006,
         n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014,
         n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022,
         n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030,
         n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038,
         n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046,
         n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054,
         n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062,
         n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
         n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
         n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086,
         n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094,
         n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
         n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110,
         n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
         n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
         n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134,
         n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142,
         n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150,
         n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158,
         n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166,
         n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174,
         n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182,
         n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190,
         n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198,
         n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206,
         n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214,
         n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222,
         n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230,
         n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238,
         n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246,
         n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254,
         n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262,
         n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270,
         n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278,
         n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286,
         n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294,
         n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302,
         n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310,
         n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318,
         n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326,
         n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334,
         n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342,
         n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350,
         n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358,
         n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366,
         n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374,
         n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382,
         n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390,
         n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398,
         n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406,
         n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414,
         n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422,
         n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430,
         n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438,
         n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446,
         n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454,
         n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462,
         n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470,
         n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478,
         n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486,
         n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494,
         n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502,
         n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510,
         n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518,
         n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526,
         n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534,
         n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542,
         n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550,
         n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558,
         n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566,
         n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574,
         n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582,
         n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590,
         n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598,
         n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606,
         n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614,
         n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622,
         n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630,
         n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638,
         n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646,
         n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654,
         n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662,
         n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670,
         n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678,
         n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686,
         n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694,
         n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702,
         n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710,
         n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718,
         n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726,
         n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734,
         n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742,
         n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750,
         n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758,
         n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766,
         n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774,
         n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782,
         n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790,
         n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798,
         n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806,
         n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814,
         n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822,
         n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830,
         n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838,
         n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846,
         n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854,
         n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862,
         n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870,
         n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878,
         n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886,
         n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894,
         n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902,
         n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910,
         n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918,
         n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926,
         n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934,
         n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942,
         n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950,
         n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958,
         n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966,
         n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974,
         n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982,
         n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990,
         n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998,
         n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006,
         n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014,
         n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022,
         n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030,
         n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038,
         n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046,
         n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054,
         n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062,
         n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070,
         n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078,
         n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086,
         n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094,
         n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102,
         n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110,
         n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118,
         n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126,
         n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134,
         n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142,
         n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150,
         n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158,
         n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166,
         n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174,
         n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182,
         n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190,
         n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198,
         n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206,
         n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214,
         n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222,
         n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230,
         n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238,
         n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246,
         n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254,
         n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262,
         n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270,
         n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278,
         n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286,
         n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294,
         n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302,
         n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310,
         n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318,
         n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326,
         n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334,
         n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342,
         n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350,
         n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358,
         n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366,
         n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374,
         n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382,
         n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390,
         n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398,
         n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406,
         n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414,
         n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422,
         n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430,
         n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438,
         n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446,
         n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454,
         n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462,
         n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470,
         n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478,
         n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486,
         n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494,
         n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502,
         n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510,
         n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518,
         n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526,
         n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534,
         n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542,
         n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550,
         n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558,
         n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566,
         n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574,
         n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582,
         n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590,
         n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598,
         n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606,
         n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614,
         n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622,
         n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630,
         n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638,
         n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646,
         n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654,
         n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662,
         n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670,
         n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678,
         n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686,
         n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694,
         n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702,
         n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710,
         n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718,
         n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726,
         n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734,
         n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742,
         n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750,
         n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758,
         n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766,
         n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774,
         n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782,
         n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790,
         n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798,
         n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806,
         n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814,
         n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822,
         n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830,
         n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838,
         n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846,
         n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854,
         n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862,
         n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870,
         n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878,
         n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886,
         n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894,
         n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902,
         n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910,
         n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918,
         n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926,
         n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934,
         n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942,
         n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950,
         n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958,
         n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966,
         n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974,
         n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982,
         n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990,
         n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998,
         n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006,
         n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014,
         n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022,
         n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030,
         n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038,
         n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046,
         n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054,
         n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062,
         n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070,
         n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078,
         n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086,
         n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094,
         n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102,
         n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110,
         n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118,
         n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126,
         n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134,
         n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142,
         n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150,
         n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158,
         n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166,
         n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174,
         n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182,
         n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190,
         n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198,
         n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206,
         n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214,
         n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222,
         n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230,
         n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238,
         n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246,
         n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254,
         n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262,
         n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270,
         n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278,
         n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286,
         n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294,
         n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302,
         n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310,
         n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318,
         n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326,
         n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334,
         n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342,
         n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350,
         n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358,
         n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366,
         n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374,
         n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382,
         n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390,
         n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398,
         n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406,
         n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414,
         n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422,
         n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430,
         n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438,
         n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446,
         n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454,
         n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462,
         n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470,
         n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478,
         n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486,
         n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494,
         n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502,
         n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510,
         n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518,
         n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526,
         n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534,
         n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542,
         n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550,
         n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558,
         n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566,
         n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574,
         n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582,
         n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590,
         n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598,
         n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606,
         n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614,
         n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622,
         n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630,
         n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638,
         n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646,
         n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654,
         n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662,
         n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670,
         n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678,
         n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686,
         n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694,
         n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702,
         n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710,
         n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718,
         n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726,
         n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734,
         n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742,
         n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750,
         n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758,
         n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766,
         n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774,
         n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782,
         n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790,
         n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798,
         n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806,
         n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814,
         n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822,
         n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830,
         n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838,
         n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846,
         n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854,
         n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862,
         n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870,
         n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878,
         n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886,
         n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894,
         n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902,
         n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910,
         n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918,
         n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926,
         n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934,
         n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942,
         n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950,
         n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958,
         n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966,
         n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974,
         n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982,
         n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990,
         n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998,
         n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006,
         n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014,
         n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022,
         n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030,
         n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038,
         n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046,
         n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054,
         n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062,
         n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070,
         n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078,
         n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086,
         n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094,
         n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102,
         n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110,
         n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118,
         n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126,
         n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134,
         n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142,
         n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150,
         n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158,
         n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166,
         n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174,
         n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182,
         n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190,
         n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198,
         n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206,
         n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214,
         n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222,
         n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230,
         n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238,
         n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246,
         n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254,
         n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262,
         n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270,
         n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278,
         n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286,
         n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294,
         n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302,
         n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310,
         n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318,
         n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326,
         n37327, n37328, n37329, n37330, n37331, n37332, n37333, n37334,
         n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342,
         n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350,
         n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358,
         n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366,
         n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374,
         n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382,
         n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390,
         n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398,
         n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406,
         n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414,
         n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422,
         n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430,
         n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438,
         n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446,
         n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454,
         n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462,
         n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470,
         n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478,
         n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486,
         n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494,
         n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502,
         n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510,
         n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518,
         n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526,
         n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534,
         n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542,
         n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550,
         n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558,
         n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566,
         n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574,
         n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582,
         n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590,
         n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598,
         n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606,
         n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614,
         n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622,
         n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630,
         n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638,
         n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646,
         n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654,
         n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662,
         n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670,
         n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678,
         n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686,
         n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694,
         n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702,
         n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710,
         n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718,
         n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726,
         n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734,
         n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742,
         n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750,
         n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758,
         n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766,
         n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774,
         n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782,
         n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790,
         n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798,
         n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806,
         n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814,
         n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822,
         n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830,
         n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838,
         n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846,
         n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854,
         n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862,
         n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870,
         n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878,
         n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886,
         n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894,
         n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902,
         n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910,
         n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918,
         n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926,
         n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934,
         n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942,
         n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950,
         n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958,
         n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966,
         n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974,
         n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982,
         n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990,
         n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998,
         n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006,
         n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014,
         n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022,
         n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030,
         n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038,
         n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046,
         n38047, n38048, n38049, n38050, n38051, n38052, n38053, n38054,
         n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062,
         n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070,
         n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078,
         n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086,
         n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094,
         n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102,
         n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110,
         n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118,
         n38119, n38120, n38121, n38122, n38123, n38124, n38125, n38126,
         n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134,
         n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142,
         n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150,
         n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158,
         n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166,
         n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174,
         n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182,
         n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190,
         n38191, n38192, n38193, n38194, n38195, n38196, n38197, n38198,
         n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206,
         n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214,
         n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222,
         n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230,
         n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238,
         n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246,
         n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254,
         n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262,
         n38263, n38264, n38265, n38266, n38267, n38268, n38269, n38270,
         n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278,
         n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286,
         n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294,
         n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302,
         n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310,
         n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318,
         n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326,
         n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334,
         n38335, n38336, n38337, n38338, n38339, n38340, n38341, n38342,
         n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350,
         n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358,
         n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366,
         n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374,
         n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382,
         n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390,
         n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398,
         n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406,
         n38407, n38408, n38409, n38410, n38411, n38412, n38413, n38414,
         n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422,
         n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430,
         n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438,
         n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446,
         n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454,
         n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462,
         n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470,
         n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478,
         n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486,
         n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494,
         n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502,
         n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510,
         n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518,
         n38519, n38520, n38521, n38522, n38523, n38524, n38525, n38526,
         n38527, n38528, n38529, n38530, n38531, n38532, n38533, n38534,
         n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542,
         n38543, n38544, n38545, n38546, n38547, n38548, n38549, n38550,
         n38551, n38552, n38553, n38554, n38555, n38556, n38557, n38558,
         n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566,
         n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574,
         n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582,
         n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590,
         n38591, n38592, n38593, n38594, n38595, n38596, n38597, n38598,
         n38599, n38600, n38601, n38602, n38603, n38604, n38605, n38606,
         n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614,
         n38615, n38616, n38617, n38618, n38619, n38620, n38621, n38622,
         n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630,
         n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638,
         n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646,
         n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654,
         n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662,
         n38663, n38664, n38665, n38666, n38667, n38668, n38669, n38670,
         n38671, n38672, n38673, n38674, n38675, n38676, n38677, n38678,
         n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686,
         n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694,
         n38695, n38696, n38697, n38698, n38699, n38700, n38701, n38702,
         n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710,
         n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718,
         n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726,
         n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734,
         n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742,
         n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750,
         n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758,
         n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766,
         n38767, n38768, n38769, n38770, n38771, n38772, n38773, n38774,
         n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782,
         n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790,
         n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798,
         n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806,
         n38807, n38808, n38809, n38810, n38811, n38812, n38813, n38814,
         n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822,
         n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830,
         n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838,
         n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846,
         n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854,
         n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862,
         n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870,
         n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878,
         n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886,
         n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894,
         n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902,
         n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910,
         n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918,
         n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926,
         n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934,
         n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942,
         n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950,
         n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958,
         n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966,
         n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974,
         n38975, n38976, n38977, n38978, n38979, n38980, n38981, n38982,
         n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990,
         n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998,
         n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006,
         n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014,
         n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022,
         n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030,
         n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038,
         n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046,
         n39047, n39048, n39049, n39050, n39051, n39052, n39053, n39054,
         n39055, n39056, n39057, n39058, n39059, n39060, n39061, n39062,
         n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070,
         n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078,
         n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086,
         n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094,
         n39095, n39096, n39097, n39098, n39099, n39100, n39101, n39102,
         n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110,
         n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118,
         n39119, n39120, n39121, n39122, n39123, n39124, n39125, n39126,
         n39127, n39128, n39129, n39130, n39131, n39132, n39133, n39134,
         n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142,
         n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150,
         n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158,
         n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166,
         n39167, n39168, n39169, n39170, n39171, n39172, n39173, n39174,
         n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182,
         n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190,
         n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198,
         n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206,
         n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214,
         n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222,
         n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230,
         n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238,
         n39239, n39240, n39241, n39242, n39243, n39244, n39245, n39246,
         n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254,
         n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262,
         n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270,
         n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278,
         n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286,
         n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294,
         n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302,
         n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310,
         n39311, n39312, n39313, n39314, n39315, n39316, n39317, n39318,
         n39319, n39320, n39321, n39322, n39323, n39324, n39325, n39326,
         n39327, n39328, n39329, n39330, n39331, n39332, n39333, n39334,
         n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342,
         n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350,
         n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358,
         n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366,
         n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374,
         n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382,
         n39383, n39384, n39385, n39386, n39387, n39388, n39389, n39390,
         n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398,
         n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406,
         n39407, n39408, n39409, n39410, n39411, n39412, n39413, n39414,
         n39415, n39416, n39417, n39418, n39419, n39420, n39421, n39422,
         n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430,
         n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438,
         n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446,
         n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454,
         n39455, n39456, n39457, n39458, n39459, n39460, n39461, n39462,
         n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470,
         n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478,
         n39479, n39480, n39481, n39482, n39483, n39484, n39485, n39486,
         n39487, n39488, n39489, n39490, n39491, n39492, n39493, n39494,
         n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502,
         n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510,
         n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518,
         n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526,
         n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534,
         n39535, n39536, n39537, n39538, n39539, n39540, n39541, n39542,
         n39543, n39544, n39545, n39546, n39547, n39548, n39549, n39550,
         n39551, n39552, n39553, n39554, n39555, n39556, n39557, n39558,
         n39559, n39560, n39561, n39562, n39563, n39564, n39565, n39566,
         n39567, n39568, n39569, n39570, n39571, n39572, n39573, n39574,
         n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582,
         n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590,
         n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598,
         n39599, n39600, n39601, n39602, n39603, n39604, n39605, n39606,
         n39607, n39608, n39609, n39610, n39611, n39612, n39613, n39614,
         n39615, n39616, n39617, n39618, n39619, n39620, n39621, n39622,
         n39623, n39624, n39625, n39626, n39627, n39628, n39629, n39630,
         n39631, n39632, n39633, n39634, n39635, n39636, n39637, n39638,
         n39639, n39640, n39641, n39642, n39643, n39644, n39645, n39646,
         n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654,
         n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662,
         n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670,
         n39671, n39672, n39673, n39674, n39675, n39676, n39677, n39678,
         n39679, n39680, n39681, n39682, n39683, n39684, n39685, n39686,
         n39687, n39688, n39689, n39690, n39691, n39692, n39693, n39694,
         n39695, n39696, n39697, n39698, n39699, n39700, n39701, n39702,
         n39703, n39704, n39705, n39706, n39707, n39708, n39709, n39710,
         n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718,
         n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726,
         n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734,
         n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742,
         n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750,
         n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758,
         n39759, n39760, n39761, n39762, n39763, n39764, n39765, n39766,
         n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774,
         n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782,
         n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790,
         n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798,
         n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806,
         n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814,
         n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822,
         n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830,
         n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838,
         n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846,
         n39847, n39848, n39849, n39850, n39851, n39852, n39853, n39854,
         n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862,
         n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870,
         n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878,
         n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886,
         n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894,
         n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902,
         n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910,
         n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918,
         n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926,
         n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934,
         n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942,
         n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950,
         n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958,
         n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966,
         n39967, n39968, n39969, n39970, n39971, n39972, n39973, n39974,
         n39975, n39976, n39977, n39978, n39979, n39980, n39981, n39982,
         n39983, n39984, n39985, n39986, n39987, n39988, n39989, n39990,
         n39991, n39992, n39993, n39994, n39995, n39996, n39997, n39998,
         n39999, n40000, n40001, n40002, n40003, n40004, n40005, n40006,
         n40007, n40008, n40009, n40010, n40011, n40012, n40013, n40014,
         n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022,
         n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030,
         n40031, n40032, n40033, n40034, n40035, n40036, n40037, n40038,
         n40039, n40040, n40041, n40042, n40043, n40044, n40045, n40046,
         n40047, n40048, n40049, n40050, n40051, n40052, n40053, n40054,
         n40055, n40056, n40057, n40058, n40059, n40060, n40061, n40062,
         n40063, n40064, n40065, n40066, n40067, n40068, n40069, n40070,
         n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078,
         n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086,
         n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094,
         n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102,
         n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110,
         n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118,
         n40119, n40120, n40121, n40122, n40123, n40124, n40125, n40126,
         n40127, n40128, n40129, n40130, n40131, n40132, n40133, n40134,
         n40135, n40136, n40137, n40138, n40139, n40140, n40141, n40142,
         n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150,
         n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158,
         n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166,
         n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174,
         n40175, n40176, n40177, n40178, n40179, n40180, n40181, n40182,
         n40183, n40184, n40185, n40186, n40187, n40188, n40189, n40190,
         n40191, n40192, n40193, n40194, n40195, n40196, n40197, n40198,
         n40199, n40200, n40201, n40202, n40203, n40204, n40205, n40206,
         n40207, n40208, n40209, n40210, n40211, n40212, n40213, n40214,
         n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222,
         n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230,
         n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238,
         n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246,
         n40247, n40248, n40249, n40250, n40251, n40252, n40253, n40254,
         n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40262,
         n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270,
         n40271, n40272, n40273, n40274, n40275, n40276, n40277, n40278,
         n40279, n40280, n40281, n40282, n40283, n40284, n40285, n40286,
         n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294,
         n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302,
         n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310,
         n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318,
         n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326,
         n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334,
         n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342,
         n40343, n40344, n40345, n40346, n40347, n40348, n40349, n40350,
         n40351, n40352, n40353, n40354, n40355, n40356, n40357, n40358,
         n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366,
         n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374,
         n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382,
         n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390,
         n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398,
         n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406,
         n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414,
         n40415, n40416, n40417, n40418, n40419, n40420, n40421, n40422,
         n40423, n40424, n40425, n40426, n40427, n40428, n40429, n40430,
         n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438,
         n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446,
         n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454,
         n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462,
         n40463, n40464, n40465, n40466, n40467, n40468, n40469, n40470,
         n40471, n40472, n40473, n40474, n40475, n40476, n40477, n40478,
         n40479, n40480, n40481, n40482, n40483, n40484, n40485, n40486,
         n40487, n40488, n40489, n40490, n40491, n40492, n40493, n40494,
         n40495, n40496, n40497, n40498, n40499, n40500, n40501, n40502,
         n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510,
         n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518,
         n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526,
         n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534,
         n40535, n40536, n40537, n40538, n40539, n40540, n40541, n40542,
         n40543, n40544, n40545, n40546, n40547, n40548, n40549, n40550,
         n40551, n40552, n40553, n40554, n40555, n40556, n40557, n40558,
         n40559, n40560, n40561, n40562, n40563, n40564, n40565, n40566,
         n40567, n40568, n40569, n40570, n40571, n40572, n40573, n40574,
         n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582,
         n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590,
         n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598,
         n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606,
         n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614,
         n40615, n40616, n40617, n40618, n40619, n40620, n40621, n40622,
         n40623, n40624, n40625, n40626, n40627, n40628, n40629, n40630,
         n40631, n40632, n40633, n40634, n40635, n40636, n40637, n40638,
         n40639, n40640, n40641, n40642, n40643, n40644, n40645, n40646,
         n40647, n40648, n40649, n40650, n40651, n40652, n40653, n40654,
         n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662,
         n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670,
         n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678,
         n40679, n40680, n40681, n40682, n40683, n40684, n40685, n40686,
         n40687, n40688, n40689, n40690, n40691, n40692, n40693, n40694,
         n40695, n40696, n40697, n40698, n40699, n40700, n40701, n40702,
         n40703, n40704, n40705, n40706, n40707, n40708, n40709, n40710,
         n40711, n40712, n40713, n40714, n40715, n40716, n40717, n40718,
         n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726,
         n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734,
         n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742,
         n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750,
         n40751, n40752, n40753, n40754, n40755, n40756, n40757, n40758,
         n40759, n40760, n40761, n40762, n40763, n40764, n40765, n40766,
         n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774,
         n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782,
         n40783, n40784, n40785, n40786, n40787, n40788, n40789, n40790,
         n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798,
         n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806,
         n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814,
         n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822,
         n40823, n40824, n40825, n40826, n40827, n40828, n40829, n40830,
         n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838,
         n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846,
         n40847, n40848, n40849, n40850, n40851, n40852, n40853, n40854,
         n40855, n40856, n40857, n40858, n40859, n40860, n40861, n40862,
         n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870,
         n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878,
         n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886,
         n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894,
         n40895, n40896, n40897, n40898, n40899, n40900, n40901, n40902,
         n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910,
         n40911, n40912, n40913, n40914, n40915, n40916, n40917, n40918,
         n40919, n40920, n40921, n40922, n40923, n40924, n40925, n40926,
         n40927, n40928, n40929, n40930, n40931, n40932, n40933, n40934,
         n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942,
         n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950,
         n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958,
         n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966,
         n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974,
         n40975, n40976, n40977, n40978, n40979, n40980, n40981, n40982,
         n40983, n40984, n40985, n40986, n40987, n40988, n40989, n40990,
         n40991, n40992, n40993, n40994, n40995, n40996, n40997, n40998,
         n40999, n41000, n41001, n41002, n41003, n41004, n41005, n41006,
         n41007, n41008, n41009, n41010, n41011, n41012, n41013, n41014,
         n41015, n41016, n41017, n41018, n41019, n41020, n41021, n41022,
         n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030,
         n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038,
         n41039, n41040, n41041, n41042, n41043, n41044, n41045, n41046,
         n41047, n41048, n41049, n41050, n41051, n41052, n41053, n41054,
         n41055, n41056, n41057, n41058, n41059, n41060, n41061, n41062,
         n41063, n41064, n41065, n41066, n41067, n41068, n41069, n41070,
         n41071, n41072, n41073, n41074, n41075, n41076, n41077, n41078,
         n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086,
         n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094,
         n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102,
         n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110,
         n41111, n41112, n41113, n41114, n41115, n41116, n41117, n41118,
         n41119, n41120, n41121, n41122, n41123, n41124, n41125, n41126,
         n41127, n41128, n41129, n41130, n41131, n41132, n41133, n41134,
         n41135, n41136, n41137, n41138, n41139, n41140, n41141, n41142,
         n41143, n41144, n41145, n41146, n41147, n41148, n41149, n41150,
         n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158,
         n41159, n41160, n41161, n41162, n41163, n41164, n41165, n41166,
         n41167, n41168, n41169, n41170, n41171, n41172, n41173, n41174,
         n41175, n41176, n41177, n41178, n41179, n41180, n41181, n41182,
         n41183, n41184, n41185, n41186, n41187, n41188, n41189, n41190,
         n41191, n41192, n41193, n41194, n41195, n41196, n41197, n41198,
         n41199, n41200, n41201, n41202, n41203, n41204, n41205, n41206,
         n41207, n41208, n41209, n41210, n41211, n41212, n41213, n41214,
         n41215, n41216, n41217, n41218, n41219, n41220, n41221, n41222,
         n41223, n41224, n41225, n41226, n41227, n41228, n41229, n41230,
         n41231, n41232, n41233, n41234, n41235, n41236, n41237, n41238,
         n41239, n41240, n41241, n41242, n41243, n41244, n41245, n41246,
         n41247, n41248, n41249, n41250, n41251, n41252, n41253, n41254,
         n41255, n41256, n41257, n41258, n41259, n41260, n41261, n41262,
         n41263, n41264, n41265, n41266, n41267, n41268, n41269, n41270,
         n41271, n41272, n41273, n41274, n41275, n41276, n41277, n41278,
         n41279, n41280, n41281, n41282, n41283, n41284, n41285, n41286,
         n41287, n41288, n41289, n41290, n41291, n41292, n41293, n41294,
         n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302,
         n41303, n41304, n41305, n41306, n41307, n41308, n41309, n41310,
         n41311, n41312, n41313, n41314, n41315, n41316, n41317, n41318,
         n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326,
         n41327, n41328, n41329, n41330, n41331, n41332, n41333, n41334,
         n41335, n41336, n41337, n41338, n41339, n41340, n41341, n41342,
         n41343, n41344, n41345, n41346, n41347, n41348, n41349, n41350,
         n41351, n41352, n41353, n41354, n41355, n41356, n41357, n41358,
         n41359, n41360, n41361, n41362, n41363, n41364, n41365, n41366,
         n41367, n41368, n41369, n41370, n41371, n41372, n41373, n41374,
         n41375, n41376, n41377, n41378, n41379, n41380, n41381, n41382,
         n41383, n41384, n41385, n41386, n41387, n41388, n41389, n41390,
         n41391, n41392, n41393, n41394, n41395, n41396, n41397, n41398,
         n41399, n41400, n41401, n41402, n41403, n41404, n41405, n41406,
         n41407, n41408, n41409, n41410, n41411, n41412, n41413, n41414,
         n41415, n41416, n41417, n41418, n41419, n41420, n41421, n41422,
         n41423, n41424, n41425, n41426, n41427, n41428, n41429, n41430,
         n41431, n41432, n41433, n41434, n41435, n41436, n41437, n41438,
         n41439, n41440, n41441, n41442, n41443, n41444, n41445, n41446,
         n41447, n41448, n41449, n41450, n41451, n41452, n41453, n41454,
         n41455, n41456, n41457, n41458, n41459, n41460, n41461, n41462,
         n41463, n41464, n41465, n41466, n41467, n41468, n41469, n41470,
         n41471, n41472, n41473, n41474, n41475, n41476, n41477, n41478,
         n41479, n41480, n41481, n41482, n41483, n41484, n41485, n41486,
         n41487, n41488, n41489, n41490, n41491, n41492, n41493, n41494,
         n41495, n41496, n41497, n41498, n41499, n41500, n41501, n41502,
         n41503, n41504, n41505, n41506, n41507, n41508, n41509, n41510,
         n41511, n41512, n41513, n41514, n41515, n41516, n41517, n41518,
         n41519, n41520, n41521, n41522, n41523, n41524, n41525, n41526,
         n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534,
         n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542,
         n41543, n41544, n41545, n41546, n41547, n41548, n41549, n41550,
         n41551, n41552, n41553, n41554, n41555, n41556, n41557, n41558,
         n41559, n41560, n41561, n41562, n41563, n41564, n41565, n41566,
         n41567, n41568, n41569, n41570, n41571, n41572, n41573, n41574,
         n41575, n41576, n41577, n41578, n41579, n41580, n41581, n41582,
         n41583, n41584, n41585, n41586, n41587, n41588, n41589, n41590,
         n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598,
         n41599, n41600, n41601, n41602, n41603, n41604, n41605, n41606,
         n41607, n41608, n41609, n41610, n41611, n41612, n41613, n41614,
         n41615, n41616, n41617, n41618, n41619, n41620, n41621, n41622,
         n41623, n41624, n41625, n41626, n41627, n41628, n41629, n41630,
         n41631, n41632, n41633, n41634, n41635, n41636, n41637, n41638,
         n41639, n41640, n41641, n41642, n41643, n41644, n41645, n41646,
         n41647, n41648, n41649, n41650, n41651, n41652, n41653, n41654,
         n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662,
         n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670,
         n41671, n41672, n41673, n41674, n41675, n41676, n41677, n41678,
         n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686,
         n41687, n41688, n41689, n41690, n41691, n41692, n41693, n41694,
         n41695, n41696, n41697, n41698, n41699, n41700, n41701, n41702,
         n41703, n41704, n41705, n41706, n41707, n41708, n41709, n41710,
         n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718,
         n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41726,
         n41727, n41728, n41729, n41730, n41731, n41732, n41733, n41734,
         n41735, n41736, n41737, n41738, n41739, n41740, n41741, n41742,
         n41743, n41744, n41745, n41746, n41747, n41748, n41749, n41750,
         n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758,
         n41759, n41760, n41761, n41762, n41763, n41764, n41765, n41766,
         n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774,
         n41775, n41776, n41777, n41778, n41779, n41780, n41781, n41782,
         n41783, n41784, n41785, n41786, n41787, n41788, n41789, n41790,
         n41791, n41792, n41793, n41794, n41795, n41796, n41797, n41798,
         n41799, n41800, n41801, n41802, n41803, n41804, n41805, n41806,
         n41807, n41808, n41809, n41810, n41811, n41812, n41813, n41814,
         n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822,
         n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830,
         n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838,
         n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846,
         n41847, n41848, n41849, n41850, n41851, n41852, n41853, n41854,
         n41855, n41856, n41857, n41858, n41859, n41860, n41861, n41862,
         n41863, n41864, n41865, n41866, n41867, n41868, n41869, n41870,
         n41871, n41872, n41873, n41874, n41875, n41876, n41877, n41878,
         n41879, n41880, n41881, n41882, n41883, n41884, n41885, n41886,
         n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894,
         n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902,
         n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910,
         n41911, n41912, n41913, n41914, n41915, n41916, n41917, n41918,
         n41919, n41920, n41921, n41922, n41923, n41924, n41925, n41926,
         n41927, n41928, n41929, n41930, n41931, n41932, n41933, n41934,
         n41935, n41936, n41937, n41938, n41939, n41940, n41941, n41942,
         n41943, n41944, n41945, n41946, n41947, n41948, n41949, n41950,
         n41951, n41952, n41953, n41954, n41955, n41956, n41957, n41958,
         n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966,
         n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974,
         n41975, n41976, n41977, n41978, n41979, n41980, n41981, n41982,
         n41983, n41984, n41985, n41986, n41987, n41988, n41989, n41990,
         n41991, n41992, n41993, n41994, n41995, n41996, n41997, n41998,
         n41999, n42000, n42001, n42002, n42003, n42004, n42005, n42006,
         n42007, n42008, n42009, n42010, n42011, n42012, n42013, n42014,
         n42015, n42016, n42017, n42018, n42019, n42020, n42021, n42022,
         n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030,
         n42031, n42032, n42033, n42034, n42035, n42036, n42037, n42038,
         n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046,
         n42047, n42048, n42049, n42050, n42051, n42052, n42053, n42054,
         n42055, n42056, n42057, n42058, n42059, n42060, n42061, n42062,
         n42063, n42064, n42065, n42066, n42067, n42068, n42069, n42070,
         n42071, n42072, n42073, n42074, n42075, n42076, n42077, n42078,
         n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42086,
         n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094,
         n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102,
         n42103, n42104, n42105, n42106, n42107, n42108, n42109, n42110,
         n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118,
         n42119, n42120, n42121, n42122, n42123, n42124, n42125, n42126,
         n42127, n42128, n42129, n42130, n42131, n42132, n42133, n42134,
         n42135, n42136, n42137, n42138, n42139, n42140, n42141, n42142,
         n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150,
         n42151, n42152, n42153, n42154, n42155, n42156, n42157, n42158,
         n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166,
         n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174,
         n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182,
         n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190,
         n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198,
         n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206,
         n42207, n42208, n42209, n42210, n42211, n42212, n42213, n42214,
         n42215, n42216, n42217, n42218, n42219, n42220, n42221, n42222,
         n42223, n42224, n42225, n42226, n42227, n42228, n42229, n42230,
         n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238,
         n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246,
         n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254,
         n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262,
         n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270,
         n42271, n42272, n42273, n42274, n42275, n42276, n42277, n42278,
         n42279, n42280, n42281, n42282, n42283, n42284, n42285, n42286,
         n42287, n42288, n42289, n42290, n42291, n42292, n42293, n42294,
         n42295, n42296, n42297, n42298, n42299, n42300, n42301, n42302,
         n42303, n42304, n42305, n42306, n42307, n42308, n42309, n42310,
         n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318,
         n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326,
         n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334,
         n42335, n42336, n42337, n42338, n42339, n42340, n42341, n42342,
         n42343, n42344, n42345, n42346, n42347, n42348, n42349, n42350,
         n42351, n42352, n42353, n42354, n42355, n42356, n42357, n42358,
         n42359, n42360, n42361, n42362, n42363, n42364, n42365, n42366,
         n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374,
         n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382,
         n42383, n42384, n42385, n42386, n42387, n42388, n42389, n42390,
         n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398,
         n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406,
         n42407, n42408, n42409, n42410, n42411, n42412, n42413, n42414,
         n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42422,
         n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430,
         n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438,
         n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446,
         n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454,
         n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462,
         n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470,
         n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478,
         n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486,
         n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494,
         n42495, n42496, n42497, n42498, n42499, n42500, n42501, n42502,
         n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510,
         n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518,
         n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42526,
         n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534,
         n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542,
         n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550,
         n42551, n42552, n42553, n42554, n42555, n42556, n42557, n42558,
         n42559, n42560, n42561, n42562, n42563, n42564, n42565, n42566,
         n42567, n42568, n42569, n42570, n42571, n42572, n42573, n42574,
         n42575, n42576, n42577, n42578, n42579, n42580, n42581, n42582,
         n42583, n42584, n42585, n42586, n42587, n42588, n42589, n42590,
         n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598,
         n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606,
         n42607, n42608, n42609, n42610, n42611, n42612, n42613, n42614,
         n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622,
         n42623, n42624, n42625, n42626, n42627, n42628, n42629, n42630,
         n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638,
         n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646,
         n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654,
         n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662,
         n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670,
         n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678,
         n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686,
         n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694,
         n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702,
         n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710,
         n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718,
         n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726,
         n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734,
         n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742,
         n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750,
         n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758,
         n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766,
         n42767, n42768, n42769, n42770, n42771, n42772, n42773, n42774,
         n42775, n42776, n42777, n42778, n42779, n42780, n42781, n42782,
         n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790,
         n42791, n42792, n42793, n42794, n42795, n42796, n42797, n42798,
         n42799, n42800, n42801, n42802, n42803, n42804, n42805, n42806,
         n42807, n42808, n42809, n42810, n42811, n42812, n42813, n42814,
         n42815, n42816, n42817, n42818, n42819, n42820, n42821, n42822,
         n42823, n42824, n42825, n42826, n42827, n42828, n42829, n42830,
         n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838,
         n42839, n42840, n42841, n42842, n42843, n42844, n42845, n42846,
         n42847, n42848, n42849, n42850, n42851, n42852, n42853, n42854,
         n42855, n42856, n42857, n42858, n42859, n42860, n42861, n42862,
         n42863, n42864, n42865, n42866, n42867, n42868, n42869, n42870,
         n42871, n42872, n42873, n42874, n42875, n42876, n42877, n42878,
         n42879, n42880, n42881, n42882, n42883, n42884, n42885, n42886,
         n42887, n42888, n42889, n42890, n42891, n42892, n42893, n42894,
         n42895, n42896, n42897, n42898, n42899, n42900, n42901, n42902,
         n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910,
         n42911, n42912, n42913, n42914, n42915, n42916, n42917, n42918,
         n42919, n42920, n42921, n42922, n42923, n42924, n42925, n42926,
         n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934,
         n42935, n42936, n42937, n42938, n42939, n42940, n42941, n42942,
         n42943, n42944, n42945, n42946, n42947, n42948, n42949, n42950,
         n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958,
         n42959, n42960, n42961, n42962, n42963, n42964, n42965, n42966,
         n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974,
         n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982,
         n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990,
         n42991, n42992, n42993, n42994, n42995, n42996, n42997, n42998,
         n42999, n43000, n43001, n43002, n43003, n43004, n43005, n43006,
         n43007, n43008, n43009, n43010, n43011, n43012, n43013, n43014,
         n43015, n43016, n43017, n43018, n43019, n43020, n43021, n43022,
         n43023, n43024, n43025, n43026, n43027, n43028, n43029, n43030,
         n43031, n43032, n43033, n43034, n43035, n43036, n43037, n43038,
         n43039, n43040, n43041, n43042, n43043, n43044, n43045, n43046,
         n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054,
         n43055, n43056, n43057, n43058, n43059, n43060, n43061, n43062,
         n43063, n43064, n43065, n43066, n43067, n43068, n43069, n43070,
         n43071, n43072, n43073, n43074, n43075, n43076, n43077, n43078,
         n43079, n43080, n43081, n43082, n43083, n43084, n43085, n43086,
         n43087, n43088, n43089, n43090, n43091, n43092, n43093, n43094,
         n43095, n43096, n43097, n43098, n43099, n43100, n43101, n43102,
         n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110,
         n43111, n43112, n43113, n43114, n43115, n43116, n43117, n43118,
         n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126,
         n43127, n43128, n43129, n43130, n43131, n43132, n43133, n43134,
         n43135, n43136, n43137, n43138, n43139, n43140, n43141, n43142,
         n43143, n43144, n43145, n43146, n43147, n43148, n43149, n43150,
         n43151, n43152, n43153, n43154, n43155, n43156, n43157, n43158,
         n43159, n43160, n43161, n43162, n43163, n43164, n43165, n43166,
         n43167, n43168, n43169, n43170, n43171, n43172, n43173, n43174,
         n43175, n43176, n43177, n43178, n43179, n43180, n43181, n43182,
         n43183, n43184, n43185, n43186, n43187, n43188, n43189, n43190,
         n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198,
         n43199, n43200, n43201, n43202, n43203, n43204, n43205, n43206,
         n43207, n43208, n43209, n43210, n43211, n43212, n43213, n43214,
         n43215, n43216, n43217, n43218, n43219, n43220, n43221, n43222,
         n43223, n43224, n43225, n43226, n43227, n43228, n43229, n43230,
         n43231, n43232, n43233, n43234, n43235, n43236, n43237, n43238,
         n43239, n43240, n43241, n43242, n43243, n43244, n43245, n43246,
         n43247, n43248, n43249, n43250, n43251, n43252, n43253, n43254,
         n43255, n43256, n43257, n43258, n43259, n43260, n43261, n43262,
         n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270,
         n43271, n43272, n43273, n43274, n43275, n43276, n43277, n43278,
         n43279, n43280, n43281, n43282, n43283, n43284, n43285, n43286,
         n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294,
         n43295, n43296, n43297, n43298, n43299, n43300, n43301, n43302,
         n43303, n43304, n43305, n43306, n43307, n43308, n43309, n43310,
         n43311, n43312, n43313, n43314, n43315, n43316, n43317, n43318,
         n43319, n43320, n43321, n43322, n43323, n43324, n43325, n43326,
         n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334,
         n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342,
         n43343, n43344, n43345, n43346, n43347, n43348, n43349, n43350,
         n43351, n43352, n43353, n43354, n43355, n43356, n43357, n43358,
         n43359, n43360, n43361, n43362, n43363, n43364, n43365, n43366,
         n43367, n43368, n43369, n43370, n43371, n43372, n43373, n43374,
         n43375, n43376, n43377, n43378, n43379, n43380, n43381, n43382,
         n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390,
         n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398,
         n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406,
         n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414,
         n43415, n43416, n43417, n43418, n43419, n43420, n43421, n43422,
         n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430,
         n43431, n43432, n43433, n43434, n43435, n43436, n43437, n43438,
         n43439, n43440, n43441, n43442, n43443, n43444, n43445, n43446,
         n43447, n43448, n43449, n43450, n43451, n43452, n43453, n43454,
         n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462,
         n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470,
         n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478,
         n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486,
         n43487, n43488, n43489, n43490, n43491, n43492, n43493, n43494,
         n43495, n43496, n43497, n43498, n43499, n43500, n43501, n43502,
         n43503, n43504, n43505, n43506, n43507, n43508, n43509, n43510,
         n43511, n43512, n43513, n43514, n43515, n43516, n43517, n43518,
         n43519, n43520, n43521, n43522, n43523, n43524, n43525, n43526,
         n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534,
         n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542,
         n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550,
         n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558,
         n43559, n43560, n43561, n43562, n43563, n43564, n43565, n43566,
         n43567, n43568, n43569, n43570, n43571, n43572, n43573, n43574,
         n43575, n43576, n43577, n43578, n43579, n43580, n43581, n43582,
         n43583, n43584, n43585, n43586, n43587, n43588, n43589, n43590,
         n43591, n43592, n43593, n43594, n43595, n43596, n43597, n43598,
         n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606,
         n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614,
         n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622,
         n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630,
         n43631, n43632, n43633, n43634, n43635, n43636, n43637, n43638,
         n43639, n43640, n43641, n43642, n43643, n43644, n43645, n43646,
         n43647, n43648, n43649, n43650, n43651, n43652, n43653, n43654,
         n43655, n43656, n43657, n43658, n43659, n43660, n43661, n43662,
         n43663, n43664, n43665, n43666, n43667, n43668, n43669, n43670,
         n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678,
         n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686,
         n43687, n43688, n43689, n43690, n43691, n43692, n43693, n43694,
         n43695, n43696, n43697, n43698, n43699, n43700, n43701, n43702,
         n43703, n43704, n43705, n43706, n43707, n43708, n43709, n43710,
         n43711, n43712, n43713, n43714, n43715, n43716, n43717, n43718,
         n43719, n43720, n43721, n43722, n43723, n43724, n43725, n43726,
         n43727, n43728, n43729, n43730, n43731, n43732, n43733, n43734,
         n43735, n43736, n43737, n43738, n43739, n43740, n43741, n43742,
         n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750,
         n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758,
         n43759, n43760, n43761, n43762, n43763, n43764, n43765, n43766,
         n43767, n43768, n43769, n43770, n43771, n43772, n43773, n43774,
         n43775, n43776, n43777, n43778, n43779, n43780, n43781, n43782,
         n43783, n43784, n43785, n43786, n43787, n43788, n43789, n43790,
         n43791, n43792, n43793, n43794, n43795, n43796, n43797, n43798,
         n43799, n43800, n43801, n43802, n43803, n43804, n43805, n43806,
         n43807, n43808, n43809, n43810, n43811, n43812, n43813, n43814,
         n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822,
         n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830,
         n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838,
         n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846,
         n43847, n43848, n43849, n43850, n43851, n43852, n43853, n43854,
         n43855, n43856, n43857, n43858, n43859, n43860, n43861, n43862,
         n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870,
         n43871, n43872, n43873, n43874, n43875, n43876, n43877, n43878,
         n43879, n43880, n43881, n43882, n43883, n43884, n43885, n43886,
         n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894,
         n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902,
         n43903, n43904, n43905, n43906, n43907, n43908, n43909, n43910,
         n43911, n43912, n43913, n43914, n43915, n43916, n43917, n43918,
         n43919, n43920, n43921, n43922, n43923, n43924, n43925, n43926,
         n43927, n43928, n43929, n43930, n43931, n43932, n43933, n43934,
         n43935, n43936, n43937, n43938, n43939, n43940, n43941, n43942,
         n43943, n43944, n43945, n43946, n43947, n43948, n43949, n43950,
         n43951, n43952, n43953, n43954, n43955, n43956, n43957, n43958,
         n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966,
         n43967, n43968, n43969, n43970, n43971, n43972, n43973, n43974,
         n43975, n43976, n43977, n43978, n43979, n43980, n43981, n43982,
         n43983, n43984, n43985, n43986, n43987, n43988, n43989, n43990,
         n43991, n43992, n43993, n43994, n43995, n43996, n43997, n43998,
         n43999, n44000, n44001, n44002, n44003, n44004, n44005, n44006,
         n44007, n44008, n44009, n44010, n44011, n44012, n44013, n44014,
         n44015, n44016, n44017, n44018, n44019, n44020, n44021, n44022,
         n44023, n44024, n44025, n44026, n44027, n44028, n44029, n44030,
         n44031, n44032, n44033, n44034, n44035, n44036, n44037, n44038,
         n44039, n44040, n44041, n44042, n44043, n44044, n44045, n44046,
         n44047, n44048, n44049, n44050, n44051, n44052, n44053, n44054,
         n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062,
         n44063, n44064, n44065, n44066, n44067, n44068, n44069, n44070,
         n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078,
         n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086,
         n44087, n44088, n44089, n44090, n44091, n44092, n44093, n44094,
         n44095, n44096, n44097, n44098, n44099, n44100, n44101, n44102,
         n44103, n44104, n44105, n44106, n44107, n44108, n44109, n44110,
         n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118,
         n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126,
         n44127, n44128, n44129, n44130, n44131, n44132, n44133, n44134,
         n44135, n44136, n44137, n44138, n44139, n44140, n44141, n44142,
         n44143, n44144, n44145, n44146, n44147, n44148, n44149, n44150,
         n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158,
         n44159, n44160, n44161, n44162, n44163, n44164, n44165, n44166,
         n44167, n44168, n44169, n44170, n44171, n44172, n44173, n44174,
         n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182,
         n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190,
         n44191, n44192, n44193, n44194, n44195, n44196, n44197, n44198,
         n44199, n44200, n44201, n44202, n44203, n44204, n44205, n44206,
         n44207, n44208, n44209, n44210, n44211, n44212, n44213, n44214,
         n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222,
         n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230,
         n44231, n44232, n44233, n44234, n44235, n44236, n44237, n44238,
         n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246,
         n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254,
         n44255, n44256, n44257, n44258, n44259, n44260, n44261, n44262,
         n44263, n44264, n44265, n44266, n44267, n44268, n44269, n44270,
         n44271, n44272, n44273, n44274, n44275, n44276, n44277, n44278,
         n44279, n44280, n44281, n44282, n44283, n44284, n44285, n44286,
         n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294,
         n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302,
         n44303, n44304, n44305, n44306, n44307, n44308, n44309, n44310,
         n44311, n44312, n44313, n44314, n44315, n44316, n44317, n44318,
         n44319, n44320, n44321, n44322, n44323, n44324, n44325, n44326,
         n44327, n44328, n44329, n44330, n44331, n44332, n44333, n44334,
         n44335, n44336, n44337, n44338, n44339, n44340, n44341, n44342,
         n44343, n44344, n44345, n44346, n44347, n44348, n44349, n44350,
         n44351, n44352, n44353, n44354, n44355, n44356, n44357, n44358,
         n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366,
         n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374,
         n44375, n44376, n44377, n44378, n44379, n44380, n44381, n44382,
         n44383, n44384, n44385, n44386, n44387, n44388, n44389, n44390,
         n44391, n44392, n44393, n44394, n44395, n44396, n44397, n44398,
         n44399, n44400, n44401, n44402, n44403, n44404, n44405, n44406,
         n44407, n44408, n44409, n44410, n44411, n44412, n44413, n44414,
         n44415, n44416, n44417, n44418, n44419, n44420, n44421, n44422,
         n44423, n44424, n44425, n44426, n44427, n44428, n44429, n44430,
         n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438,
         n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446,
         n44447, n44448, n44449, n44450, n44451, n44452, n44453, n44454,
         n44455, n44456, n44457, n44458, n44459, n44460, n44461, n44462,
         n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470,
         n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478,
         n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486,
         n44487, n44488, n44489, n44490, n44491, n44492, n44493, n44494,
         n44495, n44496, n44497, n44498, n44499, n44500, n44501, n44502,
         n44503, n44504, n44505, n44506, n44507, n44508, n44509, n44510,
         n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518,
         n44519, n44520, n44521, n44522, n44523, n44524, n44525, n44526,
         n44527, n44528, n44529, n44530, n44531, n44532, n44533, n44534,
         n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542,
         n44543, n44544, n44545, n44546, n44547, n44548, n44549, n44550,
         n44551, n44552, n44553, n44554, n44555, n44556, n44557, n44558,
         n44559, n44560, n44561, n44562, n44563, n44564, n44565, n44566,
         n44567, n44568, n44569, n44570, n44571, n44572, n44573, n44574,
         n44575, n44576, n44577, n44578, n44579, n44580, n44581, n44582,
         n44583, n44584, n44585, n44586, n44587, n44588, n44589, n44590,
         n44591, n44592, n44593, n44594, n44595, n44596, n44597, n44598,
         n44599, n44600, n44601, n44602, n44603, n44604, n44605, n44606,
         n44607, n44608, n44609, n44610, n44611, n44612, n44613, n44614,
         n44615, n44616, n44617, n44618, n44619, n44620, n44621, n44622,
         n44623, n44624, n44625, n44626, n44627, n44628, n44629, n44630,
         n44631, n44632, n44633, n44634, n44635, n44636, n44637, n44638,
         n44639, n44640, n44641, n44642, n44643, n44644, n44645, n44646,
         n44647, n44648, n44649, n44650, n44651, n44652, n44653, n44654,
         n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662,
         n44663, n44664, n44665, n44666, n44667, n44668, n44669, n44670,
         n44671, n44672, n44673, n44674, n44675, n44676, n44677, n44678,
         n44679, n44680, n44681, n44682, n44683, n44684, n44685, n44686,
         n44687, n44688, n44689, n44690, n44691, n44692, n44693, n44694,
         n44695, n44696, n44697, n44698, n44699, n44700, n44701, n44702,
         n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710,
         n44711, n44712, n44713, n44714, n44715, n44716, n44717, n44718,
         n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726,
         n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734,
         n44735, n44736, n44737, n44738, n44739, n44740, n44741, n44742,
         n44743, n44744, n44745, n44746, n44747, n44748, n44749, n44750,
         n44751, n44752, n44753, n44754, n44755, n44756, n44757, n44758,
         n44759, n44760, n44761, n44762, n44763, n44764, n44765, n44766,
         n44767, n44768, n44769, n44770, n44771, n44772, n44773, n44774,
         n44775, n44776, n44777, n44778, n44779, n44780, n44781, n44782,
         n44783, n44784, n44785, n44786, n44787, n44788, n44789, n44790,
         n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798,
         n44799, n44800, n44801, n44802, n44803, n44804, n44805, n44806,
         n44807, n44808, n44809, n44810, n44811, n44812, n44813, n44814,
         n44815, n44816, n44817, n44818, n44819, n44820, n44821, n44822,
         n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830,
         n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838,
         n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846,
         n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854,
         n44855, n44856, n44857, n44858, n44859, n44860, n44861, n44862,
         n44863, n44864, n44865, n44866, n44867, n44868, n44869, n44870,
         n44871, n44872, n44873, n44874, n44875, n44876, n44877, n44878,
         n44879, n44880, n44881, n44882, n44883, n44884, n44885, n44886,
         n44887, n44888, n44889, n44890, n44891, n44892, n44893, n44894,
         n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902,
         n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910,
         n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918,
         n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926,
         n44927, n44928, n44929, n44930, n44931, n44932, n44933, n44934,
         n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942,
         n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950,
         n44951, n44952, n44953, n44954, n44955, n44956, n44957, n44958,
         n44959, n44960, n44961, n44962, n44963, n44964, n44965, n44966,
         n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974,
         n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982,
         n44983, n44984, n44985, n44986, n44987, n44988, n44989, n44990,
         n44991, n44992, n44993, n44994, n44995, n44996, n44997, n44998,
         n44999, n45000, n45001, n45002, n45003, n45004, n45005, n45006,
         n45007, n45008, n45009, n45010, n45011, n45012, n45013, n45014,
         n45015, n45016, n45017, n45018, n45019, n45020, n45021, n45022,
         n45023, n45024, n45025, n45026, n45027, n45028, n45029, n45030,
         n45031, n45032, n45033, n45034, n45035, n45036, n45037, n45038,
         n45039, n45040, n45041, n45042, n45043, n45044, n45045, n45046,
         n45047, n45048, n45049, n45050, n45051, n45052, n45053, n45054,
         n45055, n45056, n45057, n45058, n45059, n45060, n45061, n45062,
         n45063, n45064, n45065, n45066, n45067, n45068, n45069, n45070,
         n45071, n45072, n45073, n45074, n45075, n45076, n45077, n45078,
         n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086,
         n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094,
         n45095, n45096, n45097, n45098, n45099, n45100, n45101, n45102,
         n45103, n45104, n45105, n45106, n45107, n45108, n45109, n45110,
         n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118,
         n45119, n45120, n45121, n45122, n45123, n45124, n45125, n45126,
         n45127, n45128, n45129, n45130, n45131, n45132, n45133, n45134,
         n45135, n45136, n45137, n45138, n45139, n45140, n45141, n45142,
         n45143, n45144, n45145, n45146, n45147, n45148, n45149, n45150,
         n45151, n45152, n45153, n45154, n45155, n45156, n45157, n45158,
         n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166,
         n45167, n45168, n45169, n45170, n45171, n45172, n45173, n45174,
         n45175, n45176, n45177, n45178, n45179, n45180, n45181, n45182,
         n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190,
         n45191, n45192, n45193, n45194, n45195, n45196, n45197, n45198,
         n45199, n45200, n45201, n45202, n45203, n45204, n45205, n45206,
         n45207, n45208, n45209, n45210, n45211, n45212, n45213, n45214,
         n45215, n45216, n45217, n45218, n45219, n45220, n45221, n45222,
         n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230,
         n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238,
         n45239, n45240, n45241, n45242, n45243, n45244, n45245, n45246,
         n45247, n45248, n45249, n45250, n45251, n45252, n45253, n45254,
         n45255, n45256, n45257, n45258, n45259, n45260, n45261, n45262,
         n45263, n45264, n45265, n45266, n45267, n45268, n45269, n45270,
         n45271, n45272, n45273, n45274, n45275, n45276, n45277, n45278,
         n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286,
         n45287, n45288, n45289, n45290, n45291, n45292, n45293, n45294,
         n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302,
         n45303, n45304, n45305, n45306, n45307, n45308, n45309, n45310,
         n45311, n45312, n45313, n45314, n45315, n45316, n45317, n45318,
         n45319, n45320, n45321, n45322, n45323, n45324, n45325, n45326,
         n45327, n45328, n45329, n45330, n45331, n45332, n45333, n45334,
         n45335, n45336, n45337, n45338, n45339, n45340, n45341, n45342,
         n45343, n45344, n45345, n45346, n45347, n45348, n45349, n45350,
         n45351, n45352, n45353, n45354, n45355, n45356, n45357, n45358,
         n45359, n45360, n45361, n45362, n45363, n45364, n45365, n45366,
         n45367, n45368, n45369, n45370, n45371, n45372, n45373, n45374,
         n45375, n45376, n45377, n45378, n45379, n45380, n45381, n45382,
         n45383, n45384, n45385, n45386, n45387, n45388, n45389, n45390,
         n45391, n45392, n45393, n45394, n45395, n45396, n45397, n45398,
         n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406,
         n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414,
         n45415, n45416, n45417, n45418, n45419, n45420, n45421, n45422,
         n45423, n45424, n45425, n45426, n45427, n45428, n45429, n45430,
         n45431, n45432, n45433, n45434, n45435, n45436, n45437, n45438,
         n45439, n45440, n45441, n45442, n45443, n45444, n45445, n45446,
         n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454,
         n45455, n45456, n45457, n45458, n45459, n45460, n45461, n45462,
         n45463, n45464, n45465, n45466, n45467, n45468, n45469, n45470,
         n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478,
         n45479, n45480, n45481, n45482, n45483, n45484, n45485, n45486,
         n45487, n45488, n45489, n45490, n45491, n45492, n45493, n45494,
         n45495, n45496, n45497, n45498, n45499, n45500, n45501, n45502,
         n45503, n45504, n45505, n45506, n45507, n45508, n45509, n45510,
         n45511, n45512, n45513, n45514, n45515, n45516, n45517, n45518,
         n45519, n45520, n45521, n45522, n45523, n45524, n45525, n45526,
         n45527, n45528, n45529, n45530, n45531, n45532, n45533, n45534,
         n45535, n45536, n45537, n45538, n45539, n45540, n45541, n45542,
         n45543, n45544, n45545, n45546, n45547, n45548, n45549, n45550,
         n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558,
         n45559, n45560, n45561, n45562, n45563, n45564, n45565, n45566,
         n45567, n45568, n45569, n45570, n45571, n45572, n45573, n45574,
         n45575, n45576, n45577, n45578, n45579, n45580, n45581, n45582,
         n45583, n45584, n45585, n45586, n45587, n45588, n45589, n45590,
         n45591, n45592, n45593, n45594, n45595, n45596, n45597, n45598,
         n45599, n45600, n45601, n45602, n45603, n45604, n45605, n45606,
         n45607, n45608, n45609, n45610, n45611, n45612, n45613, n45614,
         n45615, n45616, n45617, n45618, n45619, n45620, n45621, n45622,
         n45623, n45624, n45625, n45626, n45627, n45628, n45629, n45630,
         n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638,
         n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646,
         n45647, n45648, n45649, n45650, n45651, n45652, n45653, n45654,
         n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662,
         n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670,
         n45671, n45672, n45673, n45674, n45675, n45676, n45677, n45678,
         n45679, n45680, n45681, n45682, n45683, n45684, n45685, n45686,
         n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694,
         n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702,
         n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710,
         n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718,
         n45719, n45720, n45721, n45722, n45723, n45724, n45725, n45726,
         n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734,
         n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742,
         n45743, n45744, n45745, n45746, n45747, n45748, n45749, n45750,
         n45751, n45752, n45753, n45754, n45755, n45756, n45757, n45758,
         n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766,
         n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774,
         n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782,
         n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790,
         n45791, n45792, n45793, n45794, n45795, n45796, n45797, n45798,
         n45799, n45800, n45801, n45802, n45803, n45804, n45805, n45806,
         n45807, n45808, n45809, n45810, n45811, n45812, n45813, n45814,
         n45815, n45816, n45817, n45818, n45819, n45820, n45821, n45822,
         n45823, n45824, n45825, n45826, n45827, n45828, n45829, n45830,
         n45831, n45832, n45833, n45834, n45835, n45836, n45837, n45838,
         n45839, n45840, n45841, n45842, n45843, n45844, n45845, n45846,
         n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854,
         n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862,
         n45863, n45864, n45865, n45866, n45867, n45868, n45869, n45870,
         n45871, n45872, n45873, n45874, n45875, n45876, n45877, n45878,
         n45879, n45880, n45881, n45882, n45883, n45884, n45885, n45886,
         n45887, n45888, n45889, n45890, n45891, n45892, n45893, n45894,
         n45895, n45896, n45897, n45898, n45899, n45900, n45901, n45902,
         n45903, n45904, n45905, n45906, n45907, n45908, n45909, n45910,
         n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918,
         n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926,
         n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934,
         n45935, n45936, n45937, n45938, n45939, n45940, n45941, n45942,
         n45943, n45944, n45945, n45946, n45947, n45948, n45949, n45950,
         n45951, n45952, n45953, n45954, n45955, n45956, n45957, n45958,
         n45959, n45960, n45961, n45962, n45963, n45964, n45965, n45966,
         n45967, n45968, n45969, n45970, n45971, n45972, n45973, n45974,
         n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982,
         n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990,
         n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998,
         n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006,
         n46007, n46008, n46009, n46010, n46011, n46012, n46013, n46014,
         n46015, n46016, n46017, n46018, n46019, n46020, n46021, n46022,
         n46023, n46024, n46025, n46026, n46027, n46028, n46029, n46030,
         n46031, n46032, n46033, n46034, n46035, n46036, n46037, n46038,
         n46039, n46040, n46041, n46042, n46043, n46044, n46045, n46046,
         n46047, n46048, n46049, n46050, n46051, n46052, n46053, n46054,
         n46055, n46056, n46057, n46058, n46059, n46060, n46061, n46062,
         n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070,
         n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078,
         n46079, n46080, n46081, n46082, n46083, n46084, n46085, n46086,
         n46087, n46088, n46089, n46090, n46091, n46092, n46093, n46094,
         n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102,
         n46103, n46104, n46105, n46106, n46107, n46108, n46109, n46110,
         n46111, n46112, n46113, n46114, n46115, n46116, n46117, n46118,
         n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126,
         n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134,
         n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142,
         n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150,
         n46151, n46152, n46153, n46154, n46155, n46156, n46157, n46158,
         n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166,
         n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174,
         n46175, n46176, n46177, n46178, n46179, n46180, n46181, n46182,
         n46183, n46184, n46185, n46186, n46187, n46188, n46189, n46190,
         n46191, n46192, n46193, n46194, n46195, n46196, n46197, n46198,
         n46199, n46200, n46201, n46202, n46203, n46204, n46205, n46206,
         n46207, n46208, n46209, n46210, n46211, n46212, n46213, n46214,
         n46215, n46216, n46217, n46218, n46219, n46220, n46221, n46222,
         n46223, n46224, n46225, n46226, n46227, n46228, n46229, n46230,
         n46231, n46232, n46233, n46234, n46235, n46236, n46237, n46238,
         n46239, n46240, n46241, n46242, n46243, n46244, n46245, n46246,
         n46247, n46248, n46249, n46250, n46251, n46252, n46253, n46254,
         n46255, n46256, n46257, n46258, n46259, n46260, n46261, n46262,
         n46263, n46264, n46265, n46266, n46267, n46268, n46269, n46270,
         n46271, n46272, n46273, n46274, n46275, n46276, n46277, n46278,
         n46279, n46280, n46281, n46282, n46283, n46284, n46285, n46286,
         n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294,
         n46295, n46296, n46297, n46298, n46299, n46300, n46301, n46302,
         n46303, n46304, n46305, n46306, n46307, n46308, n46309, n46310,
         n46311, n46312, n46313, n46314, n46315, n46316, n46317, n46318,
         n46319, n46320, n46321, n46322, n46323, n46324, n46325, n46326,
         n46327, n46328, n46329, n46330, n46331, n46332, n46333, n46334,
         n46335, n46336, n46337, n46338, n46339, n46340, n46341, n46342,
         n46343, n46344, n46345, n46346, n46347, n46348, n46349, n46350,
         n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358,
         n46359, n46360, n46361, n46362, n46363, n46364, n46365, n46366,
         n46367, n46368, n46369, n46370, n46371, n46372, n46373, n46374,
         n46375, n46376, n46377, n46378, n46379, n46380, n46381, n46382,
         n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46390,
         n46391, n46392, n46393, n46394, n46395, n46396, n46397, n46398,
         n46399, n46400, n46401, n46402, n46403, n46404, n46405, n46406,
         n46407, n46408, n46409, n46410, n46411, n46412, n46413, n46414,
         n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422,
         n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430,
         n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438,
         n46439, n46440, n46441, n46442, n46443, n46444, n46445, n46446,
         n46447, n46448, n46449, n46450, n46451, n46452, n46453, n46454,
         n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462,
         n46463, n46464, n46465, n46466, n46467, n46468, n46469, n46470,
         n46471, n46472, n46473, n46474, n46475, n46476, n46477, n46478,
         n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486,
         n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494,
         n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502,
         n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510,
         n46511, n46512, n46513, n46514, n46515, n46516, n46517, n46518,
         n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526,
         n46527, n46528, n46529, n46530, n46531, n46532, n46533, n46534,
         n46535, n46536, n46537, n46538, n46539, n46540, n46541, n46542,
         n46543, n46544, n46545, n46546, n46547, n46548, n46549, n46550,
         n46551, n46552, n46553, n46554, n46555, n46556, n46557, n46558,
         n46559, n46560, n46561, n46562, n46563, n46564, n46565, n46566,
         n46567, n46568, n46569, n46570, n46571, n46572, n46573, n46574,
         n46575, n46576, n46577, n46578, n46579, n46580, n46581, n46582,
         n46583, n46584, n46585, n46586, n46587, n46588, n46589, n46590,
         n46591, n46592, n46593, n46594, n46595, n46596, n46597, n46598,
         n46599, n46600, n46601, n46602, n46603, n46604, n46605, n46606,
         n46607, n46608, n46609, n46610, n46611, n46612, n46613, n46614,
         n46615, n46616, n46617, n46618, n46619, n46620, n46621, n46622,
         n46623, n46624, n46625, n46626, n46627, n46628, n46629, n46630,
         n46631, n46632, n46633, n46634, n46635, n46636, n46637, n46638,
         n46639, n46640, n46641, n46642, n46643, n46644, n46645, n46646,
         n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654,
         n46655, n46656, n46657, n46658, n46659, n46660, n46661, n46662,
         n46663, n46664, n46665, n46666, n46667, n46668, n46669, n46670,
         n46671, n46672, n46673, n46674, n46675, n46676, n46677, n46678,
         n46679, n46680, n46681, n46682, n46683, n46684, n46685, n46686,
         n46687, n46688, n46689, n46690, n46691, n46692, n46693, n46694,
         n46695, n46696, n46697, n46698, n46699, n46700, n46701, n46702,
         n46703, n46704, n46705, n46706, n46707, n46708, n46709, n46710,
         n46711, n46712, n46713, n46714, n46715, n46716, n46717, n46718,
         n46719, n46720, n46721, n46722, n46723, n46724, n46725, n46726,
         n46727, n46728, n46729, n46730, n46731, n46732, n46733, n46734,
         n46735, n46736, n46737, n46738, n46739, n46740, n46741, n46742,
         n46743, n46744, n46745, n46746, n46747, n46748, n46749, n46750,
         n46751, n46752, n46753, n46754, n46755, n46756, n46757, n46758,
         n46759, n46760, n46761, n46762, n46763, n46764, n46765, n46766,
         n46767, n46768, n46769, n46770, n46771, n46772, n46773, n46774,
         n46775, n46776, n46777, n46778, n46779, n46780, n46781, n46782,
         n46783, n46784, n46785, n46786, n46787, n46788, n46789, n46790,
         n46791, n46792, n46793, n46794, n46795, n46796, n46797, n46798,
         n46799, n46800, n46801, n46802, n46803, n46804, n46805, n46806,
         n46807, n46808, n46809, n46810, n46811, n46812, n46813, n46814,
         n46815, n46816, n46817, n46818, n46819, n46820, n46821, n46822,
         n46823, n46824, n46825, n46826, n46827, n46828, n46829, n46830,
         n46831, n46832, n46833, n46834, n46835, n46836, n46837, n46838,
         n46839, n46840, n46841, n46842, n46843, n46844, n46845, n46846,
         n46847, n46848, n46849, n46850, n46851, n46852, n46853, n46854,
         n46855, n46856, n46857, n46858, n46859, n46860, n46861, n46862,
         n46863, n46864, n46865, n46866, n46867, n46868, n46869, n46870,
         n46871, n46872, n46873, n46874, n46875, n46876, n46877, n46878,
         n46879, n46880, n46881, n46882, n46883, n46884, n46885, n46886,
         n46887, n46888, n46889, n46890, n46891, n46892, n46893, n46894,
         n46895, n46896, n46897, n46898, n46899, n46900, n46901, n46902,
         n46903, n46904, n46905, n46906, n46907, n46908, n46909, n46910,
         n46911, n46912, n46913, n46914, n46915, n46916, n46917, n46918,
         n46919, n46920, n46921, n46922, n46923, n46924, n46925, n46926,
         n46927, n46928, n46929, n46930, n46931, n46932, n46933, n46934,
         n46935, n46936, n46937, n46938, n46939, n46940, n46941, n46942,
         n46943, n46944, n46945, n46946, n46947, n46948, n46949, n46950,
         n46951, n46952, n46953, n46954, n46955, n46956, n46957, n46958,
         n46959, n46960, n46961, n46962, n46963, n46964, n46965, n46966,
         n46967, n46968, n46969, n46970, n46971, n46972, n46973, n46974,
         n46975, n46976, n46977, n46978, n46979, n46980, n46981, n46982,
         n46983, n46984, n46985, n46986, n46987, n46988, n46989, n46990,
         n46991, n46992, n46993, n46994, n46995, n46996, n46997, n46998,
         n46999, n47000, n47001, n47002, n47003, n47004, n47005, n47006,
         n47007, n47008, n47009, n47010, n47011, n47012, n47013, n47014,
         n47015, n47016, n47017, n47018, n47019, n47020, n47021, n47022,
         n47023, n47024, n47025, n47026, n47027, n47028, n47029, n47030,
         n47031, n47032, n47033, n47034, n47035, n47036, n47037, n47038,
         n47039, n47040, n47041, n47042, n47043, n47044, n47045, n47046,
         n47047, n47048, n47049, n47050, n47051, n47052, n47053, n47054,
         n47055, n47056, n47057, n47058, n47059, n47060, n47061, n47062,
         n47063, n47064, n47065, n47066, n47067, n47068, n47069, n47070,
         n47071, n47072, n47073, n47074, n47075, n47076, n47077, n47078,
         n47079, n47080, n47081, n47082, n47083, n47084, n47085, n47086,
         n47087, n47088, n47089, n47090, n47091, n47092, n47093, n47094,
         n47095, n47096, n47097, n47098, n47099, n47100, n47101, n47102,
         n47103, n47104, n47105, n47106, n47107, n47108, n47109, n47110,
         n47111, n47112, n47113, n47114, n47115, n47116, n47117, n47118,
         n47119, n47120, n47121, n47122, n47123, n47124, n47125, n47126,
         n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134,
         n47135, n47136, n47137, n47138, n47139, n47140, n47141, n47142,
         n47143, n47144, n47145, n47146, n47147, n47148, n47149, n47150,
         n47151, n47152, n47153, n47154, n47155, n47156, n47157, n47158,
         n47159, n47160, n47161, n47162, n47163, n47164, n47165, n47166,
         n47167, n47168, n47169, n47170, n47171, n47172, n47173, n47174,
         n47175, n47176, n47177, n47178, n47179, n47180, n47181, n47182,
         n47183, n47184, n47185, n47186, n47187, n47188, n47189, n47190,
         n47191, n47192, n47193, n47194, n47195, n47196, n47197, n47198,
         n47199, n47200, n47201, n47202, n47203, n47204, n47205, n47206,
         n47207, n47208, n47209, n47210, n47211, n47212, n47213, n47214,
         n47215, n47216, n47217, n47218, n47219, n47220, n47221, n47222,
         n47223, n47224, n47225, n47226, n47227, n47228, n47229, n47230,
         n47231, n47232, n47233, n47234, n47235, n47236, n47237, n47238,
         n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246,
         n47247, n47248, n47249, n47250, n47251, n47252, n47253, n47254,
         n47255, n47256, n47257, n47258, n47259, n47260, n47261, n47262,
         n47263, n47264, n47265, n47266, n47267, n47268, n47269, n47270,
         n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278,
         n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286,
         n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294,
         n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302,
         n47303, n47304, n47305, n47306, n47307, n47308, n47309, n47310,
         n47311, n47312, n47313, n47314, n47315, n47316, n47317, n47318,
         n47319, n47320, n47321, n47322, n47323, n47324, n47325, n47326,
         n47327, n47328, n47329, n47330, n47331, n47332, n47333, n47334,
         n47335, n47336, n47337, n47338, n47339, n47340, n47341, n47342,
         n47343, n47344, n47345, n47346, n47347, n47348, n47349, n47350,
         n47351, n47352, n47353, n47354, n47355, n47356, n47357, n47358,
         n47359, n47360, n47361, n47362, n47363, n47364, n47365, n47366,
         n47367, n47368, n47369, n47370, n47371, n47372, n47373, n47374,
         n47375, n47376, n47377, n47378, n47379, n47380, n47381, n47382,
         n47383, n47384, n47385, n47386, n47387, n47388, n47389, n47390,
         n47391, n47392, n47393, n47394, n47395, n47396, n47397, n47398,
         n47399, n47400, n47401, n47402, n47403, n47404, n47405, n47406,
         n47407, n47408, n47409, n47410, n47411, n47412, n47413, n47414,
         n47415, n47416, n47417, n47418, n47419, n47420, n47421, n47422,
         n47423, n47424, n47425, n47426, n47427, n47428, n47429, n47430,
         n47431, n47432, n47433, n47434, n47435, n47436, n47437, n47438,
         n47439, n47440, n47441, n47442, n47443, n47444, n47445, n47446,
         n47447, n47448, n47449, n47450, n47451, n47452, n47453, n47454,
         n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462,
         n47463, n47464, n47465, n47466, n47467, n47468, n47469, n47470,
         n47471, n47472, n47473, n47474, n47475, n47476, n47477, n47478,
         n47479, n47480, n47481, n47482, n47483, n47484, n47485, n47486,
         n47487, n47488, n47489, n47490, n47491, n47492, n47493, n47494,
         n47495, n47496, n47497, n47498, n47499, n47500, n47501, n47502,
         n47503, n47504, n47505, n47506, n47507, n47508, n47509, n47510,
         n47511, n47512, n47513, n47514, n47515, n47516, n47517, n47518,
         n47519, n47520, n47521, n47522, n47523, n47524, n47525, n47526,
         n47527, n47528, n47529, n47530, n47531, n47532, n47533, n47534,
         n47535, n47536, n47537, n47538, n47539, n47540, n47541, n47542,
         n47543, n47544, n47545, n47546, n47547, n47548, n47549, n47550,
         n47551, n47552, n47553, n47554, n47555, n47556, n47557, n47558,
         n47559, n47560, n47561, n47562, n47563, n47564, n47565, n47566,
         n47567, n47568, n47569, n47570, n47571, n47572, n47573, n47574,
         n47575, n47576, n47577, n47578, n47579, n47580, n47581, n47582,
         n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590,
         n47591, n47592, n47593, n47594, n47595, n47596, n47597, n47598,
         n47599, n47600, n47601, n47602, n47603, n47604, n47605, n47606,
         n47607, n47608, n47609, n47610, n47611, n47612, n47613, n47614,
         n47615, n47616, n47617, n47618, n47619, n47620, n47621, n47622,
         n47623, n47624, n47625, n47626, n47627, n47628, n47629, n47630,
         n47631, n47632, n47633, n47634, n47635, n47636, n47637, n47638,
         n47639, n47640, n47641, n47642, n47643, n47644, n47645, n47646,
         n47647, n47648, n47649, n47650, n47651, n47652, n47653, n47654,
         n47655, n47656, n47657, n47658, n47659, n47660, n47661, n47662,
         n47663, n47664, n47665, n47666, n47667, n47668, n47669, n47670,
         n47671, n47672, n47673, n47674, n47675, n47676, n47677, n47678,
         n47679, n47680, n47681, n47682, n47683, n47684, n47685, n47686,
         n47687, n47688, n47689, n47690, n47691, n47692, n47693, n47694,
         n47695, n47696, n47697, n47698, n47699, n47700, n47701, n47702,
         n47703, n47704, n47705, n47706, n47707, n47708, n47709, n47710,
         n47711, n47712, n47713, n47714, n47715, n47716, n47717, n47718,
         n47719, n47720, n47721, n47722, n47723, n47724, n47725, n47726,
         n47727, n47728, n47729, n47730, n47731, n47732, n47733, n47734,
         n47735, n47736, n47737, n47738, n47739, n47740, n47741, n47742,
         n47743, n47744, n47745, n47746, n47747, n47748, n47749, n47750,
         n47751, n47752, n47753, n47754, n47755, n47756, n47757, n47758,
         n47759, n47760, n47761, n47762, n47763, n47764, n47765, n47766,
         n47767, n47768, n47769, n47770, n47771, n47772, n47773, n47774,
         n47775, n47776, n47777, n47778, n47779, n47780, n47781, n47782,
         n47783, n47784, n47785, n47786, n47787, n47788, n47789, n47790,
         n47791, n47792, n47793, n47794, n47795, n47796, n47797, n47798,
         n47799, n47800, n47801, n47802, n47803, n47804, n47805, n47806,
         n47807, n47808, n47809, n47810, n47811, n47812, n47813, n47814,
         n47815, n47816, n47817, n47818, n47819, n47820, n47821, n47822,
         n47823, n47824, n47825, n47826, n47827, n47828, n47829, n47830,
         n47831, n47832, n47833, n47834, n47835, n47836, n47837, n47838,
         n47839, n47840, n47841, n47842, n47843, n47844, n47845, n47846,
         n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854,
         n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862,
         n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870,
         n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878,
         n47879, n47880, n47881, n47882, n47883, n47884, n47885, n47886,
         n47887, n47888, n47889, n47890, n47891, n47892, n47893, n47894,
         n47895, n47896, n47897, n47898, n47899, n47900, n47901, n47902,
         n47903, n47904, n47905, n47906, n47907, n47908, n47909, n47910,
         n47911, n47912, n47913, n47914, n47915, n47916, n47917, n47918,
         n47919, n47920, n47921, n47922, n47923, n47924, n47925, n47926,
         n47927, n47928, n47929, n47930, n47931, n47932, n47933, n47934,
         n47935, n47936, n47937, n47938, n47939, n47940, n47941, n47942,
         n47943, n47944, n47945, n47946, n47947, n47948, n47949, n47950,
         n47951, n47952, n47953, n47954, n47955, n47956, n47957, n47958,
         n47959, n47960, n47961, n47962, n47963, n47964, n47965, n47966,
         n47967, n47968, n47969, n47970, n47971, n47972, n47973, n47974,
         n47975, n47976, n47977, n47978, n47979, n47980, n47981, n47982,
         n47983, n47984, n47985, n47986, n47987, n47988, n47989, n47990,
         n47991, n47992, n47993, n47994, n47995, n47996, n47997, n47998,
         n47999, n48000, n48001, n48002, n48003, n48004, n48005, n48006,
         n48007, n48008, n48009, n48010, n48011, n48012, n48013, n48014,
         n48015, n48016, n48017, n48018, n48019, n48020, n48021, n48022,
         n48023, n48024, n48025, n48026, n48027, n48028, n48029, n48030,
         n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038,
         n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046,
         n48047, n48048, n48049, n48050, n48051, n48052, n48053, n48054,
         n48055, n48056, n48057, n48058, n48059, n48060, n48061, n48062,
         n48063, n48064, n48065, n48066, n48067, n48068, n48069, n48070,
         n48071, n48072, n48073, n48074, n48075, n48076, n48077, n48078,
         n48079, n48080, n48081, n48082, n48083, n48084, n48085, n48086,
         n48087, n48088, n48089, n48090, n48091, n48092, n48093, n48094,
         n48095, n48096, n48097, n48098, n48099, n48100, n48101, n48102,
         n48103, n48104, n48105, n48106, n48107, n48108, n48109, n48110,
         n48111, n48112, n48113, n48114, n48115, n48116, n48117, n48118,
         n48119, n48120, n48121, n48122, n48123, n48124, n48125, n48126,
         n48127, n48128, n48129, n48130, n48131, n48132, n48133, n48134,
         n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142,
         n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150,
         n48151, n48152, n48153, n48154, n48155, n48156, n48157, n48158,
         n48159, n48160, n48161, n48162, n48163, n48164, n48165, n48166,
         n48167, n48168, n48169, n48170, n48171, n48172, n48173, n48174,
         n48175, n48176, n48177, n48178, n48179, n48180, n48181, n48182,
         n48183, n48184, n48185, n48186, n48187, n48188, n48189, n48190,
         n48191, n48192, n48193, n48194, n48195, n48196, n48197, n48198,
         n48199, n48200, n48201, n48202, n48203, n48204, n48205, n48206,
         n48207, n48208, n48209, n48210, n48211, n48212, n48213, n48214,
         n48215, n48216, n48217, n48218, n48219, n48220, n48221, n48222,
         n48223, n48224, n48225, n48226, n48227, n48228, n48229, n48230,
         n48231, n48232, n48233, n48234, n48235, n48236, n48237, n48238,
         n48239, n48240, n48241, n48242, n48243, n48244, n48245, n48246,
         n48247, n48248, n48249, n48250, n48251, n48252, n48253, n48254,
         n48255, n48256, n48257, n48258, n48259, n48260, n48261, n48262,
         n48263, n48264, n48265, n48266, n48267, n48268, n48269, n48270,
         n48271, n48272, n48273, n48274, n48275, n48276, n48277, n48278,
         n48279, n48280, n48281, n48282, n48283, n48284, n48285, n48286,
         n48287, n48288, n48289, n48290, n48291, n48292, n48293, n48294,
         n48295, n48296, n48297, n48298, n48299, n48300, n48301, n48302,
         n48303, n48304, n48305, n48306, n48307, n48308, n48309, n48310,
         n48311, n48312, n48313, n48314, n48315, n48316, n48317, n48318,
         n48319, n48320, n48321, n48322, n48323, n48324, n48325, n48326,
         n48327, n48328, n48329, n48330, n48331, n48332, n48333, n48334,
         n48335, n48336, n48337, n48338, n48339, n48340, n48341, n48342,
         n48343, n48344, n48345, n48346, n48347, n48348, n48349, n48350,
         n48351, n48352, n48353, n48354, n48355, n48356, n48357, n48358,
         n48359, n48360, n48361, n48362, n48363, n48364, n48365, n48366,
         n48367, n48368, n48369, n48370, n48371, n48372, n48373, n48374,
         n48375, n48376, n48377, n48378, n48379, n48380, n48381, n48382,
         n48383, n48384, n48385, n48386, n48387, n48388, n48389, n48390,
         n48391, n48392, n48393, n48394, n48395, n48396, n48397, n48398,
         n48399, n48400, n48401, n48402, n48403, n48404, n48405, n48406,
         n48407, n48408, n48409, n48410, n48411, n48412, n48413, n48414,
         n48415, n48416, n48417, n48418, n48419, n48420, n48421, n48422,
         n48423, n48424, n48425, n48426, n48427, n48428, n48429, n48430,
         n48431, n48432, n48433, n48434, n48435, n48436, n48437, n48438,
         n48439, n48440, n48441, n48442, n48443, n48444, n48445, n48446,
         n48447, n48448, n48449, n48450, n48451, n48452, n48453, n48454,
         n48455, n48456, n48457, n48458, n48459, n48460, n48461, n48462,
         n48463, n48464, n48465, n48466, n48467, n48468, n48469, n48470,
         n48471, n48472, n48473, n48474, n48475, n48476, n48477, n48478,
         n48479, n48480, n48481, n48482, n48483, n48484, n48485, n48486,
         n48487, n48488, n48489, n48490, n48491, n48492, n48493, n48494,
         n48495, n48496, n48497, n48498, n48499, n48500, n48501, n48502,
         n48503, n48504, n48505, n48506, n48507, n48508, n48509, n48510,
         n48511, n48512, n48513, n48514, n48515, n48516, n48517, n48518,
         n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526,
         n48527, n48528, n48529, n48530, n48531, n48532, n48533, n48534,
         n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542,
         n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550,
         n48551, n48552, n48553, n48554, n48555, n48556, n48557, n48558,
         n48559, n48560, n48561, n48562, n48563, n48564, n48565, n48566,
         n48567, n48568, n48569, n48570, n48571, n48572, n48573, n48574,
         n48575, n48576, n48577, n48578, n48579, n48580, n48581, n48582,
         n48583, n48584, n48585, n48586, n48587, n48588, n48589, n48590,
         n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598,
         n48599, n48600, n48601, n48602, n48603, n48604, n48605, n48606,
         n48607, n48608, n48609, n48610, n48611, n48612, n48613, n48614,
         n48615, n48616, n48617, n48618, n48619, n48620, n48621, n48622,
         n48623, n48624, n48625, n48626, n48627, n48628, n48629, n48630,
         n48631, n48632, n48633, n48634, n48635, n48636, n48637, n48638,
         n48639, n48640, n48641, n48642, n48643, n48644, n48645, n48646,
         n48647, n48648, n48649, n48650, n48651, n48652, n48653, n48654,
         n48655, n48656, n48657, n48658, n48659, n48660, n48661, n48662,
         n48663, n48664, n48665, n48666, n48667, n48668, n48669, n48670,
         n48671, n48672, n48673, n48674, n48675, n48676, n48677, n48678,
         n48679, n48680, n48681, n48682, n48683, n48684, n48685, n48686,
         n48687, n48688, n48689, n48690, n48691, n48692, n48693, n48694,
         n48695, n48696, n48697, n48698, n48699, n48700, n48701, n48702,
         n48703, n48704, n48705, n48706, n48707, n48708, n48709, n48710,
         n48711, n48712, n48713, n48714, n48715, n48716, n48717, n48718,
         n48719, n48720, n48721, n48722, n48723, n48724, n48725, n48726,
         n48727, n48728, n48729, n48730, n48731, n48732, n48733, n48734,
         n48735, n48736, n48737, n48738, n48739, n48740, n48741, n48742,
         n48743, n48744, n48745, n48746, n48747, n48748, n48749, n48750,
         n48751, n48752, n48753, n48754, n48755, n48756, n48757, n48758,
         n48759, n48760, n48761, n48762, n48763, n48764, n48765, n48766,
         n48767, n48768, n48769, n48770, n48771, n48772, n48773, n48774,
         n48775, n48776, n48777, n48778, n48779, n48780, n48781, n48782,
         n48783, n48784, n48785, n48786, n48787, n48788, n48789, n48790,
         n48791, n48792, n48793, n48794, n48795, n48796, n48797, n48798,
         n48799, n48800, n48801, n48802, n48803, n48804, n48805, n48806,
         n48807, n48808, n48809, n48810, n48811, n48812, n48813, n48814,
         n48815, n48816, n48817, n48818, n48819, n48820, n48821, n48822,
         n48823, n48824, n48825, n48826, n48827, n48828, n48829, n48830,
         n48831, n48832, n48833, n48834, n48835, n48836, n48837, n48838,
         n48839, n48840, n48841, n48842, n48843, n48844, n48845, n48846,
         n48847, n48848, n48849, n48850, n48851, n48852, n48853, n48854,
         n48855, n48856, n48857, n48858, n48859, n48860, n48861, n48862,
         n48863, n48864, n48865, n48866, n48867, n48868, n48869, n48870,
         n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878,
         n48879, n48880, n48881, n48882, n48883, n48884, n48885, n48886,
         n48887, n48888, n48889, n48890, n48891, n48892, n48893, n48894,
         n48895, n48896, n48897, n48898, n48899, n48900, n48901, n48902,
         n48903, n48904, n48905, n48906, n48907, n48908, n48909, n48910,
         n48911, n48912, n48913, n48914, n48915, n48916, n48917, n48918,
         n48919, n48920, n48921, n48922, n48923, n48924, n48925, n48926,
         n48927, n48928, n48929, n48930, n48931, n48932, n48933, n48934,
         n48935, n48936, n48937, n48938, n48939, n48940, n48941, n48942,
         n48943, n48944, n48945, n48946, n48947, n48948, n48949, n48950,
         n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958,
         n48959, n48960, n48961, n48962, n48963, n48964, n48965, n48966,
         n48967, n48968, n48969, n48970, n48971, n48972, n48973, n48974,
         n48975, n48976, n48977, n48978, n48979, n48980, n48981, n48982,
         n48983, n48984, n48985, n48986, n48987, n48988, n48989, n48990,
         n48991, n48992, n48993, n48994, n48995, n48996, n48997, n48998,
         n48999, n49000, n49001, n49002, n49003, n49004, n49005, n49006,
         n49007, n49008, n49009, n49010, n49011, n49012, n49013, n49014,
         n49015, n49016, n49017, n49018, n49019, n49020, n49021, n49022,
         n49023, n49024, n49025, n49026, n49027, n49028, n49029, n49030,
         n49031, n49032, n49033, n49034, n49035, n49036, n49037, n49038,
         n49039, n49040, n49041, n49042, n49043, n49044, n49045, n49046,
         n49047, n49048, n49049, n49050, n49051, n49052, n49053, n49054,
         n49055, n49056, n49057, n49058, n49059, n49060, n49061, n49062,
         n49063, n49064, n49065, n49066, n49067, n49068, n49069, n49070,
         n49071, n49072, n49073, n49074, n49075, n49076, n49077, n49078,
         n49079, n49080, n49081, n49082, n49083, n49084, n49085, n49086,
         n49087, n49088, n49089, n49090, n49091, n49092, n49093, n49094,
         n49095, n49096, n49097, n49098, n49099, n49100, n49101, n49102,
         n49103, n49104, n49105, n49106, n49107, n49108, n49109, n49110,
         n49111, n49112, n49113, n49114, n49115, n49116, n49117, n49118,
         n49119, n49120, n49121, n49122, n49123, n49124, n49125, n49126,
         n49127, n49128, n49129, n49130, n49131, n49132, n49133, n49134,
         n49135, n49136, n49137, n49138, n49139, n49140, n49141, n49142,
         n49143, n49144, n49145, n49146, n49147, n49148, n49149, n49150,
         n49151, n49152, n49153, n49154, n49155, n49156, n49157, n49158,
         n49159, n49160, n49161, n49162, n49163, n49164, n49165, n49166,
         n49167, n49168, n49169, n49170, n49171, n49172, n49173, n49174,
         n49175, n49176, n49177, n49178, n49179, n49180, n49181, n49182,
         n49183, n49184, n49185, n49186, n49187, n49188, n49189, n49190,
         n49191, n49192, n49193, n49194, n49195, n49196, n49197, n49198,
         n49199, n49200, n49201, n49202, n49203, n49204, n49205, n49206,
         n49207, n49208, n49209, n49210, n49211, n49212, n49213, n49214,
         n49215, n49216, n49217, n49218, n49219, n49220, n49221, n49222,
         n49223, n49224, n49225, n49226, n49227, n49228, n49229, n49230,
         n49231, n49232, n49233, n49234, n49235, n49236, n49237, n49238,
         n49239, n49240, n49241, n49242, n49243, n49244, n49245, n49246,
         n49247, n49248, n49249, n49250, n49251, n49252, n49253, n49254,
         n49255, n49256, n49257, n49258, n49259, n49260, n49261, n49262,
         n49263, n49264, n49265, n49266, n49267, n49268, n49269, n49270,
         n49271, n49272, n49273, n49274, n49275, n49276, n49277, n49278,
         n49279, n49280, n49281, n49282, n49283, n49284, n49285, n49286,
         n49287, n49288, n49289, n49290, n49291, n49292, n49293, n49294,
         n49295, n49296, n49297, n49298, n49299, n49300, n49301, n49302,
         n49303, n49304, n49305, n49306, n49307, n49308, n49309, n49310,
         n49311, n49312, n49313, n49314, n49315, n49316, n49317, n49318,
         n49319, n49320, n49321, n49322, n49323, n49324, n49325, n49326,
         n49327, n49328, n49329, n49330, n49331, n49332, n49333, n49334,
         n49335, n49336, n49337, n49338, n49339, n49340, n49341, n49342,
         n49343, n49344, n49345, n49346, n49347, n49348, n49349, n49350,
         n49351, n49352, n49353, n49354, n49355, n49356, n49357, n49358,
         n49359, n49360, n49361, n49362, n49363, n49364, n49365, n49366,
         n49367, n49368, n49369, n49370, n49371, n49372, n49373, n49374,
         n49375, n49376, n49377, n49378, n49379, n49380, n49381, n49382,
         n49383, n49384, n49385, n49386, n49387, n49388, n49389, n49390,
         n49391, n49392, n49393, n49394, n49395, n49396, n49397, n49398,
         n49399, n49400, n49401, n49402, n49403, n49404, n49405, n49406,
         n49407, n49408, n49409, n49410, n49411, n49412, n49413, n49414,
         n49415, n49416, n49417, n49418, n49419, n49420, n49421, n49422,
         n49423, n49424, n49425, n49426, n49427, n49428, n49429, n49430,
         n49431, n49432, n49433, n49434, n49435, n49436, n49437, n49438,
         n49439, n49440, n49441, n49442, n49443, n49444, n49445, n49446,
         n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454,
         n49455, n49456, n49457, n49458, n49459, n49460, n49461, n49462,
         n49463, n49464, n49465, n49466, n49467, n49468, n49469, n49470,
         n49471, n49472, n49473, n49474, n49475, n49476, n49477, n49478,
         n49479, n49480, n49481, n49482, n49483, n49484, n49485, n49486,
         n49487, n49488, n49489, n49490, n49491, n49492, n49493, n49494,
         n49495, n49496, n49497, n49498, n49499, n49500, n49501, n49502,
         n49503, n49504, n49505, n49506, n49507, n49508, n49509, n49510,
         n49511, n49512, n49513, n49514, n49515, n49516, n49517, n49518,
         n49519, n49520, n49521, n49522, n49523, n49524, n49525, n49526,
         n49527, n49528, n49529, n49530, n49531, n49532, n49533, n49534,
         n49535, n49536, n49537, n49538, n49539, n49540, n49541, n49542,
         n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550,
         n49551, n49552, n49553, n49554, n49555, n49556, n49557, n49558,
         n49559, n49560, n49561, n49562, n49563, n49564, n49565, n49566,
         n49567, n49568, n49569, n49570, n49571, n49572, n49573, n49574,
         n49575, n49576, n49577, n49578, n49579, n49580, n49581, n49582,
         n49583, n49584, n49585, n49586, n49587, n49588, n49589, n49590,
         n49591, n49592, n49593, n49594, n49595, n49596, n49597, n49598,
         n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606,
         n49607, n49608, n49609, n49610, n49611, n49612, n49613, n49614,
         n49615, n49616, n49617, n49618, n49619, n49620, n49621, n49622,
         n49623, n49624, n49625, n49626, n49627, n49628, n49629, n49630,
         n49631, n49632, n49633, n49634, n49635, n49636, n49637, n49638,
         n49639, n49640, n49641, n49642, n49643, n49644, n49645, n49646,
         n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654,
         n49655, n49656, n49657, n49658, n49659, n49660, n49661, n49662,
         n49663, n49664, n49665, n49666, n49667, n49668, n49669, n49670,
         n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678,
         n49679, n49680, n49681, n49682, n49683, n49684, n49685, n49686,
         n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694,
         n49695, n49696, n49697, n49698, n49699, n49700, n49701, n49702,
         n49703, n49704, n49705, n49706, n49707, n49708, n49709, n49710,
         n49711, n49712, n49713, n49714, n49715, n49716, n49717, n49718,
         n49719, n49720, n49721, n49722, n49723, n49724, n49725, n49726,
         n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734,
         n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742,
         n49743, n49744, n49745, n49746, n49747, n49748, n49749, n49750,
         n49751, n49752, n49753, n49754, n49755, n49756, n49757, n49758,
         n49759, n49760, n49761, n49762, n49763, n49764, n49765, n49766,
         n49767, n49768, n49769, n49770, n49771, n49772, n49773, n49774,
         n49775, n49776, n49777, n49778, n49779, n49780, n49781, n49782,
         n49783, n49784, n49785, n49786, n49787, n49788, n49789, n49790,
         n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798,
         n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806,
         n49807, n49808, n49809, n49810, n49811, n49812, n49813, n49814,
         n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822,
         n49823, n49824, n49825, n49826, n49827, n49828, n49829, n49830,
         n49831, n49832, n49833, n49834, n49835, n49836, n49837, n49838,
         n49839, n49840, n49841, n49842, n49843, n49844, n49845, n49846,
         n49847, n49848, n49849, n49850, n49851, n49852, n49853, n49854,
         n49855, n49856, n49857, n49858, n49859, n49860, n49861, n49862,
         n49863, n49864, n49865, n49866, n49867, n49868, n49869, n49870,
         n49871, n49872, n49873, n49874, n49875, n49876, n49877, n49878,
         n49879, n49880, n49881, n49882, n49883, n49884, n49885, n49886,
         n49887, n49888, n49889, n49890, n49891, n49892, n49893, n49894,
         n49895, n49896, n49897, n49898, n49899, n49900, n49901, n49902,
         n49903, n49904, n49905, n49906, n49907, n49908, n49909, n49910,
         n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918,
         n49919, n49920, n49921, n49922, n49923, n49924, n49925, n49926,
         n49927, n49928, n49929, n49930, n49931, n49932, n49933, n49934,
         n49935, n49936, n49937, n49938, n49939, n49940, n49941, n49942,
         n49943, n49944, n49945, n49946, n49947, n49948, n49949, n49950,
         n49951, n49952, n49953, n49954, n49955, n49956, n49957, n49958,
         n49959, n49960, n49961, n49962, n49963, n49964, n49965, n49966,
         n49967, n49968, n49969, n49970, n49971, n49972, n49973, n49974,
         n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982,
         n49983, n49984, n49985, n49986, n49987, n49988, n49989, n49990,
         n49991, n49992, n49993, n49994, n49995, n49996, n49997, n49998,
         n49999, n50000, n50001, n50002, n50003, n50004, n50005, n50006,
         n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014,
         n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022,
         n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030,
         n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038,
         n50039, n50040, n50041, n50042, n50043, n50044, n50045, n50046,
         n50047, n50048, n50049, n50050, n50051, n50052, n50053, n50054,
         n50055, n50056, n50057, n50058, n50059, n50060, n50061, n50062,
         n50063, n50064, n50065, n50066, n50067, n50068, n50069, n50070,
         n50071, n50072, n50073, n50074, n50075, n50076, n50077, n50078,
         n50079, n50080, n50081, n50082, n50083, n50084, n50085, n50086,
         n50087, n50088, n50089, n50090, n50091, n50092, n50093, n50094,
         n50095, n50096, n50097, n50098, n50099, n50100, n50101, n50102,
         n50103, n50104, n50105, n50106, n50107, n50108, n50109, n50110,
         n50111, n50112, n50113, n50114, n50115, n50116, n50117, n50118,
         n50119, n50120, n50121, n50122, n50123, n50124, n50125, n50126,
         n50127, n50128, n50129, n50130, n50131, n50132, n50133, n50134,
         n50135, n50136, n50137, n50138, n50139, n50140, n50141, n50142,
         n50143, n50144, n50145, n50146, n50147, n50148, n50149, n50150,
         n50151, n50152, n50153, n50154, n50155, n50156, n50157, n50158,
         n50159, n50160, n50161, n50162, n50163, n50164, n50165, n50166,
         n50167, n50168, n50169, n50170, n50171, n50172, n50173, n50174,
         n50175, n50176, n50177, n50178, n50179, n50180, n50181, n50182,
         n50183, n50184, n50185, n50186, n50187, n50188, n50189, n50190,
         n50191, n50192, n50193, n50194, n50195, n50196, n50197, n50198,
         n50199, n50200, n50201, n50202, n50203, n50204, n50205, n50206,
         n50207, n50208, n50209, n50210, n50211, n50212, n50213, n50214,
         n50215, n50216, n50217, n50218, n50219, n50220, n50221, n50222,
         n50223, n50224, n50225, n50226, n50227, n50228, n50229, n50230,
         n50231, n50232, n50233, n50234, n50235, n50236, n50237, n50238,
         n50239, n50240, n50241, n50242, n50243, n50244, n50245, n50246,
         n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254,
         n50255, n50256, n50257, n50258, n50259, n50260, n50261, n50262,
         n50263, n50264, n50265, n50266, n50267, n50268, n50269, n50270,
         n50271, n50272, n50273, n50274, n50275, n50276, n50277, n50278,
         n50279, n50280, n50281, n50282, n50283, n50284, n50285, n50286,
         n50287, n50288, n50289, n50290, n50291, n50292, n50293, n50294,
         n50295, n50296, n50297, n50298, n50299, n50300, n50301, n50302,
         n50303, n50304, n50305, n50306, n50307, n50308, n50309, n50310,
         n50311, n50312, n50313, n50314, n50315, n50316, n50317, n50318,
         n50319, n50320, n50321, n50322, n50323, n50324, n50325, n50326,
         n50327, n50328, n50329, n50330, n50331, n50332, n50333, n50334,
         n50335, n50336, n50337, n50338, n50339, n50340, n50341, n50342,
         n50343, n50344, n50345, n50346, n50347, n50348, n50349, n50350,
         n50351, n50352, n50353, n50354, n50355, n50356, n50357, n50358,
         n50359, n50360, n50361, n50362, n50363, n50364, n50365, n50366,
         n50367, n50368, n50369, n50370, n50371, n50372, n50373, n50374,
         n50375, n50376, n50377, n50378, n50379, n50380, n50381, n50382,
         n50383, n50384, n50385, n50386, n50387, n50388, n50389, n50390,
         n50391, n50392, n50393, n50394, n50395, n50396, n50397, n50398,
         n50399, n50400, n50401, n50402, n50403, n50404, n50405, n50406,
         n50407, n50408, n50409, n50410, n50411, n50412, n50413, n50414,
         n50415, n50416, n50417, n50418, n50419, n50420, n50421, n50422,
         n50423, n50424, n50425, n50426, n50427, n50428, n50429, n50430,
         n50431, n50432, n50433, n50434, n50435, n50436, n50437, n50438,
         n50439, n50440, n50441, n50442, n50443, n50444, n50445, n50446,
         n50447, n50448, n50449, n50450, n50451, n50452, n50453, n50454,
         n50455, n50456, n50457, n50458, n50459, n50460, n50461, n50462,
         n50463, n50464, n50465, n50466, n50467, n50468, n50469, n50470,
         n50471, n50472, n50473, n50474, n50475, n50476, n50477, n50478,
         n50479, n50480, n50481, n50482, n50483, n50484, n50485, n50486,
         n50487, n50488, n50489, n50490, n50491, n50492, n50493, n50494,
         n50495, n50496, n50497, n50498, n50499, n50500, n50501, n50502,
         n50503, n50504, n50505, n50506, n50507, n50508, n50509, n50510,
         n50511, n50512, n50513, n50514, n50515, n50516, n50517, n50518,
         n50519, n50520, n50521, n50522, n50523, n50524, n50525, n50526,
         n50527, n50528, n50529, n50530, n50531, n50532, n50533, n50534,
         n50535, n50536, n50537, n50538, n50539, n50540, n50541, n50542,
         n50543, n50544, n50545, n50546, n50547, n50548, n50549, n50550,
         n50551, n50552, n50553, n50554, n50555, n50556, n50557, n50558,
         n50559, n50560, n50561, n50562, n50563, n50564, n50565, n50566,
         n50567, n50568, n50569, n50570, n50571, n50572, n50573, n50574,
         n50575, n50576, n50577, n50578, n50579, n50580, n50581, n50582,
         n50583, n50584, n50585, n50586, n50587, n50588, n50589, n50590,
         n50591, n50592, n50593, n50594, n50595, n50596, n50597, n50598,
         n50599, n50600, n50601, n50602, n50603, n50604, n50605, n50606,
         n50607, n50608, n50609, n50610, n50611, n50612, n50613, n50614,
         n50615, n50616, n50617, n50618, n50619, n50620, n50621, n50622,
         n50623, n50624, n50625, n50626, n50627, n50628, n50629, n50630,
         n50631, n50632, n50633, n50634, n50635, n50636, n50637, n50638,
         n50639, n50640, n50641, n50642, n50643, n50644, n50645, n50646,
         n50647, n50648, n50649, n50650, n50651, n50652, n50653, n50654,
         n50655, n50656, n50657, n50658, n50659, n50660, n50661, n50662,
         n50663, n50664, n50665, n50666, n50667, n50668, n50669, n50670,
         n50671, n50672, n50673, n50674, n50675, n50676, n50677, n50678,
         n50679, n50680, n50681, n50682, n50683, n50684, n50685, n50686,
         n50687, n50688, n50689, n50690, n50691, n50692, n50693, n50694,
         n50695, n50696, n50697, n50698, n50699, n50700, n50701, n50702,
         n50703, n50704, n50705, n50706, n50707, n50708, n50709, n50710,
         n50711, n50712, n50713, n50714, n50715, n50716, n50717, n50718,
         n50719, n50720, n50721, n50722, n50723, n50724, n50725, n50726,
         n50727, n50728, n50729, n50730, n50731, n50732, n50733, n50734,
         n50735, n50736, n50737, n50738, n50739, n50740, n50741, n50742,
         n50743, n50744, n50745, n50746, n50747, n50748, n50749, n50750,
         n50751, n50752, n50753, n50754, n50755, n50756, n50757, n50758,
         n50759, n50760, n50761, n50762, n50763, n50764, n50765, n50766,
         n50767, n50768, n50769, n50770, n50771, n50772, n50773, n50774,
         n50775, n50776, n50777, n50778, n50779, n50780, n50781, n50782,
         n50783, n50784, n50785, n50786, n50787, n50788, n50789, n50790,
         n50791, n50792, n50793, n50794, n50795, n50796, n50797, n50798,
         n50799, n50800, n50801, n50802, n50803, n50804, n50805, n50806,
         n50807, n50808, n50809, n50810, n50811, n50812, n50813, n50814,
         n50815, n50816, n50817, n50818, n50819, n50820, n50821, n50822,
         n50823, n50824, n50825, n50826, n50827, n50828, n50829, n50830,
         n50831, n50832, n50833, n50834, n50835, n50836, n50837, n50838,
         n50839, n50840, n50841, n50842, n50843, n50844, n50845, n50846,
         n50847, n50848, n50849, n50850, n50851, n50852, n50853, n50854,
         n50855, n50856, n50857, n50858, n50859, n50860, n50861, n50862,
         n50863, n50864, n50865, n50866, n50867, n50868, n50869, n50870,
         n50871, n50872, n50873, n50874, n50875, n50876, n50877, n50878,
         n50879, n50880, n50881, n50882, n50883, n50884, n50885, n50886,
         n50887, n50888, n50889, n50890, n50891, n50892, n50893, n50894,
         n50895, n50896, n50897, n50898, n50899, n50900, n50901, n50902,
         n50903, n50904, n50905, n50906, n50907, n50908, n50909, n50910,
         n50911, n50912, n50913, n50914, n50915, n50916, n50917, n50918,
         n50919, n50920, n50921, n50922, n50923, n50924, n50925, n50926,
         n50927, n50928, n50929, n50930, n50931, n50932, n50933, n50934,
         n50935, n50936, n50937, n50938, n50939, n50940, n50941, n50942,
         n50943, n50944, n50945, n50946, n50947, n50948, n50949, n50950,
         n50951, n50952, n50953, n50954, n50955, n50956, n50957, n50958,
         n50959, n50960, n50961, n50962, n50963, n50964, n50965, n50966,
         n50967, n50968, n50969, n50970, n50971, n50972, n50973, n50974,
         n50975, n50976, n50977, n50978, n50979, n50980, n50981, n50982,
         n50983, n50984, n50985, n50986, n50987, n50988, n50989, n50990,
         n50991, n50992, n50993, n50994, n50995, n50996, n50997, n50998,
         n50999, n51000, n51001, n51002, n51003, n51004, n51005, n51006,
         n51007, n51008, n51009, n51010, n51011, n51012, n51013, n51014,
         n51015, n51016, n51017, n51018, n51019, n51020, n51021, n51022,
         n51023, n51024, n51025, n51026, n51027, n51028, n51029, n51030,
         n51031, n51032, n51033, n51034, n51035, n51036, n51037, n51038,
         n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046,
         n51047, n51048, n51049, n51050, n51051, n51052, n51053, n51054,
         n51055, n51056, n51057, n51058, n51059, n51060, n51061, n51062,
         n51063, n51064, n51065, n51066, n51067, n51068, n51069, n51070,
         n51071, n51072, n51073, n51074, n51075, n51076, n51077, n51078,
         n51079, n51080, n51081, n51082, n51083, n51084, n51085, n51086,
         n51087, n51088, n51089, n51090, n51091, n51092, n51093, n51094,
         n51095, n51096, n51097, n51098, n51099, n51100, n51101, n51102,
         n51103, n51104, n51105, n51106, n51107, n51108, n51109, n51110,
         n51111, n51112, n51113, n51114, n51115, n51116, n51117, n51118,
         n51119, n51120, n51121, n51122, n51123, n51124, n51125, n51126,
         n51127, n51128, n51129, n51130, n51131, n51132, n51133, n51134,
         n51135, n51136, n51137, n51138, n51139, n51140, n51141, n51142,
         n51143, n51144, n51145, n51146, n51147, n51148, n51149, n51150,
         n51151, n51152, n51153, n51154, n51155, n51156, n51157, n51158,
         n51159, n51160, n51161, n51162, n51163, n51164, n51165, n51166,
         n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174,
         n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51182,
         n51183, n51184, n51185, n51186, n51187, n51188, n51189, n51190,
         n51191, n51192, n51193, n51194, n51195, n51196, n51197, n51198,
         n51199, n51200, n51201, n51202, n51203, n51204, n51205, n51206,
         n51207, n51208, n51209, n51210, n51211, n51212, n51213, n51214,
         n51215, n51216, n51217, n51218, n51219, n51220, n51221, n51222,
         n51223, n51224, n51225, n51226, n51227, n51228, n51229, n51230,
         n51231, n51232, n51233, n51234, n51235, n51236, n51237, n51238,
         n51239, n51240, n51241, n51242, n51243, n51244, n51245, n51246,
         n51247, n51248, n51249, n51250, n51251, n51252, n51253, n51254,
         n51255, n51256, n51257, n51258, n51259, n51260, n51261, n51262,
         n51263, n51264, n51265, n51266, n51267, n51268, n51269, n51270,
         n51271, n51272, n51273, n51274, n51275, n51276, n51277, n51278,
         n51279, n51280, n51281, n51282, n51283, n51284, n51285, n51286,
         n51287, n51288, n51289, n51290, n51291, n51292, n51293, n51294,
         n51295, n51296, n51297, n51298, n51299, n51300, n51301, n51302,
         n51303, n51304, n51305, n51306, n51307, n51308, n51309, n51310,
         n51311, n51312, n51313, n51314, n51315, n51316, n51317, n51318,
         n51319, n51320, n51321, n51322, n51323, n51324, n51325, n51326,
         n51327, n51328, n51329, n51330, n51331, n51332, n51333, n51334,
         n51335, n51336, n51337, n51338, n51339, n51340, n51341, n51342,
         n51343, n51344, n51345, n51346, n51347, n51348, n51349, n51350,
         n51351, n51352, n51353, n51354, n51355, n51356, n51357, n51358,
         n51359, n51360, n51361, n51362, n51363, n51364, n51365, n51366,
         n51367, n51368, n51369, n51370, n51371, n51372, n51373, n51374,
         n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51382,
         n51383, n51384, n51385, n51386, n51387, n51388, n51389, n51390,
         n51391, n51392, n51393, n51394, n51395, n51396, n51397, n51398,
         n51399, n51400, n51401, n51402, n51403, n51404, n51405, n51406,
         n51407, n51408, n51409, n51410, n51411, n51412, n51413, n51414,
         n51415, n51416, n51417, n51418, n51419, n51420, n51421, n51422,
         n51423, n51424, n51425, n51426, n51427, n51428, n51429, n51430,
         n51431, n51432, n51433, n51434, n51435, n51436, n51437, n51438,
         n51439, n51440, n51441, n51442, n51443, n51444, n51445, n51446,
         n51447, n51448, n51449, n51450, n51451, n51452, n51453, n51454,
         n51455, n51456, n51457, n51458, n51459, n51460, n51461, n51462,
         n51463, n51464, n51465, n51466, n51467, n51468, n51469, n51470,
         n51471, n51472, n51473, n51474, n51475, n51476, n51477, n51478,
         n51479, n51480, n51481, n51482, n51483, n51484, n51485, n51486,
         n51487, n51488, n51489, n51490, n51491, n51492, n51493, n51494,
         n51495, n51496, n51497, n51498, n51499, n51500, n51501, n51502,
         n51503, n51504, n51505, n51506, n51507, n51508, n51509, n51510,
         n51511, n51512, n51513, n51514, n51515, n51516, n51517, n51518,
         n51519, n51520, n51521, n51522, n51523, n51524, n51525, n51526,
         n51527, n51528, n51529, n51530, n51531, n51532, n51533, n51534,
         n51535, n51536, n51537, n51538, n51539, n51540, n51541, n51542,
         n51543, n51544, n51545, n51546, n51547, n51548, n51549, n51550,
         n51551, n51552, n51553, n51554, n51555, n51556, n51557, n51558,
         n51559, n51560, n51561, n51562, n51563, n51564, n51565, n51566,
         n51567, n51568, n51569, n51570, n51571, n51572, n51573, n51574,
         n51575, n51576, n51577, n51578, n51579, n51580, n51581, n51582,
         n51583, n51584, n51585, n51586, n51587, n51588, n51589, n51590,
         n51591, n51592, n51593, n51594, n51595, n51596, n51597, n51598,
         n51599, n51600, n51601, n51602, n51603, n51604, n51605, n51606,
         n51607, n51608, n51609, n51610, n51611, n51612, n51613, n51614,
         n51615, n51616, n51617, n51618, n51619, n51620, n51621, n51622,
         n51623, n51624, n51625, n51626, n51627, n51628, n51629, n51630,
         n51631, n51632, n51633, n51634, n51635, n51636, n51637, n51638,
         n51639, n51640, n51641, n51642, n51643, n51644, n51645, n51646,
         n51647, n51648, n51649, n51650, n51651, n51652, n51653, n51654,
         n51655, n51656, n51657, n51658, n51659, n51660, n51661, n51662,
         n51663, n51664, n51665, n51666, n51667, n51668, n51669, n51670,
         n51671, n51672, n51673, n51674, n51675, n51676, n51677, n51678,
         n51679, n51680, n51681, n51682, n51683, n51684, n51685, n51686,
         n51687, n51688, n51689, n51690, n51691, n51692, n51693, n51694,
         n51695, n51696, n51697, n51698, n51699, n51700, n51701, n51702,
         n51703, n51704, n51705, n51706, n51707, n51708, n51709, n51710,
         n51711, n51712, n51713, n51714, n51715, n51716, n51717, n51718,
         n51719, n51720, n51721, n51722, n51723, n51724, n51725, n51726,
         n51727, n51728, n51729, n51730, n51731, n51732, n51733, n51734,
         n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742,
         n51743, n51744, n51745, n51746, n51747, n51748, n51749, n51750,
         n51751, n51752, n51753, n51754, n51755, n51756, n51757, n51758,
         n51759, n51760, n51761, n51762, n51763, n51764, n51765, n51766,
         n51767, n51768, n51769, n51770, n51771, n51772, n51773, n51774,
         n51775, n51776, n51777, n51778, n51779, n51780, n51781, n51782,
         n51783, n51784, n51785, n51786, n51787, n51788, n51789, n51790,
         n51791, n51792, n51793, n51794, n51795, n51796, n51797, n51798,
         n51799, n51800, n51801, n51802, n51803, n51804, n51805, n51806,
         n51807, n51808, n51809, n51810, n51811, n51812, n51813, n51814,
         n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51822,
         n51823, n51824, n51825, n51826, n51827, n51828, n51829, n51830,
         n51831, n51832, n51833, n51834, n51835, n51836, n51837, n51838,
         n51839, n51840, n51841, n51842, n51843, n51844, n51845, n51846,
         n51847, n51848, n51849, n51850, n51851, n51852, n51853, n51854,
         n51855, n51856, n51857, n51858, n51859, n51860, n51861, n51862,
         n51863, n51864, n51865, n51866, n51867, n51868, n51869, n51870,
         n51871, n51872, n51873, n51874, n51875, n51876, n51877, n51878,
         n51879, n51880, n51881, n51882, n51883, n51884, n51885, n51886,
         n51887, n51888, n51889, n51890, n51891, n51892, n51893, n51894,
         n51895, n51896, n51897, n51898, n51899, n51900, n51901, n51902,
         n51903, n51904, n51905, n51906, n51907, n51908, n51909, n51910,
         n51911, n51912, n51913, n51914, n51915, n51916, n51917, n51918,
         n51919, n51920, n51921, n51922, n51923, n51924, n51925, n51926,
         n51927, n51928, n51929, n51930, n51931, n51932, n51933, n51934,
         n51935, n51936, n51937, n51938, n51939, n51940, n51941, n51942,
         n51943, n51944, n51945, n51946, n51947, n51948, n51949, n51950,
         n51951, n51952, n51953, n51954, n51955, n51956, n51957, n51958,
         n51959, n51960, n51961, n51962, n51963, n51964, n51965, n51966,
         n51967, n51968, n51969, n51970, n51971, n51972, n51973, n51974,
         n51975, n51976, n51977, n51978, n51979, n51980, n51981, n51982,
         n51983, n51984, n51985, n51986, n51987, n51988, n51989, n51990,
         n51991, n51992, n51993, n51994, n51995, n51996, n51997, n51998,
         n51999, n52000, n52001, n52002, n52003, n52004, n52005, n52006,
         n52007, n52008, n52009, n52010, n52011, n52012, n52013, n52014,
         n52015, n52016, n52017, n52018, n52019, n52020, n52021, n52022,
         n52023, n52024, n52025, n52026, n52027, n52028, n52029, n52030,
         n52031, n52032, n52033, n52034, n52035, n52036, n52037, n52038,
         n52039, n52040, n52041, n52042, n52043, n52044, n52045, n52046,
         n52047, n52048, n52049, n52050, n52051, n52052, n52053, n52054,
         n52055, n52056, n52057, n52058, n52059, n52060, n52061, n52062,
         n52063, n52064, n52065, n52066, n52067, n52068, n52069, n52070,
         n52071, n52072, n52073, n52074, n52075, n52076, n52077, n52078,
         n52079, n52080, n52081, n52082, n52083, n52084, n52085, n52086,
         n52087, n52088, n52089, n52090, n52091, n52092, n52093, n52094,
         n52095, n52096, n52097, n52098, n52099, n52100, n52101, n52102,
         n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110,
         n52111, n52112, n52113, n52114, n52115, n52116, n52117, n52118,
         n52119, n52120, n52121, n52122, n52123, n52124, n52125, n52126,
         n52127, n52128, n52129, n52130, n52131, n52132, n52133, n52134,
         n52135, n52136, n52137, n52138, n52139, n52140, n52141, n52142,
         n52143, n52144, n52145, n52146, n52147, n52148, n52149, n52150,
         n52151, n52152, n52153, n52154, n52155, n52156, n52157, n52158,
         n52159, n52160, n52161, n52162, n52163, n52164, n52165, n52166,
         n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52174,
         n52175, n52176, n52177, n52178, n52179, n52180, n52181, n52182,
         n52183, n52184, n52185, n52186, n52187, n52188, n52189, n52190,
         n52191, n52192, n52193, n52194, n52195, n52196, n52197, n52198,
         n52199, n52200, n52201, n52202, n52203, n52204, n52205, n52206,
         n52207, n52208, n52209, n52210, n52211, n52212, n52213, n52214,
         n52215, n52216, n52217, n52218, n52219, n52220, n52221, n52222,
         n52223, n52224, n52225, n52226, n52227, n52228, n52229, n52230,
         n52231, n52232, n52233, n52234, n52235, n52236, n52237, n52238,
         n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246,
         n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254,
         n52255, n52256, n52257, n52258, n52259, n52260, n52261, n52262,
         n52263, n52264, n52265, n52266, n52267, n52268, n52269, n52270,
         n52271, n52272, n52273, n52274, n52275, n52276, n52277, n52278,
         n52279, n52280, n52281, n52282, n52283, n52284, n52285, n52286,
         n52287, n52288, n52289, n52290, n52291, n52292, n52293, n52294,
         n52295, n52296, n52297, n52298, n52299, n52300, n52301, n52302,
         n52303, n52304, n52305, n52306, n52307, n52308, n52309, n52310,
         n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318,
         n52319, n52320, n52321, n52322, n52323, n52324, n52325, n52326,
         n52327, n52328, n52329, n52330, n52331, n52332, n52333, n52334,
         n52335, n52336, n52337, n52338, n52339, n52340, n52341, n52342,
         n52343, n52344, n52345, n52346, n52347, n52348, n52349, n52350,
         n52351, n52352, n52353, n52354, n52355, n52356, n52357, n52358,
         n52359, n52360, n52361, n52362, n52363, n52364, n52365, n52366,
         n52367, n52368, n52369, n52370, n52371, n52372, n52373, n52374,
         n52375, n52376, n52377, n52378, n52379, n52380, n52381, n52382,
         n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390,
         n52391, n52392, n52393, n52394, n52395, n52396, n52397, n52398,
         n52399, n52400, n52401, n52402, n52403, n52404, n52405, n52406,
         n52407, n52408, n52409, n52410, n52411, n52412, n52413, n52414,
         n52415, n52416, n52417, n52418, n52419, n52420, n52421, n52422,
         n52423, n52424, n52425, n52426, n52427, n52428, n52429, n52430,
         n52431, n52432, n52433, n52434, n52435, n52436, n52437, n52438,
         n52439, n52440, n52441, n52442, n52443, n52444, n52445, n52446,
         n52447, n52448, n52449, n52450, n52451, n52452, n52453, n52454,
         n52455, n52456, n52457, n52458, n52459, n52460, n52461, n52462,
         n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470,
         n52471, n52472, n52473, n52474, n52475, n52476, n52477, n52478,
         n52479, n52480, n52481, n52482, n52483, n52484, n52485, n52486,
         n52487, n52488, n52489, n52490, n52491, n52492, n52493, n52494,
         n52495, n52496, n52497, n52498, n52499, n52500, n52501, n52502,
         n52503, n52504, n52505, n52506, n52507, n52508, n52509, n52510,
         n52511, n52512, n52513, n52514, n52515, n52516, n52517, n52518,
         n52519, n52520, n52521, n52522, n52523, n52524, n52525, n52526,
         n52527, n52528, n52529, n52530, n52531, n52532, n52533, n52534,
         n52535, n52536, n52537, n52538, n52539, n52540, n52541, n52542,
         n52543, n52544, n52545, n52546, n52547, n52548, n52549, n52550,
         n52551, n52552, n52553, n52554, n52555, n52556, n52557, n52558,
         n52559, n52560, n52561, n52562, n52563, n52564, n52565, n52566,
         n52567, n52568, n52569, n52570, n52571, n52572, n52573, n52574,
         n52575, n52576, n52577, n52578, n52579, n52580, n52581, n52582,
         n52583, n52584, n52585, n52586, n52587, n52588, n52589, n52590,
         n52591, n52592, n52593, n52594, n52595, n52596, n52597, n52598,
         n52599, n52600, n52601, n52602, n52603, n52604, n52605, n52606,
         n52607, n52608, n52609, n52610, n52611, n52612, n52613, n52614,
         n52615, n52616, n52617, n52618, n52619, n52620, n52621, n52622,
         n52623, n52624, n52625, n52626, n52627, n52628, n52629, n52630,
         n52631, n52632, n52633, n52634, n52635, n52636, n52637, n52638,
         n52639, n52640, n52641, n52642, n52643, n52644, n52645, n52646,
         n52647, n52648, n52649, n52650, n52651, n52652, n52653, n52654,
         n52655, n52656, n52657, n52658, n52659, n52660, n52661, n52662,
         n52663, n52664, n52665, n52666, n52667, n52668, n52669, n52670,
         n52671, n52672, n52673, n52674, n52675, n52676, n52677, n52678,
         n52679, n52680, n52681, n52682, n52683, n52684, n52685, n52686,
         n52687, n52688, n52689, n52690, n52691, n52692, n52693, n52694,
         n52695, n52696, n52697, n52698, n52699, n52700, n52701, n52702,
         n52703, n52704, n52705, n52706, n52707, n52708, n52709, n52710,
         n52711, n52712, n52713, n52714, n52715, n52716, n52717, n52718,
         n52719, n52720, n52721, n52722, n52723, n52724, n52725, n52726,
         n52727, n52728, n52729, n52730, n52731, n52732, n52733, n52734,
         n52735, n52736, n52737, n52738, n52739, n52740, n52741, n52742,
         n52743, n52744, n52745, n52746, n52747, n52748, n52749, n52750,
         n52751, n52752, n52753, n52754, n52755, n52756, n52757, n52758,
         n52759, n52760, n52761, n52762, n52763, n52764, n52765, n52766,
         n52767, n52768, n52769, n52770, n52771, n52772, n52773, n52774,
         n52775, n52776, n52777, n52778, n52779, n52780, n52781, n52782,
         n52783, n52784, n52785, n52786, n52787, n52788, n52789, n52790,
         n52791, n52792, n52793, n52794, n52795, n52796, n52797, n52798,
         n52799, n52800, n52801, n52802, n52803, n52804, n52805, n52806,
         n52807, n52808, n52809, n52810, n52811, n52812, n52813, n52814,
         n52815, n52816, n52817, n52818, n52819, n52820, n52821, n52822,
         n52823, n52824, n52825, n52826, n52827, n52828, n52829, n52830,
         n52831, n52832, n52833, n52834, n52835, n52836, n52837, n52838,
         n52839, n52840, n52841, n52842, n52843, n52844, n52845, n52846,
         n52847, n52848, n52849, n52850, n52851, n52852, n52853, n52854,
         n52855, n52856, n52857, n52858, n52859, n52860, n52861, n52862,
         n52863, n52864, n52865, n52866, n52867, n52868, n52869, n52870,
         n52871, n52872, n52873, n52874, n52875, n52876, n52877, n52878,
         n52879, n52880, n52881, n52882, n52883, n52884, n52885, n52886,
         n52887, n52888, n52889, n52890, n52891, n52892, n52893, n52894,
         n52895, n52896, n52897, n52898, n52899, n52900, n52901, n52902,
         n52903, n52904, n52905, n52906, n52907, n52908, n52909, n52910,
         n52911, n52912, n52913, n52914, n52915, n52916, n52917, n52918,
         n52919, n52920, n52921, n52922, n52923, n52924, n52925, n52926,
         n52927, n52928, n52929, n52930, n52931, n52932, n52933, n52934,
         n52935, n52936, n52937, n52938, n52939, n52940, n52941, n52942,
         n52943, n52944, n52945, n52946, n52947, n52948, n52949, n52950,
         n52951, n52952, n52953, n52954, n52955, n52956, n52957, n52958,
         n52959, n52960, n52961, n52962, n52963, n52964, n52965, n52966,
         n52967, n52968, n52969, n52970, n52971, n52972, n52973, n52974,
         n52975, n52976, n52977, n52978, n52979, n52980, n52981, n52982,
         n52983, n52984, n52985, n52986, n52987, n52988, n52989, n52990,
         n52991, n52992, n52993, n52994, n52995, n52996, n52997, n52998,
         n52999, n53000, n53001, n53002, n53003, n53004, n53005, n53006,
         n53007, n53008, n53009, n53010, n53011, n53012, n53013, n53014,
         n53015, n53016, n53017, n53018, n53019, n53020, n53021, n53022,
         n53023, n53024, n53025, n53026, n53027, n53028, n53029, n53030,
         n53031, n53032, n53033, n53034, n53035, n53036, n53037, n53038,
         n53039, n53040, n53041, n53042, n53043, n53044, n53045, n53046,
         n53047, n53048, n53049, n53050, n53051, n53052, n53053, n53054,
         n53055, n53056, n53057, n53058, n53059, n53060, n53061, n53062,
         n53063, n53064, n53065, n53066, n53067, n53068, n53069, n53070,
         n53071, n53072, n53073, n53074, n53075, n53076, n53077, n53078,
         n53079, n53080, n53081, n53082, n53083, n53084, n53085, n53086,
         n53087, n53088, n53089, n53090, n53091, n53092, n53093, n53094,
         n53095, n53096, n53097, n53098, n53099, n53100, n53101, n53102,
         n53103, n53104, n53105, n53106, n53107, n53108, n53109, n53110,
         n53111, n53112, n53113, n53114, n53115, n53116, n53117, n53118,
         n53119, n53120, n53121, n53122, n53123, n53124, n53125, n53126,
         n53127, n53128, n53129, n53130, n53131, n53132, n53133, n53134,
         n53135, n53136, n53137, n53138, n53139, n53140, n53141, n53142,
         n53143, n53144, n53145, n53146, n53147, n53148, n53149, n53150,
         n53151, n53152, n53153, n53154, n53155, n53156, n53157, n53158,
         n53159, n53160, n53161, n53162, n53163, n53164, n53165, n53166,
         n53167, n53168, n53169, n53170, n53171, n53172, n53173, n53174,
         n53175, n53176, n53177, n53178, n53179, n53180, n53181, n53182,
         n53183, n53184, n53185, n53186, n53187, n53188, n53189, n53190,
         n53191, n53192, n53193, n53194, n53195, n53196, n53197, n53198,
         n53199, n53200, n53201, n53202, n53203, n53204, n53205, n53206,
         n53207, n53208, n53209, n53210, n53211, n53212, n53213, n53214,
         n53215, n53216, n53217, n53218, n53219, n53220, n53221, n53222,
         n53223, n53224, n53225, n53226, n53227, n53228, n53229, n53230,
         n53231, n53232, n53233, n53234, n53235, n53236, n53237, n53238,
         n53239, n53240, n53241, n53242, n53243, n53244, n53245, n53246,
         n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254,
         n53255, n53256, n53257, n53258, n53259, n53260, n53261, n53262,
         n53263, n53264, n53265, n53266, n53267, n53268, n53269, n53270,
         n53271, n53272, n53273, n53274, n53275, n53276, n53277, n53278,
         n53279, n53280, n53281, n53282, n53283, n53284, n53285, n53286,
         n53287, n53288, n53289, n53290, n53291, n53292, n53293, n53294,
         n53295, n53296, n53297, n53298, n53299, n53300, n53301, n53302,
         n53303, n53304, n53305, n53306, n53307, n53308, n53309, n53310,
         n53311, n53312, n53313, n53314, n53315, n53316, n53317, n53318,
         n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326,
         n53327, n53328, n53329, n53330, n53331, n53332, n53333, n53334,
         n53335, n53336, n53337, n53338, n53339, n53340, n53341, n53342,
         n53343, n53344, n53345, n53346, n53347, n53348, n53349, n53350,
         n53351, n53352, n53353, n53354, n53355, n53356, n53357, n53358,
         n53359, n53360, n53361, n53362, n53363, n53364, n53365, n53366,
         n53367, n53368, n53369, n53370, n53371, n53372, n53373, n53374,
         n53375, n53376, n53377, n53378, n53379, n53380, n53381, n53382,
         n53383, n53384, n53385, n53386, n53387, n53388, n53389, n53390,
         n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398,
         n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406,
         n53407, n53408, n53409, n53410, n53411, n53412, n53413, n53414,
         n53415, n53416, n53417, n53418, n53419, n53420, n53421, n53422,
         n53423, n53424, n53425, n53426, n53427, n53428, n53429, n53430,
         n53431, n53432, n53433, n53434, n53435, n53436, n53437, n53438,
         n53439, n53440, n53441, n53442, n53443, n53444, n53445, n53446,
         n53447, n53448, n53449, n53450, n53451, n53452, n53453, n53454,
         n53455, n53456, n53457, n53458, n53459, n53460, n53461, n53462,
         n53463, n53464, n53465, n53466, n53467, n53468, n53469, n53470,
         n53471, n53472, n53473, n53474, n53475, n53476, n53477, n53478,
         n53479, n53480, n53481, n53482, n53483, n53484, n53485, n53486,
         n53487, n53488, n53489, n53490, n53491, n53492, n53493, n53494,
         n53495, n53496, n53497, n53498, n53499, n53500, n53501, n53502,
         n53503, n53504, n53505, n53506, n53507, n53508, n53509, n53510,
         n53511, n53512, n53513, n53514, n53515, n53516, n53517, n53518,
         n53519, n53520, n53521, n53522, n53523, n53524, n53525, n53526,
         n53527, n53528, n53529, n53530, n53531, n53532, n53533, n53534,
         n53535, n53536, n53537, n53538, n53539, n53540, n53541, n53542,
         n53543, n53544, n53545, n53546, n53547, n53548, n53549, n53550,
         n53551, n53552, n53553, n53554, n53555, n53556, n53557, n53558,
         n53559, n53560, n53561, n53562, n53563, n53564, n53565, n53566,
         n53567, n53568, n53569, n53570, n53571, n53572, n53573, n53574,
         n53575, n53576, n53577, n53578, n53579, n53580, n53581, n53582,
         n53583, n53584, n53585, n53586, n53587, n53588, n53589, n53590,
         n53591, n53592, n53593, n53594, n53595, n53596, n53597, n53598,
         n53599, n53600, n53601, n53602, n53603, n53604, n53605, n53606,
         n53607, n53608, n53609, n53610, n53611, n53612, n53613, n53614,
         n53615, n53616, n53617, n53618, n53619, n53620, n53621, n53622,
         n53623, n53624, n53625, n53626, n53627, n53628, n53629, n53630,
         n53631, n53632, n53633, n53634, n53635, n53636, n53637, n53638,
         n53639, n53640, n53641, n53642, n53643, n53644, n53645, n53646,
         n53647, n53648, n53649, n53650, n53651, n53652, n53653, n53654,
         n53655, n53656, n53657, n53658, n53659, n53660, n53661, n53662,
         n53663, n53664, n53665, n53666, n53667, n53668, n53669, n53670,
         n53671, n53672, n53673, n53674, n53675, n53676, n53677, n53678,
         n53679, n53680, n53681, n53682, n53683, n53684, n53685, n53686,
         n53687, n53688, n53689, n53690, n53691, n53692, n53693, n53694,
         n53695, n53696, n53697, n53698, n53699, n53700, n53701, n53702,
         n53703, n53704, n53705, n53706, n53707, n53708, n53709, n53710,
         n53711, n53712, n53713, n53714, n53715, n53716, n53717, n53718,
         n53719, n53720, n53721, n53722, n53723, n53724, n53725, n53726,
         n53727, n53728, n53729, n53730, n53731, n53732, n53733, n53734,
         n53735, n53736, n53737, n53738, n53739, n53740, n53741, n53742,
         n53743, n53744, n53745, n53746, n53747, n53748, n53749, n53750,
         n53751, n53752, n53753, n53754, n53755, n53756, n53757, n53758,
         n53759, n53760, n53761, n53762, n53763, n53764, n53765, n53766,
         n53767, n53768, n53769, n53770, n53771, n53772, n53773, n53774,
         n53775, n53776, n53777, n53778, n53779, n53780, n53781, n53782,
         n53783, n53784, n53785, n53786, n53787, n53788, n53789, n53790,
         n53791, n53792, n53793, n53794, n53795, n53796, n53797, n53798,
         n53799, n53800, n53801, n53802, n53803, n53804, n53805, n53806,
         n53807, n53808, n53809, n53810, n53811, n53812, n53813, n53814,
         n53815, n53816, n53817, n53818, n53819, n53820, n53821, n53822,
         n53823, n53824, n53825, n53826, n53827, n53828, n53829, n53830,
         n53831, n53832, n53833, n53834, n53835, n53836, n53837, n53838,
         n53839, n53840, n53841, n53842, n53843, n53844, n53845, n53846,
         n53847, n53848, n53849, n53850, n53851, n53852, n53853, n53854,
         n53855, n53856, n53857, n53858, n53859, n53860, n53861, n53862,
         n53863, n53864, n53865, n53866, n53867, n53868, n53869, n53870,
         n53871, n53872, n53873, n53874, n53875, n53876, n53877, n53878,
         n53879, n53880, n53881, n53882, n53883, n53884, n53885, n53886,
         n53887, n53888, n53889, n53890, n53891, n53892, n53893, n53894,
         n53895, n53896, n53897, n53898, n53899, n53900, n53901, n53902,
         n53903, n53904, n53905, n53906, n53907, n53908, n53909, n53910,
         n53911, n53912, n53913, n53914, n53915, n53916, n53917, n53918,
         n53919, n53920, n53921, n53922, n53923, n53924, n53925, n53926,
         n53927, n53928, n53929, n53930, n53931, n53932, n53933, n53934,
         n53935, n53936, n53937, n53938, n53939, n53940, n53941, n53942,
         n53943, n53944, n53945, n53946, n53947, n53948, n53949, n53950,
         n53951, n53952, n53953, n53954, n53955, n53956, n53957, n53958,
         n53959, n53960, n53961, n53962, n53963, n53964, n53965, n53966,
         n53967, n53968, n53969, n53970, n53971, n53972, n53973, n53974,
         n53975, n53976, n53977, n53978, n53979, n53980, n53981, n53982,
         n53983, n53984, n53985, n53986, n53987, n53988, n53989, n53990,
         n53991, n53992, n53993, n53994, n53995, n53996, n53997, n53998,
         n53999, n54000, n54001, n54002, n54003, n54004, n54005, n54006,
         n54007, n54008, n54009, n54010, n54011, n54012, n54013, n54014,
         n54015, n54016, n54017, n54018, n54019, n54020, n54021, n54022,
         n54023, n54024, n54025, n54026, n54027, n54028, n54029, n54030,
         n54031, n54032, n54033, n54034, n54035, n54036, n54037, n54038,
         n54039, n54040, n54041, n54042, n54043, n54044, n54045, n54046,
         n54047, n54048, n54049, n54050, n54051, n54052, n54053, n54054,
         n54055, n54056, n54057, n54058, n54059, n54060, n54061, n54062,
         n54063, n54064, n54065, n54066, n54067, n54068, n54069, n54070,
         n54071, n54072, n54073, n54074, n54075, n54076, n54077, n54078,
         n54079, n54080, n54081, n54082, n54083, n54084, n54085, n54086,
         n54087, n54088, n54089, n54090, n54091, n54092, n54093, n54094,
         n54095, n54096, n54097, n54098, n54099, n54100, n54101, n54102,
         n54103, n54104, n54105, n54106, n54107, n54108, n54109, n54110,
         n54111, n54112, n54113, n54114, n54115, n54116, n54117, n54118,
         n54119, n54120, n54121, n54122, n54123, n54124, n54125, n54126,
         n54127, n54128, n54129, n54130, n54131, n54132, n54133, n54134,
         n54135, n54136, n54137, n54138, n54139, n54140, n54141, n54142,
         n54143, n54144, n54145, n54146, n54147, n54148, n54149, n54150,
         n54151, n54152, n54153, n54154, n54155, n54156, n54157, n54158,
         n54159, n54160, n54161, n54162, n54163, n54164, n54165, n54166,
         n54167, n54168, n54169, n54170, n54171, n54172, n54173, n54174,
         n54175, n54176, n54177, n54178, n54179, n54180, n54181, n54182,
         n54183, n54184, n54185, n54186, n54187, n54188, n54189, n54190,
         n54191, n54192, n54193, n54194, n54195, n54196, n54197, n54198,
         n54199, n54200, n54201, n54202, n54203, n54204, n54205, n54206,
         n54207, n54208, n54209, n54210, n54211, n54212, n54213, n54214,
         n54215, n54216, n54217, n54218, n54219, n54220, n54221, n54222,
         n54223, n54224, n54225, n54226, n54227, n54228, n54229, n54230,
         n54231, n54232, n54233, n54234, n54235, n54236, n54237, n54238,
         n54239, n54240, n54241, n54242, n54243, n54244, n54245, n54246,
         n54247, n54248, n54249, n54250, n54251, n54252, n54253, n54254,
         n54255, n54256, n54257, n54258, n54259, n54260, n54261, n54262,
         n54263, n54264, n54265, n54266, n54267, n54268, n54269, n54270,
         n54271, n54272, n54273, n54274, n54275, n54276, n54277, n54278,
         n54279, n54280, n54281, n54282, n54283, n54284, n54285, n54286,
         n54287, n54288, n54289, n54290, n54291, n54292, n54293, n54294,
         n54295, n54296, n54297, n54298, n54299, n54300, n54301, n54302,
         n54303, n54304, n54305, n54306, n54307, n54308, n54309, n54310,
         n54311, n54312, n54313, n54314, n54315, n54316, n54317, n54318,
         n54319, n54320, n54321, n54322, n54323, n54324, n54325, n54326,
         n54327, n54328, n54329, n54330, n54331, n54332, n54333, n54334,
         n54335, n54336, n54337, n54338;
  wire   [12:0] olocal;
  wire   [13:0] oglobal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, 
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, 
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, 
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        SYNOPSYS_UNCONNECTED__352, SYNOPSYS_UNCONNECTED__353, 
        SYNOPSYS_UNCONNECTED__354, SYNOPSYS_UNCONNECTED__355, 
        SYNOPSYS_UNCONNECTED__356, SYNOPSYS_UNCONNECTED__357, 
        SYNOPSYS_UNCONNECTED__358, SYNOPSYS_UNCONNECTED__359, 
        SYNOPSYS_UNCONNECTED__360, SYNOPSYS_UNCONNECTED__361, 
        SYNOPSYS_UNCONNECTED__362, SYNOPSYS_UNCONNECTED__363, 
        SYNOPSYS_UNCONNECTED__364, SYNOPSYS_UNCONNECTED__365, 
        SYNOPSYS_UNCONNECTED__366, SYNOPSYS_UNCONNECTED__367, 
        SYNOPSYS_UNCONNECTED__368, SYNOPSYS_UNCONNECTED__369, 
        SYNOPSYS_UNCONNECTED__370, SYNOPSYS_UNCONNECTED__371, 
        SYNOPSYS_UNCONNECTED__372, SYNOPSYS_UNCONNECTED__373, 
        SYNOPSYS_UNCONNECTED__374, SYNOPSYS_UNCONNECTED__375, 
        SYNOPSYS_UNCONNECTED__376, SYNOPSYS_UNCONNECTED__377, 
        SYNOPSYS_UNCONNECTED__378, SYNOPSYS_UNCONNECTED__379, 
        SYNOPSYS_UNCONNECTED__380, SYNOPSYS_UNCONNECTED__381, 
        SYNOPSYS_UNCONNECTED__382, SYNOPSYS_UNCONNECTED__383, 
        SYNOPSYS_UNCONNECTED__384, SYNOPSYS_UNCONNECTED__385, 
        SYNOPSYS_UNCONNECTED__386, SYNOPSYS_UNCONNECTED__387, 
        SYNOPSYS_UNCONNECTED__388, SYNOPSYS_UNCONNECTED__389, 
        SYNOPSYS_UNCONNECTED__390, SYNOPSYS_UNCONNECTED__391, 
        SYNOPSYS_UNCONNECTED__392, SYNOPSYS_UNCONNECTED__393, 
        SYNOPSYS_UNCONNECTED__394, SYNOPSYS_UNCONNECTED__395, 
        SYNOPSYS_UNCONNECTED__396, SYNOPSYS_UNCONNECTED__397, 
        SYNOPSYS_UNCONNECTED__398, SYNOPSYS_UNCONNECTED__399, 
        SYNOPSYS_UNCONNECTED__400, SYNOPSYS_UNCONNECTED__401, 
        SYNOPSYS_UNCONNECTED__402, SYNOPSYS_UNCONNECTED__403, 
        SYNOPSYS_UNCONNECTED__404, SYNOPSYS_UNCONNECTED__405, 
        SYNOPSYS_UNCONNECTED__406, SYNOPSYS_UNCONNECTED__407, 
        SYNOPSYS_UNCONNECTED__408, SYNOPSYS_UNCONNECTED__409, 
        SYNOPSYS_UNCONNECTED__410, SYNOPSYS_UNCONNECTED__411, 
        SYNOPSYS_UNCONNECTED__412, SYNOPSYS_UNCONNECTED__413, 
        SYNOPSYS_UNCONNECTED__414, SYNOPSYS_UNCONNECTED__415, 
        SYNOPSYS_UNCONNECTED__416, SYNOPSYS_UNCONNECTED__417, 
        SYNOPSYS_UNCONNECTED__418, SYNOPSYS_UNCONNECTED__419, 
        SYNOPSYS_UNCONNECTED__420, SYNOPSYS_UNCONNECTED__421, 
        SYNOPSYS_UNCONNECTED__422, SYNOPSYS_UNCONNECTED__423, 
        SYNOPSYS_UNCONNECTED__424, SYNOPSYS_UNCONNECTED__425, 
        SYNOPSYS_UNCONNECTED__426, SYNOPSYS_UNCONNECTED__427, 
        SYNOPSYS_UNCONNECTED__428, SYNOPSYS_UNCONNECTED__429, 
        SYNOPSYS_UNCONNECTED__430, SYNOPSYS_UNCONNECTED__431, 
        SYNOPSYS_UNCONNECTED__432, SYNOPSYS_UNCONNECTED__433, 
        SYNOPSYS_UNCONNECTED__434, SYNOPSYS_UNCONNECTED__435, 
        SYNOPSYS_UNCONNECTED__436, SYNOPSYS_UNCONNECTED__437, 
        SYNOPSYS_UNCONNECTED__438, SYNOPSYS_UNCONNECTED__439, 
        SYNOPSYS_UNCONNECTED__440, SYNOPSYS_UNCONNECTED__441, 
        SYNOPSYS_UNCONNECTED__442, SYNOPSYS_UNCONNECTED__443, 
        SYNOPSYS_UNCONNECTED__444, SYNOPSYS_UNCONNECTED__445, 
        SYNOPSYS_UNCONNECTED__446, SYNOPSYS_UNCONNECTED__447, 
        SYNOPSYS_UNCONNECTED__448, SYNOPSYS_UNCONNECTED__449, 
        SYNOPSYS_UNCONNECTED__450, SYNOPSYS_UNCONNECTED__451, 
        SYNOPSYS_UNCONNECTED__452, SYNOPSYS_UNCONNECTED__453, 
        SYNOPSYS_UNCONNECTED__454, SYNOPSYS_UNCONNECTED__455, 
        SYNOPSYS_UNCONNECTED__456, SYNOPSYS_UNCONNECTED__457, 
        SYNOPSYS_UNCONNECTED__458, SYNOPSYS_UNCONNECTED__459, 
        SYNOPSYS_UNCONNECTED__460, SYNOPSYS_UNCONNECTED__461, 
        SYNOPSYS_UNCONNECTED__462, SYNOPSYS_UNCONNECTED__463, 
        SYNOPSYS_UNCONNECTED__464, SYNOPSYS_UNCONNECTED__465, 
        SYNOPSYS_UNCONNECTED__466, SYNOPSYS_UNCONNECTED__467, 
        SYNOPSYS_UNCONNECTED__468, SYNOPSYS_UNCONNECTED__469, 
        SYNOPSYS_UNCONNECTED__470, SYNOPSYS_UNCONNECTED__471, 
        SYNOPSYS_UNCONNECTED__472, SYNOPSYS_UNCONNECTED__473, 
        SYNOPSYS_UNCONNECTED__474, SYNOPSYS_UNCONNECTED__475, 
        SYNOPSYS_UNCONNECTED__476, SYNOPSYS_UNCONNECTED__477, 
        SYNOPSYS_UNCONNECTED__478, SYNOPSYS_UNCONNECTED__479, 
        SYNOPSYS_UNCONNECTED__480, SYNOPSYS_UNCONNECTED__481, 
        SYNOPSYS_UNCONNECTED__482, SYNOPSYS_UNCONNECTED__483, 
        SYNOPSYS_UNCONNECTED__484, SYNOPSYS_UNCONNECTED__485, 
        SYNOPSYS_UNCONNECTED__486, SYNOPSYS_UNCONNECTED__487, 
        SYNOPSYS_UNCONNECTED__488, SYNOPSYS_UNCONNECTED__489, 
        SYNOPSYS_UNCONNECTED__490, SYNOPSYS_UNCONNECTED__491, 
        SYNOPSYS_UNCONNECTED__492, SYNOPSYS_UNCONNECTED__493, 
        SYNOPSYS_UNCONNECTED__494, SYNOPSYS_UNCONNECTED__495, 
        SYNOPSYS_UNCONNECTED__496, SYNOPSYS_UNCONNECTED__497, 
        SYNOPSYS_UNCONNECTED__498, SYNOPSYS_UNCONNECTED__499, 
        SYNOPSYS_UNCONNECTED__500, SYNOPSYS_UNCONNECTED__501, 
        SYNOPSYS_UNCONNECTED__502, SYNOPSYS_UNCONNECTED__503, 
        SYNOPSYS_UNCONNECTED__504, SYNOPSYS_UNCONNECTED__505, 
        SYNOPSYS_UNCONNECTED__506, SYNOPSYS_UNCONNECTED__507, 
        SYNOPSYS_UNCONNECTED__508, SYNOPSYS_UNCONNECTED__509, 
        SYNOPSYS_UNCONNECTED__510, SYNOPSYS_UNCONNECTED__511, 
        SYNOPSYS_UNCONNECTED__512, SYNOPSYS_UNCONNECTED__513, 
        SYNOPSYS_UNCONNECTED__514, SYNOPSYS_UNCONNECTED__515, 
        SYNOPSYS_UNCONNECTED__516, SYNOPSYS_UNCONNECTED__517, 
        SYNOPSYS_UNCONNECTED__518, SYNOPSYS_UNCONNECTED__519, 
        SYNOPSYS_UNCONNECTED__520, SYNOPSYS_UNCONNECTED__521, 
        SYNOPSYS_UNCONNECTED__522, SYNOPSYS_UNCONNECTED__523, 
        SYNOPSYS_UNCONNECTED__524, SYNOPSYS_UNCONNECTED__525, 
        SYNOPSYS_UNCONNECTED__526, SYNOPSYS_UNCONNECTED__527, 
        SYNOPSYS_UNCONNECTED__528, SYNOPSYS_UNCONNECTED__529, 
        SYNOPSYS_UNCONNECTED__530, SYNOPSYS_UNCONNECTED__531, 
        SYNOPSYS_UNCONNECTED__532, SYNOPSYS_UNCONNECTED__533, 
        SYNOPSYS_UNCONNECTED__534, SYNOPSYS_UNCONNECTED__535, 
        SYNOPSYS_UNCONNECTED__536, SYNOPSYS_UNCONNECTED__537, 
        SYNOPSYS_UNCONNECTED__538, SYNOPSYS_UNCONNECTED__539, 
        SYNOPSYS_UNCONNECTED__540, SYNOPSYS_UNCONNECTED__541, 
        SYNOPSYS_UNCONNECTED__542, SYNOPSYS_UNCONNECTED__543, 
        SYNOPSYS_UNCONNECTED__544, SYNOPSYS_UNCONNECTED__545, 
        SYNOPSYS_UNCONNECTED__546, SYNOPSYS_UNCONNECTED__547, 
        SYNOPSYS_UNCONNECTED__548, SYNOPSYS_UNCONNECTED__549, 
        SYNOPSYS_UNCONNECTED__550, SYNOPSYS_UNCONNECTED__551, 
        SYNOPSYS_UNCONNECTED__552, SYNOPSYS_UNCONNECTED__553, 
        SYNOPSYS_UNCONNECTED__554, SYNOPSYS_UNCONNECTED__555, 
        SYNOPSYS_UNCONNECTED__556, SYNOPSYS_UNCONNECTED__557, 
        SYNOPSYS_UNCONNECTED__558, SYNOPSYS_UNCONNECTED__559, 
        SYNOPSYS_UNCONNECTED__560, SYNOPSYS_UNCONNECTED__561, 
        SYNOPSYS_UNCONNECTED__562, SYNOPSYS_UNCONNECTED__563, 
        SYNOPSYS_UNCONNECTED__564, SYNOPSYS_UNCONNECTED__565, 
        SYNOPSYS_UNCONNECTED__566, SYNOPSYS_UNCONNECTED__567, 
        SYNOPSYS_UNCONNECTED__568, SYNOPSYS_UNCONNECTED__569, 
        SYNOPSYS_UNCONNECTED__570, SYNOPSYS_UNCONNECTED__571, 
        SYNOPSYS_UNCONNECTED__572, SYNOPSYS_UNCONNECTED__573, 
        SYNOPSYS_UNCONNECTED__574, SYNOPSYS_UNCONNECTED__575, 
        SYNOPSYS_UNCONNECTED__576, SYNOPSYS_UNCONNECTED__577, 
        SYNOPSYS_UNCONNECTED__578, SYNOPSYS_UNCONNECTED__579, 
        SYNOPSYS_UNCONNECTED__580, SYNOPSYS_UNCONNECTED__581, 
        SYNOPSYS_UNCONNECTED__582, SYNOPSYS_UNCONNECTED__583, 
        SYNOPSYS_UNCONNECTED__584, SYNOPSYS_UNCONNECTED__585, 
        SYNOPSYS_UNCONNECTED__586, SYNOPSYS_UNCONNECTED__587, 
        SYNOPSYS_UNCONNECTED__588, SYNOPSYS_UNCONNECTED__589, 
        SYNOPSYS_UNCONNECTED__590, SYNOPSYS_UNCONNECTED__591, 
        SYNOPSYS_UNCONNECTED__592, SYNOPSYS_UNCONNECTED__593, 
        SYNOPSYS_UNCONNECTED__594, SYNOPSYS_UNCONNECTED__595, 
        SYNOPSYS_UNCONNECTED__596, SYNOPSYS_UNCONNECTED__597, 
        SYNOPSYS_UNCONNECTED__598, SYNOPSYS_UNCONNECTED__599, 
        SYNOPSYS_UNCONNECTED__600, SYNOPSYS_UNCONNECTED__601, 
        SYNOPSYS_UNCONNECTED__602, SYNOPSYS_UNCONNECTED__603, 
        SYNOPSYS_UNCONNECTED__604, SYNOPSYS_UNCONNECTED__605, 
        SYNOPSYS_UNCONNECTED__606, SYNOPSYS_UNCONNECTED__607, 
        SYNOPSYS_UNCONNECTED__608, SYNOPSYS_UNCONNECTED__609, 
        SYNOPSYS_UNCONNECTED__610, SYNOPSYS_UNCONNECTED__611, 
        SYNOPSYS_UNCONNECTED__612, SYNOPSYS_UNCONNECTED__613, 
        SYNOPSYS_UNCONNECTED__614, SYNOPSYS_UNCONNECTED__615, 
        SYNOPSYS_UNCONNECTED__616, SYNOPSYS_UNCONNECTED__617, 
        SYNOPSYS_UNCONNECTED__618, SYNOPSYS_UNCONNECTED__619, 
        SYNOPSYS_UNCONNECTED__620, SYNOPSYS_UNCONNECTED__621, 
        SYNOPSYS_UNCONNECTED__622, SYNOPSYS_UNCONNECTED__623, 
        SYNOPSYS_UNCONNECTED__624, SYNOPSYS_UNCONNECTED__625, 
        SYNOPSYS_UNCONNECTED__626, SYNOPSYS_UNCONNECTED__627, 
        SYNOPSYS_UNCONNECTED__628, SYNOPSYS_UNCONNECTED__629, 
        SYNOPSYS_UNCONNECTED__630, SYNOPSYS_UNCONNECTED__631, 
        SYNOPSYS_UNCONNECTED__632, SYNOPSYS_UNCONNECTED__633, 
        SYNOPSYS_UNCONNECTED__634, SYNOPSYS_UNCONNECTED__635, 
        SYNOPSYS_UNCONNECTED__636, SYNOPSYS_UNCONNECTED__637, 
        SYNOPSYS_UNCONNECTED__638, SYNOPSYS_UNCONNECTED__639, 
        SYNOPSYS_UNCONNECTED__640, SYNOPSYS_UNCONNECTED__641, 
        SYNOPSYS_UNCONNECTED__642, SYNOPSYS_UNCONNECTED__643, 
        SYNOPSYS_UNCONNECTED__644, SYNOPSYS_UNCONNECTED__645, 
        SYNOPSYS_UNCONNECTED__646, SYNOPSYS_UNCONNECTED__647, 
        SYNOPSYS_UNCONNECTED__648, SYNOPSYS_UNCONNECTED__649, 
        SYNOPSYS_UNCONNECTED__650, SYNOPSYS_UNCONNECTED__651, 
        SYNOPSYS_UNCONNECTED__652, SYNOPSYS_UNCONNECTED__653, 
        SYNOPSYS_UNCONNECTED__654, SYNOPSYS_UNCONNECTED__655, 
        SYNOPSYS_UNCONNECTED__656, SYNOPSYS_UNCONNECTED__657, 
        SYNOPSYS_UNCONNECTED__658, SYNOPSYS_UNCONNECTED__659, 
        SYNOPSYS_UNCONNECTED__660, SYNOPSYS_UNCONNECTED__661, 
        SYNOPSYS_UNCONNECTED__662, SYNOPSYS_UNCONNECTED__663, 
        SYNOPSYS_UNCONNECTED__664, SYNOPSYS_UNCONNECTED__665, 
        SYNOPSYS_UNCONNECTED__666, SYNOPSYS_UNCONNECTED__667, 
        SYNOPSYS_UNCONNECTED__668, SYNOPSYS_UNCONNECTED__669, 
        SYNOPSYS_UNCONNECTED__670, SYNOPSYS_UNCONNECTED__671, 
        SYNOPSYS_UNCONNECTED__672, SYNOPSYS_UNCONNECTED__673, 
        SYNOPSYS_UNCONNECTED__674, SYNOPSYS_UNCONNECTED__675, 
        SYNOPSYS_UNCONNECTED__676, SYNOPSYS_UNCONNECTED__677, 
        SYNOPSYS_UNCONNECTED__678, SYNOPSYS_UNCONNECTED__679, 
        SYNOPSYS_UNCONNECTED__680, SYNOPSYS_UNCONNECTED__681, 
        SYNOPSYS_UNCONNECTED__682, SYNOPSYS_UNCONNECTED__683, 
        SYNOPSYS_UNCONNECTED__684, SYNOPSYS_UNCONNECTED__685, 
        SYNOPSYS_UNCONNECTED__686, SYNOPSYS_UNCONNECTED__687, 
        SYNOPSYS_UNCONNECTED__688, SYNOPSYS_UNCONNECTED__689, 
        SYNOPSYS_UNCONNECTED__690, SYNOPSYS_UNCONNECTED__691, 
        SYNOPSYS_UNCONNECTED__692, SYNOPSYS_UNCONNECTED__693, 
        SYNOPSYS_UNCONNECTED__694, SYNOPSYS_UNCONNECTED__695, 
        SYNOPSYS_UNCONNECTED__696, SYNOPSYS_UNCONNECTED__697, 
        SYNOPSYS_UNCONNECTED__698, SYNOPSYS_UNCONNECTED__699, 
        SYNOPSYS_UNCONNECTED__700, SYNOPSYS_UNCONNECTED__701, 
        SYNOPSYS_UNCONNECTED__702, SYNOPSYS_UNCONNECTED__703, 
        SYNOPSYS_UNCONNECTED__704, SYNOPSYS_UNCONNECTED__705, 
        SYNOPSYS_UNCONNECTED__706, SYNOPSYS_UNCONNECTED__707, 
        SYNOPSYS_UNCONNECTED__708, SYNOPSYS_UNCONNECTED__709, 
        SYNOPSYS_UNCONNECTED__710, SYNOPSYS_UNCONNECTED__711, 
        SYNOPSYS_UNCONNECTED__712, SYNOPSYS_UNCONNECTED__713, 
        SYNOPSYS_UNCONNECTED__714, SYNOPSYS_UNCONNECTED__715, 
        SYNOPSYS_UNCONNECTED__716, SYNOPSYS_UNCONNECTED__717, 
        SYNOPSYS_UNCONNECTED__718, SYNOPSYS_UNCONNECTED__719, 
        SYNOPSYS_UNCONNECTED__720, SYNOPSYS_UNCONNECTED__721, 
        SYNOPSYS_UNCONNECTED__722, SYNOPSYS_UNCONNECTED__723, 
        SYNOPSYS_UNCONNECTED__724, SYNOPSYS_UNCONNECTED__725, 
        SYNOPSYS_UNCONNECTED__726, SYNOPSYS_UNCONNECTED__727, 
        SYNOPSYS_UNCONNECTED__728, SYNOPSYS_UNCONNECTED__729, 
        SYNOPSYS_UNCONNECTED__730, SYNOPSYS_UNCONNECTED__731, 
        SYNOPSYS_UNCONNECTED__732, SYNOPSYS_UNCONNECTED__733, 
        SYNOPSYS_UNCONNECTED__734, SYNOPSYS_UNCONNECTED__735, 
        SYNOPSYS_UNCONNECTED__736, SYNOPSYS_UNCONNECTED__737, 
        SYNOPSYS_UNCONNECTED__738, SYNOPSYS_UNCONNECTED__739, 
        SYNOPSYS_UNCONNECTED__740, SYNOPSYS_UNCONNECTED__741, 
        SYNOPSYS_UNCONNECTED__742, SYNOPSYS_UNCONNECTED__743, 
        SYNOPSYS_UNCONNECTED__744, SYNOPSYS_UNCONNECTED__745, 
        SYNOPSYS_UNCONNECTED__746, SYNOPSYS_UNCONNECTED__747, 
        SYNOPSYS_UNCONNECTED__748, SYNOPSYS_UNCONNECTED__749, 
        SYNOPSYS_UNCONNECTED__750, SYNOPSYS_UNCONNECTED__751, 
        SYNOPSYS_UNCONNECTED__752, SYNOPSYS_UNCONNECTED__753, 
        SYNOPSYS_UNCONNECTED__754, SYNOPSYS_UNCONNECTED__755, 
        SYNOPSYS_UNCONNECTED__756, SYNOPSYS_UNCONNECTED__757, 
        SYNOPSYS_UNCONNECTED__758, SYNOPSYS_UNCONNECTED__759, 
        SYNOPSYS_UNCONNECTED__760, SYNOPSYS_UNCONNECTED__761, 
        SYNOPSYS_UNCONNECTED__762, SYNOPSYS_UNCONNECTED__763, 
        SYNOPSYS_UNCONNECTED__764, SYNOPSYS_UNCONNECTED__765, 
        SYNOPSYS_UNCONNECTED__766, SYNOPSYS_UNCONNECTED__767, 
        SYNOPSYS_UNCONNECTED__768, SYNOPSYS_UNCONNECTED__769, 
        SYNOPSYS_UNCONNECTED__770, SYNOPSYS_UNCONNECTED__771, 
        SYNOPSYS_UNCONNECTED__772, SYNOPSYS_UNCONNECTED__773, 
        SYNOPSYS_UNCONNECTED__774, SYNOPSYS_UNCONNECTED__775, 
        SYNOPSYS_UNCONNECTED__776, SYNOPSYS_UNCONNECTED__777, 
        SYNOPSYS_UNCONNECTED__778, SYNOPSYS_UNCONNECTED__779, 
        SYNOPSYS_UNCONNECTED__780, SYNOPSYS_UNCONNECTED__781, 
        SYNOPSYS_UNCONNECTED__782, SYNOPSYS_UNCONNECTED__783, 
        SYNOPSYS_UNCONNECTED__784, SYNOPSYS_UNCONNECTED__785, 
        SYNOPSYS_UNCONNECTED__786, SYNOPSYS_UNCONNECTED__787, 
        SYNOPSYS_UNCONNECTED__788, SYNOPSYS_UNCONNECTED__789, 
        SYNOPSYS_UNCONNECTED__790, SYNOPSYS_UNCONNECTED__791, 
        SYNOPSYS_UNCONNECTED__792, SYNOPSYS_UNCONNECTED__793, 
        SYNOPSYS_UNCONNECTED__794, SYNOPSYS_UNCONNECTED__795, 
        SYNOPSYS_UNCONNECTED__796, SYNOPSYS_UNCONNECTED__797, 
        SYNOPSYS_UNCONNECTED__798, SYNOPSYS_UNCONNECTED__799, 
        SYNOPSYS_UNCONNECTED__800, SYNOPSYS_UNCONNECTED__801, 
        SYNOPSYS_UNCONNECTED__802, SYNOPSYS_UNCONNECTED__803, 
        SYNOPSYS_UNCONNECTED__804, SYNOPSYS_UNCONNECTED__805, 
        SYNOPSYS_UNCONNECTED__806, SYNOPSYS_UNCONNECTED__807, 
        SYNOPSYS_UNCONNECTED__808, SYNOPSYS_UNCONNECTED__809, 
        SYNOPSYS_UNCONNECTED__810, SYNOPSYS_UNCONNECTED__811, 
        SYNOPSYS_UNCONNECTED__812, SYNOPSYS_UNCONNECTED__813, 
        SYNOPSYS_UNCONNECTED__814, SYNOPSYS_UNCONNECTED__815, 
        SYNOPSYS_UNCONNECTED__816, SYNOPSYS_UNCONNECTED__817, 
        SYNOPSYS_UNCONNECTED__818, SYNOPSYS_UNCONNECTED__819, 
        SYNOPSYS_UNCONNECTED__820, SYNOPSYS_UNCONNECTED__821, 
        SYNOPSYS_UNCONNECTED__822, SYNOPSYS_UNCONNECTED__823, 
        SYNOPSYS_UNCONNECTED__824, SYNOPSYS_UNCONNECTED__825, 
        SYNOPSYS_UNCONNECTED__826, SYNOPSYS_UNCONNECTED__827, 
        SYNOPSYS_UNCONNECTED__828, SYNOPSYS_UNCONNECTED__829, 
        SYNOPSYS_UNCONNECTED__830, SYNOPSYS_UNCONNECTED__831, 
        SYNOPSYS_UNCONNECTED__832, SYNOPSYS_UNCONNECTED__833, 
        SYNOPSYS_UNCONNECTED__834, SYNOPSYS_UNCONNECTED__835, 
        SYNOPSYS_UNCONNECTED__836, SYNOPSYS_UNCONNECTED__837, 
        SYNOPSYS_UNCONNECTED__838, SYNOPSYS_UNCONNECTED__839, 
        SYNOPSYS_UNCONNECTED__840, SYNOPSYS_UNCONNECTED__841, 
        SYNOPSYS_UNCONNECTED__842, SYNOPSYS_UNCONNECTED__843, 
        SYNOPSYS_UNCONNECTED__844, SYNOPSYS_UNCONNECTED__845, 
        SYNOPSYS_UNCONNECTED__846, SYNOPSYS_UNCONNECTED__847, 
        SYNOPSYS_UNCONNECTED__848, SYNOPSYS_UNCONNECTED__849, 
        SYNOPSYS_UNCONNECTED__850, SYNOPSYS_UNCONNECTED__851, 
        SYNOPSYS_UNCONNECTED__852, SYNOPSYS_UNCONNECTED__853, 
        SYNOPSYS_UNCONNECTED__854, SYNOPSYS_UNCONNECTED__855, 
        SYNOPSYS_UNCONNECTED__856, SYNOPSYS_UNCONNECTED__857, 
        SYNOPSYS_UNCONNECTED__858, SYNOPSYS_UNCONNECTED__859, 
        SYNOPSYS_UNCONNECTED__860, SYNOPSYS_UNCONNECTED__861, 
        SYNOPSYS_UNCONNECTED__862, SYNOPSYS_UNCONNECTED__863, 
        SYNOPSYS_UNCONNECTED__864, SYNOPSYS_UNCONNECTED__865, 
        SYNOPSYS_UNCONNECTED__866, SYNOPSYS_UNCONNECTED__867, 
        SYNOPSYS_UNCONNECTED__868, SYNOPSYS_UNCONNECTED__869, 
        SYNOPSYS_UNCONNECTED__870, SYNOPSYS_UNCONNECTED__871, 
        SYNOPSYS_UNCONNECTED__872, SYNOPSYS_UNCONNECTED__873, 
        SYNOPSYS_UNCONNECTED__874, SYNOPSYS_UNCONNECTED__875, 
        SYNOPSYS_UNCONNECTED__876, SYNOPSYS_UNCONNECTED__877, 
        SYNOPSYS_UNCONNECTED__878, SYNOPSYS_UNCONNECTED__879, 
        SYNOPSYS_UNCONNECTED__880, SYNOPSYS_UNCONNECTED__881, 
        SYNOPSYS_UNCONNECTED__882, SYNOPSYS_UNCONNECTED__883, 
        SYNOPSYS_UNCONNECTED__884, SYNOPSYS_UNCONNECTED__885, 
        SYNOPSYS_UNCONNECTED__886, SYNOPSYS_UNCONNECTED__887, 
        SYNOPSYS_UNCONNECTED__888, SYNOPSYS_UNCONNECTED__889, 
        SYNOPSYS_UNCONNECTED__890, SYNOPSYS_UNCONNECTED__891, 
        SYNOPSYS_UNCONNECTED__892, SYNOPSYS_UNCONNECTED__893, 
        SYNOPSYS_UNCONNECTED__894, SYNOPSYS_UNCONNECTED__895, 
        SYNOPSYS_UNCONNECTED__896, SYNOPSYS_UNCONNECTED__897, 
        SYNOPSYS_UNCONNECTED__898, SYNOPSYS_UNCONNECTED__899, 
        SYNOPSYS_UNCONNECTED__900, SYNOPSYS_UNCONNECTED__901, 
        SYNOPSYS_UNCONNECTED__902, SYNOPSYS_UNCONNECTED__903, 
        SYNOPSYS_UNCONNECTED__904, SYNOPSYS_UNCONNECTED__905, 
        SYNOPSYS_UNCONNECTED__906, SYNOPSYS_UNCONNECTED__907, 
        SYNOPSYS_UNCONNECTED__908, SYNOPSYS_UNCONNECTED__909, 
        SYNOPSYS_UNCONNECTED__910, SYNOPSYS_UNCONNECTED__911, 
        SYNOPSYS_UNCONNECTED__912, SYNOPSYS_UNCONNECTED__913, 
        SYNOPSYS_UNCONNECTED__914, SYNOPSYS_UNCONNECTED__915, 
        SYNOPSYS_UNCONNECTED__916, SYNOPSYS_UNCONNECTED__917, 
        SYNOPSYS_UNCONNECTED__918, SYNOPSYS_UNCONNECTED__919, 
        SYNOPSYS_UNCONNECTED__920, SYNOPSYS_UNCONNECTED__921, 
        SYNOPSYS_UNCONNECTED__922, SYNOPSYS_UNCONNECTED__923, 
        SYNOPSYS_UNCONNECTED__924, SYNOPSYS_UNCONNECTED__925, 
        SYNOPSYS_UNCONNECTED__926, SYNOPSYS_UNCONNECTED__927, 
        SYNOPSYS_UNCONNECTED__928, SYNOPSYS_UNCONNECTED__929, 
        SYNOPSYS_UNCONNECTED__930, SYNOPSYS_UNCONNECTED__931, 
        SYNOPSYS_UNCONNECTED__932, SYNOPSYS_UNCONNECTED__933, 
        SYNOPSYS_UNCONNECTED__934, SYNOPSYS_UNCONNECTED__935, 
        SYNOPSYS_UNCONNECTED__936, SYNOPSYS_UNCONNECTED__937, 
        SYNOPSYS_UNCONNECTED__938, SYNOPSYS_UNCONNECTED__939, 
        SYNOPSYS_UNCONNECTED__940, SYNOPSYS_UNCONNECTED__941, 
        SYNOPSYS_UNCONNECTED__942, SYNOPSYS_UNCONNECTED__943, 
        SYNOPSYS_UNCONNECTED__944, SYNOPSYS_UNCONNECTED__945, 
        SYNOPSYS_UNCONNECTED__946, SYNOPSYS_UNCONNECTED__947, 
        SYNOPSYS_UNCONNECTED__948, SYNOPSYS_UNCONNECTED__949, 
        SYNOPSYS_UNCONNECTED__950, SYNOPSYS_UNCONNECTED__951, 
        SYNOPSYS_UNCONNECTED__952, SYNOPSYS_UNCONNECTED__953, 
        SYNOPSYS_UNCONNECTED__954, SYNOPSYS_UNCONNECTED__955, 
        SYNOPSYS_UNCONNECTED__956, SYNOPSYS_UNCONNECTED__957, 
        SYNOPSYS_UNCONNECTED__958, SYNOPSYS_UNCONNECTED__959, 
        SYNOPSYS_UNCONNECTED__960, SYNOPSYS_UNCONNECTED__961, 
        SYNOPSYS_UNCONNECTED__962, SYNOPSYS_UNCONNECTED__963, 
        SYNOPSYS_UNCONNECTED__964, SYNOPSYS_UNCONNECTED__965, 
        SYNOPSYS_UNCONNECTED__966, SYNOPSYS_UNCONNECTED__967, 
        SYNOPSYS_UNCONNECTED__968, SYNOPSYS_UNCONNECTED__969, 
        SYNOPSYS_UNCONNECTED__970, SYNOPSYS_UNCONNECTED__971, 
        SYNOPSYS_UNCONNECTED__972, SYNOPSYS_UNCONNECTED__973, 
        SYNOPSYS_UNCONNECTED__974, SYNOPSYS_UNCONNECTED__975, 
        SYNOPSYS_UNCONNECTED__976, SYNOPSYS_UNCONNECTED__977, 
        SYNOPSYS_UNCONNECTED__978, SYNOPSYS_UNCONNECTED__979, 
        SYNOPSYS_UNCONNECTED__980, SYNOPSYS_UNCONNECTED__981, 
        SYNOPSYS_UNCONNECTED__982, SYNOPSYS_UNCONNECTED__983, 
        SYNOPSYS_UNCONNECTED__984, SYNOPSYS_UNCONNECTED__985, 
        SYNOPSYS_UNCONNECTED__986, SYNOPSYS_UNCONNECTED__987, 
        SYNOPSYS_UNCONNECTED__988, SYNOPSYS_UNCONNECTED__989, 
        SYNOPSYS_UNCONNECTED__990, SYNOPSYS_UNCONNECTED__991, 
        SYNOPSYS_UNCONNECTED__992, SYNOPSYS_UNCONNECTED__993, 
        SYNOPSYS_UNCONNECTED__994, SYNOPSYS_UNCONNECTED__995, 
        SYNOPSYS_UNCONNECTED__996, SYNOPSYS_UNCONNECTED__997, 
        SYNOPSYS_UNCONNECTED__998, SYNOPSYS_UNCONNECTED__999, 
        SYNOPSYS_UNCONNECTED__1000, SYNOPSYS_UNCONNECTED__1001, 
        SYNOPSYS_UNCONNECTED__1002, SYNOPSYS_UNCONNECTED__1003, 
        SYNOPSYS_UNCONNECTED__1004, SYNOPSYS_UNCONNECTED__1005, 
        SYNOPSYS_UNCONNECTED__1006, SYNOPSYS_UNCONNECTED__1007, 
        SYNOPSYS_UNCONNECTED__1008, SYNOPSYS_UNCONNECTED__1009, 
        SYNOPSYS_UNCONNECTED__1010, SYNOPSYS_UNCONNECTED__1011, 
        SYNOPSYS_UNCONNECTED__1012, SYNOPSYS_UNCONNECTED__1013, 
        SYNOPSYS_UNCONNECTED__1014, SYNOPSYS_UNCONNECTED__1015, 
        SYNOPSYS_UNCONNECTED__1016, SYNOPSYS_UNCONNECTED__1017, 
        SYNOPSYS_UNCONNECTED__1018, SYNOPSYS_UNCONNECTED__1019, 
        SYNOPSYS_UNCONNECTED__1020, SYNOPSYS_UNCONNECTED__1021, 
        SYNOPSYS_UNCONNECTED__1022, SYNOPSYS_UNCONNECTED__1023, 
        SYNOPSYS_UNCONNECTED__1024, SYNOPSYS_UNCONNECTED__1025, 
        SYNOPSYS_UNCONNECTED__1026, SYNOPSYS_UNCONNECTED__1027, 
        SYNOPSYS_UNCONNECTED__1028, SYNOPSYS_UNCONNECTED__1029, 
        SYNOPSYS_UNCONNECTED__1030, SYNOPSYS_UNCONNECTED__1031, 
        SYNOPSYS_UNCONNECTED__1032, SYNOPSYS_UNCONNECTED__1033, 
        SYNOPSYS_UNCONNECTED__1034, SYNOPSYS_UNCONNECTED__1035, 
        SYNOPSYS_UNCONNECTED__1036, SYNOPSYS_UNCONNECTED__1037, 
        SYNOPSYS_UNCONNECTED__1038, SYNOPSYS_UNCONNECTED__1039, 
        SYNOPSYS_UNCONNECTED__1040, SYNOPSYS_UNCONNECTED__1041, 
        SYNOPSYS_UNCONNECTED__1042, SYNOPSYS_UNCONNECTED__1043, 
        SYNOPSYS_UNCONNECTED__1044, SYNOPSYS_UNCONNECTED__1045, 
        SYNOPSYS_UNCONNECTED__1046, SYNOPSYS_UNCONNECTED__1047, 
        SYNOPSYS_UNCONNECTED__1048, SYNOPSYS_UNCONNECTED__1049, 
        SYNOPSYS_UNCONNECTED__1050, SYNOPSYS_UNCONNECTED__1051, 
        SYNOPSYS_UNCONNECTED__1052, SYNOPSYS_UNCONNECTED__1053, 
        SYNOPSYS_UNCONNECTED__1054, SYNOPSYS_UNCONNECTED__1055, 
        SYNOPSYS_UNCONNECTED__1056, SYNOPSYS_UNCONNECTED__1057, 
        SYNOPSYS_UNCONNECTED__1058, SYNOPSYS_UNCONNECTED__1059, 
        SYNOPSYS_UNCONNECTED__1060, SYNOPSYS_UNCONNECTED__1061, 
        SYNOPSYS_UNCONNECTED__1062, SYNOPSYS_UNCONNECTED__1063, 
        SYNOPSYS_UNCONNECTED__1064, SYNOPSYS_UNCONNECTED__1065, 
        SYNOPSYS_UNCONNECTED__1066, SYNOPSYS_UNCONNECTED__1067, 
        SYNOPSYS_UNCONNECTED__1068, SYNOPSYS_UNCONNECTED__1069, 
        SYNOPSYS_UNCONNECTED__1070, SYNOPSYS_UNCONNECTED__1071, 
        SYNOPSYS_UNCONNECTED__1072, SYNOPSYS_UNCONNECTED__1073, 
        SYNOPSYS_UNCONNECTED__1074, SYNOPSYS_UNCONNECTED__1075, 
        SYNOPSYS_UNCONNECTED__1076, SYNOPSYS_UNCONNECTED__1077, 
        SYNOPSYS_UNCONNECTED__1078, SYNOPSYS_UNCONNECTED__1079, 
        SYNOPSYS_UNCONNECTED__1080, SYNOPSYS_UNCONNECTED__1081, 
        SYNOPSYS_UNCONNECTED__1082, SYNOPSYS_UNCONNECTED__1083, 
        SYNOPSYS_UNCONNECTED__1084, SYNOPSYS_UNCONNECTED__1085, 
        SYNOPSYS_UNCONNECTED__1086, SYNOPSYS_UNCONNECTED__1087, 
        SYNOPSYS_UNCONNECTED__1088, SYNOPSYS_UNCONNECTED__1089, 
        SYNOPSYS_UNCONNECTED__1090, SYNOPSYS_UNCONNECTED__1091, 
        SYNOPSYS_UNCONNECTED__1092, SYNOPSYS_UNCONNECTED__1093, 
        SYNOPSYS_UNCONNECTED__1094, SYNOPSYS_UNCONNECTED__1095, 
        SYNOPSYS_UNCONNECTED__1096, SYNOPSYS_UNCONNECTED__1097, 
        SYNOPSYS_UNCONNECTED__1098, SYNOPSYS_UNCONNECTED__1099, 
        SYNOPSYS_UNCONNECTED__1100, SYNOPSYS_UNCONNECTED__1101, 
        SYNOPSYS_UNCONNECTED__1102, SYNOPSYS_UNCONNECTED__1103, 
        SYNOPSYS_UNCONNECTED__1104, SYNOPSYS_UNCONNECTED__1105, 
        SYNOPSYS_UNCONNECTED__1106, SYNOPSYS_UNCONNECTED__1107, 
        SYNOPSYS_UNCONNECTED__1108, SYNOPSYS_UNCONNECTED__1109, 
        SYNOPSYS_UNCONNECTED__1110, SYNOPSYS_UNCONNECTED__1111, 
        SYNOPSYS_UNCONNECTED__1112, SYNOPSYS_UNCONNECTED__1113, 
        SYNOPSYS_UNCONNECTED__1114, SYNOPSYS_UNCONNECTED__1115, 
        SYNOPSYS_UNCONNECTED__1116, SYNOPSYS_UNCONNECTED__1117, 
        SYNOPSYS_UNCONNECTED__1118, SYNOPSYS_UNCONNECTED__1119, 
        SYNOPSYS_UNCONNECTED__1120, SYNOPSYS_UNCONNECTED__1121, 
        SYNOPSYS_UNCONNECTED__1122, SYNOPSYS_UNCONNECTED__1123, 
        SYNOPSYS_UNCONNECTED__1124, SYNOPSYS_UNCONNECTED__1125, 
        SYNOPSYS_UNCONNECTED__1126, SYNOPSYS_UNCONNECTED__1127, 
        SYNOPSYS_UNCONNECTED__1128, SYNOPSYS_UNCONNECTED__1129, 
        SYNOPSYS_UNCONNECTED__1130, SYNOPSYS_UNCONNECTED__1131, 
        SYNOPSYS_UNCONNECTED__1132, SYNOPSYS_UNCONNECTED__1133, 
        SYNOPSYS_UNCONNECTED__1134, SYNOPSYS_UNCONNECTED__1135, 
        SYNOPSYS_UNCONNECTED__1136, SYNOPSYS_UNCONNECTED__1137, 
        SYNOPSYS_UNCONNECTED__1138, SYNOPSYS_UNCONNECTED__1139, 
        SYNOPSYS_UNCONNECTED__1140, SYNOPSYS_UNCONNECTED__1141, 
        SYNOPSYS_UNCONNECTED__1142, SYNOPSYS_UNCONNECTED__1143, 
        SYNOPSYS_UNCONNECTED__1144, SYNOPSYS_UNCONNECTED__1145, 
        SYNOPSYS_UNCONNECTED__1146, SYNOPSYS_UNCONNECTED__1147, 
        SYNOPSYS_UNCONNECTED__1148, SYNOPSYS_UNCONNECTED__1149, 
        SYNOPSYS_UNCONNECTED__1150, SYNOPSYS_UNCONNECTED__1151, 
        SYNOPSYS_UNCONNECTED__1152, SYNOPSYS_UNCONNECTED__1153, 
        SYNOPSYS_UNCONNECTED__1154, SYNOPSYS_UNCONNECTED__1155, 
        SYNOPSYS_UNCONNECTED__1156, SYNOPSYS_UNCONNECTED__1157, 
        SYNOPSYS_UNCONNECTED__1158, SYNOPSYS_UNCONNECTED__1159, 
        SYNOPSYS_UNCONNECTED__1160, SYNOPSYS_UNCONNECTED__1161, 
        SYNOPSYS_UNCONNECTED__1162, SYNOPSYS_UNCONNECTED__1163, 
        SYNOPSYS_UNCONNECTED__1164, SYNOPSYS_UNCONNECTED__1165, 
        SYNOPSYS_UNCONNECTED__1166, SYNOPSYS_UNCONNECTED__1167, 
        SYNOPSYS_UNCONNECTED__1168, SYNOPSYS_UNCONNECTED__1169, 
        SYNOPSYS_UNCONNECTED__1170, SYNOPSYS_UNCONNECTED__1171, 
        SYNOPSYS_UNCONNECTED__1172, SYNOPSYS_UNCONNECTED__1173, 
        SYNOPSYS_UNCONNECTED__1174, SYNOPSYS_UNCONNECTED__1175, 
        SYNOPSYS_UNCONNECTED__1176, SYNOPSYS_UNCONNECTED__1177, 
        SYNOPSYS_UNCONNECTED__1178, SYNOPSYS_UNCONNECTED__1179, 
        SYNOPSYS_UNCONNECTED__1180, SYNOPSYS_UNCONNECTED__1181, 
        SYNOPSYS_UNCONNECTED__1182, SYNOPSYS_UNCONNECTED__1183, 
        SYNOPSYS_UNCONNECTED__1184, SYNOPSYS_UNCONNECTED__1185, 
        SYNOPSYS_UNCONNECTED__1186, SYNOPSYS_UNCONNECTED__1187, 
        SYNOPSYS_UNCONNECTED__1188, SYNOPSYS_UNCONNECTED__1189, 
        SYNOPSYS_UNCONNECTED__1190, SYNOPSYS_UNCONNECTED__1191, 
        SYNOPSYS_UNCONNECTED__1192, SYNOPSYS_UNCONNECTED__1193, 
        SYNOPSYS_UNCONNECTED__1194, SYNOPSYS_UNCONNECTED__1195, 
        SYNOPSYS_UNCONNECTED__1196, SYNOPSYS_UNCONNECTED__1197, 
        SYNOPSYS_UNCONNECTED__1198, SYNOPSYS_UNCONNECTED__1199, 
        SYNOPSYS_UNCONNECTED__1200, SYNOPSYS_UNCONNECTED__1201, 
        SYNOPSYS_UNCONNECTED__1202, SYNOPSYS_UNCONNECTED__1203, 
        SYNOPSYS_UNCONNECTED__1204, SYNOPSYS_UNCONNECTED__1205, 
        SYNOPSYS_UNCONNECTED__1206, SYNOPSYS_UNCONNECTED__1207, 
        SYNOPSYS_UNCONNECTED__1208, SYNOPSYS_UNCONNECTED__1209, 
        SYNOPSYS_UNCONNECTED__1210, SYNOPSYS_UNCONNECTED__1211, 
        SYNOPSYS_UNCONNECTED__1212, SYNOPSYS_UNCONNECTED__1213, 
        SYNOPSYS_UNCONNECTED__1214, SYNOPSYS_UNCONNECTED__1215, 
        SYNOPSYS_UNCONNECTED__1216, SYNOPSYS_UNCONNECTED__1217, 
        SYNOPSYS_UNCONNECTED__1218, SYNOPSYS_UNCONNECTED__1219, 
        SYNOPSYS_UNCONNECTED__1220, SYNOPSYS_UNCONNECTED__1221, 
        SYNOPSYS_UNCONNECTED__1222, SYNOPSYS_UNCONNECTED__1223, 
        SYNOPSYS_UNCONNECTED__1224, SYNOPSYS_UNCONNECTED__1225, 
        SYNOPSYS_UNCONNECTED__1226, SYNOPSYS_UNCONNECTED__1227, 
        SYNOPSYS_UNCONNECTED__1228, SYNOPSYS_UNCONNECTED__1229, 
        SYNOPSYS_UNCONNECTED__1230, SYNOPSYS_UNCONNECTED__1231, 
        SYNOPSYS_UNCONNECTED__1232, SYNOPSYS_UNCONNECTED__1233, 
        SYNOPSYS_UNCONNECTED__1234, SYNOPSYS_UNCONNECTED__1235, 
        SYNOPSYS_UNCONNECTED__1236, SYNOPSYS_UNCONNECTED__1237, 
        SYNOPSYS_UNCONNECTED__1238, SYNOPSYS_UNCONNECTED__1239, 
        SYNOPSYS_UNCONNECTED__1240, SYNOPSYS_UNCONNECTED__1241, 
        SYNOPSYS_UNCONNECTED__1242, SYNOPSYS_UNCONNECTED__1243, 
        SYNOPSYS_UNCONNECTED__1244, SYNOPSYS_UNCONNECTED__1245, 
        SYNOPSYS_UNCONNECTED__1246, SYNOPSYS_UNCONNECTED__1247, 
        SYNOPSYS_UNCONNECTED__1248, SYNOPSYS_UNCONNECTED__1249, 
        SYNOPSYS_UNCONNECTED__1250, SYNOPSYS_UNCONNECTED__1251, 
        SYNOPSYS_UNCONNECTED__1252, SYNOPSYS_UNCONNECTED__1253, 
        SYNOPSYS_UNCONNECTED__1254, SYNOPSYS_UNCONNECTED__1255, 
        SYNOPSYS_UNCONNECTED__1256, SYNOPSYS_UNCONNECTED__1257, 
        SYNOPSYS_UNCONNECTED__1258, SYNOPSYS_UNCONNECTED__1259, 
        SYNOPSYS_UNCONNECTED__1260, SYNOPSYS_UNCONNECTED__1261, 
        SYNOPSYS_UNCONNECTED__1262, SYNOPSYS_UNCONNECTED__1263, 
        SYNOPSYS_UNCONNECTED__1264, SYNOPSYS_UNCONNECTED__1265, 
        SYNOPSYS_UNCONNECTED__1266, SYNOPSYS_UNCONNECTED__1267, 
        SYNOPSYS_UNCONNECTED__1268, SYNOPSYS_UNCONNECTED__1269, 
        SYNOPSYS_UNCONNECTED__1270, SYNOPSYS_UNCONNECTED__1271, 
        SYNOPSYS_UNCONNECTED__1272, SYNOPSYS_UNCONNECTED__1273, 
        SYNOPSYS_UNCONNECTED__1274, SYNOPSYS_UNCONNECTED__1275, 
        SYNOPSYS_UNCONNECTED__1276, SYNOPSYS_UNCONNECTED__1277, 
        SYNOPSYS_UNCONNECTED__1278, SYNOPSYS_UNCONNECTED__1279, 
        SYNOPSYS_UNCONNECTED__1280, SYNOPSYS_UNCONNECTED__1281, 
        SYNOPSYS_UNCONNECTED__1282, SYNOPSYS_UNCONNECTED__1283, 
        SYNOPSYS_UNCONNECTED__1284, SYNOPSYS_UNCONNECTED__1285, 
        SYNOPSYS_UNCONNECTED__1286, SYNOPSYS_UNCONNECTED__1287, 
        SYNOPSYS_UNCONNECTED__1288, SYNOPSYS_UNCONNECTED__1289, 
        SYNOPSYS_UNCONNECTED__1290, SYNOPSYS_UNCONNECTED__1291, 
        SYNOPSYS_UNCONNECTED__1292, SYNOPSYS_UNCONNECTED__1293, 
        SYNOPSYS_UNCONNECTED__1294, SYNOPSYS_UNCONNECTED__1295, 
        SYNOPSYS_UNCONNECTED__1296, SYNOPSYS_UNCONNECTED__1297, 
        SYNOPSYS_UNCONNECTED__1298, SYNOPSYS_UNCONNECTED__1299, 
        SYNOPSYS_UNCONNECTED__1300, SYNOPSYS_UNCONNECTED__1301, 
        SYNOPSYS_UNCONNECTED__1302, SYNOPSYS_UNCONNECTED__1303, 
        SYNOPSYS_UNCONNECTED__1304, SYNOPSYS_UNCONNECTED__1305, 
        SYNOPSYS_UNCONNECTED__1306, SYNOPSYS_UNCONNECTED__1307, 
        SYNOPSYS_UNCONNECTED__1308, SYNOPSYS_UNCONNECTED__1309, 
        SYNOPSYS_UNCONNECTED__1310, SYNOPSYS_UNCONNECTED__1311, 
        SYNOPSYS_UNCONNECTED__1312, SYNOPSYS_UNCONNECTED__1313, 
        SYNOPSYS_UNCONNECTED__1314, SYNOPSYS_UNCONNECTED__1315, 
        SYNOPSYS_UNCONNECTED__1316, SYNOPSYS_UNCONNECTED__1317, 
        SYNOPSYS_UNCONNECTED__1318, SYNOPSYS_UNCONNECTED__1319, 
        SYNOPSYS_UNCONNECTED__1320, SYNOPSYS_UNCONNECTED__1321, 
        SYNOPSYS_UNCONNECTED__1322, SYNOPSYS_UNCONNECTED__1323, 
        SYNOPSYS_UNCONNECTED__1324, SYNOPSYS_UNCONNECTED__1325, 
        SYNOPSYS_UNCONNECTED__1326, SYNOPSYS_UNCONNECTED__1327, 
        SYNOPSYS_UNCONNECTED__1328, SYNOPSYS_UNCONNECTED__1329, 
        SYNOPSYS_UNCONNECTED__1330, SYNOPSYS_UNCONNECTED__1331, 
        SYNOPSYS_UNCONNECTED__1332, SYNOPSYS_UNCONNECTED__1333, 
        SYNOPSYS_UNCONNECTED__1334, SYNOPSYS_UNCONNECTED__1335, 
        SYNOPSYS_UNCONNECTED__1336, SYNOPSYS_UNCONNECTED__1337, 
        SYNOPSYS_UNCONNECTED__1338, SYNOPSYS_UNCONNECTED__1339, 
        SYNOPSYS_UNCONNECTED__1340, SYNOPSYS_UNCONNECTED__1341, 
        SYNOPSYS_UNCONNECTED__1342, SYNOPSYS_UNCONNECTED__1343, 
        SYNOPSYS_UNCONNECTED__1344, SYNOPSYS_UNCONNECTED__1345, 
        SYNOPSYS_UNCONNECTED__1346, SYNOPSYS_UNCONNECTED__1347, 
        SYNOPSYS_UNCONNECTED__1348, SYNOPSYS_UNCONNECTED__1349, 
        SYNOPSYS_UNCONNECTED__1350, SYNOPSYS_UNCONNECTED__1351, 
        SYNOPSYS_UNCONNECTED__1352, SYNOPSYS_UNCONNECTED__1353, 
        SYNOPSYS_UNCONNECTED__1354, SYNOPSYS_UNCONNECTED__1355, 
        SYNOPSYS_UNCONNECTED__1356, SYNOPSYS_UNCONNECTED__1357, 
        SYNOPSYS_UNCONNECTED__1358, SYNOPSYS_UNCONNECTED__1359, 
        SYNOPSYS_UNCONNECTED__1360, SYNOPSYS_UNCONNECTED__1361, 
        SYNOPSYS_UNCONNECTED__1362, SYNOPSYS_UNCONNECTED__1363, 
        SYNOPSYS_UNCONNECTED__1364, SYNOPSYS_UNCONNECTED__1365, 
        SYNOPSYS_UNCONNECTED__1366, SYNOPSYS_UNCONNECTED__1367, 
        SYNOPSYS_UNCONNECTED__1368, SYNOPSYS_UNCONNECTED__1369, 
        SYNOPSYS_UNCONNECTED__1370, SYNOPSYS_UNCONNECTED__1371, 
        SYNOPSYS_UNCONNECTED__1372, SYNOPSYS_UNCONNECTED__1373, 
        SYNOPSYS_UNCONNECTED__1374, SYNOPSYS_UNCONNECTED__1375, 
        SYNOPSYS_UNCONNECTED__1376, SYNOPSYS_UNCONNECTED__1377, 
        SYNOPSYS_UNCONNECTED__1378, SYNOPSYS_UNCONNECTED__1379, 
        SYNOPSYS_UNCONNECTED__1380, SYNOPSYS_UNCONNECTED__1381, 
        SYNOPSYS_UNCONNECTED__1382, SYNOPSYS_UNCONNECTED__1383, 
        SYNOPSYS_UNCONNECTED__1384, SYNOPSYS_UNCONNECTED__1385, 
        SYNOPSYS_UNCONNECTED__1386, SYNOPSYS_UNCONNECTED__1387, 
        SYNOPSYS_UNCONNECTED__1388, SYNOPSYS_UNCONNECTED__1389, 
        SYNOPSYS_UNCONNECTED__1390, SYNOPSYS_UNCONNECTED__1391, 
        SYNOPSYS_UNCONNECTED__1392, SYNOPSYS_UNCONNECTED__1393, 
        SYNOPSYS_UNCONNECTED__1394, SYNOPSYS_UNCONNECTED__1395, 
        SYNOPSYS_UNCONNECTED__1396, SYNOPSYS_UNCONNECTED__1397, 
        SYNOPSYS_UNCONNECTED__1398, SYNOPSYS_UNCONNECTED__1399, 
        SYNOPSYS_UNCONNECTED__1400, SYNOPSYS_UNCONNECTED__1401, 
        SYNOPSYS_UNCONNECTED__1402, SYNOPSYS_UNCONNECTED__1403, 
        SYNOPSYS_UNCONNECTED__1404, SYNOPSYS_UNCONNECTED__1405, 
        SYNOPSYS_UNCONNECTED__1406, SYNOPSYS_UNCONNECTED__1407, 
        SYNOPSYS_UNCONNECTED__1408, SYNOPSYS_UNCONNECTED__1409, 
        SYNOPSYS_UNCONNECTED__1410, SYNOPSYS_UNCONNECTED__1411, 
        SYNOPSYS_UNCONNECTED__1412, SYNOPSYS_UNCONNECTED__1413, 
        SYNOPSYS_UNCONNECTED__1414, SYNOPSYS_UNCONNECTED__1415, 
        SYNOPSYS_UNCONNECTED__1416, SYNOPSYS_UNCONNECTED__1417, 
        SYNOPSYS_UNCONNECTED__1418, SYNOPSYS_UNCONNECTED__1419, 
        SYNOPSYS_UNCONNECTED__1420, SYNOPSYS_UNCONNECTED__1421, 
        SYNOPSYS_UNCONNECTED__1422, SYNOPSYS_UNCONNECTED__1423, 
        SYNOPSYS_UNCONNECTED__1424, SYNOPSYS_UNCONNECTED__1425, 
        SYNOPSYS_UNCONNECTED__1426, SYNOPSYS_UNCONNECTED__1427, 
        SYNOPSYS_UNCONNECTED__1428, SYNOPSYS_UNCONNECTED__1429, 
        SYNOPSYS_UNCONNECTED__1430, SYNOPSYS_UNCONNECTED__1431, 
        SYNOPSYS_UNCONNECTED__1432, SYNOPSYS_UNCONNECTED__1433, 
        SYNOPSYS_UNCONNECTED__1434, SYNOPSYS_UNCONNECTED__1435, 
        SYNOPSYS_UNCONNECTED__1436, SYNOPSYS_UNCONNECTED__1437, 
        SYNOPSYS_UNCONNECTED__1438, SYNOPSYS_UNCONNECTED__1439, 
        SYNOPSYS_UNCONNECTED__1440, SYNOPSYS_UNCONNECTED__1441, 
        SYNOPSYS_UNCONNECTED__1442, SYNOPSYS_UNCONNECTED__1443, 
        SYNOPSYS_UNCONNECTED__1444, SYNOPSYS_UNCONNECTED__1445, 
        SYNOPSYS_UNCONNECTED__1446, SYNOPSYS_UNCONNECTED__1447, 
        SYNOPSYS_UNCONNECTED__1448, SYNOPSYS_UNCONNECTED__1449, 
        SYNOPSYS_UNCONNECTED__1450, SYNOPSYS_UNCONNECTED__1451, 
        SYNOPSYS_UNCONNECTED__1452, SYNOPSYS_UNCONNECTED__1453, 
        SYNOPSYS_UNCONNECTED__1454, SYNOPSYS_UNCONNECTED__1455, 
        SYNOPSYS_UNCONNECTED__1456, SYNOPSYS_UNCONNECTED__1457, 
        SYNOPSYS_UNCONNECTED__1458, SYNOPSYS_UNCONNECTED__1459, 
        SYNOPSYS_UNCONNECTED__1460, SYNOPSYS_UNCONNECTED__1461, 
        SYNOPSYS_UNCONNECTED__1462, SYNOPSYS_UNCONNECTED__1463, 
        SYNOPSYS_UNCONNECTED__1464, SYNOPSYS_UNCONNECTED__1465, 
        SYNOPSYS_UNCONNECTED__1466, SYNOPSYS_UNCONNECTED__1467, 
        SYNOPSYS_UNCONNECTED__1468, SYNOPSYS_UNCONNECTED__1469, 
        SYNOPSYS_UNCONNECTED__1470, SYNOPSYS_UNCONNECTED__1471, 
        SYNOPSYS_UNCONNECTED__1472, SYNOPSYS_UNCONNECTED__1473, 
        SYNOPSYS_UNCONNECTED__1474, SYNOPSYS_UNCONNECTED__1475, 
        SYNOPSYS_UNCONNECTED__1476, SYNOPSYS_UNCONNECTED__1477, 
        SYNOPSYS_UNCONNECTED__1478, SYNOPSYS_UNCONNECTED__1479, 
        SYNOPSYS_UNCONNECTED__1480, SYNOPSYS_UNCONNECTED__1481, 
        SYNOPSYS_UNCONNECTED__1482, SYNOPSYS_UNCONNECTED__1483, 
        SYNOPSYS_UNCONNECTED__1484, SYNOPSYS_UNCONNECTED__1485, 
        SYNOPSYS_UNCONNECTED__1486, SYNOPSYS_UNCONNECTED__1487, 
        SYNOPSYS_UNCONNECTED__1488, SYNOPSYS_UNCONNECTED__1489, 
        SYNOPSYS_UNCONNECTED__1490, SYNOPSYS_UNCONNECTED__1491, 
        SYNOPSYS_UNCONNECTED__1492, SYNOPSYS_UNCONNECTED__1493, 
        SYNOPSYS_UNCONNECTED__1494, SYNOPSYS_UNCONNECTED__1495, 
        SYNOPSYS_UNCONNECTED__1496, SYNOPSYS_UNCONNECTED__1497, 
        SYNOPSYS_UNCONNECTED__1498, SYNOPSYS_UNCONNECTED__1499, 
        SYNOPSYS_UNCONNECTED__1500, SYNOPSYS_UNCONNECTED__1501, 
        SYNOPSYS_UNCONNECTED__1502, SYNOPSYS_UNCONNECTED__1503, 
        SYNOPSYS_UNCONNECTED__1504, SYNOPSYS_UNCONNECTED__1505, 
        SYNOPSYS_UNCONNECTED__1506, SYNOPSYS_UNCONNECTED__1507, 
        SYNOPSYS_UNCONNECTED__1508, SYNOPSYS_UNCONNECTED__1509, 
        SYNOPSYS_UNCONNECTED__1510, SYNOPSYS_UNCONNECTED__1511, 
        SYNOPSYS_UNCONNECTED__1512, SYNOPSYS_UNCONNECTED__1513, 
        SYNOPSYS_UNCONNECTED__1514, SYNOPSYS_UNCONNECTED__1515, 
        SYNOPSYS_UNCONNECTED__1516, SYNOPSYS_UNCONNECTED__1517, 
        SYNOPSYS_UNCONNECTED__1518, SYNOPSYS_UNCONNECTED__1519, 
        SYNOPSYS_UNCONNECTED__1520, SYNOPSYS_UNCONNECTED__1521, 
        SYNOPSYS_UNCONNECTED__1522, SYNOPSYS_UNCONNECTED__1523, 
        SYNOPSYS_UNCONNECTED__1524, SYNOPSYS_UNCONNECTED__1525, 
        SYNOPSYS_UNCONNECTED__1526, SYNOPSYS_UNCONNECTED__1527, 
        SYNOPSYS_UNCONNECTED__1528, SYNOPSYS_UNCONNECTED__1529, 
        SYNOPSYS_UNCONNECTED__1530, SYNOPSYS_UNCONNECTED__1531, 
        SYNOPSYS_UNCONNECTED__1532, SYNOPSYS_UNCONNECTED__1533, 
        SYNOPSYS_UNCONNECTED__1534, SYNOPSYS_UNCONNECTED__1535, 
        SYNOPSYS_UNCONNECTED__1536, SYNOPSYS_UNCONNECTED__1537, 
        SYNOPSYS_UNCONNECTED__1538, SYNOPSYS_UNCONNECTED__1539, 
        SYNOPSYS_UNCONNECTED__1540, SYNOPSYS_UNCONNECTED__1541, 
        SYNOPSYS_UNCONNECTED__1542, SYNOPSYS_UNCONNECTED__1543, 
        SYNOPSYS_UNCONNECTED__1544, SYNOPSYS_UNCONNECTED__1545, 
        SYNOPSYS_UNCONNECTED__1546, SYNOPSYS_UNCONNECTED__1547, 
        SYNOPSYS_UNCONNECTED__1548, SYNOPSYS_UNCONNECTED__1549, 
        SYNOPSYS_UNCONNECTED__1550, SYNOPSYS_UNCONNECTED__1551, 
        SYNOPSYS_UNCONNECTED__1552, SYNOPSYS_UNCONNECTED__1553, 
        SYNOPSYS_UNCONNECTED__1554, SYNOPSYS_UNCONNECTED__1555, 
        SYNOPSYS_UNCONNECTED__1556, SYNOPSYS_UNCONNECTED__1557, 
        SYNOPSYS_UNCONNECTED__1558, SYNOPSYS_UNCONNECTED__1559, 
        SYNOPSYS_UNCONNECTED__1560, SYNOPSYS_UNCONNECTED__1561, 
        SYNOPSYS_UNCONNECTED__1562, SYNOPSYS_UNCONNECTED__1563, 
        SYNOPSYS_UNCONNECTED__1564, SYNOPSYS_UNCONNECTED__1565, 
        SYNOPSYS_UNCONNECTED__1566, SYNOPSYS_UNCONNECTED__1567, 
        SYNOPSYS_UNCONNECTED__1568, SYNOPSYS_UNCONNECTED__1569, 
        SYNOPSYS_UNCONNECTED__1570, SYNOPSYS_UNCONNECTED__1571, 
        SYNOPSYS_UNCONNECTED__1572, SYNOPSYS_UNCONNECTED__1573, 
        SYNOPSYS_UNCONNECTED__1574, SYNOPSYS_UNCONNECTED__1575, 
        SYNOPSYS_UNCONNECTED__1576, SYNOPSYS_UNCONNECTED__1577, 
        SYNOPSYS_UNCONNECTED__1578, SYNOPSYS_UNCONNECTED__1579, 
        SYNOPSYS_UNCONNECTED__1580, SYNOPSYS_UNCONNECTED__1581, 
        SYNOPSYS_UNCONNECTED__1582, SYNOPSYS_UNCONNECTED__1583, 
        SYNOPSYS_UNCONNECTED__1584, SYNOPSYS_UNCONNECTED__1585, 
        SYNOPSYS_UNCONNECTED__1586, SYNOPSYS_UNCONNECTED__1587, 
        SYNOPSYS_UNCONNECTED__1588, SYNOPSYS_UNCONNECTED__1589, 
        SYNOPSYS_UNCONNECTED__1590, SYNOPSYS_UNCONNECTED__1591, 
        SYNOPSYS_UNCONNECTED__1592, SYNOPSYS_UNCONNECTED__1593, 
        SYNOPSYS_UNCONNECTED__1594, SYNOPSYS_UNCONNECTED__1595, 
        SYNOPSYS_UNCONNECTED__1596, SYNOPSYS_UNCONNECTED__1597, 
        SYNOPSYS_UNCONNECTED__1598, SYNOPSYS_UNCONNECTED__1599, 
        SYNOPSYS_UNCONNECTED__1600, SYNOPSYS_UNCONNECTED__1601, 
        SYNOPSYS_UNCONNECTED__1602, SYNOPSYS_UNCONNECTED__1603, 
        SYNOPSYS_UNCONNECTED__1604, SYNOPSYS_UNCONNECTED__1605, 
        SYNOPSYS_UNCONNECTED__1606, SYNOPSYS_UNCONNECTED__1607, 
        SYNOPSYS_UNCONNECTED__1608, SYNOPSYS_UNCONNECTED__1609, 
        SYNOPSYS_UNCONNECTED__1610, SYNOPSYS_UNCONNECTED__1611, 
        SYNOPSYS_UNCONNECTED__1612, SYNOPSYS_UNCONNECTED__1613, 
        SYNOPSYS_UNCONNECTED__1614, SYNOPSYS_UNCONNECTED__1615, 
        SYNOPSYS_UNCONNECTED__1616, SYNOPSYS_UNCONNECTED__1617, 
        SYNOPSYS_UNCONNECTED__1618, SYNOPSYS_UNCONNECTED__1619, 
        SYNOPSYS_UNCONNECTED__1620, SYNOPSYS_UNCONNECTED__1621, 
        SYNOPSYS_UNCONNECTED__1622, SYNOPSYS_UNCONNECTED__1623, 
        SYNOPSYS_UNCONNECTED__1624, SYNOPSYS_UNCONNECTED__1625, 
        SYNOPSYS_UNCONNECTED__1626, SYNOPSYS_UNCONNECTED__1627, 
        SYNOPSYS_UNCONNECTED__1628, SYNOPSYS_UNCONNECTED__1629, 
        SYNOPSYS_UNCONNECTED__1630, SYNOPSYS_UNCONNECTED__1631, 
        SYNOPSYS_UNCONNECTED__1632, SYNOPSYS_UNCONNECTED__1633, 
        SYNOPSYS_UNCONNECTED__1634, SYNOPSYS_UNCONNECTED__1635, 
        SYNOPSYS_UNCONNECTED__1636, SYNOPSYS_UNCONNECTED__1637, 
        SYNOPSYS_UNCONNECTED__1638, SYNOPSYS_UNCONNECTED__1639, 
        SYNOPSYS_UNCONNECTED__1640, SYNOPSYS_UNCONNECTED__1641, 
        SYNOPSYS_UNCONNECTED__1642, SYNOPSYS_UNCONNECTED__1643, 
        SYNOPSYS_UNCONNECTED__1644, SYNOPSYS_UNCONNECTED__1645, 
        SYNOPSYS_UNCONNECTED__1646, SYNOPSYS_UNCONNECTED__1647, 
        SYNOPSYS_UNCONNECTED__1648, SYNOPSYS_UNCONNECTED__1649, 
        SYNOPSYS_UNCONNECTED__1650, SYNOPSYS_UNCONNECTED__1651, 
        SYNOPSYS_UNCONNECTED__1652, SYNOPSYS_UNCONNECTED__1653, 
        SYNOPSYS_UNCONNECTED__1654, SYNOPSYS_UNCONNECTED__1655, 
        SYNOPSYS_UNCONNECTED__1656, SYNOPSYS_UNCONNECTED__1657, 
        SYNOPSYS_UNCONNECTED__1658, SYNOPSYS_UNCONNECTED__1659, 
        SYNOPSYS_UNCONNECTED__1660, SYNOPSYS_UNCONNECTED__1661, 
        SYNOPSYS_UNCONNECTED__1662, SYNOPSYS_UNCONNECTED__1663, 
        SYNOPSYS_UNCONNECTED__1664, SYNOPSYS_UNCONNECTED__1665, 
        SYNOPSYS_UNCONNECTED__1666, SYNOPSYS_UNCONNECTED__1667, 
        SYNOPSYS_UNCONNECTED__1668, SYNOPSYS_UNCONNECTED__1669, 
        SYNOPSYS_UNCONNECTED__1670, SYNOPSYS_UNCONNECTED__1671, 
        SYNOPSYS_UNCONNECTED__1672, SYNOPSYS_UNCONNECTED__1673, 
        SYNOPSYS_UNCONNECTED__1674, SYNOPSYS_UNCONNECTED__1675, 
        SYNOPSYS_UNCONNECTED__1676, SYNOPSYS_UNCONNECTED__1677, 
        SYNOPSYS_UNCONNECTED__1678, SYNOPSYS_UNCONNECTED__1679, 
        SYNOPSYS_UNCONNECTED__1680, SYNOPSYS_UNCONNECTED__1681, 
        SYNOPSYS_UNCONNECTED__1682, SYNOPSYS_UNCONNECTED__1683, 
        SYNOPSYS_UNCONNECTED__1684, SYNOPSYS_UNCONNECTED__1685, 
        SYNOPSYS_UNCONNECTED__1686, SYNOPSYS_UNCONNECTED__1687, 
        SYNOPSYS_UNCONNECTED__1688, SYNOPSYS_UNCONNECTED__1689, 
        SYNOPSYS_UNCONNECTED__1690, SYNOPSYS_UNCONNECTED__1691, 
        SYNOPSYS_UNCONNECTED__1692, SYNOPSYS_UNCONNECTED__1693, 
        SYNOPSYS_UNCONNECTED__1694, SYNOPSYS_UNCONNECTED__1695, 
        SYNOPSYS_UNCONNECTED__1696, SYNOPSYS_UNCONNECTED__1697, 
        SYNOPSYS_UNCONNECTED__1698, SYNOPSYS_UNCONNECTED__1699, 
        SYNOPSYS_UNCONNECTED__1700, SYNOPSYS_UNCONNECTED__1701, 
        SYNOPSYS_UNCONNECTED__1702, SYNOPSYS_UNCONNECTED__1703, 
        SYNOPSYS_UNCONNECTED__1704, SYNOPSYS_UNCONNECTED__1705, 
        SYNOPSYS_UNCONNECTED__1706, SYNOPSYS_UNCONNECTED__1707, 
        SYNOPSYS_UNCONNECTED__1708, SYNOPSYS_UNCONNECTED__1709, 
        SYNOPSYS_UNCONNECTED__1710, SYNOPSYS_UNCONNECTED__1711, 
        SYNOPSYS_UNCONNECTED__1712, SYNOPSYS_UNCONNECTED__1713, 
        SYNOPSYS_UNCONNECTED__1714, SYNOPSYS_UNCONNECTED__1715, 
        SYNOPSYS_UNCONNECTED__1716, SYNOPSYS_UNCONNECTED__1717, 
        SYNOPSYS_UNCONNECTED__1718, SYNOPSYS_UNCONNECTED__1719, 
        SYNOPSYS_UNCONNECTED__1720, SYNOPSYS_UNCONNECTED__1721, 
        SYNOPSYS_UNCONNECTED__1722, SYNOPSYS_UNCONNECTED__1723, 
        SYNOPSYS_UNCONNECTED__1724, SYNOPSYS_UNCONNECTED__1725, 
        SYNOPSYS_UNCONNECTED__1726, SYNOPSYS_UNCONNECTED__1727, 
        SYNOPSYS_UNCONNECTED__1728, SYNOPSYS_UNCONNECTED__1729, 
        SYNOPSYS_UNCONNECTED__1730, SYNOPSYS_UNCONNECTED__1731, 
        SYNOPSYS_UNCONNECTED__1732, SYNOPSYS_UNCONNECTED__1733, 
        SYNOPSYS_UNCONNECTED__1734, SYNOPSYS_UNCONNECTED__1735, 
        SYNOPSYS_UNCONNECTED__1736, SYNOPSYS_UNCONNECTED__1737, 
        SYNOPSYS_UNCONNECTED__1738, SYNOPSYS_UNCONNECTED__1739, 
        SYNOPSYS_UNCONNECTED__1740, SYNOPSYS_UNCONNECTED__1741, 
        SYNOPSYS_UNCONNECTED__1742, SYNOPSYS_UNCONNECTED__1743, 
        SYNOPSYS_UNCONNECTED__1744, SYNOPSYS_UNCONNECTED__1745, 
        SYNOPSYS_UNCONNECTED__1746, SYNOPSYS_UNCONNECTED__1747, 
        SYNOPSYS_UNCONNECTED__1748, SYNOPSYS_UNCONNECTED__1749, 
        SYNOPSYS_UNCONNECTED__1750, SYNOPSYS_UNCONNECTED__1751, 
        SYNOPSYS_UNCONNECTED__1752, SYNOPSYS_UNCONNECTED__1753, 
        SYNOPSYS_UNCONNECTED__1754, SYNOPSYS_UNCONNECTED__1755, 
        SYNOPSYS_UNCONNECTED__1756, SYNOPSYS_UNCONNECTED__1757, 
        SYNOPSYS_UNCONNECTED__1758, SYNOPSYS_UNCONNECTED__1759, 
        SYNOPSYS_UNCONNECTED__1760, SYNOPSYS_UNCONNECTED__1761, 
        SYNOPSYS_UNCONNECTED__1762, SYNOPSYS_UNCONNECTED__1763, 
        SYNOPSYS_UNCONNECTED__1764, SYNOPSYS_UNCONNECTED__1765, 
        SYNOPSYS_UNCONNECTED__1766, SYNOPSYS_UNCONNECTED__1767, 
        SYNOPSYS_UNCONNECTED__1768, SYNOPSYS_UNCONNECTED__1769, 
        SYNOPSYS_UNCONNECTED__1770, SYNOPSYS_UNCONNECTED__1771, 
        SYNOPSYS_UNCONNECTED__1772, SYNOPSYS_UNCONNECTED__1773, 
        SYNOPSYS_UNCONNECTED__1774, SYNOPSYS_UNCONNECTED__1775, 
        SYNOPSYS_UNCONNECTED__1776, SYNOPSYS_UNCONNECTED__1777, 
        SYNOPSYS_UNCONNECTED__1778, SYNOPSYS_UNCONNECTED__1779, 
        SYNOPSYS_UNCONNECTED__1780, SYNOPSYS_UNCONNECTED__1781, 
        SYNOPSYS_UNCONNECTED__1782, SYNOPSYS_UNCONNECTED__1783, 
        SYNOPSYS_UNCONNECTED__1784, SYNOPSYS_UNCONNECTED__1785, 
        SYNOPSYS_UNCONNECTED__1786, SYNOPSYS_UNCONNECTED__1787, 
        SYNOPSYS_UNCONNECTED__1788, SYNOPSYS_UNCONNECTED__1789, 
        SYNOPSYS_UNCONNECTED__1790, SYNOPSYS_UNCONNECTED__1791, 
        SYNOPSYS_UNCONNECTED__1792, SYNOPSYS_UNCONNECTED__1793, 
        SYNOPSYS_UNCONNECTED__1794, SYNOPSYS_UNCONNECTED__1795, 
        SYNOPSYS_UNCONNECTED__1796, SYNOPSYS_UNCONNECTED__1797, 
        SYNOPSYS_UNCONNECTED__1798, SYNOPSYS_UNCONNECTED__1799, 
        SYNOPSYS_UNCONNECTED__1800, SYNOPSYS_UNCONNECTED__1801, 
        SYNOPSYS_UNCONNECTED__1802, SYNOPSYS_UNCONNECTED__1803, 
        SYNOPSYS_UNCONNECTED__1804, SYNOPSYS_UNCONNECTED__1805, 
        SYNOPSYS_UNCONNECTED__1806, SYNOPSYS_UNCONNECTED__1807, 
        SYNOPSYS_UNCONNECTED__1808, SYNOPSYS_UNCONNECTED__1809, 
        SYNOPSYS_UNCONNECTED__1810, SYNOPSYS_UNCONNECTED__1811, 
        SYNOPSYS_UNCONNECTED__1812, SYNOPSYS_UNCONNECTED__1813, 
        SYNOPSYS_UNCONNECTED__1814, SYNOPSYS_UNCONNECTED__1815, 
        SYNOPSYS_UNCONNECTED__1816, SYNOPSYS_UNCONNECTED__1817, 
        SYNOPSYS_UNCONNECTED__1818, SYNOPSYS_UNCONNECTED__1819, 
        SYNOPSYS_UNCONNECTED__1820, SYNOPSYS_UNCONNECTED__1821, 
        SYNOPSYS_UNCONNECTED__1822, SYNOPSYS_UNCONNECTED__1823, 
        SYNOPSYS_UNCONNECTED__1824, SYNOPSYS_UNCONNECTED__1825, 
        SYNOPSYS_UNCONNECTED__1826, SYNOPSYS_UNCONNECTED__1827, 
        SYNOPSYS_UNCONNECTED__1828, SYNOPSYS_UNCONNECTED__1829, 
        SYNOPSYS_UNCONNECTED__1830, SYNOPSYS_UNCONNECTED__1831, 
        SYNOPSYS_UNCONNECTED__1832, SYNOPSYS_UNCONNECTED__1833, 
        SYNOPSYS_UNCONNECTED__1834, SYNOPSYS_UNCONNECTED__1835, 
        SYNOPSYS_UNCONNECTED__1836, SYNOPSYS_UNCONNECTED__1837, 
        SYNOPSYS_UNCONNECTED__1838, SYNOPSYS_UNCONNECTED__1839, 
        SYNOPSYS_UNCONNECTED__1840, SYNOPSYS_UNCONNECTED__1841, 
        SYNOPSYS_UNCONNECTED__1842, SYNOPSYS_UNCONNECTED__1843, 
        SYNOPSYS_UNCONNECTED__1844, SYNOPSYS_UNCONNECTED__1845, 
        SYNOPSYS_UNCONNECTED__1846, SYNOPSYS_UNCONNECTED__1847, 
        SYNOPSYS_UNCONNECTED__1848, SYNOPSYS_UNCONNECTED__1849, 
        SYNOPSYS_UNCONNECTED__1850, SYNOPSYS_UNCONNECTED__1851, 
        SYNOPSYS_UNCONNECTED__1852, SYNOPSYS_UNCONNECTED__1853, 
        SYNOPSYS_UNCONNECTED__1854, SYNOPSYS_UNCONNECTED__1855, 
        SYNOPSYS_UNCONNECTED__1856, SYNOPSYS_UNCONNECTED__1857, 
        SYNOPSYS_UNCONNECTED__1858, SYNOPSYS_UNCONNECTED__1859, 
        SYNOPSYS_UNCONNECTED__1860, SYNOPSYS_UNCONNECTED__1861, 
        SYNOPSYS_UNCONNECTED__1862, SYNOPSYS_UNCONNECTED__1863, 
        SYNOPSYS_UNCONNECTED__1864, SYNOPSYS_UNCONNECTED__1865, 
        SYNOPSYS_UNCONNECTED__1866, SYNOPSYS_UNCONNECTED__1867, 
        SYNOPSYS_UNCONNECTED__1868, SYNOPSYS_UNCONNECTED__1869, 
        SYNOPSYS_UNCONNECTED__1870, SYNOPSYS_UNCONNECTED__1871, 
        SYNOPSYS_UNCONNECTED__1872, SYNOPSYS_UNCONNECTED__1873, 
        SYNOPSYS_UNCONNECTED__1874, SYNOPSYS_UNCONNECTED__1875, 
        SYNOPSYS_UNCONNECTED__1876, SYNOPSYS_UNCONNECTED__1877, 
        SYNOPSYS_UNCONNECTED__1878, SYNOPSYS_UNCONNECTED__1879, 
        SYNOPSYS_UNCONNECTED__1880, SYNOPSYS_UNCONNECTED__1881, 
        SYNOPSYS_UNCONNECTED__1882, SYNOPSYS_UNCONNECTED__1883, 
        SYNOPSYS_UNCONNECTED__1884, SYNOPSYS_UNCONNECTED__1885, 
        SYNOPSYS_UNCONNECTED__1886, SYNOPSYS_UNCONNECTED__1887, 
        SYNOPSYS_UNCONNECTED__1888, SYNOPSYS_UNCONNECTED__1889, 
        SYNOPSYS_UNCONNECTED__1890, SYNOPSYS_UNCONNECTED__1891, 
        SYNOPSYS_UNCONNECTED__1892, SYNOPSYS_UNCONNECTED__1893, 
        SYNOPSYS_UNCONNECTED__1894, SYNOPSYS_UNCONNECTED__1895, 
        SYNOPSYS_UNCONNECTED__1896, SYNOPSYS_UNCONNECTED__1897, 
        SYNOPSYS_UNCONNECTED__1898, SYNOPSYS_UNCONNECTED__1899, 
        SYNOPSYS_UNCONNECTED__1900, SYNOPSYS_UNCONNECTED__1901, 
        SYNOPSYS_UNCONNECTED__1902, SYNOPSYS_UNCONNECTED__1903, 
        SYNOPSYS_UNCONNECTED__1904, SYNOPSYS_UNCONNECTED__1905, 
        SYNOPSYS_UNCONNECTED__1906, SYNOPSYS_UNCONNECTED__1907, 
        SYNOPSYS_UNCONNECTED__1908, SYNOPSYS_UNCONNECTED__1909, 
        SYNOPSYS_UNCONNECTED__1910, SYNOPSYS_UNCONNECTED__1911, 
        SYNOPSYS_UNCONNECTED__1912, SYNOPSYS_UNCONNECTED__1913, 
        SYNOPSYS_UNCONNECTED__1914, SYNOPSYS_UNCONNECTED__1915, 
        SYNOPSYS_UNCONNECTED__1916, SYNOPSYS_UNCONNECTED__1917, 
        SYNOPSYS_UNCONNECTED__1918, SYNOPSYS_UNCONNECTED__1919, 
        SYNOPSYS_UNCONNECTED__1920, SYNOPSYS_UNCONNECTED__1921, 
        SYNOPSYS_UNCONNECTED__1922, SYNOPSYS_UNCONNECTED__1923, 
        SYNOPSYS_UNCONNECTED__1924, SYNOPSYS_UNCONNECTED__1925, 
        SYNOPSYS_UNCONNECTED__1926, SYNOPSYS_UNCONNECTED__1927, 
        SYNOPSYS_UNCONNECTED__1928, SYNOPSYS_UNCONNECTED__1929, 
        SYNOPSYS_UNCONNECTED__1930, SYNOPSYS_UNCONNECTED__1931, 
        SYNOPSYS_UNCONNECTED__1932, SYNOPSYS_UNCONNECTED__1933, 
        SYNOPSYS_UNCONNECTED__1934, SYNOPSYS_UNCONNECTED__1935, 
        SYNOPSYS_UNCONNECTED__1936, SYNOPSYS_UNCONNECTED__1937, 
        SYNOPSYS_UNCONNECTED__1938, SYNOPSYS_UNCONNECTED__1939, 
        SYNOPSYS_UNCONNECTED__1940, SYNOPSYS_UNCONNECTED__1941, 
        SYNOPSYS_UNCONNECTED__1942, SYNOPSYS_UNCONNECTED__1943, 
        SYNOPSYS_UNCONNECTED__1944, SYNOPSYS_UNCONNECTED__1945, 
        SYNOPSYS_UNCONNECTED__1946, SYNOPSYS_UNCONNECTED__1947, 
        SYNOPSYS_UNCONNECTED__1948, SYNOPSYS_UNCONNECTED__1949, 
        SYNOPSYS_UNCONNECTED__1950, SYNOPSYS_UNCONNECTED__1951, 
        SYNOPSYS_UNCONNECTED__1952, SYNOPSYS_UNCONNECTED__1953, 
        SYNOPSYS_UNCONNECTED__1954, SYNOPSYS_UNCONNECTED__1955, 
        SYNOPSYS_UNCONNECTED__1956, SYNOPSYS_UNCONNECTED__1957, 
        SYNOPSYS_UNCONNECTED__1958, SYNOPSYS_UNCONNECTED__1959, 
        SYNOPSYS_UNCONNECTED__1960, SYNOPSYS_UNCONNECTED__1961, 
        SYNOPSYS_UNCONNECTED__1962, SYNOPSYS_UNCONNECTED__1963, 
        SYNOPSYS_UNCONNECTED__1964, SYNOPSYS_UNCONNECTED__1965, 
        SYNOPSYS_UNCONNECTED__1966, SYNOPSYS_UNCONNECTED__1967, 
        SYNOPSYS_UNCONNECTED__1968, SYNOPSYS_UNCONNECTED__1969, 
        SYNOPSYS_UNCONNECTED__1970, SYNOPSYS_UNCONNECTED__1971, 
        SYNOPSYS_UNCONNECTED__1972, SYNOPSYS_UNCONNECTED__1973, 
        SYNOPSYS_UNCONNECTED__1974, SYNOPSYS_UNCONNECTED__1975, 
        SYNOPSYS_UNCONNECTED__1976, SYNOPSYS_UNCONNECTED__1977, 
        SYNOPSYS_UNCONNECTED__1978, SYNOPSYS_UNCONNECTED__1979, 
        SYNOPSYS_UNCONNECTED__1980, SYNOPSYS_UNCONNECTED__1981, 
        SYNOPSYS_UNCONNECTED__1982, SYNOPSYS_UNCONNECTED__1983, 
        SYNOPSYS_UNCONNECTED__1984, SYNOPSYS_UNCONNECTED__1985, 
        SYNOPSYS_UNCONNECTED__1986, SYNOPSYS_UNCONNECTED__1987, 
        SYNOPSYS_UNCONNECTED__1988, SYNOPSYS_UNCONNECTED__1989, 
        SYNOPSYS_UNCONNECTED__1990, SYNOPSYS_UNCONNECTED__1991, 
        SYNOPSYS_UNCONNECTED__1992, SYNOPSYS_UNCONNECTED__1993, 
        SYNOPSYS_UNCONNECTED__1994, SYNOPSYS_UNCONNECTED__1995, 
        SYNOPSYS_UNCONNECTED__1996, SYNOPSYS_UNCONNECTED__1997, 
        SYNOPSYS_UNCONNECTED__1998, SYNOPSYS_UNCONNECTED__1999, 
        SYNOPSYS_UNCONNECTED__2000, SYNOPSYS_UNCONNECTED__2001, 
        SYNOPSYS_UNCONNECTED__2002, SYNOPSYS_UNCONNECTED__2003;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  hamming_N16000_CC2_DW01_add_0 add_97 ( .A(oglobal), .B({1'b0, olocal}), .CI(
        1'b0), .SUM(o) );
  hamming_N16000_CC2_DW01_add_1 add_2667_root_add_71_I832 ( .A({1'b0, N69222, 
        N69221, N69220, N69219, N69218, N69217, N69216, N69215, N69214, N69213, 
        N69212, N69211}), .B({N69236, N69235, N69234, N69233, N69232, N69231, 
        N69230, N69229, N69228, N69227, N69226, N69225, N69224}), .CI(1'b0), 
        .SUM(olocal) );
  hamming_N16000_CC2_DW01_add_2 add_2668_root_add_71_I832 ( .A({1'b0, N69196, 
        N69195, N69194, N69193, N69192, N69191, N69190, N69189, N69188, N69187, 
        N69186, N69185}), .B({1'b0, N69209, N69208, N69207, N69206, N69205, 
        N69204, N69203, N69202, N69201, N69200, N69199, N69198}), .CI(1'b0), 
        .SUM({N69236, N69235, N69234, N69233, N69232, N69231, N69230, N69229, 
        N69228, N69227, N69226, N69225, N69224}) );
  hamming_N16000_CC2_DW01_add_3 add_2669_root_add_71_I832 ( .A({1'b0, 1'b0, 
        N69169, N69168, N69167, N69166, N69165, N69164, N69163, N69162, N69161, 
        N69160, N69159}), .B({1'b0, 1'b0, N69182, N69181, N69180, N69179, 
        N69178, N69177, N69176, N69175, N69174, N69173, N69172}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N69222, N69221, N69220, N69219, N69218, 
        N69217, N69216, N69215, N69214, N69213, N69212, N69211}) );
  hamming_N16000_CC2_DW01_add_4 add_2670_root_add_71_I832 ( .A({1'b0, 1'b0, 
        N69143, N69142, N69141, N69140, N69139, N69138, N69137, N69136, N69135, 
        N69134, N69133}), .B({1'b0, 1'b0, N69156, N69155, N69154, N69153, 
        N69152, N69151, N69150, N69149, N69148, N69147, N69146}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__1, N69209, N69208, N69207, N69206, N69205, 
        N69204, N69203, N69202, N69201, N69200, N69199, N69198}) );
  hamming_N16000_CC2_DW01_add_5 add_2671_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, N69116, N69115, N69114, N69113, N69112, N69111, N69110, N69109, 
        N69108, N69107}), .B({1'b0, 1'b0, N69130, N69129, N69128, N69127, 
        N69126, N69125, N69124, N69123, N69122, N69121, N69120}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__2, N69196, N69195, N69194, N69193, N69192, 
        N69191, N69190, N69189, N69188, N69187, N69186, N69185}) );
  hamming_N16000_CC2_DW01_add_6 add_2672_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, N69090, N69089, N69088, N69087, N69086, N69085, N69084, N69083, 
        N69082, N69081}), .B({1'b0, 1'b0, 1'b0, N69103, N69102, N69101, N69100, 
        N69099, N69098, N69097, N69096, N69095, N69094}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, N69182, N69181, 
        N69180, N69179, N69178, N69177, N69176, N69175, N69174, N69173, N69172}) );
  hamming_N16000_CC2_DW01_add_7 add_2673_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, N69064, N69063, N69062, N69061, N69060, N69059, N69058, N69057, 
        N69056, N69055}), .B({1'b0, 1'b0, 1'b0, N69077, N69076, N69075, N69074, 
        N69073, N69072, N69071, N69070, N69069, N69068}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, N69169, N69168, 
        N69167, N69166, N69165, N69164, N69163, N69162, N69161, N69160, N69159}) );
  hamming_N16000_CC2_DW01_add_8 add_2674_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, N69038, N69037, N69036, N69035, N69034, N69033, N69032, N69031, 
        N69030, N69029}), .B({1'b0, 1'b0, 1'b0, N69051, N69050, N69049, N69048, 
        N69047, N69046, N69045, N69044, N69043, N69042}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, N69156, N69155, 
        N69154, N69153, N69152, N69151, N69150, N69149, N69148, N69147, N69146}) );
  hamming_N16000_CC2_DW01_add_9 add_2675_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, N69012, N69011, N69010, N69009, N69008, N69007, N69006, N69005, 
        N69004, N69003}), .B({1'b0, 1'b0, 1'b0, N69025, N69024, N69023, N69022, 
        N69021, N69020, N69019, N69018, N69017, N69016}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, N69143, N69142, 
        N69141, N69140, N69139, N69138, N69137, N69136, N69135, N69134, N69133}) );
  hamming_N16000_CC2_DW01_add_10 add_2676_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68985, N68984, N68983, N68982, N68981, N68980, N68979, 
        N68978, N68977}), .B({1'b0, 1'b0, 1'b0, N68999, N68998, N68997, N68996, 
        N68995, N68994, N68993, N68992, N68991, N68990}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, N69130, N69129, 
        N69128, N69127, N69126, N69125, N69124, N69123, N69122, N69121, N69120}) );
  hamming_N16000_CC2_DW01_add_11 add_2677_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68959, N68958, N68957, N68956, N68955, N68954, N68953, 
        N68952, N68951}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68972, N68971, N68970, 
        N68969, N68968, N68967, N68966, N68965, N68964}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N69116, N69115, N69114, N69113, N69112, 
        N69111, N69110, N69109, N69108, N69107}) );
  hamming_N16000_CC2_DW01_add_12 add_2678_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68933, N68932, N68931, N68930, N68929, N68928, N68927, 
        N68926, N68925}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68946, N68945, N68944, 
        N68943, N68942, N68941, N68940, N68939, N68938}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, N69103, N69102, N69101, N69100, N69099, 
        N69098, N69097, N69096, N69095, N69094}) );
  hamming_N16000_CC2_DW01_add_13 add_2679_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68907, N68906, N68905, N68904, N68903, N68902, N68901, 
        N68900, N68899}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68920, N68919, N68918, 
        N68917, N68916, N68915, N68914, N68913, N68912}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, N69090, N69089, N69088, N69087, N69086, 
        N69085, N69084, N69083, N69082, N69081}) );
  hamming_N16000_CC2_DW01_add_14 add_2680_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68881, N68880, N68879, N68878, N68877, N68876, N68875, 
        N68874, N68873}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68894, N68893, N68892, 
        N68891, N68890, N68889, N68888, N68887, N68886}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, N69077, N69076, N69075, N69074, N69073, 
        N69072, N69071, N69070, N69069, N69068}) );
  hamming_N16000_CC2_DW01_add_15 add_2681_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68855, N68854, N68853, N68852, N68851, N68850, N68849, 
        N68848, N68847}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68868, N68867, N68866, 
        N68865, N68864, N68863, N68862, N68861, N68860}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, N69064, N69063, N69062, N69061, N69060, 
        N69059, N69058, N69057, N69056, N69055}) );
  hamming_N16000_CC2_DW01_add_16 add_2682_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68829, N68828, N68827, N68826, N68825, N68824, N68823, 
        N68822, N68821}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68842, N68841, N68840, 
        N68839, N68838, N68837, N68836, N68835, N68834}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, N69051, N69050, N69049, N69048, N69047, 
        N69046, N69045, N69044, N69043, N69042}) );
  hamming_N16000_CC2_DW01_add_17 add_2683_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68803, N68802, N68801, N68800, N68799, N68798, N68797, 
        N68796, N68795}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68816, N68815, N68814, 
        N68813, N68812, N68811, N68810, N68809, N68808}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, N69038, N69037, N69036, N69035, N69034, 
        N69033, N69032, N69031, N69030, N69029}) );
  hamming_N16000_CC2_DW01_add_18 add_2684_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68777, N68776, N68775, N68774, N68773, N68772, N68771, 
        N68770, N68769}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68790, N68789, N68788, 
        N68787, N68786, N68785, N68784, N68783, N68782}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, N69025, N69024, N69023, N69022, N69021, 
        N69020, N69019, N69018, N69017, N69016}) );
  hamming_N16000_CC2_DW01_add_19 add_2685_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68751, N68750, N68749, N68748, N68747, N68746, N68745, 
        N68744, N68743}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68764, N68763, N68762, 
        N68761, N68760, N68759, N68758, N68757, N68756}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, N69012, N69011, N69010, N69009, N69008, 
        N69007, N69006, N69005, N69004, N69003}) );
  hamming_N16000_CC2_DW01_add_20 add_2686_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68725, N68724, N68723, N68722, N68721, N68720, N68719, 
        N68718, N68717}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68738, N68737, N68736, 
        N68735, N68734, N68733, N68732, N68731, N68730}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, N68999, N68998, N68997, N68996, N68995, 
        N68994, N68993, N68992, N68991, N68990}) );
  hamming_N16000_CC2_DW01_add_21 add_2687_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68698, N68697, N68696, N68695, N68694, N68693, 
        N68692, N68691}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68711, N68710, 
        N68709, N68708, N68707, N68706, N68705, N68704}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, N68985, N68984, 
        N68983, N68982, N68981, N68980, N68979, N68978, N68977}) );
  hamming_N16000_CC2_DW01_add_22 add_2688_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68672, N68671, N68670, N68669, N68668, N68667, 
        N68666, N68665}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68685, N68684, 
        N68683, N68682, N68681, N68680, N68679, N68678}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, N68972, N68971, 
        N68970, N68969, N68968, N68967, N68966, N68965, N68964}) );
  hamming_N16000_CC2_DW01_add_23 add_2689_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68646, N68645, N68644, N68643, N68642, N68641, 
        N68640, N68639}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68659, N68658, 
        N68657, N68656, N68655, N68654, N68653, N68652}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, N68959, N68958, 
        N68957, N68956, N68955, N68954, N68953, N68952, N68951}) );
  hamming_N16000_CC2_DW01_add_24 add_2690_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68620, N68619, N68618, N68617, N68616, N68615, 
        N68614, N68613}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68633, N68632, 
        N68631, N68630, N68629, N68628, N68627, N68626}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, N68946, N68945, 
        N68944, N68943, N68942, N68941, N68940, N68939, N68938}) );
  hamming_N16000_CC2_DW01_add_25 add_2691_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68594, N68593, N68592, N68591, N68590, N68589, 
        N68588, N68587}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68607, N68606, 
        N68605, N68604, N68603, N68602, N68601, N68600}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, N68933, N68932, 
        N68931, N68930, N68929, N68928, N68927, N68926, N68925}) );
  hamming_N16000_CC2_DW01_add_26 add_2692_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68568, N68567, N68566, N68565, N68564, N68563, 
        N68562, N68561}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68581, N68580, 
        N68579, N68578, N68577, N68576, N68575, N68574}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, N68920, N68919, 
        N68918, N68917, N68916, N68915, N68914, N68913, N68912}) );
  hamming_N16000_CC2_DW01_add_27 add_2693_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68542, N68541, N68540, N68539, N68538, N68537, 
        N68536, N68535}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68555, N68554, 
        N68553, N68552, N68551, N68550, N68549, N68548}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, N68907, N68906, 
        N68905, N68904, N68903, N68902, N68901, N68900, N68899}) );
  hamming_N16000_CC2_DW01_add_28 add_2694_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68516, N68515, N68514, N68513, N68512, N68511, 
        N68510, N68509}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68529, N68528, 
        N68527, N68526, N68525, N68524, N68523, N68522}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, N68894, N68893, 
        N68892, N68891, N68890, N68889, N68888, N68887, N68886}) );
  hamming_N16000_CC2_DW01_add_29 add_2695_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68490, N68489, N68488, N68487, N68486, N68485, 
        N68484, N68483}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68503, N68502, 
        N68501, N68500, N68499, N68498, N68497, N68496}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, N68881, N68880, 
        N68879, N68878, N68877, N68876, N68875, N68874, N68873}) );
  hamming_N16000_CC2_DW01_add_30 add_2696_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68464, N68463, N68462, N68461, N68460, N68459, 
        N68458, N68457}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68477, N68476, 
        N68475, N68474, N68473, N68472, N68471, N68470}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, N68868, N68867, 
        N68866, N68865, N68864, N68863, N68862, N68861, N68860}) );
  hamming_N16000_CC2_DW01_add_31 add_2697_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68438, N68437, N68436, N68435, N68434, N68433, 
        N68432, N68431}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68451, N68450, 
        N68449, N68448, N68447, N68446, N68445, N68444}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, N68855, N68854, 
        N68853, N68852, N68851, N68850, N68849, N68848, N68847}) );
  hamming_N16000_CC2_DW01_add_32 add_2698_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68412, N68411, N68410, N68409, N68408, N68407, 
        N68406, N68405}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68425, N68424, 
        N68423, N68422, N68421, N68420, N68419, N68418}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, N68842, N68841, 
        N68840, N68839, N68838, N68837, N68836, N68835, N68834}) );
  hamming_N16000_CC2_DW01_add_33 add_2699_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68386, N68385, N68384, N68383, N68382, N68381, 
        N68380, N68379}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68399, N68398, 
        N68397, N68396, N68395, N68394, N68393, N68392}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, N68829, N68828, 
        N68827, N68826, N68825, N68824, N68823, N68822, N68821}) );
  hamming_N16000_CC2_DW01_add_34 add_2700_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68360, N68359, N68358, N68357, N68356, N68355, 
        N68354, N68353}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68373, N68372, 
        N68371, N68370, N68369, N68368, N68367, N68366}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, N68816, N68815, 
        N68814, N68813, N68812, N68811, N68810, N68809, N68808}) );
  hamming_N16000_CC2_DW01_add_35 add_2701_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68334, N68333, N68332, N68331, N68330, N68329, 
        N68328, N68327}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68347, N68346, 
        N68345, N68344, N68343, N68342, N68341, N68340}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, N68803, N68802, 
        N68801, N68800, N68799, N68798, N68797, N68796, N68795}) );
  hamming_N16000_CC2_DW01_add_36 add_2702_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68308, N68307, N68306, N68305, N68304, N68303, 
        N68302, N68301}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68321, N68320, 
        N68319, N68318, N68317, N68316, N68315, N68314}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, N68790, N68789, 
        N68788, N68787, N68786, N68785, N68784, N68783, N68782}) );
  hamming_N16000_CC2_DW01_add_37 add_2703_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68282, N68281, N68280, N68279, N68278, N68277, 
        N68276, N68275}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68295, N68294, 
        N68293, N68292, N68291, N68290, N68289, N68288}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, N68777, N68776, 
        N68775, N68774, N68773, N68772, N68771, N68770, N68769}) );
  hamming_N16000_CC2_DW01_add_38 add_2704_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68256, N68255, N68254, N68253, N68252, N68251, 
        N68250, N68249}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68269, N68268, 
        N68267, N68266, N68265, N68264, N68263, N68262}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, N68764, N68763, 
        N68762, N68761, N68760, N68759, N68758, N68757, N68756}) );
  hamming_N16000_CC2_DW01_add_39 add_2705_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68230, N68229, N68228, N68227, N68226, N68225, 
        N68224, N68223}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68243, N68242, 
        N68241, N68240, N68239, N68238, N68237, N68236}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, N68751, N68750, 
        N68749, N68748, N68747, N68746, N68745, N68744, N68743}) );
  hamming_N16000_CC2_DW01_add_40 add_2706_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68204, N68203, N68202, N68201, N68200, N68199, 
        N68198, N68197}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68217, N68216, 
        N68215, N68214, N68213, N68212, N68211, N68210}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, N68738, N68737, 
        N68736, N68735, N68734, N68733, N68732, N68731, N68730}) );
  hamming_N16000_CC2_DW01_add_41 add_2707_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68178, N68177, N68176, N68175, N68174, N68173, 
        N68172, N68171}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68191, N68190, 
        N68189, N68188, N68187, N68186, N68185, N68184}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, N68725, N68724, 
        N68723, N68722, N68721, N68720, N68719, N68718, N68717}) );
  hamming_N16000_CC2_DW01_add_42 add_2708_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68151, N68150, N68149, N68148, N68147, N68146, 
        N68145}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68164, N68163, 
        N68162, N68161, N68160, N68159, N68158}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, N68711, N68710, N68709, N68708, N68707, 
        N68706, N68705, N68704}) );
  hamming_N16000_CC2_DW01_add_43 add_2709_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68125, N68124, N68123, N68122, N68121, N68120, 
        N68119}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68138, N68137, 
        N68136, N68135, N68134, N68133, N68132}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, N68698, N68697, N68696, N68695, N68694, 
        N68693, N68692, N68691}) );
  hamming_N16000_CC2_DW01_add_44 add_2710_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68099, N68098, N68097, N68096, N68095, N68094, 
        N68093}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68112, N68111, 
        N68110, N68109, N68108, N68107, N68106}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__137, SYNOPSYS_UNCONNECTED__138, 
        SYNOPSYS_UNCONNECTED__139, SYNOPSYS_UNCONNECTED__140, 
        SYNOPSYS_UNCONNECTED__141, N68685, N68684, N68683, N68682, N68681, 
        N68680, N68679, N68678}) );
  hamming_N16000_CC2_DW01_add_45 add_2711_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68073, N68072, N68071, N68070, N68069, N68068, 
        N68067}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68086, N68085, 
        N68084, N68083, N68082, N68081, N68080}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, N68672, N68671, N68670, N68669, N68668, 
        N68667, N68666, N68665}) );
  hamming_N16000_CC2_DW01_add_46 add_2712_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68047, N68046, N68045, N68044, N68043, N68042, 
        N68041}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68060, N68059, 
        N68058, N68057, N68056, N68055, N68054}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__147, SYNOPSYS_UNCONNECTED__148, 
        SYNOPSYS_UNCONNECTED__149, SYNOPSYS_UNCONNECTED__150, 
        SYNOPSYS_UNCONNECTED__151, N68659, N68658, N68657, N68656, N68655, 
        N68654, N68653, N68652}) );
  hamming_N16000_CC2_DW01_add_47 add_2713_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68021, N68020, N68019, N68018, N68017, N68016, 
        N68015}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68034, N68033, 
        N68032, N68031, N68030, N68029, N68028}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, N68646, N68645, N68644, N68643, N68642, 
        N68641, N68640, N68639}) );
  hamming_N16000_CC2_DW01_add_48 add_2714_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67995, N67994, N67993, N67992, N67991, N67990, 
        N67989}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68008, N68007, 
        N68006, N68005, N68004, N68003, N68002}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, 
        SYNOPSYS_UNCONNECTED__159, SYNOPSYS_UNCONNECTED__160, 
        SYNOPSYS_UNCONNECTED__161, N68633, N68632, N68631, N68630, N68629, 
        N68628, N68627, N68626}) );
  hamming_N16000_CC2_DW01_add_49 add_2715_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67969, N67968, N67967, N67966, N67965, N67964, 
        N67963}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67982, N67981, 
        N67980, N67979, N67978, N67977, N67976}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, N68620, N68619, N68618, N68617, N68616, 
        N68615, N68614, N68613}) );
  hamming_N16000_CC2_DW01_add_50 add_2716_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67943, N67942, N67941, N67940, N67939, N67938, 
        N67937}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67956, N67955, 
        N67954, N67953, N67952, N67951, N67950}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__167, SYNOPSYS_UNCONNECTED__168, 
        SYNOPSYS_UNCONNECTED__169, SYNOPSYS_UNCONNECTED__170, 
        SYNOPSYS_UNCONNECTED__171, N68607, N68606, N68605, N68604, N68603, 
        N68602, N68601, N68600}) );
  hamming_N16000_CC2_DW01_add_51 add_2717_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67917, N67916, N67915, N67914, N67913, N67912, 
        N67911}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67930, N67929, 
        N67928, N67927, N67926, N67925, N67924}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, N68594, N68593, N68592, N68591, N68590, 
        N68589, N68588, N68587}) );
  hamming_N16000_CC2_DW01_add_52 add_2718_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67891, N67890, N67889, N67888, N67887, N67886, 
        N67885}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67904, N67903, 
        N67902, N67901, N67900, N67899, N67898}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__177, SYNOPSYS_UNCONNECTED__178, 
        SYNOPSYS_UNCONNECTED__179, SYNOPSYS_UNCONNECTED__180, 
        SYNOPSYS_UNCONNECTED__181, N68581, N68580, N68579, N68578, N68577, 
        N68576, N68575, N68574}) );
  hamming_N16000_CC2_DW01_add_53 add_2719_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67865, N67864, N67863, N67862, N67861, N67860, 
        N67859}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67878, N67877, 
        N67876, N67875, N67874, N67873, N67872}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, N68568, N68567, N68566, N68565, N68564, 
        N68563, N68562, N68561}) );
  hamming_N16000_CC2_DW01_add_54 add_2720_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67839, N67838, N67837, N67836, N67835, N67834, 
        N67833}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67852, N67851, 
        N67850, N67849, N67848, N67847, N67846}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__187, SYNOPSYS_UNCONNECTED__188, 
        SYNOPSYS_UNCONNECTED__189, SYNOPSYS_UNCONNECTED__190, 
        SYNOPSYS_UNCONNECTED__191, N68555, N68554, N68553, N68552, N68551, 
        N68550, N68549, N68548}) );
  hamming_N16000_CC2_DW01_add_55 add_2721_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67813, N67812, N67811, N67810, N67809, N67808, 
        N67807}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67826, N67825, 
        N67824, N67823, N67822, N67821, N67820}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, N68542, N68541, N68540, N68539, N68538, 
        N68537, N68536, N68535}) );
  hamming_N16000_CC2_DW01_add_56 add_2722_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67787, N67786, N67785, N67784, N67783, N67782, 
        N67781}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67800, N67799, 
        N67798, N67797, N67796, N67795, N67794}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__197, SYNOPSYS_UNCONNECTED__198, 
        SYNOPSYS_UNCONNECTED__199, SYNOPSYS_UNCONNECTED__200, 
        SYNOPSYS_UNCONNECTED__201, N68529, N68528, N68527, N68526, N68525, 
        N68524, N68523, N68522}) );
  hamming_N16000_CC2_DW01_add_57 add_2723_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67761, N67760, N67759, N67758, N67757, N67756, 
        N67755}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67774, N67773, 
        N67772, N67771, N67770, N67769, N67768}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, N68516, N68515, N68514, N68513, N68512, 
        N68511, N68510, N68509}) );
  hamming_N16000_CC2_DW01_add_58 add_2724_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67735, N67734, N67733, N67732, N67731, N67730, 
        N67729}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67748, N67747, 
        N67746, N67745, N67744, N67743, N67742}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__207, SYNOPSYS_UNCONNECTED__208, 
        SYNOPSYS_UNCONNECTED__209, SYNOPSYS_UNCONNECTED__210, 
        SYNOPSYS_UNCONNECTED__211, N68503, N68502, N68501, N68500, N68499, 
        N68498, N68497, N68496}) );
  hamming_N16000_CC2_DW01_add_59 add_2725_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67709, N67708, N67707, N67706, N67705, N67704, 
        N67703}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67722, N67721, 
        N67720, N67719, N67718, N67717, N67716}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, N68490, N68489, N68488, N68487, N68486, 
        N68485, N68484, N68483}) );
  hamming_N16000_CC2_DW01_add_60 add_2726_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67683, N67682, N67681, N67680, N67679, N67678, 
        N67677}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67696, N67695, 
        N67694, N67693, N67692, N67691, N67690}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__217, SYNOPSYS_UNCONNECTED__218, 
        SYNOPSYS_UNCONNECTED__219, SYNOPSYS_UNCONNECTED__220, 
        SYNOPSYS_UNCONNECTED__221, N68477, N68476, N68475, N68474, N68473, 
        N68472, N68471, N68470}) );
  hamming_N16000_CC2_DW01_add_61 add_2727_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67657, N67656, N67655, N67654, N67653, N67652, 
        N67651}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67670, N67669, 
        N67668, N67667, N67666, N67665, N67664}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, N68464, N68463, N68462, N68461, N68460, 
        N68459, N68458, N68457}) );
  hamming_N16000_CC2_DW01_add_62 add_2728_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67631, N67630, N67629, N67628, N67627, N67626, 
        N67625}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67644, N67643, 
        N67642, N67641, N67640, N67639, N67638}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__227, SYNOPSYS_UNCONNECTED__228, 
        SYNOPSYS_UNCONNECTED__229, SYNOPSYS_UNCONNECTED__230, 
        SYNOPSYS_UNCONNECTED__231, N68451, N68450, N68449, N68448, N68447, 
        N68446, N68445, N68444}) );
  hamming_N16000_CC2_DW01_add_63 add_2729_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67605, N67604, N67603, N67602, N67601, N67600, 
        N67599}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67618, N67617, 
        N67616, N67615, N67614, N67613, N67612}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, N68438, N68437, N68436, N68435, N68434, 
        N68433, N68432, N68431}) );
  hamming_N16000_CC2_DW01_add_64 add_2730_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67579, N67578, N67577, N67576, N67575, N67574, 
        N67573}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67592, N67591, 
        N67590, N67589, N67588, N67587, N67586}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__237, SYNOPSYS_UNCONNECTED__238, 
        SYNOPSYS_UNCONNECTED__239, SYNOPSYS_UNCONNECTED__240, 
        SYNOPSYS_UNCONNECTED__241, N68425, N68424, N68423, N68422, N68421, 
        N68420, N68419, N68418}) );
  hamming_N16000_CC2_DW01_add_65 add_2731_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67553, N67552, N67551, N67550, N67549, N67548, 
        N67547}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67566, N67565, 
        N67564, N67563, N67562, N67561, N67560}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, N68412, N68411, N68410, N68409, N68408, 
        N68407, N68406, N68405}) );
  hamming_N16000_CC2_DW01_add_66 add_2732_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67527, N67526, N67525, N67524, N67523, N67522, 
        N67521}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67540, N67539, 
        N67538, N67537, N67536, N67535, N67534}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__247, SYNOPSYS_UNCONNECTED__248, 
        SYNOPSYS_UNCONNECTED__249, SYNOPSYS_UNCONNECTED__250, 
        SYNOPSYS_UNCONNECTED__251, N68399, N68398, N68397, N68396, N68395, 
        N68394, N68393, N68392}) );
  hamming_N16000_CC2_DW01_add_67 add_2733_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67501, N67500, N67499, N67498, N67497, N67496, 
        N67495}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67514, N67513, 
        N67512, N67511, N67510, N67509, N67508}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, N68386, N68385, N68384, N68383, N68382, 
        N68381, N68380, N68379}) );
  hamming_N16000_CC2_DW01_add_68 add_2734_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67475, N67474, N67473, N67472, N67471, N67470, 
        N67469}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67488, N67487, 
        N67486, N67485, N67484, N67483, N67482}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__257, SYNOPSYS_UNCONNECTED__258, 
        SYNOPSYS_UNCONNECTED__259, SYNOPSYS_UNCONNECTED__260, 
        SYNOPSYS_UNCONNECTED__261, N68373, N68372, N68371, N68370, N68369, 
        N68368, N68367, N68366}) );
  hamming_N16000_CC2_DW01_add_69 add_2735_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67449, N67448, N67447, N67446, N67445, N67444, 
        N67443}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67462, N67461, 
        N67460, N67459, N67458, N67457, N67456}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, N68360, N68359, N68358, N68357, N68356, 
        N68355, N68354, N68353}) );
  hamming_N16000_CC2_DW01_add_70 add_2736_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67423, N67422, N67421, N67420, N67419, N67418, 
        N67417}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67436, N67435, 
        N67434, N67433, N67432, N67431, N67430}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__267, SYNOPSYS_UNCONNECTED__268, 
        SYNOPSYS_UNCONNECTED__269, SYNOPSYS_UNCONNECTED__270, 
        SYNOPSYS_UNCONNECTED__271, N68347, N68346, N68345, N68344, N68343, 
        N68342, N68341, N68340}) );
  hamming_N16000_CC2_DW01_add_71 add_2737_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67397, N67396, N67395, N67394, N67393, N67392, 
        N67391}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67410, N67409, 
        N67408, N67407, N67406, N67405, N67404}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, N68334, N68333, N68332, N68331, N68330, 
        N68329, N68328, N68327}) );
  hamming_N16000_CC2_DW01_add_72 add_2738_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67371, N67370, N67369, N67368, N67367, N67366, 
        N67365}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67384, N67383, 
        N67382, N67381, N67380, N67379, N67378}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__277, SYNOPSYS_UNCONNECTED__278, 
        SYNOPSYS_UNCONNECTED__279, SYNOPSYS_UNCONNECTED__280, 
        SYNOPSYS_UNCONNECTED__281, N68321, N68320, N68319, N68318, N68317, 
        N68316, N68315, N68314}) );
  hamming_N16000_CC2_DW01_add_73 add_2739_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67345, N67344, N67343, N67342, N67341, N67340, 
        N67339}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67358, N67357, 
        N67356, N67355, N67354, N67353, N67352}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, N68308, N68307, N68306, N68305, N68304, 
        N68303, N68302, N68301}) );
  hamming_N16000_CC2_DW01_add_74 add_2740_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67319, N67318, N67317, N67316, N67315, N67314, 
        N67313}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67332, N67331, 
        N67330, N67329, N67328, N67327, N67326}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__287, SYNOPSYS_UNCONNECTED__288, 
        SYNOPSYS_UNCONNECTED__289, SYNOPSYS_UNCONNECTED__290, 
        SYNOPSYS_UNCONNECTED__291, N68295, N68294, N68293, N68292, N68291, 
        N68290, N68289, N68288}) );
  hamming_N16000_CC2_DW01_add_75 add_2741_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67293, N67292, N67291, N67290, N67289, N67288, 
        N67287}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67306, N67305, 
        N67304, N67303, N67302, N67301, N67300}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, N68282, N68281, N68280, N68279, N68278, 
        N68277, N68276, N68275}) );
  hamming_N16000_CC2_DW01_add_76 add_2742_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67267, N67266, N67265, N67264, N67263, N67262, 
        N67261}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67280, N67279, 
        N67278, N67277, N67276, N67275, N67274}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__297, SYNOPSYS_UNCONNECTED__298, 
        SYNOPSYS_UNCONNECTED__299, SYNOPSYS_UNCONNECTED__300, 
        SYNOPSYS_UNCONNECTED__301, N68269, N68268, N68267, N68266, N68265, 
        N68264, N68263, N68262}) );
  hamming_N16000_CC2_DW01_add_77 add_2743_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67241, N67240, N67239, N67238, N67237, N67236, 
        N67235}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67254, N67253, 
        N67252, N67251, N67250, N67249, N67248}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, N68256, N68255, N68254, N68253, N68252, 
        N68251, N68250, N68249}) );
  hamming_N16000_CC2_DW01_add_78 add_2744_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67215, N67214, N67213, N67212, N67211, N67210, 
        N67209}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67228, N67227, 
        N67226, N67225, N67224, N67223, N67222}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__307, SYNOPSYS_UNCONNECTED__308, 
        SYNOPSYS_UNCONNECTED__309, SYNOPSYS_UNCONNECTED__310, 
        SYNOPSYS_UNCONNECTED__311, N68243, N68242, N68241, N68240, N68239, 
        N68238, N68237, N68236}) );
  hamming_N16000_CC2_DW01_add_79 add_2745_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67189, N67188, N67187, N67186, N67185, N67184, 
        N67183}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67202, N67201, 
        N67200, N67199, N67198, N67197, N67196}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, N68230, N68229, N68228, N68227, N68226, 
        N68225, N68224, N68223}) );
  hamming_N16000_CC2_DW01_add_80 add_2746_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67163, N67162, N67161, N67160, N67159, N67158, 
        N67157}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67176, N67175, 
        N67174, N67173, N67172, N67171, N67170}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__317, SYNOPSYS_UNCONNECTED__318, 
        SYNOPSYS_UNCONNECTED__319, SYNOPSYS_UNCONNECTED__320, 
        SYNOPSYS_UNCONNECTED__321, N68217, N68216, N68215, N68214, N68213, 
        N68212, N68211, N68210}) );
  hamming_N16000_CC2_DW01_add_81 add_2747_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67137, N67136, N67135, N67134, N67133, N67132, 
        N67131}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67150, N67149, 
        N67148, N67147, N67146, N67145, N67144}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, N68204, N68203, N68202, N68201, N68200, 
        N68199, N68198, N68197}) );
  hamming_N16000_CC2_DW01_add_82 add_2748_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67111, N67110, N67109, N67108, N67107, N67106, 
        N67105}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67124, N67123, 
        N67122, N67121, N67120, N67119, N67118}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__327, SYNOPSYS_UNCONNECTED__328, 
        SYNOPSYS_UNCONNECTED__329, SYNOPSYS_UNCONNECTED__330, 
        SYNOPSYS_UNCONNECTED__331, N68191, N68190, N68189, N68188, N68187, 
        N68186, N68185, N68184}) );
  hamming_N16000_CC2_DW01_add_83 add_2749_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67084, N67083, N67082, N67081, N67080, 
        N67079}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67098, N67097, 
        N67096, N67095, N67094, N67093, N67092}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, N68178, N68177, N68176, N68175, N68174, 
        N68173, N68172, N68171}) );
  hamming_N16000_CC2_DW01_add_84 add_2750_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67058, N67057, N67056, N67055, N67054, 
        N67053}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67071, N67070, 
        N67069, N67068, N67067, N67066}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__337, SYNOPSYS_UNCONNECTED__338, 
        SYNOPSYS_UNCONNECTED__339, SYNOPSYS_UNCONNECTED__340, 
        SYNOPSYS_UNCONNECTED__341, SYNOPSYS_UNCONNECTED__342, N68164, N68163, 
        N68162, N68161, N68160, N68159, N68158}) );
  hamming_N16000_CC2_DW01_add_85 add_2751_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67032, N67031, N67030, N67029, N67028, 
        N67027}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67045, N67044, 
        N67043, N67042, N67041, N67040}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__343, SYNOPSYS_UNCONNECTED__344, 
        SYNOPSYS_UNCONNECTED__345, SYNOPSYS_UNCONNECTED__346, 
        SYNOPSYS_UNCONNECTED__347, SYNOPSYS_UNCONNECTED__348, N68151, N68150, 
        N68149, N68148, N68147, N68146, N68145}) );
  hamming_N16000_CC2_DW01_add_86 add_2752_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67006, N67005, N67004, N67003, N67002, 
        N67001}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67019, N67018, 
        N67017, N67016, N67015, N67014}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__349, SYNOPSYS_UNCONNECTED__350, 
        SYNOPSYS_UNCONNECTED__351, SYNOPSYS_UNCONNECTED__352, 
        SYNOPSYS_UNCONNECTED__353, SYNOPSYS_UNCONNECTED__354, N68138, N68137, 
        N68136, N68135, N68134, N68133, N68132}) );
  hamming_N16000_CC2_DW01_add_87 add_2753_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66980, N66979, N66978, N66977, N66976, 
        N66975}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66993, N66992, 
        N66991, N66990, N66989, N66988}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__355, SYNOPSYS_UNCONNECTED__356, 
        SYNOPSYS_UNCONNECTED__357, SYNOPSYS_UNCONNECTED__358, 
        SYNOPSYS_UNCONNECTED__359, SYNOPSYS_UNCONNECTED__360, N68125, N68124, 
        N68123, N68122, N68121, N68120, N68119}) );
  hamming_N16000_CC2_DW01_add_88 add_2754_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66954, N66953, N66952, N66951, N66950, 
        N66949}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66967, N66966, 
        N66965, N66964, N66963, N66962}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__361, SYNOPSYS_UNCONNECTED__362, 
        SYNOPSYS_UNCONNECTED__363, SYNOPSYS_UNCONNECTED__364, 
        SYNOPSYS_UNCONNECTED__365, SYNOPSYS_UNCONNECTED__366, N68112, N68111, 
        N68110, N68109, N68108, N68107, N68106}) );
  hamming_N16000_CC2_DW01_add_89 add_2755_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66928, N66927, N66926, N66925, N66924, 
        N66923}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66941, N66940, 
        N66939, N66938, N66937, N66936}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__367, SYNOPSYS_UNCONNECTED__368, 
        SYNOPSYS_UNCONNECTED__369, SYNOPSYS_UNCONNECTED__370, 
        SYNOPSYS_UNCONNECTED__371, SYNOPSYS_UNCONNECTED__372, N68099, N68098, 
        N68097, N68096, N68095, N68094, N68093}) );
  hamming_N16000_CC2_DW01_add_90 add_2756_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66902, N66901, N66900, N66899, N66898, 
        N66897}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66915, N66914, 
        N66913, N66912, N66911, N66910}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__373, SYNOPSYS_UNCONNECTED__374, 
        SYNOPSYS_UNCONNECTED__375, SYNOPSYS_UNCONNECTED__376, 
        SYNOPSYS_UNCONNECTED__377, SYNOPSYS_UNCONNECTED__378, N68086, N68085, 
        N68084, N68083, N68082, N68081, N68080}) );
  hamming_N16000_CC2_DW01_add_91 add_2757_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66876, N66875, N66874, N66873, N66872, 
        N66871}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66889, N66888, 
        N66887, N66886, N66885, N66884}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__379, SYNOPSYS_UNCONNECTED__380, 
        SYNOPSYS_UNCONNECTED__381, SYNOPSYS_UNCONNECTED__382, 
        SYNOPSYS_UNCONNECTED__383, SYNOPSYS_UNCONNECTED__384, N68073, N68072, 
        N68071, N68070, N68069, N68068, N68067}) );
  hamming_N16000_CC2_DW01_add_92 add_2758_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66850, N66849, N66848, N66847, N66846, 
        N66845}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66863, N66862, 
        N66861, N66860, N66859, N66858}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__385, SYNOPSYS_UNCONNECTED__386, 
        SYNOPSYS_UNCONNECTED__387, SYNOPSYS_UNCONNECTED__388, 
        SYNOPSYS_UNCONNECTED__389, SYNOPSYS_UNCONNECTED__390, N68060, N68059, 
        N68058, N68057, N68056, N68055, N68054}) );
  hamming_N16000_CC2_DW01_add_93 add_2759_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66824, N66823, N66822, N66821, N66820, 
        N66819}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66837, N66836, 
        N66835, N66834, N66833, N66832}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__391, SYNOPSYS_UNCONNECTED__392, 
        SYNOPSYS_UNCONNECTED__393, SYNOPSYS_UNCONNECTED__394, 
        SYNOPSYS_UNCONNECTED__395, SYNOPSYS_UNCONNECTED__396, N68047, N68046, 
        N68045, N68044, N68043, N68042, N68041}) );
  hamming_N16000_CC2_DW01_add_94 add_2760_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66798, N66797, N66796, N66795, N66794, 
        N66793}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66811, N66810, 
        N66809, N66808, N66807, N66806}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__397, SYNOPSYS_UNCONNECTED__398, 
        SYNOPSYS_UNCONNECTED__399, SYNOPSYS_UNCONNECTED__400, 
        SYNOPSYS_UNCONNECTED__401, SYNOPSYS_UNCONNECTED__402, N68034, N68033, 
        N68032, N68031, N68030, N68029, N68028}) );
  hamming_N16000_CC2_DW01_add_95 add_2761_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66772, N66771, N66770, N66769, N66768, 
        N66767}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66785, N66784, 
        N66783, N66782, N66781, N66780}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__403, SYNOPSYS_UNCONNECTED__404, 
        SYNOPSYS_UNCONNECTED__405, SYNOPSYS_UNCONNECTED__406, 
        SYNOPSYS_UNCONNECTED__407, SYNOPSYS_UNCONNECTED__408, N68021, N68020, 
        N68019, N68018, N68017, N68016, N68015}) );
  hamming_N16000_CC2_DW01_add_96 add_2762_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66746, N66745, N66744, N66743, N66742, 
        N66741}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66759, N66758, 
        N66757, N66756, N66755, N66754}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__409, SYNOPSYS_UNCONNECTED__410, 
        SYNOPSYS_UNCONNECTED__411, SYNOPSYS_UNCONNECTED__412, 
        SYNOPSYS_UNCONNECTED__413, SYNOPSYS_UNCONNECTED__414, N68008, N68007, 
        N68006, N68005, N68004, N68003, N68002}) );
  hamming_N16000_CC2_DW01_add_97 add_2763_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66720, N66719, N66718, N66717, N66716, 
        N66715}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66733, N66732, 
        N66731, N66730, N66729, N66728}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__415, SYNOPSYS_UNCONNECTED__416, 
        SYNOPSYS_UNCONNECTED__417, SYNOPSYS_UNCONNECTED__418, 
        SYNOPSYS_UNCONNECTED__419, SYNOPSYS_UNCONNECTED__420, N67995, N67994, 
        N67993, N67992, N67991, N67990, N67989}) );
  hamming_N16000_CC2_DW01_add_98 add_2764_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66694, N66693, N66692, N66691, N66690, 
        N66689}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66707, N66706, 
        N66705, N66704, N66703, N66702}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__421, SYNOPSYS_UNCONNECTED__422, 
        SYNOPSYS_UNCONNECTED__423, SYNOPSYS_UNCONNECTED__424, 
        SYNOPSYS_UNCONNECTED__425, SYNOPSYS_UNCONNECTED__426, N67982, N67981, 
        N67980, N67979, N67978, N67977, N67976}) );
  hamming_N16000_CC2_DW01_add_99 add_2765_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66668, N66667, N66666, N66665, N66664, 
        N66663}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66681, N66680, 
        N66679, N66678, N66677, N66676}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__427, SYNOPSYS_UNCONNECTED__428, 
        SYNOPSYS_UNCONNECTED__429, SYNOPSYS_UNCONNECTED__430, 
        SYNOPSYS_UNCONNECTED__431, SYNOPSYS_UNCONNECTED__432, N67969, N67968, 
        N67967, N67966, N67965, N67964, N67963}) );
  hamming_N16000_CC2_DW01_add_100 add_2766_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66642, N66641, N66640, N66639, N66638, 
        N66637}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66655, N66654, 
        N66653, N66652, N66651, N66650}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__433, SYNOPSYS_UNCONNECTED__434, 
        SYNOPSYS_UNCONNECTED__435, SYNOPSYS_UNCONNECTED__436, 
        SYNOPSYS_UNCONNECTED__437, SYNOPSYS_UNCONNECTED__438, N67956, N67955, 
        N67954, N67953, N67952, N67951, N67950}) );
  hamming_N16000_CC2_DW01_add_101 add_2767_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66616, N66615, N66614, N66613, N66612, 
        N66611}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66629, N66628, 
        N66627, N66626, N66625, N66624}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__439, SYNOPSYS_UNCONNECTED__440, 
        SYNOPSYS_UNCONNECTED__441, SYNOPSYS_UNCONNECTED__442, 
        SYNOPSYS_UNCONNECTED__443, SYNOPSYS_UNCONNECTED__444, N67943, N67942, 
        N67941, N67940, N67939, N67938, N67937}) );
  hamming_N16000_CC2_DW01_add_102 add_2768_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66590, N66589, N66588, N66587, N66586, 
        N66585}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66603, N66602, 
        N66601, N66600, N66599, N66598}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__445, SYNOPSYS_UNCONNECTED__446, 
        SYNOPSYS_UNCONNECTED__447, SYNOPSYS_UNCONNECTED__448, 
        SYNOPSYS_UNCONNECTED__449, SYNOPSYS_UNCONNECTED__450, N67930, N67929, 
        N67928, N67927, N67926, N67925, N67924}) );
  hamming_N16000_CC2_DW01_add_103 add_2769_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66564, N66563, N66562, N66561, N66560, 
        N66559}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66577, N66576, 
        N66575, N66574, N66573, N66572}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__451, SYNOPSYS_UNCONNECTED__452, 
        SYNOPSYS_UNCONNECTED__453, SYNOPSYS_UNCONNECTED__454, 
        SYNOPSYS_UNCONNECTED__455, SYNOPSYS_UNCONNECTED__456, N67917, N67916, 
        N67915, N67914, N67913, N67912, N67911}) );
  hamming_N16000_CC2_DW01_add_104 add_2770_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66538, N66537, N66536, N66535, N66534, 
        N66533}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66551, N66550, 
        N66549, N66548, N66547, N66546}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__457, SYNOPSYS_UNCONNECTED__458, 
        SYNOPSYS_UNCONNECTED__459, SYNOPSYS_UNCONNECTED__460, 
        SYNOPSYS_UNCONNECTED__461, SYNOPSYS_UNCONNECTED__462, N67904, N67903, 
        N67902, N67901, N67900, N67899, N67898}) );
  hamming_N16000_CC2_DW01_add_105 add_2771_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66512, N66511, N66510, N66509, N66508, 
        N66507}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66525, N66524, 
        N66523, N66522, N66521, N66520}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__463, SYNOPSYS_UNCONNECTED__464, 
        SYNOPSYS_UNCONNECTED__465, SYNOPSYS_UNCONNECTED__466, 
        SYNOPSYS_UNCONNECTED__467, SYNOPSYS_UNCONNECTED__468, N67891, N67890, 
        N67889, N67888, N67887, N67886, N67885}) );
  hamming_N16000_CC2_DW01_add_106 add_2772_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66486, N66485, N66484, N66483, N66482, 
        N66481}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66499, N66498, 
        N66497, N66496, N66495, N66494}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__469, SYNOPSYS_UNCONNECTED__470, 
        SYNOPSYS_UNCONNECTED__471, SYNOPSYS_UNCONNECTED__472, 
        SYNOPSYS_UNCONNECTED__473, SYNOPSYS_UNCONNECTED__474, N67878, N67877, 
        N67876, N67875, N67874, N67873, N67872}) );
  hamming_N16000_CC2_DW01_add_107 add_2773_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66460, N66459, N66458, N66457, N66456, 
        N66455}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66473, N66472, 
        N66471, N66470, N66469, N66468}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__475, SYNOPSYS_UNCONNECTED__476, 
        SYNOPSYS_UNCONNECTED__477, SYNOPSYS_UNCONNECTED__478, 
        SYNOPSYS_UNCONNECTED__479, SYNOPSYS_UNCONNECTED__480, N67865, N67864, 
        N67863, N67862, N67861, N67860, N67859}) );
  hamming_N16000_CC2_DW01_add_108 add_2774_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66434, N66433, N66432, N66431, N66430, 
        N66429}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66447, N66446, 
        N66445, N66444, N66443, N66442}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__481, SYNOPSYS_UNCONNECTED__482, 
        SYNOPSYS_UNCONNECTED__483, SYNOPSYS_UNCONNECTED__484, 
        SYNOPSYS_UNCONNECTED__485, SYNOPSYS_UNCONNECTED__486, N67852, N67851, 
        N67850, N67849, N67848, N67847, N67846}) );
  hamming_N16000_CC2_DW01_add_109 add_2775_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66408, N66407, N66406, N66405, N66404, 
        N66403}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66421, N66420, 
        N66419, N66418, N66417, N66416}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__487, SYNOPSYS_UNCONNECTED__488, 
        SYNOPSYS_UNCONNECTED__489, SYNOPSYS_UNCONNECTED__490, 
        SYNOPSYS_UNCONNECTED__491, SYNOPSYS_UNCONNECTED__492, N67839, N67838, 
        N67837, N67836, N67835, N67834, N67833}) );
  hamming_N16000_CC2_DW01_add_110 add_2776_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66382, N66381, N66380, N66379, N66378, 
        N66377}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66395, N66394, 
        N66393, N66392, N66391, N66390}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__493, SYNOPSYS_UNCONNECTED__494, 
        SYNOPSYS_UNCONNECTED__495, SYNOPSYS_UNCONNECTED__496, 
        SYNOPSYS_UNCONNECTED__497, SYNOPSYS_UNCONNECTED__498, N67826, N67825, 
        N67824, N67823, N67822, N67821, N67820}) );
  hamming_N16000_CC2_DW01_add_111 add_2777_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66356, N66355, N66354, N66353, N66352, 
        N66351}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66369, N66368, 
        N66367, N66366, N66365, N66364}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__499, SYNOPSYS_UNCONNECTED__500, 
        SYNOPSYS_UNCONNECTED__501, SYNOPSYS_UNCONNECTED__502, 
        SYNOPSYS_UNCONNECTED__503, SYNOPSYS_UNCONNECTED__504, N67813, N67812, 
        N67811, N67810, N67809, N67808, N67807}) );
  hamming_N16000_CC2_DW01_add_112 add_2778_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66330, N66329, N66328, N66327, N66326, 
        N66325}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66343, N66342, 
        N66341, N66340, N66339, N66338}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__505, SYNOPSYS_UNCONNECTED__506, 
        SYNOPSYS_UNCONNECTED__507, SYNOPSYS_UNCONNECTED__508, 
        SYNOPSYS_UNCONNECTED__509, SYNOPSYS_UNCONNECTED__510, N67800, N67799, 
        N67798, N67797, N67796, N67795, N67794}) );
  hamming_N16000_CC2_DW01_add_113 add_2779_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66304, N66303, N66302, N66301, N66300, 
        N66299}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66317, N66316, 
        N66315, N66314, N66313, N66312}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__511, SYNOPSYS_UNCONNECTED__512, 
        SYNOPSYS_UNCONNECTED__513, SYNOPSYS_UNCONNECTED__514, 
        SYNOPSYS_UNCONNECTED__515, SYNOPSYS_UNCONNECTED__516, N67787, N67786, 
        N67785, N67784, N67783, N67782, N67781}) );
  hamming_N16000_CC2_DW01_add_114 add_2780_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66278, N66277, N66276, N66275, N66274, 
        N66273}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66291, N66290, 
        N66289, N66288, N66287, N66286}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__517, SYNOPSYS_UNCONNECTED__518, 
        SYNOPSYS_UNCONNECTED__519, SYNOPSYS_UNCONNECTED__520, 
        SYNOPSYS_UNCONNECTED__521, SYNOPSYS_UNCONNECTED__522, N67774, N67773, 
        N67772, N67771, N67770, N67769, N67768}) );
  hamming_N16000_CC2_DW01_add_115 add_2781_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66252, N66251, N66250, N66249, N66248, 
        N66247}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66265, N66264, 
        N66263, N66262, N66261, N66260}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__523, SYNOPSYS_UNCONNECTED__524, 
        SYNOPSYS_UNCONNECTED__525, SYNOPSYS_UNCONNECTED__526, 
        SYNOPSYS_UNCONNECTED__527, SYNOPSYS_UNCONNECTED__528, N67761, N67760, 
        N67759, N67758, N67757, N67756, N67755}) );
  hamming_N16000_CC2_DW01_add_116 add_2782_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66226, N66225, N66224, N66223, N66222, 
        N66221}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66239, N66238, 
        N66237, N66236, N66235, N66234}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__529, SYNOPSYS_UNCONNECTED__530, 
        SYNOPSYS_UNCONNECTED__531, SYNOPSYS_UNCONNECTED__532, 
        SYNOPSYS_UNCONNECTED__533, SYNOPSYS_UNCONNECTED__534, N67748, N67747, 
        N67746, N67745, N67744, N67743, N67742}) );
  hamming_N16000_CC2_DW01_add_117 add_2783_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66200, N66199, N66198, N66197, N66196, 
        N66195}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66213, N66212, 
        N66211, N66210, N66209, N66208}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__535, SYNOPSYS_UNCONNECTED__536, 
        SYNOPSYS_UNCONNECTED__537, SYNOPSYS_UNCONNECTED__538, 
        SYNOPSYS_UNCONNECTED__539, SYNOPSYS_UNCONNECTED__540, N67735, N67734, 
        N67733, N67732, N67731, N67730, N67729}) );
  hamming_N16000_CC2_DW01_add_118 add_2784_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66174, N66173, N66172, N66171, N66170, 
        N66169}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66187, N66186, 
        N66185, N66184, N66183, N66182}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__541, SYNOPSYS_UNCONNECTED__542, 
        SYNOPSYS_UNCONNECTED__543, SYNOPSYS_UNCONNECTED__544, 
        SYNOPSYS_UNCONNECTED__545, SYNOPSYS_UNCONNECTED__546, N67722, N67721, 
        N67720, N67719, N67718, N67717, N67716}) );
  hamming_N16000_CC2_DW01_add_119 add_2785_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66148, N66147, N66146, N66145, N66144, 
        N66143}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66161, N66160, 
        N66159, N66158, N66157, N66156}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__547, SYNOPSYS_UNCONNECTED__548, 
        SYNOPSYS_UNCONNECTED__549, SYNOPSYS_UNCONNECTED__550, 
        SYNOPSYS_UNCONNECTED__551, SYNOPSYS_UNCONNECTED__552, N67709, N67708, 
        N67707, N67706, N67705, N67704, N67703}) );
  hamming_N16000_CC2_DW01_add_120 add_2786_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66122, N66121, N66120, N66119, N66118, 
        N66117}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66135, N66134, 
        N66133, N66132, N66131, N66130}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__553, SYNOPSYS_UNCONNECTED__554, 
        SYNOPSYS_UNCONNECTED__555, SYNOPSYS_UNCONNECTED__556, 
        SYNOPSYS_UNCONNECTED__557, SYNOPSYS_UNCONNECTED__558, N67696, N67695, 
        N67694, N67693, N67692, N67691, N67690}) );
  hamming_N16000_CC2_DW01_add_121 add_2787_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66096, N66095, N66094, N66093, N66092, 
        N66091}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66109, N66108, 
        N66107, N66106, N66105, N66104}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__559, SYNOPSYS_UNCONNECTED__560, 
        SYNOPSYS_UNCONNECTED__561, SYNOPSYS_UNCONNECTED__562, 
        SYNOPSYS_UNCONNECTED__563, SYNOPSYS_UNCONNECTED__564, N67683, N67682, 
        N67681, N67680, N67679, N67678, N67677}) );
  hamming_N16000_CC2_DW01_add_122 add_2788_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66070, N66069, N66068, N66067, N66066, 
        N66065}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66083, N66082, 
        N66081, N66080, N66079, N66078}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__565, SYNOPSYS_UNCONNECTED__566, 
        SYNOPSYS_UNCONNECTED__567, SYNOPSYS_UNCONNECTED__568, 
        SYNOPSYS_UNCONNECTED__569, SYNOPSYS_UNCONNECTED__570, N67670, N67669, 
        N67668, N67667, N67666, N67665, N67664}) );
  hamming_N16000_CC2_DW01_add_123 add_2789_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66044, N66043, N66042, N66041, N66040, 
        N66039}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66057, N66056, 
        N66055, N66054, N66053, N66052}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__571, SYNOPSYS_UNCONNECTED__572, 
        SYNOPSYS_UNCONNECTED__573, SYNOPSYS_UNCONNECTED__574, 
        SYNOPSYS_UNCONNECTED__575, SYNOPSYS_UNCONNECTED__576, N67657, N67656, 
        N67655, N67654, N67653, N67652, N67651}) );
  hamming_N16000_CC2_DW01_add_124 add_2790_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66018, N66017, N66016, N66015, N66014, 
        N66013}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66031, N66030, 
        N66029, N66028, N66027, N66026}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__577, SYNOPSYS_UNCONNECTED__578, 
        SYNOPSYS_UNCONNECTED__579, SYNOPSYS_UNCONNECTED__580, 
        SYNOPSYS_UNCONNECTED__581, SYNOPSYS_UNCONNECTED__582, N67644, N67643, 
        N67642, N67641, N67640, N67639, N67638}) );
  hamming_N16000_CC2_DW01_add_125 add_2791_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65992, N65991, N65990, N65989, N65988, 
        N65987}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66005, N66004, 
        N66003, N66002, N66001, N66000}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__583, SYNOPSYS_UNCONNECTED__584, 
        SYNOPSYS_UNCONNECTED__585, SYNOPSYS_UNCONNECTED__586, 
        SYNOPSYS_UNCONNECTED__587, SYNOPSYS_UNCONNECTED__588, N67631, N67630, 
        N67629, N67628, N67627, N67626, N67625}) );
  hamming_N16000_CC2_DW01_add_126 add_2792_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65966, N65965, N65964, N65963, N65962, 
        N65961}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65979, N65978, 
        N65977, N65976, N65975, N65974}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__589, SYNOPSYS_UNCONNECTED__590, 
        SYNOPSYS_UNCONNECTED__591, SYNOPSYS_UNCONNECTED__592, 
        SYNOPSYS_UNCONNECTED__593, SYNOPSYS_UNCONNECTED__594, N67618, N67617, 
        N67616, N67615, N67614, N67613, N67612}) );
  hamming_N16000_CC2_DW01_add_127 add_2793_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65940, N65939, N65938, N65937, N65936, 
        N65935}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65953, N65952, 
        N65951, N65950, N65949, N65948}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__595, SYNOPSYS_UNCONNECTED__596, 
        SYNOPSYS_UNCONNECTED__597, SYNOPSYS_UNCONNECTED__598, 
        SYNOPSYS_UNCONNECTED__599, SYNOPSYS_UNCONNECTED__600, N67605, N67604, 
        N67603, N67602, N67601, N67600, N67599}) );
  hamming_N16000_CC2_DW01_add_128 add_2794_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65914, N65913, N65912, N65911, N65910, 
        N65909}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65927, N65926, 
        N65925, N65924, N65923, N65922}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__601, SYNOPSYS_UNCONNECTED__602, 
        SYNOPSYS_UNCONNECTED__603, SYNOPSYS_UNCONNECTED__604, 
        SYNOPSYS_UNCONNECTED__605, SYNOPSYS_UNCONNECTED__606, N67592, N67591, 
        N67590, N67589, N67588, N67587, N67586}) );
  hamming_N16000_CC2_DW01_add_129 add_2795_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65888, N65887, N65886, N65885, N65884, 
        N65883}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65901, N65900, 
        N65899, N65898, N65897, N65896}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__607, SYNOPSYS_UNCONNECTED__608, 
        SYNOPSYS_UNCONNECTED__609, SYNOPSYS_UNCONNECTED__610, 
        SYNOPSYS_UNCONNECTED__611, SYNOPSYS_UNCONNECTED__612, N67579, N67578, 
        N67577, N67576, N67575, N67574, N67573}) );
  hamming_N16000_CC2_DW01_add_130 add_2796_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65862, N65861, N65860, N65859, N65858, 
        N65857}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65875, N65874, 
        N65873, N65872, N65871, N65870}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__613, SYNOPSYS_UNCONNECTED__614, 
        SYNOPSYS_UNCONNECTED__615, SYNOPSYS_UNCONNECTED__616, 
        SYNOPSYS_UNCONNECTED__617, SYNOPSYS_UNCONNECTED__618, N67566, N67565, 
        N67564, N67563, N67562, N67561, N67560}) );
  hamming_N16000_CC2_DW01_add_131 add_2797_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65836, N65835, N65834, N65833, N65832, 
        N65831}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65849, N65848, 
        N65847, N65846, N65845, N65844}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__619, SYNOPSYS_UNCONNECTED__620, 
        SYNOPSYS_UNCONNECTED__621, SYNOPSYS_UNCONNECTED__622, 
        SYNOPSYS_UNCONNECTED__623, SYNOPSYS_UNCONNECTED__624, N67553, N67552, 
        N67551, N67550, N67549, N67548, N67547}) );
  hamming_N16000_CC2_DW01_add_132 add_2798_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65810, N65809, N65808, N65807, N65806, 
        N65805}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65823, N65822, 
        N65821, N65820, N65819, N65818}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__625, SYNOPSYS_UNCONNECTED__626, 
        SYNOPSYS_UNCONNECTED__627, SYNOPSYS_UNCONNECTED__628, 
        SYNOPSYS_UNCONNECTED__629, SYNOPSYS_UNCONNECTED__630, N67540, N67539, 
        N67538, N67537, N67536, N67535, N67534}) );
  hamming_N16000_CC2_DW01_add_133 add_2799_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65784, N65783, N65782, N65781, N65780, 
        N65779}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65797, N65796, 
        N65795, N65794, N65793, N65792}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__631, SYNOPSYS_UNCONNECTED__632, 
        SYNOPSYS_UNCONNECTED__633, SYNOPSYS_UNCONNECTED__634, 
        SYNOPSYS_UNCONNECTED__635, SYNOPSYS_UNCONNECTED__636, N67527, N67526, 
        N67525, N67524, N67523, N67522, N67521}) );
  hamming_N16000_CC2_DW01_add_134 add_2800_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65758, N65757, N65756, N65755, N65754, 
        N65753}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65771, N65770, 
        N65769, N65768, N65767, N65766}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__637, SYNOPSYS_UNCONNECTED__638, 
        SYNOPSYS_UNCONNECTED__639, SYNOPSYS_UNCONNECTED__640, 
        SYNOPSYS_UNCONNECTED__641, SYNOPSYS_UNCONNECTED__642, N67514, N67513, 
        N67512, N67511, N67510, N67509, N67508}) );
  hamming_N16000_CC2_DW01_add_135 add_2801_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65732, N65731, N65730, N65729, N65728, 
        N65727}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65745, N65744, 
        N65743, N65742, N65741, N65740}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__643, SYNOPSYS_UNCONNECTED__644, 
        SYNOPSYS_UNCONNECTED__645, SYNOPSYS_UNCONNECTED__646, 
        SYNOPSYS_UNCONNECTED__647, SYNOPSYS_UNCONNECTED__648, N67501, N67500, 
        N67499, N67498, N67497, N67496, N67495}) );
  hamming_N16000_CC2_DW01_add_136 add_2802_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65706, N65705, N65704, N65703, N65702, 
        N65701}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65719, N65718, 
        N65717, N65716, N65715, N65714}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__649, SYNOPSYS_UNCONNECTED__650, 
        SYNOPSYS_UNCONNECTED__651, SYNOPSYS_UNCONNECTED__652, 
        SYNOPSYS_UNCONNECTED__653, SYNOPSYS_UNCONNECTED__654, N67488, N67487, 
        N67486, N67485, N67484, N67483, N67482}) );
  hamming_N16000_CC2_DW01_add_137 add_2803_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65680, N65679, N65678, N65677, N65676, 
        N65675}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65693, N65692, 
        N65691, N65690, N65689, N65688}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__655, SYNOPSYS_UNCONNECTED__656, 
        SYNOPSYS_UNCONNECTED__657, SYNOPSYS_UNCONNECTED__658, 
        SYNOPSYS_UNCONNECTED__659, SYNOPSYS_UNCONNECTED__660, N67475, N67474, 
        N67473, N67472, N67471, N67470, N67469}) );
  hamming_N16000_CC2_DW01_add_138 add_2804_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65654, N65653, N65652, N65651, N65650, 
        N65649}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65667, N65666, 
        N65665, N65664, N65663, N65662}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__661, SYNOPSYS_UNCONNECTED__662, 
        SYNOPSYS_UNCONNECTED__663, SYNOPSYS_UNCONNECTED__664, 
        SYNOPSYS_UNCONNECTED__665, SYNOPSYS_UNCONNECTED__666, N67462, N67461, 
        N67460, N67459, N67458, N67457, N67456}) );
  hamming_N16000_CC2_DW01_add_139 add_2805_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65628, N65627, N65626, N65625, N65624, 
        N65623}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65641, N65640, 
        N65639, N65638, N65637, N65636}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__667, SYNOPSYS_UNCONNECTED__668, 
        SYNOPSYS_UNCONNECTED__669, SYNOPSYS_UNCONNECTED__670, 
        SYNOPSYS_UNCONNECTED__671, SYNOPSYS_UNCONNECTED__672, N67449, N67448, 
        N67447, N67446, N67445, N67444, N67443}) );
  hamming_N16000_CC2_DW01_add_140 add_2806_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65602, N65601, N65600, N65599, N65598, 
        N65597}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65615, N65614, 
        N65613, N65612, N65611, N65610}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__673, SYNOPSYS_UNCONNECTED__674, 
        SYNOPSYS_UNCONNECTED__675, SYNOPSYS_UNCONNECTED__676, 
        SYNOPSYS_UNCONNECTED__677, SYNOPSYS_UNCONNECTED__678, N67436, N67435, 
        N67434, N67433, N67432, N67431, N67430}) );
  hamming_N16000_CC2_DW01_add_141 add_2807_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65576, N65575, N65574, N65573, N65572, 
        N65571}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65589, N65588, 
        N65587, N65586, N65585, N65584}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__679, SYNOPSYS_UNCONNECTED__680, 
        SYNOPSYS_UNCONNECTED__681, SYNOPSYS_UNCONNECTED__682, 
        SYNOPSYS_UNCONNECTED__683, SYNOPSYS_UNCONNECTED__684, N67423, N67422, 
        N67421, N67420, N67419, N67418, N67417}) );
  hamming_N16000_CC2_DW01_add_142 add_2808_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65550, N65549, N65548, N65547, N65546, 
        N65545}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65563, N65562, 
        N65561, N65560, N65559, N65558}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__685, SYNOPSYS_UNCONNECTED__686, 
        SYNOPSYS_UNCONNECTED__687, SYNOPSYS_UNCONNECTED__688, 
        SYNOPSYS_UNCONNECTED__689, SYNOPSYS_UNCONNECTED__690, N67410, N67409, 
        N67408, N67407, N67406, N67405, N67404}) );
  hamming_N16000_CC2_DW01_add_143 add_2809_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65524, N65523, N65522, N65521, N65520, 
        N65519}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65537, N65536, 
        N65535, N65534, N65533, N65532}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__691, SYNOPSYS_UNCONNECTED__692, 
        SYNOPSYS_UNCONNECTED__693, SYNOPSYS_UNCONNECTED__694, 
        SYNOPSYS_UNCONNECTED__695, SYNOPSYS_UNCONNECTED__696, N67397, N67396, 
        N67395, N67394, N67393, N67392, N67391}) );
  hamming_N16000_CC2_DW01_add_144 add_2810_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65498, N65497, N65496, N65495, N65494, 
        N65493}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65511, N65510, 
        N65509, N65508, N65507, N65506}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__697, SYNOPSYS_UNCONNECTED__698, 
        SYNOPSYS_UNCONNECTED__699, SYNOPSYS_UNCONNECTED__700, 
        SYNOPSYS_UNCONNECTED__701, SYNOPSYS_UNCONNECTED__702, N67384, N67383, 
        N67382, N67381, N67380, N67379, N67378}) );
  hamming_N16000_CC2_DW01_add_145 add_2811_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65472, N65471, N65470, N65469, N65468, 
        N65467}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65485, N65484, 
        N65483, N65482, N65481, N65480}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__703, SYNOPSYS_UNCONNECTED__704, 
        SYNOPSYS_UNCONNECTED__705, SYNOPSYS_UNCONNECTED__706, 
        SYNOPSYS_UNCONNECTED__707, SYNOPSYS_UNCONNECTED__708, N67371, N67370, 
        N67369, N67368, N67367, N67366, N67365}) );
  hamming_N16000_CC2_DW01_add_146 add_2812_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65446, N65445, N65444, N65443, N65442, 
        N65441}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65459, N65458, 
        N65457, N65456, N65455, N65454}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__709, SYNOPSYS_UNCONNECTED__710, 
        SYNOPSYS_UNCONNECTED__711, SYNOPSYS_UNCONNECTED__712, 
        SYNOPSYS_UNCONNECTED__713, SYNOPSYS_UNCONNECTED__714, N67358, N67357, 
        N67356, N67355, N67354, N67353, N67352}) );
  hamming_N16000_CC2_DW01_add_147 add_2813_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65420, N65419, N65418, N65417, N65416, 
        N65415}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65433, N65432, 
        N65431, N65430, N65429, N65428}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__715, SYNOPSYS_UNCONNECTED__716, 
        SYNOPSYS_UNCONNECTED__717, SYNOPSYS_UNCONNECTED__718, 
        SYNOPSYS_UNCONNECTED__719, SYNOPSYS_UNCONNECTED__720, N67345, N67344, 
        N67343, N67342, N67341, N67340, N67339}) );
  hamming_N16000_CC2_DW01_add_148 add_2814_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65394, N65393, N65392, N65391, N65390, 
        N65389}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65407, N65406, 
        N65405, N65404, N65403, N65402}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__721, SYNOPSYS_UNCONNECTED__722, 
        SYNOPSYS_UNCONNECTED__723, SYNOPSYS_UNCONNECTED__724, 
        SYNOPSYS_UNCONNECTED__725, SYNOPSYS_UNCONNECTED__726, N67332, N67331, 
        N67330, N67329, N67328, N67327, N67326}) );
  hamming_N16000_CC2_DW01_add_149 add_2815_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65368, N65367, N65366, N65365, N65364, 
        N65363}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65381, N65380, 
        N65379, N65378, N65377, N65376}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__727, SYNOPSYS_UNCONNECTED__728, 
        SYNOPSYS_UNCONNECTED__729, SYNOPSYS_UNCONNECTED__730, 
        SYNOPSYS_UNCONNECTED__731, SYNOPSYS_UNCONNECTED__732, N67319, N67318, 
        N67317, N67316, N67315, N67314, N67313}) );
  hamming_N16000_CC2_DW01_add_150 add_2816_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65342, N65341, N65340, N65339, N65338, 
        N65337}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65355, N65354, 
        N65353, N65352, N65351, N65350}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__733, SYNOPSYS_UNCONNECTED__734, 
        SYNOPSYS_UNCONNECTED__735, SYNOPSYS_UNCONNECTED__736, 
        SYNOPSYS_UNCONNECTED__737, SYNOPSYS_UNCONNECTED__738, N67306, N67305, 
        N67304, N67303, N67302, N67301, N67300}) );
  hamming_N16000_CC2_DW01_add_151 add_2817_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65316, N65315, N65314, N65313, N65312, 
        N65311}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65329, N65328, 
        N65327, N65326, N65325, N65324}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__739, SYNOPSYS_UNCONNECTED__740, 
        SYNOPSYS_UNCONNECTED__741, SYNOPSYS_UNCONNECTED__742, 
        SYNOPSYS_UNCONNECTED__743, SYNOPSYS_UNCONNECTED__744, N67293, N67292, 
        N67291, N67290, N67289, N67288, N67287}) );
  hamming_N16000_CC2_DW01_add_152 add_2818_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65290, N65289, N65288, N65287, N65286, 
        N65285}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65303, N65302, 
        N65301, N65300, N65299, N65298}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__745, SYNOPSYS_UNCONNECTED__746, 
        SYNOPSYS_UNCONNECTED__747, SYNOPSYS_UNCONNECTED__748, 
        SYNOPSYS_UNCONNECTED__749, SYNOPSYS_UNCONNECTED__750, N67280, N67279, 
        N67278, N67277, N67276, N67275, N67274}) );
  hamming_N16000_CC2_DW01_add_153 add_2819_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65264, N65263, N65262, N65261, N65260, 
        N65259}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65277, N65276, 
        N65275, N65274, N65273, N65272}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__751, SYNOPSYS_UNCONNECTED__752, 
        SYNOPSYS_UNCONNECTED__753, SYNOPSYS_UNCONNECTED__754, 
        SYNOPSYS_UNCONNECTED__755, SYNOPSYS_UNCONNECTED__756, N67267, N67266, 
        N67265, N67264, N67263, N67262, N67261}) );
  hamming_N16000_CC2_DW01_add_154 add_2820_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65238, N65237, N65236, N65235, N65234, 
        N65233}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65251, N65250, 
        N65249, N65248, N65247, N65246}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__757, SYNOPSYS_UNCONNECTED__758, 
        SYNOPSYS_UNCONNECTED__759, SYNOPSYS_UNCONNECTED__760, 
        SYNOPSYS_UNCONNECTED__761, SYNOPSYS_UNCONNECTED__762, N67254, N67253, 
        N67252, N67251, N67250, N67249, N67248}) );
  hamming_N16000_CC2_DW01_add_155 add_2821_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65212, N65211, N65210, N65209, N65208, 
        N65207}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65225, N65224, 
        N65223, N65222, N65221, N65220}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__763, SYNOPSYS_UNCONNECTED__764, 
        SYNOPSYS_UNCONNECTED__765, SYNOPSYS_UNCONNECTED__766, 
        SYNOPSYS_UNCONNECTED__767, SYNOPSYS_UNCONNECTED__768, N67241, N67240, 
        N67239, N67238, N67237, N67236, N67235}) );
  hamming_N16000_CC2_DW01_add_156 add_2822_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65186, N65185, N65184, N65183, N65182, 
        N65181}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65199, N65198, 
        N65197, N65196, N65195, N65194}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__769, SYNOPSYS_UNCONNECTED__770, 
        SYNOPSYS_UNCONNECTED__771, SYNOPSYS_UNCONNECTED__772, 
        SYNOPSYS_UNCONNECTED__773, SYNOPSYS_UNCONNECTED__774, N67228, N67227, 
        N67226, N67225, N67224, N67223, N67222}) );
  hamming_N16000_CC2_DW01_add_157 add_2823_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65160, N65159, N65158, N65157, N65156, 
        N65155}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65173, N65172, 
        N65171, N65170, N65169, N65168}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__775, SYNOPSYS_UNCONNECTED__776, 
        SYNOPSYS_UNCONNECTED__777, SYNOPSYS_UNCONNECTED__778, 
        SYNOPSYS_UNCONNECTED__779, SYNOPSYS_UNCONNECTED__780, N67215, N67214, 
        N67213, N67212, N67211, N67210, N67209}) );
  hamming_N16000_CC2_DW01_add_158 add_2824_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65134, N65133, N65132, N65131, N65130, 
        N65129}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65147, N65146, 
        N65145, N65144, N65143, N65142}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__781, SYNOPSYS_UNCONNECTED__782, 
        SYNOPSYS_UNCONNECTED__783, SYNOPSYS_UNCONNECTED__784, 
        SYNOPSYS_UNCONNECTED__785, SYNOPSYS_UNCONNECTED__786, N67202, N67201, 
        N67200, N67199, N67198, N67197, N67196}) );
  hamming_N16000_CC2_DW01_add_159 add_2825_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65108, N65107, N65106, N65105, N65104, 
        N65103}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65121, N65120, 
        N65119, N65118, N65117, N65116}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__787, SYNOPSYS_UNCONNECTED__788, 
        SYNOPSYS_UNCONNECTED__789, SYNOPSYS_UNCONNECTED__790, 
        SYNOPSYS_UNCONNECTED__791, SYNOPSYS_UNCONNECTED__792, N67189, N67188, 
        N67187, N67186, N67185, N67184, N67183}) );
  hamming_N16000_CC2_DW01_add_160 add_2826_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65082, N65081, N65080, N65079, N65078, 
        N65077}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65095, N65094, 
        N65093, N65092, N65091, N65090}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__793, SYNOPSYS_UNCONNECTED__794, 
        SYNOPSYS_UNCONNECTED__795, SYNOPSYS_UNCONNECTED__796, 
        SYNOPSYS_UNCONNECTED__797, SYNOPSYS_UNCONNECTED__798, N67176, N67175, 
        N67174, N67173, N67172, N67171, N67170}) );
  hamming_N16000_CC2_DW01_add_161 add_2827_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65056, N65055, N65054, N65053, N65052, 
        N65051}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65069, N65068, 
        N65067, N65066, N65065, N65064}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__799, SYNOPSYS_UNCONNECTED__800, 
        SYNOPSYS_UNCONNECTED__801, SYNOPSYS_UNCONNECTED__802, 
        SYNOPSYS_UNCONNECTED__803, SYNOPSYS_UNCONNECTED__804, N67163, N67162, 
        N67161, N67160, N67159, N67158, N67157}) );
  hamming_N16000_CC2_DW01_add_162 add_2828_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65030, N65029, N65028, N65027, N65026, 
        N65025}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65043, N65042, 
        N65041, N65040, N65039, N65038}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__805, SYNOPSYS_UNCONNECTED__806, 
        SYNOPSYS_UNCONNECTED__807, SYNOPSYS_UNCONNECTED__808, 
        SYNOPSYS_UNCONNECTED__809, SYNOPSYS_UNCONNECTED__810, N67150, N67149, 
        N67148, N67147, N67146, N67145, N67144}) );
  hamming_N16000_CC2_DW01_add_163 add_2829_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65004, N65003, N65002, N65001, N65000, 
        N64999}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65017, N65016, 
        N65015, N65014, N65013, N65012}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__811, SYNOPSYS_UNCONNECTED__812, 
        SYNOPSYS_UNCONNECTED__813, SYNOPSYS_UNCONNECTED__814, 
        SYNOPSYS_UNCONNECTED__815, SYNOPSYS_UNCONNECTED__816, N67137, N67136, 
        N67135, N67134, N67133, N67132, N67131}) );
  hamming_N16000_CC2_DW01_add_164 add_2830_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64978, N64977, N64976, N64975, N64974, 
        N64973}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64991, N64990, 
        N64989, N64988, N64987, N64986}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__817, SYNOPSYS_UNCONNECTED__818, 
        SYNOPSYS_UNCONNECTED__819, SYNOPSYS_UNCONNECTED__820, 
        SYNOPSYS_UNCONNECTED__821, SYNOPSYS_UNCONNECTED__822, N67124, N67123, 
        N67122, N67121, N67120, N67119, N67118}) );
  hamming_N16000_CC2_DW01_add_165 add_2831_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64952, N64951, N64950, N64949, N64948, 
        N64947}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64965, N64964, 
        N64963, N64962, N64961, N64960}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__823, SYNOPSYS_UNCONNECTED__824, 
        SYNOPSYS_UNCONNECTED__825, SYNOPSYS_UNCONNECTED__826, 
        SYNOPSYS_UNCONNECTED__827, SYNOPSYS_UNCONNECTED__828, N67111, N67110, 
        N67109, N67108, N67107, N67106, N67105}) );
  hamming_N16000_CC2_DW01_add_166 add_2832_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64926, N64925, N64924, N64923, N64922, 
        N64921}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64939, N64938, 
        N64937, N64936, N64935, N64934}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__829, SYNOPSYS_UNCONNECTED__830, 
        SYNOPSYS_UNCONNECTED__831, SYNOPSYS_UNCONNECTED__832, 
        SYNOPSYS_UNCONNECTED__833, SYNOPSYS_UNCONNECTED__834, N67098, N67097, 
        N67096, N67095, N67094, N67093, N67092}) );
  hamming_N16000_CC2_DW01_add_167 add_2833_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64899, N64898, N64897, N64896, 
        N64895}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64912, 
        N64911, N64910, N64909, N64908}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__835, SYNOPSYS_UNCONNECTED__836, 
        SYNOPSYS_UNCONNECTED__837, SYNOPSYS_UNCONNECTED__838, 
        SYNOPSYS_UNCONNECTED__839, SYNOPSYS_UNCONNECTED__840, 
        SYNOPSYS_UNCONNECTED__841, N67084, N67083, N67082, N67081, N67080, 
        N67079}) );
  hamming_N16000_CC2_DW01_add_168 add_2834_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64873, N64872, N64871, N64870, 
        N64869}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64886, 
        N64885, N64884, N64883, N64882}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__842, SYNOPSYS_UNCONNECTED__843, 
        SYNOPSYS_UNCONNECTED__844, SYNOPSYS_UNCONNECTED__845, 
        SYNOPSYS_UNCONNECTED__846, SYNOPSYS_UNCONNECTED__847, 
        SYNOPSYS_UNCONNECTED__848, N67071, N67070, N67069, N67068, N67067, 
        N67066}) );
  hamming_N16000_CC2_DW01_add_169 add_2835_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64847, N64846, N64845, N64844, 
        N64843}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64860, 
        N64859, N64858, N64857, N64856}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__849, SYNOPSYS_UNCONNECTED__850, 
        SYNOPSYS_UNCONNECTED__851, SYNOPSYS_UNCONNECTED__852, 
        SYNOPSYS_UNCONNECTED__853, SYNOPSYS_UNCONNECTED__854, 
        SYNOPSYS_UNCONNECTED__855, N67058, N67057, N67056, N67055, N67054, 
        N67053}) );
  hamming_N16000_CC2_DW01_add_170 add_2836_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64821, N64820, N64819, N64818, 
        N64817}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64834, 
        N64833, N64832, N64831, N64830}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__856, SYNOPSYS_UNCONNECTED__857, 
        SYNOPSYS_UNCONNECTED__858, SYNOPSYS_UNCONNECTED__859, 
        SYNOPSYS_UNCONNECTED__860, SYNOPSYS_UNCONNECTED__861, 
        SYNOPSYS_UNCONNECTED__862, N67045, N67044, N67043, N67042, N67041, 
        N67040}) );
  hamming_N16000_CC2_DW01_add_171 add_2837_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64795, N64794, N64793, N64792, 
        N64791}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64808, 
        N64807, N64806, N64805, N64804}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__863, SYNOPSYS_UNCONNECTED__864, 
        SYNOPSYS_UNCONNECTED__865, SYNOPSYS_UNCONNECTED__866, 
        SYNOPSYS_UNCONNECTED__867, SYNOPSYS_UNCONNECTED__868, 
        SYNOPSYS_UNCONNECTED__869, N67032, N67031, N67030, N67029, N67028, 
        N67027}) );
  hamming_N16000_CC2_DW01_add_172 add_2838_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64769, N64768, N64767, N64766, 
        N64765}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64782, 
        N64781, N64780, N64779, N64778}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__870, SYNOPSYS_UNCONNECTED__871, 
        SYNOPSYS_UNCONNECTED__872, SYNOPSYS_UNCONNECTED__873, 
        SYNOPSYS_UNCONNECTED__874, SYNOPSYS_UNCONNECTED__875, 
        SYNOPSYS_UNCONNECTED__876, N67019, N67018, N67017, N67016, N67015, 
        N67014}) );
  hamming_N16000_CC2_DW01_add_173 add_2839_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64743, N64742, N64741, N64740, 
        N64739}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64756, 
        N64755, N64754, N64753, N64752}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__877, SYNOPSYS_UNCONNECTED__878, 
        SYNOPSYS_UNCONNECTED__879, SYNOPSYS_UNCONNECTED__880, 
        SYNOPSYS_UNCONNECTED__881, SYNOPSYS_UNCONNECTED__882, 
        SYNOPSYS_UNCONNECTED__883, N67006, N67005, N67004, N67003, N67002, 
        N67001}) );
  hamming_N16000_CC2_DW01_add_174 add_2840_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64717, N64716, N64715, N64714, 
        N64713}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64730, 
        N64729, N64728, N64727, N64726}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__884, SYNOPSYS_UNCONNECTED__885, 
        SYNOPSYS_UNCONNECTED__886, SYNOPSYS_UNCONNECTED__887, 
        SYNOPSYS_UNCONNECTED__888, SYNOPSYS_UNCONNECTED__889, 
        SYNOPSYS_UNCONNECTED__890, N66993, N66992, N66991, N66990, N66989, 
        N66988}) );
  hamming_N16000_CC2_DW01_add_175 add_2841_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64691, N64690, N64689, N64688, 
        N64687}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64704, 
        N64703, N64702, N64701, N64700}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__891, SYNOPSYS_UNCONNECTED__892, 
        SYNOPSYS_UNCONNECTED__893, SYNOPSYS_UNCONNECTED__894, 
        SYNOPSYS_UNCONNECTED__895, SYNOPSYS_UNCONNECTED__896, 
        SYNOPSYS_UNCONNECTED__897, N66980, N66979, N66978, N66977, N66976, 
        N66975}) );
  hamming_N16000_CC2_DW01_add_176 add_2842_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64665, N64664, N64663, N64662, 
        N64661}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64678, 
        N64677, N64676, N64675, N64674}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__898, SYNOPSYS_UNCONNECTED__899, 
        SYNOPSYS_UNCONNECTED__900, SYNOPSYS_UNCONNECTED__901, 
        SYNOPSYS_UNCONNECTED__902, SYNOPSYS_UNCONNECTED__903, 
        SYNOPSYS_UNCONNECTED__904, N66967, N66966, N66965, N66964, N66963, 
        N66962}) );
  hamming_N16000_CC2_DW01_add_177 add_2843_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64639, N64638, N64637, N64636, 
        N64635}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64652, 
        N64651, N64650, N64649, N64648}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__905, SYNOPSYS_UNCONNECTED__906, 
        SYNOPSYS_UNCONNECTED__907, SYNOPSYS_UNCONNECTED__908, 
        SYNOPSYS_UNCONNECTED__909, SYNOPSYS_UNCONNECTED__910, 
        SYNOPSYS_UNCONNECTED__911, N66954, N66953, N66952, N66951, N66950, 
        N66949}) );
  hamming_N16000_CC2_DW01_add_178 add_2844_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64613, N64612, N64611, N64610, 
        N64609}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64626, 
        N64625, N64624, N64623, N64622}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__912, SYNOPSYS_UNCONNECTED__913, 
        SYNOPSYS_UNCONNECTED__914, SYNOPSYS_UNCONNECTED__915, 
        SYNOPSYS_UNCONNECTED__916, SYNOPSYS_UNCONNECTED__917, 
        SYNOPSYS_UNCONNECTED__918, N66941, N66940, N66939, N66938, N66937, 
        N66936}) );
  hamming_N16000_CC2_DW01_add_179 add_2845_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64587, N64586, N64585, N64584, 
        N64583}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64600, 
        N64599, N64598, N64597, N64596}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__919, SYNOPSYS_UNCONNECTED__920, 
        SYNOPSYS_UNCONNECTED__921, SYNOPSYS_UNCONNECTED__922, 
        SYNOPSYS_UNCONNECTED__923, SYNOPSYS_UNCONNECTED__924, 
        SYNOPSYS_UNCONNECTED__925, N66928, N66927, N66926, N66925, N66924, 
        N66923}) );
  hamming_N16000_CC2_DW01_add_180 add_2846_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64561, N64560, N64559, N64558, 
        N64557}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64574, 
        N64573, N64572, N64571, N64570}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__926, SYNOPSYS_UNCONNECTED__927, 
        SYNOPSYS_UNCONNECTED__928, SYNOPSYS_UNCONNECTED__929, 
        SYNOPSYS_UNCONNECTED__930, SYNOPSYS_UNCONNECTED__931, 
        SYNOPSYS_UNCONNECTED__932, N66915, N66914, N66913, N66912, N66911, 
        N66910}) );
  hamming_N16000_CC2_DW01_add_181 add_2847_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64535, N64534, N64533, N64532, 
        N64531}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64548, 
        N64547, N64546, N64545, N64544}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__933, SYNOPSYS_UNCONNECTED__934, 
        SYNOPSYS_UNCONNECTED__935, SYNOPSYS_UNCONNECTED__936, 
        SYNOPSYS_UNCONNECTED__937, SYNOPSYS_UNCONNECTED__938, 
        SYNOPSYS_UNCONNECTED__939, N66902, N66901, N66900, N66899, N66898, 
        N66897}) );
  hamming_N16000_CC2_DW01_add_182 add_2848_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64509, N64508, N64507, N64506, 
        N64505}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64522, 
        N64521, N64520, N64519, N64518}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__940, SYNOPSYS_UNCONNECTED__941, 
        SYNOPSYS_UNCONNECTED__942, SYNOPSYS_UNCONNECTED__943, 
        SYNOPSYS_UNCONNECTED__944, SYNOPSYS_UNCONNECTED__945, 
        SYNOPSYS_UNCONNECTED__946, N66889, N66888, N66887, N66886, N66885, 
        N66884}) );
  hamming_N16000_CC2_DW01_add_183 add_2849_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64483, N64482, N64481, N64480, 
        N64479}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64496, 
        N64495, N64494, N64493, N64492}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__947, SYNOPSYS_UNCONNECTED__948, 
        SYNOPSYS_UNCONNECTED__949, SYNOPSYS_UNCONNECTED__950, 
        SYNOPSYS_UNCONNECTED__951, SYNOPSYS_UNCONNECTED__952, 
        SYNOPSYS_UNCONNECTED__953, N66876, N66875, N66874, N66873, N66872, 
        N66871}) );
  hamming_N16000_CC2_DW01_add_184 add_2850_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64457, N64456, N64455, N64454, 
        N64453}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64470, 
        N64469, N64468, N64467, N64466}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__954, SYNOPSYS_UNCONNECTED__955, 
        SYNOPSYS_UNCONNECTED__956, SYNOPSYS_UNCONNECTED__957, 
        SYNOPSYS_UNCONNECTED__958, SYNOPSYS_UNCONNECTED__959, 
        SYNOPSYS_UNCONNECTED__960, N66863, N66862, N66861, N66860, N66859, 
        N66858}) );
  hamming_N16000_CC2_DW01_add_185 add_2851_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64431, N64430, N64429, N64428, 
        N64427}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64444, 
        N64443, N64442, N64441, N64440}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__961, SYNOPSYS_UNCONNECTED__962, 
        SYNOPSYS_UNCONNECTED__963, SYNOPSYS_UNCONNECTED__964, 
        SYNOPSYS_UNCONNECTED__965, SYNOPSYS_UNCONNECTED__966, 
        SYNOPSYS_UNCONNECTED__967, N66850, N66849, N66848, N66847, N66846, 
        N66845}) );
  hamming_N16000_CC2_DW01_add_186 add_2852_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64405, N64404, N64403, N64402, 
        N64401}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64418, 
        N64417, N64416, N64415, N64414}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__968, SYNOPSYS_UNCONNECTED__969, 
        SYNOPSYS_UNCONNECTED__970, SYNOPSYS_UNCONNECTED__971, 
        SYNOPSYS_UNCONNECTED__972, SYNOPSYS_UNCONNECTED__973, 
        SYNOPSYS_UNCONNECTED__974, N66837, N66836, N66835, N66834, N66833, 
        N66832}) );
  hamming_N16000_CC2_DW01_add_187 add_2853_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64379, N64378, N64377, N64376, 
        N64375}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64392, 
        N64391, N64390, N64389, N64388}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__975, SYNOPSYS_UNCONNECTED__976, 
        SYNOPSYS_UNCONNECTED__977, SYNOPSYS_UNCONNECTED__978, 
        SYNOPSYS_UNCONNECTED__979, SYNOPSYS_UNCONNECTED__980, 
        SYNOPSYS_UNCONNECTED__981, N66824, N66823, N66822, N66821, N66820, 
        N66819}) );
  hamming_N16000_CC2_DW01_add_188 add_2854_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64353, N64352, N64351, N64350, 
        N64349}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64366, 
        N64365, N64364, N64363, N64362}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__982, SYNOPSYS_UNCONNECTED__983, 
        SYNOPSYS_UNCONNECTED__984, SYNOPSYS_UNCONNECTED__985, 
        SYNOPSYS_UNCONNECTED__986, SYNOPSYS_UNCONNECTED__987, 
        SYNOPSYS_UNCONNECTED__988, N66811, N66810, N66809, N66808, N66807, 
        N66806}) );
  hamming_N16000_CC2_DW01_add_189 add_2855_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64327, N64326, N64325, N64324, 
        N64323}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64340, 
        N64339, N64338, N64337, N64336}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__989, SYNOPSYS_UNCONNECTED__990, 
        SYNOPSYS_UNCONNECTED__991, SYNOPSYS_UNCONNECTED__992, 
        SYNOPSYS_UNCONNECTED__993, SYNOPSYS_UNCONNECTED__994, 
        SYNOPSYS_UNCONNECTED__995, N66798, N66797, N66796, N66795, N66794, 
        N66793}) );
  hamming_N16000_CC2_DW01_add_190 add_2856_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64301, N64300, N64299, N64298, 
        N64297}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64314, 
        N64313, N64312, N64311, N64310}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__996, SYNOPSYS_UNCONNECTED__997, 
        SYNOPSYS_UNCONNECTED__998, SYNOPSYS_UNCONNECTED__999, 
        SYNOPSYS_UNCONNECTED__1000, SYNOPSYS_UNCONNECTED__1001, 
        SYNOPSYS_UNCONNECTED__1002, N66785, N66784, N66783, N66782, N66781, 
        N66780}) );
  hamming_N16000_CC2_DW01_add_191 add_2857_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64275, N64274, N64273, N64272, 
        N64271}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64288, 
        N64287, N64286, N64285, N64284}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1003, SYNOPSYS_UNCONNECTED__1004, 
        SYNOPSYS_UNCONNECTED__1005, SYNOPSYS_UNCONNECTED__1006, 
        SYNOPSYS_UNCONNECTED__1007, SYNOPSYS_UNCONNECTED__1008, 
        SYNOPSYS_UNCONNECTED__1009, N66772, N66771, N66770, N66769, N66768, 
        N66767}) );
  hamming_N16000_CC2_DW01_add_192 add_2858_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64249, N64248, N64247, N64246, 
        N64245}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64262, 
        N64261, N64260, N64259, N64258}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1010, SYNOPSYS_UNCONNECTED__1011, 
        SYNOPSYS_UNCONNECTED__1012, SYNOPSYS_UNCONNECTED__1013, 
        SYNOPSYS_UNCONNECTED__1014, SYNOPSYS_UNCONNECTED__1015, 
        SYNOPSYS_UNCONNECTED__1016, N66759, N66758, N66757, N66756, N66755, 
        N66754}) );
  hamming_N16000_CC2_DW01_add_193 add_2859_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64223, N64222, N64221, N64220, 
        N64219}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64236, 
        N64235, N64234, N64233, N64232}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1017, SYNOPSYS_UNCONNECTED__1018, 
        SYNOPSYS_UNCONNECTED__1019, SYNOPSYS_UNCONNECTED__1020, 
        SYNOPSYS_UNCONNECTED__1021, SYNOPSYS_UNCONNECTED__1022, 
        SYNOPSYS_UNCONNECTED__1023, N66746, N66745, N66744, N66743, N66742, 
        N66741}) );
  hamming_N16000_CC2_DW01_add_194 add_2860_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64197, N64196, N64195, N64194, 
        N64193}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64210, 
        N64209, N64208, N64207, N64206}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1024, SYNOPSYS_UNCONNECTED__1025, 
        SYNOPSYS_UNCONNECTED__1026, SYNOPSYS_UNCONNECTED__1027, 
        SYNOPSYS_UNCONNECTED__1028, SYNOPSYS_UNCONNECTED__1029, 
        SYNOPSYS_UNCONNECTED__1030, N66733, N66732, N66731, N66730, N66729, 
        N66728}) );
  hamming_N16000_CC2_DW01_add_195 add_2861_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64171, N64170, N64169, N64168, 
        N64167}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64184, 
        N64183, N64182, N64181, N64180}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1031, SYNOPSYS_UNCONNECTED__1032, 
        SYNOPSYS_UNCONNECTED__1033, SYNOPSYS_UNCONNECTED__1034, 
        SYNOPSYS_UNCONNECTED__1035, SYNOPSYS_UNCONNECTED__1036, 
        SYNOPSYS_UNCONNECTED__1037, N66720, N66719, N66718, N66717, N66716, 
        N66715}) );
  hamming_N16000_CC2_DW01_add_196 add_2862_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64145, N64144, N64143, N64142, 
        N64141}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64158, 
        N64157, N64156, N64155, N64154}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1038, SYNOPSYS_UNCONNECTED__1039, 
        SYNOPSYS_UNCONNECTED__1040, SYNOPSYS_UNCONNECTED__1041, 
        SYNOPSYS_UNCONNECTED__1042, SYNOPSYS_UNCONNECTED__1043, 
        SYNOPSYS_UNCONNECTED__1044, N66707, N66706, N66705, N66704, N66703, 
        N66702}) );
  hamming_N16000_CC2_DW01_add_197 add_2863_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64119, N64118, N64117, N64116, 
        N64115}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64132, 
        N64131, N64130, N64129, N64128}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1045, SYNOPSYS_UNCONNECTED__1046, 
        SYNOPSYS_UNCONNECTED__1047, SYNOPSYS_UNCONNECTED__1048, 
        SYNOPSYS_UNCONNECTED__1049, SYNOPSYS_UNCONNECTED__1050, 
        SYNOPSYS_UNCONNECTED__1051, N66694, N66693, N66692, N66691, N66690, 
        N66689}) );
  hamming_N16000_CC2_DW01_add_198 add_2864_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64093, N64092, N64091, N64090, 
        N64089}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64106, 
        N64105, N64104, N64103, N64102}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1052, SYNOPSYS_UNCONNECTED__1053, 
        SYNOPSYS_UNCONNECTED__1054, SYNOPSYS_UNCONNECTED__1055, 
        SYNOPSYS_UNCONNECTED__1056, SYNOPSYS_UNCONNECTED__1057, 
        SYNOPSYS_UNCONNECTED__1058, N66681, N66680, N66679, N66678, N66677, 
        N66676}) );
  hamming_N16000_CC2_DW01_add_199 add_2865_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64067, N64066, N64065, N64064, 
        N64063}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64080, 
        N64079, N64078, N64077, N64076}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1059, SYNOPSYS_UNCONNECTED__1060, 
        SYNOPSYS_UNCONNECTED__1061, SYNOPSYS_UNCONNECTED__1062, 
        SYNOPSYS_UNCONNECTED__1063, SYNOPSYS_UNCONNECTED__1064, 
        SYNOPSYS_UNCONNECTED__1065, N66668, N66667, N66666, N66665, N66664, 
        N66663}) );
  hamming_N16000_CC2_DW01_add_200 add_2866_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64041, N64040, N64039, N64038, 
        N64037}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64054, 
        N64053, N64052, N64051, N64050}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1066, SYNOPSYS_UNCONNECTED__1067, 
        SYNOPSYS_UNCONNECTED__1068, SYNOPSYS_UNCONNECTED__1069, 
        SYNOPSYS_UNCONNECTED__1070, SYNOPSYS_UNCONNECTED__1071, 
        SYNOPSYS_UNCONNECTED__1072, N66655, N66654, N66653, N66652, N66651, 
        N66650}) );
  hamming_N16000_CC2_DW01_add_201 add_2867_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64015, N64014, N64013, N64012, 
        N64011}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64028, 
        N64027, N64026, N64025, N64024}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1073, SYNOPSYS_UNCONNECTED__1074, 
        SYNOPSYS_UNCONNECTED__1075, SYNOPSYS_UNCONNECTED__1076, 
        SYNOPSYS_UNCONNECTED__1077, SYNOPSYS_UNCONNECTED__1078, 
        SYNOPSYS_UNCONNECTED__1079, N66642, N66641, N66640, N66639, N66638, 
        N66637}) );
  hamming_N16000_CC2_DW01_add_202 add_2868_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63989, N63988, N63987, N63986, 
        N63985}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64002, 
        N64001, N64000, N63999, N63998}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1080, SYNOPSYS_UNCONNECTED__1081, 
        SYNOPSYS_UNCONNECTED__1082, SYNOPSYS_UNCONNECTED__1083, 
        SYNOPSYS_UNCONNECTED__1084, SYNOPSYS_UNCONNECTED__1085, 
        SYNOPSYS_UNCONNECTED__1086, N66629, N66628, N66627, N66626, N66625, 
        N66624}) );
  hamming_N16000_CC2_DW01_add_203 add_2869_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63963, N63962, N63961, N63960, 
        N63959}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63976, 
        N63975, N63974, N63973, N63972}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1087, SYNOPSYS_UNCONNECTED__1088, 
        SYNOPSYS_UNCONNECTED__1089, SYNOPSYS_UNCONNECTED__1090, 
        SYNOPSYS_UNCONNECTED__1091, SYNOPSYS_UNCONNECTED__1092, 
        SYNOPSYS_UNCONNECTED__1093, N66616, N66615, N66614, N66613, N66612, 
        N66611}) );
  hamming_N16000_CC2_DW01_add_204 add_2870_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63937, N63936, N63935, N63934, 
        N63933}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63950, 
        N63949, N63948, N63947, N63946}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1094, SYNOPSYS_UNCONNECTED__1095, 
        SYNOPSYS_UNCONNECTED__1096, SYNOPSYS_UNCONNECTED__1097, 
        SYNOPSYS_UNCONNECTED__1098, SYNOPSYS_UNCONNECTED__1099, 
        SYNOPSYS_UNCONNECTED__1100, N66603, N66602, N66601, N66600, N66599, 
        N66598}) );
  hamming_N16000_CC2_DW01_add_205 add_2871_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63911, N63910, N63909, N63908, 
        N63907}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63924, 
        N63923, N63922, N63921, N63920}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1101, SYNOPSYS_UNCONNECTED__1102, 
        SYNOPSYS_UNCONNECTED__1103, SYNOPSYS_UNCONNECTED__1104, 
        SYNOPSYS_UNCONNECTED__1105, SYNOPSYS_UNCONNECTED__1106, 
        SYNOPSYS_UNCONNECTED__1107, N66590, N66589, N66588, N66587, N66586, 
        N66585}) );
  hamming_N16000_CC2_DW01_add_206 add_2872_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63885, N63884, N63883, N63882, 
        N63881}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63898, 
        N63897, N63896, N63895, N63894}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1108, SYNOPSYS_UNCONNECTED__1109, 
        SYNOPSYS_UNCONNECTED__1110, SYNOPSYS_UNCONNECTED__1111, 
        SYNOPSYS_UNCONNECTED__1112, SYNOPSYS_UNCONNECTED__1113, 
        SYNOPSYS_UNCONNECTED__1114, N66577, N66576, N66575, N66574, N66573, 
        N66572}) );
  hamming_N16000_CC2_DW01_add_207 add_2873_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63859, N63858, N63857, N63856, 
        N63855}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63872, 
        N63871, N63870, N63869, N63868}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1115, SYNOPSYS_UNCONNECTED__1116, 
        SYNOPSYS_UNCONNECTED__1117, SYNOPSYS_UNCONNECTED__1118, 
        SYNOPSYS_UNCONNECTED__1119, SYNOPSYS_UNCONNECTED__1120, 
        SYNOPSYS_UNCONNECTED__1121, N66564, N66563, N66562, N66561, N66560, 
        N66559}) );
  hamming_N16000_CC2_DW01_add_208 add_2874_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63833, N63832, N63831, N63830, 
        N63829}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63846, 
        N63845, N63844, N63843, N63842}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1122, SYNOPSYS_UNCONNECTED__1123, 
        SYNOPSYS_UNCONNECTED__1124, SYNOPSYS_UNCONNECTED__1125, 
        SYNOPSYS_UNCONNECTED__1126, SYNOPSYS_UNCONNECTED__1127, 
        SYNOPSYS_UNCONNECTED__1128, N66551, N66550, N66549, N66548, N66547, 
        N66546}) );
  hamming_N16000_CC2_DW01_add_209 add_2875_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63807, N63806, N63805, N63804, 
        N63803}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63820, 
        N63819, N63818, N63817, N63816}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1129, SYNOPSYS_UNCONNECTED__1130, 
        SYNOPSYS_UNCONNECTED__1131, SYNOPSYS_UNCONNECTED__1132, 
        SYNOPSYS_UNCONNECTED__1133, SYNOPSYS_UNCONNECTED__1134, 
        SYNOPSYS_UNCONNECTED__1135, N66538, N66537, N66536, N66535, N66534, 
        N66533}) );
  hamming_N16000_CC2_DW01_add_210 add_2876_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63781, N63780, N63779, N63778, 
        N63777}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63794, 
        N63793, N63792, N63791, N63790}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1136, SYNOPSYS_UNCONNECTED__1137, 
        SYNOPSYS_UNCONNECTED__1138, SYNOPSYS_UNCONNECTED__1139, 
        SYNOPSYS_UNCONNECTED__1140, SYNOPSYS_UNCONNECTED__1141, 
        SYNOPSYS_UNCONNECTED__1142, N66525, N66524, N66523, N66522, N66521, 
        N66520}) );
  hamming_N16000_CC2_DW01_add_211 add_2877_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63755, N63754, N63753, N63752, 
        N63751}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63768, 
        N63767, N63766, N63765, N63764}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1143, SYNOPSYS_UNCONNECTED__1144, 
        SYNOPSYS_UNCONNECTED__1145, SYNOPSYS_UNCONNECTED__1146, 
        SYNOPSYS_UNCONNECTED__1147, SYNOPSYS_UNCONNECTED__1148, 
        SYNOPSYS_UNCONNECTED__1149, N66512, N66511, N66510, N66509, N66508, 
        N66507}) );
  hamming_N16000_CC2_DW01_add_212 add_2878_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63729, N63728, N63727, N63726, 
        N63725}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63742, 
        N63741, N63740, N63739, N63738}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1150, SYNOPSYS_UNCONNECTED__1151, 
        SYNOPSYS_UNCONNECTED__1152, SYNOPSYS_UNCONNECTED__1153, 
        SYNOPSYS_UNCONNECTED__1154, SYNOPSYS_UNCONNECTED__1155, 
        SYNOPSYS_UNCONNECTED__1156, N66499, N66498, N66497, N66496, N66495, 
        N66494}) );
  hamming_N16000_CC2_DW01_add_213 add_2879_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63703, N63702, N63701, N63700, 
        N63699}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63716, 
        N63715, N63714, N63713, N63712}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1157, SYNOPSYS_UNCONNECTED__1158, 
        SYNOPSYS_UNCONNECTED__1159, SYNOPSYS_UNCONNECTED__1160, 
        SYNOPSYS_UNCONNECTED__1161, SYNOPSYS_UNCONNECTED__1162, 
        SYNOPSYS_UNCONNECTED__1163, N66486, N66485, N66484, N66483, N66482, 
        N66481}) );
  hamming_N16000_CC2_DW01_add_214 add_2880_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63677, N63676, N63675, N63674, 
        N63673}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63690, 
        N63689, N63688, N63687, N63686}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1164, SYNOPSYS_UNCONNECTED__1165, 
        SYNOPSYS_UNCONNECTED__1166, SYNOPSYS_UNCONNECTED__1167, 
        SYNOPSYS_UNCONNECTED__1168, SYNOPSYS_UNCONNECTED__1169, 
        SYNOPSYS_UNCONNECTED__1170, N66473, N66472, N66471, N66470, N66469, 
        N66468}) );
  hamming_N16000_CC2_DW01_add_215 add_2881_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63651, N63650, N63649, N63648, 
        N63647}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63664, 
        N63663, N63662, N63661, N63660}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1171, SYNOPSYS_UNCONNECTED__1172, 
        SYNOPSYS_UNCONNECTED__1173, SYNOPSYS_UNCONNECTED__1174, 
        SYNOPSYS_UNCONNECTED__1175, SYNOPSYS_UNCONNECTED__1176, 
        SYNOPSYS_UNCONNECTED__1177, N66460, N66459, N66458, N66457, N66456, 
        N66455}) );
  hamming_N16000_CC2_DW01_add_216 add_2882_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63625, N63624, N63623, N63622, 
        N63621}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63638, 
        N63637, N63636, N63635, N63634}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1178, SYNOPSYS_UNCONNECTED__1179, 
        SYNOPSYS_UNCONNECTED__1180, SYNOPSYS_UNCONNECTED__1181, 
        SYNOPSYS_UNCONNECTED__1182, SYNOPSYS_UNCONNECTED__1183, 
        SYNOPSYS_UNCONNECTED__1184, N66447, N66446, N66445, N66444, N66443, 
        N66442}) );
  hamming_N16000_CC2_DW01_add_217 add_2883_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63599, N63598, N63597, N63596, 
        N63595}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63612, 
        N63611, N63610, N63609, N63608}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1185, SYNOPSYS_UNCONNECTED__1186, 
        SYNOPSYS_UNCONNECTED__1187, SYNOPSYS_UNCONNECTED__1188, 
        SYNOPSYS_UNCONNECTED__1189, SYNOPSYS_UNCONNECTED__1190, 
        SYNOPSYS_UNCONNECTED__1191, N66434, N66433, N66432, N66431, N66430, 
        N66429}) );
  hamming_N16000_CC2_DW01_add_218 add_2884_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63573, N63572, N63571, N63570, 
        N63569}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63586, 
        N63585, N63584, N63583, N63582}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1192, SYNOPSYS_UNCONNECTED__1193, 
        SYNOPSYS_UNCONNECTED__1194, SYNOPSYS_UNCONNECTED__1195, 
        SYNOPSYS_UNCONNECTED__1196, SYNOPSYS_UNCONNECTED__1197, 
        SYNOPSYS_UNCONNECTED__1198, N66421, N66420, N66419, N66418, N66417, 
        N66416}) );
  hamming_N16000_CC2_DW01_add_219 add_2885_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63547, N63546, N63545, N63544, 
        N63543}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63560, 
        N63559, N63558, N63557, N63556}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1199, SYNOPSYS_UNCONNECTED__1200, 
        SYNOPSYS_UNCONNECTED__1201, SYNOPSYS_UNCONNECTED__1202, 
        SYNOPSYS_UNCONNECTED__1203, SYNOPSYS_UNCONNECTED__1204, 
        SYNOPSYS_UNCONNECTED__1205, N66408, N66407, N66406, N66405, N66404, 
        N66403}) );
  hamming_N16000_CC2_DW01_add_220 add_2886_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63521, N63520, N63519, N63518, 
        N63517}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63534, 
        N63533, N63532, N63531, N63530}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1206, SYNOPSYS_UNCONNECTED__1207, 
        SYNOPSYS_UNCONNECTED__1208, SYNOPSYS_UNCONNECTED__1209, 
        SYNOPSYS_UNCONNECTED__1210, SYNOPSYS_UNCONNECTED__1211, 
        SYNOPSYS_UNCONNECTED__1212, N66395, N66394, N66393, N66392, N66391, 
        N66390}) );
  hamming_N16000_CC2_DW01_add_221 add_2887_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63495, N63494, N63493, N63492, 
        N63491}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63508, 
        N63507, N63506, N63505, N63504}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1213, SYNOPSYS_UNCONNECTED__1214, 
        SYNOPSYS_UNCONNECTED__1215, SYNOPSYS_UNCONNECTED__1216, 
        SYNOPSYS_UNCONNECTED__1217, SYNOPSYS_UNCONNECTED__1218, 
        SYNOPSYS_UNCONNECTED__1219, N66382, N66381, N66380, N66379, N66378, 
        N66377}) );
  hamming_N16000_CC2_DW01_add_222 add_2888_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63469, N63468, N63467, N63466, 
        N63465}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63482, 
        N63481, N63480, N63479, N63478}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1220, SYNOPSYS_UNCONNECTED__1221, 
        SYNOPSYS_UNCONNECTED__1222, SYNOPSYS_UNCONNECTED__1223, 
        SYNOPSYS_UNCONNECTED__1224, SYNOPSYS_UNCONNECTED__1225, 
        SYNOPSYS_UNCONNECTED__1226, N66369, N66368, N66367, N66366, N66365, 
        N66364}) );
  hamming_N16000_CC2_DW01_add_223 add_2889_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63443, N63442, N63441, N63440, 
        N63439}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63456, 
        N63455, N63454, N63453, N63452}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1227, SYNOPSYS_UNCONNECTED__1228, 
        SYNOPSYS_UNCONNECTED__1229, SYNOPSYS_UNCONNECTED__1230, 
        SYNOPSYS_UNCONNECTED__1231, SYNOPSYS_UNCONNECTED__1232, 
        SYNOPSYS_UNCONNECTED__1233, N66356, N66355, N66354, N66353, N66352, 
        N66351}) );
  hamming_N16000_CC2_DW01_add_224 add_2890_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63417, N63416, N63415, N63414, 
        N63413}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63430, 
        N63429, N63428, N63427, N63426}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1234, SYNOPSYS_UNCONNECTED__1235, 
        SYNOPSYS_UNCONNECTED__1236, SYNOPSYS_UNCONNECTED__1237, 
        SYNOPSYS_UNCONNECTED__1238, SYNOPSYS_UNCONNECTED__1239, 
        SYNOPSYS_UNCONNECTED__1240, N66343, N66342, N66341, N66340, N66339, 
        N66338}) );
  hamming_N16000_CC2_DW01_add_225 add_2891_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63391, N63390, N63389, N63388, 
        N63387}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63404, 
        N63403, N63402, N63401, N63400}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1241, SYNOPSYS_UNCONNECTED__1242, 
        SYNOPSYS_UNCONNECTED__1243, SYNOPSYS_UNCONNECTED__1244, 
        SYNOPSYS_UNCONNECTED__1245, SYNOPSYS_UNCONNECTED__1246, 
        SYNOPSYS_UNCONNECTED__1247, N66330, N66329, N66328, N66327, N66326, 
        N66325}) );
  hamming_N16000_CC2_DW01_add_226 add_2892_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63365, N63364, N63363, N63362, 
        N63361}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63378, 
        N63377, N63376, N63375, N63374}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1248, SYNOPSYS_UNCONNECTED__1249, 
        SYNOPSYS_UNCONNECTED__1250, SYNOPSYS_UNCONNECTED__1251, 
        SYNOPSYS_UNCONNECTED__1252, SYNOPSYS_UNCONNECTED__1253, 
        SYNOPSYS_UNCONNECTED__1254, N66317, N66316, N66315, N66314, N66313, 
        N66312}) );
  hamming_N16000_CC2_DW01_add_227 add_2893_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63339, N63338, N63337, N63336, 
        N63335}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63352, 
        N63351, N63350, N63349, N63348}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1255, SYNOPSYS_UNCONNECTED__1256, 
        SYNOPSYS_UNCONNECTED__1257, SYNOPSYS_UNCONNECTED__1258, 
        SYNOPSYS_UNCONNECTED__1259, SYNOPSYS_UNCONNECTED__1260, 
        SYNOPSYS_UNCONNECTED__1261, N66304, N66303, N66302, N66301, N66300, 
        N66299}) );
  hamming_N16000_CC2_DW01_add_228 add_2894_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63313, N63312, N63311, N63310, 
        N63309}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63326, 
        N63325, N63324, N63323, N63322}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1262, SYNOPSYS_UNCONNECTED__1263, 
        SYNOPSYS_UNCONNECTED__1264, SYNOPSYS_UNCONNECTED__1265, 
        SYNOPSYS_UNCONNECTED__1266, SYNOPSYS_UNCONNECTED__1267, 
        SYNOPSYS_UNCONNECTED__1268, N66291, N66290, N66289, N66288, N66287, 
        N66286}) );
  hamming_N16000_CC2_DW01_add_229 add_2895_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63287, N63286, N63285, N63284, 
        N63283}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63300, 
        N63299, N63298, N63297, N63296}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1269, SYNOPSYS_UNCONNECTED__1270, 
        SYNOPSYS_UNCONNECTED__1271, SYNOPSYS_UNCONNECTED__1272, 
        SYNOPSYS_UNCONNECTED__1273, SYNOPSYS_UNCONNECTED__1274, 
        SYNOPSYS_UNCONNECTED__1275, N66278, N66277, N66276, N66275, N66274, 
        N66273}) );
  hamming_N16000_CC2_DW01_add_230 add_2896_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63261, N63260, N63259, N63258, 
        N63257}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63274, 
        N63273, N63272, N63271, N63270}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1276, SYNOPSYS_UNCONNECTED__1277, 
        SYNOPSYS_UNCONNECTED__1278, SYNOPSYS_UNCONNECTED__1279, 
        SYNOPSYS_UNCONNECTED__1280, SYNOPSYS_UNCONNECTED__1281, 
        SYNOPSYS_UNCONNECTED__1282, N66265, N66264, N66263, N66262, N66261, 
        N66260}) );
  hamming_N16000_CC2_DW01_add_231 add_2897_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63235, N63234, N63233, N63232, 
        N63231}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63248, 
        N63247, N63246, N63245, N63244}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1283, SYNOPSYS_UNCONNECTED__1284, 
        SYNOPSYS_UNCONNECTED__1285, SYNOPSYS_UNCONNECTED__1286, 
        SYNOPSYS_UNCONNECTED__1287, SYNOPSYS_UNCONNECTED__1288, 
        SYNOPSYS_UNCONNECTED__1289, N66252, N66251, N66250, N66249, N66248, 
        N66247}) );
  hamming_N16000_CC2_DW01_add_232 add_2898_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63209, N63208, N63207, N63206, 
        N63205}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63222, 
        N63221, N63220, N63219, N63218}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1290, SYNOPSYS_UNCONNECTED__1291, 
        SYNOPSYS_UNCONNECTED__1292, SYNOPSYS_UNCONNECTED__1293, 
        SYNOPSYS_UNCONNECTED__1294, SYNOPSYS_UNCONNECTED__1295, 
        SYNOPSYS_UNCONNECTED__1296, N66239, N66238, N66237, N66236, N66235, 
        N66234}) );
  hamming_N16000_CC2_DW01_add_233 add_2899_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63183, N63182, N63181, N63180, 
        N63179}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63196, 
        N63195, N63194, N63193, N63192}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1297, SYNOPSYS_UNCONNECTED__1298, 
        SYNOPSYS_UNCONNECTED__1299, SYNOPSYS_UNCONNECTED__1300, 
        SYNOPSYS_UNCONNECTED__1301, SYNOPSYS_UNCONNECTED__1302, 
        SYNOPSYS_UNCONNECTED__1303, N66226, N66225, N66224, N66223, N66222, 
        N66221}) );
  hamming_N16000_CC2_DW01_add_234 add_2900_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63157, N63156, N63155, N63154, 
        N63153}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63170, 
        N63169, N63168, N63167, N63166}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1304, SYNOPSYS_UNCONNECTED__1305, 
        SYNOPSYS_UNCONNECTED__1306, SYNOPSYS_UNCONNECTED__1307, 
        SYNOPSYS_UNCONNECTED__1308, SYNOPSYS_UNCONNECTED__1309, 
        SYNOPSYS_UNCONNECTED__1310, N66213, N66212, N66211, N66210, N66209, 
        N66208}) );
  hamming_N16000_CC2_DW01_add_235 add_2901_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63131, N63130, N63129, N63128, 
        N63127}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63144, 
        N63143, N63142, N63141, N63140}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1311, SYNOPSYS_UNCONNECTED__1312, 
        SYNOPSYS_UNCONNECTED__1313, SYNOPSYS_UNCONNECTED__1314, 
        SYNOPSYS_UNCONNECTED__1315, SYNOPSYS_UNCONNECTED__1316, 
        SYNOPSYS_UNCONNECTED__1317, N66200, N66199, N66198, N66197, N66196, 
        N66195}) );
  hamming_N16000_CC2_DW01_add_236 add_2902_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63105, N63104, N63103, N63102, 
        N63101}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63118, 
        N63117, N63116, N63115, N63114}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1318, SYNOPSYS_UNCONNECTED__1319, 
        SYNOPSYS_UNCONNECTED__1320, SYNOPSYS_UNCONNECTED__1321, 
        SYNOPSYS_UNCONNECTED__1322, SYNOPSYS_UNCONNECTED__1323, 
        SYNOPSYS_UNCONNECTED__1324, N66187, N66186, N66185, N66184, N66183, 
        N66182}) );
  hamming_N16000_CC2_DW01_add_237 add_2903_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63079, N63078, N63077, N63076, 
        N63075}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63092, 
        N63091, N63090, N63089, N63088}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1325, SYNOPSYS_UNCONNECTED__1326, 
        SYNOPSYS_UNCONNECTED__1327, SYNOPSYS_UNCONNECTED__1328, 
        SYNOPSYS_UNCONNECTED__1329, SYNOPSYS_UNCONNECTED__1330, 
        SYNOPSYS_UNCONNECTED__1331, N66174, N66173, N66172, N66171, N66170, 
        N66169}) );
  hamming_N16000_CC2_DW01_add_238 add_2904_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63053, N63052, N63051, N63050, 
        N63049}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63066, 
        N63065, N63064, N63063, N63062}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1332, SYNOPSYS_UNCONNECTED__1333, 
        SYNOPSYS_UNCONNECTED__1334, SYNOPSYS_UNCONNECTED__1335, 
        SYNOPSYS_UNCONNECTED__1336, SYNOPSYS_UNCONNECTED__1337, 
        SYNOPSYS_UNCONNECTED__1338, N66161, N66160, N66159, N66158, N66157, 
        N66156}) );
  hamming_N16000_CC2_DW01_add_239 add_2905_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63027, N63026, N63025, N63024, 
        N63023}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63040, 
        N63039, N63038, N63037, N63036}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1339, SYNOPSYS_UNCONNECTED__1340, 
        SYNOPSYS_UNCONNECTED__1341, SYNOPSYS_UNCONNECTED__1342, 
        SYNOPSYS_UNCONNECTED__1343, SYNOPSYS_UNCONNECTED__1344, 
        SYNOPSYS_UNCONNECTED__1345, N66148, N66147, N66146, N66145, N66144, 
        N66143}) );
  hamming_N16000_CC2_DW01_add_240 add_2906_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63001, N63000, N62999, N62998, 
        N62997}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63014, 
        N63013, N63012, N63011, N63010}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1346, SYNOPSYS_UNCONNECTED__1347, 
        SYNOPSYS_UNCONNECTED__1348, SYNOPSYS_UNCONNECTED__1349, 
        SYNOPSYS_UNCONNECTED__1350, SYNOPSYS_UNCONNECTED__1351, 
        SYNOPSYS_UNCONNECTED__1352, N66135, N66134, N66133, N66132, N66131, 
        N66130}) );
  hamming_N16000_CC2_DW01_add_241 add_2907_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62975, N62974, N62973, N62972, 
        N62971}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62988, 
        N62987, N62986, N62985, N62984}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1353, SYNOPSYS_UNCONNECTED__1354, 
        SYNOPSYS_UNCONNECTED__1355, SYNOPSYS_UNCONNECTED__1356, 
        SYNOPSYS_UNCONNECTED__1357, SYNOPSYS_UNCONNECTED__1358, 
        SYNOPSYS_UNCONNECTED__1359, N66122, N66121, N66120, N66119, N66118, 
        N66117}) );
  hamming_N16000_CC2_DW01_add_242 add_2908_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62949, N62948, N62947, N62946, 
        N62945}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62962, 
        N62961, N62960, N62959, N62958}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1360, SYNOPSYS_UNCONNECTED__1361, 
        SYNOPSYS_UNCONNECTED__1362, SYNOPSYS_UNCONNECTED__1363, 
        SYNOPSYS_UNCONNECTED__1364, SYNOPSYS_UNCONNECTED__1365, 
        SYNOPSYS_UNCONNECTED__1366, N66109, N66108, N66107, N66106, N66105, 
        N66104}) );
  hamming_N16000_CC2_DW01_add_243 add_2909_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62923, N62922, N62921, N62920, 
        N62919}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62936, 
        N62935, N62934, N62933, N62932}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1367, SYNOPSYS_UNCONNECTED__1368, 
        SYNOPSYS_UNCONNECTED__1369, SYNOPSYS_UNCONNECTED__1370, 
        SYNOPSYS_UNCONNECTED__1371, SYNOPSYS_UNCONNECTED__1372, 
        SYNOPSYS_UNCONNECTED__1373, N66096, N66095, N66094, N66093, N66092, 
        N66091}) );
  hamming_N16000_CC2_DW01_add_244 add_2910_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62897, N62896, N62895, N62894, 
        N62893}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62910, 
        N62909, N62908, N62907, N62906}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1374, SYNOPSYS_UNCONNECTED__1375, 
        SYNOPSYS_UNCONNECTED__1376, SYNOPSYS_UNCONNECTED__1377, 
        SYNOPSYS_UNCONNECTED__1378, SYNOPSYS_UNCONNECTED__1379, 
        SYNOPSYS_UNCONNECTED__1380, N66083, N66082, N66081, N66080, N66079, 
        N66078}) );
  hamming_N16000_CC2_DW01_add_245 add_2911_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62871, N62870, N62869, N62868, 
        N62867}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62884, 
        N62883, N62882, N62881, N62880}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1381, SYNOPSYS_UNCONNECTED__1382, 
        SYNOPSYS_UNCONNECTED__1383, SYNOPSYS_UNCONNECTED__1384, 
        SYNOPSYS_UNCONNECTED__1385, SYNOPSYS_UNCONNECTED__1386, 
        SYNOPSYS_UNCONNECTED__1387, N66070, N66069, N66068, N66067, N66066, 
        N66065}) );
  hamming_N16000_CC2_DW01_add_246 add_2912_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62845, N62844, N62843, N62842, 
        N62841}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62858, 
        N62857, N62856, N62855, N62854}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1388, SYNOPSYS_UNCONNECTED__1389, 
        SYNOPSYS_UNCONNECTED__1390, SYNOPSYS_UNCONNECTED__1391, 
        SYNOPSYS_UNCONNECTED__1392, SYNOPSYS_UNCONNECTED__1393, 
        SYNOPSYS_UNCONNECTED__1394, N66057, N66056, N66055, N66054, N66053, 
        N66052}) );
  hamming_N16000_CC2_DW01_add_247 add_2913_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62819, N62818, N62817, N62816, 
        N62815}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62832, 
        N62831, N62830, N62829, N62828}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1395, SYNOPSYS_UNCONNECTED__1396, 
        SYNOPSYS_UNCONNECTED__1397, SYNOPSYS_UNCONNECTED__1398, 
        SYNOPSYS_UNCONNECTED__1399, SYNOPSYS_UNCONNECTED__1400, 
        SYNOPSYS_UNCONNECTED__1401, N66044, N66043, N66042, N66041, N66040, 
        N66039}) );
  hamming_N16000_CC2_DW01_add_248 add_2914_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62793, N62792, N62791, N62790, 
        N62789}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62806, 
        N62805, N62804, N62803, N62802}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1402, SYNOPSYS_UNCONNECTED__1403, 
        SYNOPSYS_UNCONNECTED__1404, SYNOPSYS_UNCONNECTED__1405, 
        SYNOPSYS_UNCONNECTED__1406, SYNOPSYS_UNCONNECTED__1407, 
        SYNOPSYS_UNCONNECTED__1408, N66031, N66030, N66029, N66028, N66027, 
        N66026}) );
  hamming_N16000_CC2_DW01_add_249 add_2915_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62767, N62766, N62765, N62764, 
        N62763}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62780, 
        N62779, N62778, N62777, N62776}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1409, SYNOPSYS_UNCONNECTED__1410, 
        SYNOPSYS_UNCONNECTED__1411, SYNOPSYS_UNCONNECTED__1412, 
        SYNOPSYS_UNCONNECTED__1413, SYNOPSYS_UNCONNECTED__1414, 
        SYNOPSYS_UNCONNECTED__1415, N66018, N66017, N66016, N66015, N66014, 
        N66013}) );
  hamming_N16000_CC2_DW01_add_250 add_2916_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62741, N62740, N62739, N62738, 
        N62737}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62754, 
        N62753, N62752, N62751, N62750}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1416, SYNOPSYS_UNCONNECTED__1417, 
        SYNOPSYS_UNCONNECTED__1418, SYNOPSYS_UNCONNECTED__1419, 
        SYNOPSYS_UNCONNECTED__1420, SYNOPSYS_UNCONNECTED__1421, 
        SYNOPSYS_UNCONNECTED__1422, N66005, N66004, N66003, N66002, N66001, 
        N66000}) );
  hamming_N16000_CC2_DW01_add_251 add_2917_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62715, N62714, N62713, N62712, 
        N62711}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62728, 
        N62727, N62726, N62725, N62724}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1423, SYNOPSYS_UNCONNECTED__1424, 
        SYNOPSYS_UNCONNECTED__1425, SYNOPSYS_UNCONNECTED__1426, 
        SYNOPSYS_UNCONNECTED__1427, SYNOPSYS_UNCONNECTED__1428, 
        SYNOPSYS_UNCONNECTED__1429, N65992, N65991, N65990, N65989, N65988, 
        N65987}) );
  hamming_N16000_CC2_DW01_add_252 add_2918_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62689, N62688, N62687, N62686, 
        N62685}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62702, 
        N62701, N62700, N62699, N62698}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1430, SYNOPSYS_UNCONNECTED__1431, 
        SYNOPSYS_UNCONNECTED__1432, SYNOPSYS_UNCONNECTED__1433, 
        SYNOPSYS_UNCONNECTED__1434, SYNOPSYS_UNCONNECTED__1435, 
        SYNOPSYS_UNCONNECTED__1436, N65979, N65978, N65977, N65976, N65975, 
        N65974}) );
  hamming_N16000_CC2_DW01_add_253 add_2919_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62663, N62662, N62661, N62660, 
        N62659}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62676, 
        N62675, N62674, N62673, N62672}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1437, SYNOPSYS_UNCONNECTED__1438, 
        SYNOPSYS_UNCONNECTED__1439, SYNOPSYS_UNCONNECTED__1440, 
        SYNOPSYS_UNCONNECTED__1441, SYNOPSYS_UNCONNECTED__1442, 
        SYNOPSYS_UNCONNECTED__1443, N65966, N65965, N65964, N65963, N65962, 
        N65961}) );
  hamming_N16000_CC2_DW01_add_254 add_2920_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62637, N62636, N62635, N62634, 
        N62633}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62650, 
        N62649, N62648, N62647, N62646}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1444, SYNOPSYS_UNCONNECTED__1445, 
        SYNOPSYS_UNCONNECTED__1446, SYNOPSYS_UNCONNECTED__1447, 
        SYNOPSYS_UNCONNECTED__1448, SYNOPSYS_UNCONNECTED__1449, 
        SYNOPSYS_UNCONNECTED__1450, N65953, N65952, N65951, N65950, N65949, 
        N65948}) );
  hamming_N16000_CC2_DW01_add_255 add_2921_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62611, N62610, N62609, N62608, 
        N62607}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62624, 
        N62623, N62622, N62621, N62620}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1451, SYNOPSYS_UNCONNECTED__1452, 
        SYNOPSYS_UNCONNECTED__1453, SYNOPSYS_UNCONNECTED__1454, 
        SYNOPSYS_UNCONNECTED__1455, SYNOPSYS_UNCONNECTED__1456, 
        SYNOPSYS_UNCONNECTED__1457, N65940, N65939, N65938, N65937, N65936, 
        N65935}) );
  hamming_N16000_CC2_DW01_add_256 add_2922_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62585, N62584, N62583, N62582, 
        N62581}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62598, 
        N62597, N62596, N62595, N62594}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1458, SYNOPSYS_UNCONNECTED__1459, 
        SYNOPSYS_UNCONNECTED__1460, SYNOPSYS_UNCONNECTED__1461, 
        SYNOPSYS_UNCONNECTED__1462, SYNOPSYS_UNCONNECTED__1463, 
        SYNOPSYS_UNCONNECTED__1464, N65927, N65926, N65925, N65924, N65923, 
        N65922}) );
  hamming_N16000_CC2_DW01_add_257 add_2923_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62559, N62558, N62557, N62556, 
        N62555}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62572, 
        N62571, N62570, N62569, N62568}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1465, SYNOPSYS_UNCONNECTED__1466, 
        SYNOPSYS_UNCONNECTED__1467, SYNOPSYS_UNCONNECTED__1468, 
        SYNOPSYS_UNCONNECTED__1469, SYNOPSYS_UNCONNECTED__1470, 
        SYNOPSYS_UNCONNECTED__1471, N65914, N65913, N65912, N65911, N65910, 
        N65909}) );
  hamming_N16000_CC2_DW01_add_258 add_2924_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62533, N62532, N62531, N62530, 
        N62529}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62546, 
        N62545, N62544, N62543, N62542}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1472, SYNOPSYS_UNCONNECTED__1473, 
        SYNOPSYS_UNCONNECTED__1474, SYNOPSYS_UNCONNECTED__1475, 
        SYNOPSYS_UNCONNECTED__1476, SYNOPSYS_UNCONNECTED__1477, 
        SYNOPSYS_UNCONNECTED__1478, N65901, N65900, N65899, N65898, N65897, 
        N65896}) );
  hamming_N16000_CC2_DW01_add_259 add_2925_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62507, N62506, N62505, N62504, 
        N62503}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62520, 
        N62519, N62518, N62517, N62516}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1479, SYNOPSYS_UNCONNECTED__1480, 
        SYNOPSYS_UNCONNECTED__1481, SYNOPSYS_UNCONNECTED__1482, 
        SYNOPSYS_UNCONNECTED__1483, SYNOPSYS_UNCONNECTED__1484, 
        SYNOPSYS_UNCONNECTED__1485, N65888, N65887, N65886, N65885, N65884, 
        N65883}) );
  hamming_N16000_CC2_DW01_add_260 add_2926_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62481, N62480, N62479, N62478, 
        N62477}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62494, 
        N62493, N62492, N62491, N62490}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1486, SYNOPSYS_UNCONNECTED__1487, 
        SYNOPSYS_UNCONNECTED__1488, SYNOPSYS_UNCONNECTED__1489, 
        SYNOPSYS_UNCONNECTED__1490, SYNOPSYS_UNCONNECTED__1491, 
        SYNOPSYS_UNCONNECTED__1492, N65875, N65874, N65873, N65872, N65871, 
        N65870}) );
  hamming_N16000_CC2_DW01_add_261 add_2927_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62455, N62454, N62453, N62452, 
        N62451}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62468, 
        N62467, N62466, N62465, N62464}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1493, SYNOPSYS_UNCONNECTED__1494, 
        SYNOPSYS_UNCONNECTED__1495, SYNOPSYS_UNCONNECTED__1496, 
        SYNOPSYS_UNCONNECTED__1497, SYNOPSYS_UNCONNECTED__1498, 
        SYNOPSYS_UNCONNECTED__1499, N65862, N65861, N65860, N65859, N65858, 
        N65857}) );
  hamming_N16000_CC2_DW01_add_262 add_2928_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62429, N62428, N62427, N62426, 
        N62425}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62442, 
        N62441, N62440, N62439, N62438}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1500, SYNOPSYS_UNCONNECTED__1501, 
        SYNOPSYS_UNCONNECTED__1502, SYNOPSYS_UNCONNECTED__1503, 
        SYNOPSYS_UNCONNECTED__1504, SYNOPSYS_UNCONNECTED__1505, 
        SYNOPSYS_UNCONNECTED__1506, N65849, N65848, N65847, N65846, N65845, 
        N65844}) );
  hamming_N16000_CC2_DW01_add_263 add_2929_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62403, N62402, N62401, N62400, 
        N62399}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62416, 
        N62415, N62414, N62413, N62412}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1507, SYNOPSYS_UNCONNECTED__1508, 
        SYNOPSYS_UNCONNECTED__1509, SYNOPSYS_UNCONNECTED__1510, 
        SYNOPSYS_UNCONNECTED__1511, SYNOPSYS_UNCONNECTED__1512, 
        SYNOPSYS_UNCONNECTED__1513, N65836, N65835, N65834, N65833, N65832, 
        N65831}) );
  hamming_N16000_CC2_DW01_add_264 add_2930_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62377, N62376, N62375, N62374, 
        N62373}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62390, 
        N62389, N62388, N62387, N62386}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1514, SYNOPSYS_UNCONNECTED__1515, 
        SYNOPSYS_UNCONNECTED__1516, SYNOPSYS_UNCONNECTED__1517, 
        SYNOPSYS_UNCONNECTED__1518, SYNOPSYS_UNCONNECTED__1519, 
        SYNOPSYS_UNCONNECTED__1520, N65823, N65822, N65821, N65820, N65819, 
        N65818}) );
  hamming_N16000_CC2_DW01_add_265 add_2931_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62351, N62350, N62349, N62348, 
        N62347}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62364, 
        N62363, N62362, N62361, N62360}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1521, SYNOPSYS_UNCONNECTED__1522, 
        SYNOPSYS_UNCONNECTED__1523, SYNOPSYS_UNCONNECTED__1524, 
        SYNOPSYS_UNCONNECTED__1525, SYNOPSYS_UNCONNECTED__1526, 
        SYNOPSYS_UNCONNECTED__1527, N65810, N65809, N65808, N65807, N65806, 
        N65805}) );
  hamming_N16000_CC2_DW01_add_266 add_2932_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62325, N62324, N62323, N62322, 
        N62321}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62338, 
        N62337, N62336, N62335, N62334}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1528, SYNOPSYS_UNCONNECTED__1529, 
        SYNOPSYS_UNCONNECTED__1530, SYNOPSYS_UNCONNECTED__1531, 
        SYNOPSYS_UNCONNECTED__1532, SYNOPSYS_UNCONNECTED__1533, 
        SYNOPSYS_UNCONNECTED__1534, N65797, N65796, N65795, N65794, N65793, 
        N65792}) );
  hamming_N16000_CC2_DW01_add_267 add_2933_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62299, N62298, N62297, N62296, 
        N62295}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62312, 
        N62311, N62310, N62309, N62308}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1535, SYNOPSYS_UNCONNECTED__1536, 
        SYNOPSYS_UNCONNECTED__1537, SYNOPSYS_UNCONNECTED__1538, 
        SYNOPSYS_UNCONNECTED__1539, SYNOPSYS_UNCONNECTED__1540, 
        SYNOPSYS_UNCONNECTED__1541, N65784, N65783, N65782, N65781, N65780, 
        N65779}) );
  hamming_N16000_CC2_DW01_add_268 add_2934_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62273, N62272, N62271, N62270, 
        N62269}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62286, 
        N62285, N62284, N62283, N62282}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1542, SYNOPSYS_UNCONNECTED__1543, 
        SYNOPSYS_UNCONNECTED__1544, SYNOPSYS_UNCONNECTED__1545, 
        SYNOPSYS_UNCONNECTED__1546, SYNOPSYS_UNCONNECTED__1547, 
        SYNOPSYS_UNCONNECTED__1548, N65771, N65770, N65769, N65768, N65767, 
        N65766}) );
  hamming_N16000_CC2_DW01_add_269 add_2935_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62247, N62246, N62245, N62244, 
        N62243}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62260, 
        N62259, N62258, N62257, N62256}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1549, SYNOPSYS_UNCONNECTED__1550, 
        SYNOPSYS_UNCONNECTED__1551, SYNOPSYS_UNCONNECTED__1552, 
        SYNOPSYS_UNCONNECTED__1553, SYNOPSYS_UNCONNECTED__1554, 
        SYNOPSYS_UNCONNECTED__1555, N65758, N65757, N65756, N65755, N65754, 
        N65753}) );
  hamming_N16000_CC2_DW01_add_270 add_2936_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62221, N62220, N62219, N62218, 
        N62217}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62234, 
        N62233, N62232, N62231, N62230}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1556, SYNOPSYS_UNCONNECTED__1557, 
        SYNOPSYS_UNCONNECTED__1558, SYNOPSYS_UNCONNECTED__1559, 
        SYNOPSYS_UNCONNECTED__1560, SYNOPSYS_UNCONNECTED__1561, 
        SYNOPSYS_UNCONNECTED__1562, N65745, N65744, N65743, N65742, N65741, 
        N65740}) );
  hamming_N16000_CC2_DW01_add_271 add_2937_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62195, N62194, N62193, N62192, 
        N62191}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62208, 
        N62207, N62206, N62205, N62204}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1563, SYNOPSYS_UNCONNECTED__1564, 
        SYNOPSYS_UNCONNECTED__1565, SYNOPSYS_UNCONNECTED__1566, 
        SYNOPSYS_UNCONNECTED__1567, SYNOPSYS_UNCONNECTED__1568, 
        SYNOPSYS_UNCONNECTED__1569, N65732, N65731, N65730, N65729, N65728, 
        N65727}) );
  hamming_N16000_CC2_DW01_add_272 add_2938_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62169, N62168, N62167, N62166, 
        N62165}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62182, 
        N62181, N62180, N62179, N62178}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1570, SYNOPSYS_UNCONNECTED__1571, 
        SYNOPSYS_UNCONNECTED__1572, SYNOPSYS_UNCONNECTED__1573, 
        SYNOPSYS_UNCONNECTED__1574, SYNOPSYS_UNCONNECTED__1575, 
        SYNOPSYS_UNCONNECTED__1576, N65719, N65718, N65717, N65716, N65715, 
        N65714}) );
  hamming_N16000_CC2_DW01_add_273 add_2939_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62143, N62142, N62141, N62140, 
        N62139}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62156, 
        N62155, N62154, N62153, N62152}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1577, SYNOPSYS_UNCONNECTED__1578, 
        SYNOPSYS_UNCONNECTED__1579, SYNOPSYS_UNCONNECTED__1580, 
        SYNOPSYS_UNCONNECTED__1581, SYNOPSYS_UNCONNECTED__1582, 
        SYNOPSYS_UNCONNECTED__1583, N65706, N65705, N65704, N65703, N65702, 
        N65701}) );
  hamming_N16000_CC2_DW01_add_274 add_2940_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62117, N62116, N62115, N62114, 
        N62113}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62130, 
        N62129, N62128, N62127, N62126}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1584, SYNOPSYS_UNCONNECTED__1585, 
        SYNOPSYS_UNCONNECTED__1586, SYNOPSYS_UNCONNECTED__1587, 
        SYNOPSYS_UNCONNECTED__1588, SYNOPSYS_UNCONNECTED__1589, 
        SYNOPSYS_UNCONNECTED__1590, N65693, N65692, N65691, N65690, N65689, 
        N65688}) );
  hamming_N16000_CC2_DW01_add_275 add_2941_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62091, N62090, N62089, N62088, 
        N62087}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62104, 
        N62103, N62102, N62101, N62100}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1591, SYNOPSYS_UNCONNECTED__1592, 
        SYNOPSYS_UNCONNECTED__1593, SYNOPSYS_UNCONNECTED__1594, 
        SYNOPSYS_UNCONNECTED__1595, SYNOPSYS_UNCONNECTED__1596, 
        SYNOPSYS_UNCONNECTED__1597, N65680, N65679, N65678, N65677, N65676, 
        N65675}) );
  hamming_N16000_CC2_DW01_add_276 add_2942_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62065, N62064, N62063, N62062, 
        N62061}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62078, 
        N62077, N62076, N62075, N62074}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1598, SYNOPSYS_UNCONNECTED__1599, 
        SYNOPSYS_UNCONNECTED__1600, SYNOPSYS_UNCONNECTED__1601, 
        SYNOPSYS_UNCONNECTED__1602, SYNOPSYS_UNCONNECTED__1603, 
        SYNOPSYS_UNCONNECTED__1604, N65667, N65666, N65665, N65664, N65663, 
        N65662}) );
  hamming_N16000_CC2_DW01_add_277 add_2943_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62039, N62038, N62037, N62036, 
        N62035}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62052, 
        N62051, N62050, N62049, N62048}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1605, SYNOPSYS_UNCONNECTED__1606, 
        SYNOPSYS_UNCONNECTED__1607, SYNOPSYS_UNCONNECTED__1608, 
        SYNOPSYS_UNCONNECTED__1609, SYNOPSYS_UNCONNECTED__1610, 
        SYNOPSYS_UNCONNECTED__1611, N65654, N65653, N65652, N65651, N65650, 
        N65649}) );
  hamming_N16000_CC2_DW01_add_278 add_2944_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62013, N62012, N62011, N62010, 
        N62009}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62026, 
        N62025, N62024, N62023, N62022}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1612, SYNOPSYS_UNCONNECTED__1613, 
        SYNOPSYS_UNCONNECTED__1614, SYNOPSYS_UNCONNECTED__1615, 
        SYNOPSYS_UNCONNECTED__1616, SYNOPSYS_UNCONNECTED__1617, 
        SYNOPSYS_UNCONNECTED__1618, N65641, N65640, N65639, N65638, N65637, 
        N65636}) );
  hamming_N16000_CC2_DW01_add_279 add_2945_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61987, N61986, N61985, N61984, 
        N61983}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62000, 
        N61999, N61998, N61997, N61996}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1619, SYNOPSYS_UNCONNECTED__1620, 
        SYNOPSYS_UNCONNECTED__1621, SYNOPSYS_UNCONNECTED__1622, 
        SYNOPSYS_UNCONNECTED__1623, SYNOPSYS_UNCONNECTED__1624, 
        SYNOPSYS_UNCONNECTED__1625, N65628, N65627, N65626, N65625, N65624, 
        N65623}) );
  hamming_N16000_CC2_DW01_add_280 add_2946_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61961, N61960, N61959, N61958, 
        N61957}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61974, 
        N61973, N61972, N61971, N61970}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1626, SYNOPSYS_UNCONNECTED__1627, 
        SYNOPSYS_UNCONNECTED__1628, SYNOPSYS_UNCONNECTED__1629, 
        SYNOPSYS_UNCONNECTED__1630, SYNOPSYS_UNCONNECTED__1631, 
        SYNOPSYS_UNCONNECTED__1632, N65615, N65614, N65613, N65612, N65611, 
        N65610}) );
  hamming_N16000_CC2_DW01_add_281 add_2947_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61935, N61934, N61933, N61932, 
        N61931}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61948, 
        N61947, N61946, N61945, N61944}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1633, SYNOPSYS_UNCONNECTED__1634, 
        SYNOPSYS_UNCONNECTED__1635, SYNOPSYS_UNCONNECTED__1636, 
        SYNOPSYS_UNCONNECTED__1637, SYNOPSYS_UNCONNECTED__1638, 
        SYNOPSYS_UNCONNECTED__1639, N65602, N65601, N65600, N65599, N65598, 
        N65597}) );
  hamming_N16000_CC2_DW01_add_282 add_2948_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61909, N61908, N61907, N61906, 
        N61905}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61922, 
        N61921, N61920, N61919, N61918}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1640, SYNOPSYS_UNCONNECTED__1641, 
        SYNOPSYS_UNCONNECTED__1642, SYNOPSYS_UNCONNECTED__1643, 
        SYNOPSYS_UNCONNECTED__1644, SYNOPSYS_UNCONNECTED__1645, 
        SYNOPSYS_UNCONNECTED__1646, N65589, N65588, N65587, N65586, N65585, 
        N65584}) );
  hamming_N16000_CC2_DW01_add_283 add_2949_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61883, N61882, N61881, N61880, 
        N61879}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61896, 
        N61895, N61894, N61893, N61892}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1647, SYNOPSYS_UNCONNECTED__1648, 
        SYNOPSYS_UNCONNECTED__1649, SYNOPSYS_UNCONNECTED__1650, 
        SYNOPSYS_UNCONNECTED__1651, SYNOPSYS_UNCONNECTED__1652, 
        SYNOPSYS_UNCONNECTED__1653, N65576, N65575, N65574, N65573, N65572, 
        N65571}) );
  hamming_N16000_CC2_DW01_add_284 add_2950_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61857, N61856, N61855, N61854, 
        N61853}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61870, 
        N61869, N61868, N61867, N61866}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1654, SYNOPSYS_UNCONNECTED__1655, 
        SYNOPSYS_UNCONNECTED__1656, SYNOPSYS_UNCONNECTED__1657, 
        SYNOPSYS_UNCONNECTED__1658, SYNOPSYS_UNCONNECTED__1659, 
        SYNOPSYS_UNCONNECTED__1660, N65563, N65562, N65561, N65560, N65559, 
        N65558}) );
  hamming_N16000_CC2_DW01_add_285 add_2951_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61831, N61830, N61829, N61828, 
        N61827}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61844, 
        N61843, N61842, N61841, N61840}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1661, SYNOPSYS_UNCONNECTED__1662, 
        SYNOPSYS_UNCONNECTED__1663, SYNOPSYS_UNCONNECTED__1664, 
        SYNOPSYS_UNCONNECTED__1665, SYNOPSYS_UNCONNECTED__1666, 
        SYNOPSYS_UNCONNECTED__1667, N65550, N65549, N65548, N65547, N65546, 
        N65545}) );
  hamming_N16000_CC2_DW01_add_286 add_2952_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61805, N61804, N61803, N61802, 
        N61801}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61818, 
        N61817, N61816, N61815, N61814}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1668, SYNOPSYS_UNCONNECTED__1669, 
        SYNOPSYS_UNCONNECTED__1670, SYNOPSYS_UNCONNECTED__1671, 
        SYNOPSYS_UNCONNECTED__1672, SYNOPSYS_UNCONNECTED__1673, 
        SYNOPSYS_UNCONNECTED__1674, N65537, N65536, N65535, N65534, N65533, 
        N65532}) );
  hamming_N16000_CC2_DW01_add_287 add_2953_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61779, N61778, N61777, N61776, 
        N61775}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61792, 
        N61791, N61790, N61789, N61788}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1675, SYNOPSYS_UNCONNECTED__1676, 
        SYNOPSYS_UNCONNECTED__1677, SYNOPSYS_UNCONNECTED__1678, 
        SYNOPSYS_UNCONNECTED__1679, SYNOPSYS_UNCONNECTED__1680, 
        SYNOPSYS_UNCONNECTED__1681, N65524, N65523, N65522, N65521, N65520, 
        N65519}) );
  hamming_N16000_CC2_DW01_add_288 add_2954_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61753, N61752, N61751, N61750, 
        N61749}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61766, 
        N61765, N61764, N61763, N61762}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1682, SYNOPSYS_UNCONNECTED__1683, 
        SYNOPSYS_UNCONNECTED__1684, SYNOPSYS_UNCONNECTED__1685, 
        SYNOPSYS_UNCONNECTED__1686, SYNOPSYS_UNCONNECTED__1687, 
        SYNOPSYS_UNCONNECTED__1688, N65511, N65510, N65509, N65508, N65507, 
        N65506}) );
  hamming_N16000_CC2_DW01_add_289 add_2955_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61727, N61726, N61725, N61724, 
        N61723}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61740, 
        N61739, N61738, N61737, N61736}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1689, SYNOPSYS_UNCONNECTED__1690, 
        SYNOPSYS_UNCONNECTED__1691, SYNOPSYS_UNCONNECTED__1692, 
        SYNOPSYS_UNCONNECTED__1693, SYNOPSYS_UNCONNECTED__1694, 
        SYNOPSYS_UNCONNECTED__1695, N65498, N65497, N65496, N65495, N65494, 
        N65493}) );
  hamming_N16000_CC2_DW01_add_290 add_2956_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61701, N61700, N61699, N61698, 
        N61697}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61714, 
        N61713, N61712, N61711, N61710}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1696, SYNOPSYS_UNCONNECTED__1697, 
        SYNOPSYS_UNCONNECTED__1698, SYNOPSYS_UNCONNECTED__1699, 
        SYNOPSYS_UNCONNECTED__1700, SYNOPSYS_UNCONNECTED__1701, 
        SYNOPSYS_UNCONNECTED__1702, N65485, N65484, N65483, N65482, N65481, 
        N65480}) );
  hamming_N16000_CC2_DW01_add_291 add_2957_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61675, N61674, N61673, N61672, 
        N61671}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61688, 
        N61687, N61686, N61685, N61684}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1703, SYNOPSYS_UNCONNECTED__1704, 
        SYNOPSYS_UNCONNECTED__1705, SYNOPSYS_UNCONNECTED__1706, 
        SYNOPSYS_UNCONNECTED__1707, SYNOPSYS_UNCONNECTED__1708, 
        SYNOPSYS_UNCONNECTED__1709, N65472, N65471, N65470, N65469, N65468, 
        N65467}) );
  hamming_N16000_CC2_DW01_add_292 add_2958_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61649, N61648, N61647, N61646, 
        N61645}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61662, 
        N61661, N61660, N61659, N61658}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1710, SYNOPSYS_UNCONNECTED__1711, 
        SYNOPSYS_UNCONNECTED__1712, SYNOPSYS_UNCONNECTED__1713, 
        SYNOPSYS_UNCONNECTED__1714, SYNOPSYS_UNCONNECTED__1715, 
        SYNOPSYS_UNCONNECTED__1716, N65459, N65458, N65457, N65456, N65455, 
        N65454}) );
  hamming_N16000_CC2_DW01_add_293 add_2959_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61623, N61622, N61621, N61620, 
        N61619}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61636, 
        N61635, N61634, N61633, N61632}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1717, SYNOPSYS_UNCONNECTED__1718, 
        SYNOPSYS_UNCONNECTED__1719, SYNOPSYS_UNCONNECTED__1720, 
        SYNOPSYS_UNCONNECTED__1721, SYNOPSYS_UNCONNECTED__1722, 
        SYNOPSYS_UNCONNECTED__1723, N65446, N65445, N65444, N65443, N65442, 
        N65441}) );
  hamming_N16000_CC2_DW01_add_294 add_2960_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61597, N61596, N61595, N61594, 
        N61593}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61610, 
        N61609, N61608, N61607, N61606}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1724, SYNOPSYS_UNCONNECTED__1725, 
        SYNOPSYS_UNCONNECTED__1726, SYNOPSYS_UNCONNECTED__1727, 
        SYNOPSYS_UNCONNECTED__1728, SYNOPSYS_UNCONNECTED__1729, 
        SYNOPSYS_UNCONNECTED__1730, N65433, N65432, N65431, N65430, N65429, 
        N65428}) );
  hamming_N16000_CC2_DW01_add_295 add_2961_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61571, N61570, N61569, N61568, 
        N61567}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61584, 
        N61583, N61582, N61581, N61580}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1731, SYNOPSYS_UNCONNECTED__1732, 
        SYNOPSYS_UNCONNECTED__1733, SYNOPSYS_UNCONNECTED__1734, 
        SYNOPSYS_UNCONNECTED__1735, SYNOPSYS_UNCONNECTED__1736, 
        SYNOPSYS_UNCONNECTED__1737, N65420, N65419, N65418, N65417, N65416, 
        N65415}) );
  hamming_N16000_CC2_DW01_add_296 add_2962_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61545, N61544, N61543, N61542, 
        N61541}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61558, 
        N61557, N61556, N61555, N61554}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1738, SYNOPSYS_UNCONNECTED__1739, 
        SYNOPSYS_UNCONNECTED__1740, SYNOPSYS_UNCONNECTED__1741, 
        SYNOPSYS_UNCONNECTED__1742, SYNOPSYS_UNCONNECTED__1743, 
        SYNOPSYS_UNCONNECTED__1744, N65407, N65406, N65405, N65404, N65403, 
        N65402}) );
  hamming_N16000_CC2_DW01_add_297 add_2963_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61519, N61518, N61517, N61516, 
        N61515}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61532, 
        N61531, N61530, N61529, N61528}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1745, SYNOPSYS_UNCONNECTED__1746, 
        SYNOPSYS_UNCONNECTED__1747, SYNOPSYS_UNCONNECTED__1748, 
        SYNOPSYS_UNCONNECTED__1749, SYNOPSYS_UNCONNECTED__1750, 
        SYNOPSYS_UNCONNECTED__1751, N65394, N65393, N65392, N65391, N65390, 
        N65389}) );
  hamming_N16000_CC2_DW01_add_298 add_2964_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61493, N61492, N61491, N61490, 
        N61489}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61506, 
        N61505, N61504, N61503, N61502}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1752, SYNOPSYS_UNCONNECTED__1753, 
        SYNOPSYS_UNCONNECTED__1754, SYNOPSYS_UNCONNECTED__1755, 
        SYNOPSYS_UNCONNECTED__1756, SYNOPSYS_UNCONNECTED__1757, 
        SYNOPSYS_UNCONNECTED__1758, N65381, N65380, N65379, N65378, N65377, 
        N65376}) );
  hamming_N16000_CC2_DW01_add_299 add_2965_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61467, N61466, N61465, N61464, 
        N61463}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61480, 
        N61479, N61478, N61477, N61476}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1759, SYNOPSYS_UNCONNECTED__1760, 
        SYNOPSYS_UNCONNECTED__1761, SYNOPSYS_UNCONNECTED__1762, 
        SYNOPSYS_UNCONNECTED__1763, SYNOPSYS_UNCONNECTED__1764, 
        SYNOPSYS_UNCONNECTED__1765, N65368, N65367, N65366, N65365, N65364, 
        N65363}) );
  hamming_N16000_CC2_DW01_add_300 add_2966_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61441, N61440, N61439, N61438, 
        N61437}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61454, 
        N61453, N61452, N61451, N61450}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1766, SYNOPSYS_UNCONNECTED__1767, 
        SYNOPSYS_UNCONNECTED__1768, SYNOPSYS_UNCONNECTED__1769, 
        SYNOPSYS_UNCONNECTED__1770, SYNOPSYS_UNCONNECTED__1771, 
        SYNOPSYS_UNCONNECTED__1772, N65355, N65354, N65353, N65352, N65351, 
        N65350}) );
  hamming_N16000_CC2_DW01_add_301 add_2967_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61415, N61414, N61413, N61412, 
        N61411}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61428, 
        N61427, N61426, N61425, N61424}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1773, SYNOPSYS_UNCONNECTED__1774, 
        SYNOPSYS_UNCONNECTED__1775, SYNOPSYS_UNCONNECTED__1776, 
        SYNOPSYS_UNCONNECTED__1777, SYNOPSYS_UNCONNECTED__1778, 
        SYNOPSYS_UNCONNECTED__1779, N65342, N65341, N65340, N65339, N65338, 
        N65337}) );
  hamming_N16000_CC2_DW01_add_302 add_2968_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61389, N61388, N61387, N61386, 
        N61385}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61402, 
        N61401, N61400, N61399, N61398}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1780, SYNOPSYS_UNCONNECTED__1781, 
        SYNOPSYS_UNCONNECTED__1782, SYNOPSYS_UNCONNECTED__1783, 
        SYNOPSYS_UNCONNECTED__1784, SYNOPSYS_UNCONNECTED__1785, 
        SYNOPSYS_UNCONNECTED__1786, N65329, N65328, N65327, N65326, N65325, 
        N65324}) );
  hamming_N16000_CC2_DW01_add_303 add_2969_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61363, N61362, N61361, N61360, 
        N61359}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61376, 
        N61375, N61374, N61373, N61372}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1787, SYNOPSYS_UNCONNECTED__1788, 
        SYNOPSYS_UNCONNECTED__1789, SYNOPSYS_UNCONNECTED__1790, 
        SYNOPSYS_UNCONNECTED__1791, SYNOPSYS_UNCONNECTED__1792, 
        SYNOPSYS_UNCONNECTED__1793, N65316, N65315, N65314, N65313, N65312, 
        N65311}) );
  hamming_N16000_CC2_DW01_add_304 add_2970_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61337, N61336, N61335, N61334, 
        N61333}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61350, 
        N61349, N61348, N61347, N61346}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1794, SYNOPSYS_UNCONNECTED__1795, 
        SYNOPSYS_UNCONNECTED__1796, SYNOPSYS_UNCONNECTED__1797, 
        SYNOPSYS_UNCONNECTED__1798, SYNOPSYS_UNCONNECTED__1799, 
        SYNOPSYS_UNCONNECTED__1800, N65303, N65302, N65301, N65300, N65299, 
        N65298}) );
  hamming_N16000_CC2_DW01_add_305 add_2971_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61311, N61310, N61309, N61308, 
        N61307}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61324, 
        N61323, N61322, N61321, N61320}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1801, SYNOPSYS_UNCONNECTED__1802, 
        SYNOPSYS_UNCONNECTED__1803, SYNOPSYS_UNCONNECTED__1804, 
        SYNOPSYS_UNCONNECTED__1805, SYNOPSYS_UNCONNECTED__1806, 
        SYNOPSYS_UNCONNECTED__1807, N65290, N65289, N65288, N65287, N65286, 
        N65285}) );
  hamming_N16000_CC2_DW01_add_306 add_2972_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61285, N61284, N61283, N61282, 
        N61281}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61298, 
        N61297, N61296, N61295, N61294}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1808, SYNOPSYS_UNCONNECTED__1809, 
        SYNOPSYS_UNCONNECTED__1810, SYNOPSYS_UNCONNECTED__1811, 
        SYNOPSYS_UNCONNECTED__1812, SYNOPSYS_UNCONNECTED__1813, 
        SYNOPSYS_UNCONNECTED__1814, N65277, N65276, N65275, N65274, N65273, 
        N65272}) );
  hamming_N16000_CC2_DW01_add_307 add_2973_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61259, N61258, N61257, N61256, 
        N61255}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61272, 
        N61271, N61270, N61269, N61268}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1815, SYNOPSYS_UNCONNECTED__1816, 
        SYNOPSYS_UNCONNECTED__1817, SYNOPSYS_UNCONNECTED__1818, 
        SYNOPSYS_UNCONNECTED__1819, SYNOPSYS_UNCONNECTED__1820, 
        SYNOPSYS_UNCONNECTED__1821, N65264, N65263, N65262, N65261, N65260, 
        N65259}) );
  hamming_N16000_CC2_DW01_add_308 add_2974_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61233, N61232, N61231, N61230, 
        N61229}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61246, 
        N61245, N61244, N61243, N61242}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1822, SYNOPSYS_UNCONNECTED__1823, 
        SYNOPSYS_UNCONNECTED__1824, SYNOPSYS_UNCONNECTED__1825, 
        SYNOPSYS_UNCONNECTED__1826, SYNOPSYS_UNCONNECTED__1827, 
        SYNOPSYS_UNCONNECTED__1828, N65251, N65250, N65249, N65248, N65247, 
        N65246}) );
  hamming_N16000_CC2_DW01_add_309 add_2975_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61207, N61206, N61205, N61204, 
        N61203}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61220, 
        N61219, N61218, N61217, N61216}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1829, SYNOPSYS_UNCONNECTED__1830, 
        SYNOPSYS_UNCONNECTED__1831, SYNOPSYS_UNCONNECTED__1832, 
        SYNOPSYS_UNCONNECTED__1833, SYNOPSYS_UNCONNECTED__1834, 
        SYNOPSYS_UNCONNECTED__1835, N65238, N65237, N65236, N65235, N65234, 
        N65233}) );
  hamming_N16000_CC2_DW01_add_310 add_2976_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61181, N61180, N61179, N61178, 
        N61177}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61194, 
        N61193, N61192, N61191, N61190}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1836, SYNOPSYS_UNCONNECTED__1837, 
        SYNOPSYS_UNCONNECTED__1838, SYNOPSYS_UNCONNECTED__1839, 
        SYNOPSYS_UNCONNECTED__1840, SYNOPSYS_UNCONNECTED__1841, 
        SYNOPSYS_UNCONNECTED__1842, N65225, N65224, N65223, N65222, N65221, 
        N65220}) );
  hamming_N16000_CC2_DW01_add_311 add_2977_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61155, N61154, N61153, N61152, 
        N61151}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61168, 
        N61167, N61166, N61165, N61164}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1843, SYNOPSYS_UNCONNECTED__1844, 
        SYNOPSYS_UNCONNECTED__1845, SYNOPSYS_UNCONNECTED__1846, 
        SYNOPSYS_UNCONNECTED__1847, SYNOPSYS_UNCONNECTED__1848, 
        SYNOPSYS_UNCONNECTED__1849, N65212, N65211, N65210, N65209, N65208, 
        N65207}) );
  hamming_N16000_CC2_DW01_add_312 add_2978_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61129, N61128, N61127, N61126, 
        N61125}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61142, 
        N61141, N61140, N61139, N61138}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1850, SYNOPSYS_UNCONNECTED__1851, 
        SYNOPSYS_UNCONNECTED__1852, SYNOPSYS_UNCONNECTED__1853, 
        SYNOPSYS_UNCONNECTED__1854, SYNOPSYS_UNCONNECTED__1855, 
        SYNOPSYS_UNCONNECTED__1856, N65199, N65198, N65197, N65196, N65195, 
        N65194}) );
  hamming_N16000_CC2_DW01_add_313 add_2979_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61103, N61102, N61101, N61100, 
        N61099}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61116, 
        N61115, N61114, N61113, N61112}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1857, SYNOPSYS_UNCONNECTED__1858, 
        SYNOPSYS_UNCONNECTED__1859, SYNOPSYS_UNCONNECTED__1860, 
        SYNOPSYS_UNCONNECTED__1861, SYNOPSYS_UNCONNECTED__1862, 
        SYNOPSYS_UNCONNECTED__1863, N65186, N65185, N65184, N65183, N65182, 
        N65181}) );
  hamming_N16000_CC2_DW01_add_314 add_2980_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61077, N61076, N61075, N61074, 
        N61073}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61090, 
        N61089, N61088, N61087, N61086}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1864, SYNOPSYS_UNCONNECTED__1865, 
        SYNOPSYS_UNCONNECTED__1866, SYNOPSYS_UNCONNECTED__1867, 
        SYNOPSYS_UNCONNECTED__1868, SYNOPSYS_UNCONNECTED__1869, 
        SYNOPSYS_UNCONNECTED__1870, N65173, N65172, N65171, N65170, N65169, 
        N65168}) );
  hamming_N16000_CC2_DW01_add_315 add_2981_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61051, N61050, N61049, N61048, 
        N61047}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61064, 
        N61063, N61062, N61061, N61060}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1871, SYNOPSYS_UNCONNECTED__1872, 
        SYNOPSYS_UNCONNECTED__1873, SYNOPSYS_UNCONNECTED__1874, 
        SYNOPSYS_UNCONNECTED__1875, SYNOPSYS_UNCONNECTED__1876, 
        SYNOPSYS_UNCONNECTED__1877, N65160, N65159, N65158, N65157, N65156, 
        N65155}) );
  hamming_N16000_CC2_DW01_add_316 add_2982_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61025, N61024, N61023, N61022, 
        N61021}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61038, 
        N61037, N61036, N61035, N61034}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1878, SYNOPSYS_UNCONNECTED__1879, 
        SYNOPSYS_UNCONNECTED__1880, SYNOPSYS_UNCONNECTED__1881, 
        SYNOPSYS_UNCONNECTED__1882, SYNOPSYS_UNCONNECTED__1883, 
        SYNOPSYS_UNCONNECTED__1884, N65147, N65146, N65145, N65144, N65143, 
        N65142}) );
  hamming_N16000_CC2_DW01_add_317 add_2983_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60999, N60998, N60997, N60996, 
        N60995}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61012, 
        N61011, N61010, N61009, N61008}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1885, SYNOPSYS_UNCONNECTED__1886, 
        SYNOPSYS_UNCONNECTED__1887, SYNOPSYS_UNCONNECTED__1888, 
        SYNOPSYS_UNCONNECTED__1889, SYNOPSYS_UNCONNECTED__1890, 
        SYNOPSYS_UNCONNECTED__1891, N65134, N65133, N65132, N65131, N65130, 
        N65129}) );
  hamming_N16000_CC2_DW01_add_318 add_2984_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60973, N60972, N60971, N60970, 
        N60969}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60986, 
        N60985, N60984, N60983, N60982}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1892, SYNOPSYS_UNCONNECTED__1893, 
        SYNOPSYS_UNCONNECTED__1894, SYNOPSYS_UNCONNECTED__1895, 
        SYNOPSYS_UNCONNECTED__1896, SYNOPSYS_UNCONNECTED__1897, 
        SYNOPSYS_UNCONNECTED__1898, N65121, N65120, N65119, N65118, N65117, 
        N65116}) );
  hamming_N16000_CC2_DW01_add_319 add_2985_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60947, N60946, N60945, N60944, 
        N60943}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60960, 
        N60959, N60958, N60957, N60956}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1899, SYNOPSYS_UNCONNECTED__1900, 
        SYNOPSYS_UNCONNECTED__1901, SYNOPSYS_UNCONNECTED__1902, 
        SYNOPSYS_UNCONNECTED__1903, SYNOPSYS_UNCONNECTED__1904, 
        SYNOPSYS_UNCONNECTED__1905, N65108, N65107, N65106, N65105, N65104, 
        N65103}) );
  hamming_N16000_CC2_DW01_add_320 add_2986_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60921, N60920, N60919, N60918, 
        N60917}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60934, 
        N60933, N60932, N60931, N60930}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1906, SYNOPSYS_UNCONNECTED__1907, 
        SYNOPSYS_UNCONNECTED__1908, SYNOPSYS_UNCONNECTED__1909, 
        SYNOPSYS_UNCONNECTED__1910, SYNOPSYS_UNCONNECTED__1911, 
        SYNOPSYS_UNCONNECTED__1912, N65095, N65094, N65093, N65092, N65091, 
        N65090}) );
  hamming_N16000_CC2_DW01_add_321 add_2987_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60895, N60894, N60893, N60892, 
        N60891}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60908, 
        N60907, N60906, N60905, N60904}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1913, SYNOPSYS_UNCONNECTED__1914, 
        SYNOPSYS_UNCONNECTED__1915, SYNOPSYS_UNCONNECTED__1916, 
        SYNOPSYS_UNCONNECTED__1917, SYNOPSYS_UNCONNECTED__1918, 
        SYNOPSYS_UNCONNECTED__1919, N65082, N65081, N65080, N65079, N65078, 
        N65077}) );
  hamming_N16000_CC2_DW01_add_322 add_2988_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60869, N60868, N60867, N60866, 
        N60865}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60882, 
        N60881, N60880, N60879, N60878}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1920, SYNOPSYS_UNCONNECTED__1921, 
        SYNOPSYS_UNCONNECTED__1922, SYNOPSYS_UNCONNECTED__1923, 
        SYNOPSYS_UNCONNECTED__1924, SYNOPSYS_UNCONNECTED__1925, 
        SYNOPSYS_UNCONNECTED__1926, N65069, N65068, N65067, N65066, N65065, 
        N65064}) );
  hamming_N16000_CC2_DW01_add_323 add_2989_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60843, N60842, N60841, N60840, 
        N60839}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60856, 
        N60855, N60854, N60853, N60852}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1927, SYNOPSYS_UNCONNECTED__1928, 
        SYNOPSYS_UNCONNECTED__1929, SYNOPSYS_UNCONNECTED__1930, 
        SYNOPSYS_UNCONNECTED__1931, SYNOPSYS_UNCONNECTED__1932, 
        SYNOPSYS_UNCONNECTED__1933, N65056, N65055, N65054, N65053, N65052, 
        N65051}) );
  hamming_N16000_CC2_DW01_add_324 add_2990_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60817, N60816, N60815, N60814, 
        N60813}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60830, 
        N60829, N60828, N60827, N60826}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1934, SYNOPSYS_UNCONNECTED__1935, 
        SYNOPSYS_UNCONNECTED__1936, SYNOPSYS_UNCONNECTED__1937, 
        SYNOPSYS_UNCONNECTED__1938, SYNOPSYS_UNCONNECTED__1939, 
        SYNOPSYS_UNCONNECTED__1940, N65043, N65042, N65041, N65040, N65039, 
        N65038}) );
  hamming_N16000_CC2_DW01_add_325 add_2991_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60791, N60790, N60789, N60788, 
        N60787}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60804, 
        N60803, N60802, N60801, N60800}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1941, SYNOPSYS_UNCONNECTED__1942, 
        SYNOPSYS_UNCONNECTED__1943, SYNOPSYS_UNCONNECTED__1944, 
        SYNOPSYS_UNCONNECTED__1945, SYNOPSYS_UNCONNECTED__1946, 
        SYNOPSYS_UNCONNECTED__1947, N65030, N65029, N65028, N65027, N65026, 
        N65025}) );
  hamming_N16000_CC2_DW01_add_326 add_2992_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60765, N60764, N60763, N60762, 
        N60761}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60778, 
        N60777, N60776, N60775, N60774}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1948, SYNOPSYS_UNCONNECTED__1949, 
        SYNOPSYS_UNCONNECTED__1950, SYNOPSYS_UNCONNECTED__1951, 
        SYNOPSYS_UNCONNECTED__1952, SYNOPSYS_UNCONNECTED__1953, 
        SYNOPSYS_UNCONNECTED__1954, N65017, N65016, N65015, N65014, N65013, 
        N65012}) );
  hamming_N16000_CC2_DW01_add_327 add_2993_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60739, N60738, N60737, N60736, 
        N60735}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60752, 
        N60751, N60750, N60749, N60748}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1955, SYNOPSYS_UNCONNECTED__1956, 
        SYNOPSYS_UNCONNECTED__1957, SYNOPSYS_UNCONNECTED__1958, 
        SYNOPSYS_UNCONNECTED__1959, SYNOPSYS_UNCONNECTED__1960, 
        SYNOPSYS_UNCONNECTED__1961, N65004, N65003, N65002, N65001, N65000, 
        N64999}) );
  hamming_N16000_CC2_DW01_add_328 add_2994_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60713, N60712, N60711, N60710, 
        N60709}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60726, 
        N60725, N60724, N60723, N60722}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1962, SYNOPSYS_UNCONNECTED__1963, 
        SYNOPSYS_UNCONNECTED__1964, SYNOPSYS_UNCONNECTED__1965, 
        SYNOPSYS_UNCONNECTED__1966, SYNOPSYS_UNCONNECTED__1967, 
        SYNOPSYS_UNCONNECTED__1968, N64991, N64990, N64989, N64988, N64987, 
        N64986}) );
  hamming_N16000_CC2_DW01_add_329 add_2995_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60687, N60686, N60685, N60684, 
        N60683}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60700, 
        N60699, N60698, N60697, N60696}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1969, SYNOPSYS_UNCONNECTED__1970, 
        SYNOPSYS_UNCONNECTED__1971, SYNOPSYS_UNCONNECTED__1972, 
        SYNOPSYS_UNCONNECTED__1973, SYNOPSYS_UNCONNECTED__1974, 
        SYNOPSYS_UNCONNECTED__1975, N64978, N64977, N64976, N64975, N64974, 
        N64973}) );
  hamming_N16000_CC2_DW01_add_330 add_2996_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60661, N60660, N60659, N60658, 
        N60657}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60674, 
        N60673, N60672, N60671, N60670}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1976, SYNOPSYS_UNCONNECTED__1977, 
        SYNOPSYS_UNCONNECTED__1978, SYNOPSYS_UNCONNECTED__1979, 
        SYNOPSYS_UNCONNECTED__1980, SYNOPSYS_UNCONNECTED__1981, 
        SYNOPSYS_UNCONNECTED__1982, N64965, N64964, N64963, N64962, N64961, 
        N64960}) );
  hamming_N16000_CC2_DW01_add_331 add_2997_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60635, N60634, N60633, N60632, 
        N60631}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60648, 
        N60647, N60646, N60645, N60644}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1983, SYNOPSYS_UNCONNECTED__1984, 
        SYNOPSYS_UNCONNECTED__1985, SYNOPSYS_UNCONNECTED__1986, 
        SYNOPSYS_UNCONNECTED__1987, SYNOPSYS_UNCONNECTED__1988, 
        SYNOPSYS_UNCONNECTED__1989, N64952, N64951, N64950, N64949, N64948, 
        N64947}) );
  hamming_N16000_CC2_DW01_add_332 add_2998_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60609, N60608, N60607, N60606, 
        N60605}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60622, 
        N60621, N60620, N60619, N60618}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1990, SYNOPSYS_UNCONNECTED__1991, 
        SYNOPSYS_UNCONNECTED__1992, SYNOPSYS_UNCONNECTED__1993, 
        SYNOPSYS_UNCONNECTED__1994, SYNOPSYS_UNCONNECTED__1995, 
        SYNOPSYS_UNCONNECTED__1996, N64939, N64938, N64937, N64936, N64935, 
        N64934}) );
  hamming_N16000_CC2_DW01_add_333 add_2999_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60582, N60581, N60580, 
        N60579}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60596, 
        N60595, N60594, N60593, N60592}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1997, SYNOPSYS_UNCONNECTED__1998, 
        SYNOPSYS_UNCONNECTED__1999, SYNOPSYS_UNCONNECTED__2000, 
        SYNOPSYS_UNCONNECTED__2001, SYNOPSYS_UNCONNECTED__2002, 
        SYNOPSYS_UNCONNECTED__2003, N64926, N64925, N64924, N64923, N64922, 
        N64921}) );
  NAND U13353 ( .A(n5354), .B(n5355), .Z(N64912) );
  NANDN U13354 ( .A(n5356), .B(n5357), .Z(n5355) );
  OR U13355 ( .A(n5358), .B(n5359), .Z(n5357) );
  NAND U13356 ( .A(n5358), .B(n5359), .Z(n5354) );
  XOR U13357 ( .A(n5358), .B(n5360), .Z(N64911) );
  XNOR U13358 ( .A(n5356), .B(n5359), .Z(n5360) );
  AND U13359 ( .A(n5361), .B(n5362), .Z(n5359) );
  NANDN U13360 ( .A(n5363), .B(n5364), .Z(n5362) );
  NANDN U13361 ( .A(n5365), .B(n5366), .Z(n5364) );
  NANDN U13362 ( .A(n5366), .B(n5365), .Z(n5361) );
  NAND U13363 ( .A(n5367), .B(n5368), .Z(n5356) );
  NANDN U13364 ( .A(n5369), .B(n5370), .Z(n5368) );
  OR U13365 ( .A(n5371), .B(n5372), .Z(n5370) );
  NAND U13366 ( .A(n5372), .B(n5371), .Z(n5367) );
  AND U13367 ( .A(n5373), .B(n5374), .Z(n5358) );
  NANDN U13368 ( .A(n5375), .B(n5376), .Z(n5374) );
  NANDN U13369 ( .A(n5377), .B(n5378), .Z(n5376) );
  NANDN U13370 ( .A(n5378), .B(n5377), .Z(n5373) );
  XOR U13371 ( .A(n5372), .B(n5379), .Z(N64910) );
  XOR U13372 ( .A(n5369), .B(n5371), .Z(n5379) );
  XNOR U13373 ( .A(n5365), .B(n5380), .Z(n5371) );
  XNOR U13374 ( .A(n5363), .B(n5366), .Z(n5380) );
  NAND U13375 ( .A(n5381), .B(n5382), .Z(n5366) );
  NAND U13376 ( .A(n5383), .B(n5384), .Z(n5382) );
  OR U13377 ( .A(n5385), .B(n5386), .Z(n5383) );
  NANDN U13378 ( .A(n5387), .B(n5385), .Z(n5381) );
  IV U13379 ( .A(n5386), .Z(n5387) );
  NAND U13380 ( .A(n5388), .B(n5389), .Z(n5363) );
  NAND U13381 ( .A(n5390), .B(n5391), .Z(n5389) );
  NANDN U13382 ( .A(n5392), .B(n5393), .Z(n5390) );
  NANDN U13383 ( .A(n5393), .B(n5392), .Z(n5388) );
  AND U13384 ( .A(n5394), .B(n5395), .Z(n5365) );
  NAND U13385 ( .A(n5396), .B(n5397), .Z(n5395) );
  OR U13386 ( .A(n5398), .B(n5399), .Z(n5396) );
  NANDN U13387 ( .A(n5400), .B(n5398), .Z(n5394) );
  NAND U13388 ( .A(n5401), .B(n5402), .Z(n5369) );
  NANDN U13389 ( .A(n5403), .B(n5404), .Z(n5402) );
  OR U13390 ( .A(n5405), .B(n5406), .Z(n5404) );
  NANDN U13391 ( .A(n5407), .B(n5405), .Z(n5401) );
  IV U13392 ( .A(n5406), .Z(n5407) );
  XNOR U13393 ( .A(n5377), .B(n5408), .Z(n5372) );
  XNOR U13394 ( .A(n5375), .B(n5378), .Z(n5408) );
  NAND U13395 ( .A(n5409), .B(n5410), .Z(n5378) );
  NAND U13396 ( .A(n5411), .B(n5412), .Z(n5410) );
  OR U13397 ( .A(n5413), .B(n5414), .Z(n5411) );
  NANDN U13398 ( .A(n5415), .B(n5413), .Z(n5409) );
  IV U13399 ( .A(n5414), .Z(n5415) );
  NAND U13400 ( .A(n5416), .B(n5417), .Z(n5375) );
  NAND U13401 ( .A(n5418), .B(n5419), .Z(n5417) );
  NANDN U13402 ( .A(n5420), .B(n5421), .Z(n5418) );
  NANDN U13403 ( .A(n5421), .B(n5420), .Z(n5416) );
  AND U13404 ( .A(n5422), .B(n5423), .Z(n5377) );
  NAND U13405 ( .A(n5424), .B(n5425), .Z(n5423) );
  OR U13406 ( .A(n5426), .B(n5427), .Z(n5424) );
  NANDN U13407 ( .A(n5428), .B(n5426), .Z(n5422) );
  XNOR U13408 ( .A(n5403), .B(n5429), .Z(N64909) );
  XOR U13409 ( .A(n5405), .B(n5406), .Z(n5429) );
  XNOR U13410 ( .A(n5419), .B(n5430), .Z(n5406) );
  XOR U13411 ( .A(n5420), .B(n5421), .Z(n5430) );
  XOR U13412 ( .A(n5426), .B(n5431), .Z(n5421) );
  XOR U13413 ( .A(n5425), .B(n5428), .Z(n5431) );
  IV U13414 ( .A(n5427), .Z(n5428) );
  NAND U13415 ( .A(n5432), .B(n5433), .Z(n5427) );
  OR U13416 ( .A(n5434), .B(n5435), .Z(n5433) );
  OR U13417 ( .A(n5436), .B(n5437), .Z(n5432) );
  NAND U13418 ( .A(n5438), .B(n5439), .Z(n5425) );
  OR U13419 ( .A(n5440), .B(n5441), .Z(n5439) );
  OR U13420 ( .A(n5442), .B(n5443), .Z(n5438) );
  NOR U13421 ( .A(n5444), .B(n5445), .Z(n5426) );
  ANDN U13422 ( .B(n5446), .A(n5447), .Z(n5420) );
  XNOR U13423 ( .A(n5413), .B(n5448), .Z(n5419) );
  XNOR U13424 ( .A(n5412), .B(n5414), .Z(n5448) );
  NAND U13425 ( .A(n5449), .B(n5450), .Z(n5414) );
  OR U13426 ( .A(n5451), .B(n5452), .Z(n5450) );
  OR U13427 ( .A(n5453), .B(n5454), .Z(n5449) );
  NAND U13428 ( .A(n5455), .B(n5456), .Z(n5412) );
  OR U13429 ( .A(n5457), .B(n5458), .Z(n5456) );
  OR U13430 ( .A(n5459), .B(n5460), .Z(n5455) );
  ANDN U13431 ( .B(n5461), .A(n5462), .Z(n5413) );
  IV U13432 ( .A(n5463), .Z(n5461) );
  ANDN U13433 ( .B(n5464), .A(n5465), .Z(n5405) );
  XOR U13434 ( .A(n5391), .B(n5466), .Z(n5403) );
  XOR U13435 ( .A(n5392), .B(n5393), .Z(n5466) );
  XOR U13436 ( .A(n5398), .B(n5467), .Z(n5393) );
  XOR U13437 ( .A(n5397), .B(n5400), .Z(n5467) );
  IV U13438 ( .A(n5399), .Z(n5400) );
  NAND U13439 ( .A(n5468), .B(n5469), .Z(n5399) );
  OR U13440 ( .A(n5470), .B(n5471), .Z(n5469) );
  OR U13441 ( .A(n5472), .B(n5473), .Z(n5468) );
  NAND U13442 ( .A(n5474), .B(n5475), .Z(n5397) );
  OR U13443 ( .A(n5476), .B(n5477), .Z(n5475) );
  OR U13444 ( .A(n5478), .B(n5479), .Z(n5474) );
  NOR U13445 ( .A(n5480), .B(n5481), .Z(n5398) );
  ANDN U13446 ( .B(n5482), .A(n5483), .Z(n5392) );
  IV U13447 ( .A(n5484), .Z(n5482) );
  XNOR U13448 ( .A(n5385), .B(n5485), .Z(n5391) );
  XNOR U13449 ( .A(n5384), .B(n5386), .Z(n5485) );
  NAND U13450 ( .A(n5486), .B(n5487), .Z(n5386) );
  OR U13451 ( .A(n5488), .B(n5489), .Z(n5487) );
  OR U13452 ( .A(n5490), .B(n5491), .Z(n5486) );
  NAND U13453 ( .A(n5492), .B(n5493), .Z(n5384) );
  OR U13454 ( .A(n5494), .B(n5495), .Z(n5493) );
  OR U13455 ( .A(n5496), .B(n5497), .Z(n5492) );
  ANDN U13456 ( .B(n5498), .A(n5499), .Z(n5385) );
  IV U13457 ( .A(n5500), .Z(n5498) );
  XNOR U13458 ( .A(n5465), .B(n5464), .Z(N64908) );
  XOR U13459 ( .A(n5484), .B(n5483), .Z(n5464) );
  XNOR U13460 ( .A(n5499), .B(n5500), .Z(n5483) );
  XNOR U13461 ( .A(n5494), .B(n5495), .Z(n5500) );
  XNOR U13462 ( .A(n5496), .B(n5497), .Z(n5495) );
  XNOR U13463 ( .A(y[7981]), .B(x[7981]), .Z(n5497) );
  XNOR U13464 ( .A(y[7982]), .B(x[7982]), .Z(n5496) );
  XNOR U13465 ( .A(y[7980]), .B(x[7980]), .Z(n5494) );
  XNOR U13466 ( .A(n5488), .B(n5489), .Z(n5499) );
  XNOR U13467 ( .A(y[7977]), .B(x[7977]), .Z(n5489) );
  XNOR U13468 ( .A(n5490), .B(n5491), .Z(n5488) );
  XNOR U13469 ( .A(y[7978]), .B(x[7978]), .Z(n5491) );
  XNOR U13470 ( .A(y[7979]), .B(x[7979]), .Z(n5490) );
  XNOR U13471 ( .A(n5481), .B(n5480), .Z(n5484) );
  XNOR U13472 ( .A(n5476), .B(n5477), .Z(n5480) );
  XNOR U13473 ( .A(y[7974]), .B(x[7974]), .Z(n5477) );
  XNOR U13474 ( .A(n5478), .B(n5479), .Z(n5476) );
  XNOR U13475 ( .A(y[7975]), .B(x[7975]), .Z(n5479) );
  XNOR U13476 ( .A(y[7976]), .B(x[7976]), .Z(n5478) );
  XNOR U13477 ( .A(n5470), .B(n5471), .Z(n5481) );
  XNOR U13478 ( .A(y[7971]), .B(x[7971]), .Z(n5471) );
  XNOR U13479 ( .A(n5472), .B(n5473), .Z(n5470) );
  XNOR U13480 ( .A(y[7972]), .B(x[7972]), .Z(n5473) );
  XNOR U13481 ( .A(y[7973]), .B(x[7973]), .Z(n5472) );
  XOR U13482 ( .A(n5446), .B(n5447), .Z(n5465) );
  XNOR U13483 ( .A(n5462), .B(n5463), .Z(n5447) );
  XNOR U13484 ( .A(n5457), .B(n5458), .Z(n5463) );
  XNOR U13485 ( .A(n5459), .B(n5460), .Z(n5458) );
  XNOR U13486 ( .A(y[7969]), .B(x[7969]), .Z(n5460) );
  XNOR U13487 ( .A(y[7970]), .B(x[7970]), .Z(n5459) );
  XNOR U13488 ( .A(y[7968]), .B(x[7968]), .Z(n5457) );
  XNOR U13489 ( .A(n5451), .B(n5452), .Z(n5462) );
  XNOR U13490 ( .A(y[7965]), .B(x[7965]), .Z(n5452) );
  XNOR U13491 ( .A(n5453), .B(n5454), .Z(n5451) );
  XNOR U13492 ( .A(y[7966]), .B(x[7966]), .Z(n5454) );
  XNOR U13493 ( .A(y[7967]), .B(x[7967]), .Z(n5453) );
  XOR U13494 ( .A(n5445), .B(n5444), .Z(n5446) );
  XNOR U13495 ( .A(n5440), .B(n5441), .Z(n5444) );
  XNOR U13496 ( .A(y[7962]), .B(x[7962]), .Z(n5441) );
  XNOR U13497 ( .A(n5442), .B(n5443), .Z(n5440) );
  XNOR U13498 ( .A(y[7963]), .B(x[7963]), .Z(n5443) );
  XNOR U13499 ( .A(y[7964]), .B(x[7964]), .Z(n5442) );
  XNOR U13500 ( .A(n5434), .B(n5435), .Z(n5445) );
  XNOR U13501 ( .A(y[7959]), .B(x[7959]), .Z(n5435) );
  XNOR U13502 ( .A(n5436), .B(n5437), .Z(n5434) );
  XNOR U13503 ( .A(y[7960]), .B(x[7960]), .Z(n5437) );
  XNOR U13504 ( .A(y[7961]), .B(x[7961]), .Z(n5436) );
  NAND U13505 ( .A(n5501), .B(n5502), .Z(N64899) );
  NANDN U13506 ( .A(n5503), .B(n5504), .Z(n5502) );
  OR U13507 ( .A(n5505), .B(n5506), .Z(n5504) );
  NAND U13508 ( .A(n5505), .B(n5506), .Z(n5501) );
  XOR U13509 ( .A(n5505), .B(n5507), .Z(N64898) );
  XNOR U13510 ( .A(n5503), .B(n5506), .Z(n5507) );
  AND U13511 ( .A(n5508), .B(n5509), .Z(n5506) );
  NANDN U13512 ( .A(n5510), .B(n5511), .Z(n5509) );
  NANDN U13513 ( .A(n5512), .B(n5513), .Z(n5511) );
  NANDN U13514 ( .A(n5513), .B(n5512), .Z(n5508) );
  NAND U13515 ( .A(n5514), .B(n5515), .Z(n5503) );
  NANDN U13516 ( .A(n5516), .B(n5517), .Z(n5515) );
  OR U13517 ( .A(n5518), .B(n5519), .Z(n5517) );
  NAND U13518 ( .A(n5519), .B(n5518), .Z(n5514) );
  AND U13519 ( .A(n5520), .B(n5521), .Z(n5505) );
  NANDN U13520 ( .A(n5522), .B(n5523), .Z(n5521) );
  NANDN U13521 ( .A(n5524), .B(n5525), .Z(n5523) );
  NANDN U13522 ( .A(n5525), .B(n5524), .Z(n5520) );
  XOR U13523 ( .A(n5519), .B(n5526), .Z(N64897) );
  XOR U13524 ( .A(n5516), .B(n5518), .Z(n5526) );
  XNOR U13525 ( .A(n5512), .B(n5527), .Z(n5518) );
  XNOR U13526 ( .A(n5510), .B(n5513), .Z(n5527) );
  NAND U13527 ( .A(n5528), .B(n5529), .Z(n5513) );
  NAND U13528 ( .A(n5530), .B(n5531), .Z(n5529) );
  OR U13529 ( .A(n5532), .B(n5533), .Z(n5530) );
  NANDN U13530 ( .A(n5534), .B(n5532), .Z(n5528) );
  IV U13531 ( .A(n5533), .Z(n5534) );
  NAND U13532 ( .A(n5535), .B(n5536), .Z(n5510) );
  NAND U13533 ( .A(n5537), .B(n5538), .Z(n5536) );
  NANDN U13534 ( .A(n5539), .B(n5540), .Z(n5537) );
  NANDN U13535 ( .A(n5540), .B(n5539), .Z(n5535) );
  AND U13536 ( .A(n5541), .B(n5542), .Z(n5512) );
  NAND U13537 ( .A(n5543), .B(n5544), .Z(n5542) );
  OR U13538 ( .A(n5545), .B(n5546), .Z(n5543) );
  NANDN U13539 ( .A(n5547), .B(n5545), .Z(n5541) );
  NAND U13540 ( .A(n5548), .B(n5549), .Z(n5516) );
  NANDN U13541 ( .A(n5550), .B(n5551), .Z(n5549) );
  OR U13542 ( .A(n5552), .B(n5553), .Z(n5551) );
  NANDN U13543 ( .A(n5554), .B(n5552), .Z(n5548) );
  IV U13544 ( .A(n5553), .Z(n5554) );
  XNOR U13545 ( .A(n5524), .B(n5555), .Z(n5519) );
  XNOR U13546 ( .A(n5522), .B(n5525), .Z(n5555) );
  NAND U13547 ( .A(n5556), .B(n5557), .Z(n5525) );
  NAND U13548 ( .A(n5558), .B(n5559), .Z(n5557) );
  OR U13549 ( .A(n5560), .B(n5561), .Z(n5558) );
  NANDN U13550 ( .A(n5562), .B(n5560), .Z(n5556) );
  IV U13551 ( .A(n5561), .Z(n5562) );
  NAND U13552 ( .A(n5563), .B(n5564), .Z(n5522) );
  NAND U13553 ( .A(n5565), .B(n5566), .Z(n5564) );
  NANDN U13554 ( .A(n5567), .B(n5568), .Z(n5565) );
  NANDN U13555 ( .A(n5568), .B(n5567), .Z(n5563) );
  AND U13556 ( .A(n5569), .B(n5570), .Z(n5524) );
  NAND U13557 ( .A(n5571), .B(n5572), .Z(n5570) );
  OR U13558 ( .A(n5573), .B(n5574), .Z(n5571) );
  NANDN U13559 ( .A(n5575), .B(n5573), .Z(n5569) );
  XNOR U13560 ( .A(n5550), .B(n5576), .Z(N64896) );
  XOR U13561 ( .A(n5552), .B(n5553), .Z(n5576) );
  XNOR U13562 ( .A(n5566), .B(n5577), .Z(n5553) );
  XOR U13563 ( .A(n5567), .B(n5568), .Z(n5577) );
  XOR U13564 ( .A(n5573), .B(n5578), .Z(n5568) );
  XOR U13565 ( .A(n5572), .B(n5575), .Z(n5578) );
  IV U13566 ( .A(n5574), .Z(n5575) );
  NAND U13567 ( .A(n5579), .B(n5580), .Z(n5574) );
  OR U13568 ( .A(n5581), .B(n5582), .Z(n5580) );
  OR U13569 ( .A(n5583), .B(n5584), .Z(n5579) );
  NAND U13570 ( .A(n5585), .B(n5586), .Z(n5572) );
  OR U13571 ( .A(n5587), .B(n5588), .Z(n5586) );
  OR U13572 ( .A(n5589), .B(n5590), .Z(n5585) );
  NOR U13573 ( .A(n5591), .B(n5592), .Z(n5573) );
  ANDN U13574 ( .B(n5593), .A(n5594), .Z(n5567) );
  XNOR U13575 ( .A(n5560), .B(n5595), .Z(n5566) );
  XNOR U13576 ( .A(n5559), .B(n5561), .Z(n5595) );
  NAND U13577 ( .A(n5596), .B(n5597), .Z(n5561) );
  OR U13578 ( .A(n5598), .B(n5599), .Z(n5597) );
  OR U13579 ( .A(n5600), .B(n5601), .Z(n5596) );
  NAND U13580 ( .A(n5602), .B(n5603), .Z(n5559) );
  OR U13581 ( .A(n5604), .B(n5605), .Z(n5603) );
  OR U13582 ( .A(n5606), .B(n5607), .Z(n5602) );
  ANDN U13583 ( .B(n5608), .A(n5609), .Z(n5560) );
  IV U13584 ( .A(n5610), .Z(n5608) );
  ANDN U13585 ( .B(n5611), .A(n5612), .Z(n5552) );
  XOR U13586 ( .A(n5538), .B(n5613), .Z(n5550) );
  XOR U13587 ( .A(n5539), .B(n5540), .Z(n5613) );
  XOR U13588 ( .A(n5545), .B(n5614), .Z(n5540) );
  XOR U13589 ( .A(n5544), .B(n5547), .Z(n5614) );
  IV U13590 ( .A(n5546), .Z(n5547) );
  NAND U13591 ( .A(n5615), .B(n5616), .Z(n5546) );
  OR U13592 ( .A(n5617), .B(n5618), .Z(n5616) );
  OR U13593 ( .A(n5619), .B(n5620), .Z(n5615) );
  NAND U13594 ( .A(n5621), .B(n5622), .Z(n5544) );
  OR U13595 ( .A(n5623), .B(n5624), .Z(n5622) );
  OR U13596 ( .A(n5625), .B(n5626), .Z(n5621) );
  NOR U13597 ( .A(n5627), .B(n5628), .Z(n5545) );
  ANDN U13598 ( .B(n5629), .A(n5630), .Z(n5539) );
  IV U13599 ( .A(n5631), .Z(n5629) );
  XNOR U13600 ( .A(n5532), .B(n5632), .Z(n5538) );
  XNOR U13601 ( .A(n5531), .B(n5533), .Z(n5632) );
  NAND U13602 ( .A(n5633), .B(n5634), .Z(n5533) );
  OR U13603 ( .A(n5635), .B(n5636), .Z(n5634) );
  OR U13604 ( .A(n5637), .B(n5638), .Z(n5633) );
  NAND U13605 ( .A(n5639), .B(n5640), .Z(n5531) );
  OR U13606 ( .A(n5641), .B(n5642), .Z(n5640) );
  OR U13607 ( .A(n5643), .B(n5644), .Z(n5639) );
  ANDN U13608 ( .B(n5645), .A(n5646), .Z(n5532) );
  IV U13609 ( .A(n5647), .Z(n5645) );
  XNOR U13610 ( .A(n5612), .B(n5611), .Z(N64895) );
  XOR U13611 ( .A(n5631), .B(n5630), .Z(n5611) );
  XNOR U13612 ( .A(n5646), .B(n5647), .Z(n5630) );
  XNOR U13613 ( .A(n5641), .B(n5642), .Z(n5647) );
  XNOR U13614 ( .A(n5643), .B(n5644), .Z(n5642) );
  XNOR U13615 ( .A(y[7957]), .B(x[7957]), .Z(n5644) );
  XNOR U13616 ( .A(y[7958]), .B(x[7958]), .Z(n5643) );
  XNOR U13617 ( .A(y[7956]), .B(x[7956]), .Z(n5641) );
  XNOR U13618 ( .A(n5635), .B(n5636), .Z(n5646) );
  XNOR U13619 ( .A(y[7953]), .B(x[7953]), .Z(n5636) );
  XNOR U13620 ( .A(n5637), .B(n5638), .Z(n5635) );
  XNOR U13621 ( .A(y[7954]), .B(x[7954]), .Z(n5638) );
  XNOR U13622 ( .A(y[7955]), .B(x[7955]), .Z(n5637) );
  XNOR U13623 ( .A(n5628), .B(n5627), .Z(n5631) );
  XNOR U13624 ( .A(n5623), .B(n5624), .Z(n5627) );
  XNOR U13625 ( .A(y[7950]), .B(x[7950]), .Z(n5624) );
  XNOR U13626 ( .A(n5625), .B(n5626), .Z(n5623) );
  XNOR U13627 ( .A(y[7951]), .B(x[7951]), .Z(n5626) );
  XNOR U13628 ( .A(y[7952]), .B(x[7952]), .Z(n5625) );
  XNOR U13629 ( .A(n5617), .B(n5618), .Z(n5628) );
  XNOR U13630 ( .A(y[7947]), .B(x[7947]), .Z(n5618) );
  XNOR U13631 ( .A(n5619), .B(n5620), .Z(n5617) );
  XNOR U13632 ( .A(y[7948]), .B(x[7948]), .Z(n5620) );
  XNOR U13633 ( .A(y[7949]), .B(x[7949]), .Z(n5619) );
  XOR U13634 ( .A(n5593), .B(n5594), .Z(n5612) );
  XNOR U13635 ( .A(n5609), .B(n5610), .Z(n5594) );
  XNOR U13636 ( .A(n5604), .B(n5605), .Z(n5610) );
  XNOR U13637 ( .A(n5606), .B(n5607), .Z(n5605) );
  XNOR U13638 ( .A(y[7945]), .B(x[7945]), .Z(n5607) );
  XNOR U13639 ( .A(y[7946]), .B(x[7946]), .Z(n5606) );
  XNOR U13640 ( .A(y[7944]), .B(x[7944]), .Z(n5604) );
  XNOR U13641 ( .A(n5598), .B(n5599), .Z(n5609) );
  XNOR U13642 ( .A(y[7941]), .B(x[7941]), .Z(n5599) );
  XNOR U13643 ( .A(n5600), .B(n5601), .Z(n5598) );
  XNOR U13644 ( .A(y[7942]), .B(x[7942]), .Z(n5601) );
  XNOR U13645 ( .A(y[7943]), .B(x[7943]), .Z(n5600) );
  XOR U13646 ( .A(n5592), .B(n5591), .Z(n5593) );
  XNOR U13647 ( .A(n5587), .B(n5588), .Z(n5591) );
  XNOR U13648 ( .A(y[7938]), .B(x[7938]), .Z(n5588) );
  XNOR U13649 ( .A(n5589), .B(n5590), .Z(n5587) );
  XNOR U13650 ( .A(y[7939]), .B(x[7939]), .Z(n5590) );
  XNOR U13651 ( .A(y[7940]), .B(x[7940]), .Z(n5589) );
  XNOR U13652 ( .A(n5581), .B(n5582), .Z(n5592) );
  XNOR U13653 ( .A(y[7935]), .B(x[7935]), .Z(n5582) );
  XNOR U13654 ( .A(n5583), .B(n5584), .Z(n5581) );
  XNOR U13655 ( .A(y[7936]), .B(x[7936]), .Z(n5584) );
  XNOR U13656 ( .A(y[7937]), .B(x[7937]), .Z(n5583) );
  NAND U13657 ( .A(n5648), .B(n5649), .Z(N64886) );
  NANDN U13658 ( .A(n5650), .B(n5651), .Z(n5649) );
  OR U13659 ( .A(n5652), .B(n5653), .Z(n5651) );
  NAND U13660 ( .A(n5652), .B(n5653), .Z(n5648) );
  XOR U13661 ( .A(n5652), .B(n5654), .Z(N64885) );
  XNOR U13662 ( .A(n5650), .B(n5653), .Z(n5654) );
  AND U13663 ( .A(n5655), .B(n5656), .Z(n5653) );
  NANDN U13664 ( .A(n5657), .B(n5658), .Z(n5656) );
  NANDN U13665 ( .A(n5659), .B(n5660), .Z(n5658) );
  NANDN U13666 ( .A(n5660), .B(n5659), .Z(n5655) );
  NAND U13667 ( .A(n5661), .B(n5662), .Z(n5650) );
  NANDN U13668 ( .A(n5663), .B(n5664), .Z(n5662) );
  OR U13669 ( .A(n5665), .B(n5666), .Z(n5664) );
  NAND U13670 ( .A(n5666), .B(n5665), .Z(n5661) );
  AND U13671 ( .A(n5667), .B(n5668), .Z(n5652) );
  NANDN U13672 ( .A(n5669), .B(n5670), .Z(n5668) );
  NANDN U13673 ( .A(n5671), .B(n5672), .Z(n5670) );
  NANDN U13674 ( .A(n5672), .B(n5671), .Z(n5667) );
  XOR U13675 ( .A(n5666), .B(n5673), .Z(N64884) );
  XOR U13676 ( .A(n5663), .B(n5665), .Z(n5673) );
  XNOR U13677 ( .A(n5659), .B(n5674), .Z(n5665) );
  XNOR U13678 ( .A(n5657), .B(n5660), .Z(n5674) );
  NAND U13679 ( .A(n5675), .B(n5676), .Z(n5660) );
  NAND U13680 ( .A(n5677), .B(n5678), .Z(n5676) );
  OR U13681 ( .A(n5679), .B(n5680), .Z(n5677) );
  NANDN U13682 ( .A(n5681), .B(n5679), .Z(n5675) );
  IV U13683 ( .A(n5680), .Z(n5681) );
  NAND U13684 ( .A(n5682), .B(n5683), .Z(n5657) );
  NAND U13685 ( .A(n5684), .B(n5685), .Z(n5683) );
  NANDN U13686 ( .A(n5686), .B(n5687), .Z(n5684) );
  NANDN U13687 ( .A(n5687), .B(n5686), .Z(n5682) );
  AND U13688 ( .A(n5688), .B(n5689), .Z(n5659) );
  NAND U13689 ( .A(n5690), .B(n5691), .Z(n5689) );
  OR U13690 ( .A(n5692), .B(n5693), .Z(n5690) );
  NANDN U13691 ( .A(n5694), .B(n5692), .Z(n5688) );
  NAND U13692 ( .A(n5695), .B(n5696), .Z(n5663) );
  NANDN U13693 ( .A(n5697), .B(n5698), .Z(n5696) );
  OR U13694 ( .A(n5699), .B(n5700), .Z(n5698) );
  NANDN U13695 ( .A(n5701), .B(n5699), .Z(n5695) );
  IV U13696 ( .A(n5700), .Z(n5701) );
  XNOR U13697 ( .A(n5671), .B(n5702), .Z(n5666) );
  XNOR U13698 ( .A(n5669), .B(n5672), .Z(n5702) );
  NAND U13699 ( .A(n5703), .B(n5704), .Z(n5672) );
  NAND U13700 ( .A(n5705), .B(n5706), .Z(n5704) );
  OR U13701 ( .A(n5707), .B(n5708), .Z(n5705) );
  NANDN U13702 ( .A(n5709), .B(n5707), .Z(n5703) );
  IV U13703 ( .A(n5708), .Z(n5709) );
  NAND U13704 ( .A(n5710), .B(n5711), .Z(n5669) );
  NAND U13705 ( .A(n5712), .B(n5713), .Z(n5711) );
  NANDN U13706 ( .A(n5714), .B(n5715), .Z(n5712) );
  NANDN U13707 ( .A(n5715), .B(n5714), .Z(n5710) );
  AND U13708 ( .A(n5716), .B(n5717), .Z(n5671) );
  NAND U13709 ( .A(n5718), .B(n5719), .Z(n5717) );
  OR U13710 ( .A(n5720), .B(n5721), .Z(n5718) );
  NANDN U13711 ( .A(n5722), .B(n5720), .Z(n5716) );
  XNOR U13712 ( .A(n5697), .B(n5723), .Z(N64883) );
  XOR U13713 ( .A(n5699), .B(n5700), .Z(n5723) );
  XNOR U13714 ( .A(n5713), .B(n5724), .Z(n5700) );
  XOR U13715 ( .A(n5714), .B(n5715), .Z(n5724) );
  XOR U13716 ( .A(n5720), .B(n5725), .Z(n5715) );
  XOR U13717 ( .A(n5719), .B(n5722), .Z(n5725) );
  IV U13718 ( .A(n5721), .Z(n5722) );
  NAND U13719 ( .A(n5726), .B(n5727), .Z(n5721) );
  OR U13720 ( .A(n5728), .B(n5729), .Z(n5727) );
  OR U13721 ( .A(n5730), .B(n5731), .Z(n5726) );
  NAND U13722 ( .A(n5732), .B(n5733), .Z(n5719) );
  OR U13723 ( .A(n5734), .B(n5735), .Z(n5733) );
  OR U13724 ( .A(n5736), .B(n5737), .Z(n5732) );
  NOR U13725 ( .A(n5738), .B(n5739), .Z(n5720) );
  ANDN U13726 ( .B(n5740), .A(n5741), .Z(n5714) );
  XNOR U13727 ( .A(n5707), .B(n5742), .Z(n5713) );
  XNOR U13728 ( .A(n5706), .B(n5708), .Z(n5742) );
  NAND U13729 ( .A(n5743), .B(n5744), .Z(n5708) );
  OR U13730 ( .A(n5745), .B(n5746), .Z(n5744) );
  OR U13731 ( .A(n5747), .B(n5748), .Z(n5743) );
  NAND U13732 ( .A(n5749), .B(n5750), .Z(n5706) );
  OR U13733 ( .A(n5751), .B(n5752), .Z(n5750) );
  OR U13734 ( .A(n5753), .B(n5754), .Z(n5749) );
  ANDN U13735 ( .B(n5755), .A(n5756), .Z(n5707) );
  IV U13736 ( .A(n5757), .Z(n5755) );
  ANDN U13737 ( .B(n5758), .A(n5759), .Z(n5699) );
  XOR U13738 ( .A(n5685), .B(n5760), .Z(n5697) );
  XOR U13739 ( .A(n5686), .B(n5687), .Z(n5760) );
  XOR U13740 ( .A(n5692), .B(n5761), .Z(n5687) );
  XOR U13741 ( .A(n5691), .B(n5694), .Z(n5761) );
  IV U13742 ( .A(n5693), .Z(n5694) );
  NAND U13743 ( .A(n5762), .B(n5763), .Z(n5693) );
  OR U13744 ( .A(n5764), .B(n5765), .Z(n5763) );
  OR U13745 ( .A(n5766), .B(n5767), .Z(n5762) );
  NAND U13746 ( .A(n5768), .B(n5769), .Z(n5691) );
  OR U13747 ( .A(n5770), .B(n5771), .Z(n5769) );
  OR U13748 ( .A(n5772), .B(n5773), .Z(n5768) );
  NOR U13749 ( .A(n5774), .B(n5775), .Z(n5692) );
  ANDN U13750 ( .B(n5776), .A(n5777), .Z(n5686) );
  IV U13751 ( .A(n5778), .Z(n5776) );
  XNOR U13752 ( .A(n5679), .B(n5779), .Z(n5685) );
  XNOR U13753 ( .A(n5678), .B(n5680), .Z(n5779) );
  NAND U13754 ( .A(n5780), .B(n5781), .Z(n5680) );
  OR U13755 ( .A(n5782), .B(n5783), .Z(n5781) );
  OR U13756 ( .A(n5784), .B(n5785), .Z(n5780) );
  NAND U13757 ( .A(n5786), .B(n5787), .Z(n5678) );
  OR U13758 ( .A(n5788), .B(n5789), .Z(n5787) );
  OR U13759 ( .A(n5790), .B(n5791), .Z(n5786) );
  ANDN U13760 ( .B(n5792), .A(n5793), .Z(n5679) );
  IV U13761 ( .A(n5794), .Z(n5792) );
  XNOR U13762 ( .A(n5759), .B(n5758), .Z(N64882) );
  XOR U13763 ( .A(n5778), .B(n5777), .Z(n5758) );
  XNOR U13764 ( .A(n5793), .B(n5794), .Z(n5777) );
  XNOR U13765 ( .A(n5788), .B(n5789), .Z(n5794) );
  XNOR U13766 ( .A(n5790), .B(n5791), .Z(n5789) );
  XNOR U13767 ( .A(y[7933]), .B(x[7933]), .Z(n5791) );
  XNOR U13768 ( .A(y[7934]), .B(x[7934]), .Z(n5790) );
  XNOR U13769 ( .A(y[7932]), .B(x[7932]), .Z(n5788) );
  XNOR U13770 ( .A(n5782), .B(n5783), .Z(n5793) );
  XNOR U13771 ( .A(y[7929]), .B(x[7929]), .Z(n5783) );
  XNOR U13772 ( .A(n5784), .B(n5785), .Z(n5782) );
  XNOR U13773 ( .A(y[7930]), .B(x[7930]), .Z(n5785) );
  XNOR U13774 ( .A(y[7931]), .B(x[7931]), .Z(n5784) );
  XNOR U13775 ( .A(n5775), .B(n5774), .Z(n5778) );
  XNOR U13776 ( .A(n5770), .B(n5771), .Z(n5774) );
  XNOR U13777 ( .A(y[7926]), .B(x[7926]), .Z(n5771) );
  XNOR U13778 ( .A(n5772), .B(n5773), .Z(n5770) );
  XNOR U13779 ( .A(y[7927]), .B(x[7927]), .Z(n5773) );
  XNOR U13780 ( .A(y[7928]), .B(x[7928]), .Z(n5772) );
  XNOR U13781 ( .A(n5764), .B(n5765), .Z(n5775) );
  XNOR U13782 ( .A(y[7923]), .B(x[7923]), .Z(n5765) );
  XNOR U13783 ( .A(n5766), .B(n5767), .Z(n5764) );
  XNOR U13784 ( .A(y[7924]), .B(x[7924]), .Z(n5767) );
  XNOR U13785 ( .A(y[7925]), .B(x[7925]), .Z(n5766) );
  XOR U13786 ( .A(n5740), .B(n5741), .Z(n5759) );
  XNOR U13787 ( .A(n5756), .B(n5757), .Z(n5741) );
  XNOR U13788 ( .A(n5751), .B(n5752), .Z(n5757) );
  XNOR U13789 ( .A(n5753), .B(n5754), .Z(n5752) );
  XNOR U13790 ( .A(y[7921]), .B(x[7921]), .Z(n5754) );
  XNOR U13791 ( .A(y[7922]), .B(x[7922]), .Z(n5753) );
  XNOR U13792 ( .A(y[7920]), .B(x[7920]), .Z(n5751) );
  XNOR U13793 ( .A(n5745), .B(n5746), .Z(n5756) );
  XNOR U13794 ( .A(y[7917]), .B(x[7917]), .Z(n5746) );
  XNOR U13795 ( .A(n5747), .B(n5748), .Z(n5745) );
  XNOR U13796 ( .A(y[7918]), .B(x[7918]), .Z(n5748) );
  XNOR U13797 ( .A(y[7919]), .B(x[7919]), .Z(n5747) );
  XOR U13798 ( .A(n5739), .B(n5738), .Z(n5740) );
  XNOR U13799 ( .A(n5734), .B(n5735), .Z(n5738) );
  XNOR U13800 ( .A(y[7914]), .B(x[7914]), .Z(n5735) );
  XNOR U13801 ( .A(n5736), .B(n5737), .Z(n5734) );
  XNOR U13802 ( .A(y[7915]), .B(x[7915]), .Z(n5737) );
  XNOR U13803 ( .A(y[7916]), .B(x[7916]), .Z(n5736) );
  XNOR U13804 ( .A(n5728), .B(n5729), .Z(n5739) );
  XNOR U13805 ( .A(y[7911]), .B(x[7911]), .Z(n5729) );
  XNOR U13806 ( .A(n5730), .B(n5731), .Z(n5728) );
  XNOR U13807 ( .A(y[7912]), .B(x[7912]), .Z(n5731) );
  XNOR U13808 ( .A(y[7913]), .B(x[7913]), .Z(n5730) );
  NAND U13809 ( .A(n5795), .B(n5796), .Z(N64873) );
  NANDN U13810 ( .A(n5797), .B(n5798), .Z(n5796) );
  OR U13811 ( .A(n5799), .B(n5800), .Z(n5798) );
  NAND U13812 ( .A(n5799), .B(n5800), .Z(n5795) );
  XOR U13813 ( .A(n5799), .B(n5801), .Z(N64872) );
  XNOR U13814 ( .A(n5797), .B(n5800), .Z(n5801) );
  AND U13815 ( .A(n5802), .B(n5803), .Z(n5800) );
  NANDN U13816 ( .A(n5804), .B(n5805), .Z(n5803) );
  NANDN U13817 ( .A(n5806), .B(n5807), .Z(n5805) );
  NANDN U13818 ( .A(n5807), .B(n5806), .Z(n5802) );
  NAND U13819 ( .A(n5808), .B(n5809), .Z(n5797) );
  NANDN U13820 ( .A(n5810), .B(n5811), .Z(n5809) );
  OR U13821 ( .A(n5812), .B(n5813), .Z(n5811) );
  NAND U13822 ( .A(n5813), .B(n5812), .Z(n5808) );
  AND U13823 ( .A(n5814), .B(n5815), .Z(n5799) );
  NANDN U13824 ( .A(n5816), .B(n5817), .Z(n5815) );
  NANDN U13825 ( .A(n5818), .B(n5819), .Z(n5817) );
  NANDN U13826 ( .A(n5819), .B(n5818), .Z(n5814) );
  XOR U13827 ( .A(n5813), .B(n5820), .Z(N64871) );
  XOR U13828 ( .A(n5810), .B(n5812), .Z(n5820) );
  XNOR U13829 ( .A(n5806), .B(n5821), .Z(n5812) );
  XNOR U13830 ( .A(n5804), .B(n5807), .Z(n5821) );
  NAND U13831 ( .A(n5822), .B(n5823), .Z(n5807) );
  NAND U13832 ( .A(n5824), .B(n5825), .Z(n5823) );
  OR U13833 ( .A(n5826), .B(n5827), .Z(n5824) );
  NANDN U13834 ( .A(n5828), .B(n5826), .Z(n5822) );
  IV U13835 ( .A(n5827), .Z(n5828) );
  NAND U13836 ( .A(n5829), .B(n5830), .Z(n5804) );
  NAND U13837 ( .A(n5831), .B(n5832), .Z(n5830) );
  NANDN U13838 ( .A(n5833), .B(n5834), .Z(n5831) );
  NANDN U13839 ( .A(n5834), .B(n5833), .Z(n5829) );
  AND U13840 ( .A(n5835), .B(n5836), .Z(n5806) );
  NAND U13841 ( .A(n5837), .B(n5838), .Z(n5836) );
  OR U13842 ( .A(n5839), .B(n5840), .Z(n5837) );
  NANDN U13843 ( .A(n5841), .B(n5839), .Z(n5835) );
  NAND U13844 ( .A(n5842), .B(n5843), .Z(n5810) );
  NANDN U13845 ( .A(n5844), .B(n5845), .Z(n5843) );
  OR U13846 ( .A(n5846), .B(n5847), .Z(n5845) );
  NANDN U13847 ( .A(n5848), .B(n5846), .Z(n5842) );
  IV U13848 ( .A(n5847), .Z(n5848) );
  XNOR U13849 ( .A(n5818), .B(n5849), .Z(n5813) );
  XNOR U13850 ( .A(n5816), .B(n5819), .Z(n5849) );
  NAND U13851 ( .A(n5850), .B(n5851), .Z(n5819) );
  NAND U13852 ( .A(n5852), .B(n5853), .Z(n5851) );
  OR U13853 ( .A(n5854), .B(n5855), .Z(n5852) );
  NANDN U13854 ( .A(n5856), .B(n5854), .Z(n5850) );
  IV U13855 ( .A(n5855), .Z(n5856) );
  NAND U13856 ( .A(n5857), .B(n5858), .Z(n5816) );
  NAND U13857 ( .A(n5859), .B(n5860), .Z(n5858) );
  NANDN U13858 ( .A(n5861), .B(n5862), .Z(n5859) );
  NANDN U13859 ( .A(n5862), .B(n5861), .Z(n5857) );
  AND U13860 ( .A(n5863), .B(n5864), .Z(n5818) );
  NAND U13861 ( .A(n5865), .B(n5866), .Z(n5864) );
  OR U13862 ( .A(n5867), .B(n5868), .Z(n5865) );
  NANDN U13863 ( .A(n5869), .B(n5867), .Z(n5863) );
  XNOR U13864 ( .A(n5844), .B(n5870), .Z(N64870) );
  XOR U13865 ( .A(n5846), .B(n5847), .Z(n5870) );
  XNOR U13866 ( .A(n5860), .B(n5871), .Z(n5847) );
  XOR U13867 ( .A(n5861), .B(n5862), .Z(n5871) );
  XOR U13868 ( .A(n5867), .B(n5872), .Z(n5862) );
  XOR U13869 ( .A(n5866), .B(n5869), .Z(n5872) );
  IV U13870 ( .A(n5868), .Z(n5869) );
  NAND U13871 ( .A(n5873), .B(n5874), .Z(n5868) );
  OR U13872 ( .A(n5875), .B(n5876), .Z(n5874) );
  OR U13873 ( .A(n5877), .B(n5878), .Z(n5873) );
  NAND U13874 ( .A(n5879), .B(n5880), .Z(n5866) );
  OR U13875 ( .A(n5881), .B(n5882), .Z(n5880) );
  OR U13876 ( .A(n5883), .B(n5884), .Z(n5879) );
  NOR U13877 ( .A(n5885), .B(n5886), .Z(n5867) );
  ANDN U13878 ( .B(n5887), .A(n5888), .Z(n5861) );
  XNOR U13879 ( .A(n5854), .B(n5889), .Z(n5860) );
  XNOR U13880 ( .A(n5853), .B(n5855), .Z(n5889) );
  NAND U13881 ( .A(n5890), .B(n5891), .Z(n5855) );
  OR U13882 ( .A(n5892), .B(n5893), .Z(n5891) );
  OR U13883 ( .A(n5894), .B(n5895), .Z(n5890) );
  NAND U13884 ( .A(n5896), .B(n5897), .Z(n5853) );
  OR U13885 ( .A(n5898), .B(n5899), .Z(n5897) );
  OR U13886 ( .A(n5900), .B(n5901), .Z(n5896) );
  ANDN U13887 ( .B(n5902), .A(n5903), .Z(n5854) );
  IV U13888 ( .A(n5904), .Z(n5902) );
  ANDN U13889 ( .B(n5905), .A(n5906), .Z(n5846) );
  XOR U13890 ( .A(n5832), .B(n5907), .Z(n5844) );
  XOR U13891 ( .A(n5833), .B(n5834), .Z(n5907) );
  XOR U13892 ( .A(n5839), .B(n5908), .Z(n5834) );
  XOR U13893 ( .A(n5838), .B(n5841), .Z(n5908) );
  IV U13894 ( .A(n5840), .Z(n5841) );
  NAND U13895 ( .A(n5909), .B(n5910), .Z(n5840) );
  OR U13896 ( .A(n5911), .B(n5912), .Z(n5910) );
  OR U13897 ( .A(n5913), .B(n5914), .Z(n5909) );
  NAND U13898 ( .A(n5915), .B(n5916), .Z(n5838) );
  OR U13899 ( .A(n5917), .B(n5918), .Z(n5916) );
  OR U13900 ( .A(n5919), .B(n5920), .Z(n5915) );
  NOR U13901 ( .A(n5921), .B(n5922), .Z(n5839) );
  ANDN U13902 ( .B(n5923), .A(n5924), .Z(n5833) );
  IV U13903 ( .A(n5925), .Z(n5923) );
  XNOR U13904 ( .A(n5826), .B(n5926), .Z(n5832) );
  XNOR U13905 ( .A(n5825), .B(n5827), .Z(n5926) );
  NAND U13906 ( .A(n5927), .B(n5928), .Z(n5827) );
  OR U13907 ( .A(n5929), .B(n5930), .Z(n5928) );
  OR U13908 ( .A(n5931), .B(n5932), .Z(n5927) );
  NAND U13909 ( .A(n5933), .B(n5934), .Z(n5825) );
  OR U13910 ( .A(n5935), .B(n5936), .Z(n5934) );
  OR U13911 ( .A(n5937), .B(n5938), .Z(n5933) );
  ANDN U13912 ( .B(n5939), .A(n5940), .Z(n5826) );
  IV U13913 ( .A(n5941), .Z(n5939) );
  XNOR U13914 ( .A(n5906), .B(n5905), .Z(N64869) );
  XOR U13915 ( .A(n5925), .B(n5924), .Z(n5905) );
  XNOR U13916 ( .A(n5940), .B(n5941), .Z(n5924) );
  XNOR U13917 ( .A(n5935), .B(n5936), .Z(n5941) );
  XNOR U13918 ( .A(n5937), .B(n5938), .Z(n5936) );
  XNOR U13919 ( .A(y[7909]), .B(x[7909]), .Z(n5938) );
  XNOR U13920 ( .A(y[7910]), .B(x[7910]), .Z(n5937) );
  XNOR U13921 ( .A(y[7908]), .B(x[7908]), .Z(n5935) );
  XNOR U13922 ( .A(n5929), .B(n5930), .Z(n5940) );
  XNOR U13923 ( .A(y[7905]), .B(x[7905]), .Z(n5930) );
  XNOR U13924 ( .A(n5931), .B(n5932), .Z(n5929) );
  XNOR U13925 ( .A(y[7906]), .B(x[7906]), .Z(n5932) );
  XNOR U13926 ( .A(y[7907]), .B(x[7907]), .Z(n5931) );
  XNOR U13927 ( .A(n5922), .B(n5921), .Z(n5925) );
  XNOR U13928 ( .A(n5917), .B(n5918), .Z(n5921) );
  XNOR U13929 ( .A(y[7902]), .B(x[7902]), .Z(n5918) );
  XNOR U13930 ( .A(n5919), .B(n5920), .Z(n5917) );
  XNOR U13931 ( .A(y[7903]), .B(x[7903]), .Z(n5920) );
  XNOR U13932 ( .A(y[7904]), .B(x[7904]), .Z(n5919) );
  XNOR U13933 ( .A(n5911), .B(n5912), .Z(n5922) );
  XNOR U13934 ( .A(y[7899]), .B(x[7899]), .Z(n5912) );
  XNOR U13935 ( .A(n5913), .B(n5914), .Z(n5911) );
  XNOR U13936 ( .A(y[7900]), .B(x[7900]), .Z(n5914) );
  XNOR U13937 ( .A(y[7901]), .B(x[7901]), .Z(n5913) );
  XOR U13938 ( .A(n5887), .B(n5888), .Z(n5906) );
  XNOR U13939 ( .A(n5903), .B(n5904), .Z(n5888) );
  XNOR U13940 ( .A(n5898), .B(n5899), .Z(n5904) );
  XNOR U13941 ( .A(n5900), .B(n5901), .Z(n5899) );
  XNOR U13942 ( .A(y[7897]), .B(x[7897]), .Z(n5901) );
  XNOR U13943 ( .A(y[7898]), .B(x[7898]), .Z(n5900) );
  XNOR U13944 ( .A(y[7896]), .B(x[7896]), .Z(n5898) );
  XNOR U13945 ( .A(n5892), .B(n5893), .Z(n5903) );
  XNOR U13946 ( .A(y[7893]), .B(x[7893]), .Z(n5893) );
  XNOR U13947 ( .A(n5894), .B(n5895), .Z(n5892) );
  XNOR U13948 ( .A(y[7894]), .B(x[7894]), .Z(n5895) );
  XNOR U13949 ( .A(y[7895]), .B(x[7895]), .Z(n5894) );
  XOR U13950 ( .A(n5886), .B(n5885), .Z(n5887) );
  XNOR U13951 ( .A(n5881), .B(n5882), .Z(n5885) );
  XNOR U13952 ( .A(y[7890]), .B(x[7890]), .Z(n5882) );
  XNOR U13953 ( .A(n5883), .B(n5884), .Z(n5881) );
  XNOR U13954 ( .A(y[7891]), .B(x[7891]), .Z(n5884) );
  XNOR U13955 ( .A(y[7892]), .B(x[7892]), .Z(n5883) );
  XNOR U13956 ( .A(n5875), .B(n5876), .Z(n5886) );
  XNOR U13957 ( .A(y[7887]), .B(x[7887]), .Z(n5876) );
  XNOR U13958 ( .A(n5877), .B(n5878), .Z(n5875) );
  XNOR U13959 ( .A(y[7888]), .B(x[7888]), .Z(n5878) );
  XNOR U13960 ( .A(y[7889]), .B(x[7889]), .Z(n5877) );
  NAND U13961 ( .A(n5942), .B(n5943), .Z(N64860) );
  NANDN U13962 ( .A(n5944), .B(n5945), .Z(n5943) );
  OR U13963 ( .A(n5946), .B(n5947), .Z(n5945) );
  NAND U13964 ( .A(n5946), .B(n5947), .Z(n5942) );
  XOR U13965 ( .A(n5946), .B(n5948), .Z(N64859) );
  XNOR U13966 ( .A(n5944), .B(n5947), .Z(n5948) );
  AND U13967 ( .A(n5949), .B(n5950), .Z(n5947) );
  NANDN U13968 ( .A(n5951), .B(n5952), .Z(n5950) );
  NANDN U13969 ( .A(n5953), .B(n5954), .Z(n5952) );
  NANDN U13970 ( .A(n5954), .B(n5953), .Z(n5949) );
  NAND U13971 ( .A(n5955), .B(n5956), .Z(n5944) );
  NANDN U13972 ( .A(n5957), .B(n5958), .Z(n5956) );
  OR U13973 ( .A(n5959), .B(n5960), .Z(n5958) );
  NAND U13974 ( .A(n5960), .B(n5959), .Z(n5955) );
  AND U13975 ( .A(n5961), .B(n5962), .Z(n5946) );
  NANDN U13976 ( .A(n5963), .B(n5964), .Z(n5962) );
  NANDN U13977 ( .A(n5965), .B(n5966), .Z(n5964) );
  NANDN U13978 ( .A(n5966), .B(n5965), .Z(n5961) );
  XOR U13979 ( .A(n5960), .B(n5967), .Z(N64858) );
  XOR U13980 ( .A(n5957), .B(n5959), .Z(n5967) );
  XNOR U13981 ( .A(n5953), .B(n5968), .Z(n5959) );
  XNOR U13982 ( .A(n5951), .B(n5954), .Z(n5968) );
  NAND U13983 ( .A(n5969), .B(n5970), .Z(n5954) );
  NAND U13984 ( .A(n5971), .B(n5972), .Z(n5970) );
  OR U13985 ( .A(n5973), .B(n5974), .Z(n5971) );
  NANDN U13986 ( .A(n5975), .B(n5973), .Z(n5969) );
  IV U13987 ( .A(n5974), .Z(n5975) );
  NAND U13988 ( .A(n5976), .B(n5977), .Z(n5951) );
  NAND U13989 ( .A(n5978), .B(n5979), .Z(n5977) );
  NANDN U13990 ( .A(n5980), .B(n5981), .Z(n5978) );
  NANDN U13991 ( .A(n5981), .B(n5980), .Z(n5976) );
  AND U13992 ( .A(n5982), .B(n5983), .Z(n5953) );
  NAND U13993 ( .A(n5984), .B(n5985), .Z(n5983) );
  OR U13994 ( .A(n5986), .B(n5987), .Z(n5984) );
  NANDN U13995 ( .A(n5988), .B(n5986), .Z(n5982) );
  NAND U13996 ( .A(n5989), .B(n5990), .Z(n5957) );
  NANDN U13997 ( .A(n5991), .B(n5992), .Z(n5990) );
  OR U13998 ( .A(n5993), .B(n5994), .Z(n5992) );
  NANDN U13999 ( .A(n5995), .B(n5993), .Z(n5989) );
  IV U14000 ( .A(n5994), .Z(n5995) );
  XNOR U14001 ( .A(n5965), .B(n5996), .Z(n5960) );
  XNOR U14002 ( .A(n5963), .B(n5966), .Z(n5996) );
  NAND U14003 ( .A(n5997), .B(n5998), .Z(n5966) );
  NAND U14004 ( .A(n5999), .B(n6000), .Z(n5998) );
  OR U14005 ( .A(n6001), .B(n6002), .Z(n5999) );
  NANDN U14006 ( .A(n6003), .B(n6001), .Z(n5997) );
  IV U14007 ( .A(n6002), .Z(n6003) );
  NAND U14008 ( .A(n6004), .B(n6005), .Z(n5963) );
  NAND U14009 ( .A(n6006), .B(n6007), .Z(n6005) );
  NANDN U14010 ( .A(n6008), .B(n6009), .Z(n6006) );
  NANDN U14011 ( .A(n6009), .B(n6008), .Z(n6004) );
  AND U14012 ( .A(n6010), .B(n6011), .Z(n5965) );
  NAND U14013 ( .A(n6012), .B(n6013), .Z(n6011) );
  OR U14014 ( .A(n6014), .B(n6015), .Z(n6012) );
  NANDN U14015 ( .A(n6016), .B(n6014), .Z(n6010) );
  XNOR U14016 ( .A(n5991), .B(n6017), .Z(N64857) );
  XOR U14017 ( .A(n5993), .B(n5994), .Z(n6017) );
  XNOR U14018 ( .A(n6007), .B(n6018), .Z(n5994) );
  XOR U14019 ( .A(n6008), .B(n6009), .Z(n6018) );
  XOR U14020 ( .A(n6014), .B(n6019), .Z(n6009) );
  XOR U14021 ( .A(n6013), .B(n6016), .Z(n6019) );
  IV U14022 ( .A(n6015), .Z(n6016) );
  NAND U14023 ( .A(n6020), .B(n6021), .Z(n6015) );
  OR U14024 ( .A(n6022), .B(n6023), .Z(n6021) );
  OR U14025 ( .A(n6024), .B(n6025), .Z(n6020) );
  NAND U14026 ( .A(n6026), .B(n6027), .Z(n6013) );
  OR U14027 ( .A(n6028), .B(n6029), .Z(n6027) );
  OR U14028 ( .A(n6030), .B(n6031), .Z(n6026) );
  NOR U14029 ( .A(n6032), .B(n6033), .Z(n6014) );
  ANDN U14030 ( .B(n6034), .A(n6035), .Z(n6008) );
  XNOR U14031 ( .A(n6001), .B(n6036), .Z(n6007) );
  XNOR U14032 ( .A(n6000), .B(n6002), .Z(n6036) );
  NAND U14033 ( .A(n6037), .B(n6038), .Z(n6002) );
  OR U14034 ( .A(n6039), .B(n6040), .Z(n6038) );
  OR U14035 ( .A(n6041), .B(n6042), .Z(n6037) );
  NAND U14036 ( .A(n6043), .B(n6044), .Z(n6000) );
  OR U14037 ( .A(n6045), .B(n6046), .Z(n6044) );
  OR U14038 ( .A(n6047), .B(n6048), .Z(n6043) );
  ANDN U14039 ( .B(n6049), .A(n6050), .Z(n6001) );
  IV U14040 ( .A(n6051), .Z(n6049) );
  ANDN U14041 ( .B(n6052), .A(n6053), .Z(n5993) );
  XOR U14042 ( .A(n5979), .B(n6054), .Z(n5991) );
  XOR U14043 ( .A(n5980), .B(n5981), .Z(n6054) );
  XOR U14044 ( .A(n5986), .B(n6055), .Z(n5981) );
  XOR U14045 ( .A(n5985), .B(n5988), .Z(n6055) );
  IV U14046 ( .A(n5987), .Z(n5988) );
  NAND U14047 ( .A(n6056), .B(n6057), .Z(n5987) );
  OR U14048 ( .A(n6058), .B(n6059), .Z(n6057) );
  OR U14049 ( .A(n6060), .B(n6061), .Z(n6056) );
  NAND U14050 ( .A(n6062), .B(n6063), .Z(n5985) );
  OR U14051 ( .A(n6064), .B(n6065), .Z(n6063) );
  OR U14052 ( .A(n6066), .B(n6067), .Z(n6062) );
  NOR U14053 ( .A(n6068), .B(n6069), .Z(n5986) );
  ANDN U14054 ( .B(n6070), .A(n6071), .Z(n5980) );
  IV U14055 ( .A(n6072), .Z(n6070) );
  XNOR U14056 ( .A(n5973), .B(n6073), .Z(n5979) );
  XNOR U14057 ( .A(n5972), .B(n5974), .Z(n6073) );
  NAND U14058 ( .A(n6074), .B(n6075), .Z(n5974) );
  OR U14059 ( .A(n6076), .B(n6077), .Z(n6075) );
  OR U14060 ( .A(n6078), .B(n6079), .Z(n6074) );
  NAND U14061 ( .A(n6080), .B(n6081), .Z(n5972) );
  OR U14062 ( .A(n6082), .B(n6083), .Z(n6081) );
  OR U14063 ( .A(n6084), .B(n6085), .Z(n6080) );
  ANDN U14064 ( .B(n6086), .A(n6087), .Z(n5973) );
  IV U14065 ( .A(n6088), .Z(n6086) );
  XNOR U14066 ( .A(n6053), .B(n6052), .Z(N64856) );
  XOR U14067 ( .A(n6072), .B(n6071), .Z(n6052) );
  XNOR U14068 ( .A(n6087), .B(n6088), .Z(n6071) );
  XNOR U14069 ( .A(n6082), .B(n6083), .Z(n6088) );
  XNOR U14070 ( .A(n6084), .B(n6085), .Z(n6083) );
  XNOR U14071 ( .A(y[7885]), .B(x[7885]), .Z(n6085) );
  XNOR U14072 ( .A(y[7886]), .B(x[7886]), .Z(n6084) );
  XNOR U14073 ( .A(y[7884]), .B(x[7884]), .Z(n6082) );
  XNOR U14074 ( .A(n6076), .B(n6077), .Z(n6087) );
  XNOR U14075 ( .A(y[7881]), .B(x[7881]), .Z(n6077) );
  XNOR U14076 ( .A(n6078), .B(n6079), .Z(n6076) );
  XNOR U14077 ( .A(y[7882]), .B(x[7882]), .Z(n6079) );
  XNOR U14078 ( .A(y[7883]), .B(x[7883]), .Z(n6078) );
  XNOR U14079 ( .A(n6069), .B(n6068), .Z(n6072) );
  XNOR U14080 ( .A(n6064), .B(n6065), .Z(n6068) );
  XNOR U14081 ( .A(y[7878]), .B(x[7878]), .Z(n6065) );
  XNOR U14082 ( .A(n6066), .B(n6067), .Z(n6064) );
  XNOR U14083 ( .A(y[7879]), .B(x[7879]), .Z(n6067) );
  XNOR U14084 ( .A(y[7880]), .B(x[7880]), .Z(n6066) );
  XNOR U14085 ( .A(n6058), .B(n6059), .Z(n6069) );
  XNOR U14086 ( .A(y[7875]), .B(x[7875]), .Z(n6059) );
  XNOR U14087 ( .A(n6060), .B(n6061), .Z(n6058) );
  XNOR U14088 ( .A(y[7876]), .B(x[7876]), .Z(n6061) );
  XNOR U14089 ( .A(y[7877]), .B(x[7877]), .Z(n6060) );
  XOR U14090 ( .A(n6034), .B(n6035), .Z(n6053) );
  XNOR U14091 ( .A(n6050), .B(n6051), .Z(n6035) );
  XNOR U14092 ( .A(n6045), .B(n6046), .Z(n6051) );
  XNOR U14093 ( .A(n6047), .B(n6048), .Z(n6046) );
  XNOR U14094 ( .A(y[7873]), .B(x[7873]), .Z(n6048) );
  XNOR U14095 ( .A(y[7874]), .B(x[7874]), .Z(n6047) );
  XNOR U14096 ( .A(y[7872]), .B(x[7872]), .Z(n6045) );
  XNOR U14097 ( .A(n6039), .B(n6040), .Z(n6050) );
  XNOR U14098 ( .A(y[7869]), .B(x[7869]), .Z(n6040) );
  XNOR U14099 ( .A(n6041), .B(n6042), .Z(n6039) );
  XNOR U14100 ( .A(y[7870]), .B(x[7870]), .Z(n6042) );
  XNOR U14101 ( .A(y[7871]), .B(x[7871]), .Z(n6041) );
  XOR U14102 ( .A(n6033), .B(n6032), .Z(n6034) );
  XNOR U14103 ( .A(n6028), .B(n6029), .Z(n6032) );
  XNOR U14104 ( .A(y[7866]), .B(x[7866]), .Z(n6029) );
  XNOR U14105 ( .A(n6030), .B(n6031), .Z(n6028) );
  XNOR U14106 ( .A(y[7867]), .B(x[7867]), .Z(n6031) );
  XNOR U14107 ( .A(y[7868]), .B(x[7868]), .Z(n6030) );
  XNOR U14108 ( .A(n6022), .B(n6023), .Z(n6033) );
  XNOR U14109 ( .A(y[7863]), .B(x[7863]), .Z(n6023) );
  XNOR U14110 ( .A(n6024), .B(n6025), .Z(n6022) );
  XNOR U14111 ( .A(y[7864]), .B(x[7864]), .Z(n6025) );
  XNOR U14112 ( .A(y[7865]), .B(x[7865]), .Z(n6024) );
  NAND U14113 ( .A(n6089), .B(n6090), .Z(N64847) );
  NANDN U14114 ( .A(n6091), .B(n6092), .Z(n6090) );
  OR U14115 ( .A(n6093), .B(n6094), .Z(n6092) );
  NAND U14116 ( .A(n6093), .B(n6094), .Z(n6089) );
  XOR U14117 ( .A(n6093), .B(n6095), .Z(N64846) );
  XNOR U14118 ( .A(n6091), .B(n6094), .Z(n6095) );
  AND U14119 ( .A(n6096), .B(n6097), .Z(n6094) );
  NANDN U14120 ( .A(n6098), .B(n6099), .Z(n6097) );
  NANDN U14121 ( .A(n6100), .B(n6101), .Z(n6099) );
  NANDN U14122 ( .A(n6101), .B(n6100), .Z(n6096) );
  NAND U14123 ( .A(n6102), .B(n6103), .Z(n6091) );
  NANDN U14124 ( .A(n6104), .B(n6105), .Z(n6103) );
  OR U14125 ( .A(n6106), .B(n6107), .Z(n6105) );
  NAND U14126 ( .A(n6107), .B(n6106), .Z(n6102) );
  AND U14127 ( .A(n6108), .B(n6109), .Z(n6093) );
  NANDN U14128 ( .A(n6110), .B(n6111), .Z(n6109) );
  NANDN U14129 ( .A(n6112), .B(n6113), .Z(n6111) );
  NANDN U14130 ( .A(n6113), .B(n6112), .Z(n6108) );
  XOR U14131 ( .A(n6107), .B(n6114), .Z(N64845) );
  XOR U14132 ( .A(n6104), .B(n6106), .Z(n6114) );
  XNOR U14133 ( .A(n6100), .B(n6115), .Z(n6106) );
  XNOR U14134 ( .A(n6098), .B(n6101), .Z(n6115) );
  NAND U14135 ( .A(n6116), .B(n6117), .Z(n6101) );
  NAND U14136 ( .A(n6118), .B(n6119), .Z(n6117) );
  OR U14137 ( .A(n6120), .B(n6121), .Z(n6118) );
  NANDN U14138 ( .A(n6122), .B(n6120), .Z(n6116) );
  IV U14139 ( .A(n6121), .Z(n6122) );
  NAND U14140 ( .A(n6123), .B(n6124), .Z(n6098) );
  NAND U14141 ( .A(n6125), .B(n6126), .Z(n6124) );
  NANDN U14142 ( .A(n6127), .B(n6128), .Z(n6125) );
  NANDN U14143 ( .A(n6128), .B(n6127), .Z(n6123) );
  AND U14144 ( .A(n6129), .B(n6130), .Z(n6100) );
  NAND U14145 ( .A(n6131), .B(n6132), .Z(n6130) );
  OR U14146 ( .A(n6133), .B(n6134), .Z(n6131) );
  NANDN U14147 ( .A(n6135), .B(n6133), .Z(n6129) );
  NAND U14148 ( .A(n6136), .B(n6137), .Z(n6104) );
  NANDN U14149 ( .A(n6138), .B(n6139), .Z(n6137) );
  OR U14150 ( .A(n6140), .B(n6141), .Z(n6139) );
  NANDN U14151 ( .A(n6142), .B(n6140), .Z(n6136) );
  IV U14152 ( .A(n6141), .Z(n6142) );
  XNOR U14153 ( .A(n6112), .B(n6143), .Z(n6107) );
  XNOR U14154 ( .A(n6110), .B(n6113), .Z(n6143) );
  NAND U14155 ( .A(n6144), .B(n6145), .Z(n6113) );
  NAND U14156 ( .A(n6146), .B(n6147), .Z(n6145) );
  OR U14157 ( .A(n6148), .B(n6149), .Z(n6146) );
  NANDN U14158 ( .A(n6150), .B(n6148), .Z(n6144) );
  IV U14159 ( .A(n6149), .Z(n6150) );
  NAND U14160 ( .A(n6151), .B(n6152), .Z(n6110) );
  NAND U14161 ( .A(n6153), .B(n6154), .Z(n6152) );
  NANDN U14162 ( .A(n6155), .B(n6156), .Z(n6153) );
  NANDN U14163 ( .A(n6156), .B(n6155), .Z(n6151) );
  AND U14164 ( .A(n6157), .B(n6158), .Z(n6112) );
  NAND U14165 ( .A(n6159), .B(n6160), .Z(n6158) );
  OR U14166 ( .A(n6161), .B(n6162), .Z(n6159) );
  NANDN U14167 ( .A(n6163), .B(n6161), .Z(n6157) );
  XNOR U14168 ( .A(n6138), .B(n6164), .Z(N64844) );
  XOR U14169 ( .A(n6140), .B(n6141), .Z(n6164) );
  XNOR U14170 ( .A(n6154), .B(n6165), .Z(n6141) );
  XOR U14171 ( .A(n6155), .B(n6156), .Z(n6165) );
  XOR U14172 ( .A(n6161), .B(n6166), .Z(n6156) );
  XOR U14173 ( .A(n6160), .B(n6163), .Z(n6166) );
  IV U14174 ( .A(n6162), .Z(n6163) );
  NAND U14175 ( .A(n6167), .B(n6168), .Z(n6162) );
  OR U14176 ( .A(n6169), .B(n6170), .Z(n6168) );
  OR U14177 ( .A(n6171), .B(n6172), .Z(n6167) );
  NAND U14178 ( .A(n6173), .B(n6174), .Z(n6160) );
  OR U14179 ( .A(n6175), .B(n6176), .Z(n6174) );
  OR U14180 ( .A(n6177), .B(n6178), .Z(n6173) );
  NOR U14181 ( .A(n6179), .B(n6180), .Z(n6161) );
  ANDN U14182 ( .B(n6181), .A(n6182), .Z(n6155) );
  XNOR U14183 ( .A(n6148), .B(n6183), .Z(n6154) );
  XNOR U14184 ( .A(n6147), .B(n6149), .Z(n6183) );
  NAND U14185 ( .A(n6184), .B(n6185), .Z(n6149) );
  OR U14186 ( .A(n6186), .B(n6187), .Z(n6185) );
  OR U14187 ( .A(n6188), .B(n6189), .Z(n6184) );
  NAND U14188 ( .A(n6190), .B(n6191), .Z(n6147) );
  OR U14189 ( .A(n6192), .B(n6193), .Z(n6191) );
  OR U14190 ( .A(n6194), .B(n6195), .Z(n6190) );
  ANDN U14191 ( .B(n6196), .A(n6197), .Z(n6148) );
  IV U14192 ( .A(n6198), .Z(n6196) );
  ANDN U14193 ( .B(n6199), .A(n6200), .Z(n6140) );
  XOR U14194 ( .A(n6126), .B(n6201), .Z(n6138) );
  XOR U14195 ( .A(n6127), .B(n6128), .Z(n6201) );
  XOR U14196 ( .A(n6133), .B(n6202), .Z(n6128) );
  XOR U14197 ( .A(n6132), .B(n6135), .Z(n6202) );
  IV U14198 ( .A(n6134), .Z(n6135) );
  NAND U14199 ( .A(n6203), .B(n6204), .Z(n6134) );
  OR U14200 ( .A(n6205), .B(n6206), .Z(n6204) );
  OR U14201 ( .A(n6207), .B(n6208), .Z(n6203) );
  NAND U14202 ( .A(n6209), .B(n6210), .Z(n6132) );
  OR U14203 ( .A(n6211), .B(n6212), .Z(n6210) );
  OR U14204 ( .A(n6213), .B(n6214), .Z(n6209) );
  NOR U14205 ( .A(n6215), .B(n6216), .Z(n6133) );
  ANDN U14206 ( .B(n6217), .A(n6218), .Z(n6127) );
  IV U14207 ( .A(n6219), .Z(n6217) );
  XNOR U14208 ( .A(n6120), .B(n6220), .Z(n6126) );
  XNOR U14209 ( .A(n6119), .B(n6121), .Z(n6220) );
  NAND U14210 ( .A(n6221), .B(n6222), .Z(n6121) );
  OR U14211 ( .A(n6223), .B(n6224), .Z(n6222) );
  OR U14212 ( .A(n6225), .B(n6226), .Z(n6221) );
  NAND U14213 ( .A(n6227), .B(n6228), .Z(n6119) );
  OR U14214 ( .A(n6229), .B(n6230), .Z(n6228) );
  OR U14215 ( .A(n6231), .B(n6232), .Z(n6227) );
  ANDN U14216 ( .B(n6233), .A(n6234), .Z(n6120) );
  IV U14217 ( .A(n6235), .Z(n6233) );
  XNOR U14218 ( .A(n6200), .B(n6199), .Z(N64843) );
  XOR U14219 ( .A(n6219), .B(n6218), .Z(n6199) );
  XNOR U14220 ( .A(n6234), .B(n6235), .Z(n6218) );
  XNOR U14221 ( .A(n6229), .B(n6230), .Z(n6235) );
  XNOR U14222 ( .A(n6231), .B(n6232), .Z(n6230) );
  XNOR U14223 ( .A(y[7861]), .B(x[7861]), .Z(n6232) );
  XNOR U14224 ( .A(y[7862]), .B(x[7862]), .Z(n6231) );
  XNOR U14225 ( .A(y[7860]), .B(x[7860]), .Z(n6229) );
  XNOR U14226 ( .A(n6223), .B(n6224), .Z(n6234) );
  XNOR U14227 ( .A(y[7857]), .B(x[7857]), .Z(n6224) );
  XNOR U14228 ( .A(n6225), .B(n6226), .Z(n6223) );
  XNOR U14229 ( .A(y[7858]), .B(x[7858]), .Z(n6226) );
  XNOR U14230 ( .A(y[7859]), .B(x[7859]), .Z(n6225) );
  XNOR U14231 ( .A(n6216), .B(n6215), .Z(n6219) );
  XNOR U14232 ( .A(n6211), .B(n6212), .Z(n6215) );
  XNOR U14233 ( .A(y[7854]), .B(x[7854]), .Z(n6212) );
  XNOR U14234 ( .A(n6213), .B(n6214), .Z(n6211) );
  XNOR U14235 ( .A(y[7855]), .B(x[7855]), .Z(n6214) );
  XNOR U14236 ( .A(y[7856]), .B(x[7856]), .Z(n6213) );
  XNOR U14237 ( .A(n6205), .B(n6206), .Z(n6216) );
  XNOR U14238 ( .A(y[7851]), .B(x[7851]), .Z(n6206) );
  XNOR U14239 ( .A(n6207), .B(n6208), .Z(n6205) );
  XNOR U14240 ( .A(y[7852]), .B(x[7852]), .Z(n6208) );
  XNOR U14241 ( .A(y[7853]), .B(x[7853]), .Z(n6207) );
  XOR U14242 ( .A(n6181), .B(n6182), .Z(n6200) );
  XNOR U14243 ( .A(n6197), .B(n6198), .Z(n6182) );
  XNOR U14244 ( .A(n6192), .B(n6193), .Z(n6198) );
  XNOR U14245 ( .A(n6194), .B(n6195), .Z(n6193) );
  XNOR U14246 ( .A(y[7849]), .B(x[7849]), .Z(n6195) );
  XNOR U14247 ( .A(y[7850]), .B(x[7850]), .Z(n6194) );
  XNOR U14248 ( .A(y[7848]), .B(x[7848]), .Z(n6192) );
  XNOR U14249 ( .A(n6186), .B(n6187), .Z(n6197) );
  XNOR U14250 ( .A(y[7845]), .B(x[7845]), .Z(n6187) );
  XNOR U14251 ( .A(n6188), .B(n6189), .Z(n6186) );
  XNOR U14252 ( .A(y[7846]), .B(x[7846]), .Z(n6189) );
  XNOR U14253 ( .A(y[7847]), .B(x[7847]), .Z(n6188) );
  XOR U14254 ( .A(n6180), .B(n6179), .Z(n6181) );
  XNOR U14255 ( .A(n6175), .B(n6176), .Z(n6179) );
  XNOR U14256 ( .A(y[7842]), .B(x[7842]), .Z(n6176) );
  XNOR U14257 ( .A(n6177), .B(n6178), .Z(n6175) );
  XNOR U14258 ( .A(y[7843]), .B(x[7843]), .Z(n6178) );
  XNOR U14259 ( .A(y[7844]), .B(x[7844]), .Z(n6177) );
  XNOR U14260 ( .A(n6169), .B(n6170), .Z(n6180) );
  XNOR U14261 ( .A(y[7839]), .B(x[7839]), .Z(n6170) );
  XNOR U14262 ( .A(n6171), .B(n6172), .Z(n6169) );
  XNOR U14263 ( .A(y[7840]), .B(x[7840]), .Z(n6172) );
  XNOR U14264 ( .A(y[7841]), .B(x[7841]), .Z(n6171) );
  NAND U14265 ( .A(n6236), .B(n6237), .Z(N64834) );
  NANDN U14266 ( .A(n6238), .B(n6239), .Z(n6237) );
  OR U14267 ( .A(n6240), .B(n6241), .Z(n6239) );
  NAND U14268 ( .A(n6240), .B(n6241), .Z(n6236) );
  XOR U14269 ( .A(n6240), .B(n6242), .Z(N64833) );
  XNOR U14270 ( .A(n6238), .B(n6241), .Z(n6242) );
  AND U14271 ( .A(n6243), .B(n6244), .Z(n6241) );
  NANDN U14272 ( .A(n6245), .B(n6246), .Z(n6244) );
  NANDN U14273 ( .A(n6247), .B(n6248), .Z(n6246) );
  NANDN U14274 ( .A(n6248), .B(n6247), .Z(n6243) );
  NAND U14275 ( .A(n6249), .B(n6250), .Z(n6238) );
  NANDN U14276 ( .A(n6251), .B(n6252), .Z(n6250) );
  OR U14277 ( .A(n6253), .B(n6254), .Z(n6252) );
  NAND U14278 ( .A(n6254), .B(n6253), .Z(n6249) );
  AND U14279 ( .A(n6255), .B(n6256), .Z(n6240) );
  NANDN U14280 ( .A(n6257), .B(n6258), .Z(n6256) );
  NANDN U14281 ( .A(n6259), .B(n6260), .Z(n6258) );
  NANDN U14282 ( .A(n6260), .B(n6259), .Z(n6255) );
  XOR U14283 ( .A(n6254), .B(n6261), .Z(N64832) );
  XOR U14284 ( .A(n6251), .B(n6253), .Z(n6261) );
  XNOR U14285 ( .A(n6247), .B(n6262), .Z(n6253) );
  XNOR U14286 ( .A(n6245), .B(n6248), .Z(n6262) );
  NAND U14287 ( .A(n6263), .B(n6264), .Z(n6248) );
  NAND U14288 ( .A(n6265), .B(n6266), .Z(n6264) );
  OR U14289 ( .A(n6267), .B(n6268), .Z(n6265) );
  NANDN U14290 ( .A(n6269), .B(n6267), .Z(n6263) );
  IV U14291 ( .A(n6268), .Z(n6269) );
  NAND U14292 ( .A(n6270), .B(n6271), .Z(n6245) );
  NAND U14293 ( .A(n6272), .B(n6273), .Z(n6271) );
  NANDN U14294 ( .A(n6274), .B(n6275), .Z(n6272) );
  NANDN U14295 ( .A(n6275), .B(n6274), .Z(n6270) );
  AND U14296 ( .A(n6276), .B(n6277), .Z(n6247) );
  NAND U14297 ( .A(n6278), .B(n6279), .Z(n6277) );
  OR U14298 ( .A(n6280), .B(n6281), .Z(n6278) );
  NANDN U14299 ( .A(n6282), .B(n6280), .Z(n6276) );
  NAND U14300 ( .A(n6283), .B(n6284), .Z(n6251) );
  NANDN U14301 ( .A(n6285), .B(n6286), .Z(n6284) );
  OR U14302 ( .A(n6287), .B(n6288), .Z(n6286) );
  NANDN U14303 ( .A(n6289), .B(n6287), .Z(n6283) );
  IV U14304 ( .A(n6288), .Z(n6289) );
  XNOR U14305 ( .A(n6259), .B(n6290), .Z(n6254) );
  XNOR U14306 ( .A(n6257), .B(n6260), .Z(n6290) );
  NAND U14307 ( .A(n6291), .B(n6292), .Z(n6260) );
  NAND U14308 ( .A(n6293), .B(n6294), .Z(n6292) );
  OR U14309 ( .A(n6295), .B(n6296), .Z(n6293) );
  NANDN U14310 ( .A(n6297), .B(n6295), .Z(n6291) );
  IV U14311 ( .A(n6296), .Z(n6297) );
  NAND U14312 ( .A(n6298), .B(n6299), .Z(n6257) );
  NAND U14313 ( .A(n6300), .B(n6301), .Z(n6299) );
  NANDN U14314 ( .A(n6302), .B(n6303), .Z(n6300) );
  NANDN U14315 ( .A(n6303), .B(n6302), .Z(n6298) );
  AND U14316 ( .A(n6304), .B(n6305), .Z(n6259) );
  NAND U14317 ( .A(n6306), .B(n6307), .Z(n6305) );
  OR U14318 ( .A(n6308), .B(n6309), .Z(n6306) );
  NANDN U14319 ( .A(n6310), .B(n6308), .Z(n6304) );
  XNOR U14320 ( .A(n6285), .B(n6311), .Z(N64831) );
  XOR U14321 ( .A(n6287), .B(n6288), .Z(n6311) );
  XNOR U14322 ( .A(n6301), .B(n6312), .Z(n6288) );
  XOR U14323 ( .A(n6302), .B(n6303), .Z(n6312) );
  XOR U14324 ( .A(n6308), .B(n6313), .Z(n6303) );
  XOR U14325 ( .A(n6307), .B(n6310), .Z(n6313) );
  IV U14326 ( .A(n6309), .Z(n6310) );
  NAND U14327 ( .A(n6314), .B(n6315), .Z(n6309) );
  OR U14328 ( .A(n6316), .B(n6317), .Z(n6315) );
  OR U14329 ( .A(n6318), .B(n6319), .Z(n6314) );
  NAND U14330 ( .A(n6320), .B(n6321), .Z(n6307) );
  OR U14331 ( .A(n6322), .B(n6323), .Z(n6321) );
  OR U14332 ( .A(n6324), .B(n6325), .Z(n6320) );
  NOR U14333 ( .A(n6326), .B(n6327), .Z(n6308) );
  ANDN U14334 ( .B(n6328), .A(n6329), .Z(n6302) );
  XNOR U14335 ( .A(n6295), .B(n6330), .Z(n6301) );
  XNOR U14336 ( .A(n6294), .B(n6296), .Z(n6330) );
  NAND U14337 ( .A(n6331), .B(n6332), .Z(n6296) );
  OR U14338 ( .A(n6333), .B(n6334), .Z(n6332) );
  OR U14339 ( .A(n6335), .B(n6336), .Z(n6331) );
  NAND U14340 ( .A(n6337), .B(n6338), .Z(n6294) );
  OR U14341 ( .A(n6339), .B(n6340), .Z(n6338) );
  OR U14342 ( .A(n6341), .B(n6342), .Z(n6337) );
  ANDN U14343 ( .B(n6343), .A(n6344), .Z(n6295) );
  IV U14344 ( .A(n6345), .Z(n6343) );
  ANDN U14345 ( .B(n6346), .A(n6347), .Z(n6287) );
  XOR U14346 ( .A(n6273), .B(n6348), .Z(n6285) );
  XOR U14347 ( .A(n6274), .B(n6275), .Z(n6348) );
  XOR U14348 ( .A(n6280), .B(n6349), .Z(n6275) );
  XOR U14349 ( .A(n6279), .B(n6282), .Z(n6349) );
  IV U14350 ( .A(n6281), .Z(n6282) );
  NAND U14351 ( .A(n6350), .B(n6351), .Z(n6281) );
  OR U14352 ( .A(n6352), .B(n6353), .Z(n6351) );
  OR U14353 ( .A(n6354), .B(n6355), .Z(n6350) );
  NAND U14354 ( .A(n6356), .B(n6357), .Z(n6279) );
  OR U14355 ( .A(n6358), .B(n6359), .Z(n6357) );
  OR U14356 ( .A(n6360), .B(n6361), .Z(n6356) );
  NOR U14357 ( .A(n6362), .B(n6363), .Z(n6280) );
  ANDN U14358 ( .B(n6364), .A(n6365), .Z(n6274) );
  IV U14359 ( .A(n6366), .Z(n6364) );
  XNOR U14360 ( .A(n6267), .B(n6367), .Z(n6273) );
  XNOR U14361 ( .A(n6266), .B(n6268), .Z(n6367) );
  NAND U14362 ( .A(n6368), .B(n6369), .Z(n6268) );
  OR U14363 ( .A(n6370), .B(n6371), .Z(n6369) );
  OR U14364 ( .A(n6372), .B(n6373), .Z(n6368) );
  NAND U14365 ( .A(n6374), .B(n6375), .Z(n6266) );
  OR U14366 ( .A(n6376), .B(n6377), .Z(n6375) );
  OR U14367 ( .A(n6378), .B(n6379), .Z(n6374) );
  ANDN U14368 ( .B(n6380), .A(n6381), .Z(n6267) );
  IV U14369 ( .A(n6382), .Z(n6380) );
  XNOR U14370 ( .A(n6347), .B(n6346), .Z(N64830) );
  XOR U14371 ( .A(n6366), .B(n6365), .Z(n6346) );
  XNOR U14372 ( .A(n6381), .B(n6382), .Z(n6365) );
  XNOR U14373 ( .A(n6376), .B(n6377), .Z(n6382) );
  XNOR U14374 ( .A(n6378), .B(n6379), .Z(n6377) );
  XNOR U14375 ( .A(y[7837]), .B(x[7837]), .Z(n6379) );
  XNOR U14376 ( .A(y[7838]), .B(x[7838]), .Z(n6378) );
  XNOR U14377 ( .A(y[7836]), .B(x[7836]), .Z(n6376) );
  XNOR U14378 ( .A(n6370), .B(n6371), .Z(n6381) );
  XNOR U14379 ( .A(y[7833]), .B(x[7833]), .Z(n6371) );
  XNOR U14380 ( .A(n6372), .B(n6373), .Z(n6370) );
  XNOR U14381 ( .A(y[7834]), .B(x[7834]), .Z(n6373) );
  XNOR U14382 ( .A(y[7835]), .B(x[7835]), .Z(n6372) );
  XNOR U14383 ( .A(n6363), .B(n6362), .Z(n6366) );
  XNOR U14384 ( .A(n6358), .B(n6359), .Z(n6362) );
  XNOR U14385 ( .A(y[7830]), .B(x[7830]), .Z(n6359) );
  XNOR U14386 ( .A(n6360), .B(n6361), .Z(n6358) );
  XNOR U14387 ( .A(y[7831]), .B(x[7831]), .Z(n6361) );
  XNOR U14388 ( .A(y[7832]), .B(x[7832]), .Z(n6360) );
  XNOR U14389 ( .A(n6352), .B(n6353), .Z(n6363) );
  XNOR U14390 ( .A(y[7827]), .B(x[7827]), .Z(n6353) );
  XNOR U14391 ( .A(n6354), .B(n6355), .Z(n6352) );
  XNOR U14392 ( .A(y[7828]), .B(x[7828]), .Z(n6355) );
  XNOR U14393 ( .A(y[7829]), .B(x[7829]), .Z(n6354) );
  XOR U14394 ( .A(n6328), .B(n6329), .Z(n6347) );
  XNOR U14395 ( .A(n6344), .B(n6345), .Z(n6329) );
  XNOR U14396 ( .A(n6339), .B(n6340), .Z(n6345) );
  XNOR U14397 ( .A(n6341), .B(n6342), .Z(n6340) );
  XNOR U14398 ( .A(y[7825]), .B(x[7825]), .Z(n6342) );
  XNOR U14399 ( .A(y[7826]), .B(x[7826]), .Z(n6341) );
  XNOR U14400 ( .A(y[7824]), .B(x[7824]), .Z(n6339) );
  XNOR U14401 ( .A(n6333), .B(n6334), .Z(n6344) );
  XNOR U14402 ( .A(y[7821]), .B(x[7821]), .Z(n6334) );
  XNOR U14403 ( .A(n6335), .B(n6336), .Z(n6333) );
  XNOR U14404 ( .A(y[7822]), .B(x[7822]), .Z(n6336) );
  XNOR U14405 ( .A(y[7823]), .B(x[7823]), .Z(n6335) );
  XOR U14406 ( .A(n6327), .B(n6326), .Z(n6328) );
  XNOR U14407 ( .A(n6322), .B(n6323), .Z(n6326) );
  XNOR U14408 ( .A(y[7818]), .B(x[7818]), .Z(n6323) );
  XNOR U14409 ( .A(n6324), .B(n6325), .Z(n6322) );
  XNOR U14410 ( .A(y[7819]), .B(x[7819]), .Z(n6325) );
  XNOR U14411 ( .A(y[7820]), .B(x[7820]), .Z(n6324) );
  XNOR U14412 ( .A(n6316), .B(n6317), .Z(n6327) );
  XNOR U14413 ( .A(y[7815]), .B(x[7815]), .Z(n6317) );
  XNOR U14414 ( .A(n6318), .B(n6319), .Z(n6316) );
  XNOR U14415 ( .A(y[7816]), .B(x[7816]), .Z(n6319) );
  XNOR U14416 ( .A(y[7817]), .B(x[7817]), .Z(n6318) );
  NAND U14417 ( .A(n6383), .B(n6384), .Z(N64821) );
  NANDN U14418 ( .A(n6385), .B(n6386), .Z(n6384) );
  OR U14419 ( .A(n6387), .B(n6388), .Z(n6386) );
  NAND U14420 ( .A(n6387), .B(n6388), .Z(n6383) );
  XOR U14421 ( .A(n6387), .B(n6389), .Z(N64820) );
  XNOR U14422 ( .A(n6385), .B(n6388), .Z(n6389) );
  AND U14423 ( .A(n6390), .B(n6391), .Z(n6388) );
  NANDN U14424 ( .A(n6392), .B(n6393), .Z(n6391) );
  NANDN U14425 ( .A(n6394), .B(n6395), .Z(n6393) );
  NANDN U14426 ( .A(n6395), .B(n6394), .Z(n6390) );
  NAND U14427 ( .A(n6396), .B(n6397), .Z(n6385) );
  NANDN U14428 ( .A(n6398), .B(n6399), .Z(n6397) );
  OR U14429 ( .A(n6400), .B(n6401), .Z(n6399) );
  NAND U14430 ( .A(n6401), .B(n6400), .Z(n6396) );
  AND U14431 ( .A(n6402), .B(n6403), .Z(n6387) );
  NANDN U14432 ( .A(n6404), .B(n6405), .Z(n6403) );
  NANDN U14433 ( .A(n6406), .B(n6407), .Z(n6405) );
  NANDN U14434 ( .A(n6407), .B(n6406), .Z(n6402) );
  XOR U14435 ( .A(n6401), .B(n6408), .Z(N64819) );
  XOR U14436 ( .A(n6398), .B(n6400), .Z(n6408) );
  XNOR U14437 ( .A(n6394), .B(n6409), .Z(n6400) );
  XNOR U14438 ( .A(n6392), .B(n6395), .Z(n6409) );
  NAND U14439 ( .A(n6410), .B(n6411), .Z(n6395) );
  NAND U14440 ( .A(n6412), .B(n6413), .Z(n6411) );
  OR U14441 ( .A(n6414), .B(n6415), .Z(n6412) );
  NANDN U14442 ( .A(n6416), .B(n6414), .Z(n6410) );
  IV U14443 ( .A(n6415), .Z(n6416) );
  NAND U14444 ( .A(n6417), .B(n6418), .Z(n6392) );
  NAND U14445 ( .A(n6419), .B(n6420), .Z(n6418) );
  NANDN U14446 ( .A(n6421), .B(n6422), .Z(n6419) );
  NANDN U14447 ( .A(n6422), .B(n6421), .Z(n6417) );
  AND U14448 ( .A(n6423), .B(n6424), .Z(n6394) );
  NAND U14449 ( .A(n6425), .B(n6426), .Z(n6424) );
  OR U14450 ( .A(n6427), .B(n6428), .Z(n6425) );
  NANDN U14451 ( .A(n6429), .B(n6427), .Z(n6423) );
  NAND U14452 ( .A(n6430), .B(n6431), .Z(n6398) );
  NANDN U14453 ( .A(n6432), .B(n6433), .Z(n6431) );
  OR U14454 ( .A(n6434), .B(n6435), .Z(n6433) );
  NANDN U14455 ( .A(n6436), .B(n6434), .Z(n6430) );
  IV U14456 ( .A(n6435), .Z(n6436) );
  XNOR U14457 ( .A(n6406), .B(n6437), .Z(n6401) );
  XNOR U14458 ( .A(n6404), .B(n6407), .Z(n6437) );
  NAND U14459 ( .A(n6438), .B(n6439), .Z(n6407) );
  NAND U14460 ( .A(n6440), .B(n6441), .Z(n6439) );
  OR U14461 ( .A(n6442), .B(n6443), .Z(n6440) );
  NANDN U14462 ( .A(n6444), .B(n6442), .Z(n6438) );
  IV U14463 ( .A(n6443), .Z(n6444) );
  NAND U14464 ( .A(n6445), .B(n6446), .Z(n6404) );
  NAND U14465 ( .A(n6447), .B(n6448), .Z(n6446) );
  NANDN U14466 ( .A(n6449), .B(n6450), .Z(n6447) );
  NANDN U14467 ( .A(n6450), .B(n6449), .Z(n6445) );
  AND U14468 ( .A(n6451), .B(n6452), .Z(n6406) );
  NAND U14469 ( .A(n6453), .B(n6454), .Z(n6452) );
  OR U14470 ( .A(n6455), .B(n6456), .Z(n6453) );
  NANDN U14471 ( .A(n6457), .B(n6455), .Z(n6451) );
  XNOR U14472 ( .A(n6432), .B(n6458), .Z(N64818) );
  XOR U14473 ( .A(n6434), .B(n6435), .Z(n6458) );
  XNOR U14474 ( .A(n6448), .B(n6459), .Z(n6435) );
  XOR U14475 ( .A(n6449), .B(n6450), .Z(n6459) );
  XOR U14476 ( .A(n6455), .B(n6460), .Z(n6450) );
  XOR U14477 ( .A(n6454), .B(n6457), .Z(n6460) );
  IV U14478 ( .A(n6456), .Z(n6457) );
  NAND U14479 ( .A(n6461), .B(n6462), .Z(n6456) );
  OR U14480 ( .A(n6463), .B(n6464), .Z(n6462) );
  OR U14481 ( .A(n6465), .B(n6466), .Z(n6461) );
  NAND U14482 ( .A(n6467), .B(n6468), .Z(n6454) );
  OR U14483 ( .A(n6469), .B(n6470), .Z(n6468) );
  OR U14484 ( .A(n6471), .B(n6472), .Z(n6467) );
  NOR U14485 ( .A(n6473), .B(n6474), .Z(n6455) );
  ANDN U14486 ( .B(n6475), .A(n6476), .Z(n6449) );
  XNOR U14487 ( .A(n6442), .B(n6477), .Z(n6448) );
  XNOR U14488 ( .A(n6441), .B(n6443), .Z(n6477) );
  NAND U14489 ( .A(n6478), .B(n6479), .Z(n6443) );
  OR U14490 ( .A(n6480), .B(n6481), .Z(n6479) );
  OR U14491 ( .A(n6482), .B(n6483), .Z(n6478) );
  NAND U14492 ( .A(n6484), .B(n6485), .Z(n6441) );
  OR U14493 ( .A(n6486), .B(n6487), .Z(n6485) );
  OR U14494 ( .A(n6488), .B(n6489), .Z(n6484) );
  ANDN U14495 ( .B(n6490), .A(n6491), .Z(n6442) );
  IV U14496 ( .A(n6492), .Z(n6490) );
  ANDN U14497 ( .B(n6493), .A(n6494), .Z(n6434) );
  XOR U14498 ( .A(n6420), .B(n6495), .Z(n6432) );
  XOR U14499 ( .A(n6421), .B(n6422), .Z(n6495) );
  XOR U14500 ( .A(n6427), .B(n6496), .Z(n6422) );
  XOR U14501 ( .A(n6426), .B(n6429), .Z(n6496) );
  IV U14502 ( .A(n6428), .Z(n6429) );
  NAND U14503 ( .A(n6497), .B(n6498), .Z(n6428) );
  OR U14504 ( .A(n6499), .B(n6500), .Z(n6498) );
  OR U14505 ( .A(n6501), .B(n6502), .Z(n6497) );
  NAND U14506 ( .A(n6503), .B(n6504), .Z(n6426) );
  OR U14507 ( .A(n6505), .B(n6506), .Z(n6504) );
  OR U14508 ( .A(n6507), .B(n6508), .Z(n6503) );
  NOR U14509 ( .A(n6509), .B(n6510), .Z(n6427) );
  ANDN U14510 ( .B(n6511), .A(n6512), .Z(n6421) );
  IV U14511 ( .A(n6513), .Z(n6511) );
  XNOR U14512 ( .A(n6414), .B(n6514), .Z(n6420) );
  XNOR U14513 ( .A(n6413), .B(n6415), .Z(n6514) );
  NAND U14514 ( .A(n6515), .B(n6516), .Z(n6415) );
  OR U14515 ( .A(n6517), .B(n6518), .Z(n6516) );
  OR U14516 ( .A(n6519), .B(n6520), .Z(n6515) );
  NAND U14517 ( .A(n6521), .B(n6522), .Z(n6413) );
  OR U14518 ( .A(n6523), .B(n6524), .Z(n6522) );
  OR U14519 ( .A(n6525), .B(n6526), .Z(n6521) );
  ANDN U14520 ( .B(n6527), .A(n6528), .Z(n6414) );
  IV U14521 ( .A(n6529), .Z(n6527) );
  XNOR U14522 ( .A(n6494), .B(n6493), .Z(N64817) );
  XOR U14523 ( .A(n6513), .B(n6512), .Z(n6493) );
  XNOR U14524 ( .A(n6528), .B(n6529), .Z(n6512) );
  XNOR U14525 ( .A(n6523), .B(n6524), .Z(n6529) );
  XNOR U14526 ( .A(n6525), .B(n6526), .Z(n6524) );
  XNOR U14527 ( .A(y[7813]), .B(x[7813]), .Z(n6526) );
  XNOR U14528 ( .A(y[7814]), .B(x[7814]), .Z(n6525) );
  XNOR U14529 ( .A(y[7812]), .B(x[7812]), .Z(n6523) );
  XNOR U14530 ( .A(n6517), .B(n6518), .Z(n6528) );
  XNOR U14531 ( .A(y[7809]), .B(x[7809]), .Z(n6518) );
  XNOR U14532 ( .A(n6519), .B(n6520), .Z(n6517) );
  XNOR U14533 ( .A(y[7810]), .B(x[7810]), .Z(n6520) );
  XNOR U14534 ( .A(y[7811]), .B(x[7811]), .Z(n6519) );
  XNOR U14535 ( .A(n6510), .B(n6509), .Z(n6513) );
  XNOR U14536 ( .A(n6505), .B(n6506), .Z(n6509) );
  XNOR U14537 ( .A(y[7806]), .B(x[7806]), .Z(n6506) );
  XNOR U14538 ( .A(n6507), .B(n6508), .Z(n6505) );
  XNOR U14539 ( .A(y[7807]), .B(x[7807]), .Z(n6508) );
  XNOR U14540 ( .A(y[7808]), .B(x[7808]), .Z(n6507) );
  XNOR U14541 ( .A(n6499), .B(n6500), .Z(n6510) );
  XNOR U14542 ( .A(y[7803]), .B(x[7803]), .Z(n6500) );
  XNOR U14543 ( .A(n6501), .B(n6502), .Z(n6499) );
  XNOR U14544 ( .A(y[7804]), .B(x[7804]), .Z(n6502) );
  XNOR U14545 ( .A(y[7805]), .B(x[7805]), .Z(n6501) );
  XOR U14546 ( .A(n6475), .B(n6476), .Z(n6494) );
  XNOR U14547 ( .A(n6491), .B(n6492), .Z(n6476) );
  XNOR U14548 ( .A(n6486), .B(n6487), .Z(n6492) );
  XNOR U14549 ( .A(n6488), .B(n6489), .Z(n6487) );
  XNOR U14550 ( .A(y[7801]), .B(x[7801]), .Z(n6489) );
  XNOR U14551 ( .A(y[7802]), .B(x[7802]), .Z(n6488) );
  XNOR U14552 ( .A(y[7800]), .B(x[7800]), .Z(n6486) );
  XNOR U14553 ( .A(n6480), .B(n6481), .Z(n6491) );
  XNOR U14554 ( .A(y[7797]), .B(x[7797]), .Z(n6481) );
  XNOR U14555 ( .A(n6482), .B(n6483), .Z(n6480) );
  XNOR U14556 ( .A(y[7798]), .B(x[7798]), .Z(n6483) );
  XNOR U14557 ( .A(y[7799]), .B(x[7799]), .Z(n6482) );
  XOR U14558 ( .A(n6474), .B(n6473), .Z(n6475) );
  XNOR U14559 ( .A(n6469), .B(n6470), .Z(n6473) );
  XNOR U14560 ( .A(y[7794]), .B(x[7794]), .Z(n6470) );
  XNOR U14561 ( .A(n6471), .B(n6472), .Z(n6469) );
  XNOR U14562 ( .A(y[7795]), .B(x[7795]), .Z(n6472) );
  XNOR U14563 ( .A(y[7796]), .B(x[7796]), .Z(n6471) );
  XNOR U14564 ( .A(n6463), .B(n6464), .Z(n6474) );
  XNOR U14565 ( .A(y[7791]), .B(x[7791]), .Z(n6464) );
  XNOR U14566 ( .A(n6465), .B(n6466), .Z(n6463) );
  XNOR U14567 ( .A(y[7792]), .B(x[7792]), .Z(n6466) );
  XNOR U14568 ( .A(y[7793]), .B(x[7793]), .Z(n6465) );
  NAND U14569 ( .A(n6530), .B(n6531), .Z(N64808) );
  NANDN U14570 ( .A(n6532), .B(n6533), .Z(n6531) );
  OR U14571 ( .A(n6534), .B(n6535), .Z(n6533) );
  NAND U14572 ( .A(n6534), .B(n6535), .Z(n6530) );
  XOR U14573 ( .A(n6534), .B(n6536), .Z(N64807) );
  XNOR U14574 ( .A(n6532), .B(n6535), .Z(n6536) );
  AND U14575 ( .A(n6537), .B(n6538), .Z(n6535) );
  NANDN U14576 ( .A(n6539), .B(n6540), .Z(n6538) );
  NANDN U14577 ( .A(n6541), .B(n6542), .Z(n6540) );
  NANDN U14578 ( .A(n6542), .B(n6541), .Z(n6537) );
  NAND U14579 ( .A(n6543), .B(n6544), .Z(n6532) );
  NANDN U14580 ( .A(n6545), .B(n6546), .Z(n6544) );
  OR U14581 ( .A(n6547), .B(n6548), .Z(n6546) );
  NAND U14582 ( .A(n6548), .B(n6547), .Z(n6543) );
  AND U14583 ( .A(n6549), .B(n6550), .Z(n6534) );
  NANDN U14584 ( .A(n6551), .B(n6552), .Z(n6550) );
  NANDN U14585 ( .A(n6553), .B(n6554), .Z(n6552) );
  NANDN U14586 ( .A(n6554), .B(n6553), .Z(n6549) );
  XOR U14587 ( .A(n6548), .B(n6555), .Z(N64806) );
  XOR U14588 ( .A(n6545), .B(n6547), .Z(n6555) );
  XNOR U14589 ( .A(n6541), .B(n6556), .Z(n6547) );
  XNOR U14590 ( .A(n6539), .B(n6542), .Z(n6556) );
  NAND U14591 ( .A(n6557), .B(n6558), .Z(n6542) );
  NAND U14592 ( .A(n6559), .B(n6560), .Z(n6558) );
  OR U14593 ( .A(n6561), .B(n6562), .Z(n6559) );
  NANDN U14594 ( .A(n6563), .B(n6561), .Z(n6557) );
  IV U14595 ( .A(n6562), .Z(n6563) );
  NAND U14596 ( .A(n6564), .B(n6565), .Z(n6539) );
  NAND U14597 ( .A(n6566), .B(n6567), .Z(n6565) );
  NANDN U14598 ( .A(n6568), .B(n6569), .Z(n6566) );
  NANDN U14599 ( .A(n6569), .B(n6568), .Z(n6564) );
  AND U14600 ( .A(n6570), .B(n6571), .Z(n6541) );
  NAND U14601 ( .A(n6572), .B(n6573), .Z(n6571) );
  OR U14602 ( .A(n6574), .B(n6575), .Z(n6572) );
  NANDN U14603 ( .A(n6576), .B(n6574), .Z(n6570) );
  NAND U14604 ( .A(n6577), .B(n6578), .Z(n6545) );
  NANDN U14605 ( .A(n6579), .B(n6580), .Z(n6578) );
  OR U14606 ( .A(n6581), .B(n6582), .Z(n6580) );
  NANDN U14607 ( .A(n6583), .B(n6581), .Z(n6577) );
  IV U14608 ( .A(n6582), .Z(n6583) );
  XNOR U14609 ( .A(n6553), .B(n6584), .Z(n6548) );
  XNOR U14610 ( .A(n6551), .B(n6554), .Z(n6584) );
  NAND U14611 ( .A(n6585), .B(n6586), .Z(n6554) );
  NAND U14612 ( .A(n6587), .B(n6588), .Z(n6586) );
  OR U14613 ( .A(n6589), .B(n6590), .Z(n6587) );
  NANDN U14614 ( .A(n6591), .B(n6589), .Z(n6585) );
  IV U14615 ( .A(n6590), .Z(n6591) );
  NAND U14616 ( .A(n6592), .B(n6593), .Z(n6551) );
  NAND U14617 ( .A(n6594), .B(n6595), .Z(n6593) );
  NANDN U14618 ( .A(n6596), .B(n6597), .Z(n6594) );
  NANDN U14619 ( .A(n6597), .B(n6596), .Z(n6592) );
  AND U14620 ( .A(n6598), .B(n6599), .Z(n6553) );
  NAND U14621 ( .A(n6600), .B(n6601), .Z(n6599) );
  OR U14622 ( .A(n6602), .B(n6603), .Z(n6600) );
  NANDN U14623 ( .A(n6604), .B(n6602), .Z(n6598) );
  XNOR U14624 ( .A(n6579), .B(n6605), .Z(N64805) );
  XOR U14625 ( .A(n6581), .B(n6582), .Z(n6605) );
  XNOR U14626 ( .A(n6595), .B(n6606), .Z(n6582) );
  XOR U14627 ( .A(n6596), .B(n6597), .Z(n6606) );
  XOR U14628 ( .A(n6602), .B(n6607), .Z(n6597) );
  XOR U14629 ( .A(n6601), .B(n6604), .Z(n6607) );
  IV U14630 ( .A(n6603), .Z(n6604) );
  NAND U14631 ( .A(n6608), .B(n6609), .Z(n6603) );
  OR U14632 ( .A(n6610), .B(n6611), .Z(n6609) );
  OR U14633 ( .A(n6612), .B(n6613), .Z(n6608) );
  NAND U14634 ( .A(n6614), .B(n6615), .Z(n6601) );
  OR U14635 ( .A(n6616), .B(n6617), .Z(n6615) );
  OR U14636 ( .A(n6618), .B(n6619), .Z(n6614) );
  NOR U14637 ( .A(n6620), .B(n6621), .Z(n6602) );
  ANDN U14638 ( .B(n6622), .A(n6623), .Z(n6596) );
  XNOR U14639 ( .A(n6589), .B(n6624), .Z(n6595) );
  XNOR U14640 ( .A(n6588), .B(n6590), .Z(n6624) );
  NAND U14641 ( .A(n6625), .B(n6626), .Z(n6590) );
  OR U14642 ( .A(n6627), .B(n6628), .Z(n6626) );
  OR U14643 ( .A(n6629), .B(n6630), .Z(n6625) );
  NAND U14644 ( .A(n6631), .B(n6632), .Z(n6588) );
  OR U14645 ( .A(n6633), .B(n6634), .Z(n6632) );
  OR U14646 ( .A(n6635), .B(n6636), .Z(n6631) );
  ANDN U14647 ( .B(n6637), .A(n6638), .Z(n6589) );
  IV U14648 ( .A(n6639), .Z(n6637) );
  ANDN U14649 ( .B(n6640), .A(n6641), .Z(n6581) );
  XOR U14650 ( .A(n6567), .B(n6642), .Z(n6579) );
  XOR U14651 ( .A(n6568), .B(n6569), .Z(n6642) );
  XOR U14652 ( .A(n6574), .B(n6643), .Z(n6569) );
  XOR U14653 ( .A(n6573), .B(n6576), .Z(n6643) );
  IV U14654 ( .A(n6575), .Z(n6576) );
  NAND U14655 ( .A(n6644), .B(n6645), .Z(n6575) );
  OR U14656 ( .A(n6646), .B(n6647), .Z(n6645) );
  OR U14657 ( .A(n6648), .B(n6649), .Z(n6644) );
  NAND U14658 ( .A(n6650), .B(n6651), .Z(n6573) );
  OR U14659 ( .A(n6652), .B(n6653), .Z(n6651) );
  OR U14660 ( .A(n6654), .B(n6655), .Z(n6650) );
  NOR U14661 ( .A(n6656), .B(n6657), .Z(n6574) );
  ANDN U14662 ( .B(n6658), .A(n6659), .Z(n6568) );
  IV U14663 ( .A(n6660), .Z(n6658) );
  XNOR U14664 ( .A(n6561), .B(n6661), .Z(n6567) );
  XNOR U14665 ( .A(n6560), .B(n6562), .Z(n6661) );
  NAND U14666 ( .A(n6662), .B(n6663), .Z(n6562) );
  OR U14667 ( .A(n6664), .B(n6665), .Z(n6663) );
  OR U14668 ( .A(n6666), .B(n6667), .Z(n6662) );
  NAND U14669 ( .A(n6668), .B(n6669), .Z(n6560) );
  OR U14670 ( .A(n6670), .B(n6671), .Z(n6669) );
  OR U14671 ( .A(n6672), .B(n6673), .Z(n6668) );
  ANDN U14672 ( .B(n6674), .A(n6675), .Z(n6561) );
  IV U14673 ( .A(n6676), .Z(n6674) );
  XNOR U14674 ( .A(n6641), .B(n6640), .Z(N64804) );
  XOR U14675 ( .A(n6660), .B(n6659), .Z(n6640) );
  XNOR U14676 ( .A(n6675), .B(n6676), .Z(n6659) );
  XNOR U14677 ( .A(n6670), .B(n6671), .Z(n6676) );
  XNOR U14678 ( .A(n6672), .B(n6673), .Z(n6671) );
  XNOR U14679 ( .A(y[7789]), .B(x[7789]), .Z(n6673) );
  XNOR U14680 ( .A(y[7790]), .B(x[7790]), .Z(n6672) );
  XNOR U14681 ( .A(y[7788]), .B(x[7788]), .Z(n6670) );
  XNOR U14682 ( .A(n6664), .B(n6665), .Z(n6675) );
  XNOR U14683 ( .A(y[7785]), .B(x[7785]), .Z(n6665) );
  XNOR U14684 ( .A(n6666), .B(n6667), .Z(n6664) );
  XNOR U14685 ( .A(y[7786]), .B(x[7786]), .Z(n6667) );
  XNOR U14686 ( .A(y[7787]), .B(x[7787]), .Z(n6666) );
  XNOR U14687 ( .A(n6657), .B(n6656), .Z(n6660) );
  XNOR U14688 ( .A(n6652), .B(n6653), .Z(n6656) );
  XNOR U14689 ( .A(y[7782]), .B(x[7782]), .Z(n6653) );
  XNOR U14690 ( .A(n6654), .B(n6655), .Z(n6652) );
  XNOR U14691 ( .A(y[7783]), .B(x[7783]), .Z(n6655) );
  XNOR U14692 ( .A(y[7784]), .B(x[7784]), .Z(n6654) );
  XNOR U14693 ( .A(n6646), .B(n6647), .Z(n6657) );
  XNOR U14694 ( .A(y[7779]), .B(x[7779]), .Z(n6647) );
  XNOR U14695 ( .A(n6648), .B(n6649), .Z(n6646) );
  XNOR U14696 ( .A(y[7780]), .B(x[7780]), .Z(n6649) );
  XNOR U14697 ( .A(y[7781]), .B(x[7781]), .Z(n6648) );
  XOR U14698 ( .A(n6622), .B(n6623), .Z(n6641) );
  XNOR U14699 ( .A(n6638), .B(n6639), .Z(n6623) );
  XNOR U14700 ( .A(n6633), .B(n6634), .Z(n6639) );
  XNOR U14701 ( .A(n6635), .B(n6636), .Z(n6634) );
  XNOR U14702 ( .A(y[7777]), .B(x[7777]), .Z(n6636) );
  XNOR U14703 ( .A(y[7778]), .B(x[7778]), .Z(n6635) );
  XNOR U14704 ( .A(y[7776]), .B(x[7776]), .Z(n6633) );
  XNOR U14705 ( .A(n6627), .B(n6628), .Z(n6638) );
  XNOR U14706 ( .A(y[7773]), .B(x[7773]), .Z(n6628) );
  XNOR U14707 ( .A(n6629), .B(n6630), .Z(n6627) );
  XNOR U14708 ( .A(y[7774]), .B(x[7774]), .Z(n6630) );
  XNOR U14709 ( .A(y[7775]), .B(x[7775]), .Z(n6629) );
  XOR U14710 ( .A(n6621), .B(n6620), .Z(n6622) );
  XNOR U14711 ( .A(n6616), .B(n6617), .Z(n6620) );
  XNOR U14712 ( .A(y[7770]), .B(x[7770]), .Z(n6617) );
  XNOR U14713 ( .A(n6618), .B(n6619), .Z(n6616) );
  XNOR U14714 ( .A(y[7771]), .B(x[7771]), .Z(n6619) );
  XNOR U14715 ( .A(y[7772]), .B(x[7772]), .Z(n6618) );
  XNOR U14716 ( .A(n6610), .B(n6611), .Z(n6621) );
  XNOR U14717 ( .A(y[7767]), .B(x[7767]), .Z(n6611) );
  XNOR U14718 ( .A(n6612), .B(n6613), .Z(n6610) );
  XNOR U14719 ( .A(y[7768]), .B(x[7768]), .Z(n6613) );
  XNOR U14720 ( .A(y[7769]), .B(x[7769]), .Z(n6612) );
  NAND U14721 ( .A(n6677), .B(n6678), .Z(N64795) );
  NANDN U14722 ( .A(n6679), .B(n6680), .Z(n6678) );
  OR U14723 ( .A(n6681), .B(n6682), .Z(n6680) );
  NAND U14724 ( .A(n6681), .B(n6682), .Z(n6677) );
  XOR U14725 ( .A(n6681), .B(n6683), .Z(N64794) );
  XNOR U14726 ( .A(n6679), .B(n6682), .Z(n6683) );
  AND U14727 ( .A(n6684), .B(n6685), .Z(n6682) );
  NANDN U14728 ( .A(n6686), .B(n6687), .Z(n6685) );
  NANDN U14729 ( .A(n6688), .B(n6689), .Z(n6687) );
  NANDN U14730 ( .A(n6689), .B(n6688), .Z(n6684) );
  NAND U14731 ( .A(n6690), .B(n6691), .Z(n6679) );
  NANDN U14732 ( .A(n6692), .B(n6693), .Z(n6691) );
  OR U14733 ( .A(n6694), .B(n6695), .Z(n6693) );
  NAND U14734 ( .A(n6695), .B(n6694), .Z(n6690) );
  AND U14735 ( .A(n6696), .B(n6697), .Z(n6681) );
  NANDN U14736 ( .A(n6698), .B(n6699), .Z(n6697) );
  NANDN U14737 ( .A(n6700), .B(n6701), .Z(n6699) );
  NANDN U14738 ( .A(n6701), .B(n6700), .Z(n6696) );
  XOR U14739 ( .A(n6695), .B(n6702), .Z(N64793) );
  XOR U14740 ( .A(n6692), .B(n6694), .Z(n6702) );
  XNOR U14741 ( .A(n6688), .B(n6703), .Z(n6694) );
  XNOR U14742 ( .A(n6686), .B(n6689), .Z(n6703) );
  NAND U14743 ( .A(n6704), .B(n6705), .Z(n6689) );
  NAND U14744 ( .A(n6706), .B(n6707), .Z(n6705) );
  OR U14745 ( .A(n6708), .B(n6709), .Z(n6706) );
  NANDN U14746 ( .A(n6710), .B(n6708), .Z(n6704) );
  IV U14747 ( .A(n6709), .Z(n6710) );
  NAND U14748 ( .A(n6711), .B(n6712), .Z(n6686) );
  NAND U14749 ( .A(n6713), .B(n6714), .Z(n6712) );
  NANDN U14750 ( .A(n6715), .B(n6716), .Z(n6713) );
  NANDN U14751 ( .A(n6716), .B(n6715), .Z(n6711) );
  AND U14752 ( .A(n6717), .B(n6718), .Z(n6688) );
  NAND U14753 ( .A(n6719), .B(n6720), .Z(n6718) );
  OR U14754 ( .A(n6721), .B(n6722), .Z(n6719) );
  NANDN U14755 ( .A(n6723), .B(n6721), .Z(n6717) );
  NAND U14756 ( .A(n6724), .B(n6725), .Z(n6692) );
  NANDN U14757 ( .A(n6726), .B(n6727), .Z(n6725) );
  OR U14758 ( .A(n6728), .B(n6729), .Z(n6727) );
  NANDN U14759 ( .A(n6730), .B(n6728), .Z(n6724) );
  IV U14760 ( .A(n6729), .Z(n6730) );
  XNOR U14761 ( .A(n6700), .B(n6731), .Z(n6695) );
  XNOR U14762 ( .A(n6698), .B(n6701), .Z(n6731) );
  NAND U14763 ( .A(n6732), .B(n6733), .Z(n6701) );
  NAND U14764 ( .A(n6734), .B(n6735), .Z(n6733) );
  OR U14765 ( .A(n6736), .B(n6737), .Z(n6734) );
  NANDN U14766 ( .A(n6738), .B(n6736), .Z(n6732) );
  IV U14767 ( .A(n6737), .Z(n6738) );
  NAND U14768 ( .A(n6739), .B(n6740), .Z(n6698) );
  NAND U14769 ( .A(n6741), .B(n6742), .Z(n6740) );
  NANDN U14770 ( .A(n6743), .B(n6744), .Z(n6741) );
  NANDN U14771 ( .A(n6744), .B(n6743), .Z(n6739) );
  AND U14772 ( .A(n6745), .B(n6746), .Z(n6700) );
  NAND U14773 ( .A(n6747), .B(n6748), .Z(n6746) );
  OR U14774 ( .A(n6749), .B(n6750), .Z(n6747) );
  NANDN U14775 ( .A(n6751), .B(n6749), .Z(n6745) );
  XNOR U14776 ( .A(n6726), .B(n6752), .Z(N64792) );
  XOR U14777 ( .A(n6728), .B(n6729), .Z(n6752) );
  XNOR U14778 ( .A(n6742), .B(n6753), .Z(n6729) );
  XOR U14779 ( .A(n6743), .B(n6744), .Z(n6753) );
  XOR U14780 ( .A(n6749), .B(n6754), .Z(n6744) );
  XOR U14781 ( .A(n6748), .B(n6751), .Z(n6754) );
  IV U14782 ( .A(n6750), .Z(n6751) );
  NAND U14783 ( .A(n6755), .B(n6756), .Z(n6750) );
  OR U14784 ( .A(n6757), .B(n6758), .Z(n6756) );
  OR U14785 ( .A(n6759), .B(n6760), .Z(n6755) );
  NAND U14786 ( .A(n6761), .B(n6762), .Z(n6748) );
  OR U14787 ( .A(n6763), .B(n6764), .Z(n6762) );
  OR U14788 ( .A(n6765), .B(n6766), .Z(n6761) );
  NOR U14789 ( .A(n6767), .B(n6768), .Z(n6749) );
  ANDN U14790 ( .B(n6769), .A(n6770), .Z(n6743) );
  XNOR U14791 ( .A(n6736), .B(n6771), .Z(n6742) );
  XNOR U14792 ( .A(n6735), .B(n6737), .Z(n6771) );
  NAND U14793 ( .A(n6772), .B(n6773), .Z(n6737) );
  OR U14794 ( .A(n6774), .B(n6775), .Z(n6773) );
  OR U14795 ( .A(n6776), .B(n6777), .Z(n6772) );
  NAND U14796 ( .A(n6778), .B(n6779), .Z(n6735) );
  OR U14797 ( .A(n6780), .B(n6781), .Z(n6779) );
  OR U14798 ( .A(n6782), .B(n6783), .Z(n6778) );
  ANDN U14799 ( .B(n6784), .A(n6785), .Z(n6736) );
  IV U14800 ( .A(n6786), .Z(n6784) );
  ANDN U14801 ( .B(n6787), .A(n6788), .Z(n6728) );
  XOR U14802 ( .A(n6714), .B(n6789), .Z(n6726) );
  XOR U14803 ( .A(n6715), .B(n6716), .Z(n6789) );
  XOR U14804 ( .A(n6721), .B(n6790), .Z(n6716) );
  XOR U14805 ( .A(n6720), .B(n6723), .Z(n6790) );
  IV U14806 ( .A(n6722), .Z(n6723) );
  NAND U14807 ( .A(n6791), .B(n6792), .Z(n6722) );
  OR U14808 ( .A(n6793), .B(n6794), .Z(n6792) );
  OR U14809 ( .A(n6795), .B(n6796), .Z(n6791) );
  NAND U14810 ( .A(n6797), .B(n6798), .Z(n6720) );
  OR U14811 ( .A(n6799), .B(n6800), .Z(n6798) );
  OR U14812 ( .A(n6801), .B(n6802), .Z(n6797) );
  NOR U14813 ( .A(n6803), .B(n6804), .Z(n6721) );
  ANDN U14814 ( .B(n6805), .A(n6806), .Z(n6715) );
  IV U14815 ( .A(n6807), .Z(n6805) );
  XNOR U14816 ( .A(n6708), .B(n6808), .Z(n6714) );
  XNOR U14817 ( .A(n6707), .B(n6709), .Z(n6808) );
  NAND U14818 ( .A(n6809), .B(n6810), .Z(n6709) );
  OR U14819 ( .A(n6811), .B(n6812), .Z(n6810) );
  OR U14820 ( .A(n6813), .B(n6814), .Z(n6809) );
  NAND U14821 ( .A(n6815), .B(n6816), .Z(n6707) );
  OR U14822 ( .A(n6817), .B(n6818), .Z(n6816) );
  OR U14823 ( .A(n6819), .B(n6820), .Z(n6815) );
  ANDN U14824 ( .B(n6821), .A(n6822), .Z(n6708) );
  IV U14825 ( .A(n6823), .Z(n6821) );
  XNOR U14826 ( .A(n6788), .B(n6787), .Z(N64791) );
  XOR U14827 ( .A(n6807), .B(n6806), .Z(n6787) );
  XNOR U14828 ( .A(n6822), .B(n6823), .Z(n6806) );
  XNOR U14829 ( .A(n6817), .B(n6818), .Z(n6823) );
  XNOR U14830 ( .A(n6819), .B(n6820), .Z(n6818) );
  XNOR U14831 ( .A(y[7765]), .B(x[7765]), .Z(n6820) );
  XNOR U14832 ( .A(y[7766]), .B(x[7766]), .Z(n6819) );
  XNOR U14833 ( .A(y[7764]), .B(x[7764]), .Z(n6817) );
  XNOR U14834 ( .A(n6811), .B(n6812), .Z(n6822) );
  XNOR U14835 ( .A(y[7761]), .B(x[7761]), .Z(n6812) );
  XNOR U14836 ( .A(n6813), .B(n6814), .Z(n6811) );
  XNOR U14837 ( .A(y[7762]), .B(x[7762]), .Z(n6814) );
  XNOR U14838 ( .A(y[7763]), .B(x[7763]), .Z(n6813) );
  XNOR U14839 ( .A(n6804), .B(n6803), .Z(n6807) );
  XNOR U14840 ( .A(n6799), .B(n6800), .Z(n6803) );
  XNOR U14841 ( .A(y[7758]), .B(x[7758]), .Z(n6800) );
  XNOR U14842 ( .A(n6801), .B(n6802), .Z(n6799) );
  XNOR U14843 ( .A(y[7759]), .B(x[7759]), .Z(n6802) );
  XNOR U14844 ( .A(y[7760]), .B(x[7760]), .Z(n6801) );
  XNOR U14845 ( .A(n6793), .B(n6794), .Z(n6804) );
  XNOR U14846 ( .A(y[7755]), .B(x[7755]), .Z(n6794) );
  XNOR U14847 ( .A(n6795), .B(n6796), .Z(n6793) );
  XNOR U14848 ( .A(y[7756]), .B(x[7756]), .Z(n6796) );
  XNOR U14849 ( .A(y[7757]), .B(x[7757]), .Z(n6795) );
  XOR U14850 ( .A(n6769), .B(n6770), .Z(n6788) );
  XNOR U14851 ( .A(n6785), .B(n6786), .Z(n6770) );
  XNOR U14852 ( .A(n6780), .B(n6781), .Z(n6786) );
  XNOR U14853 ( .A(n6782), .B(n6783), .Z(n6781) );
  XNOR U14854 ( .A(y[7753]), .B(x[7753]), .Z(n6783) );
  XNOR U14855 ( .A(y[7754]), .B(x[7754]), .Z(n6782) );
  XNOR U14856 ( .A(y[7752]), .B(x[7752]), .Z(n6780) );
  XNOR U14857 ( .A(n6774), .B(n6775), .Z(n6785) );
  XNOR U14858 ( .A(y[7749]), .B(x[7749]), .Z(n6775) );
  XNOR U14859 ( .A(n6776), .B(n6777), .Z(n6774) );
  XNOR U14860 ( .A(y[7750]), .B(x[7750]), .Z(n6777) );
  XNOR U14861 ( .A(y[7751]), .B(x[7751]), .Z(n6776) );
  XOR U14862 ( .A(n6768), .B(n6767), .Z(n6769) );
  XNOR U14863 ( .A(n6763), .B(n6764), .Z(n6767) );
  XNOR U14864 ( .A(y[7746]), .B(x[7746]), .Z(n6764) );
  XNOR U14865 ( .A(n6765), .B(n6766), .Z(n6763) );
  XNOR U14866 ( .A(y[7747]), .B(x[7747]), .Z(n6766) );
  XNOR U14867 ( .A(y[7748]), .B(x[7748]), .Z(n6765) );
  XNOR U14868 ( .A(n6757), .B(n6758), .Z(n6768) );
  XNOR U14869 ( .A(y[7743]), .B(x[7743]), .Z(n6758) );
  XNOR U14870 ( .A(n6759), .B(n6760), .Z(n6757) );
  XNOR U14871 ( .A(y[7744]), .B(x[7744]), .Z(n6760) );
  XNOR U14872 ( .A(y[7745]), .B(x[7745]), .Z(n6759) );
  NAND U14873 ( .A(n6824), .B(n6825), .Z(N64782) );
  NANDN U14874 ( .A(n6826), .B(n6827), .Z(n6825) );
  OR U14875 ( .A(n6828), .B(n6829), .Z(n6827) );
  NAND U14876 ( .A(n6828), .B(n6829), .Z(n6824) );
  XOR U14877 ( .A(n6828), .B(n6830), .Z(N64781) );
  XNOR U14878 ( .A(n6826), .B(n6829), .Z(n6830) );
  AND U14879 ( .A(n6831), .B(n6832), .Z(n6829) );
  NANDN U14880 ( .A(n6833), .B(n6834), .Z(n6832) );
  NANDN U14881 ( .A(n6835), .B(n6836), .Z(n6834) );
  NANDN U14882 ( .A(n6836), .B(n6835), .Z(n6831) );
  NAND U14883 ( .A(n6837), .B(n6838), .Z(n6826) );
  NANDN U14884 ( .A(n6839), .B(n6840), .Z(n6838) );
  OR U14885 ( .A(n6841), .B(n6842), .Z(n6840) );
  NAND U14886 ( .A(n6842), .B(n6841), .Z(n6837) );
  AND U14887 ( .A(n6843), .B(n6844), .Z(n6828) );
  NANDN U14888 ( .A(n6845), .B(n6846), .Z(n6844) );
  NANDN U14889 ( .A(n6847), .B(n6848), .Z(n6846) );
  NANDN U14890 ( .A(n6848), .B(n6847), .Z(n6843) );
  XOR U14891 ( .A(n6842), .B(n6849), .Z(N64780) );
  XOR U14892 ( .A(n6839), .B(n6841), .Z(n6849) );
  XNOR U14893 ( .A(n6835), .B(n6850), .Z(n6841) );
  XNOR U14894 ( .A(n6833), .B(n6836), .Z(n6850) );
  NAND U14895 ( .A(n6851), .B(n6852), .Z(n6836) );
  NAND U14896 ( .A(n6853), .B(n6854), .Z(n6852) );
  OR U14897 ( .A(n6855), .B(n6856), .Z(n6853) );
  NANDN U14898 ( .A(n6857), .B(n6855), .Z(n6851) );
  IV U14899 ( .A(n6856), .Z(n6857) );
  NAND U14900 ( .A(n6858), .B(n6859), .Z(n6833) );
  NAND U14901 ( .A(n6860), .B(n6861), .Z(n6859) );
  NANDN U14902 ( .A(n6862), .B(n6863), .Z(n6860) );
  NANDN U14903 ( .A(n6863), .B(n6862), .Z(n6858) );
  AND U14904 ( .A(n6864), .B(n6865), .Z(n6835) );
  NAND U14905 ( .A(n6866), .B(n6867), .Z(n6865) );
  OR U14906 ( .A(n6868), .B(n6869), .Z(n6866) );
  NANDN U14907 ( .A(n6870), .B(n6868), .Z(n6864) );
  NAND U14908 ( .A(n6871), .B(n6872), .Z(n6839) );
  NANDN U14909 ( .A(n6873), .B(n6874), .Z(n6872) );
  OR U14910 ( .A(n6875), .B(n6876), .Z(n6874) );
  NANDN U14911 ( .A(n6877), .B(n6875), .Z(n6871) );
  IV U14912 ( .A(n6876), .Z(n6877) );
  XNOR U14913 ( .A(n6847), .B(n6878), .Z(n6842) );
  XNOR U14914 ( .A(n6845), .B(n6848), .Z(n6878) );
  NAND U14915 ( .A(n6879), .B(n6880), .Z(n6848) );
  NAND U14916 ( .A(n6881), .B(n6882), .Z(n6880) );
  OR U14917 ( .A(n6883), .B(n6884), .Z(n6881) );
  NANDN U14918 ( .A(n6885), .B(n6883), .Z(n6879) );
  IV U14919 ( .A(n6884), .Z(n6885) );
  NAND U14920 ( .A(n6886), .B(n6887), .Z(n6845) );
  NAND U14921 ( .A(n6888), .B(n6889), .Z(n6887) );
  NANDN U14922 ( .A(n6890), .B(n6891), .Z(n6888) );
  NANDN U14923 ( .A(n6891), .B(n6890), .Z(n6886) );
  AND U14924 ( .A(n6892), .B(n6893), .Z(n6847) );
  NAND U14925 ( .A(n6894), .B(n6895), .Z(n6893) );
  OR U14926 ( .A(n6896), .B(n6897), .Z(n6894) );
  NANDN U14927 ( .A(n6898), .B(n6896), .Z(n6892) );
  XNOR U14928 ( .A(n6873), .B(n6899), .Z(N64779) );
  XOR U14929 ( .A(n6875), .B(n6876), .Z(n6899) );
  XNOR U14930 ( .A(n6889), .B(n6900), .Z(n6876) );
  XOR U14931 ( .A(n6890), .B(n6891), .Z(n6900) );
  XOR U14932 ( .A(n6896), .B(n6901), .Z(n6891) );
  XOR U14933 ( .A(n6895), .B(n6898), .Z(n6901) );
  IV U14934 ( .A(n6897), .Z(n6898) );
  NAND U14935 ( .A(n6902), .B(n6903), .Z(n6897) );
  OR U14936 ( .A(n6904), .B(n6905), .Z(n6903) );
  OR U14937 ( .A(n6906), .B(n6907), .Z(n6902) );
  NAND U14938 ( .A(n6908), .B(n6909), .Z(n6895) );
  OR U14939 ( .A(n6910), .B(n6911), .Z(n6909) );
  OR U14940 ( .A(n6912), .B(n6913), .Z(n6908) );
  NOR U14941 ( .A(n6914), .B(n6915), .Z(n6896) );
  ANDN U14942 ( .B(n6916), .A(n6917), .Z(n6890) );
  XNOR U14943 ( .A(n6883), .B(n6918), .Z(n6889) );
  XNOR U14944 ( .A(n6882), .B(n6884), .Z(n6918) );
  NAND U14945 ( .A(n6919), .B(n6920), .Z(n6884) );
  OR U14946 ( .A(n6921), .B(n6922), .Z(n6920) );
  OR U14947 ( .A(n6923), .B(n6924), .Z(n6919) );
  NAND U14948 ( .A(n6925), .B(n6926), .Z(n6882) );
  OR U14949 ( .A(n6927), .B(n6928), .Z(n6926) );
  OR U14950 ( .A(n6929), .B(n6930), .Z(n6925) );
  ANDN U14951 ( .B(n6931), .A(n6932), .Z(n6883) );
  IV U14952 ( .A(n6933), .Z(n6931) );
  ANDN U14953 ( .B(n6934), .A(n6935), .Z(n6875) );
  XOR U14954 ( .A(n6861), .B(n6936), .Z(n6873) );
  XOR U14955 ( .A(n6862), .B(n6863), .Z(n6936) );
  XOR U14956 ( .A(n6868), .B(n6937), .Z(n6863) );
  XOR U14957 ( .A(n6867), .B(n6870), .Z(n6937) );
  IV U14958 ( .A(n6869), .Z(n6870) );
  NAND U14959 ( .A(n6938), .B(n6939), .Z(n6869) );
  OR U14960 ( .A(n6940), .B(n6941), .Z(n6939) );
  OR U14961 ( .A(n6942), .B(n6943), .Z(n6938) );
  NAND U14962 ( .A(n6944), .B(n6945), .Z(n6867) );
  OR U14963 ( .A(n6946), .B(n6947), .Z(n6945) );
  OR U14964 ( .A(n6948), .B(n6949), .Z(n6944) );
  NOR U14965 ( .A(n6950), .B(n6951), .Z(n6868) );
  ANDN U14966 ( .B(n6952), .A(n6953), .Z(n6862) );
  IV U14967 ( .A(n6954), .Z(n6952) );
  XNOR U14968 ( .A(n6855), .B(n6955), .Z(n6861) );
  XNOR U14969 ( .A(n6854), .B(n6856), .Z(n6955) );
  NAND U14970 ( .A(n6956), .B(n6957), .Z(n6856) );
  OR U14971 ( .A(n6958), .B(n6959), .Z(n6957) );
  OR U14972 ( .A(n6960), .B(n6961), .Z(n6956) );
  NAND U14973 ( .A(n6962), .B(n6963), .Z(n6854) );
  OR U14974 ( .A(n6964), .B(n6965), .Z(n6963) );
  OR U14975 ( .A(n6966), .B(n6967), .Z(n6962) );
  ANDN U14976 ( .B(n6968), .A(n6969), .Z(n6855) );
  IV U14977 ( .A(n6970), .Z(n6968) );
  XNOR U14978 ( .A(n6935), .B(n6934), .Z(N64778) );
  XOR U14979 ( .A(n6954), .B(n6953), .Z(n6934) );
  XNOR U14980 ( .A(n6969), .B(n6970), .Z(n6953) );
  XNOR U14981 ( .A(n6964), .B(n6965), .Z(n6970) );
  XNOR U14982 ( .A(n6966), .B(n6967), .Z(n6965) );
  XNOR U14983 ( .A(y[7741]), .B(x[7741]), .Z(n6967) );
  XNOR U14984 ( .A(y[7742]), .B(x[7742]), .Z(n6966) );
  XNOR U14985 ( .A(y[7740]), .B(x[7740]), .Z(n6964) );
  XNOR U14986 ( .A(n6958), .B(n6959), .Z(n6969) );
  XNOR U14987 ( .A(y[7737]), .B(x[7737]), .Z(n6959) );
  XNOR U14988 ( .A(n6960), .B(n6961), .Z(n6958) );
  XNOR U14989 ( .A(y[7738]), .B(x[7738]), .Z(n6961) );
  XNOR U14990 ( .A(y[7739]), .B(x[7739]), .Z(n6960) );
  XNOR U14991 ( .A(n6951), .B(n6950), .Z(n6954) );
  XNOR U14992 ( .A(n6946), .B(n6947), .Z(n6950) );
  XNOR U14993 ( .A(y[7734]), .B(x[7734]), .Z(n6947) );
  XNOR U14994 ( .A(n6948), .B(n6949), .Z(n6946) );
  XNOR U14995 ( .A(y[7735]), .B(x[7735]), .Z(n6949) );
  XNOR U14996 ( .A(y[7736]), .B(x[7736]), .Z(n6948) );
  XNOR U14997 ( .A(n6940), .B(n6941), .Z(n6951) );
  XNOR U14998 ( .A(y[7731]), .B(x[7731]), .Z(n6941) );
  XNOR U14999 ( .A(n6942), .B(n6943), .Z(n6940) );
  XNOR U15000 ( .A(y[7732]), .B(x[7732]), .Z(n6943) );
  XNOR U15001 ( .A(y[7733]), .B(x[7733]), .Z(n6942) );
  XOR U15002 ( .A(n6916), .B(n6917), .Z(n6935) );
  XNOR U15003 ( .A(n6932), .B(n6933), .Z(n6917) );
  XNOR U15004 ( .A(n6927), .B(n6928), .Z(n6933) );
  XNOR U15005 ( .A(n6929), .B(n6930), .Z(n6928) );
  XNOR U15006 ( .A(y[7729]), .B(x[7729]), .Z(n6930) );
  XNOR U15007 ( .A(y[7730]), .B(x[7730]), .Z(n6929) );
  XNOR U15008 ( .A(y[7728]), .B(x[7728]), .Z(n6927) );
  XNOR U15009 ( .A(n6921), .B(n6922), .Z(n6932) );
  XNOR U15010 ( .A(y[7725]), .B(x[7725]), .Z(n6922) );
  XNOR U15011 ( .A(n6923), .B(n6924), .Z(n6921) );
  XNOR U15012 ( .A(y[7726]), .B(x[7726]), .Z(n6924) );
  XNOR U15013 ( .A(y[7727]), .B(x[7727]), .Z(n6923) );
  XOR U15014 ( .A(n6915), .B(n6914), .Z(n6916) );
  XNOR U15015 ( .A(n6910), .B(n6911), .Z(n6914) );
  XNOR U15016 ( .A(y[7722]), .B(x[7722]), .Z(n6911) );
  XNOR U15017 ( .A(n6912), .B(n6913), .Z(n6910) );
  XNOR U15018 ( .A(y[7723]), .B(x[7723]), .Z(n6913) );
  XNOR U15019 ( .A(y[7724]), .B(x[7724]), .Z(n6912) );
  XNOR U15020 ( .A(n6904), .B(n6905), .Z(n6915) );
  XNOR U15021 ( .A(y[7719]), .B(x[7719]), .Z(n6905) );
  XNOR U15022 ( .A(n6906), .B(n6907), .Z(n6904) );
  XNOR U15023 ( .A(y[7720]), .B(x[7720]), .Z(n6907) );
  XNOR U15024 ( .A(y[7721]), .B(x[7721]), .Z(n6906) );
  NAND U15025 ( .A(n6971), .B(n6972), .Z(N64769) );
  NANDN U15026 ( .A(n6973), .B(n6974), .Z(n6972) );
  OR U15027 ( .A(n6975), .B(n6976), .Z(n6974) );
  NAND U15028 ( .A(n6975), .B(n6976), .Z(n6971) );
  XOR U15029 ( .A(n6975), .B(n6977), .Z(N64768) );
  XNOR U15030 ( .A(n6973), .B(n6976), .Z(n6977) );
  AND U15031 ( .A(n6978), .B(n6979), .Z(n6976) );
  NANDN U15032 ( .A(n6980), .B(n6981), .Z(n6979) );
  NANDN U15033 ( .A(n6982), .B(n6983), .Z(n6981) );
  NANDN U15034 ( .A(n6983), .B(n6982), .Z(n6978) );
  NAND U15035 ( .A(n6984), .B(n6985), .Z(n6973) );
  NANDN U15036 ( .A(n6986), .B(n6987), .Z(n6985) );
  OR U15037 ( .A(n6988), .B(n6989), .Z(n6987) );
  NAND U15038 ( .A(n6989), .B(n6988), .Z(n6984) );
  AND U15039 ( .A(n6990), .B(n6991), .Z(n6975) );
  NANDN U15040 ( .A(n6992), .B(n6993), .Z(n6991) );
  NANDN U15041 ( .A(n6994), .B(n6995), .Z(n6993) );
  NANDN U15042 ( .A(n6995), .B(n6994), .Z(n6990) );
  XOR U15043 ( .A(n6989), .B(n6996), .Z(N64767) );
  XOR U15044 ( .A(n6986), .B(n6988), .Z(n6996) );
  XNOR U15045 ( .A(n6982), .B(n6997), .Z(n6988) );
  XNOR U15046 ( .A(n6980), .B(n6983), .Z(n6997) );
  NAND U15047 ( .A(n6998), .B(n6999), .Z(n6983) );
  NAND U15048 ( .A(n7000), .B(n7001), .Z(n6999) );
  OR U15049 ( .A(n7002), .B(n7003), .Z(n7000) );
  NANDN U15050 ( .A(n7004), .B(n7002), .Z(n6998) );
  IV U15051 ( .A(n7003), .Z(n7004) );
  NAND U15052 ( .A(n7005), .B(n7006), .Z(n6980) );
  NAND U15053 ( .A(n7007), .B(n7008), .Z(n7006) );
  NANDN U15054 ( .A(n7009), .B(n7010), .Z(n7007) );
  NANDN U15055 ( .A(n7010), .B(n7009), .Z(n7005) );
  AND U15056 ( .A(n7011), .B(n7012), .Z(n6982) );
  NAND U15057 ( .A(n7013), .B(n7014), .Z(n7012) );
  OR U15058 ( .A(n7015), .B(n7016), .Z(n7013) );
  NANDN U15059 ( .A(n7017), .B(n7015), .Z(n7011) );
  NAND U15060 ( .A(n7018), .B(n7019), .Z(n6986) );
  NANDN U15061 ( .A(n7020), .B(n7021), .Z(n7019) );
  OR U15062 ( .A(n7022), .B(n7023), .Z(n7021) );
  NANDN U15063 ( .A(n7024), .B(n7022), .Z(n7018) );
  IV U15064 ( .A(n7023), .Z(n7024) );
  XNOR U15065 ( .A(n6994), .B(n7025), .Z(n6989) );
  XNOR U15066 ( .A(n6992), .B(n6995), .Z(n7025) );
  NAND U15067 ( .A(n7026), .B(n7027), .Z(n6995) );
  NAND U15068 ( .A(n7028), .B(n7029), .Z(n7027) );
  OR U15069 ( .A(n7030), .B(n7031), .Z(n7028) );
  NANDN U15070 ( .A(n7032), .B(n7030), .Z(n7026) );
  IV U15071 ( .A(n7031), .Z(n7032) );
  NAND U15072 ( .A(n7033), .B(n7034), .Z(n6992) );
  NAND U15073 ( .A(n7035), .B(n7036), .Z(n7034) );
  NANDN U15074 ( .A(n7037), .B(n7038), .Z(n7035) );
  NANDN U15075 ( .A(n7038), .B(n7037), .Z(n7033) );
  AND U15076 ( .A(n7039), .B(n7040), .Z(n6994) );
  NAND U15077 ( .A(n7041), .B(n7042), .Z(n7040) );
  OR U15078 ( .A(n7043), .B(n7044), .Z(n7041) );
  NANDN U15079 ( .A(n7045), .B(n7043), .Z(n7039) );
  XNOR U15080 ( .A(n7020), .B(n7046), .Z(N64766) );
  XOR U15081 ( .A(n7022), .B(n7023), .Z(n7046) );
  XNOR U15082 ( .A(n7036), .B(n7047), .Z(n7023) );
  XOR U15083 ( .A(n7037), .B(n7038), .Z(n7047) );
  XOR U15084 ( .A(n7043), .B(n7048), .Z(n7038) );
  XOR U15085 ( .A(n7042), .B(n7045), .Z(n7048) );
  IV U15086 ( .A(n7044), .Z(n7045) );
  NAND U15087 ( .A(n7049), .B(n7050), .Z(n7044) );
  OR U15088 ( .A(n7051), .B(n7052), .Z(n7050) );
  OR U15089 ( .A(n7053), .B(n7054), .Z(n7049) );
  NAND U15090 ( .A(n7055), .B(n7056), .Z(n7042) );
  OR U15091 ( .A(n7057), .B(n7058), .Z(n7056) );
  OR U15092 ( .A(n7059), .B(n7060), .Z(n7055) );
  NOR U15093 ( .A(n7061), .B(n7062), .Z(n7043) );
  ANDN U15094 ( .B(n7063), .A(n7064), .Z(n7037) );
  XNOR U15095 ( .A(n7030), .B(n7065), .Z(n7036) );
  XNOR U15096 ( .A(n7029), .B(n7031), .Z(n7065) );
  NAND U15097 ( .A(n7066), .B(n7067), .Z(n7031) );
  OR U15098 ( .A(n7068), .B(n7069), .Z(n7067) );
  OR U15099 ( .A(n7070), .B(n7071), .Z(n7066) );
  NAND U15100 ( .A(n7072), .B(n7073), .Z(n7029) );
  OR U15101 ( .A(n7074), .B(n7075), .Z(n7073) );
  OR U15102 ( .A(n7076), .B(n7077), .Z(n7072) );
  ANDN U15103 ( .B(n7078), .A(n7079), .Z(n7030) );
  IV U15104 ( .A(n7080), .Z(n7078) );
  ANDN U15105 ( .B(n7081), .A(n7082), .Z(n7022) );
  XOR U15106 ( .A(n7008), .B(n7083), .Z(n7020) );
  XOR U15107 ( .A(n7009), .B(n7010), .Z(n7083) );
  XOR U15108 ( .A(n7015), .B(n7084), .Z(n7010) );
  XOR U15109 ( .A(n7014), .B(n7017), .Z(n7084) );
  IV U15110 ( .A(n7016), .Z(n7017) );
  NAND U15111 ( .A(n7085), .B(n7086), .Z(n7016) );
  OR U15112 ( .A(n7087), .B(n7088), .Z(n7086) );
  OR U15113 ( .A(n7089), .B(n7090), .Z(n7085) );
  NAND U15114 ( .A(n7091), .B(n7092), .Z(n7014) );
  OR U15115 ( .A(n7093), .B(n7094), .Z(n7092) );
  OR U15116 ( .A(n7095), .B(n7096), .Z(n7091) );
  NOR U15117 ( .A(n7097), .B(n7098), .Z(n7015) );
  ANDN U15118 ( .B(n7099), .A(n7100), .Z(n7009) );
  IV U15119 ( .A(n7101), .Z(n7099) );
  XNOR U15120 ( .A(n7002), .B(n7102), .Z(n7008) );
  XNOR U15121 ( .A(n7001), .B(n7003), .Z(n7102) );
  NAND U15122 ( .A(n7103), .B(n7104), .Z(n7003) );
  OR U15123 ( .A(n7105), .B(n7106), .Z(n7104) );
  OR U15124 ( .A(n7107), .B(n7108), .Z(n7103) );
  NAND U15125 ( .A(n7109), .B(n7110), .Z(n7001) );
  OR U15126 ( .A(n7111), .B(n7112), .Z(n7110) );
  OR U15127 ( .A(n7113), .B(n7114), .Z(n7109) );
  ANDN U15128 ( .B(n7115), .A(n7116), .Z(n7002) );
  IV U15129 ( .A(n7117), .Z(n7115) );
  XNOR U15130 ( .A(n7082), .B(n7081), .Z(N64765) );
  XOR U15131 ( .A(n7101), .B(n7100), .Z(n7081) );
  XNOR U15132 ( .A(n7116), .B(n7117), .Z(n7100) );
  XNOR U15133 ( .A(n7111), .B(n7112), .Z(n7117) );
  XNOR U15134 ( .A(n7113), .B(n7114), .Z(n7112) );
  XNOR U15135 ( .A(y[7717]), .B(x[7717]), .Z(n7114) );
  XNOR U15136 ( .A(y[7718]), .B(x[7718]), .Z(n7113) );
  XNOR U15137 ( .A(y[7716]), .B(x[7716]), .Z(n7111) );
  XNOR U15138 ( .A(n7105), .B(n7106), .Z(n7116) );
  XNOR U15139 ( .A(y[7713]), .B(x[7713]), .Z(n7106) );
  XNOR U15140 ( .A(n7107), .B(n7108), .Z(n7105) );
  XNOR U15141 ( .A(y[7714]), .B(x[7714]), .Z(n7108) );
  XNOR U15142 ( .A(y[7715]), .B(x[7715]), .Z(n7107) );
  XNOR U15143 ( .A(n7098), .B(n7097), .Z(n7101) );
  XNOR U15144 ( .A(n7093), .B(n7094), .Z(n7097) );
  XNOR U15145 ( .A(y[7710]), .B(x[7710]), .Z(n7094) );
  XNOR U15146 ( .A(n7095), .B(n7096), .Z(n7093) );
  XNOR U15147 ( .A(y[7711]), .B(x[7711]), .Z(n7096) );
  XNOR U15148 ( .A(y[7712]), .B(x[7712]), .Z(n7095) );
  XNOR U15149 ( .A(n7087), .B(n7088), .Z(n7098) );
  XNOR U15150 ( .A(y[7707]), .B(x[7707]), .Z(n7088) );
  XNOR U15151 ( .A(n7089), .B(n7090), .Z(n7087) );
  XNOR U15152 ( .A(y[7708]), .B(x[7708]), .Z(n7090) );
  XNOR U15153 ( .A(y[7709]), .B(x[7709]), .Z(n7089) );
  XOR U15154 ( .A(n7063), .B(n7064), .Z(n7082) );
  XNOR U15155 ( .A(n7079), .B(n7080), .Z(n7064) );
  XNOR U15156 ( .A(n7074), .B(n7075), .Z(n7080) );
  XNOR U15157 ( .A(n7076), .B(n7077), .Z(n7075) );
  XNOR U15158 ( .A(y[7705]), .B(x[7705]), .Z(n7077) );
  XNOR U15159 ( .A(y[7706]), .B(x[7706]), .Z(n7076) );
  XNOR U15160 ( .A(y[7704]), .B(x[7704]), .Z(n7074) );
  XNOR U15161 ( .A(n7068), .B(n7069), .Z(n7079) );
  XNOR U15162 ( .A(y[7701]), .B(x[7701]), .Z(n7069) );
  XNOR U15163 ( .A(n7070), .B(n7071), .Z(n7068) );
  XNOR U15164 ( .A(y[7702]), .B(x[7702]), .Z(n7071) );
  XNOR U15165 ( .A(y[7703]), .B(x[7703]), .Z(n7070) );
  XOR U15166 ( .A(n7062), .B(n7061), .Z(n7063) );
  XNOR U15167 ( .A(n7057), .B(n7058), .Z(n7061) );
  XNOR U15168 ( .A(y[7698]), .B(x[7698]), .Z(n7058) );
  XNOR U15169 ( .A(n7059), .B(n7060), .Z(n7057) );
  XNOR U15170 ( .A(y[7699]), .B(x[7699]), .Z(n7060) );
  XNOR U15171 ( .A(y[7700]), .B(x[7700]), .Z(n7059) );
  XNOR U15172 ( .A(n7051), .B(n7052), .Z(n7062) );
  XNOR U15173 ( .A(y[7695]), .B(x[7695]), .Z(n7052) );
  XNOR U15174 ( .A(n7053), .B(n7054), .Z(n7051) );
  XNOR U15175 ( .A(y[7696]), .B(x[7696]), .Z(n7054) );
  XNOR U15176 ( .A(y[7697]), .B(x[7697]), .Z(n7053) );
  NAND U15177 ( .A(n7118), .B(n7119), .Z(N64756) );
  NANDN U15178 ( .A(n7120), .B(n7121), .Z(n7119) );
  OR U15179 ( .A(n7122), .B(n7123), .Z(n7121) );
  NAND U15180 ( .A(n7122), .B(n7123), .Z(n7118) );
  XOR U15181 ( .A(n7122), .B(n7124), .Z(N64755) );
  XNOR U15182 ( .A(n7120), .B(n7123), .Z(n7124) );
  AND U15183 ( .A(n7125), .B(n7126), .Z(n7123) );
  NANDN U15184 ( .A(n7127), .B(n7128), .Z(n7126) );
  NANDN U15185 ( .A(n7129), .B(n7130), .Z(n7128) );
  NANDN U15186 ( .A(n7130), .B(n7129), .Z(n7125) );
  NAND U15187 ( .A(n7131), .B(n7132), .Z(n7120) );
  NANDN U15188 ( .A(n7133), .B(n7134), .Z(n7132) );
  OR U15189 ( .A(n7135), .B(n7136), .Z(n7134) );
  NAND U15190 ( .A(n7136), .B(n7135), .Z(n7131) );
  AND U15191 ( .A(n7137), .B(n7138), .Z(n7122) );
  NANDN U15192 ( .A(n7139), .B(n7140), .Z(n7138) );
  NANDN U15193 ( .A(n7141), .B(n7142), .Z(n7140) );
  NANDN U15194 ( .A(n7142), .B(n7141), .Z(n7137) );
  XOR U15195 ( .A(n7136), .B(n7143), .Z(N64754) );
  XOR U15196 ( .A(n7133), .B(n7135), .Z(n7143) );
  XNOR U15197 ( .A(n7129), .B(n7144), .Z(n7135) );
  XNOR U15198 ( .A(n7127), .B(n7130), .Z(n7144) );
  NAND U15199 ( .A(n7145), .B(n7146), .Z(n7130) );
  NAND U15200 ( .A(n7147), .B(n7148), .Z(n7146) );
  OR U15201 ( .A(n7149), .B(n7150), .Z(n7147) );
  NANDN U15202 ( .A(n7151), .B(n7149), .Z(n7145) );
  IV U15203 ( .A(n7150), .Z(n7151) );
  NAND U15204 ( .A(n7152), .B(n7153), .Z(n7127) );
  NAND U15205 ( .A(n7154), .B(n7155), .Z(n7153) );
  NANDN U15206 ( .A(n7156), .B(n7157), .Z(n7154) );
  NANDN U15207 ( .A(n7157), .B(n7156), .Z(n7152) );
  AND U15208 ( .A(n7158), .B(n7159), .Z(n7129) );
  NAND U15209 ( .A(n7160), .B(n7161), .Z(n7159) );
  OR U15210 ( .A(n7162), .B(n7163), .Z(n7160) );
  NANDN U15211 ( .A(n7164), .B(n7162), .Z(n7158) );
  NAND U15212 ( .A(n7165), .B(n7166), .Z(n7133) );
  NANDN U15213 ( .A(n7167), .B(n7168), .Z(n7166) );
  OR U15214 ( .A(n7169), .B(n7170), .Z(n7168) );
  NANDN U15215 ( .A(n7171), .B(n7169), .Z(n7165) );
  IV U15216 ( .A(n7170), .Z(n7171) );
  XNOR U15217 ( .A(n7141), .B(n7172), .Z(n7136) );
  XNOR U15218 ( .A(n7139), .B(n7142), .Z(n7172) );
  NAND U15219 ( .A(n7173), .B(n7174), .Z(n7142) );
  NAND U15220 ( .A(n7175), .B(n7176), .Z(n7174) );
  OR U15221 ( .A(n7177), .B(n7178), .Z(n7175) );
  NANDN U15222 ( .A(n7179), .B(n7177), .Z(n7173) );
  IV U15223 ( .A(n7178), .Z(n7179) );
  NAND U15224 ( .A(n7180), .B(n7181), .Z(n7139) );
  NAND U15225 ( .A(n7182), .B(n7183), .Z(n7181) );
  NANDN U15226 ( .A(n7184), .B(n7185), .Z(n7182) );
  NANDN U15227 ( .A(n7185), .B(n7184), .Z(n7180) );
  AND U15228 ( .A(n7186), .B(n7187), .Z(n7141) );
  NAND U15229 ( .A(n7188), .B(n7189), .Z(n7187) );
  OR U15230 ( .A(n7190), .B(n7191), .Z(n7188) );
  NANDN U15231 ( .A(n7192), .B(n7190), .Z(n7186) );
  XNOR U15232 ( .A(n7167), .B(n7193), .Z(N64753) );
  XOR U15233 ( .A(n7169), .B(n7170), .Z(n7193) );
  XNOR U15234 ( .A(n7183), .B(n7194), .Z(n7170) );
  XOR U15235 ( .A(n7184), .B(n7185), .Z(n7194) );
  XOR U15236 ( .A(n7190), .B(n7195), .Z(n7185) );
  XOR U15237 ( .A(n7189), .B(n7192), .Z(n7195) );
  IV U15238 ( .A(n7191), .Z(n7192) );
  NAND U15239 ( .A(n7196), .B(n7197), .Z(n7191) );
  OR U15240 ( .A(n7198), .B(n7199), .Z(n7197) );
  OR U15241 ( .A(n7200), .B(n7201), .Z(n7196) );
  NAND U15242 ( .A(n7202), .B(n7203), .Z(n7189) );
  OR U15243 ( .A(n7204), .B(n7205), .Z(n7203) );
  OR U15244 ( .A(n7206), .B(n7207), .Z(n7202) );
  NOR U15245 ( .A(n7208), .B(n7209), .Z(n7190) );
  ANDN U15246 ( .B(n7210), .A(n7211), .Z(n7184) );
  XNOR U15247 ( .A(n7177), .B(n7212), .Z(n7183) );
  XNOR U15248 ( .A(n7176), .B(n7178), .Z(n7212) );
  NAND U15249 ( .A(n7213), .B(n7214), .Z(n7178) );
  OR U15250 ( .A(n7215), .B(n7216), .Z(n7214) );
  OR U15251 ( .A(n7217), .B(n7218), .Z(n7213) );
  NAND U15252 ( .A(n7219), .B(n7220), .Z(n7176) );
  OR U15253 ( .A(n7221), .B(n7222), .Z(n7220) );
  OR U15254 ( .A(n7223), .B(n7224), .Z(n7219) );
  ANDN U15255 ( .B(n7225), .A(n7226), .Z(n7177) );
  IV U15256 ( .A(n7227), .Z(n7225) );
  ANDN U15257 ( .B(n7228), .A(n7229), .Z(n7169) );
  XOR U15258 ( .A(n7155), .B(n7230), .Z(n7167) );
  XOR U15259 ( .A(n7156), .B(n7157), .Z(n7230) );
  XOR U15260 ( .A(n7162), .B(n7231), .Z(n7157) );
  XOR U15261 ( .A(n7161), .B(n7164), .Z(n7231) );
  IV U15262 ( .A(n7163), .Z(n7164) );
  NAND U15263 ( .A(n7232), .B(n7233), .Z(n7163) );
  OR U15264 ( .A(n7234), .B(n7235), .Z(n7233) );
  OR U15265 ( .A(n7236), .B(n7237), .Z(n7232) );
  NAND U15266 ( .A(n7238), .B(n7239), .Z(n7161) );
  OR U15267 ( .A(n7240), .B(n7241), .Z(n7239) );
  OR U15268 ( .A(n7242), .B(n7243), .Z(n7238) );
  NOR U15269 ( .A(n7244), .B(n7245), .Z(n7162) );
  ANDN U15270 ( .B(n7246), .A(n7247), .Z(n7156) );
  IV U15271 ( .A(n7248), .Z(n7246) );
  XNOR U15272 ( .A(n7149), .B(n7249), .Z(n7155) );
  XNOR U15273 ( .A(n7148), .B(n7150), .Z(n7249) );
  NAND U15274 ( .A(n7250), .B(n7251), .Z(n7150) );
  OR U15275 ( .A(n7252), .B(n7253), .Z(n7251) );
  OR U15276 ( .A(n7254), .B(n7255), .Z(n7250) );
  NAND U15277 ( .A(n7256), .B(n7257), .Z(n7148) );
  OR U15278 ( .A(n7258), .B(n7259), .Z(n7257) );
  OR U15279 ( .A(n7260), .B(n7261), .Z(n7256) );
  ANDN U15280 ( .B(n7262), .A(n7263), .Z(n7149) );
  IV U15281 ( .A(n7264), .Z(n7262) );
  XNOR U15282 ( .A(n7229), .B(n7228), .Z(N64752) );
  XOR U15283 ( .A(n7248), .B(n7247), .Z(n7228) );
  XNOR U15284 ( .A(n7263), .B(n7264), .Z(n7247) );
  XNOR U15285 ( .A(n7258), .B(n7259), .Z(n7264) );
  XNOR U15286 ( .A(n7260), .B(n7261), .Z(n7259) );
  XNOR U15287 ( .A(y[7693]), .B(x[7693]), .Z(n7261) );
  XNOR U15288 ( .A(y[7694]), .B(x[7694]), .Z(n7260) );
  XNOR U15289 ( .A(y[7692]), .B(x[7692]), .Z(n7258) );
  XNOR U15290 ( .A(n7252), .B(n7253), .Z(n7263) );
  XNOR U15291 ( .A(y[7689]), .B(x[7689]), .Z(n7253) );
  XNOR U15292 ( .A(n7254), .B(n7255), .Z(n7252) );
  XNOR U15293 ( .A(y[7690]), .B(x[7690]), .Z(n7255) );
  XNOR U15294 ( .A(y[7691]), .B(x[7691]), .Z(n7254) );
  XNOR U15295 ( .A(n7245), .B(n7244), .Z(n7248) );
  XNOR U15296 ( .A(n7240), .B(n7241), .Z(n7244) );
  XNOR U15297 ( .A(y[7686]), .B(x[7686]), .Z(n7241) );
  XNOR U15298 ( .A(n7242), .B(n7243), .Z(n7240) );
  XNOR U15299 ( .A(y[7687]), .B(x[7687]), .Z(n7243) );
  XNOR U15300 ( .A(y[7688]), .B(x[7688]), .Z(n7242) );
  XNOR U15301 ( .A(n7234), .B(n7235), .Z(n7245) );
  XNOR U15302 ( .A(y[7683]), .B(x[7683]), .Z(n7235) );
  XNOR U15303 ( .A(n7236), .B(n7237), .Z(n7234) );
  XNOR U15304 ( .A(y[7684]), .B(x[7684]), .Z(n7237) );
  XNOR U15305 ( .A(y[7685]), .B(x[7685]), .Z(n7236) );
  XOR U15306 ( .A(n7210), .B(n7211), .Z(n7229) );
  XNOR U15307 ( .A(n7226), .B(n7227), .Z(n7211) );
  XNOR U15308 ( .A(n7221), .B(n7222), .Z(n7227) );
  XNOR U15309 ( .A(n7223), .B(n7224), .Z(n7222) );
  XNOR U15310 ( .A(y[7681]), .B(x[7681]), .Z(n7224) );
  XNOR U15311 ( .A(y[7682]), .B(x[7682]), .Z(n7223) );
  XNOR U15312 ( .A(y[7680]), .B(x[7680]), .Z(n7221) );
  XNOR U15313 ( .A(n7215), .B(n7216), .Z(n7226) );
  XNOR U15314 ( .A(y[7677]), .B(x[7677]), .Z(n7216) );
  XNOR U15315 ( .A(n7217), .B(n7218), .Z(n7215) );
  XNOR U15316 ( .A(y[7678]), .B(x[7678]), .Z(n7218) );
  XNOR U15317 ( .A(y[7679]), .B(x[7679]), .Z(n7217) );
  XOR U15318 ( .A(n7209), .B(n7208), .Z(n7210) );
  XNOR U15319 ( .A(n7204), .B(n7205), .Z(n7208) );
  XNOR U15320 ( .A(y[7674]), .B(x[7674]), .Z(n7205) );
  XNOR U15321 ( .A(n7206), .B(n7207), .Z(n7204) );
  XNOR U15322 ( .A(y[7675]), .B(x[7675]), .Z(n7207) );
  XNOR U15323 ( .A(y[7676]), .B(x[7676]), .Z(n7206) );
  XNOR U15324 ( .A(n7198), .B(n7199), .Z(n7209) );
  XNOR U15325 ( .A(y[7671]), .B(x[7671]), .Z(n7199) );
  XNOR U15326 ( .A(n7200), .B(n7201), .Z(n7198) );
  XNOR U15327 ( .A(y[7672]), .B(x[7672]), .Z(n7201) );
  XNOR U15328 ( .A(y[7673]), .B(x[7673]), .Z(n7200) );
  NAND U15329 ( .A(n7265), .B(n7266), .Z(N64743) );
  NANDN U15330 ( .A(n7267), .B(n7268), .Z(n7266) );
  OR U15331 ( .A(n7269), .B(n7270), .Z(n7268) );
  NAND U15332 ( .A(n7269), .B(n7270), .Z(n7265) );
  XOR U15333 ( .A(n7269), .B(n7271), .Z(N64742) );
  XNOR U15334 ( .A(n7267), .B(n7270), .Z(n7271) );
  AND U15335 ( .A(n7272), .B(n7273), .Z(n7270) );
  NANDN U15336 ( .A(n7274), .B(n7275), .Z(n7273) );
  NANDN U15337 ( .A(n7276), .B(n7277), .Z(n7275) );
  NANDN U15338 ( .A(n7277), .B(n7276), .Z(n7272) );
  NAND U15339 ( .A(n7278), .B(n7279), .Z(n7267) );
  NANDN U15340 ( .A(n7280), .B(n7281), .Z(n7279) );
  OR U15341 ( .A(n7282), .B(n7283), .Z(n7281) );
  NAND U15342 ( .A(n7283), .B(n7282), .Z(n7278) );
  AND U15343 ( .A(n7284), .B(n7285), .Z(n7269) );
  NANDN U15344 ( .A(n7286), .B(n7287), .Z(n7285) );
  NANDN U15345 ( .A(n7288), .B(n7289), .Z(n7287) );
  NANDN U15346 ( .A(n7289), .B(n7288), .Z(n7284) );
  XOR U15347 ( .A(n7283), .B(n7290), .Z(N64741) );
  XOR U15348 ( .A(n7280), .B(n7282), .Z(n7290) );
  XNOR U15349 ( .A(n7276), .B(n7291), .Z(n7282) );
  XNOR U15350 ( .A(n7274), .B(n7277), .Z(n7291) );
  NAND U15351 ( .A(n7292), .B(n7293), .Z(n7277) );
  NAND U15352 ( .A(n7294), .B(n7295), .Z(n7293) );
  OR U15353 ( .A(n7296), .B(n7297), .Z(n7294) );
  NANDN U15354 ( .A(n7298), .B(n7296), .Z(n7292) );
  IV U15355 ( .A(n7297), .Z(n7298) );
  NAND U15356 ( .A(n7299), .B(n7300), .Z(n7274) );
  NAND U15357 ( .A(n7301), .B(n7302), .Z(n7300) );
  NANDN U15358 ( .A(n7303), .B(n7304), .Z(n7301) );
  NANDN U15359 ( .A(n7304), .B(n7303), .Z(n7299) );
  AND U15360 ( .A(n7305), .B(n7306), .Z(n7276) );
  NAND U15361 ( .A(n7307), .B(n7308), .Z(n7306) );
  OR U15362 ( .A(n7309), .B(n7310), .Z(n7307) );
  NANDN U15363 ( .A(n7311), .B(n7309), .Z(n7305) );
  NAND U15364 ( .A(n7312), .B(n7313), .Z(n7280) );
  NANDN U15365 ( .A(n7314), .B(n7315), .Z(n7313) );
  OR U15366 ( .A(n7316), .B(n7317), .Z(n7315) );
  NANDN U15367 ( .A(n7318), .B(n7316), .Z(n7312) );
  IV U15368 ( .A(n7317), .Z(n7318) );
  XNOR U15369 ( .A(n7288), .B(n7319), .Z(n7283) );
  XNOR U15370 ( .A(n7286), .B(n7289), .Z(n7319) );
  NAND U15371 ( .A(n7320), .B(n7321), .Z(n7289) );
  NAND U15372 ( .A(n7322), .B(n7323), .Z(n7321) );
  OR U15373 ( .A(n7324), .B(n7325), .Z(n7322) );
  NANDN U15374 ( .A(n7326), .B(n7324), .Z(n7320) );
  IV U15375 ( .A(n7325), .Z(n7326) );
  NAND U15376 ( .A(n7327), .B(n7328), .Z(n7286) );
  NAND U15377 ( .A(n7329), .B(n7330), .Z(n7328) );
  NANDN U15378 ( .A(n7331), .B(n7332), .Z(n7329) );
  NANDN U15379 ( .A(n7332), .B(n7331), .Z(n7327) );
  AND U15380 ( .A(n7333), .B(n7334), .Z(n7288) );
  NAND U15381 ( .A(n7335), .B(n7336), .Z(n7334) );
  OR U15382 ( .A(n7337), .B(n7338), .Z(n7335) );
  NANDN U15383 ( .A(n7339), .B(n7337), .Z(n7333) );
  XNOR U15384 ( .A(n7314), .B(n7340), .Z(N64740) );
  XOR U15385 ( .A(n7316), .B(n7317), .Z(n7340) );
  XNOR U15386 ( .A(n7330), .B(n7341), .Z(n7317) );
  XOR U15387 ( .A(n7331), .B(n7332), .Z(n7341) );
  XOR U15388 ( .A(n7337), .B(n7342), .Z(n7332) );
  XOR U15389 ( .A(n7336), .B(n7339), .Z(n7342) );
  IV U15390 ( .A(n7338), .Z(n7339) );
  NAND U15391 ( .A(n7343), .B(n7344), .Z(n7338) );
  OR U15392 ( .A(n7345), .B(n7346), .Z(n7344) );
  OR U15393 ( .A(n7347), .B(n7348), .Z(n7343) );
  NAND U15394 ( .A(n7349), .B(n7350), .Z(n7336) );
  OR U15395 ( .A(n7351), .B(n7352), .Z(n7350) );
  OR U15396 ( .A(n7353), .B(n7354), .Z(n7349) );
  NOR U15397 ( .A(n7355), .B(n7356), .Z(n7337) );
  ANDN U15398 ( .B(n7357), .A(n7358), .Z(n7331) );
  XNOR U15399 ( .A(n7324), .B(n7359), .Z(n7330) );
  XNOR U15400 ( .A(n7323), .B(n7325), .Z(n7359) );
  NAND U15401 ( .A(n7360), .B(n7361), .Z(n7325) );
  OR U15402 ( .A(n7362), .B(n7363), .Z(n7361) );
  OR U15403 ( .A(n7364), .B(n7365), .Z(n7360) );
  NAND U15404 ( .A(n7366), .B(n7367), .Z(n7323) );
  OR U15405 ( .A(n7368), .B(n7369), .Z(n7367) );
  OR U15406 ( .A(n7370), .B(n7371), .Z(n7366) );
  ANDN U15407 ( .B(n7372), .A(n7373), .Z(n7324) );
  IV U15408 ( .A(n7374), .Z(n7372) );
  ANDN U15409 ( .B(n7375), .A(n7376), .Z(n7316) );
  XOR U15410 ( .A(n7302), .B(n7377), .Z(n7314) );
  XOR U15411 ( .A(n7303), .B(n7304), .Z(n7377) );
  XOR U15412 ( .A(n7309), .B(n7378), .Z(n7304) );
  XOR U15413 ( .A(n7308), .B(n7311), .Z(n7378) );
  IV U15414 ( .A(n7310), .Z(n7311) );
  NAND U15415 ( .A(n7379), .B(n7380), .Z(n7310) );
  OR U15416 ( .A(n7381), .B(n7382), .Z(n7380) );
  OR U15417 ( .A(n7383), .B(n7384), .Z(n7379) );
  NAND U15418 ( .A(n7385), .B(n7386), .Z(n7308) );
  OR U15419 ( .A(n7387), .B(n7388), .Z(n7386) );
  OR U15420 ( .A(n7389), .B(n7390), .Z(n7385) );
  NOR U15421 ( .A(n7391), .B(n7392), .Z(n7309) );
  ANDN U15422 ( .B(n7393), .A(n7394), .Z(n7303) );
  IV U15423 ( .A(n7395), .Z(n7393) );
  XNOR U15424 ( .A(n7296), .B(n7396), .Z(n7302) );
  XNOR U15425 ( .A(n7295), .B(n7297), .Z(n7396) );
  NAND U15426 ( .A(n7397), .B(n7398), .Z(n7297) );
  OR U15427 ( .A(n7399), .B(n7400), .Z(n7398) );
  OR U15428 ( .A(n7401), .B(n7402), .Z(n7397) );
  NAND U15429 ( .A(n7403), .B(n7404), .Z(n7295) );
  OR U15430 ( .A(n7405), .B(n7406), .Z(n7404) );
  OR U15431 ( .A(n7407), .B(n7408), .Z(n7403) );
  ANDN U15432 ( .B(n7409), .A(n7410), .Z(n7296) );
  IV U15433 ( .A(n7411), .Z(n7409) );
  XNOR U15434 ( .A(n7376), .B(n7375), .Z(N64739) );
  XOR U15435 ( .A(n7395), .B(n7394), .Z(n7375) );
  XNOR U15436 ( .A(n7410), .B(n7411), .Z(n7394) );
  XNOR U15437 ( .A(n7405), .B(n7406), .Z(n7411) );
  XNOR U15438 ( .A(n7407), .B(n7408), .Z(n7406) );
  XNOR U15439 ( .A(y[7669]), .B(x[7669]), .Z(n7408) );
  XNOR U15440 ( .A(y[7670]), .B(x[7670]), .Z(n7407) );
  XNOR U15441 ( .A(y[7668]), .B(x[7668]), .Z(n7405) );
  XNOR U15442 ( .A(n7399), .B(n7400), .Z(n7410) );
  XNOR U15443 ( .A(y[7665]), .B(x[7665]), .Z(n7400) );
  XNOR U15444 ( .A(n7401), .B(n7402), .Z(n7399) );
  XNOR U15445 ( .A(y[7666]), .B(x[7666]), .Z(n7402) );
  XNOR U15446 ( .A(y[7667]), .B(x[7667]), .Z(n7401) );
  XNOR U15447 ( .A(n7392), .B(n7391), .Z(n7395) );
  XNOR U15448 ( .A(n7387), .B(n7388), .Z(n7391) );
  XNOR U15449 ( .A(y[7662]), .B(x[7662]), .Z(n7388) );
  XNOR U15450 ( .A(n7389), .B(n7390), .Z(n7387) );
  XNOR U15451 ( .A(y[7663]), .B(x[7663]), .Z(n7390) );
  XNOR U15452 ( .A(y[7664]), .B(x[7664]), .Z(n7389) );
  XNOR U15453 ( .A(n7381), .B(n7382), .Z(n7392) );
  XNOR U15454 ( .A(y[7659]), .B(x[7659]), .Z(n7382) );
  XNOR U15455 ( .A(n7383), .B(n7384), .Z(n7381) );
  XNOR U15456 ( .A(y[7660]), .B(x[7660]), .Z(n7384) );
  XNOR U15457 ( .A(y[7661]), .B(x[7661]), .Z(n7383) );
  XOR U15458 ( .A(n7357), .B(n7358), .Z(n7376) );
  XNOR U15459 ( .A(n7373), .B(n7374), .Z(n7358) );
  XNOR U15460 ( .A(n7368), .B(n7369), .Z(n7374) );
  XNOR U15461 ( .A(n7370), .B(n7371), .Z(n7369) );
  XNOR U15462 ( .A(y[7657]), .B(x[7657]), .Z(n7371) );
  XNOR U15463 ( .A(y[7658]), .B(x[7658]), .Z(n7370) );
  XNOR U15464 ( .A(y[7656]), .B(x[7656]), .Z(n7368) );
  XNOR U15465 ( .A(n7362), .B(n7363), .Z(n7373) );
  XNOR U15466 ( .A(y[7653]), .B(x[7653]), .Z(n7363) );
  XNOR U15467 ( .A(n7364), .B(n7365), .Z(n7362) );
  XNOR U15468 ( .A(y[7654]), .B(x[7654]), .Z(n7365) );
  XNOR U15469 ( .A(y[7655]), .B(x[7655]), .Z(n7364) );
  XOR U15470 ( .A(n7356), .B(n7355), .Z(n7357) );
  XNOR U15471 ( .A(n7351), .B(n7352), .Z(n7355) );
  XNOR U15472 ( .A(y[7650]), .B(x[7650]), .Z(n7352) );
  XNOR U15473 ( .A(n7353), .B(n7354), .Z(n7351) );
  XNOR U15474 ( .A(y[7651]), .B(x[7651]), .Z(n7354) );
  XNOR U15475 ( .A(y[7652]), .B(x[7652]), .Z(n7353) );
  XNOR U15476 ( .A(n7345), .B(n7346), .Z(n7356) );
  XNOR U15477 ( .A(y[7647]), .B(x[7647]), .Z(n7346) );
  XNOR U15478 ( .A(n7347), .B(n7348), .Z(n7345) );
  XNOR U15479 ( .A(y[7648]), .B(x[7648]), .Z(n7348) );
  XNOR U15480 ( .A(y[7649]), .B(x[7649]), .Z(n7347) );
  NAND U15481 ( .A(n7412), .B(n7413), .Z(N64730) );
  NANDN U15482 ( .A(n7414), .B(n7415), .Z(n7413) );
  OR U15483 ( .A(n7416), .B(n7417), .Z(n7415) );
  NAND U15484 ( .A(n7416), .B(n7417), .Z(n7412) );
  XOR U15485 ( .A(n7416), .B(n7418), .Z(N64729) );
  XNOR U15486 ( .A(n7414), .B(n7417), .Z(n7418) );
  AND U15487 ( .A(n7419), .B(n7420), .Z(n7417) );
  NANDN U15488 ( .A(n7421), .B(n7422), .Z(n7420) );
  NANDN U15489 ( .A(n7423), .B(n7424), .Z(n7422) );
  NANDN U15490 ( .A(n7424), .B(n7423), .Z(n7419) );
  NAND U15491 ( .A(n7425), .B(n7426), .Z(n7414) );
  NANDN U15492 ( .A(n7427), .B(n7428), .Z(n7426) );
  OR U15493 ( .A(n7429), .B(n7430), .Z(n7428) );
  NAND U15494 ( .A(n7430), .B(n7429), .Z(n7425) );
  AND U15495 ( .A(n7431), .B(n7432), .Z(n7416) );
  NANDN U15496 ( .A(n7433), .B(n7434), .Z(n7432) );
  NANDN U15497 ( .A(n7435), .B(n7436), .Z(n7434) );
  NANDN U15498 ( .A(n7436), .B(n7435), .Z(n7431) );
  XOR U15499 ( .A(n7430), .B(n7437), .Z(N64728) );
  XOR U15500 ( .A(n7427), .B(n7429), .Z(n7437) );
  XNOR U15501 ( .A(n7423), .B(n7438), .Z(n7429) );
  XNOR U15502 ( .A(n7421), .B(n7424), .Z(n7438) );
  NAND U15503 ( .A(n7439), .B(n7440), .Z(n7424) );
  NAND U15504 ( .A(n7441), .B(n7442), .Z(n7440) );
  OR U15505 ( .A(n7443), .B(n7444), .Z(n7441) );
  NANDN U15506 ( .A(n7445), .B(n7443), .Z(n7439) );
  IV U15507 ( .A(n7444), .Z(n7445) );
  NAND U15508 ( .A(n7446), .B(n7447), .Z(n7421) );
  NAND U15509 ( .A(n7448), .B(n7449), .Z(n7447) );
  NANDN U15510 ( .A(n7450), .B(n7451), .Z(n7448) );
  NANDN U15511 ( .A(n7451), .B(n7450), .Z(n7446) );
  AND U15512 ( .A(n7452), .B(n7453), .Z(n7423) );
  NAND U15513 ( .A(n7454), .B(n7455), .Z(n7453) );
  OR U15514 ( .A(n7456), .B(n7457), .Z(n7454) );
  NANDN U15515 ( .A(n7458), .B(n7456), .Z(n7452) );
  NAND U15516 ( .A(n7459), .B(n7460), .Z(n7427) );
  NANDN U15517 ( .A(n7461), .B(n7462), .Z(n7460) );
  OR U15518 ( .A(n7463), .B(n7464), .Z(n7462) );
  NANDN U15519 ( .A(n7465), .B(n7463), .Z(n7459) );
  IV U15520 ( .A(n7464), .Z(n7465) );
  XNOR U15521 ( .A(n7435), .B(n7466), .Z(n7430) );
  XNOR U15522 ( .A(n7433), .B(n7436), .Z(n7466) );
  NAND U15523 ( .A(n7467), .B(n7468), .Z(n7436) );
  NAND U15524 ( .A(n7469), .B(n7470), .Z(n7468) );
  OR U15525 ( .A(n7471), .B(n7472), .Z(n7469) );
  NANDN U15526 ( .A(n7473), .B(n7471), .Z(n7467) );
  IV U15527 ( .A(n7472), .Z(n7473) );
  NAND U15528 ( .A(n7474), .B(n7475), .Z(n7433) );
  NAND U15529 ( .A(n7476), .B(n7477), .Z(n7475) );
  NANDN U15530 ( .A(n7478), .B(n7479), .Z(n7476) );
  NANDN U15531 ( .A(n7479), .B(n7478), .Z(n7474) );
  AND U15532 ( .A(n7480), .B(n7481), .Z(n7435) );
  NAND U15533 ( .A(n7482), .B(n7483), .Z(n7481) );
  OR U15534 ( .A(n7484), .B(n7485), .Z(n7482) );
  NANDN U15535 ( .A(n7486), .B(n7484), .Z(n7480) );
  XNOR U15536 ( .A(n7461), .B(n7487), .Z(N64727) );
  XOR U15537 ( .A(n7463), .B(n7464), .Z(n7487) );
  XNOR U15538 ( .A(n7477), .B(n7488), .Z(n7464) );
  XOR U15539 ( .A(n7478), .B(n7479), .Z(n7488) );
  XOR U15540 ( .A(n7484), .B(n7489), .Z(n7479) );
  XOR U15541 ( .A(n7483), .B(n7486), .Z(n7489) );
  IV U15542 ( .A(n7485), .Z(n7486) );
  NAND U15543 ( .A(n7490), .B(n7491), .Z(n7485) );
  OR U15544 ( .A(n7492), .B(n7493), .Z(n7491) );
  OR U15545 ( .A(n7494), .B(n7495), .Z(n7490) );
  NAND U15546 ( .A(n7496), .B(n7497), .Z(n7483) );
  OR U15547 ( .A(n7498), .B(n7499), .Z(n7497) );
  OR U15548 ( .A(n7500), .B(n7501), .Z(n7496) );
  NOR U15549 ( .A(n7502), .B(n7503), .Z(n7484) );
  ANDN U15550 ( .B(n7504), .A(n7505), .Z(n7478) );
  XNOR U15551 ( .A(n7471), .B(n7506), .Z(n7477) );
  XNOR U15552 ( .A(n7470), .B(n7472), .Z(n7506) );
  NAND U15553 ( .A(n7507), .B(n7508), .Z(n7472) );
  OR U15554 ( .A(n7509), .B(n7510), .Z(n7508) );
  OR U15555 ( .A(n7511), .B(n7512), .Z(n7507) );
  NAND U15556 ( .A(n7513), .B(n7514), .Z(n7470) );
  OR U15557 ( .A(n7515), .B(n7516), .Z(n7514) );
  OR U15558 ( .A(n7517), .B(n7518), .Z(n7513) );
  ANDN U15559 ( .B(n7519), .A(n7520), .Z(n7471) );
  IV U15560 ( .A(n7521), .Z(n7519) );
  ANDN U15561 ( .B(n7522), .A(n7523), .Z(n7463) );
  XOR U15562 ( .A(n7449), .B(n7524), .Z(n7461) );
  XOR U15563 ( .A(n7450), .B(n7451), .Z(n7524) );
  XOR U15564 ( .A(n7456), .B(n7525), .Z(n7451) );
  XOR U15565 ( .A(n7455), .B(n7458), .Z(n7525) );
  IV U15566 ( .A(n7457), .Z(n7458) );
  NAND U15567 ( .A(n7526), .B(n7527), .Z(n7457) );
  OR U15568 ( .A(n7528), .B(n7529), .Z(n7527) );
  OR U15569 ( .A(n7530), .B(n7531), .Z(n7526) );
  NAND U15570 ( .A(n7532), .B(n7533), .Z(n7455) );
  OR U15571 ( .A(n7534), .B(n7535), .Z(n7533) );
  OR U15572 ( .A(n7536), .B(n7537), .Z(n7532) );
  NOR U15573 ( .A(n7538), .B(n7539), .Z(n7456) );
  ANDN U15574 ( .B(n7540), .A(n7541), .Z(n7450) );
  IV U15575 ( .A(n7542), .Z(n7540) );
  XNOR U15576 ( .A(n7443), .B(n7543), .Z(n7449) );
  XNOR U15577 ( .A(n7442), .B(n7444), .Z(n7543) );
  NAND U15578 ( .A(n7544), .B(n7545), .Z(n7444) );
  OR U15579 ( .A(n7546), .B(n7547), .Z(n7545) );
  OR U15580 ( .A(n7548), .B(n7549), .Z(n7544) );
  NAND U15581 ( .A(n7550), .B(n7551), .Z(n7442) );
  OR U15582 ( .A(n7552), .B(n7553), .Z(n7551) );
  OR U15583 ( .A(n7554), .B(n7555), .Z(n7550) );
  ANDN U15584 ( .B(n7556), .A(n7557), .Z(n7443) );
  IV U15585 ( .A(n7558), .Z(n7556) );
  XNOR U15586 ( .A(n7523), .B(n7522), .Z(N64726) );
  XOR U15587 ( .A(n7542), .B(n7541), .Z(n7522) );
  XNOR U15588 ( .A(n7557), .B(n7558), .Z(n7541) );
  XNOR U15589 ( .A(n7552), .B(n7553), .Z(n7558) );
  XNOR U15590 ( .A(n7554), .B(n7555), .Z(n7553) );
  XNOR U15591 ( .A(y[7645]), .B(x[7645]), .Z(n7555) );
  XNOR U15592 ( .A(y[7646]), .B(x[7646]), .Z(n7554) );
  XNOR U15593 ( .A(y[7644]), .B(x[7644]), .Z(n7552) );
  XNOR U15594 ( .A(n7546), .B(n7547), .Z(n7557) );
  XNOR U15595 ( .A(y[7641]), .B(x[7641]), .Z(n7547) );
  XNOR U15596 ( .A(n7548), .B(n7549), .Z(n7546) );
  XNOR U15597 ( .A(y[7642]), .B(x[7642]), .Z(n7549) );
  XNOR U15598 ( .A(y[7643]), .B(x[7643]), .Z(n7548) );
  XNOR U15599 ( .A(n7539), .B(n7538), .Z(n7542) );
  XNOR U15600 ( .A(n7534), .B(n7535), .Z(n7538) );
  XNOR U15601 ( .A(y[7638]), .B(x[7638]), .Z(n7535) );
  XNOR U15602 ( .A(n7536), .B(n7537), .Z(n7534) );
  XNOR U15603 ( .A(y[7639]), .B(x[7639]), .Z(n7537) );
  XNOR U15604 ( .A(y[7640]), .B(x[7640]), .Z(n7536) );
  XNOR U15605 ( .A(n7528), .B(n7529), .Z(n7539) );
  XNOR U15606 ( .A(y[7635]), .B(x[7635]), .Z(n7529) );
  XNOR U15607 ( .A(n7530), .B(n7531), .Z(n7528) );
  XNOR U15608 ( .A(y[7636]), .B(x[7636]), .Z(n7531) );
  XNOR U15609 ( .A(y[7637]), .B(x[7637]), .Z(n7530) );
  XOR U15610 ( .A(n7504), .B(n7505), .Z(n7523) );
  XNOR U15611 ( .A(n7520), .B(n7521), .Z(n7505) );
  XNOR U15612 ( .A(n7515), .B(n7516), .Z(n7521) );
  XNOR U15613 ( .A(n7517), .B(n7518), .Z(n7516) );
  XNOR U15614 ( .A(y[7633]), .B(x[7633]), .Z(n7518) );
  XNOR U15615 ( .A(y[7634]), .B(x[7634]), .Z(n7517) );
  XNOR U15616 ( .A(y[7632]), .B(x[7632]), .Z(n7515) );
  XNOR U15617 ( .A(n7509), .B(n7510), .Z(n7520) );
  XNOR U15618 ( .A(y[7629]), .B(x[7629]), .Z(n7510) );
  XNOR U15619 ( .A(n7511), .B(n7512), .Z(n7509) );
  XNOR U15620 ( .A(y[7630]), .B(x[7630]), .Z(n7512) );
  XNOR U15621 ( .A(y[7631]), .B(x[7631]), .Z(n7511) );
  XOR U15622 ( .A(n7503), .B(n7502), .Z(n7504) );
  XNOR U15623 ( .A(n7498), .B(n7499), .Z(n7502) );
  XNOR U15624 ( .A(y[7626]), .B(x[7626]), .Z(n7499) );
  XNOR U15625 ( .A(n7500), .B(n7501), .Z(n7498) );
  XNOR U15626 ( .A(y[7627]), .B(x[7627]), .Z(n7501) );
  XNOR U15627 ( .A(y[7628]), .B(x[7628]), .Z(n7500) );
  XNOR U15628 ( .A(n7492), .B(n7493), .Z(n7503) );
  XNOR U15629 ( .A(y[7623]), .B(x[7623]), .Z(n7493) );
  XNOR U15630 ( .A(n7494), .B(n7495), .Z(n7492) );
  XNOR U15631 ( .A(y[7624]), .B(x[7624]), .Z(n7495) );
  XNOR U15632 ( .A(y[7625]), .B(x[7625]), .Z(n7494) );
  NAND U15633 ( .A(n7559), .B(n7560), .Z(N64717) );
  NANDN U15634 ( .A(n7561), .B(n7562), .Z(n7560) );
  OR U15635 ( .A(n7563), .B(n7564), .Z(n7562) );
  NAND U15636 ( .A(n7563), .B(n7564), .Z(n7559) );
  XOR U15637 ( .A(n7563), .B(n7565), .Z(N64716) );
  XNOR U15638 ( .A(n7561), .B(n7564), .Z(n7565) );
  AND U15639 ( .A(n7566), .B(n7567), .Z(n7564) );
  NANDN U15640 ( .A(n7568), .B(n7569), .Z(n7567) );
  NANDN U15641 ( .A(n7570), .B(n7571), .Z(n7569) );
  NANDN U15642 ( .A(n7571), .B(n7570), .Z(n7566) );
  NAND U15643 ( .A(n7572), .B(n7573), .Z(n7561) );
  NANDN U15644 ( .A(n7574), .B(n7575), .Z(n7573) );
  OR U15645 ( .A(n7576), .B(n7577), .Z(n7575) );
  NAND U15646 ( .A(n7577), .B(n7576), .Z(n7572) );
  AND U15647 ( .A(n7578), .B(n7579), .Z(n7563) );
  NANDN U15648 ( .A(n7580), .B(n7581), .Z(n7579) );
  NANDN U15649 ( .A(n7582), .B(n7583), .Z(n7581) );
  NANDN U15650 ( .A(n7583), .B(n7582), .Z(n7578) );
  XOR U15651 ( .A(n7577), .B(n7584), .Z(N64715) );
  XOR U15652 ( .A(n7574), .B(n7576), .Z(n7584) );
  XNOR U15653 ( .A(n7570), .B(n7585), .Z(n7576) );
  XNOR U15654 ( .A(n7568), .B(n7571), .Z(n7585) );
  NAND U15655 ( .A(n7586), .B(n7587), .Z(n7571) );
  NAND U15656 ( .A(n7588), .B(n7589), .Z(n7587) );
  OR U15657 ( .A(n7590), .B(n7591), .Z(n7588) );
  NANDN U15658 ( .A(n7592), .B(n7590), .Z(n7586) );
  IV U15659 ( .A(n7591), .Z(n7592) );
  NAND U15660 ( .A(n7593), .B(n7594), .Z(n7568) );
  NAND U15661 ( .A(n7595), .B(n7596), .Z(n7594) );
  NANDN U15662 ( .A(n7597), .B(n7598), .Z(n7595) );
  NANDN U15663 ( .A(n7598), .B(n7597), .Z(n7593) );
  AND U15664 ( .A(n7599), .B(n7600), .Z(n7570) );
  NAND U15665 ( .A(n7601), .B(n7602), .Z(n7600) );
  OR U15666 ( .A(n7603), .B(n7604), .Z(n7601) );
  NANDN U15667 ( .A(n7605), .B(n7603), .Z(n7599) );
  NAND U15668 ( .A(n7606), .B(n7607), .Z(n7574) );
  NANDN U15669 ( .A(n7608), .B(n7609), .Z(n7607) );
  OR U15670 ( .A(n7610), .B(n7611), .Z(n7609) );
  NANDN U15671 ( .A(n7612), .B(n7610), .Z(n7606) );
  IV U15672 ( .A(n7611), .Z(n7612) );
  XNOR U15673 ( .A(n7582), .B(n7613), .Z(n7577) );
  XNOR U15674 ( .A(n7580), .B(n7583), .Z(n7613) );
  NAND U15675 ( .A(n7614), .B(n7615), .Z(n7583) );
  NAND U15676 ( .A(n7616), .B(n7617), .Z(n7615) );
  OR U15677 ( .A(n7618), .B(n7619), .Z(n7616) );
  NANDN U15678 ( .A(n7620), .B(n7618), .Z(n7614) );
  IV U15679 ( .A(n7619), .Z(n7620) );
  NAND U15680 ( .A(n7621), .B(n7622), .Z(n7580) );
  NAND U15681 ( .A(n7623), .B(n7624), .Z(n7622) );
  NANDN U15682 ( .A(n7625), .B(n7626), .Z(n7623) );
  NANDN U15683 ( .A(n7626), .B(n7625), .Z(n7621) );
  AND U15684 ( .A(n7627), .B(n7628), .Z(n7582) );
  NAND U15685 ( .A(n7629), .B(n7630), .Z(n7628) );
  OR U15686 ( .A(n7631), .B(n7632), .Z(n7629) );
  NANDN U15687 ( .A(n7633), .B(n7631), .Z(n7627) );
  XNOR U15688 ( .A(n7608), .B(n7634), .Z(N64714) );
  XOR U15689 ( .A(n7610), .B(n7611), .Z(n7634) );
  XNOR U15690 ( .A(n7624), .B(n7635), .Z(n7611) );
  XOR U15691 ( .A(n7625), .B(n7626), .Z(n7635) );
  XOR U15692 ( .A(n7631), .B(n7636), .Z(n7626) );
  XOR U15693 ( .A(n7630), .B(n7633), .Z(n7636) );
  IV U15694 ( .A(n7632), .Z(n7633) );
  NAND U15695 ( .A(n7637), .B(n7638), .Z(n7632) );
  OR U15696 ( .A(n7639), .B(n7640), .Z(n7638) );
  OR U15697 ( .A(n7641), .B(n7642), .Z(n7637) );
  NAND U15698 ( .A(n7643), .B(n7644), .Z(n7630) );
  OR U15699 ( .A(n7645), .B(n7646), .Z(n7644) );
  OR U15700 ( .A(n7647), .B(n7648), .Z(n7643) );
  NOR U15701 ( .A(n7649), .B(n7650), .Z(n7631) );
  ANDN U15702 ( .B(n7651), .A(n7652), .Z(n7625) );
  XNOR U15703 ( .A(n7618), .B(n7653), .Z(n7624) );
  XNOR U15704 ( .A(n7617), .B(n7619), .Z(n7653) );
  NAND U15705 ( .A(n7654), .B(n7655), .Z(n7619) );
  OR U15706 ( .A(n7656), .B(n7657), .Z(n7655) );
  OR U15707 ( .A(n7658), .B(n7659), .Z(n7654) );
  NAND U15708 ( .A(n7660), .B(n7661), .Z(n7617) );
  OR U15709 ( .A(n7662), .B(n7663), .Z(n7661) );
  OR U15710 ( .A(n7664), .B(n7665), .Z(n7660) );
  ANDN U15711 ( .B(n7666), .A(n7667), .Z(n7618) );
  IV U15712 ( .A(n7668), .Z(n7666) );
  ANDN U15713 ( .B(n7669), .A(n7670), .Z(n7610) );
  XOR U15714 ( .A(n7596), .B(n7671), .Z(n7608) );
  XOR U15715 ( .A(n7597), .B(n7598), .Z(n7671) );
  XOR U15716 ( .A(n7603), .B(n7672), .Z(n7598) );
  XOR U15717 ( .A(n7602), .B(n7605), .Z(n7672) );
  IV U15718 ( .A(n7604), .Z(n7605) );
  NAND U15719 ( .A(n7673), .B(n7674), .Z(n7604) );
  OR U15720 ( .A(n7675), .B(n7676), .Z(n7674) );
  OR U15721 ( .A(n7677), .B(n7678), .Z(n7673) );
  NAND U15722 ( .A(n7679), .B(n7680), .Z(n7602) );
  OR U15723 ( .A(n7681), .B(n7682), .Z(n7680) );
  OR U15724 ( .A(n7683), .B(n7684), .Z(n7679) );
  NOR U15725 ( .A(n7685), .B(n7686), .Z(n7603) );
  ANDN U15726 ( .B(n7687), .A(n7688), .Z(n7597) );
  IV U15727 ( .A(n7689), .Z(n7687) );
  XNOR U15728 ( .A(n7590), .B(n7690), .Z(n7596) );
  XNOR U15729 ( .A(n7589), .B(n7591), .Z(n7690) );
  NAND U15730 ( .A(n7691), .B(n7692), .Z(n7591) );
  OR U15731 ( .A(n7693), .B(n7694), .Z(n7692) );
  OR U15732 ( .A(n7695), .B(n7696), .Z(n7691) );
  NAND U15733 ( .A(n7697), .B(n7698), .Z(n7589) );
  OR U15734 ( .A(n7699), .B(n7700), .Z(n7698) );
  OR U15735 ( .A(n7701), .B(n7702), .Z(n7697) );
  ANDN U15736 ( .B(n7703), .A(n7704), .Z(n7590) );
  IV U15737 ( .A(n7705), .Z(n7703) );
  XNOR U15738 ( .A(n7670), .B(n7669), .Z(N64713) );
  XOR U15739 ( .A(n7689), .B(n7688), .Z(n7669) );
  XNOR U15740 ( .A(n7704), .B(n7705), .Z(n7688) );
  XNOR U15741 ( .A(n7699), .B(n7700), .Z(n7705) );
  XNOR U15742 ( .A(n7701), .B(n7702), .Z(n7700) );
  XNOR U15743 ( .A(y[7621]), .B(x[7621]), .Z(n7702) );
  XNOR U15744 ( .A(y[7622]), .B(x[7622]), .Z(n7701) );
  XNOR U15745 ( .A(y[7620]), .B(x[7620]), .Z(n7699) );
  XNOR U15746 ( .A(n7693), .B(n7694), .Z(n7704) );
  XNOR U15747 ( .A(y[7617]), .B(x[7617]), .Z(n7694) );
  XNOR U15748 ( .A(n7695), .B(n7696), .Z(n7693) );
  XNOR U15749 ( .A(y[7618]), .B(x[7618]), .Z(n7696) );
  XNOR U15750 ( .A(y[7619]), .B(x[7619]), .Z(n7695) );
  XNOR U15751 ( .A(n7686), .B(n7685), .Z(n7689) );
  XNOR U15752 ( .A(n7681), .B(n7682), .Z(n7685) );
  XNOR U15753 ( .A(y[7614]), .B(x[7614]), .Z(n7682) );
  XNOR U15754 ( .A(n7683), .B(n7684), .Z(n7681) );
  XNOR U15755 ( .A(y[7615]), .B(x[7615]), .Z(n7684) );
  XNOR U15756 ( .A(y[7616]), .B(x[7616]), .Z(n7683) );
  XNOR U15757 ( .A(n7675), .B(n7676), .Z(n7686) );
  XNOR U15758 ( .A(y[7611]), .B(x[7611]), .Z(n7676) );
  XNOR U15759 ( .A(n7677), .B(n7678), .Z(n7675) );
  XNOR U15760 ( .A(y[7612]), .B(x[7612]), .Z(n7678) );
  XNOR U15761 ( .A(y[7613]), .B(x[7613]), .Z(n7677) );
  XOR U15762 ( .A(n7651), .B(n7652), .Z(n7670) );
  XNOR U15763 ( .A(n7667), .B(n7668), .Z(n7652) );
  XNOR U15764 ( .A(n7662), .B(n7663), .Z(n7668) );
  XNOR U15765 ( .A(n7664), .B(n7665), .Z(n7663) );
  XNOR U15766 ( .A(y[7609]), .B(x[7609]), .Z(n7665) );
  XNOR U15767 ( .A(y[7610]), .B(x[7610]), .Z(n7664) );
  XNOR U15768 ( .A(y[7608]), .B(x[7608]), .Z(n7662) );
  XNOR U15769 ( .A(n7656), .B(n7657), .Z(n7667) );
  XNOR U15770 ( .A(y[7605]), .B(x[7605]), .Z(n7657) );
  XNOR U15771 ( .A(n7658), .B(n7659), .Z(n7656) );
  XNOR U15772 ( .A(y[7606]), .B(x[7606]), .Z(n7659) );
  XNOR U15773 ( .A(y[7607]), .B(x[7607]), .Z(n7658) );
  XOR U15774 ( .A(n7650), .B(n7649), .Z(n7651) );
  XNOR U15775 ( .A(n7645), .B(n7646), .Z(n7649) );
  XNOR U15776 ( .A(y[7602]), .B(x[7602]), .Z(n7646) );
  XNOR U15777 ( .A(n7647), .B(n7648), .Z(n7645) );
  XNOR U15778 ( .A(y[7603]), .B(x[7603]), .Z(n7648) );
  XNOR U15779 ( .A(y[7604]), .B(x[7604]), .Z(n7647) );
  XNOR U15780 ( .A(n7639), .B(n7640), .Z(n7650) );
  XNOR U15781 ( .A(y[7599]), .B(x[7599]), .Z(n7640) );
  XNOR U15782 ( .A(n7641), .B(n7642), .Z(n7639) );
  XNOR U15783 ( .A(y[7600]), .B(x[7600]), .Z(n7642) );
  XNOR U15784 ( .A(y[7601]), .B(x[7601]), .Z(n7641) );
  NAND U15785 ( .A(n7706), .B(n7707), .Z(N64704) );
  NANDN U15786 ( .A(n7708), .B(n7709), .Z(n7707) );
  OR U15787 ( .A(n7710), .B(n7711), .Z(n7709) );
  NAND U15788 ( .A(n7710), .B(n7711), .Z(n7706) );
  XOR U15789 ( .A(n7710), .B(n7712), .Z(N64703) );
  XNOR U15790 ( .A(n7708), .B(n7711), .Z(n7712) );
  AND U15791 ( .A(n7713), .B(n7714), .Z(n7711) );
  NANDN U15792 ( .A(n7715), .B(n7716), .Z(n7714) );
  NANDN U15793 ( .A(n7717), .B(n7718), .Z(n7716) );
  NANDN U15794 ( .A(n7718), .B(n7717), .Z(n7713) );
  NAND U15795 ( .A(n7719), .B(n7720), .Z(n7708) );
  NANDN U15796 ( .A(n7721), .B(n7722), .Z(n7720) );
  OR U15797 ( .A(n7723), .B(n7724), .Z(n7722) );
  NAND U15798 ( .A(n7724), .B(n7723), .Z(n7719) );
  AND U15799 ( .A(n7725), .B(n7726), .Z(n7710) );
  NANDN U15800 ( .A(n7727), .B(n7728), .Z(n7726) );
  NANDN U15801 ( .A(n7729), .B(n7730), .Z(n7728) );
  NANDN U15802 ( .A(n7730), .B(n7729), .Z(n7725) );
  XOR U15803 ( .A(n7724), .B(n7731), .Z(N64702) );
  XOR U15804 ( .A(n7721), .B(n7723), .Z(n7731) );
  XNOR U15805 ( .A(n7717), .B(n7732), .Z(n7723) );
  XNOR U15806 ( .A(n7715), .B(n7718), .Z(n7732) );
  NAND U15807 ( .A(n7733), .B(n7734), .Z(n7718) );
  NAND U15808 ( .A(n7735), .B(n7736), .Z(n7734) );
  OR U15809 ( .A(n7737), .B(n7738), .Z(n7735) );
  NANDN U15810 ( .A(n7739), .B(n7737), .Z(n7733) );
  IV U15811 ( .A(n7738), .Z(n7739) );
  NAND U15812 ( .A(n7740), .B(n7741), .Z(n7715) );
  NAND U15813 ( .A(n7742), .B(n7743), .Z(n7741) );
  NANDN U15814 ( .A(n7744), .B(n7745), .Z(n7742) );
  NANDN U15815 ( .A(n7745), .B(n7744), .Z(n7740) );
  AND U15816 ( .A(n7746), .B(n7747), .Z(n7717) );
  NAND U15817 ( .A(n7748), .B(n7749), .Z(n7747) );
  OR U15818 ( .A(n7750), .B(n7751), .Z(n7748) );
  NANDN U15819 ( .A(n7752), .B(n7750), .Z(n7746) );
  NAND U15820 ( .A(n7753), .B(n7754), .Z(n7721) );
  NANDN U15821 ( .A(n7755), .B(n7756), .Z(n7754) );
  OR U15822 ( .A(n7757), .B(n7758), .Z(n7756) );
  NANDN U15823 ( .A(n7759), .B(n7757), .Z(n7753) );
  IV U15824 ( .A(n7758), .Z(n7759) );
  XNOR U15825 ( .A(n7729), .B(n7760), .Z(n7724) );
  XNOR U15826 ( .A(n7727), .B(n7730), .Z(n7760) );
  NAND U15827 ( .A(n7761), .B(n7762), .Z(n7730) );
  NAND U15828 ( .A(n7763), .B(n7764), .Z(n7762) );
  OR U15829 ( .A(n7765), .B(n7766), .Z(n7763) );
  NANDN U15830 ( .A(n7767), .B(n7765), .Z(n7761) );
  IV U15831 ( .A(n7766), .Z(n7767) );
  NAND U15832 ( .A(n7768), .B(n7769), .Z(n7727) );
  NAND U15833 ( .A(n7770), .B(n7771), .Z(n7769) );
  NANDN U15834 ( .A(n7772), .B(n7773), .Z(n7770) );
  NANDN U15835 ( .A(n7773), .B(n7772), .Z(n7768) );
  AND U15836 ( .A(n7774), .B(n7775), .Z(n7729) );
  NAND U15837 ( .A(n7776), .B(n7777), .Z(n7775) );
  OR U15838 ( .A(n7778), .B(n7779), .Z(n7776) );
  NANDN U15839 ( .A(n7780), .B(n7778), .Z(n7774) );
  XNOR U15840 ( .A(n7755), .B(n7781), .Z(N64701) );
  XOR U15841 ( .A(n7757), .B(n7758), .Z(n7781) );
  XNOR U15842 ( .A(n7771), .B(n7782), .Z(n7758) );
  XOR U15843 ( .A(n7772), .B(n7773), .Z(n7782) );
  XOR U15844 ( .A(n7778), .B(n7783), .Z(n7773) );
  XOR U15845 ( .A(n7777), .B(n7780), .Z(n7783) );
  IV U15846 ( .A(n7779), .Z(n7780) );
  NAND U15847 ( .A(n7784), .B(n7785), .Z(n7779) );
  OR U15848 ( .A(n7786), .B(n7787), .Z(n7785) );
  OR U15849 ( .A(n7788), .B(n7789), .Z(n7784) );
  NAND U15850 ( .A(n7790), .B(n7791), .Z(n7777) );
  OR U15851 ( .A(n7792), .B(n7793), .Z(n7791) );
  OR U15852 ( .A(n7794), .B(n7795), .Z(n7790) );
  NOR U15853 ( .A(n7796), .B(n7797), .Z(n7778) );
  ANDN U15854 ( .B(n7798), .A(n7799), .Z(n7772) );
  XNOR U15855 ( .A(n7765), .B(n7800), .Z(n7771) );
  XNOR U15856 ( .A(n7764), .B(n7766), .Z(n7800) );
  NAND U15857 ( .A(n7801), .B(n7802), .Z(n7766) );
  OR U15858 ( .A(n7803), .B(n7804), .Z(n7802) );
  OR U15859 ( .A(n7805), .B(n7806), .Z(n7801) );
  NAND U15860 ( .A(n7807), .B(n7808), .Z(n7764) );
  OR U15861 ( .A(n7809), .B(n7810), .Z(n7808) );
  OR U15862 ( .A(n7811), .B(n7812), .Z(n7807) );
  ANDN U15863 ( .B(n7813), .A(n7814), .Z(n7765) );
  IV U15864 ( .A(n7815), .Z(n7813) );
  ANDN U15865 ( .B(n7816), .A(n7817), .Z(n7757) );
  XOR U15866 ( .A(n7743), .B(n7818), .Z(n7755) );
  XOR U15867 ( .A(n7744), .B(n7745), .Z(n7818) );
  XOR U15868 ( .A(n7750), .B(n7819), .Z(n7745) );
  XOR U15869 ( .A(n7749), .B(n7752), .Z(n7819) );
  IV U15870 ( .A(n7751), .Z(n7752) );
  NAND U15871 ( .A(n7820), .B(n7821), .Z(n7751) );
  OR U15872 ( .A(n7822), .B(n7823), .Z(n7821) );
  OR U15873 ( .A(n7824), .B(n7825), .Z(n7820) );
  NAND U15874 ( .A(n7826), .B(n7827), .Z(n7749) );
  OR U15875 ( .A(n7828), .B(n7829), .Z(n7827) );
  OR U15876 ( .A(n7830), .B(n7831), .Z(n7826) );
  NOR U15877 ( .A(n7832), .B(n7833), .Z(n7750) );
  ANDN U15878 ( .B(n7834), .A(n7835), .Z(n7744) );
  IV U15879 ( .A(n7836), .Z(n7834) );
  XNOR U15880 ( .A(n7737), .B(n7837), .Z(n7743) );
  XNOR U15881 ( .A(n7736), .B(n7738), .Z(n7837) );
  NAND U15882 ( .A(n7838), .B(n7839), .Z(n7738) );
  OR U15883 ( .A(n7840), .B(n7841), .Z(n7839) );
  OR U15884 ( .A(n7842), .B(n7843), .Z(n7838) );
  NAND U15885 ( .A(n7844), .B(n7845), .Z(n7736) );
  OR U15886 ( .A(n7846), .B(n7847), .Z(n7845) );
  OR U15887 ( .A(n7848), .B(n7849), .Z(n7844) );
  ANDN U15888 ( .B(n7850), .A(n7851), .Z(n7737) );
  IV U15889 ( .A(n7852), .Z(n7850) );
  XNOR U15890 ( .A(n7817), .B(n7816), .Z(N64700) );
  XOR U15891 ( .A(n7836), .B(n7835), .Z(n7816) );
  XNOR U15892 ( .A(n7851), .B(n7852), .Z(n7835) );
  XNOR U15893 ( .A(n7846), .B(n7847), .Z(n7852) );
  XNOR U15894 ( .A(n7848), .B(n7849), .Z(n7847) );
  XNOR U15895 ( .A(y[7597]), .B(x[7597]), .Z(n7849) );
  XNOR U15896 ( .A(y[7598]), .B(x[7598]), .Z(n7848) );
  XNOR U15897 ( .A(y[7596]), .B(x[7596]), .Z(n7846) );
  XNOR U15898 ( .A(n7840), .B(n7841), .Z(n7851) );
  XNOR U15899 ( .A(y[7593]), .B(x[7593]), .Z(n7841) );
  XNOR U15900 ( .A(n7842), .B(n7843), .Z(n7840) );
  XNOR U15901 ( .A(y[7594]), .B(x[7594]), .Z(n7843) );
  XNOR U15902 ( .A(y[7595]), .B(x[7595]), .Z(n7842) );
  XNOR U15903 ( .A(n7833), .B(n7832), .Z(n7836) );
  XNOR U15904 ( .A(n7828), .B(n7829), .Z(n7832) );
  XNOR U15905 ( .A(y[7590]), .B(x[7590]), .Z(n7829) );
  XNOR U15906 ( .A(n7830), .B(n7831), .Z(n7828) );
  XNOR U15907 ( .A(y[7591]), .B(x[7591]), .Z(n7831) );
  XNOR U15908 ( .A(y[7592]), .B(x[7592]), .Z(n7830) );
  XNOR U15909 ( .A(n7822), .B(n7823), .Z(n7833) );
  XNOR U15910 ( .A(y[7587]), .B(x[7587]), .Z(n7823) );
  XNOR U15911 ( .A(n7824), .B(n7825), .Z(n7822) );
  XNOR U15912 ( .A(y[7588]), .B(x[7588]), .Z(n7825) );
  XNOR U15913 ( .A(y[7589]), .B(x[7589]), .Z(n7824) );
  XOR U15914 ( .A(n7798), .B(n7799), .Z(n7817) );
  XNOR U15915 ( .A(n7814), .B(n7815), .Z(n7799) );
  XNOR U15916 ( .A(n7809), .B(n7810), .Z(n7815) );
  XNOR U15917 ( .A(n7811), .B(n7812), .Z(n7810) );
  XNOR U15918 ( .A(y[7585]), .B(x[7585]), .Z(n7812) );
  XNOR U15919 ( .A(y[7586]), .B(x[7586]), .Z(n7811) );
  XNOR U15920 ( .A(y[7584]), .B(x[7584]), .Z(n7809) );
  XNOR U15921 ( .A(n7803), .B(n7804), .Z(n7814) );
  XNOR U15922 ( .A(y[7581]), .B(x[7581]), .Z(n7804) );
  XNOR U15923 ( .A(n7805), .B(n7806), .Z(n7803) );
  XNOR U15924 ( .A(y[7582]), .B(x[7582]), .Z(n7806) );
  XNOR U15925 ( .A(y[7583]), .B(x[7583]), .Z(n7805) );
  XOR U15926 ( .A(n7797), .B(n7796), .Z(n7798) );
  XNOR U15927 ( .A(n7792), .B(n7793), .Z(n7796) );
  XNOR U15928 ( .A(y[7578]), .B(x[7578]), .Z(n7793) );
  XNOR U15929 ( .A(n7794), .B(n7795), .Z(n7792) );
  XNOR U15930 ( .A(y[7579]), .B(x[7579]), .Z(n7795) );
  XNOR U15931 ( .A(y[7580]), .B(x[7580]), .Z(n7794) );
  XNOR U15932 ( .A(n7786), .B(n7787), .Z(n7797) );
  XNOR U15933 ( .A(y[7575]), .B(x[7575]), .Z(n7787) );
  XNOR U15934 ( .A(n7788), .B(n7789), .Z(n7786) );
  XNOR U15935 ( .A(y[7576]), .B(x[7576]), .Z(n7789) );
  XNOR U15936 ( .A(y[7577]), .B(x[7577]), .Z(n7788) );
  NAND U15937 ( .A(n7853), .B(n7854), .Z(N64691) );
  NANDN U15938 ( .A(n7855), .B(n7856), .Z(n7854) );
  OR U15939 ( .A(n7857), .B(n7858), .Z(n7856) );
  NAND U15940 ( .A(n7857), .B(n7858), .Z(n7853) );
  XOR U15941 ( .A(n7857), .B(n7859), .Z(N64690) );
  XNOR U15942 ( .A(n7855), .B(n7858), .Z(n7859) );
  AND U15943 ( .A(n7860), .B(n7861), .Z(n7858) );
  NANDN U15944 ( .A(n7862), .B(n7863), .Z(n7861) );
  NANDN U15945 ( .A(n7864), .B(n7865), .Z(n7863) );
  NANDN U15946 ( .A(n7865), .B(n7864), .Z(n7860) );
  NAND U15947 ( .A(n7866), .B(n7867), .Z(n7855) );
  NANDN U15948 ( .A(n7868), .B(n7869), .Z(n7867) );
  OR U15949 ( .A(n7870), .B(n7871), .Z(n7869) );
  NAND U15950 ( .A(n7871), .B(n7870), .Z(n7866) );
  AND U15951 ( .A(n7872), .B(n7873), .Z(n7857) );
  NANDN U15952 ( .A(n7874), .B(n7875), .Z(n7873) );
  NANDN U15953 ( .A(n7876), .B(n7877), .Z(n7875) );
  NANDN U15954 ( .A(n7877), .B(n7876), .Z(n7872) );
  XOR U15955 ( .A(n7871), .B(n7878), .Z(N64689) );
  XOR U15956 ( .A(n7868), .B(n7870), .Z(n7878) );
  XNOR U15957 ( .A(n7864), .B(n7879), .Z(n7870) );
  XNOR U15958 ( .A(n7862), .B(n7865), .Z(n7879) );
  NAND U15959 ( .A(n7880), .B(n7881), .Z(n7865) );
  NAND U15960 ( .A(n7882), .B(n7883), .Z(n7881) );
  OR U15961 ( .A(n7884), .B(n7885), .Z(n7882) );
  NANDN U15962 ( .A(n7886), .B(n7884), .Z(n7880) );
  IV U15963 ( .A(n7885), .Z(n7886) );
  NAND U15964 ( .A(n7887), .B(n7888), .Z(n7862) );
  NAND U15965 ( .A(n7889), .B(n7890), .Z(n7888) );
  NANDN U15966 ( .A(n7891), .B(n7892), .Z(n7889) );
  NANDN U15967 ( .A(n7892), .B(n7891), .Z(n7887) );
  AND U15968 ( .A(n7893), .B(n7894), .Z(n7864) );
  NAND U15969 ( .A(n7895), .B(n7896), .Z(n7894) );
  OR U15970 ( .A(n7897), .B(n7898), .Z(n7895) );
  NANDN U15971 ( .A(n7899), .B(n7897), .Z(n7893) );
  NAND U15972 ( .A(n7900), .B(n7901), .Z(n7868) );
  NANDN U15973 ( .A(n7902), .B(n7903), .Z(n7901) );
  OR U15974 ( .A(n7904), .B(n7905), .Z(n7903) );
  NANDN U15975 ( .A(n7906), .B(n7904), .Z(n7900) );
  IV U15976 ( .A(n7905), .Z(n7906) );
  XNOR U15977 ( .A(n7876), .B(n7907), .Z(n7871) );
  XNOR U15978 ( .A(n7874), .B(n7877), .Z(n7907) );
  NAND U15979 ( .A(n7908), .B(n7909), .Z(n7877) );
  NAND U15980 ( .A(n7910), .B(n7911), .Z(n7909) );
  OR U15981 ( .A(n7912), .B(n7913), .Z(n7910) );
  NANDN U15982 ( .A(n7914), .B(n7912), .Z(n7908) );
  IV U15983 ( .A(n7913), .Z(n7914) );
  NAND U15984 ( .A(n7915), .B(n7916), .Z(n7874) );
  NAND U15985 ( .A(n7917), .B(n7918), .Z(n7916) );
  NANDN U15986 ( .A(n7919), .B(n7920), .Z(n7917) );
  NANDN U15987 ( .A(n7920), .B(n7919), .Z(n7915) );
  AND U15988 ( .A(n7921), .B(n7922), .Z(n7876) );
  NAND U15989 ( .A(n7923), .B(n7924), .Z(n7922) );
  OR U15990 ( .A(n7925), .B(n7926), .Z(n7923) );
  NANDN U15991 ( .A(n7927), .B(n7925), .Z(n7921) );
  XNOR U15992 ( .A(n7902), .B(n7928), .Z(N64688) );
  XOR U15993 ( .A(n7904), .B(n7905), .Z(n7928) );
  XNOR U15994 ( .A(n7918), .B(n7929), .Z(n7905) );
  XOR U15995 ( .A(n7919), .B(n7920), .Z(n7929) );
  XOR U15996 ( .A(n7925), .B(n7930), .Z(n7920) );
  XOR U15997 ( .A(n7924), .B(n7927), .Z(n7930) );
  IV U15998 ( .A(n7926), .Z(n7927) );
  NAND U15999 ( .A(n7931), .B(n7932), .Z(n7926) );
  OR U16000 ( .A(n7933), .B(n7934), .Z(n7932) );
  OR U16001 ( .A(n7935), .B(n7936), .Z(n7931) );
  NAND U16002 ( .A(n7937), .B(n7938), .Z(n7924) );
  OR U16003 ( .A(n7939), .B(n7940), .Z(n7938) );
  OR U16004 ( .A(n7941), .B(n7942), .Z(n7937) );
  NOR U16005 ( .A(n7943), .B(n7944), .Z(n7925) );
  ANDN U16006 ( .B(n7945), .A(n7946), .Z(n7919) );
  XNOR U16007 ( .A(n7912), .B(n7947), .Z(n7918) );
  XNOR U16008 ( .A(n7911), .B(n7913), .Z(n7947) );
  NAND U16009 ( .A(n7948), .B(n7949), .Z(n7913) );
  OR U16010 ( .A(n7950), .B(n7951), .Z(n7949) );
  OR U16011 ( .A(n7952), .B(n7953), .Z(n7948) );
  NAND U16012 ( .A(n7954), .B(n7955), .Z(n7911) );
  OR U16013 ( .A(n7956), .B(n7957), .Z(n7955) );
  OR U16014 ( .A(n7958), .B(n7959), .Z(n7954) );
  ANDN U16015 ( .B(n7960), .A(n7961), .Z(n7912) );
  IV U16016 ( .A(n7962), .Z(n7960) );
  ANDN U16017 ( .B(n7963), .A(n7964), .Z(n7904) );
  XOR U16018 ( .A(n7890), .B(n7965), .Z(n7902) );
  XOR U16019 ( .A(n7891), .B(n7892), .Z(n7965) );
  XOR U16020 ( .A(n7897), .B(n7966), .Z(n7892) );
  XOR U16021 ( .A(n7896), .B(n7899), .Z(n7966) );
  IV U16022 ( .A(n7898), .Z(n7899) );
  NAND U16023 ( .A(n7967), .B(n7968), .Z(n7898) );
  OR U16024 ( .A(n7969), .B(n7970), .Z(n7968) );
  OR U16025 ( .A(n7971), .B(n7972), .Z(n7967) );
  NAND U16026 ( .A(n7973), .B(n7974), .Z(n7896) );
  OR U16027 ( .A(n7975), .B(n7976), .Z(n7974) );
  OR U16028 ( .A(n7977), .B(n7978), .Z(n7973) );
  NOR U16029 ( .A(n7979), .B(n7980), .Z(n7897) );
  ANDN U16030 ( .B(n7981), .A(n7982), .Z(n7891) );
  IV U16031 ( .A(n7983), .Z(n7981) );
  XNOR U16032 ( .A(n7884), .B(n7984), .Z(n7890) );
  XNOR U16033 ( .A(n7883), .B(n7885), .Z(n7984) );
  NAND U16034 ( .A(n7985), .B(n7986), .Z(n7885) );
  OR U16035 ( .A(n7987), .B(n7988), .Z(n7986) );
  OR U16036 ( .A(n7989), .B(n7990), .Z(n7985) );
  NAND U16037 ( .A(n7991), .B(n7992), .Z(n7883) );
  OR U16038 ( .A(n7993), .B(n7994), .Z(n7992) );
  OR U16039 ( .A(n7995), .B(n7996), .Z(n7991) );
  ANDN U16040 ( .B(n7997), .A(n7998), .Z(n7884) );
  IV U16041 ( .A(n7999), .Z(n7997) );
  XNOR U16042 ( .A(n7964), .B(n7963), .Z(N64687) );
  XOR U16043 ( .A(n7983), .B(n7982), .Z(n7963) );
  XNOR U16044 ( .A(n7998), .B(n7999), .Z(n7982) );
  XNOR U16045 ( .A(n7993), .B(n7994), .Z(n7999) );
  XNOR U16046 ( .A(n7995), .B(n7996), .Z(n7994) );
  XNOR U16047 ( .A(y[7573]), .B(x[7573]), .Z(n7996) );
  XNOR U16048 ( .A(y[7574]), .B(x[7574]), .Z(n7995) );
  XNOR U16049 ( .A(y[7572]), .B(x[7572]), .Z(n7993) );
  XNOR U16050 ( .A(n7987), .B(n7988), .Z(n7998) );
  XNOR U16051 ( .A(y[7569]), .B(x[7569]), .Z(n7988) );
  XNOR U16052 ( .A(n7989), .B(n7990), .Z(n7987) );
  XNOR U16053 ( .A(y[7570]), .B(x[7570]), .Z(n7990) );
  XNOR U16054 ( .A(y[7571]), .B(x[7571]), .Z(n7989) );
  XNOR U16055 ( .A(n7980), .B(n7979), .Z(n7983) );
  XNOR U16056 ( .A(n7975), .B(n7976), .Z(n7979) );
  XNOR U16057 ( .A(y[7566]), .B(x[7566]), .Z(n7976) );
  XNOR U16058 ( .A(n7977), .B(n7978), .Z(n7975) );
  XNOR U16059 ( .A(y[7567]), .B(x[7567]), .Z(n7978) );
  XNOR U16060 ( .A(y[7568]), .B(x[7568]), .Z(n7977) );
  XNOR U16061 ( .A(n7969), .B(n7970), .Z(n7980) );
  XNOR U16062 ( .A(y[7563]), .B(x[7563]), .Z(n7970) );
  XNOR U16063 ( .A(n7971), .B(n7972), .Z(n7969) );
  XNOR U16064 ( .A(y[7564]), .B(x[7564]), .Z(n7972) );
  XNOR U16065 ( .A(y[7565]), .B(x[7565]), .Z(n7971) );
  XOR U16066 ( .A(n7945), .B(n7946), .Z(n7964) );
  XNOR U16067 ( .A(n7961), .B(n7962), .Z(n7946) );
  XNOR U16068 ( .A(n7956), .B(n7957), .Z(n7962) );
  XNOR U16069 ( .A(n7958), .B(n7959), .Z(n7957) );
  XNOR U16070 ( .A(y[7561]), .B(x[7561]), .Z(n7959) );
  XNOR U16071 ( .A(y[7562]), .B(x[7562]), .Z(n7958) );
  XNOR U16072 ( .A(y[7560]), .B(x[7560]), .Z(n7956) );
  XNOR U16073 ( .A(n7950), .B(n7951), .Z(n7961) );
  XNOR U16074 ( .A(y[7557]), .B(x[7557]), .Z(n7951) );
  XNOR U16075 ( .A(n7952), .B(n7953), .Z(n7950) );
  XNOR U16076 ( .A(y[7558]), .B(x[7558]), .Z(n7953) );
  XNOR U16077 ( .A(y[7559]), .B(x[7559]), .Z(n7952) );
  XOR U16078 ( .A(n7944), .B(n7943), .Z(n7945) );
  XNOR U16079 ( .A(n7939), .B(n7940), .Z(n7943) );
  XNOR U16080 ( .A(y[7554]), .B(x[7554]), .Z(n7940) );
  XNOR U16081 ( .A(n7941), .B(n7942), .Z(n7939) );
  XNOR U16082 ( .A(y[7555]), .B(x[7555]), .Z(n7942) );
  XNOR U16083 ( .A(y[7556]), .B(x[7556]), .Z(n7941) );
  XNOR U16084 ( .A(n7933), .B(n7934), .Z(n7944) );
  XNOR U16085 ( .A(y[7551]), .B(x[7551]), .Z(n7934) );
  XNOR U16086 ( .A(n7935), .B(n7936), .Z(n7933) );
  XNOR U16087 ( .A(y[7552]), .B(x[7552]), .Z(n7936) );
  XNOR U16088 ( .A(y[7553]), .B(x[7553]), .Z(n7935) );
  NAND U16089 ( .A(n8000), .B(n8001), .Z(N64678) );
  NANDN U16090 ( .A(n8002), .B(n8003), .Z(n8001) );
  OR U16091 ( .A(n8004), .B(n8005), .Z(n8003) );
  NAND U16092 ( .A(n8004), .B(n8005), .Z(n8000) );
  XOR U16093 ( .A(n8004), .B(n8006), .Z(N64677) );
  XNOR U16094 ( .A(n8002), .B(n8005), .Z(n8006) );
  AND U16095 ( .A(n8007), .B(n8008), .Z(n8005) );
  NANDN U16096 ( .A(n8009), .B(n8010), .Z(n8008) );
  NANDN U16097 ( .A(n8011), .B(n8012), .Z(n8010) );
  NANDN U16098 ( .A(n8012), .B(n8011), .Z(n8007) );
  NAND U16099 ( .A(n8013), .B(n8014), .Z(n8002) );
  NANDN U16100 ( .A(n8015), .B(n8016), .Z(n8014) );
  OR U16101 ( .A(n8017), .B(n8018), .Z(n8016) );
  NAND U16102 ( .A(n8018), .B(n8017), .Z(n8013) );
  AND U16103 ( .A(n8019), .B(n8020), .Z(n8004) );
  NANDN U16104 ( .A(n8021), .B(n8022), .Z(n8020) );
  NANDN U16105 ( .A(n8023), .B(n8024), .Z(n8022) );
  NANDN U16106 ( .A(n8024), .B(n8023), .Z(n8019) );
  XOR U16107 ( .A(n8018), .B(n8025), .Z(N64676) );
  XOR U16108 ( .A(n8015), .B(n8017), .Z(n8025) );
  XNOR U16109 ( .A(n8011), .B(n8026), .Z(n8017) );
  XNOR U16110 ( .A(n8009), .B(n8012), .Z(n8026) );
  NAND U16111 ( .A(n8027), .B(n8028), .Z(n8012) );
  NAND U16112 ( .A(n8029), .B(n8030), .Z(n8028) );
  OR U16113 ( .A(n8031), .B(n8032), .Z(n8029) );
  NANDN U16114 ( .A(n8033), .B(n8031), .Z(n8027) );
  IV U16115 ( .A(n8032), .Z(n8033) );
  NAND U16116 ( .A(n8034), .B(n8035), .Z(n8009) );
  NAND U16117 ( .A(n8036), .B(n8037), .Z(n8035) );
  NANDN U16118 ( .A(n8038), .B(n8039), .Z(n8036) );
  NANDN U16119 ( .A(n8039), .B(n8038), .Z(n8034) );
  AND U16120 ( .A(n8040), .B(n8041), .Z(n8011) );
  NAND U16121 ( .A(n8042), .B(n8043), .Z(n8041) );
  OR U16122 ( .A(n8044), .B(n8045), .Z(n8042) );
  NANDN U16123 ( .A(n8046), .B(n8044), .Z(n8040) );
  NAND U16124 ( .A(n8047), .B(n8048), .Z(n8015) );
  NANDN U16125 ( .A(n8049), .B(n8050), .Z(n8048) );
  OR U16126 ( .A(n8051), .B(n8052), .Z(n8050) );
  NANDN U16127 ( .A(n8053), .B(n8051), .Z(n8047) );
  IV U16128 ( .A(n8052), .Z(n8053) );
  XNOR U16129 ( .A(n8023), .B(n8054), .Z(n8018) );
  XNOR U16130 ( .A(n8021), .B(n8024), .Z(n8054) );
  NAND U16131 ( .A(n8055), .B(n8056), .Z(n8024) );
  NAND U16132 ( .A(n8057), .B(n8058), .Z(n8056) );
  OR U16133 ( .A(n8059), .B(n8060), .Z(n8057) );
  NANDN U16134 ( .A(n8061), .B(n8059), .Z(n8055) );
  IV U16135 ( .A(n8060), .Z(n8061) );
  NAND U16136 ( .A(n8062), .B(n8063), .Z(n8021) );
  NAND U16137 ( .A(n8064), .B(n8065), .Z(n8063) );
  NANDN U16138 ( .A(n8066), .B(n8067), .Z(n8064) );
  NANDN U16139 ( .A(n8067), .B(n8066), .Z(n8062) );
  AND U16140 ( .A(n8068), .B(n8069), .Z(n8023) );
  NAND U16141 ( .A(n8070), .B(n8071), .Z(n8069) );
  OR U16142 ( .A(n8072), .B(n8073), .Z(n8070) );
  NANDN U16143 ( .A(n8074), .B(n8072), .Z(n8068) );
  XNOR U16144 ( .A(n8049), .B(n8075), .Z(N64675) );
  XOR U16145 ( .A(n8051), .B(n8052), .Z(n8075) );
  XNOR U16146 ( .A(n8065), .B(n8076), .Z(n8052) );
  XOR U16147 ( .A(n8066), .B(n8067), .Z(n8076) );
  XOR U16148 ( .A(n8072), .B(n8077), .Z(n8067) );
  XOR U16149 ( .A(n8071), .B(n8074), .Z(n8077) );
  IV U16150 ( .A(n8073), .Z(n8074) );
  NAND U16151 ( .A(n8078), .B(n8079), .Z(n8073) );
  OR U16152 ( .A(n8080), .B(n8081), .Z(n8079) );
  OR U16153 ( .A(n8082), .B(n8083), .Z(n8078) );
  NAND U16154 ( .A(n8084), .B(n8085), .Z(n8071) );
  OR U16155 ( .A(n8086), .B(n8087), .Z(n8085) );
  OR U16156 ( .A(n8088), .B(n8089), .Z(n8084) );
  NOR U16157 ( .A(n8090), .B(n8091), .Z(n8072) );
  ANDN U16158 ( .B(n8092), .A(n8093), .Z(n8066) );
  XNOR U16159 ( .A(n8059), .B(n8094), .Z(n8065) );
  XNOR U16160 ( .A(n8058), .B(n8060), .Z(n8094) );
  NAND U16161 ( .A(n8095), .B(n8096), .Z(n8060) );
  OR U16162 ( .A(n8097), .B(n8098), .Z(n8096) );
  OR U16163 ( .A(n8099), .B(n8100), .Z(n8095) );
  NAND U16164 ( .A(n8101), .B(n8102), .Z(n8058) );
  OR U16165 ( .A(n8103), .B(n8104), .Z(n8102) );
  OR U16166 ( .A(n8105), .B(n8106), .Z(n8101) );
  ANDN U16167 ( .B(n8107), .A(n8108), .Z(n8059) );
  IV U16168 ( .A(n8109), .Z(n8107) );
  ANDN U16169 ( .B(n8110), .A(n8111), .Z(n8051) );
  XOR U16170 ( .A(n8037), .B(n8112), .Z(n8049) );
  XOR U16171 ( .A(n8038), .B(n8039), .Z(n8112) );
  XOR U16172 ( .A(n8044), .B(n8113), .Z(n8039) );
  XOR U16173 ( .A(n8043), .B(n8046), .Z(n8113) );
  IV U16174 ( .A(n8045), .Z(n8046) );
  NAND U16175 ( .A(n8114), .B(n8115), .Z(n8045) );
  OR U16176 ( .A(n8116), .B(n8117), .Z(n8115) );
  OR U16177 ( .A(n8118), .B(n8119), .Z(n8114) );
  NAND U16178 ( .A(n8120), .B(n8121), .Z(n8043) );
  OR U16179 ( .A(n8122), .B(n8123), .Z(n8121) );
  OR U16180 ( .A(n8124), .B(n8125), .Z(n8120) );
  NOR U16181 ( .A(n8126), .B(n8127), .Z(n8044) );
  ANDN U16182 ( .B(n8128), .A(n8129), .Z(n8038) );
  IV U16183 ( .A(n8130), .Z(n8128) );
  XNOR U16184 ( .A(n8031), .B(n8131), .Z(n8037) );
  XNOR U16185 ( .A(n8030), .B(n8032), .Z(n8131) );
  NAND U16186 ( .A(n8132), .B(n8133), .Z(n8032) );
  OR U16187 ( .A(n8134), .B(n8135), .Z(n8133) );
  OR U16188 ( .A(n8136), .B(n8137), .Z(n8132) );
  NAND U16189 ( .A(n8138), .B(n8139), .Z(n8030) );
  OR U16190 ( .A(n8140), .B(n8141), .Z(n8139) );
  OR U16191 ( .A(n8142), .B(n8143), .Z(n8138) );
  ANDN U16192 ( .B(n8144), .A(n8145), .Z(n8031) );
  IV U16193 ( .A(n8146), .Z(n8144) );
  XNOR U16194 ( .A(n8111), .B(n8110), .Z(N64674) );
  XOR U16195 ( .A(n8130), .B(n8129), .Z(n8110) );
  XNOR U16196 ( .A(n8145), .B(n8146), .Z(n8129) );
  XNOR U16197 ( .A(n8140), .B(n8141), .Z(n8146) );
  XNOR U16198 ( .A(n8142), .B(n8143), .Z(n8141) );
  XNOR U16199 ( .A(y[7549]), .B(x[7549]), .Z(n8143) );
  XNOR U16200 ( .A(y[7550]), .B(x[7550]), .Z(n8142) );
  XNOR U16201 ( .A(y[7548]), .B(x[7548]), .Z(n8140) );
  XNOR U16202 ( .A(n8134), .B(n8135), .Z(n8145) );
  XNOR U16203 ( .A(y[7545]), .B(x[7545]), .Z(n8135) );
  XNOR U16204 ( .A(n8136), .B(n8137), .Z(n8134) );
  XNOR U16205 ( .A(y[7546]), .B(x[7546]), .Z(n8137) );
  XNOR U16206 ( .A(y[7547]), .B(x[7547]), .Z(n8136) );
  XNOR U16207 ( .A(n8127), .B(n8126), .Z(n8130) );
  XNOR U16208 ( .A(n8122), .B(n8123), .Z(n8126) );
  XNOR U16209 ( .A(y[7542]), .B(x[7542]), .Z(n8123) );
  XNOR U16210 ( .A(n8124), .B(n8125), .Z(n8122) );
  XNOR U16211 ( .A(y[7543]), .B(x[7543]), .Z(n8125) );
  XNOR U16212 ( .A(y[7544]), .B(x[7544]), .Z(n8124) );
  XNOR U16213 ( .A(n8116), .B(n8117), .Z(n8127) );
  XNOR U16214 ( .A(y[7539]), .B(x[7539]), .Z(n8117) );
  XNOR U16215 ( .A(n8118), .B(n8119), .Z(n8116) );
  XNOR U16216 ( .A(y[7540]), .B(x[7540]), .Z(n8119) );
  XNOR U16217 ( .A(y[7541]), .B(x[7541]), .Z(n8118) );
  XOR U16218 ( .A(n8092), .B(n8093), .Z(n8111) );
  XNOR U16219 ( .A(n8108), .B(n8109), .Z(n8093) );
  XNOR U16220 ( .A(n8103), .B(n8104), .Z(n8109) );
  XNOR U16221 ( .A(n8105), .B(n8106), .Z(n8104) );
  XNOR U16222 ( .A(y[7537]), .B(x[7537]), .Z(n8106) );
  XNOR U16223 ( .A(y[7538]), .B(x[7538]), .Z(n8105) );
  XNOR U16224 ( .A(y[7536]), .B(x[7536]), .Z(n8103) );
  XNOR U16225 ( .A(n8097), .B(n8098), .Z(n8108) );
  XNOR U16226 ( .A(y[7533]), .B(x[7533]), .Z(n8098) );
  XNOR U16227 ( .A(n8099), .B(n8100), .Z(n8097) );
  XNOR U16228 ( .A(y[7534]), .B(x[7534]), .Z(n8100) );
  XNOR U16229 ( .A(y[7535]), .B(x[7535]), .Z(n8099) );
  XOR U16230 ( .A(n8091), .B(n8090), .Z(n8092) );
  XNOR U16231 ( .A(n8086), .B(n8087), .Z(n8090) );
  XNOR U16232 ( .A(y[7530]), .B(x[7530]), .Z(n8087) );
  XNOR U16233 ( .A(n8088), .B(n8089), .Z(n8086) );
  XNOR U16234 ( .A(y[7531]), .B(x[7531]), .Z(n8089) );
  XNOR U16235 ( .A(y[7532]), .B(x[7532]), .Z(n8088) );
  XNOR U16236 ( .A(n8080), .B(n8081), .Z(n8091) );
  XNOR U16237 ( .A(y[7527]), .B(x[7527]), .Z(n8081) );
  XNOR U16238 ( .A(n8082), .B(n8083), .Z(n8080) );
  XNOR U16239 ( .A(y[7528]), .B(x[7528]), .Z(n8083) );
  XNOR U16240 ( .A(y[7529]), .B(x[7529]), .Z(n8082) );
  NAND U16241 ( .A(n8147), .B(n8148), .Z(N64665) );
  NANDN U16242 ( .A(n8149), .B(n8150), .Z(n8148) );
  OR U16243 ( .A(n8151), .B(n8152), .Z(n8150) );
  NAND U16244 ( .A(n8151), .B(n8152), .Z(n8147) );
  XOR U16245 ( .A(n8151), .B(n8153), .Z(N64664) );
  XNOR U16246 ( .A(n8149), .B(n8152), .Z(n8153) );
  AND U16247 ( .A(n8154), .B(n8155), .Z(n8152) );
  NANDN U16248 ( .A(n8156), .B(n8157), .Z(n8155) );
  NANDN U16249 ( .A(n8158), .B(n8159), .Z(n8157) );
  NANDN U16250 ( .A(n8159), .B(n8158), .Z(n8154) );
  NAND U16251 ( .A(n8160), .B(n8161), .Z(n8149) );
  NANDN U16252 ( .A(n8162), .B(n8163), .Z(n8161) );
  OR U16253 ( .A(n8164), .B(n8165), .Z(n8163) );
  NAND U16254 ( .A(n8165), .B(n8164), .Z(n8160) );
  AND U16255 ( .A(n8166), .B(n8167), .Z(n8151) );
  NANDN U16256 ( .A(n8168), .B(n8169), .Z(n8167) );
  NANDN U16257 ( .A(n8170), .B(n8171), .Z(n8169) );
  NANDN U16258 ( .A(n8171), .B(n8170), .Z(n8166) );
  XOR U16259 ( .A(n8165), .B(n8172), .Z(N64663) );
  XOR U16260 ( .A(n8162), .B(n8164), .Z(n8172) );
  XNOR U16261 ( .A(n8158), .B(n8173), .Z(n8164) );
  XNOR U16262 ( .A(n8156), .B(n8159), .Z(n8173) );
  NAND U16263 ( .A(n8174), .B(n8175), .Z(n8159) );
  NAND U16264 ( .A(n8176), .B(n8177), .Z(n8175) );
  OR U16265 ( .A(n8178), .B(n8179), .Z(n8176) );
  NANDN U16266 ( .A(n8180), .B(n8178), .Z(n8174) );
  IV U16267 ( .A(n8179), .Z(n8180) );
  NAND U16268 ( .A(n8181), .B(n8182), .Z(n8156) );
  NAND U16269 ( .A(n8183), .B(n8184), .Z(n8182) );
  NANDN U16270 ( .A(n8185), .B(n8186), .Z(n8183) );
  NANDN U16271 ( .A(n8186), .B(n8185), .Z(n8181) );
  AND U16272 ( .A(n8187), .B(n8188), .Z(n8158) );
  NAND U16273 ( .A(n8189), .B(n8190), .Z(n8188) );
  OR U16274 ( .A(n8191), .B(n8192), .Z(n8189) );
  NANDN U16275 ( .A(n8193), .B(n8191), .Z(n8187) );
  NAND U16276 ( .A(n8194), .B(n8195), .Z(n8162) );
  NANDN U16277 ( .A(n8196), .B(n8197), .Z(n8195) );
  OR U16278 ( .A(n8198), .B(n8199), .Z(n8197) );
  NANDN U16279 ( .A(n8200), .B(n8198), .Z(n8194) );
  IV U16280 ( .A(n8199), .Z(n8200) );
  XNOR U16281 ( .A(n8170), .B(n8201), .Z(n8165) );
  XNOR U16282 ( .A(n8168), .B(n8171), .Z(n8201) );
  NAND U16283 ( .A(n8202), .B(n8203), .Z(n8171) );
  NAND U16284 ( .A(n8204), .B(n8205), .Z(n8203) );
  OR U16285 ( .A(n8206), .B(n8207), .Z(n8204) );
  NANDN U16286 ( .A(n8208), .B(n8206), .Z(n8202) );
  IV U16287 ( .A(n8207), .Z(n8208) );
  NAND U16288 ( .A(n8209), .B(n8210), .Z(n8168) );
  NAND U16289 ( .A(n8211), .B(n8212), .Z(n8210) );
  NANDN U16290 ( .A(n8213), .B(n8214), .Z(n8211) );
  NANDN U16291 ( .A(n8214), .B(n8213), .Z(n8209) );
  AND U16292 ( .A(n8215), .B(n8216), .Z(n8170) );
  NAND U16293 ( .A(n8217), .B(n8218), .Z(n8216) );
  OR U16294 ( .A(n8219), .B(n8220), .Z(n8217) );
  NANDN U16295 ( .A(n8221), .B(n8219), .Z(n8215) );
  XNOR U16296 ( .A(n8196), .B(n8222), .Z(N64662) );
  XOR U16297 ( .A(n8198), .B(n8199), .Z(n8222) );
  XNOR U16298 ( .A(n8212), .B(n8223), .Z(n8199) );
  XOR U16299 ( .A(n8213), .B(n8214), .Z(n8223) );
  XOR U16300 ( .A(n8219), .B(n8224), .Z(n8214) );
  XOR U16301 ( .A(n8218), .B(n8221), .Z(n8224) );
  IV U16302 ( .A(n8220), .Z(n8221) );
  NAND U16303 ( .A(n8225), .B(n8226), .Z(n8220) );
  OR U16304 ( .A(n8227), .B(n8228), .Z(n8226) );
  OR U16305 ( .A(n8229), .B(n8230), .Z(n8225) );
  NAND U16306 ( .A(n8231), .B(n8232), .Z(n8218) );
  OR U16307 ( .A(n8233), .B(n8234), .Z(n8232) );
  OR U16308 ( .A(n8235), .B(n8236), .Z(n8231) );
  NOR U16309 ( .A(n8237), .B(n8238), .Z(n8219) );
  ANDN U16310 ( .B(n8239), .A(n8240), .Z(n8213) );
  XNOR U16311 ( .A(n8206), .B(n8241), .Z(n8212) );
  XNOR U16312 ( .A(n8205), .B(n8207), .Z(n8241) );
  NAND U16313 ( .A(n8242), .B(n8243), .Z(n8207) );
  OR U16314 ( .A(n8244), .B(n8245), .Z(n8243) );
  OR U16315 ( .A(n8246), .B(n8247), .Z(n8242) );
  NAND U16316 ( .A(n8248), .B(n8249), .Z(n8205) );
  OR U16317 ( .A(n8250), .B(n8251), .Z(n8249) );
  OR U16318 ( .A(n8252), .B(n8253), .Z(n8248) );
  ANDN U16319 ( .B(n8254), .A(n8255), .Z(n8206) );
  IV U16320 ( .A(n8256), .Z(n8254) );
  ANDN U16321 ( .B(n8257), .A(n8258), .Z(n8198) );
  XOR U16322 ( .A(n8184), .B(n8259), .Z(n8196) );
  XOR U16323 ( .A(n8185), .B(n8186), .Z(n8259) );
  XOR U16324 ( .A(n8191), .B(n8260), .Z(n8186) );
  XOR U16325 ( .A(n8190), .B(n8193), .Z(n8260) );
  IV U16326 ( .A(n8192), .Z(n8193) );
  NAND U16327 ( .A(n8261), .B(n8262), .Z(n8192) );
  OR U16328 ( .A(n8263), .B(n8264), .Z(n8262) );
  OR U16329 ( .A(n8265), .B(n8266), .Z(n8261) );
  NAND U16330 ( .A(n8267), .B(n8268), .Z(n8190) );
  OR U16331 ( .A(n8269), .B(n8270), .Z(n8268) );
  OR U16332 ( .A(n8271), .B(n8272), .Z(n8267) );
  NOR U16333 ( .A(n8273), .B(n8274), .Z(n8191) );
  ANDN U16334 ( .B(n8275), .A(n8276), .Z(n8185) );
  IV U16335 ( .A(n8277), .Z(n8275) );
  XNOR U16336 ( .A(n8178), .B(n8278), .Z(n8184) );
  XNOR U16337 ( .A(n8177), .B(n8179), .Z(n8278) );
  NAND U16338 ( .A(n8279), .B(n8280), .Z(n8179) );
  OR U16339 ( .A(n8281), .B(n8282), .Z(n8280) );
  OR U16340 ( .A(n8283), .B(n8284), .Z(n8279) );
  NAND U16341 ( .A(n8285), .B(n8286), .Z(n8177) );
  OR U16342 ( .A(n8287), .B(n8288), .Z(n8286) );
  OR U16343 ( .A(n8289), .B(n8290), .Z(n8285) );
  ANDN U16344 ( .B(n8291), .A(n8292), .Z(n8178) );
  IV U16345 ( .A(n8293), .Z(n8291) );
  XNOR U16346 ( .A(n8258), .B(n8257), .Z(N64661) );
  XOR U16347 ( .A(n8277), .B(n8276), .Z(n8257) );
  XNOR U16348 ( .A(n8292), .B(n8293), .Z(n8276) );
  XNOR U16349 ( .A(n8287), .B(n8288), .Z(n8293) );
  XNOR U16350 ( .A(n8289), .B(n8290), .Z(n8288) );
  XNOR U16351 ( .A(y[7525]), .B(x[7525]), .Z(n8290) );
  XNOR U16352 ( .A(y[7526]), .B(x[7526]), .Z(n8289) );
  XNOR U16353 ( .A(y[7524]), .B(x[7524]), .Z(n8287) );
  XNOR U16354 ( .A(n8281), .B(n8282), .Z(n8292) );
  XNOR U16355 ( .A(y[7521]), .B(x[7521]), .Z(n8282) );
  XNOR U16356 ( .A(n8283), .B(n8284), .Z(n8281) );
  XNOR U16357 ( .A(y[7522]), .B(x[7522]), .Z(n8284) );
  XNOR U16358 ( .A(y[7523]), .B(x[7523]), .Z(n8283) );
  XNOR U16359 ( .A(n8274), .B(n8273), .Z(n8277) );
  XNOR U16360 ( .A(n8269), .B(n8270), .Z(n8273) );
  XNOR U16361 ( .A(y[7518]), .B(x[7518]), .Z(n8270) );
  XNOR U16362 ( .A(n8271), .B(n8272), .Z(n8269) );
  XNOR U16363 ( .A(y[7519]), .B(x[7519]), .Z(n8272) );
  XNOR U16364 ( .A(y[7520]), .B(x[7520]), .Z(n8271) );
  XNOR U16365 ( .A(n8263), .B(n8264), .Z(n8274) );
  XNOR U16366 ( .A(y[7515]), .B(x[7515]), .Z(n8264) );
  XNOR U16367 ( .A(n8265), .B(n8266), .Z(n8263) );
  XNOR U16368 ( .A(y[7516]), .B(x[7516]), .Z(n8266) );
  XNOR U16369 ( .A(y[7517]), .B(x[7517]), .Z(n8265) );
  XOR U16370 ( .A(n8239), .B(n8240), .Z(n8258) );
  XNOR U16371 ( .A(n8255), .B(n8256), .Z(n8240) );
  XNOR U16372 ( .A(n8250), .B(n8251), .Z(n8256) );
  XNOR U16373 ( .A(n8252), .B(n8253), .Z(n8251) );
  XNOR U16374 ( .A(y[7513]), .B(x[7513]), .Z(n8253) );
  XNOR U16375 ( .A(y[7514]), .B(x[7514]), .Z(n8252) );
  XNOR U16376 ( .A(y[7512]), .B(x[7512]), .Z(n8250) );
  XNOR U16377 ( .A(n8244), .B(n8245), .Z(n8255) );
  XNOR U16378 ( .A(y[7509]), .B(x[7509]), .Z(n8245) );
  XNOR U16379 ( .A(n8246), .B(n8247), .Z(n8244) );
  XNOR U16380 ( .A(y[7510]), .B(x[7510]), .Z(n8247) );
  XNOR U16381 ( .A(y[7511]), .B(x[7511]), .Z(n8246) );
  XOR U16382 ( .A(n8238), .B(n8237), .Z(n8239) );
  XNOR U16383 ( .A(n8233), .B(n8234), .Z(n8237) );
  XNOR U16384 ( .A(y[7506]), .B(x[7506]), .Z(n8234) );
  XNOR U16385 ( .A(n8235), .B(n8236), .Z(n8233) );
  XNOR U16386 ( .A(y[7507]), .B(x[7507]), .Z(n8236) );
  XNOR U16387 ( .A(y[7508]), .B(x[7508]), .Z(n8235) );
  XNOR U16388 ( .A(n8227), .B(n8228), .Z(n8238) );
  XNOR U16389 ( .A(y[7503]), .B(x[7503]), .Z(n8228) );
  XNOR U16390 ( .A(n8229), .B(n8230), .Z(n8227) );
  XNOR U16391 ( .A(y[7504]), .B(x[7504]), .Z(n8230) );
  XNOR U16392 ( .A(y[7505]), .B(x[7505]), .Z(n8229) );
  NAND U16393 ( .A(n8294), .B(n8295), .Z(N64652) );
  NANDN U16394 ( .A(n8296), .B(n8297), .Z(n8295) );
  OR U16395 ( .A(n8298), .B(n8299), .Z(n8297) );
  NAND U16396 ( .A(n8298), .B(n8299), .Z(n8294) );
  XOR U16397 ( .A(n8298), .B(n8300), .Z(N64651) );
  XNOR U16398 ( .A(n8296), .B(n8299), .Z(n8300) );
  AND U16399 ( .A(n8301), .B(n8302), .Z(n8299) );
  NANDN U16400 ( .A(n8303), .B(n8304), .Z(n8302) );
  NANDN U16401 ( .A(n8305), .B(n8306), .Z(n8304) );
  NANDN U16402 ( .A(n8306), .B(n8305), .Z(n8301) );
  NAND U16403 ( .A(n8307), .B(n8308), .Z(n8296) );
  NANDN U16404 ( .A(n8309), .B(n8310), .Z(n8308) );
  OR U16405 ( .A(n8311), .B(n8312), .Z(n8310) );
  NAND U16406 ( .A(n8312), .B(n8311), .Z(n8307) );
  AND U16407 ( .A(n8313), .B(n8314), .Z(n8298) );
  NANDN U16408 ( .A(n8315), .B(n8316), .Z(n8314) );
  NANDN U16409 ( .A(n8317), .B(n8318), .Z(n8316) );
  NANDN U16410 ( .A(n8318), .B(n8317), .Z(n8313) );
  XOR U16411 ( .A(n8312), .B(n8319), .Z(N64650) );
  XOR U16412 ( .A(n8309), .B(n8311), .Z(n8319) );
  XNOR U16413 ( .A(n8305), .B(n8320), .Z(n8311) );
  XNOR U16414 ( .A(n8303), .B(n8306), .Z(n8320) );
  NAND U16415 ( .A(n8321), .B(n8322), .Z(n8306) );
  NAND U16416 ( .A(n8323), .B(n8324), .Z(n8322) );
  OR U16417 ( .A(n8325), .B(n8326), .Z(n8323) );
  NANDN U16418 ( .A(n8327), .B(n8325), .Z(n8321) );
  IV U16419 ( .A(n8326), .Z(n8327) );
  NAND U16420 ( .A(n8328), .B(n8329), .Z(n8303) );
  NAND U16421 ( .A(n8330), .B(n8331), .Z(n8329) );
  NANDN U16422 ( .A(n8332), .B(n8333), .Z(n8330) );
  NANDN U16423 ( .A(n8333), .B(n8332), .Z(n8328) );
  AND U16424 ( .A(n8334), .B(n8335), .Z(n8305) );
  NAND U16425 ( .A(n8336), .B(n8337), .Z(n8335) );
  OR U16426 ( .A(n8338), .B(n8339), .Z(n8336) );
  NANDN U16427 ( .A(n8340), .B(n8338), .Z(n8334) );
  NAND U16428 ( .A(n8341), .B(n8342), .Z(n8309) );
  NANDN U16429 ( .A(n8343), .B(n8344), .Z(n8342) );
  OR U16430 ( .A(n8345), .B(n8346), .Z(n8344) );
  NANDN U16431 ( .A(n8347), .B(n8345), .Z(n8341) );
  IV U16432 ( .A(n8346), .Z(n8347) );
  XNOR U16433 ( .A(n8317), .B(n8348), .Z(n8312) );
  XNOR U16434 ( .A(n8315), .B(n8318), .Z(n8348) );
  NAND U16435 ( .A(n8349), .B(n8350), .Z(n8318) );
  NAND U16436 ( .A(n8351), .B(n8352), .Z(n8350) );
  OR U16437 ( .A(n8353), .B(n8354), .Z(n8351) );
  NANDN U16438 ( .A(n8355), .B(n8353), .Z(n8349) );
  IV U16439 ( .A(n8354), .Z(n8355) );
  NAND U16440 ( .A(n8356), .B(n8357), .Z(n8315) );
  NAND U16441 ( .A(n8358), .B(n8359), .Z(n8357) );
  NANDN U16442 ( .A(n8360), .B(n8361), .Z(n8358) );
  NANDN U16443 ( .A(n8361), .B(n8360), .Z(n8356) );
  AND U16444 ( .A(n8362), .B(n8363), .Z(n8317) );
  NAND U16445 ( .A(n8364), .B(n8365), .Z(n8363) );
  OR U16446 ( .A(n8366), .B(n8367), .Z(n8364) );
  NANDN U16447 ( .A(n8368), .B(n8366), .Z(n8362) );
  XNOR U16448 ( .A(n8343), .B(n8369), .Z(N64649) );
  XOR U16449 ( .A(n8345), .B(n8346), .Z(n8369) );
  XNOR U16450 ( .A(n8359), .B(n8370), .Z(n8346) );
  XOR U16451 ( .A(n8360), .B(n8361), .Z(n8370) );
  XOR U16452 ( .A(n8366), .B(n8371), .Z(n8361) );
  XOR U16453 ( .A(n8365), .B(n8368), .Z(n8371) );
  IV U16454 ( .A(n8367), .Z(n8368) );
  NAND U16455 ( .A(n8372), .B(n8373), .Z(n8367) );
  OR U16456 ( .A(n8374), .B(n8375), .Z(n8373) );
  OR U16457 ( .A(n8376), .B(n8377), .Z(n8372) );
  NAND U16458 ( .A(n8378), .B(n8379), .Z(n8365) );
  OR U16459 ( .A(n8380), .B(n8381), .Z(n8379) );
  OR U16460 ( .A(n8382), .B(n8383), .Z(n8378) );
  NOR U16461 ( .A(n8384), .B(n8385), .Z(n8366) );
  ANDN U16462 ( .B(n8386), .A(n8387), .Z(n8360) );
  XNOR U16463 ( .A(n8353), .B(n8388), .Z(n8359) );
  XNOR U16464 ( .A(n8352), .B(n8354), .Z(n8388) );
  NAND U16465 ( .A(n8389), .B(n8390), .Z(n8354) );
  OR U16466 ( .A(n8391), .B(n8392), .Z(n8390) );
  OR U16467 ( .A(n8393), .B(n8394), .Z(n8389) );
  NAND U16468 ( .A(n8395), .B(n8396), .Z(n8352) );
  OR U16469 ( .A(n8397), .B(n8398), .Z(n8396) );
  OR U16470 ( .A(n8399), .B(n8400), .Z(n8395) );
  ANDN U16471 ( .B(n8401), .A(n8402), .Z(n8353) );
  IV U16472 ( .A(n8403), .Z(n8401) );
  ANDN U16473 ( .B(n8404), .A(n8405), .Z(n8345) );
  XOR U16474 ( .A(n8331), .B(n8406), .Z(n8343) );
  XOR U16475 ( .A(n8332), .B(n8333), .Z(n8406) );
  XOR U16476 ( .A(n8338), .B(n8407), .Z(n8333) );
  XOR U16477 ( .A(n8337), .B(n8340), .Z(n8407) );
  IV U16478 ( .A(n8339), .Z(n8340) );
  NAND U16479 ( .A(n8408), .B(n8409), .Z(n8339) );
  OR U16480 ( .A(n8410), .B(n8411), .Z(n8409) );
  OR U16481 ( .A(n8412), .B(n8413), .Z(n8408) );
  NAND U16482 ( .A(n8414), .B(n8415), .Z(n8337) );
  OR U16483 ( .A(n8416), .B(n8417), .Z(n8415) );
  OR U16484 ( .A(n8418), .B(n8419), .Z(n8414) );
  NOR U16485 ( .A(n8420), .B(n8421), .Z(n8338) );
  ANDN U16486 ( .B(n8422), .A(n8423), .Z(n8332) );
  IV U16487 ( .A(n8424), .Z(n8422) );
  XNOR U16488 ( .A(n8325), .B(n8425), .Z(n8331) );
  XNOR U16489 ( .A(n8324), .B(n8326), .Z(n8425) );
  NAND U16490 ( .A(n8426), .B(n8427), .Z(n8326) );
  OR U16491 ( .A(n8428), .B(n8429), .Z(n8427) );
  OR U16492 ( .A(n8430), .B(n8431), .Z(n8426) );
  NAND U16493 ( .A(n8432), .B(n8433), .Z(n8324) );
  OR U16494 ( .A(n8434), .B(n8435), .Z(n8433) );
  OR U16495 ( .A(n8436), .B(n8437), .Z(n8432) );
  ANDN U16496 ( .B(n8438), .A(n8439), .Z(n8325) );
  IV U16497 ( .A(n8440), .Z(n8438) );
  XNOR U16498 ( .A(n8405), .B(n8404), .Z(N64648) );
  XOR U16499 ( .A(n8424), .B(n8423), .Z(n8404) );
  XNOR U16500 ( .A(n8439), .B(n8440), .Z(n8423) );
  XNOR U16501 ( .A(n8434), .B(n8435), .Z(n8440) );
  XNOR U16502 ( .A(n8436), .B(n8437), .Z(n8435) );
  XNOR U16503 ( .A(y[7501]), .B(x[7501]), .Z(n8437) );
  XNOR U16504 ( .A(y[7502]), .B(x[7502]), .Z(n8436) );
  XNOR U16505 ( .A(y[7500]), .B(x[7500]), .Z(n8434) );
  XNOR U16506 ( .A(n8428), .B(n8429), .Z(n8439) );
  XNOR U16507 ( .A(y[7497]), .B(x[7497]), .Z(n8429) );
  XNOR U16508 ( .A(n8430), .B(n8431), .Z(n8428) );
  XNOR U16509 ( .A(y[7498]), .B(x[7498]), .Z(n8431) );
  XNOR U16510 ( .A(y[7499]), .B(x[7499]), .Z(n8430) );
  XNOR U16511 ( .A(n8421), .B(n8420), .Z(n8424) );
  XNOR U16512 ( .A(n8416), .B(n8417), .Z(n8420) );
  XNOR U16513 ( .A(y[7494]), .B(x[7494]), .Z(n8417) );
  XNOR U16514 ( .A(n8418), .B(n8419), .Z(n8416) );
  XNOR U16515 ( .A(y[7495]), .B(x[7495]), .Z(n8419) );
  XNOR U16516 ( .A(y[7496]), .B(x[7496]), .Z(n8418) );
  XNOR U16517 ( .A(n8410), .B(n8411), .Z(n8421) );
  XNOR U16518 ( .A(y[7491]), .B(x[7491]), .Z(n8411) );
  XNOR U16519 ( .A(n8412), .B(n8413), .Z(n8410) );
  XNOR U16520 ( .A(y[7492]), .B(x[7492]), .Z(n8413) );
  XNOR U16521 ( .A(y[7493]), .B(x[7493]), .Z(n8412) );
  XOR U16522 ( .A(n8386), .B(n8387), .Z(n8405) );
  XNOR U16523 ( .A(n8402), .B(n8403), .Z(n8387) );
  XNOR U16524 ( .A(n8397), .B(n8398), .Z(n8403) );
  XNOR U16525 ( .A(n8399), .B(n8400), .Z(n8398) );
  XNOR U16526 ( .A(y[7489]), .B(x[7489]), .Z(n8400) );
  XNOR U16527 ( .A(y[7490]), .B(x[7490]), .Z(n8399) );
  XNOR U16528 ( .A(y[7488]), .B(x[7488]), .Z(n8397) );
  XNOR U16529 ( .A(n8391), .B(n8392), .Z(n8402) );
  XNOR U16530 ( .A(y[7485]), .B(x[7485]), .Z(n8392) );
  XNOR U16531 ( .A(n8393), .B(n8394), .Z(n8391) );
  XNOR U16532 ( .A(y[7486]), .B(x[7486]), .Z(n8394) );
  XNOR U16533 ( .A(y[7487]), .B(x[7487]), .Z(n8393) );
  XOR U16534 ( .A(n8385), .B(n8384), .Z(n8386) );
  XNOR U16535 ( .A(n8380), .B(n8381), .Z(n8384) );
  XNOR U16536 ( .A(y[7482]), .B(x[7482]), .Z(n8381) );
  XNOR U16537 ( .A(n8382), .B(n8383), .Z(n8380) );
  XNOR U16538 ( .A(y[7483]), .B(x[7483]), .Z(n8383) );
  XNOR U16539 ( .A(y[7484]), .B(x[7484]), .Z(n8382) );
  XNOR U16540 ( .A(n8374), .B(n8375), .Z(n8385) );
  XNOR U16541 ( .A(y[7479]), .B(x[7479]), .Z(n8375) );
  XNOR U16542 ( .A(n8376), .B(n8377), .Z(n8374) );
  XNOR U16543 ( .A(y[7480]), .B(x[7480]), .Z(n8377) );
  XNOR U16544 ( .A(y[7481]), .B(x[7481]), .Z(n8376) );
  NAND U16545 ( .A(n8441), .B(n8442), .Z(N64639) );
  NANDN U16546 ( .A(n8443), .B(n8444), .Z(n8442) );
  OR U16547 ( .A(n8445), .B(n8446), .Z(n8444) );
  NAND U16548 ( .A(n8445), .B(n8446), .Z(n8441) );
  XOR U16549 ( .A(n8445), .B(n8447), .Z(N64638) );
  XNOR U16550 ( .A(n8443), .B(n8446), .Z(n8447) );
  AND U16551 ( .A(n8448), .B(n8449), .Z(n8446) );
  NANDN U16552 ( .A(n8450), .B(n8451), .Z(n8449) );
  NANDN U16553 ( .A(n8452), .B(n8453), .Z(n8451) );
  NANDN U16554 ( .A(n8453), .B(n8452), .Z(n8448) );
  NAND U16555 ( .A(n8454), .B(n8455), .Z(n8443) );
  NANDN U16556 ( .A(n8456), .B(n8457), .Z(n8455) );
  OR U16557 ( .A(n8458), .B(n8459), .Z(n8457) );
  NAND U16558 ( .A(n8459), .B(n8458), .Z(n8454) );
  AND U16559 ( .A(n8460), .B(n8461), .Z(n8445) );
  NANDN U16560 ( .A(n8462), .B(n8463), .Z(n8461) );
  NANDN U16561 ( .A(n8464), .B(n8465), .Z(n8463) );
  NANDN U16562 ( .A(n8465), .B(n8464), .Z(n8460) );
  XOR U16563 ( .A(n8459), .B(n8466), .Z(N64637) );
  XOR U16564 ( .A(n8456), .B(n8458), .Z(n8466) );
  XNOR U16565 ( .A(n8452), .B(n8467), .Z(n8458) );
  XNOR U16566 ( .A(n8450), .B(n8453), .Z(n8467) );
  NAND U16567 ( .A(n8468), .B(n8469), .Z(n8453) );
  NAND U16568 ( .A(n8470), .B(n8471), .Z(n8469) );
  OR U16569 ( .A(n8472), .B(n8473), .Z(n8470) );
  NANDN U16570 ( .A(n8474), .B(n8472), .Z(n8468) );
  IV U16571 ( .A(n8473), .Z(n8474) );
  NAND U16572 ( .A(n8475), .B(n8476), .Z(n8450) );
  NAND U16573 ( .A(n8477), .B(n8478), .Z(n8476) );
  NANDN U16574 ( .A(n8479), .B(n8480), .Z(n8477) );
  NANDN U16575 ( .A(n8480), .B(n8479), .Z(n8475) );
  AND U16576 ( .A(n8481), .B(n8482), .Z(n8452) );
  NAND U16577 ( .A(n8483), .B(n8484), .Z(n8482) );
  OR U16578 ( .A(n8485), .B(n8486), .Z(n8483) );
  NANDN U16579 ( .A(n8487), .B(n8485), .Z(n8481) );
  NAND U16580 ( .A(n8488), .B(n8489), .Z(n8456) );
  NANDN U16581 ( .A(n8490), .B(n8491), .Z(n8489) );
  OR U16582 ( .A(n8492), .B(n8493), .Z(n8491) );
  NANDN U16583 ( .A(n8494), .B(n8492), .Z(n8488) );
  IV U16584 ( .A(n8493), .Z(n8494) );
  XNOR U16585 ( .A(n8464), .B(n8495), .Z(n8459) );
  XNOR U16586 ( .A(n8462), .B(n8465), .Z(n8495) );
  NAND U16587 ( .A(n8496), .B(n8497), .Z(n8465) );
  NAND U16588 ( .A(n8498), .B(n8499), .Z(n8497) );
  OR U16589 ( .A(n8500), .B(n8501), .Z(n8498) );
  NANDN U16590 ( .A(n8502), .B(n8500), .Z(n8496) );
  IV U16591 ( .A(n8501), .Z(n8502) );
  NAND U16592 ( .A(n8503), .B(n8504), .Z(n8462) );
  NAND U16593 ( .A(n8505), .B(n8506), .Z(n8504) );
  NANDN U16594 ( .A(n8507), .B(n8508), .Z(n8505) );
  NANDN U16595 ( .A(n8508), .B(n8507), .Z(n8503) );
  AND U16596 ( .A(n8509), .B(n8510), .Z(n8464) );
  NAND U16597 ( .A(n8511), .B(n8512), .Z(n8510) );
  OR U16598 ( .A(n8513), .B(n8514), .Z(n8511) );
  NANDN U16599 ( .A(n8515), .B(n8513), .Z(n8509) );
  XNOR U16600 ( .A(n8490), .B(n8516), .Z(N64636) );
  XOR U16601 ( .A(n8492), .B(n8493), .Z(n8516) );
  XNOR U16602 ( .A(n8506), .B(n8517), .Z(n8493) );
  XOR U16603 ( .A(n8507), .B(n8508), .Z(n8517) );
  XOR U16604 ( .A(n8513), .B(n8518), .Z(n8508) );
  XOR U16605 ( .A(n8512), .B(n8515), .Z(n8518) );
  IV U16606 ( .A(n8514), .Z(n8515) );
  NAND U16607 ( .A(n8519), .B(n8520), .Z(n8514) );
  OR U16608 ( .A(n8521), .B(n8522), .Z(n8520) );
  OR U16609 ( .A(n8523), .B(n8524), .Z(n8519) );
  NAND U16610 ( .A(n8525), .B(n8526), .Z(n8512) );
  OR U16611 ( .A(n8527), .B(n8528), .Z(n8526) );
  OR U16612 ( .A(n8529), .B(n8530), .Z(n8525) );
  NOR U16613 ( .A(n8531), .B(n8532), .Z(n8513) );
  ANDN U16614 ( .B(n8533), .A(n8534), .Z(n8507) );
  XNOR U16615 ( .A(n8500), .B(n8535), .Z(n8506) );
  XNOR U16616 ( .A(n8499), .B(n8501), .Z(n8535) );
  NAND U16617 ( .A(n8536), .B(n8537), .Z(n8501) );
  OR U16618 ( .A(n8538), .B(n8539), .Z(n8537) );
  OR U16619 ( .A(n8540), .B(n8541), .Z(n8536) );
  NAND U16620 ( .A(n8542), .B(n8543), .Z(n8499) );
  OR U16621 ( .A(n8544), .B(n8545), .Z(n8543) );
  OR U16622 ( .A(n8546), .B(n8547), .Z(n8542) );
  ANDN U16623 ( .B(n8548), .A(n8549), .Z(n8500) );
  IV U16624 ( .A(n8550), .Z(n8548) );
  ANDN U16625 ( .B(n8551), .A(n8552), .Z(n8492) );
  XOR U16626 ( .A(n8478), .B(n8553), .Z(n8490) );
  XOR U16627 ( .A(n8479), .B(n8480), .Z(n8553) );
  XOR U16628 ( .A(n8485), .B(n8554), .Z(n8480) );
  XOR U16629 ( .A(n8484), .B(n8487), .Z(n8554) );
  IV U16630 ( .A(n8486), .Z(n8487) );
  NAND U16631 ( .A(n8555), .B(n8556), .Z(n8486) );
  OR U16632 ( .A(n8557), .B(n8558), .Z(n8556) );
  OR U16633 ( .A(n8559), .B(n8560), .Z(n8555) );
  NAND U16634 ( .A(n8561), .B(n8562), .Z(n8484) );
  OR U16635 ( .A(n8563), .B(n8564), .Z(n8562) );
  OR U16636 ( .A(n8565), .B(n8566), .Z(n8561) );
  NOR U16637 ( .A(n8567), .B(n8568), .Z(n8485) );
  ANDN U16638 ( .B(n8569), .A(n8570), .Z(n8479) );
  IV U16639 ( .A(n8571), .Z(n8569) );
  XNOR U16640 ( .A(n8472), .B(n8572), .Z(n8478) );
  XNOR U16641 ( .A(n8471), .B(n8473), .Z(n8572) );
  NAND U16642 ( .A(n8573), .B(n8574), .Z(n8473) );
  OR U16643 ( .A(n8575), .B(n8576), .Z(n8574) );
  OR U16644 ( .A(n8577), .B(n8578), .Z(n8573) );
  NAND U16645 ( .A(n8579), .B(n8580), .Z(n8471) );
  OR U16646 ( .A(n8581), .B(n8582), .Z(n8580) );
  OR U16647 ( .A(n8583), .B(n8584), .Z(n8579) );
  ANDN U16648 ( .B(n8585), .A(n8586), .Z(n8472) );
  IV U16649 ( .A(n8587), .Z(n8585) );
  XNOR U16650 ( .A(n8552), .B(n8551), .Z(N64635) );
  XOR U16651 ( .A(n8571), .B(n8570), .Z(n8551) );
  XNOR U16652 ( .A(n8586), .B(n8587), .Z(n8570) );
  XNOR U16653 ( .A(n8581), .B(n8582), .Z(n8587) );
  XNOR U16654 ( .A(n8583), .B(n8584), .Z(n8582) );
  XNOR U16655 ( .A(y[7477]), .B(x[7477]), .Z(n8584) );
  XNOR U16656 ( .A(y[7478]), .B(x[7478]), .Z(n8583) );
  XNOR U16657 ( .A(y[7476]), .B(x[7476]), .Z(n8581) );
  XNOR U16658 ( .A(n8575), .B(n8576), .Z(n8586) );
  XNOR U16659 ( .A(y[7473]), .B(x[7473]), .Z(n8576) );
  XNOR U16660 ( .A(n8577), .B(n8578), .Z(n8575) );
  XNOR U16661 ( .A(y[7474]), .B(x[7474]), .Z(n8578) );
  XNOR U16662 ( .A(y[7475]), .B(x[7475]), .Z(n8577) );
  XNOR U16663 ( .A(n8568), .B(n8567), .Z(n8571) );
  XNOR U16664 ( .A(n8563), .B(n8564), .Z(n8567) );
  XNOR U16665 ( .A(y[7470]), .B(x[7470]), .Z(n8564) );
  XNOR U16666 ( .A(n8565), .B(n8566), .Z(n8563) );
  XNOR U16667 ( .A(y[7471]), .B(x[7471]), .Z(n8566) );
  XNOR U16668 ( .A(y[7472]), .B(x[7472]), .Z(n8565) );
  XNOR U16669 ( .A(n8557), .B(n8558), .Z(n8568) );
  XNOR U16670 ( .A(y[7467]), .B(x[7467]), .Z(n8558) );
  XNOR U16671 ( .A(n8559), .B(n8560), .Z(n8557) );
  XNOR U16672 ( .A(y[7468]), .B(x[7468]), .Z(n8560) );
  XNOR U16673 ( .A(y[7469]), .B(x[7469]), .Z(n8559) );
  XOR U16674 ( .A(n8533), .B(n8534), .Z(n8552) );
  XNOR U16675 ( .A(n8549), .B(n8550), .Z(n8534) );
  XNOR U16676 ( .A(n8544), .B(n8545), .Z(n8550) );
  XNOR U16677 ( .A(n8546), .B(n8547), .Z(n8545) );
  XNOR U16678 ( .A(y[7465]), .B(x[7465]), .Z(n8547) );
  XNOR U16679 ( .A(y[7466]), .B(x[7466]), .Z(n8546) );
  XNOR U16680 ( .A(y[7464]), .B(x[7464]), .Z(n8544) );
  XNOR U16681 ( .A(n8538), .B(n8539), .Z(n8549) );
  XNOR U16682 ( .A(y[7461]), .B(x[7461]), .Z(n8539) );
  XNOR U16683 ( .A(n8540), .B(n8541), .Z(n8538) );
  XNOR U16684 ( .A(y[7462]), .B(x[7462]), .Z(n8541) );
  XNOR U16685 ( .A(y[7463]), .B(x[7463]), .Z(n8540) );
  XOR U16686 ( .A(n8532), .B(n8531), .Z(n8533) );
  XNOR U16687 ( .A(n8527), .B(n8528), .Z(n8531) );
  XNOR U16688 ( .A(y[7458]), .B(x[7458]), .Z(n8528) );
  XNOR U16689 ( .A(n8529), .B(n8530), .Z(n8527) );
  XNOR U16690 ( .A(y[7459]), .B(x[7459]), .Z(n8530) );
  XNOR U16691 ( .A(y[7460]), .B(x[7460]), .Z(n8529) );
  XNOR U16692 ( .A(n8521), .B(n8522), .Z(n8532) );
  XNOR U16693 ( .A(y[7455]), .B(x[7455]), .Z(n8522) );
  XNOR U16694 ( .A(n8523), .B(n8524), .Z(n8521) );
  XNOR U16695 ( .A(y[7456]), .B(x[7456]), .Z(n8524) );
  XNOR U16696 ( .A(y[7457]), .B(x[7457]), .Z(n8523) );
  NAND U16697 ( .A(n8588), .B(n8589), .Z(N64626) );
  NANDN U16698 ( .A(n8590), .B(n8591), .Z(n8589) );
  OR U16699 ( .A(n8592), .B(n8593), .Z(n8591) );
  NAND U16700 ( .A(n8592), .B(n8593), .Z(n8588) );
  XOR U16701 ( .A(n8592), .B(n8594), .Z(N64625) );
  XNOR U16702 ( .A(n8590), .B(n8593), .Z(n8594) );
  AND U16703 ( .A(n8595), .B(n8596), .Z(n8593) );
  NANDN U16704 ( .A(n8597), .B(n8598), .Z(n8596) );
  NANDN U16705 ( .A(n8599), .B(n8600), .Z(n8598) );
  NANDN U16706 ( .A(n8600), .B(n8599), .Z(n8595) );
  NAND U16707 ( .A(n8601), .B(n8602), .Z(n8590) );
  NANDN U16708 ( .A(n8603), .B(n8604), .Z(n8602) );
  OR U16709 ( .A(n8605), .B(n8606), .Z(n8604) );
  NAND U16710 ( .A(n8606), .B(n8605), .Z(n8601) );
  AND U16711 ( .A(n8607), .B(n8608), .Z(n8592) );
  NANDN U16712 ( .A(n8609), .B(n8610), .Z(n8608) );
  NANDN U16713 ( .A(n8611), .B(n8612), .Z(n8610) );
  NANDN U16714 ( .A(n8612), .B(n8611), .Z(n8607) );
  XOR U16715 ( .A(n8606), .B(n8613), .Z(N64624) );
  XOR U16716 ( .A(n8603), .B(n8605), .Z(n8613) );
  XNOR U16717 ( .A(n8599), .B(n8614), .Z(n8605) );
  XNOR U16718 ( .A(n8597), .B(n8600), .Z(n8614) );
  NAND U16719 ( .A(n8615), .B(n8616), .Z(n8600) );
  NAND U16720 ( .A(n8617), .B(n8618), .Z(n8616) );
  OR U16721 ( .A(n8619), .B(n8620), .Z(n8617) );
  NANDN U16722 ( .A(n8621), .B(n8619), .Z(n8615) );
  IV U16723 ( .A(n8620), .Z(n8621) );
  NAND U16724 ( .A(n8622), .B(n8623), .Z(n8597) );
  NAND U16725 ( .A(n8624), .B(n8625), .Z(n8623) );
  NANDN U16726 ( .A(n8626), .B(n8627), .Z(n8624) );
  NANDN U16727 ( .A(n8627), .B(n8626), .Z(n8622) );
  AND U16728 ( .A(n8628), .B(n8629), .Z(n8599) );
  NAND U16729 ( .A(n8630), .B(n8631), .Z(n8629) );
  OR U16730 ( .A(n8632), .B(n8633), .Z(n8630) );
  NANDN U16731 ( .A(n8634), .B(n8632), .Z(n8628) );
  NAND U16732 ( .A(n8635), .B(n8636), .Z(n8603) );
  NANDN U16733 ( .A(n8637), .B(n8638), .Z(n8636) );
  OR U16734 ( .A(n8639), .B(n8640), .Z(n8638) );
  NANDN U16735 ( .A(n8641), .B(n8639), .Z(n8635) );
  IV U16736 ( .A(n8640), .Z(n8641) );
  XNOR U16737 ( .A(n8611), .B(n8642), .Z(n8606) );
  XNOR U16738 ( .A(n8609), .B(n8612), .Z(n8642) );
  NAND U16739 ( .A(n8643), .B(n8644), .Z(n8612) );
  NAND U16740 ( .A(n8645), .B(n8646), .Z(n8644) );
  OR U16741 ( .A(n8647), .B(n8648), .Z(n8645) );
  NANDN U16742 ( .A(n8649), .B(n8647), .Z(n8643) );
  IV U16743 ( .A(n8648), .Z(n8649) );
  NAND U16744 ( .A(n8650), .B(n8651), .Z(n8609) );
  NAND U16745 ( .A(n8652), .B(n8653), .Z(n8651) );
  NANDN U16746 ( .A(n8654), .B(n8655), .Z(n8652) );
  NANDN U16747 ( .A(n8655), .B(n8654), .Z(n8650) );
  AND U16748 ( .A(n8656), .B(n8657), .Z(n8611) );
  NAND U16749 ( .A(n8658), .B(n8659), .Z(n8657) );
  OR U16750 ( .A(n8660), .B(n8661), .Z(n8658) );
  NANDN U16751 ( .A(n8662), .B(n8660), .Z(n8656) );
  XNOR U16752 ( .A(n8637), .B(n8663), .Z(N64623) );
  XOR U16753 ( .A(n8639), .B(n8640), .Z(n8663) );
  XNOR U16754 ( .A(n8653), .B(n8664), .Z(n8640) );
  XOR U16755 ( .A(n8654), .B(n8655), .Z(n8664) );
  XOR U16756 ( .A(n8660), .B(n8665), .Z(n8655) );
  XOR U16757 ( .A(n8659), .B(n8662), .Z(n8665) );
  IV U16758 ( .A(n8661), .Z(n8662) );
  NAND U16759 ( .A(n8666), .B(n8667), .Z(n8661) );
  OR U16760 ( .A(n8668), .B(n8669), .Z(n8667) );
  OR U16761 ( .A(n8670), .B(n8671), .Z(n8666) );
  NAND U16762 ( .A(n8672), .B(n8673), .Z(n8659) );
  OR U16763 ( .A(n8674), .B(n8675), .Z(n8673) );
  OR U16764 ( .A(n8676), .B(n8677), .Z(n8672) );
  NOR U16765 ( .A(n8678), .B(n8679), .Z(n8660) );
  ANDN U16766 ( .B(n8680), .A(n8681), .Z(n8654) );
  XNOR U16767 ( .A(n8647), .B(n8682), .Z(n8653) );
  XNOR U16768 ( .A(n8646), .B(n8648), .Z(n8682) );
  NAND U16769 ( .A(n8683), .B(n8684), .Z(n8648) );
  OR U16770 ( .A(n8685), .B(n8686), .Z(n8684) );
  OR U16771 ( .A(n8687), .B(n8688), .Z(n8683) );
  NAND U16772 ( .A(n8689), .B(n8690), .Z(n8646) );
  OR U16773 ( .A(n8691), .B(n8692), .Z(n8690) );
  OR U16774 ( .A(n8693), .B(n8694), .Z(n8689) );
  ANDN U16775 ( .B(n8695), .A(n8696), .Z(n8647) );
  IV U16776 ( .A(n8697), .Z(n8695) );
  ANDN U16777 ( .B(n8698), .A(n8699), .Z(n8639) );
  XOR U16778 ( .A(n8625), .B(n8700), .Z(n8637) );
  XOR U16779 ( .A(n8626), .B(n8627), .Z(n8700) );
  XOR U16780 ( .A(n8632), .B(n8701), .Z(n8627) );
  XOR U16781 ( .A(n8631), .B(n8634), .Z(n8701) );
  IV U16782 ( .A(n8633), .Z(n8634) );
  NAND U16783 ( .A(n8702), .B(n8703), .Z(n8633) );
  OR U16784 ( .A(n8704), .B(n8705), .Z(n8703) );
  OR U16785 ( .A(n8706), .B(n8707), .Z(n8702) );
  NAND U16786 ( .A(n8708), .B(n8709), .Z(n8631) );
  OR U16787 ( .A(n8710), .B(n8711), .Z(n8709) );
  OR U16788 ( .A(n8712), .B(n8713), .Z(n8708) );
  NOR U16789 ( .A(n8714), .B(n8715), .Z(n8632) );
  ANDN U16790 ( .B(n8716), .A(n8717), .Z(n8626) );
  IV U16791 ( .A(n8718), .Z(n8716) );
  XNOR U16792 ( .A(n8619), .B(n8719), .Z(n8625) );
  XNOR U16793 ( .A(n8618), .B(n8620), .Z(n8719) );
  NAND U16794 ( .A(n8720), .B(n8721), .Z(n8620) );
  OR U16795 ( .A(n8722), .B(n8723), .Z(n8721) );
  OR U16796 ( .A(n8724), .B(n8725), .Z(n8720) );
  NAND U16797 ( .A(n8726), .B(n8727), .Z(n8618) );
  OR U16798 ( .A(n8728), .B(n8729), .Z(n8727) );
  OR U16799 ( .A(n8730), .B(n8731), .Z(n8726) );
  ANDN U16800 ( .B(n8732), .A(n8733), .Z(n8619) );
  IV U16801 ( .A(n8734), .Z(n8732) );
  XNOR U16802 ( .A(n8699), .B(n8698), .Z(N64622) );
  XOR U16803 ( .A(n8718), .B(n8717), .Z(n8698) );
  XNOR U16804 ( .A(n8733), .B(n8734), .Z(n8717) );
  XNOR U16805 ( .A(n8728), .B(n8729), .Z(n8734) );
  XNOR U16806 ( .A(n8730), .B(n8731), .Z(n8729) );
  XNOR U16807 ( .A(y[7453]), .B(x[7453]), .Z(n8731) );
  XNOR U16808 ( .A(y[7454]), .B(x[7454]), .Z(n8730) );
  XNOR U16809 ( .A(y[7452]), .B(x[7452]), .Z(n8728) );
  XNOR U16810 ( .A(n8722), .B(n8723), .Z(n8733) );
  XNOR U16811 ( .A(y[7449]), .B(x[7449]), .Z(n8723) );
  XNOR U16812 ( .A(n8724), .B(n8725), .Z(n8722) );
  XNOR U16813 ( .A(y[7450]), .B(x[7450]), .Z(n8725) );
  XNOR U16814 ( .A(y[7451]), .B(x[7451]), .Z(n8724) );
  XNOR U16815 ( .A(n8715), .B(n8714), .Z(n8718) );
  XNOR U16816 ( .A(n8710), .B(n8711), .Z(n8714) );
  XNOR U16817 ( .A(y[7446]), .B(x[7446]), .Z(n8711) );
  XNOR U16818 ( .A(n8712), .B(n8713), .Z(n8710) );
  XNOR U16819 ( .A(y[7447]), .B(x[7447]), .Z(n8713) );
  XNOR U16820 ( .A(y[7448]), .B(x[7448]), .Z(n8712) );
  XNOR U16821 ( .A(n8704), .B(n8705), .Z(n8715) );
  XNOR U16822 ( .A(y[7443]), .B(x[7443]), .Z(n8705) );
  XNOR U16823 ( .A(n8706), .B(n8707), .Z(n8704) );
  XNOR U16824 ( .A(y[7444]), .B(x[7444]), .Z(n8707) );
  XNOR U16825 ( .A(y[7445]), .B(x[7445]), .Z(n8706) );
  XOR U16826 ( .A(n8680), .B(n8681), .Z(n8699) );
  XNOR U16827 ( .A(n8696), .B(n8697), .Z(n8681) );
  XNOR U16828 ( .A(n8691), .B(n8692), .Z(n8697) );
  XNOR U16829 ( .A(n8693), .B(n8694), .Z(n8692) );
  XNOR U16830 ( .A(y[7441]), .B(x[7441]), .Z(n8694) );
  XNOR U16831 ( .A(y[7442]), .B(x[7442]), .Z(n8693) );
  XNOR U16832 ( .A(y[7440]), .B(x[7440]), .Z(n8691) );
  XNOR U16833 ( .A(n8685), .B(n8686), .Z(n8696) );
  XNOR U16834 ( .A(y[7437]), .B(x[7437]), .Z(n8686) );
  XNOR U16835 ( .A(n8687), .B(n8688), .Z(n8685) );
  XNOR U16836 ( .A(y[7438]), .B(x[7438]), .Z(n8688) );
  XNOR U16837 ( .A(y[7439]), .B(x[7439]), .Z(n8687) );
  XOR U16838 ( .A(n8679), .B(n8678), .Z(n8680) );
  XNOR U16839 ( .A(n8674), .B(n8675), .Z(n8678) );
  XNOR U16840 ( .A(y[7434]), .B(x[7434]), .Z(n8675) );
  XNOR U16841 ( .A(n8676), .B(n8677), .Z(n8674) );
  XNOR U16842 ( .A(y[7435]), .B(x[7435]), .Z(n8677) );
  XNOR U16843 ( .A(y[7436]), .B(x[7436]), .Z(n8676) );
  XNOR U16844 ( .A(n8668), .B(n8669), .Z(n8679) );
  XNOR U16845 ( .A(y[7431]), .B(x[7431]), .Z(n8669) );
  XNOR U16846 ( .A(n8670), .B(n8671), .Z(n8668) );
  XNOR U16847 ( .A(y[7432]), .B(x[7432]), .Z(n8671) );
  XNOR U16848 ( .A(y[7433]), .B(x[7433]), .Z(n8670) );
  NAND U16849 ( .A(n8735), .B(n8736), .Z(N64613) );
  NANDN U16850 ( .A(n8737), .B(n8738), .Z(n8736) );
  OR U16851 ( .A(n8739), .B(n8740), .Z(n8738) );
  NAND U16852 ( .A(n8739), .B(n8740), .Z(n8735) );
  XOR U16853 ( .A(n8739), .B(n8741), .Z(N64612) );
  XNOR U16854 ( .A(n8737), .B(n8740), .Z(n8741) );
  AND U16855 ( .A(n8742), .B(n8743), .Z(n8740) );
  NANDN U16856 ( .A(n8744), .B(n8745), .Z(n8743) );
  NANDN U16857 ( .A(n8746), .B(n8747), .Z(n8745) );
  NANDN U16858 ( .A(n8747), .B(n8746), .Z(n8742) );
  NAND U16859 ( .A(n8748), .B(n8749), .Z(n8737) );
  NANDN U16860 ( .A(n8750), .B(n8751), .Z(n8749) );
  OR U16861 ( .A(n8752), .B(n8753), .Z(n8751) );
  NAND U16862 ( .A(n8753), .B(n8752), .Z(n8748) );
  AND U16863 ( .A(n8754), .B(n8755), .Z(n8739) );
  NANDN U16864 ( .A(n8756), .B(n8757), .Z(n8755) );
  NANDN U16865 ( .A(n8758), .B(n8759), .Z(n8757) );
  NANDN U16866 ( .A(n8759), .B(n8758), .Z(n8754) );
  XOR U16867 ( .A(n8753), .B(n8760), .Z(N64611) );
  XOR U16868 ( .A(n8750), .B(n8752), .Z(n8760) );
  XNOR U16869 ( .A(n8746), .B(n8761), .Z(n8752) );
  XNOR U16870 ( .A(n8744), .B(n8747), .Z(n8761) );
  NAND U16871 ( .A(n8762), .B(n8763), .Z(n8747) );
  NAND U16872 ( .A(n8764), .B(n8765), .Z(n8763) );
  OR U16873 ( .A(n8766), .B(n8767), .Z(n8764) );
  NANDN U16874 ( .A(n8768), .B(n8766), .Z(n8762) );
  IV U16875 ( .A(n8767), .Z(n8768) );
  NAND U16876 ( .A(n8769), .B(n8770), .Z(n8744) );
  NAND U16877 ( .A(n8771), .B(n8772), .Z(n8770) );
  NANDN U16878 ( .A(n8773), .B(n8774), .Z(n8771) );
  NANDN U16879 ( .A(n8774), .B(n8773), .Z(n8769) );
  AND U16880 ( .A(n8775), .B(n8776), .Z(n8746) );
  NAND U16881 ( .A(n8777), .B(n8778), .Z(n8776) );
  OR U16882 ( .A(n8779), .B(n8780), .Z(n8777) );
  NANDN U16883 ( .A(n8781), .B(n8779), .Z(n8775) );
  NAND U16884 ( .A(n8782), .B(n8783), .Z(n8750) );
  NANDN U16885 ( .A(n8784), .B(n8785), .Z(n8783) );
  OR U16886 ( .A(n8786), .B(n8787), .Z(n8785) );
  NANDN U16887 ( .A(n8788), .B(n8786), .Z(n8782) );
  IV U16888 ( .A(n8787), .Z(n8788) );
  XNOR U16889 ( .A(n8758), .B(n8789), .Z(n8753) );
  XNOR U16890 ( .A(n8756), .B(n8759), .Z(n8789) );
  NAND U16891 ( .A(n8790), .B(n8791), .Z(n8759) );
  NAND U16892 ( .A(n8792), .B(n8793), .Z(n8791) );
  OR U16893 ( .A(n8794), .B(n8795), .Z(n8792) );
  NANDN U16894 ( .A(n8796), .B(n8794), .Z(n8790) );
  IV U16895 ( .A(n8795), .Z(n8796) );
  NAND U16896 ( .A(n8797), .B(n8798), .Z(n8756) );
  NAND U16897 ( .A(n8799), .B(n8800), .Z(n8798) );
  NANDN U16898 ( .A(n8801), .B(n8802), .Z(n8799) );
  NANDN U16899 ( .A(n8802), .B(n8801), .Z(n8797) );
  AND U16900 ( .A(n8803), .B(n8804), .Z(n8758) );
  NAND U16901 ( .A(n8805), .B(n8806), .Z(n8804) );
  OR U16902 ( .A(n8807), .B(n8808), .Z(n8805) );
  NANDN U16903 ( .A(n8809), .B(n8807), .Z(n8803) );
  XNOR U16904 ( .A(n8784), .B(n8810), .Z(N64610) );
  XOR U16905 ( .A(n8786), .B(n8787), .Z(n8810) );
  XNOR U16906 ( .A(n8800), .B(n8811), .Z(n8787) );
  XOR U16907 ( .A(n8801), .B(n8802), .Z(n8811) );
  XOR U16908 ( .A(n8807), .B(n8812), .Z(n8802) );
  XOR U16909 ( .A(n8806), .B(n8809), .Z(n8812) );
  IV U16910 ( .A(n8808), .Z(n8809) );
  NAND U16911 ( .A(n8813), .B(n8814), .Z(n8808) );
  OR U16912 ( .A(n8815), .B(n8816), .Z(n8814) );
  OR U16913 ( .A(n8817), .B(n8818), .Z(n8813) );
  NAND U16914 ( .A(n8819), .B(n8820), .Z(n8806) );
  OR U16915 ( .A(n8821), .B(n8822), .Z(n8820) );
  OR U16916 ( .A(n8823), .B(n8824), .Z(n8819) );
  NOR U16917 ( .A(n8825), .B(n8826), .Z(n8807) );
  ANDN U16918 ( .B(n8827), .A(n8828), .Z(n8801) );
  XNOR U16919 ( .A(n8794), .B(n8829), .Z(n8800) );
  XNOR U16920 ( .A(n8793), .B(n8795), .Z(n8829) );
  NAND U16921 ( .A(n8830), .B(n8831), .Z(n8795) );
  OR U16922 ( .A(n8832), .B(n8833), .Z(n8831) );
  OR U16923 ( .A(n8834), .B(n8835), .Z(n8830) );
  NAND U16924 ( .A(n8836), .B(n8837), .Z(n8793) );
  OR U16925 ( .A(n8838), .B(n8839), .Z(n8837) );
  OR U16926 ( .A(n8840), .B(n8841), .Z(n8836) );
  ANDN U16927 ( .B(n8842), .A(n8843), .Z(n8794) );
  IV U16928 ( .A(n8844), .Z(n8842) );
  ANDN U16929 ( .B(n8845), .A(n8846), .Z(n8786) );
  XOR U16930 ( .A(n8772), .B(n8847), .Z(n8784) );
  XOR U16931 ( .A(n8773), .B(n8774), .Z(n8847) );
  XOR U16932 ( .A(n8779), .B(n8848), .Z(n8774) );
  XOR U16933 ( .A(n8778), .B(n8781), .Z(n8848) );
  IV U16934 ( .A(n8780), .Z(n8781) );
  NAND U16935 ( .A(n8849), .B(n8850), .Z(n8780) );
  OR U16936 ( .A(n8851), .B(n8852), .Z(n8850) );
  OR U16937 ( .A(n8853), .B(n8854), .Z(n8849) );
  NAND U16938 ( .A(n8855), .B(n8856), .Z(n8778) );
  OR U16939 ( .A(n8857), .B(n8858), .Z(n8856) );
  OR U16940 ( .A(n8859), .B(n8860), .Z(n8855) );
  NOR U16941 ( .A(n8861), .B(n8862), .Z(n8779) );
  ANDN U16942 ( .B(n8863), .A(n8864), .Z(n8773) );
  IV U16943 ( .A(n8865), .Z(n8863) );
  XNOR U16944 ( .A(n8766), .B(n8866), .Z(n8772) );
  XNOR U16945 ( .A(n8765), .B(n8767), .Z(n8866) );
  NAND U16946 ( .A(n8867), .B(n8868), .Z(n8767) );
  OR U16947 ( .A(n8869), .B(n8870), .Z(n8868) );
  OR U16948 ( .A(n8871), .B(n8872), .Z(n8867) );
  NAND U16949 ( .A(n8873), .B(n8874), .Z(n8765) );
  OR U16950 ( .A(n8875), .B(n8876), .Z(n8874) );
  OR U16951 ( .A(n8877), .B(n8878), .Z(n8873) );
  ANDN U16952 ( .B(n8879), .A(n8880), .Z(n8766) );
  IV U16953 ( .A(n8881), .Z(n8879) );
  XNOR U16954 ( .A(n8846), .B(n8845), .Z(N64609) );
  XOR U16955 ( .A(n8865), .B(n8864), .Z(n8845) );
  XNOR U16956 ( .A(n8880), .B(n8881), .Z(n8864) );
  XNOR U16957 ( .A(n8875), .B(n8876), .Z(n8881) );
  XNOR U16958 ( .A(n8877), .B(n8878), .Z(n8876) );
  XNOR U16959 ( .A(y[7429]), .B(x[7429]), .Z(n8878) );
  XNOR U16960 ( .A(y[7430]), .B(x[7430]), .Z(n8877) );
  XNOR U16961 ( .A(y[7428]), .B(x[7428]), .Z(n8875) );
  XNOR U16962 ( .A(n8869), .B(n8870), .Z(n8880) );
  XNOR U16963 ( .A(y[7425]), .B(x[7425]), .Z(n8870) );
  XNOR U16964 ( .A(n8871), .B(n8872), .Z(n8869) );
  XNOR U16965 ( .A(y[7426]), .B(x[7426]), .Z(n8872) );
  XNOR U16966 ( .A(y[7427]), .B(x[7427]), .Z(n8871) );
  XNOR U16967 ( .A(n8862), .B(n8861), .Z(n8865) );
  XNOR U16968 ( .A(n8857), .B(n8858), .Z(n8861) );
  XNOR U16969 ( .A(y[7422]), .B(x[7422]), .Z(n8858) );
  XNOR U16970 ( .A(n8859), .B(n8860), .Z(n8857) );
  XNOR U16971 ( .A(y[7423]), .B(x[7423]), .Z(n8860) );
  XNOR U16972 ( .A(y[7424]), .B(x[7424]), .Z(n8859) );
  XNOR U16973 ( .A(n8851), .B(n8852), .Z(n8862) );
  XNOR U16974 ( .A(y[7419]), .B(x[7419]), .Z(n8852) );
  XNOR U16975 ( .A(n8853), .B(n8854), .Z(n8851) );
  XNOR U16976 ( .A(y[7420]), .B(x[7420]), .Z(n8854) );
  XNOR U16977 ( .A(y[7421]), .B(x[7421]), .Z(n8853) );
  XOR U16978 ( .A(n8827), .B(n8828), .Z(n8846) );
  XNOR U16979 ( .A(n8843), .B(n8844), .Z(n8828) );
  XNOR U16980 ( .A(n8838), .B(n8839), .Z(n8844) );
  XNOR U16981 ( .A(n8840), .B(n8841), .Z(n8839) );
  XNOR U16982 ( .A(y[7417]), .B(x[7417]), .Z(n8841) );
  XNOR U16983 ( .A(y[7418]), .B(x[7418]), .Z(n8840) );
  XNOR U16984 ( .A(y[7416]), .B(x[7416]), .Z(n8838) );
  XNOR U16985 ( .A(n8832), .B(n8833), .Z(n8843) );
  XNOR U16986 ( .A(y[7413]), .B(x[7413]), .Z(n8833) );
  XNOR U16987 ( .A(n8834), .B(n8835), .Z(n8832) );
  XNOR U16988 ( .A(y[7414]), .B(x[7414]), .Z(n8835) );
  XNOR U16989 ( .A(y[7415]), .B(x[7415]), .Z(n8834) );
  XOR U16990 ( .A(n8826), .B(n8825), .Z(n8827) );
  XNOR U16991 ( .A(n8821), .B(n8822), .Z(n8825) );
  XNOR U16992 ( .A(y[7410]), .B(x[7410]), .Z(n8822) );
  XNOR U16993 ( .A(n8823), .B(n8824), .Z(n8821) );
  XNOR U16994 ( .A(y[7411]), .B(x[7411]), .Z(n8824) );
  XNOR U16995 ( .A(y[7412]), .B(x[7412]), .Z(n8823) );
  XNOR U16996 ( .A(n8815), .B(n8816), .Z(n8826) );
  XNOR U16997 ( .A(y[7407]), .B(x[7407]), .Z(n8816) );
  XNOR U16998 ( .A(n8817), .B(n8818), .Z(n8815) );
  XNOR U16999 ( .A(y[7408]), .B(x[7408]), .Z(n8818) );
  XNOR U17000 ( .A(y[7409]), .B(x[7409]), .Z(n8817) );
  NAND U17001 ( .A(n8882), .B(n8883), .Z(N64600) );
  NANDN U17002 ( .A(n8884), .B(n8885), .Z(n8883) );
  OR U17003 ( .A(n8886), .B(n8887), .Z(n8885) );
  NAND U17004 ( .A(n8886), .B(n8887), .Z(n8882) );
  XOR U17005 ( .A(n8886), .B(n8888), .Z(N64599) );
  XNOR U17006 ( .A(n8884), .B(n8887), .Z(n8888) );
  AND U17007 ( .A(n8889), .B(n8890), .Z(n8887) );
  NANDN U17008 ( .A(n8891), .B(n8892), .Z(n8890) );
  NANDN U17009 ( .A(n8893), .B(n8894), .Z(n8892) );
  NANDN U17010 ( .A(n8894), .B(n8893), .Z(n8889) );
  NAND U17011 ( .A(n8895), .B(n8896), .Z(n8884) );
  NANDN U17012 ( .A(n8897), .B(n8898), .Z(n8896) );
  OR U17013 ( .A(n8899), .B(n8900), .Z(n8898) );
  NAND U17014 ( .A(n8900), .B(n8899), .Z(n8895) );
  AND U17015 ( .A(n8901), .B(n8902), .Z(n8886) );
  NANDN U17016 ( .A(n8903), .B(n8904), .Z(n8902) );
  NANDN U17017 ( .A(n8905), .B(n8906), .Z(n8904) );
  NANDN U17018 ( .A(n8906), .B(n8905), .Z(n8901) );
  XOR U17019 ( .A(n8900), .B(n8907), .Z(N64598) );
  XOR U17020 ( .A(n8897), .B(n8899), .Z(n8907) );
  XNOR U17021 ( .A(n8893), .B(n8908), .Z(n8899) );
  XNOR U17022 ( .A(n8891), .B(n8894), .Z(n8908) );
  NAND U17023 ( .A(n8909), .B(n8910), .Z(n8894) );
  NAND U17024 ( .A(n8911), .B(n8912), .Z(n8910) );
  OR U17025 ( .A(n8913), .B(n8914), .Z(n8911) );
  NANDN U17026 ( .A(n8915), .B(n8913), .Z(n8909) );
  IV U17027 ( .A(n8914), .Z(n8915) );
  NAND U17028 ( .A(n8916), .B(n8917), .Z(n8891) );
  NAND U17029 ( .A(n8918), .B(n8919), .Z(n8917) );
  NANDN U17030 ( .A(n8920), .B(n8921), .Z(n8918) );
  NANDN U17031 ( .A(n8921), .B(n8920), .Z(n8916) );
  AND U17032 ( .A(n8922), .B(n8923), .Z(n8893) );
  NAND U17033 ( .A(n8924), .B(n8925), .Z(n8923) );
  OR U17034 ( .A(n8926), .B(n8927), .Z(n8924) );
  NANDN U17035 ( .A(n8928), .B(n8926), .Z(n8922) );
  NAND U17036 ( .A(n8929), .B(n8930), .Z(n8897) );
  NANDN U17037 ( .A(n8931), .B(n8932), .Z(n8930) );
  OR U17038 ( .A(n8933), .B(n8934), .Z(n8932) );
  NANDN U17039 ( .A(n8935), .B(n8933), .Z(n8929) );
  IV U17040 ( .A(n8934), .Z(n8935) );
  XNOR U17041 ( .A(n8905), .B(n8936), .Z(n8900) );
  XNOR U17042 ( .A(n8903), .B(n8906), .Z(n8936) );
  NAND U17043 ( .A(n8937), .B(n8938), .Z(n8906) );
  NAND U17044 ( .A(n8939), .B(n8940), .Z(n8938) );
  OR U17045 ( .A(n8941), .B(n8942), .Z(n8939) );
  NANDN U17046 ( .A(n8943), .B(n8941), .Z(n8937) );
  IV U17047 ( .A(n8942), .Z(n8943) );
  NAND U17048 ( .A(n8944), .B(n8945), .Z(n8903) );
  NAND U17049 ( .A(n8946), .B(n8947), .Z(n8945) );
  NANDN U17050 ( .A(n8948), .B(n8949), .Z(n8946) );
  NANDN U17051 ( .A(n8949), .B(n8948), .Z(n8944) );
  AND U17052 ( .A(n8950), .B(n8951), .Z(n8905) );
  NAND U17053 ( .A(n8952), .B(n8953), .Z(n8951) );
  OR U17054 ( .A(n8954), .B(n8955), .Z(n8952) );
  NANDN U17055 ( .A(n8956), .B(n8954), .Z(n8950) );
  XNOR U17056 ( .A(n8931), .B(n8957), .Z(N64597) );
  XOR U17057 ( .A(n8933), .B(n8934), .Z(n8957) );
  XNOR U17058 ( .A(n8947), .B(n8958), .Z(n8934) );
  XOR U17059 ( .A(n8948), .B(n8949), .Z(n8958) );
  XOR U17060 ( .A(n8954), .B(n8959), .Z(n8949) );
  XOR U17061 ( .A(n8953), .B(n8956), .Z(n8959) );
  IV U17062 ( .A(n8955), .Z(n8956) );
  NAND U17063 ( .A(n8960), .B(n8961), .Z(n8955) );
  OR U17064 ( .A(n8962), .B(n8963), .Z(n8961) );
  OR U17065 ( .A(n8964), .B(n8965), .Z(n8960) );
  NAND U17066 ( .A(n8966), .B(n8967), .Z(n8953) );
  OR U17067 ( .A(n8968), .B(n8969), .Z(n8967) );
  OR U17068 ( .A(n8970), .B(n8971), .Z(n8966) );
  NOR U17069 ( .A(n8972), .B(n8973), .Z(n8954) );
  ANDN U17070 ( .B(n8974), .A(n8975), .Z(n8948) );
  XNOR U17071 ( .A(n8941), .B(n8976), .Z(n8947) );
  XNOR U17072 ( .A(n8940), .B(n8942), .Z(n8976) );
  NAND U17073 ( .A(n8977), .B(n8978), .Z(n8942) );
  OR U17074 ( .A(n8979), .B(n8980), .Z(n8978) );
  OR U17075 ( .A(n8981), .B(n8982), .Z(n8977) );
  NAND U17076 ( .A(n8983), .B(n8984), .Z(n8940) );
  OR U17077 ( .A(n8985), .B(n8986), .Z(n8984) );
  OR U17078 ( .A(n8987), .B(n8988), .Z(n8983) );
  ANDN U17079 ( .B(n8989), .A(n8990), .Z(n8941) );
  IV U17080 ( .A(n8991), .Z(n8989) );
  ANDN U17081 ( .B(n8992), .A(n8993), .Z(n8933) );
  XOR U17082 ( .A(n8919), .B(n8994), .Z(n8931) );
  XOR U17083 ( .A(n8920), .B(n8921), .Z(n8994) );
  XOR U17084 ( .A(n8926), .B(n8995), .Z(n8921) );
  XOR U17085 ( .A(n8925), .B(n8928), .Z(n8995) );
  IV U17086 ( .A(n8927), .Z(n8928) );
  NAND U17087 ( .A(n8996), .B(n8997), .Z(n8927) );
  OR U17088 ( .A(n8998), .B(n8999), .Z(n8997) );
  OR U17089 ( .A(n9000), .B(n9001), .Z(n8996) );
  NAND U17090 ( .A(n9002), .B(n9003), .Z(n8925) );
  OR U17091 ( .A(n9004), .B(n9005), .Z(n9003) );
  OR U17092 ( .A(n9006), .B(n9007), .Z(n9002) );
  NOR U17093 ( .A(n9008), .B(n9009), .Z(n8926) );
  ANDN U17094 ( .B(n9010), .A(n9011), .Z(n8920) );
  IV U17095 ( .A(n9012), .Z(n9010) );
  XNOR U17096 ( .A(n8913), .B(n9013), .Z(n8919) );
  XNOR U17097 ( .A(n8912), .B(n8914), .Z(n9013) );
  NAND U17098 ( .A(n9014), .B(n9015), .Z(n8914) );
  OR U17099 ( .A(n9016), .B(n9017), .Z(n9015) );
  OR U17100 ( .A(n9018), .B(n9019), .Z(n9014) );
  NAND U17101 ( .A(n9020), .B(n9021), .Z(n8912) );
  OR U17102 ( .A(n9022), .B(n9023), .Z(n9021) );
  OR U17103 ( .A(n9024), .B(n9025), .Z(n9020) );
  ANDN U17104 ( .B(n9026), .A(n9027), .Z(n8913) );
  IV U17105 ( .A(n9028), .Z(n9026) );
  XNOR U17106 ( .A(n8993), .B(n8992), .Z(N64596) );
  XOR U17107 ( .A(n9012), .B(n9011), .Z(n8992) );
  XNOR U17108 ( .A(n9027), .B(n9028), .Z(n9011) );
  XNOR U17109 ( .A(n9022), .B(n9023), .Z(n9028) );
  XNOR U17110 ( .A(n9024), .B(n9025), .Z(n9023) );
  XNOR U17111 ( .A(y[7405]), .B(x[7405]), .Z(n9025) );
  XNOR U17112 ( .A(y[7406]), .B(x[7406]), .Z(n9024) );
  XNOR U17113 ( .A(y[7404]), .B(x[7404]), .Z(n9022) );
  XNOR U17114 ( .A(n9016), .B(n9017), .Z(n9027) );
  XNOR U17115 ( .A(y[7401]), .B(x[7401]), .Z(n9017) );
  XNOR U17116 ( .A(n9018), .B(n9019), .Z(n9016) );
  XNOR U17117 ( .A(y[7402]), .B(x[7402]), .Z(n9019) );
  XNOR U17118 ( .A(y[7403]), .B(x[7403]), .Z(n9018) );
  XNOR U17119 ( .A(n9009), .B(n9008), .Z(n9012) );
  XNOR U17120 ( .A(n9004), .B(n9005), .Z(n9008) );
  XNOR U17121 ( .A(y[7398]), .B(x[7398]), .Z(n9005) );
  XNOR U17122 ( .A(n9006), .B(n9007), .Z(n9004) );
  XNOR U17123 ( .A(y[7399]), .B(x[7399]), .Z(n9007) );
  XNOR U17124 ( .A(y[7400]), .B(x[7400]), .Z(n9006) );
  XNOR U17125 ( .A(n8998), .B(n8999), .Z(n9009) );
  XNOR U17126 ( .A(y[7395]), .B(x[7395]), .Z(n8999) );
  XNOR U17127 ( .A(n9000), .B(n9001), .Z(n8998) );
  XNOR U17128 ( .A(y[7396]), .B(x[7396]), .Z(n9001) );
  XNOR U17129 ( .A(y[7397]), .B(x[7397]), .Z(n9000) );
  XOR U17130 ( .A(n8974), .B(n8975), .Z(n8993) );
  XNOR U17131 ( .A(n8990), .B(n8991), .Z(n8975) );
  XNOR U17132 ( .A(n8985), .B(n8986), .Z(n8991) );
  XNOR U17133 ( .A(n8987), .B(n8988), .Z(n8986) );
  XNOR U17134 ( .A(y[7393]), .B(x[7393]), .Z(n8988) );
  XNOR U17135 ( .A(y[7394]), .B(x[7394]), .Z(n8987) );
  XNOR U17136 ( .A(y[7392]), .B(x[7392]), .Z(n8985) );
  XNOR U17137 ( .A(n8979), .B(n8980), .Z(n8990) );
  XNOR U17138 ( .A(y[7389]), .B(x[7389]), .Z(n8980) );
  XNOR U17139 ( .A(n8981), .B(n8982), .Z(n8979) );
  XNOR U17140 ( .A(y[7390]), .B(x[7390]), .Z(n8982) );
  XNOR U17141 ( .A(y[7391]), .B(x[7391]), .Z(n8981) );
  XOR U17142 ( .A(n8973), .B(n8972), .Z(n8974) );
  XNOR U17143 ( .A(n8968), .B(n8969), .Z(n8972) );
  XNOR U17144 ( .A(y[7386]), .B(x[7386]), .Z(n8969) );
  XNOR U17145 ( .A(n8970), .B(n8971), .Z(n8968) );
  XNOR U17146 ( .A(y[7387]), .B(x[7387]), .Z(n8971) );
  XNOR U17147 ( .A(y[7388]), .B(x[7388]), .Z(n8970) );
  XNOR U17148 ( .A(n8962), .B(n8963), .Z(n8973) );
  XNOR U17149 ( .A(y[7383]), .B(x[7383]), .Z(n8963) );
  XNOR U17150 ( .A(n8964), .B(n8965), .Z(n8962) );
  XNOR U17151 ( .A(y[7384]), .B(x[7384]), .Z(n8965) );
  XNOR U17152 ( .A(y[7385]), .B(x[7385]), .Z(n8964) );
  NAND U17153 ( .A(n9029), .B(n9030), .Z(N64587) );
  NANDN U17154 ( .A(n9031), .B(n9032), .Z(n9030) );
  OR U17155 ( .A(n9033), .B(n9034), .Z(n9032) );
  NAND U17156 ( .A(n9033), .B(n9034), .Z(n9029) );
  XOR U17157 ( .A(n9033), .B(n9035), .Z(N64586) );
  XNOR U17158 ( .A(n9031), .B(n9034), .Z(n9035) );
  AND U17159 ( .A(n9036), .B(n9037), .Z(n9034) );
  NANDN U17160 ( .A(n9038), .B(n9039), .Z(n9037) );
  NANDN U17161 ( .A(n9040), .B(n9041), .Z(n9039) );
  NANDN U17162 ( .A(n9041), .B(n9040), .Z(n9036) );
  NAND U17163 ( .A(n9042), .B(n9043), .Z(n9031) );
  NANDN U17164 ( .A(n9044), .B(n9045), .Z(n9043) );
  OR U17165 ( .A(n9046), .B(n9047), .Z(n9045) );
  NAND U17166 ( .A(n9047), .B(n9046), .Z(n9042) );
  AND U17167 ( .A(n9048), .B(n9049), .Z(n9033) );
  NANDN U17168 ( .A(n9050), .B(n9051), .Z(n9049) );
  NANDN U17169 ( .A(n9052), .B(n9053), .Z(n9051) );
  NANDN U17170 ( .A(n9053), .B(n9052), .Z(n9048) );
  XOR U17171 ( .A(n9047), .B(n9054), .Z(N64585) );
  XOR U17172 ( .A(n9044), .B(n9046), .Z(n9054) );
  XNOR U17173 ( .A(n9040), .B(n9055), .Z(n9046) );
  XNOR U17174 ( .A(n9038), .B(n9041), .Z(n9055) );
  NAND U17175 ( .A(n9056), .B(n9057), .Z(n9041) );
  NAND U17176 ( .A(n9058), .B(n9059), .Z(n9057) );
  OR U17177 ( .A(n9060), .B(n9061), .Z(n9058) );
  NANDN U17178 ( .A(n9062), .B(n9060), .Z(n9056) );
  IV U17179 ( .A(n9061), .Z(n9062) );
  NAND U17180 ( .A(n9063), .B(n9064), .Z(n9038) );
  NAND U17181 ( .A(n9065), .B(n9066), .Z(n9064) );
  NANDN U17182 ( .A(n9067), .B(n9068), .Z(n9065) );
  NANDN U17183 ( .A(n9068), .B(n9067), .Z(n9063) );
  AND U17184 ( .A(n9069), .B(n9070), .Z(n9040) );
  NAND U17185 ( .A(n9071), .B(n9072), .Z(n9070) );
  OR U17186 ( .A(n9073), .B(n9074), .Z(n9071) );
  NANDN U17187 ( .A(n9075), .B(n9073), .Z(n9069) );
  NAND U17188 ( .A(n9076), .B(n9077), .Z(n9044) );
  NANDN U17189 ( .A(n9078), .B(n9079), .Z(n9077) );
  OR U17190 ( .A(n9080), .B(n9081), .Z(n9079) );
  NANDN U17191 ( .A(n9082), .B(n9080), .Z(n9076) );
  IV U17192 ( .A(n9081), .Z(n9082) );
  XNOR U17193 ( .A(n9052), .B(n9083), .Z(n9047) );
  XNOR U17194 ( .A(n9050), .B(n9053), .Z(n9083) );
  NAND U17195 ( .A(n9084), .B(n9085), .Z(n9053) );
  NAND U17196 ( .A(n9086), .B(n9087), .Z(n9085) );
  OR U17197 ( .A(n9088), .B(n9089), .Z(n9086) );
  NANDN U17198 ( .A(n9090), .B(n9088), .Z(n9084) );
  IV U17199 ( .A(n9089), .Z(n9090) );
  NAND U17200 ( .A(n9091), .B(n9092), .Z(n9050) );
  NAND U17201 ( .A(n9093), .B(n9094), .Z(n9092) );
  NANDN U17202 ( .A(n9095), .B(n9096), .Z(n9093) );
  NANDN U17203 ( .A(n9096), .B(n9095), .Z(n9091) );
  AND U17204 ( .A(n9097), .B(n9098), .Z(n9052) );
  NAND U17205 ( .A(n9099), .B(n9100), .Z(n9098) );
  OR U17206 ( .A(n9101), .B(n9102), .Z(n9099) );
  NANDN U17207 ( .A(n9103), .B(n9101), .Z(n9097) );
  XNOR U17208 ( .A(n9078), .B(n9104), .Z(N64584) );
  XOR U17209 ( .A(n9080), .B(n9081), .Z(n9104) );
  XNOR U17210 ( .A(n9094), .B(n9105), .Z(n9081) );
  XOR U17211 ( .A(n9095), .B(n9096), .Z(n9105) );
  XOR U17212 ( .A(n9101), .B(n9106), .Z(n9096) );
  XOR U17213 ( .A(n9100), .B(n9103), .Z(n9106) );
  IV U17214 ( .A(n9102), .Z(n9103) );
  NAND U17215 ( .A(n9107), .B(n9108), .Z(n9102) );
  OR U17216 ( .A(n9109), .B(n9110), .Z(n9108) );
  OR U17217 ( .A(n9111), .B(n9112), .Z(n9107) );
  NAND U17218 ( .A(n9113), .B(n9114), .Z(n9100) );
  OR U17219 ( .A(n9115), .B(n9116), .Z(n9114) );
  OR U17220 ( .A(n9117), .B(n9118), .Z(n9113) );
  NOR U17221 ( .A(n9119), .B(n9120), .Z(n9101) );
  ANDN U17222 ( .B(n9121), .A(n9122), .Z(n9095) );
  XNOR U17223 ( .A(n9088), .B(n9123), .Z(n9094) );
  XNOR U17224 ( .A(n9087), .B(n9089), .Z(n9123) );
  NAND U17225 ( .A(n9124), .B(n9125), .Z(n9089) );
  OR U17226 ( .A(n9126), .B(n9127), .Z(n9125) );
  OR U17227 ( .A(n9128), .B(n9129), .Z(n9124) );
  NAND U17228 ( .A(n9130), .B(n9131), .Z(n9087) );
  OR U17229 ( .A(n9132), .B(n9133), .Z(n9131) );
  OR U17230 ( .A(n9134), .B(n9135), .Z(n9130) );
  ANDN U17231 ( .B(n9136), .A(n9137), .Z(n9088) );
  IV U17232 ( .A(n9138), .Z(n9136) );
  ANDN U17233 ( .B(n9139), .A(n9140), .Z(n9080) );
  XOR U17234 ( .A(n9066), .B(n9141), .Z(n9078) );
  XOR U17235 ( .A(n9067), .B(n9068), .Z(n9141) );
  XOR U17236 ( .A(n9073), .B(n9142), .Z(n9068) );
  XOR U17237 ( .A(n9072), .B(n9075), .Z(n9142) );
  IV U17238 ( .A(n9074), .Z(n9075) );
  NAND U17239 ( .A(n9143), .B(n9144), .Z(n9074) );
  OR U17240 ( .A(n9145), .B(n9146), .Z(n9144) );
  OR U17241 ( .A(n9147), .B(n9148), .Z(n9143) );
  NAND U17242 ( .A(n9149), .B(n9150), .Z(n9072) );
  OR U17243 ( .A(n9151), .B(n9152), .Z(n9150) );
  OR U17244 ( .A(n9153), .B(n9154), .Z(n9149) );
  NOR U17245 ( .A(n9155), .B(n9156), .Z(n9073) );
  ANDN U17246 ( .B(n9157), .A(n9158), .Z(n9067) );
  IV U17247 ( .A(n9159), .Z(n9157) );
  XNOR U17248 ( .A(n9060), .B(n9160), .Z(n9066) );
  XNOR U17249 ( .A(n9059), .B(n9061), .Z(n9160) );
  NAND U17250 ( .A(n9161), .B(n9162), .Z(n9061) );
  OR U17251 ( .A(n9163), .B(n9164), .Z(n9162) );
  OR U17252 ( .A(n9165), .B(n9166), .Z(n9161) );
  NAND U17253 ( .A(n9167), .B(n9168), .Z(n9059) );
  OR U17254 ( .A(n9169), .B(n9170), .Z(n9168) );
  OR U17255 ( .A(n9171), .B(n9172), .Z(n9167) );
  ANDN U17256 ( .B(n9173), .A(n9174), .Z(n9060) );
  IV U17257 ( .A(n9175), .Z(n9173) );
  XNOR U17258 ( .A(n9140), .B(n9139), .Z(N64583) );
  XOR U17259 ( .A(n9159), .B(n9158), .Z(n9139) );
  XNOR U17260 ( .A(n9174), .B(n9175), .Z(n9158) );
  XNOR U17261 ( .A(n9169), .B(n9170), .Z(n9175) );
  XNOR U17262 ( .A(n9171), .B(n9172), .Z(n9170) );
  XNOR U17263 ( .A(y[7381]), .B(x[7381]), .Z(n9172) );
  XNOR U17264 ( .A(y[7382]), .B(x[7382]), .Z(n9171) );
  XNOR U17265 ( .A(y[7380]), .B(x[7380]), .Z(n9169) );
  XNOR U17266 ( .A(n9163), .B(n9164), .Z(n9174) );
  XNOR U17267 ( .A(y[7377]), .B(x[7377]), .Z(n9164) );
  XNOR U17268 ( .A(n9165), .B(n9166), .Z(n9163) );
  XNOR U17269 ( .A(y[7378]), .B(x[7378]), .Z(n9166) );
  XNOR U17270 ( .A(y[7379]), .B(x[7379]), .Z(n9165) );
  XNOR U17271 ( .A(n9156), .B(n9155), .Z(n9159) );
  XNOR U17272 ( .A(n9151), .B(n9152), .Z(n9155) );
  XNOR U17273 ( .A(y[7374]), .B(x[7374]), .Z(n9152) );
  XNOR U17274 ( .A(n9153), .B(n9154), .Z(n9151) );
  XNOR U17275 ( .A(y[7375]), .B(x[7375]), .Z(n9154) );
  XNOR U17276 ( .A(y[7376]), .B(x[7376]), .Z(n9153) );
  XNOR U17277 ( .A(n9145), .B(n9146), .Z(n9156) );
  XNOR U17278 ( .A(y[7371]), .B(x[7371]), .Z(n9146) );
  XNOR U17279 ( .A(n9147), .B(n9148), .Z(n9145) );
  XNOR U17280 ( .A(y[7372]), .B(x[7372]), .Z(n9148) );
  XNOR U17281 ( .A(y[7373]), .B(x[7373]), .Z(n9147) );
  XOR U17282 ( .A(n9121), .B(n9122), .Z(n9140) );
  XNOR U17283 ( .A(n9137), .B(n9138), .Z(n9122) );
  XNOR U17284 ( .A(n9132), .B(n9133), .Z(n9138) );
  XNOR U17285 ( .A(n9134), .B(n9135), .Z(n9133) );
  XNOR U17286 ( .A(y[7369]), .B(x[7369]), .Z(n9135) );
  XNOR U17287 ( .A(y[7370]), .B(x[7370]), .Z(n9134) );
  XNOR U17288 ( .A(y[7368]), .B(x[7368]), .Z(n9132) );
  XNOR U17289 ( .A(n9126), .B(n9127), .Z(n9137) );
  XNOR U17290 ( .A(y[7365]), .B(x[7365]), .Z(n9127) );
  XNOR U17291 ( .A(n9128), .B(n9129), .Z(n9126) );
  XNOR U17292 ( .A(y[7366]), .B(x[7366]), .Z(n9129) );
  XNOR U17293 ( .A(y[7367]), .B(x[7367]), .Z(n9128) );
  XOR U17294 ( .A(n9120), .B(n9119), .Z(n9121) );
  XNOR U17295 ( .A(n9115), .B(n9116), .Z(n9119) );
  XNOR U17296 ( .A(y[7362]), .B(x[7362]), .Z(n9116) );
  XNOR U17297 ( .A(n9117), .B(n9118), .Z(n9115) );
  XNOR U17298 ( .A(y[7363]), .B(x[7363]), .Z(n9118) );
  XNOR U17299 ( .A(y[7364]), .B(x[7364]), .Z(n9117) );
  XNOR U17300 ( .A(n9109), .B(n9110), .Z(n9120) );
  XNOR U17301 ( .A(y[7359]), .B(x[7359]), .Z(n9110) );
  XNOR U17302 ( .A(n9111), .B(n9112), .Z(n9109) );
  XNOR U17303 ( .A(y[7360]), .B(x[7360]), .Z(n9112) );
  XNOR U17304 ( .A(y[7361]), .B(x[7361]), .Z(n9111) );
  NAND U17305 ( .A(n9176), .B(n9177), .Z(N64574) );
  NANDN U17306 ( .A(n9178), .B(n9179), .Z(n9177) );
  OR U17307 ( .A(n9180), .B(n9181), .Z(n9179) );
  NAND U17308 ( .A(n9180), .B(n9181), .Z(n9176) );
  XOR U17309 ( .A(n9180), .B(n9182), .Z(N64573) );
  XNOR U17310 ( .A(n9178), .B(n9181), .Z(n9182) );
  AND U17311 ( .A(n9183), .B(n9184), .Z(n9181) );
  NANDN U17312 ( .A(n9185), .B(n9186), .Z(n9184) );
  NANDN U17313 ( .A(n9187), .B(n9188), .Z(n9186) );
  NANDN U17314 ( .A(n9188), .B(n9187), .Z(n9183) );
  NAND U17315 ( .A(n9189), .B(n9190), .Z(n9178) );
  NANDN U17316 ( .A(n9191), .B(n9192), .Z(n9190) );
  OR U17317 ( .A(n9193), .B(n9194), .Z(n9192) );
  NAND U17318 ( .A(n9194), .B(n9193), .Z(n9189) );
  AND U17319 ( .A(n9195), .B(n9196), .Z(n9180) );
  NANDN U17320 ( .A(n9197), .B(n9198), .Z(n9196) );
  NANDN U17321 ( .A(n9199), .B(n9200), .Z(n9198) );
  NANDN U17322 ( .A(n9200), .B(n9199), .Z(n9195) );
  XOR U17323 ( .A(n9194), .B(n9201), .Z(N64572) );
  XOR U17324 ( .A(n9191), .B(n9193), .Z(n9201) );
  XNOR U17325 ( .A(n9187), .B(n9202), .Z(n9193) );
  XNOR U17326 ( .A(n9185), .B(n9188), .Z(n9202) );
  NAND U17327 ( .A(n9203), .B(n9204), .Z(n9188) );
  NAND U17328 ( .A(n9205), .B(n9206), .Z(n9204) );
  OR U17329 ( .A(n9207), .B(n9208), .Z(n9205) );
  NANDN U17330 ( .A(n9209), .B(n9207), .Z(n9203) );
  IV U17331 ( .A(n9208), .Z(n9209) );
  NAND U17332 ( .A(n9210), .B(n9211), .Z(n9185) );
  NAND U17333 ( .A(n9212), .B(n9213), .Z(n9211) );
  NANDN U17334 ( .A(n9214), .B(n9215), .Z(n9212) );
  NANDN U17335 ( .A(n9215), .B(n9214), .Z(n9210) );
  AND U17336 ( .A(n9216), .B(n9217), .Z(n9187) );
  NAND U17337 ( .A(n9218), .B(n9219), .Z(n9217) );
  OR U17338 ( .A(n9220), .B(n9221), .Z(n9218) );
  NANDN U17339 ( .A(n9222), .B(n9220), .Z(n9216) );
  NAND U17340 ( .A(n9223), .B(n9224), .Z(n9191) );
  NANDN U17341 ( .A(n9225), .B(n9226), .Z(n9224) );
  OR U17342 ( .A(n9227), .B(n9228), .Z(n9226) );
  NANDN U17343 ( .A(n9229), .B(n9227), .Z(n9223) );
  IV U17344 ( .A(n9228), .Z(n9229) );
  XNOR U17345 ( .A(n9199), .B(n9230), .Z(n9194) );
  XNOR U17346 ( .A(n9197), .B(n9200), .Z(n9230) );
  NAND U17347 ( .A(n9231), .B(n9232), .Z(n9200) );
  NAND U17348 ( .A(n9233), .B(n9234), .Z(n9232) );
  OR U17349 ( .A(n9235), .B(n9236), .Z(n9233) );
  NANDN U17350 ( .A(n9237), .B(n9235), .Z(n9231) );
  IV U17351 ( .A(n9236), .Z(n9237) );
  NAND U17352 ( .A(n9238), .B(n9239), .Z(n9197) );
  NAND U17353 ( .A(n9240), .B(n9241), .Z(n9239) );
  NANDN U17354 ( .A(n9242), .B(n9243), .Z(n9240) );
  NANDN U17355 ( .A(n9243), .B(n9242), .Z(n9238) );
  AND U17356 ( .A(n9244), .B(n9245), .Z(n9199) );
  NAND U17357 ( .A(n9246), .B(n9247), .Z(n9245) );
  OR U17358 ( .A(n9248), .B(n9249), .Z(n9246) );
  NANDN U17359 ( .A(n9250), .B(n9248), .Z(n9244) );
  XNOR U17360 ( .A(n9225), .B(n9251), .Z(N64571) );
  XOR U17361 ( .A(n9227), .B(n9228), .Z(n9251) );
  XNOR U17362 ( .A(n9241), .B(n9252), .Z(n9228) );
  XOR U17363 ( .A(n9242), .B(n9243), .Z(n9252) );
  XOR U17364 ( .A(n9248), .B(n9253), .Z(n9243) );
  XOR U17365 ( .A(n9247), .B(n9250), .Z(n9253) );
  IV U17366 ( .A(n9249), .Z(n9250) );
  NAND U17367 ( .A(n9254), .B(n9255), .Z(n9249) );
  OR U17368 ( .A(n9256), .B(n9257), .Z(n9255) );
  OR U17369 ( .A(n9258), .B(n9259), .Z(n9254) );
  NAND U17370 ( .A(n9260), .B(n9261), .Z(n9247) );
  OR U17371 ( .A(n9262), .B(n9263), .Z(n9261) );
  OR U17372 ( .A(n9264), .B(n9265), .Z(n9260) );
  NOR U17373 ( .A(n9266), .B(n9267), .Z(n9248) );
  ANDN U17374 ( .B(n9268), .A(n9269), .Z(n9242) );
  XNOR U17375 ( .A(n9235), .B(n9270), .Z(n9241) );
  XNOR U17376 ( .A(n9234), .B(n9236), .Z(n9270) );
  NAND U17377 ( .A(n9271), .B(n9272), .Z(n9236) );
  OR U17378 ( .A(n9273), .B(n9274), .Z(n9272) );
  OR U17379 ( .A(n9275), .B(n9276), .Z(n9271) );
  NAND U17380 ( .A(n9277), .B(n9278), .Z(n9234) );
  OR U17381 ( .A(n9279), .B(n9280), .Z(n9278) );
  OR U17382 ( .A(n9281), .B(n9282), .Z(n9277) );
  ANDN U17383 ( .B(n9283), .A(n9284), .Z(n9235) );
  IV U17384 ( .A(n9285), .Z(n9283) );
  ANDN U17385 ( .B(n9286), .A(n9287), .Z(n9227) );
  XOR U17386 ( .A(n9213), .B(n9288), .Z(n9225) );
  XOR U17387 ( .A(n9214), .B(n9215), .Z(n9288) );
  XOR U17388 ( .A(n9220), .B(n9289), .Z(n9215) );
  XOR U17389 ( .A(n9219), .B(n9222), .Z(n9289) );
  IV U17390 ( .A(n9221), .Z(n9222) );
  NAND U17391 ( .A(n9290), .B(n9291), .Z(n9221) );
  OR U17392 ( .A(n9292), .B(n9293), .Z(n9291) );
  OR U17393 ( .A(n9294), .B(n9295), .Z(n9290) );
  NAND U17394 ( .A(n9296), .B(n9297), .Z(n9219) );
  OR U17395 ( .A(n9298), .B(n9299), .Z(n9297) );
  OR U17396 ( .A(n9300), .B(n9301), .Z(n9296) );
  NOR U17397 ( .A(n9302), .B(n9303), .Z(n9220) );
  ANDN U17398 ( .B(n9304), .A(n9305), .Z(n9214) );
  IV U17399 ( .A(n9306), .Z(n9304) );
  XNOR U17400 ( .A(n9207), .B(n9307), .Z(n9213) );
  XNOR U17401 ( .A(n9206), .B(n9208), .Z(n9307) );
  NAND U17402 ( .A(n9308), .B(n9309), .Z(n9208) );
  OR U17403 ( .A(n9310), .B(n9311), .Z(n9309) );
  OR U17404 ( .A(n9312), .B(n9313), .Z(n9308) );
  NAND U17405 ( .A(n9314), .B(n9315), .Z(n9206) );
  OR U17406 ( .A(n9316), .B(n9317), .Z(n9315) );
  OR U17407 ( .A(n9318), .B(n9319), .Z(n9314) );
  ANDN U17408 ( .B(n9320), .A(n9321), .Z(n9207) );
  IV U17409 ( .A(n9322), .Z(n9320) );
  XNOR U17410 ( .A(n9287), .B(n9286), .Z(N64570) );
  XOR U17411 ( .A(n9306), .B(n9305), .Z(n9286) );
  XNOR U17412 ( .A(n9321), .B(n9322), .Z(n9305) );
  XNOR U17413 ( .A(n9316), .B(n9317), .Z(n9322) );
  XNOR U17414 ( .A(n9318), .B(n9319), .Z(n9317) );
  XNOR U17415 ( .A(y[7357]), .B(x[7357]), .Z(n9319) );
  XNOR U17416 ( .A(y[7358]), .B(x[7358]), .Z(n9318) );
  XNOR U17417 ( .A(y[7356]), .B(x[7356]), .Z(n9316) );
  XNOR U17418 ( .A(n9310), .B(n9311), .Z(n9321) );
  XNOR U17419 ( .A(y[7353]), .B(x[7353]), .Z(n9311) );
  XNOR U17420 ( .A(n9312), .B(n9313), .Z(n9310) );
  XNOR U17421 ( .A(y[7354]), .B(x[7354]), .Z(n9313) );
  XNOR U17422 ( .A(y[7355]), .B(x[7355]), .Z(n9312) );
  XNOR U17423 ( .A(n9303), .B(n9302), .Z(n9306) );
  XNOR U17424 ( .A(n9298), .B(n9299), .Z(n9302) );
  XNOR U17425 ( .A(y[7350]), .B(x[7350]), .Z(n9299) );
  XNOR U17426 ( .A(n9300), .B(n9301), .Z(n9298) );
  XNOR U17427 ( .A(y[7351]), .B(x[7351]), .Z(n9301) );
  XNOR U17428 ( .A(y[7352]), .B(x[7352]), .Z(n9300) );
  XNOR U17429 ( .A(n9292), .B(n9293), .Z(n9303) );
  XNOR U17430 ( .A(y[7347]), .B(x[7347]), .Z(n9293) );
  XNOR U17431 ( .A(n9294), .B(n9295), .Z(n9292) );
  XNOR U17432 ( .A(y[7348]), .B(x[7348]), .Z(n9295) );
  XNOR U17433 ( .A(y[7349]), .B(x[7349]), .Z(n9294) );
  XOR U17434 ( .A(n9268), .B(n9269), .Z(n9287) );
  XNOR U17435 ( .A(n9284), .B(n9285), .Z(n9269) );
  XNOR U17436 ( .A(n9279), .B(n9280), .Z(n9285) );
  XNOR U17437 ( .A(n9281), .B(n9282), .Z(n9280) );
  XNOR U17438 ( .A(y[7345]), .B(x[7345]), .Z(n9282) );
  XNOR U17439 ( .A(y[7346]), .B(x[7346]), .Z(n9281) );
  XNOR U17440 ( .A(y[7344]), .B(x[7344]), .Z(n9279) );
  XNOR U17441 ( .A(n9273), .B(n9274), .Z(n9284) );
  XNOR U17442 ( .A(y[7341]), .B(x[7341]), .Z(n9274) );
  XNOR U17443 ( .A(n9275), .B(n9276), .Z(n9273) );
  XNOR U17444 ( .A(y[7342]), .B(x[7342]), .Z(n9276) );
  XNOR U17445 ( .A(y[7343]), .B(x[7343]), .Z(n9275) );
  XOR U17446 ( .A(n9267), .B(n9266), .Z(n9268) );
  XNOR U17447 ( .A(n9262), .B(n9263), .Z(n9266) );
  XNOR U17448 ( .A(y[7338]), .B(x[7338]), .Z(n9263) );
  XNOR U17449 ( .A(n9264), .B(n9265), .Z(n9262) );
  XNOR U17450 ( .A(y[7339]), .B(x[7339]), .Z(n9265) );
  XNOR U17451 ( .A(y[7340]), .B(x[7340]), .Z(n9264) );
  XNOR U17452 ( .A(n9256), .B(n9257), .Z(n9267) );
  XNOR U17453 ( .A(y[7335]), .B(x[7335]), .Z(n9257) );
  XNOR U17454 ( .A(n9258), .B(n9259), .Z(n9256) );
  XNOR U17455 ( .A(y[7336]), .B(x[7336]), .Z(n9259) );
  XNOR U17456 ( .A(y[7337]), .B(x[7337]), .Z(n9258) );
  NAND U17457 ( .A(n9323), .B(n9324), .Z(N64561) );
  NANDN U17458 ( .A(n9325), .B(n9326), .Z(n9324) );
  OR U17459 ( .A(n9327), .B(n9328), .Z(n9326) );
  NAND U17460 ( .A(n9327), .B(n9328), .Z(n9323) );
  XOR U17461 ( .A(n9327), .B(n9329), .Z(N64560) );
  XNOR U17462 ( .A(n9325), .B(n9328), .Z(n9329) );
  AND U17463 ( .A(n9330), .B(n9331), .Z(n9328) );
  NANDN U17464 ( .A(n9332), .B(n9333), .Z(n9331) );
  NANDN U17465 ( .A(n9334), .B(n9335), .Z(n9333) );
  NANDN U17466 ( .A(n9335), .B(n9334), .Z(n9330) );
  NAND U17467 ( .A(n9336), .B(n9337), .Z(n9325) );
  NANDN U17468 ( .A(n9338), .B(n9339), .Z(n9337) );
  OR U17469 ( .A(n9340), .B(n9341), .Z(n9339) );
  NAND U17470 ( .A(n9341), .B(n9340), .Z(n9336) );
  AND U17471 ( .A(n9342), .B(n9343), .Z(n9327) );
  NANDN U17472 ( .A(n9344), .B(n9345), .Z(n9343) );
  NANDN U17473 ( .A(n9346), .B(n9347), .Z(n9345) );
  NANDN U17474 ( .A(n9347), .B(n9346), .Z(n9342) );
  XOR U17475 ( .A(n9341), .B(n9348), .Z(N64559) );
  XOR U17476 ( .A(n9338), .B(n9340), .Z(n9348) );
  XNOR U17477 ( .A(n9334), .B(n9349), .Z(n9340) );
  XNOR U17478 ( .A(n9332), .B(n9335), .Z(n9349) );
  NAND U17479 ( .A(n9350), .B(n9351), .Z(n9335) );
  NAND U17480 ( .A(n9352), .B(n9353), .Z(n9351) );
  OR U17481 ( .A(n9354), .B(n9355), .Z(n9352) );
  NANDN U17482 ( .A(n9356), .B(n9354), .Z(n9350) );
  IV U17483 ( .A(n9355), .Z(n9356) );
  NAND U17484 ( .A(n9357), .B(n9358), .Z(n9332) );
  NAND U17485 ( .A(n9359), .B(n9360), .Z(n9358) );
  NANDN U17486 ( .A(n9361), .B(n9362), .Z(n9359) );
  NANDN U17487 ( .A(n9362), .B(n9361), .Z(n9357) );
  AND U17488 ( .A(n9363), .B(n9364), .Z(n9334) );
  NAND U17489 ( .A(n9365), .B(n9366), .Z(n9364) );
  OR U17490 ( .A(n9367), .B(n9368), .Z(n9365) );
  NANDN U17491 ( .A(n9369), .B(n9367), .Z(n9363) );
  NAND U17492 ( .A(n9370), .B(n9371), .Z(n9338) );
  NANDN U17493 ( .A(n9372), .B(n9373), .Z(n9371) );
  OR U17494 ( .A(n9374), .B(n9375), .Z(n9373) );
  NANDN U17495 ( .A(n9376), .B(n9374), .Z(n9370) );
  IV U17496 ( .A(n9375), .Z(n9376) );
  XNOR U17497 ( .A(n9346), .B(n9377), .Z(n9341) );
  XNOR U17498 ( .A(n9344), .B(n9347), .Z(n9377) );
  NAND U17499 ( .A(n9378), .B(n9379), .Z(n9347) );
  NAND U17500 ( .A(n9380), .B(n9381), .Z(n9379) );
  OR U17501 ( .A(n9382), .B(n9383), .Z(n9380) );
  NANDN U17502 ( .A(n9384), .B(n9382), .Z(n9378) );
  IV U17503 ( .A(n9383), .Z(n9384) );
  NAND U17504 ( .A(n9385), .B(n9386), .Z(n9344) );
  NAND U17505 ( .A(n9387), .B(n9388), .Z(n9386) );
  NANDN U17506 ( .A(n9389), .B(n9390), .Z(n9387) );
  NANDN U17507 ( .A(n9390), .B(n9389), .Z(n9385) );
  AND U17508 ( .A(n9391), .B(n9392), .Z(n9346) );
  NAND U17509 ( .A(n9393), .B(n9394), .Z(n9392) );
  OR U17510 ( .A(n9395), .B(n9396), .Z(n9393) );
  NANDN U17511 ( .A(n9397), .B(n9395), .Z(n9391) );
  XNOR U17512 ( .A(n9372), .B(n9398), .Z(N64558) );
  XOR U17513 ( .A(n9374), .B(n9375), .Z(n9398) );
  XNOR U17514 ( .A(n9388), .B(n9399), .Z(n9375) );
  XOR U17515 ( .A(n9389), .B(n9390), .Z(n9399) );
  XOR U17516 ( .A(n9395), .B(n9400), .Z(n9390) );
  XOR U17517 ( .A(n9394), .B(n9397), .Z(n9400) );
  IV U17518 ( .A(n9396), .Z(n9397) );
  NAND U17519 ( .A(n9401), .B(n9402), .Z(n9396) );
  OR U17520 ( .A(n9403), .B(n9404), .Z(n9402) );
  OR U17521 ( .A(n9405), .B(n9406), .Z(n9401) );
  NAND U17522 ( .A(n9407), .B(n9408), .Z(n9394) );
  OR U17523 ( .A(n9409), .B(n9410), .Z(n9408) );
  OR U17524 ( .A(n9411), .B(n9412), .Z(n9407) );
  NOR U17525 ( .A(n9413), .B(n9414), .Z(n9395) );
  ANDN U17526 ( .B(n9415), .A(n9416), .Z(n9389) );
  XNOR U17527 ( .A(n9382), .B(n9417), .Z(n9388) );
  XNOR U17528 ( .A(n9381), .B(n9383), .Z(n9417) );
  NAND U17529 ( .A(n9418), .B(n9419), .Z(n9383) );
  OR U17530 ( .A(n9420), .B(n9421), .Z(n9419) );
  OR U17531 ( .A(n9422), .B(n9423), .Z(n9418) );
  NAND U17532 ( .A(n9424), .B(n9425), .Z(n9381) );
  OR U17533 ( .A(n9426), .B(n9427), .Z(n9425) );
  OR U17534 ( .A(n9428), .B(n9429), .Z(n9424) );
  ANDN U17535 ( .B(n9430), .A(n9431), .Z(n9382) );
  IV U17536 ( .A(n9432), .Z(n9430) );
  ANDN U17537 ( .B(n9433), .A(n9434), .Z(n9374) );
  XOR U17538 ( .A(n9360), .B(n9435), .Z(n9372) );
  XOR U17539 ( .A(n9361), .B(n9362), .Z(n9435) );
  XOR U17540 ( .A(n9367), .B(n9436), .Z(n9362) );
  XOR U17541 ( .A(n9366), .B(n9369), .Z(n9436) );
  IV U17542 ( .A(n9368), .Z(n9369) );
  NAND U17543 ( .A(n9437), .B(n9438), .Z(n9368) );
  OR U17544 ( .A(n9439), .B(n9440), .Z(n9438) );
  OR U17545 ( .A(n9441), .B(n9442), .Z(n9437) );
  NAND U17546 ( .A(n9443), .B(n9444), .Z(n9366) );
  OR U17547 ( .A(n9445), .B(n9446), .Z(n9444) );
  OR U17548 ( .A(n9447), .B(n9448), .Z(n9443) );
  NOR U17549 ( .A(n9449), .B(n9450), .Z(n9367) );
  ANDN U17550 ( .B(n9451), .A(n9452), .Z(n9361) );
  IV U17551 ( .A(n9453), .Z(n9451) );
  XNOR U17552 ( .A(n9354), .B(n9454), .Z(n9360) );
  XNOR U17553 ( .A(n9353), .B(n9355), .Z(n9454) );
  NAND U17554 ( .A(n9455), .B(n9456), .Z(n9355) );
  OR U17555 ( .A(n9457), .B(n9458), .Z(n9456) );
  OR U17556 ( .A(n9459), .B(n9460), .Z(n9455) );
  NAND U17557 ( .A(n9461), .B(n9462), .Z(n9353) );
  OR U17558 ( .A(n9463), .B(n9464), .Z(n9462) );
  OR U17559 ( .A(n9465), .B(n9466), .Z(n9461) );
  ANDN U17560 ( .B(n9467), .A(n9468), .Z(n9354) );
  IV U17561 ( .A(n9469), .Z(n9467) );
  XNOR U17562 ( .A(n9434), .B(n9433), .Z(N64557) );
  XOR U17563 ( .A(n9453), .B(n9452), .Z(n9433) );
  XNOR U17564 ( .A(n9468), .B(n9469), .Z(n9452) );
  XNOR U17565 ( .A(n9463), .B(n9464), .Z(n9469) );
  XNOR U17566 ( .A(n9465), .B(n9466), .Z(n9464) );
  XNOR U17567 ( .A(y[7333]), .B(x[7333]), .Z(n9466) );
  XNOR U17568 ( .A(y[7334]), .B(x[7334]), .Z(n9465) );
  XNOR U17569 ( .A(y[7332]), .B(x[7332]), .Z(n9463) );
  XNOR U17570 ( .A(n9457), .B(n9458), .Z(n9468) );
  XNOR U17571 ( .A(y[7329]), .B(x[7329]), .Z(n9458) );
  XNOR U17572 ( .A(n9459), .B(n9460), .Z(n9457) );
  XNOR U17573 ( .A(y[7330]), .B(x[7330]), .Z(n9460) );
  XNOR U17574 ( .A(y[7331]), .B(x[7331]), .Z(n9459) );
  XNOR U17575 ( .A(n9450), .B(n9449), .Z(n9453) );
  XNOR U17576 ( .A(n9445), .B(n9446), .Z(n9449) );
  XNOR U17577 ( .A(y[7326]), .B(x[7326]), .Z(n9446) );
  XNOR U17578 ( .A(n9447), .B(n9448), .Z(n9445) );
  XNOR U17579 ( .A(y[7327]), .B(x[7327]), .Z(n9448) );
  XNOR U17580 ( .A(y[7328]), .B(x[7328]), .Z(n9447) );
  XNOR U17581 ( .A(n9439), .B(n9440), .Z(n9450) );
  XNOR U17582 ( .A(y[7323]), .B(x[7323]), .Z(n9440) );
  XNOR U17583 ( .A(n9441), .B(n9442), .Z(n9439) );
  XNOR U17584 ( .A(y[7324]), .B(x[7324]), .Z(n9442) );
  XNOR U17585 ( .A(y[7325]), .B(x[7325]), .Z(n9441) );
  XOR U17586 ( .A(n9415), .B(n9416), .Z(n9434) );
  XNOR U17587 ( .A(n9431), .B(n9432), .Z(n9416) );
  XNOR U17588 ( .A(n9426), .B(n9427), .Z(n9432) );
  XNOR U17589 ( .A(n9428), .B(n9429), .Z(n9427) );
  XNOR U17590 ( .A(y[7321]), .B(x[7321]), .Z(n9429) );
  XNOR U17591 ( .A(y[7322]), .B(x[7322]), .Z(n9428) );
  XNOR U17592 ( .A(y[7320]), .B(x[7320]), .Z(n9426) );
  XNOR U17593 ( .A(n9420), .B(n9421), .Z(n9431) );
  XNOR U17594 ( .A(y[7317]), .B(x[7317]), .Z(n9421) );
  XNOR U17595 ( .A(n9422), .B(n9423), .Z(n9420) );
  XNOR U17596 ( .A(y[7318]), .B(x[7318]), .Z(n9423) );
  XNOR U17597 ( .A(y[7319]), .B(x[7319]), .Z(n9422) );
  XOR U17598 ( .A(n9414), .B(n9413), .Z(n9415) );
  XNOR U17599 ( .A(n9409), .B(n9410), .Z(n9413) );
  XNOR U17600 ( .A(y[7314]), .B(x[7314]), .Z(n9410) );
  XNOR U17601 ( .A(n9411), .B(n9412), .Z(n9409) );
  XNOR U17602 ( .A(y[7315]), .B(x[7315]), .Z(n9412) );
  XNOR U17603 ( .A(y[7316]), .B(x[7316]), .Z(n9411) );
  XNOR U17604 ( .A(n9403), .B(n9404), .Z(n9414) );
  XNOR U17605 ( .A(y[7311]), .B(x[7311]), .Z(n9404) );
  XNOR U17606 ( .A(n9405), .B(n9406), .Z(n9403) );
  XNOR U17607 ( .A(y[7312]), .B(x[7312]), .Z(n9406) );
  XNOR U17608 ( .A(y[7313]), .B(x[7313]), .Z(n9405) );
  NAND U17609 ( .A(n9470), .B(n9471), .Z(N64548) );
  NANDN U17610 ( .A(n9472), .B(n9473), .Z(n9471) );
  OR U17611 ( .A(n9474), .B(n9475), .Z(n9473) );
  NAND U17612 ( .A(n9474), .B(n9475), .Z(n9470) );
  XOR U17613 ( .A(n9474), .B(n9476), .Z(N64547) );
  XNOR U17614 ( .A(n9472), .B(n9475), .Z(n9476) );
  AND U17615 ( .A(n9477), .B(n9478), .Z(n9475) );
  NANDN U17616 ( .A(n9479), .B(n9480), .Z(n9478) );
  NANDN U17617 ( .A(n9481), .B(n9482), .Z(n9480) );
  NANDN U17618 ( .A(n9482), .B(n9481), .Z(n9477) );
  NAND U17619 ( .A(n9483), .B(n9484), .Z(n9472) );
  NANDN U17620 ( .A(n9485), .B(n9486), .Z(n9484) );
  OR U17621 ( .A(n9487), .B(n9488), .Z(n9486) );
  NAND U17622 ( .A(n9488), .B(n9487), .Z(n9483) );
  AND U17623 ( .A(n9489), .B(n9490), .Z(n9474) );
  NANDN U17624 ( .A(n9491), .B(n9492), .Z(n9490) );
  NANDN U17625 ( .A(n9493), .B(n9494), .Z(n9492) );
  NANDN U17626 ( .A(n9494), .B(n9493), .Z(n9489) );
  XOR U17627 ( .A(n9488), .B(n9495), .Z(N64546) );
  XOR U17628 ( .A(n9485), .B(n9487), .Z(n9495) );
  XNOR U17629 ( .A(n9481), .B(n9496), .Z(n9487) );
  XNOR U17630 ( .A(n9479), .B(n9482), .Z(n9496) );
  NAND U17631 ( .A(n9497), .B(n9498), .Z(n9482) );
  NAND U17632 ( .A(n9499), .B(n9500), .Z(n9498) );
  OR U17633 ( .A(n9501), .B(n9502), .Z(n9499) );
  NANDN U17634 ( .A(n9503), .B(n9501), .Z(n9497) );
  IV U17635 ( .A(n9502), .Z(n9503) );
  NAND U17636 ( .A(n9504), .B(n9505), .Z(n9479) );
  NAND U17637 ( .A(n9506), .B(n9507), .Z(n9505) );
  NANDN U17638 ( .A(n9508), .B(n9509), .Z(n9506) );
  NANDN U17639 ( .A(n9509), .B(n9508), .Z(n9504) );
  AND U17640 ( .A(n9510), .B(n9511), .Z(n9481) );
  NAND U17641 ( .A(n9512), .B(n9513), .Z(n9511) );
  OR U17642 ( .A(n9514), .B(n9515), .Z(n9512) );
  NANDN U17643 ( .A(n9516), .B(n9514), .Z(n9510) );
  NAND U17644 ( .A(n9517), .B(n9518), .Z(n9485) );
  NANDN U17645 ( .A(n9519), .B(n9520), .Z(n9518) );
  OR U17646 ( .A(n9521), .B(n9522), .Z(n9520) );
  NANDN U17647 ( .A(n9523), .B(n9521), .Z(n9517) );
  IV U17648 ( .A(n9522), .Z(n9523) );
  XNOR U17649 ( .A(n9493), .B(n9524), .Z(n9488) );
  XNOR U17650 ( .A(n9491), .B(n9494), .Z(n9524) );
  NAND U17651 ( .A(n9525), .B(n9526), .Z(n9494) );
  NAND U17652 ( .A(n9527), .B(n9528), .Z(n9526) );
  OR U17653 ( .A(n9529), .B(n9530), .Z(n9527) );
  NANDN U17654 ( .A(n9531), .B(n9529), .Z(n9525) );
  IV U17655 ( .A(n9530), .Z(n9531) );
  NAND U17656 ( .A(n9532), .B(n9533), .Z(n9491) );
  NAND U17657 ( .A(n9534), .B(n9535), .Z(n9533) );
  NANDN U17658 ( .A(n9536), .B(n9537), .Z(n9534) );
  NANDN U17659 ( .A(n9537), .B(n9536), .Z(n9532) );
  AND U17660 ( .A(n9538), .B(n9539), .Z(n9493) );
  NAND U17661 ( .A(n9540), .B(n9541), .Z(n9539) );
  OR U17662 ( .A(n9542), .B(n9543), .Z(n9540) );
  NANDN U17663 ( .A(n9544), .B(n9542), .Z(n9538) );
  XNOR U17664 ( .A(n9519), .B(n9545), .Z(N64545) );
  XOR U17665 ( .A(n9521), .B(n9522), .Z(n9545) );
  XNOR U17666 ( .A(n9535), .B(n9546), .Z(n9522) );
  XOR U17667 ( .A(n9536), .B(n9537), .Z(n9546) );
  XOR U17668 ( .A(n9542), .B(n9547), .Z(n9537) );
  XOR U17669 ( .A(n9541), .B(n9544), .Z(n9547) );
  IV U17670 ( .A(n9543), .Z(n9544) );
  NAND U17671 ( .A(n9548), .B(n9549), .Z(n9543) );
  OR U17672 ( .A(n9550), .B(n9551), .Z(n9549) );
  OR U17673 ( .A(n9552), .B(n9553), .Z(n9548) );
  NAND U17674 ( .A(n9554), .B(n9555), .Z(n9541) );
  OR U17675 ( .A(n9556), .B(n9557), .Z(n9555) );
  OR U17676 ( .A(n9558), .B(n9559), .Z(n9554) );
  NOR U17677 ( .A(n9560), .B(n9561), .Z(n9542) );
  ANDN U17678 ( .B(n9562), .A(n9563), .Z(n9536) );
  XNOR U17679 ( .A(n9529), .B(n9564), .Z(n9535) );
  XNOR U17680 ( .A(n9528), .B(n9530), .Z(n9564) );
  NAND U17681 ( .A(n9565), .B(n9566), .Z(n9530) );
  OR U17682 ( .A(n9567), .B(n9568), .Z(n9566) );
  OR U17683 ( .A(n9569), .B(n9570), .Z(n9565) );
  NAND U17684 ( .A(n9571), .B(n9572), .Z(n9528) );
  OR U17685 ( .A(n9573), .B(n9574), .Z(n9572) );
  OR U17686 ( .A(n9575), .B(n9576), .Z(n9571) );
  ANDN U17687 ( .B(n9577), .A(n9578), .Z(n9529) );
  IV U17688 ( .A(n9579), .Z(n9577) );
  ANDN U17689 ( .B(n9580), .A(n9581), .Z(n9521) );
  XOR U17690 ( .A(n9507), .B(n9582), .Z(n9519) );
  XOR U17691 ( .A(n9508), .B(n9509), .Z(n9582) );
  XOR U17692 ( .A(n9514), .B(n9583), .Z(n9509) );
  XOR U17693 ( .A(n9513), .B(n9516), .Z(n9583) );
  IV U17694 ( .A(n9515), .Z(n9516) );
  NAND U17695 ( .A(n9584), .B(n9585), .Z(n9515) );
  OR U17696 ( .A(n9586), .B(n9587), .Z(n9585) );
  OR U17697 ( .A(n9588), .B(n9589), .Z(n9584) );
  NAND U17698 ( .A(n9590), .B(n9591), .Z(n9513) );
  OR U17699 ( .A(n9592), .B(n9593), .Z(n9591) );
  OR U17700 ( .A(n9594), .B(n9595), .Z(n9590) );
  NOR U17701 ( .A(n9596), .B(n9597), .Z(n9514) );
  ANDN U17702 ( .B(n9598), .A(n9599), .Z(n9508) );
  IV U17703 ( .A(n9600), .Z(n9598) );
  XNOR U17704 ( .A(n9501), .B(n9601), .Z(n9507) );
  XNOR U17705 ( .A(n9500), .B(n9502), .Z(n9601) );
  NAND U17706 ( .A(n9602), .B(n9603), .Z(n9502) );
  OR U17707 ( .A(n9604), .B(n9605), .Z(n9603) );
  OR U17708 ( .A(n9606), .B(n9607), .Z(n9602) );
  NAND U17709 ( .A(n9608), .B(n9609), .Z(n9500) );
  OR U17710 ( .A(n9610), .B(n9611), .Z(n9609) );
  OR U17711 ( .A(n9612), .B(n9613), .Z(n9608) );
  ANDN U17712 ( .B(n9614), .A(n9615), .Z(n9501) );
  IV U17713 ( .A(n9616), .Z(n9614) );
  XNOR U17714 ( .A(n9581), .B(n9580), .Z(N64544) );
  XOR U17715 ( .A(n9600), .B(n9599), .Z(n9580) );
  XNOR U17716 ( .A(n9615), .B(n9616), .Z(n9599) );
  XNOR U17717 ( .A(n9610), .B(n9611), .Z(n9616) );
  XNOR U17718 ( .A(n9612), .B(n9613), .Z(n9611) );
  XNOR U17719 ( .A(y[7309]), .B(x[7309]), .Z(n9613) );
  XNOR U17720 ( .A(y[7310]), .B(x[7310]), .Z(n9612) );
  XNOR U17721 ( .A(y[7308]), .B(x[7308]), .Z(n9610) );
  XNOR U17722 ( .A(n9604), .B(n9605), .Z(n9615) );
  XNOR U17723 ( .A(y[7305]), .B(x[7305]), .Z(n9605) );
  XNOR U17724 ( .A(n9606), .B(n9607), .Z(n9604) );
  XNOR U17725 ( .A(y[7306]), .B(x[7306]), .Z(n9607) );
  XNOR U17726 ( .A(y[7307]), .B(x[7307]), .Z(n9606) );
  XNOR U17727 ( .A(n9597), .B(n9596), .Z(n9600) );
  XNOR U17728 ( .A(n9592), .B(n9593), .Z(n9596) );
  XNOR U17729 ( .A(y[7302]), .B(x[7302]), .Z(n9593) );
  XNOR U17730 ( .A(n9594), .B(n9595), .Z(n9592) );
  XNOR U17731 ( .A(y[7303]), .B(x[7303]), .Z(n9595) );
  XNOR U17732 ( .A(y[7304]), .B(x[7304]), .Z(n9594) );
  XNOR U17733 ( .A(n9586), .B(n9587), .Z(n9597) );
  XNOR U17734 ( .A(y[7299]), .B(x[7299]), .Z(n9587) );
  XNOR U17735 ( .A(n9588), .B(n9589), .Z(n9586) );
  XNOR U17736 ( .A(y[7300]), .B(x[7300]), .Z(n9589) );
  XNOR U17737 ( .A(y[7301]), .B(x[7301]), .Z(n9588) );
  XOR U17738 ( .A(n9562), .B(n9563), .Z(n9581) );
  XNOR U17739 ( .A(n9578), .B(n9579), .Z(n9563) );
  XNOR U17740 ( .A(n9573), .B(n9574), .Z(n9579) );
  XNOR U17741 ( .A(n9575), .B(n9576), .Z(n9574) );
  XNOR U17742 ( .A(y[7297]), .B(x[7297]), .Z(n9576) );
  XNOR U17743 ( .A(y[7298]), .B(x[7298]), .Z(n9575) );
  XNOR U17744 ( .A(y[7296]), .B(x[7296]), .Z(n9573) );
  XNOR U17745 ( .A(n9567), .B(n9568), .Z(n9578) );
  XNOR U17746 ( .A(y[7293]), .B(x[7293]), .Z(n9568) );
  XNOR U17747 ( .A(n9569), .B(n9570), .Z(n9567) );
  XNOR U17748 ( .A(y[7294]), .B(x[7294]), .Z(n9570) );
  XNOR U17749 ( .A(y[7295]), .B(x[7295]), .Z(n9569) );
  XOR U17750 ( .A(n9561), .B(n9560), .Z(n9562) );
  XNOR U17751 ( .A(n9556), .B(n9557), .Z(n9560) );
  XNOR U17752 ( .A(y[7290]), .B(x[7290]), .Z(n9557) );
  XNOR U17753 ( .A(n9558), .B(n9559), .Z(n9556) );
  XNOR U17754 ( .A(y[7291]), .B(x[7291]), .Z(n9559) );
  XNOR U17755 ( .A(y[7292]), .B(x[7292]), .Z(n9558) );
  XNOR U17756 ( .A(n9550), .B(n9551), .Z(n9561) );
  XNOR U17757 ( .A(y[7287]), .B(x[7287]), .Z(n9551) );
  XNOR U17758 ( .A(n9552), .B(n9553), .Z(n9550) );
  XNOR U17759 ( .A(y[7288]), .B(x[7288]), .Z(n9553) );
  XNOR U17760 ( .A(y[7289]), .B(x[7289]), .Z(n9552) );
  NAND U17761 ( .A(n9617), .B(n9618), .Z(N64535) );
  NANDN U17762 ( .A(n9619), .B(n9620), .Z(n9618) );
  OR U17763 ( .A(n9621), .B(n9622), .Z(n9620) );
  NAND U17764 ( .A(n9621), .B(n9622), .Z(n9617) );
  XOR U17765 ( .A(n9621), .B(n9623), .Z(N64534) );
  XNOR U17766 ( .A(n9619), .B(n9622), .Z(n9623) );
  AND U17767 ( .A(n9624), .B(n9625), .Z(n9622) );
  NANDN U17768 ( .A(n9626), .B(n9627), .Z(n9625) );
  NANDN U17769 ( .A(n9628), .B(n9629), .Z(n9627) );
  NANDN U17770 ( .A(n9629), .B(n9628), .Z(n9624) );
  NAND U17771 ( .A(n9630), .B(n9631), .Z(n9619) );
  NANDN U17772 ( .A(n9632), .B(n9633), .Z(n9631) );
  OR U17773 ( .A(n9634), .B(n9635), .Z(n9633) );
  NAND U17774 ( .A(n9635), .B(n9634), .Z(n9630) );
  AND U17775 ( .A(n9636), .B(n9637), .Z(n9621) );
  NANDN U17776 ( .A(n9638), .B(n9639), .Z(n9637) );
  NANDN U17777 ( .A(n9640), .B(n9641), .Z(n9639) );
  NANDN U17778 ( .A(n9641), .B(n9640), .Z(n9636) );
  XOR U17779 ( .A(n9635), .B(n9642), .Z(N64533) );
  XOR U17780 ( .A(n9632), .B(n9634), .Z(n9642) );
  XNOR U17781 ( .A(n9628), .B(n9643), .Z(n9634) );
  XNOR U17782 ( .A(n9626), .B(n9629), .Z(n9643) );
  NAND U17783 ( .A(n9644), .B(n9645), .Z(n9629) );
  NAND U17784 ( .A(n9646), .B(n9647), .Z(n9645) );
  OR U17785 ( .A(n9648), .B(n9649), .Z(n9646) );
  NANDN U17786 ( .A(n9650), .B(n9648), .Z(n9644) );
  IV U17787 ( .A(n9649), .Z(n9650) );
  NAND U17788 ( .A(n9651), .B(n9652), .Z(n9626) );
  NAND U17789 ( .A(n9653), .B(n9654), .Z(n9652) );
  NANDN U17790 ( .A(n9655), .B(n9656), .Z(n9653) );
  NANDN U17791 ( .A(n9656), .B(n9655), .Z(n9651) );
  AND U17792 ( .A(n9657), .B(n9658), .Z(n9628) );
  NAND U17793 ( .A(n9659), .B(n9660), .Z(n9658) );
  OR U17794 ( .A(n9661), .B(n9662), .Z(n9659) );
  NANDN U17795 ( .A(n9663), .B(n9661), .Z(n9657) );
  NAND U17796 ( .A(n9664), .B(n9665), .Z(n9632) );
  NANDN U17797 ( .A(n9666), .B(n9667), .Z(n9665) );
  OR U17798 ( .A(n9668), .B(n9669), .Z(n9667) );
  NANDN U17799 ( .A(n9670), .B(n9668), .Z(n9664) );
  IV U17800 ( .A(n9669), .Z(n9670) );
  XNOR U17801 ( .A(n9640), .B(n9671), .Z(n9635) );
  XNOR U17802 ( .A(n9638), .B(n9641), .Z(n9671) );
  NAND U17803 ( .A(n9672), .B(n9673), .Z(n9641) );
  NAND U17804 ( .A(n9674), .B(n9675), .Z(n9673) );
  OR U17805 ( .A(n9676), .B(n9677), .Z(n9674) );
  NANDN U17806 ( .A(n9678), .B(n9676), .Z(n9672) );
  IV U17807 ( .A(n9677), .Z(n9678) );
  NAND U17808 ( .A(n9679), .B(n9680), .Z(n9638) );
  NAND U17809 ( .A(n9681), .B(n9682), .Z(n9680) );
  NANDN U17810 ( .A(n9683), .B(n9684), .Z(n9681) );
  NANDN U17811 ( .A(n9684), .B(n9683), .Z(n9679) );
  AND U17812 ( .A(n9685), .B(n9686), .Z(n9640) );
  NAND U17813 ( .A(n9687), .B(n9688), .Z(n9686) );
  OR U17814 ( .A(n9689), .B(n9690), .Z(n9687) );
  NANDN U17815 ( .A(n9691), .B(n9689), .Z(n9685) );
  XNOR U17816 ( .A(n9666), .B(n9692), .Z(N64532) );
  XOR U17817 ( .A(n9668), .B(n9669), .Z(n9692) );
  XNOR U17818 ( .A(n9682), .B(n9693), .Z(n9669) );
  XOR U17819 ( .A(n9683), .B(n9684), .Z(n9693) );
  XOR U17820 ( .A(n9689), .B(n9694), .Z(n9684) );
  XOR U17821 ( .A(n9688), .B(n9691), .Z(n9694) );
  IV U17822 ( .A(n9690), .Z(n9691) );
  NAND U17823 ( .A(n9695), .B(n9696), .Z(n9690) );
  OR U17824 ( .A(n9697), .B(n9698), .Z(n9696) );
  OR U17825 ( .A(n9699), .B(n9700), .Z(n9695) );
  NAND U17826 ( .A(n9701), .B(n9702), .Z(n9688) );
  OR U17827 ( .A(n9703), .B(n9704), .Z(n9702) );
  OR U17828 ( .A(n9705), .B(n9706), .Z(n9701) );
  NOR U17829 ( .A(n9707), .B(n9708), .Z(n9689) );
  ANDN U17830 ( .B(n9709), .A(n9710), .Z(n9683) );
  XNOR U17831 ( .A(n9676), .B(n9711), .Z(n9682) );
  XNOR U17832 ( .A(n9675), .B(n9677), .Z(n9711) );
  NAND U17833 ( .A(n9712), .B(n9713), .Z(n9677) );
  OR U17834 ( .A(n9714), .B(n9715), .Z(n9713) );
  OR U17835 ( .A(n9716), .B(n9717), .Z(n9712) );
  NAND U17836 ( .A(n9718), .B(n9719), .Z(n9675) );
  OR U17837 ( .A(n9720), .B(n9721), .Z(n9719) );
  OR U17838 ( .A(n9722), .B(n9723), .Z(n9718) );
  ANDN U17839 ( .B(n9724), .A(n9725), .Z(n9676) );
  IV U17840 ( .A(n9726), .Z(n9724) );
  ANDN U17841 ( .B(n9727), .A(n9728), .Z(n9668) );
  XOR U17842 ( .A(n9654), .B(n9729), .Z(n9666) );
  XOR U17843 ( .A(n9655), .B(n9656), .Z(n9729) );
  XOR U17844 ( .A(n9661), .B(n9730), .Z(n9656) );
  XOR U17845 ( .A(n9660), .B(n9663), .Z(n9730) );
  IV U17846 ( .A(n9662), .Z(n9663) );
  NAND U17847 ( .A(n9731), .B(n9732), .Z(n9662) );
  OR U17848 ( .A(n9733), .B(n9734), .Z(n9732) );
  OR U17849 ( .A(n9735), .B(n9736), .Z(n9731) );
  NAND U17850 ( .A(n9737), .B(n9738), .Z(n9660) );
  OR U17851 ( .A(n9739), .B(n9740), .Z(n9738) );
  OR U17852 ( .A(n9741), .B(n9742), .Z(n9737) );
  NOR U17853 ( .A(n9743), .B(n9744), .Z(n9661) );
  ANDN U17854 ( .B(n9745), .A(n9746), .Z(n9655) );
  IV U17855 ( .A(n9747), .Z(n9745) );
  XNOR U17856 ( .A(n9648), .B(n9748), .Z(n9654) );
  XNOR U17857 ( .A(n9647), .B(n9649), .Z(n9748) );
  NAND U17858 ( .A(n9749), .B(n9750), .Z(n9649) );
  OR U17859 ( .A(n9751), .B(n9752), .Z(n9750) );
  OR U17860 ( .A(n9753), .B(n9754), .Z(n9749) );
  NAND U17861 ( .A(n9755), .B(n9756), .Z(n9647) );
  OR U17862 ( .A(n9757), .B(n9758), .Z(n9756) );
  OR U17863 ( .A(n9759), .B(n9760), .Z(n9755) );
  ANDN U17864 ( .B(n9761), .A(n9762), .Z(n9648) );
  IV U17865 ( .A(n9763), .Z(n9761) );
  XNOR U17866 ( .A(n9728), .B(n9727), .Z(N64531) );
  XOR U17867 ( .A(n9747), .B(n9746), .Z(n9727) );
  XNOR U17868 ( .A(n9762), .B(n9763), .Z(n9746) );
  XNOR U17869 ( .A(n9757), .B(n9758), .Z(n9763) );
  XNOR U17870 ( .A(n9759), .B(n9760), .Z(n9758) );
  XNOR U17871 ( .A(y[7285]), .B(x[7285]), .Z(n9760) );
  XNOR U17872 ( .A(y[7286]), .B(x[7286]), .Z(n9759) );
  XNOR U17873 ( .A(y[7284]), .B(x[7284]), .Z(n9757) );
  XNOR U17874 ( .A(n9751), .B(n9752), .Z(n9762) );
  XNOR U17875 ( .A(y[7281]), .B(x[7281]), .Z(n9752) );
  XNOR U17876 ( .A(n9753), .B(n9754), .Z(n9751) );
  XNOR U17877 ( .A(y[7282]), .B(x[7282]), .Z(n9754) );
  XNOR U17878 ( .A(y[7283]), .B(x[7283]), .Z(n9753) );
  XNOR U17879 ( .A(n9744), .B(n9743), .Z(n9747) );
  XNOR U17880 ( .A(n9739), .B(n9740), .Z(n9743) );
  XNOR U17881 ( .A(y[7278]), .B(x[7278]), .Z(n9740) );
  XNOR U17882 ( .A(n9741), .B(n9742), .Z(n9739) );
  XNOR U17883 ( .A(y[7279]), .B(x[7279]), .Z(n9742) );
  XNOR U17884 ( .A(y[7280]), .B(x[7280]), .Z(n9741) );
  XNOR U17885 ( .A(n9733), .B(n9734), .Z(n9744) );
  XNOR U17886 ( .A(y[7275]), .B(x[7275]), .Z(n9734) );
  XNOR U17887 ( .A(n9735), .B(n9736), .Z(n9733) );
  XNOR U17888 ( .A(y[7276]), .B(x[7276]), .Z(n9736) );
  XNOR U17889 ( .A(y[7277]), .B(x[7277]), .Z(n9735) );
  XOR U17890 ( .A(n9709), .B(n9710), .Z(n9728) );
  XNOR U17891 ( .A(n9725), .B(n9726), .Z(n9710) );
  XNOR U17892 ( .A(n9720), .B(n9721), .Z(n9726) );
  XNOR U17893 ( .A(n9722), .B(n9723), .Z(n9721) );
  XNOR U17894 ( .A(y[7273]), .B(x[7273]), .Z(n9723) );
  XNOR U17895 ( .A(y[7274]), .B(x[7274]), .Z(n9722) );
  XNOR U17896 ( .A(y[7272]), .B(x[7272]), .Z(n9720) );
  XNOR U17897 ( .A(n9714), .B(n9715), .Z(n9725) );
  XNOR U17898 ( .A(y[7269]), .B(x[7269]), .Z(n9715) );
  XNOR U17899 ( .A(n9716), .B(n9717), .Z(n9714) );
  XNOR U17900 ( .A(y[7270]), .B(x[7270]), .Z(n9717) );
  XNOR U17901 ( .A(y[7271]), .B(x[7271]), .Z(n9716) );
  XOR U17902 ( .A(n9708), .B(n9707), .Z(n9709) );
  XNOR U17903 ( .A(n9703), .B(n9704), .Z(n9707) );
  XNOR U17904 ( .A(y[7266]), .B(x[7266]), .Z(n9704) );
  XNOR U17905 ( .A(n9705), .B(n9706), .Z(n9703) );
  XNOR U17906 ( .A(y[7267]), .B(x[7267]), .Z(n9706) );
  XNOR U17907 ( .A(y[7268]), .B(x[7268]), .Z(n9705) );
  XNOR U17908 ( .A(n9697), .B(n9698), .Z(n9708) );
  XNOR U17909 ( .A(y[7263]), .B(x[7263]), .Z(n9698) );
  XNOR U17910 ( .A(n9699), .B(n9700), .Z(n9697) );
  XNOR U17911 ( .A(y[7264]), .B(x[7264]), .Z(n9700) );
  XNOR U17912 ( .A(y[7265]), .B(x[7265]), .Z(n9699) );
  NAND U17913 ( .A(n9764), .B(n9765), .Z(N64522) );
  NANDN U17914 ( .A(n9766), .B(n9767), .Z(n9765) );
  OR U17915 ( .A(n9768), .B(n9769), .Z(n9767) );
  NAND U17916 ( .A(n9768), .B(n9769), .Z(n9764) );
  XOR U17917 ( .A(n9768), .B(n9770), .Z(N64521) );
  XNOR U17918 ( .A(n9766), .B(n9769), .Z(n9770) );
  AND U17919 ( .A(n9771), .B(n9772), .Z(n9769) );
  NANDN U17920 ( .A(n9773), .B(n9774), .Z(n9772) );
  NANDN U17921 ( .A(n9775), .B(n9776), .Z(n9774) );
  NANDN U17922 ( .A(n9776), .B(n9775), .Z(n9771) );
  NAND U17923 ( .A(n9777), .B(n9778), .Z(n9766) );
  NANDN U17924 ( .A(n9779), .B(n9780), .Z(n9778) );
  OR U17925 ( .A(n9781), .B(n9782), .Z(n9780) );
  NAND U17926 ( .A(n9782), .B(n9781), .Z(n9777) );
  AND U17927 ( .A(n9783), .B(n9784), .Z(n9768) );
  NANDN U17928 ( .A(n9785), .B(n9786), .Z(n9784) );
  NANDN U17929 ( .A(n9787), .B(n9788), .Z(n9786) );
  NANDN U17930 ( .A(n9788), .B(n9787), .Z(n9783) );
  XOR U17931 ( .A(n9782), .B(n9789), .Z(N64520) );
  XOR U17932 ( .A(n9779), .B(n9781), .Z(n9789) );
  XNOR U17933 ( .A(n9775), .B(n9790), .Z(n9781) );
  XNOR U17934 ( .A(n9773), .B(n9776), .Z(n9790) );
  NAND U17935 ( .A(n9791), .B(n9792), .Z(n9776) );
  NAND U17936 ( .A(n9793), .B(n9794), .Z(n9792) );
  OR U17937 ( .A(n9795), .B(n9796), .Z(n9793) );
  NANDN U17938 ( .A(n9797), .B(n9795), .Z(n9791) );
  IV U17939 ( .A(n9796), .Z(n9797) );
  NAND U17940 ( .A(n9798), .B(n9799), .Z(n9773) );
  NAND U17941 ( .A(n9800), .B(n9801), .Z(n9799) );
  NANDN U17942 ( .A(n9802), .B(n9803), .Z(n9800) );
  NANDN U17943 ( .A(n9803), .B(n9802), .Z(n9798) );
  AND U17944 ( .A(n9804), .B(n9805), .Z(n9775) );
  NAND U17945 ( .A(n9806), .B(n9807), .Z(n9805) );
  OR U17946 ( .A(n9808), .B(n9809), .Z(n9806) );
  NANDN U17947 ( .A(n9810), .B(n9808), .Z(n9804) );
  NAND U17948 ( .A(n9811), .B(n9812), .Z(n9779) );
  NANDN U17949 ( .A(n9813), .B(n9814), .Z(n9812) );
  OR U17950 ( .A(n9815), .B(n9816), .Z(n9814) );
  NANDN U17951 ( .A(n9817), .B(n9815), .Z(n9811) );
  IV U17952 ( .A(n9816), .Z(n9817) );
  XNOR U17953 ( .A(n9787), .B(n9818), .Z(n9782) );
  XNOR U17954 ( .A(n9785), .B(n9788), .Z(n9818) );
  NAND U17955 ( .A(n9819), .B(n9820), .Z(n9788) );
  NAND U17956 ( .A(n9821), .B(n9822), .Z(n9820) );
  OR U17957 ( .A(n9823), .B(n9824), .Z(n9821) );
  NANDN U17958 ( .A(n9825), .B(n9823), .Z(n9819) );
  IV U17959 ( .A(n9824), .Z(n9825) );
  NAND U17960 ( .A(n9826), .B(n9827), .Z(n9785) );
  NAND U17961 ( .A(n9828), .B(n9829), .Z(n9827) );
  NANDN U17962 ( .A(n9830), .B(n9831), .Z(n9828) );
  NANDN U17963 ( .A(n9831), .B(n9830), .Z(n9826) );
  AND U17964 ( .A(n9832), .B(n9833), .Z(n9787) );
  NAND U17965 ( .A(n9834), .B(n9835), .Z(n9833) );
  OR U17966 ( .A(n9836), .B(n9837), .Z(n9834) );
  NANDN U17967 ( .A(n9838), .B(n9836), .Z(n9832) );
  XNOR U17968 ( .A(n9813), .B(n9839), .Z(N64519) );
  XOR U17969 ( .A(n9815), .B(n9816), .Z(n9839) );
  XNOR U17970 ( .A(n9829), .B(n9840), .Z(n9816) );
  XOR U17971 ( .A(n9830), .B(n9831), .Z(n9840) );
  XOR U17972 ( .A(n9836), .B(n9841), .Z(n9831) );
  XOR U17973 ( .A(n9835), .B(n9838), .Z(n9841) );
  IV U17974 ( .A(n9837), .Z(n9838) );
  NAND U17975 ( .A(n9842), .B(n9843), .Z(n9837) );
  OR U17976 ( .A(n9844), .B(n9845), .Z(n9843) );
  OR U17977 ( .A(n9846), .B(n9847), .Z(n9842) );
  NAND U17978 ( .A(n9848), .B(n9849), .Z(n9835) );
  OR U17979 ( .A(n9850), .B(n9851), .Z(n9849) );
  OR U17980 ( .A(n9852), .B(n9853), .Z(n9848) );
  NOR U17981 ( .A(n9854), .B(n9855), .Z(n9836) );
  ANDN U17982 ( .B(n9856), .A(n9857), .Z(n9830) );
  XNOR U17983 ( .A(n9823), .B(n9858), .Z(n9829) );
  XNOR U17984 ( .A(n9822), .B(n9824), .Z(n9858) );
  NAND U17985 ( .A(n9859), .B(n9860), .Z(n9824) );
  OR U17986 ( .A(n9861), .B(n9862), .Z(n9860) );
  OR U17987 ( .A(n9863), .B(n9864), .Z(n9859) );
  NAND U17988 ( .A(n9865), .B(n9866), .Z(n9822) );
  OR U17989 ( .A(n9867), .B(n9868), .Z(n9866) );
  OR U17990 ( .A(n9869), .B(n9870), .Z(n9865) );
  ANDN U17991 ( .B(n9871), .A(n9872), .Z(n9823) );
  IV U17992 ( .A(n9873), .Z(n9871) );
  ANDN U17993 ( .B(n9874), .A(n9875), .Z(n9815) );
  XOR U17994 ( .A(n9801), .B(n9876), .Z(n9813) );
  XOR U17995 ( .A(n9802), .B(n9803), .Z(n9876) );
  XOR U17996 ( .A(n9808), .B(n9877), .Z(n9803) );
  XOR U17997 ( .A(n9807), .B(n9810), .Z(n9877) );
  IV U17998 ( .A(n9809), .Z(n9810) );
  NAND U17999 ( .A(n9878), .B(n9879), .Z(n9809) );
  OR U18000 ( .A(n9880), .B(n9881), .Z(n9879) );
  OR U18001 ( .A(n9882), .B(n9883), .Z(n9878) );
  NAND U18002 ( .A(n9884), .B(n9885), .Z(n9807) );
  OR U18003 ( .A(n9886), .B(n9887), .Z(n9885) );
  OR U18004 ( .A(n9888), .B(n9889), .Z(n9884) );
  NOR U18005 ( .A(n9890), .B(n9891), .Z(n9808) );
  ANDN U18006 ( .B(n9892), .A(n9893), .Z(n9802) );
  IV U18007 ( .A(n9894), .Z(n9892) );
  XNOR U18008 ( .A(n9795), .B(n9895), .Z(n9801) );
  XNOR U18009 ( .A(n9794), .B(n9796), .Z(n9895) );
  NAND U18010 ( .A(n9896), .B(n9897), .Z(n9796) );
  OR U18011 ( .A(n9898), .B(n9899), .Z(n9897) );
  OR U18012 ( .A(n9900), .B(n9901), .Z(n9896) );
  NAND U18013 ( .A(n9902), .B(n9903), .Z(n9794) );
  OR U18014 ( .A(n9904), .B(n9905), .Z(n9903) );
  OR U18015 ( .A(n9906), .B(n9907), .Z(n9902) );
  ANDN U18016 ( .B(n9908), .A(n9909), .Z(n9795) );
  IV U18017 ( .A(n9910), .Z(n9908) );
  XNOR U18018 ( .A(n9875), .B(n9874), .Z(N64518) );
  XOR U18019 ( .A(n9894), .B(n9893), .Z(n9874) );
  XNOR U18020 ( .A(n9909), .B(n9910), .Z(n9893) );
  XNOR U18021 ( .A(n9904), .B(n9905), .Z(n9910) );
  XNOR U18022 ( .A(n9906), .B(n9907), .Z(n9905) );
  XNOR U18023 ( .A(y[7261]), .B(x[7261]), .Z(n9907) );
  XNOR U18024 ( .A(y[7262]), .B(x[7262]), .Z(n9906) );
  XNOR U18025 ( .A(y[7260]), .B(x[7260]), .Z(n9904) );
  XNOR U18026 ( .A(n9898), .B(n9899), .Z(n9909) );
  XNOR U18027 ( .A(y[7257]), .B(x[7257]), .Z(n9899) );
  XNOR U18028 ( .A(n9900), .B(n9901), .Z(n9898) );
  XNOR U18029 ( .A(y[7258]), .B(x[7258]), .Z(n9901) );
  XNOR U18030 ( .A(y[7259]), .B(x[7259]), .Z(n9900) );
  XNOR U18031 ( .A(n9891), .B(n9890), .Z(n9894) );
  XNOR U18032 ( .A(n9886), .B(n9887), .Z(n9890) );
  XNOR U18033 ( .A(y[7254]), .B(x[7254]), .Z(n9887) );
  XNOR U18034 ( .A(n9888), .B(n9889), .Z(n9886) );
  XNOR U18035 ( .A(y[7255]), .B(x[7255]), .Z(n9889) );
  XNOR U18036 ( .A(y[7256]), .B(x[7256]), .Z(n9888) );
  XNOR U18037 ( .A(n9880), .B(n9881), .Z(n9891) );
  XNOR U18038 ( .A(y[7251]), .B(x[7251]), .Z(n9881) );
  XNOR U18039 ( .A(n9882), .B(n9883), .Z(n9880) );
  XNOR U18040 ( .A(y[7252]), .B(x[7252]), .Z(n9883) );
  XNOR U18041 ( .A(y[7253]), .B(x[7253]), .Z(n9882) );
  XOR U18042 ( .A(n9856), .B(n9857), .Z(n9875) );
  XNOR U18043 ( .A(n9872), .B(n9873), .Z(n9857) );
  XNOR U18044 ( .A(n9867), .B(n9868), .Z(n9873) );
  XNOR U18045 ( .A(n9869), .B(n9870), .Z(n9868) );
  XNOR U18046 ( .A(y[7249]), .B(x[7249]), .Z(n9870) );
  XNOR U18047 ( .A(y[7250]), .B(x[7250]), .Z(n9869) );
  XNOR U18048 ( .A(y[7248]), .B(x[7248]), .Z(n9867) );
  XNOR U18049 ( .A(n9861), .B(n9862), .Z(n9872) );
  XNOR U18050 ( .A(y[7245]), .B(x[7245]), .Z(n9862) );
  XNOR U18051 ( .A(n9863), .B(n9864), .Z(n9861) );
  XNOR U18052 ( .A(y[7246]), .B(x[7246]), .Z(n9864) );
  XNOR U18053 ( .A(y[7247]), .B(x[7247]), .Z(n9863) );
  XOR U18054 ( .A(n9855), .B(n9854), .Z(n9856) );
  XNOR U18055 ( .A(n9850), .B(n9851), .Z(n9854) );
  XNOR U18056 ( .A(y[7242]), .B(x[7242]), .Z(n9851) );
  XNOR U18057 ( .A(n9852), .B(n9853), .Z(n9850) );
  XNOR U18058 ( .A(y[7243]), .B(x[7243]), .Z(n9853) );
  XNOR U18059 ( .A(y[7244]), .B(x[7244]), .Z(n9852) );
  XNOR U18060 ( .A(n9844), .B(n9845), .Z(n9855) );
  XNOR U18061 ( .A(y[7239]), .B(x[7239]), .Z(n9845) );
  XNOR U18062 ( .A(n9846), .B(n9847), .Z(n9844) );
  XNOR U18063 ( .A(y[7240]), .B(x[7240]), .Z(n9847) );
  XNOR U18064 ( .A(y[7241]), .B(x[7241]), .Z(n9846) );
  NAND U18065 ( .A(n9911), .B(n9912), .Z(N64509) );
  NANDN U18066 ( .A(n9913), .B(n9914), .Z(n9912) );
  OR U18067 ( .A(n9915), .B(n9916), .Z(n9914) );
  NAND U18068 ( .A(n9915), .B(n9916), .Z(n9911) );
  XOR U18069 ( .A(n9915), .B(n9917), .Z(N64508) );
  XNOR U18070 ( .A(n9913), .B(n9916), .Z(n9917) );
  AND U18071 ( .A(n9918), .B(n9919), .Z(n9916) );
  NANDN U18072 ( .A(n9920), .B(n9921), .Z(n9919) );
  NANDN U18073 ( .A(n9922), .B(n9923), .Z(n9921) );
  NANDN U18074 ( .A(n9923), .B(n9922), .Z(n9918) );
  NAND U18075 ( .A(n9924), .B(n9925), .Z(n9913) );
  NANDN U18076 ( .A(n9926), .B(n9927), .Z(n9925) );
  OR U18077 ( .A(n9928), .B(n9929), .Z(n9927) );
  NAND U18078 ( .A(n9929), .B(n9928), .Z(n9924) );
  AND U18079 ( .A(n9930), .B(n9931), .Z(n9915) );
  NANDN U18080 ( .A(n9932), .B(n9933), .Z(n9931) );
  NANDN U18081 ( .A(n9934), .B(n9935), .Z(n9933) );
  NANDN U18082 ( .A(n9935), .B(n9934), .Z(n9930) );
  XOR U18083 ( .A(n9929), .B(n9936), .Z(N64507) );
  XOR U18084 ( .A(n9926), .B(n9928), .Z(n9936) );
  XNOR U18085 ( .A(n9922), .B(n9937), .Z(n9928) );
  XNOR U18086 ( .A(n9920), .B(n9923), .Z(n9937) );
  NAND U18087 ( .A(n9938), .B(n9939), .Z(n9923) );
  NAND U18088 ( .A(n9940), .B(n9941), .Z(n9939) );
  OR U18089 ( .A(n9942), .B(n9943), .Z(n9940) );
  NANDN U18090 ( .A(n9944), .B(n9942), .Z(n9938) );
  IV U18091 ( .A(n9943), .Z(n9944) );
  NAND U18092 ( .A(n9945), .B(n9946), .Z(n9920) );
  NAND U18093 ( .A(n9947), .B(n9948), .Z(n9946) );
  NANDN U18094 ( .A(n9949), .B(n9950), .Z(n9947) );
  NANDN U18095 ( .A(n9950), .B(n9949), .Z(n9945) );
  AND U18096 ( .A(n9951), .B(n9952), .Z(n9922) );
  NAND U18097 ( .A(n9953), .B(n9954), .Z(n9952) );
  OR U18098 ( .A(n9955), .B(n9956), .Z(n9953) );
  NANDN U18099 ( .A(n9957), .B(n9955), .Z(n9951) );
  NAND U18100 ( .A(n9958), .B(n9959), .Z(n9926) );
  NANDN U18101 ( .A(n9960), .B(n9961), .Z(n9959) );
  OR U18102 ( .A(n9962), .B(n9963), .Z(n9961) );
  NANDN U18103 ( .A(n9964), .B(n9962), .Z(n9958) );
  IV U18104 ( .A(n9963), .Z(n9964) );
  XNOR U18105 ( .A(n9934), .B(n9965), .Z(n9929) );
  XNOR U18106 ( .A(n9932), .B(n9935), .Z(n9965) );
  NAND U18107 ( .A(n9966), .B(n9967), .Z(n9935) );
  NAND U18108 ( .A(n9968), .B(n9969), .Z(n9967) );
  OR U18109 ( .A(n9970), .B(n9971), .Z(n9968) );
  NANDN U18110 ( .A(n9972), .B(n9970), .Z(n9966) );
  IV U18111 ( .A(n9971), .Z(n9972) );
  NAND U18112 ( .A(n9973), .B(n9974), .Z(n9932) );
  NAND U18113 ( .A(n9975), .B(n9976), .Z(n9974) );
  NANDN U18114 ( .A(n9977), .B(n9978), .Z(n9975) );
  NANDN U18115 ( .A(n9978), .B(n9977), .Z(n9973) );
  AND U18116 ( .A(n9979), .B(n9980), .Z(n9934) );
  NAND U18117 ( .A(n9981), .B(n9982), .Z(n9980) );
  OR U18118 ( .A(n9983), .B(n9984), .Z(n9981) );
  NANDN U18119 ( .A(n9985), .B(n9983), .Z(n9979) );
  XNOR U18120 ( .A(n9960), .B(n9986), .Z(N64506) );
  XOR U18121 ( .A(n9962), .B(n9963), .Z(n9986) );
  XNOR U18122 ( .A(n9976), .B(n9987), .Z(n9963) );
  XOR U18123 ( .A(n9977), .B(n9978), .Z(n9987) );
  XOR U18124 ( .A(n9983), .B(n9988), .Z(n9978) );
  XOR U18125 ( .A(n9982), .B(n9985), .Z(n9988) );
  IV U18126 ( .A(n9984), .Z(n9985) );
  NAND U18127 ( .A(n9989), .B(n9990), .Z(n9984) );
  OR U18128 ( .A(n9991), .B(n9992), .Z(n9990) );
  OR U18129 ( .A(n9993), .B(n9994), .Z(n9989) );
  NAND U18130 ( .A(n9995), .B(n9996), .Z(n9982) );
  OR U18131 ( .A(n9997), .B(n9998), .Z(n9996) );
  OR U18132 ( .A(n9999), .B(n10000), .Z(n9995) );
  NOR U18133 ( .A(n10001), .B(n10002), .Z(n9983) );
  ANDN U18134 ( .B(n10003), .A(n10004), .Z(n9977) );
  XNOR U18135 ( .A(n9970), .B(n10005), .Z(n9976) );
  XNOR U18136 ( .A(n9969), .B(n9971), .Z(n10005) );
  NAND U18137 ( .A(n10006), .B(n10007), .Z(n9971) );
  OR U18138 ( .A(n10008), .B(n10009), .Z(n10007) );
  OR U18139 ( .A(n10010), .B(n10011), .Z(n10006) );
  NAND U18140 ( .A(n10012), .B(n10013), .Z(n9969) );
  OR U18141 ( .A(n10014), .B(n10015), .Z(n10013) );
  OR U18142 ( .A(n10016), .B(n10017), .Z(n10012) );
  ANDN U18143 ( .B(n10018), .A(n10019), .Z(n9970) );
  IV U18144 ( .A(n10020), .Z(n10018) );
  ANDN U18145 ( .B(n10021), .A(n10022), .Z(n9962) );
  XOR U18146 ( .A(n9948), .B(n10023), .Z(n9960) );
  XOR U18147 ( .A(n9949), .B(n9950), .Z(n10023) );
  XOR U18148 ( .A(n9955), .B(n10024), .Z(n9950) );
  XOR U18149 ( .A(n9954), .B(n9957), .Z(n10024) );
  IV U18150 ( .A(n9956), .Z(n9957) );
  NAND U18151 ( .A(n10025), .B(n10026), .Z(n9956) );
  OR U18152 ( .A(n10027), .B(n10028), .Z(n10026) );
  OR U18153 ( .A(n10029), .B(n10030), .Z(n10025) );
  NAND U18154 ( .A(n10031), .B(n10032), .Z(n9954) );
  OR U18155 ( .A(n10033), .B(n10034), .Z(n10032) );
  OR U18156 ( .A(n10035), .B(n10036), .Z(n10031) );
  NOR U18157 ( .A(n10037), .B(n10038), .Z(n9955) );
  ANDN U18158 ( .B(n10039), .A(n10040), .Z(n9949) );
  IV U18159 ( .A(n10041), .Z(n10039) );
  XNOR U18160 ( .A(n9942), .B(n10042), .Z(n9948) );
  XNOR U18161 ( .A(n9941), .B(n9943), .Z(n10042) );
  NAND U18162 ( .A(n10043), .B(n10044), .Z(n9943) );
  OR U18163 ( .A(n10045), .B(n10046), .Z(n10044) );
  OR U18164 ( .A(n10047), .B(n10048), .Z(n10043) );
  NAND U18165 ( .A(n10049), .B(n10050), .Z(n9941) );
  OR U18166 ( .A(n10051), .B(n10052), .Z(n10050) );
  OR U18167 ( .A(n10053), .B(n10054), .Z(n10049) );
  ANDN U18168 ( .B(n10055), .A(n10056), .Z(n9942) );
  IV U18169 ( .A(n10057), .Z(n10055) );
  XNOR U18170 ( .A(n10022), .B(n10021), .Z(N64505) );
  XOR U18171 ( .A(n10041), .B(n10040), .Z(n10021) );
  XNOR U18172 ( .A(n10056), .B(n10057), .Z(n10040) );
  XNOR U18173 ( .A(n10051), .B(n10052), .Z(n10057) );
  XNOR U18174 ( .A(n10053), .B(n10054), .Z(n10052) );
  XNOR U18175 ( .A(y[7237]), .B(x[7237]), .Z(n10054) );
  XNOR U18176 ( .A(y[7238]), .B(x[7238]), .Z(n10053) );
  XNOR U18177 ( .A(y[7236]), .B(x[7236]), .Z(n10051) );
  XNOR U18178 ( .A(n10045), .B(n10046), .Z(n10056) );
  XNOR U18179 ( .A(y[7233]), .B(x[7233]), .Z(n10046) );
  XNOR U18180 ( .A(n10047), .B(n10048), .Z(n10045) );
  XNOR U18181 ( .A(y[7234]), .B(x[7234]), .Z(n10048) );
  XNOR U18182 ( .A(y[7235]), .B(x[7235]), .Z(n10047) );
  XNOR U18183 ( .A(n10038), .B(n10037), .Z(n10041) );
  XNOR U18184 ( .A(n10033), .B(n10034), .Z(n10037) );
  XNOR U18185 ( .A(y[7230]), .B(x[7230]), .Z(n10034) );
  XNOR U18186 ( .A(n10035), .B(n10036), .Z(n10033) );
  XNOR U18187 ( .A(y[7231]), .B(x[7231]), .Z(n10036) );
  XNOR U18188 ( .A(y[7232]), .B(x[7232]), .Z(n10035) );
  XNOR U18189 ( .A(n10027), .B(n10028), .Z(n10038) );
  XNOR U18190 ( .A(y[7227]), .B(x[7227]), .Z(n10028) );
  XNOR U18191 ( .A(n10029), .B(n10030), .Z(n10027) );
  XNOR U18192 ( .A(y[7228]), .B(x[7228]), .Z(n10030) );
  XNOR U18193 ( .A(y[7229]), .B(x[7229]), .Z(n10029) );
  XOR U18194 ( .A(n10003), .B(n10004), .Z(n10022) );
  XNOR U18195 ( .A(n10019), .B(n10020), .Z(n10004) );
  XNOR U18196 ( .A(n10014), .B(n10015), .Z(n10020) );
  XNOR U18197 ( .A(n10016), .B(n10017), .Z(n10015) );
  XNOR U18198 ( .A(y[7225]), .B(x[7225]), .Z(n10017) );
  XNOR U18199 ( .A(y[7226]), .B(x[7226]), .Z(n10016) );
  XNOR U18200 ( .A(y[7224]), .B(x[7224]), .Z(n10014) );
  XNOR U18201 ( .A(n10008), .B(n10009), .Z(n10019) );
  XNOR U18202 ( .A(y[7221]), .B(x[7221]), .Z(n10009) );
  XNOR U18203 ( .A(n10010), .B(n10011), .Z(n10008) );
  XNOR U18204 ( .A(y[7222]), .B(x[7222]), .Z(n10011) );
  XNOR U18205 ( .A(y[7223]), .B(x[7223]), .Z(n10010) );
  XOR U18206 ( .A(n10002), .B(n10001), .Z(n10003) );
  XNOR U18207 ( .A(n9997), .B(n9998), .Z(n10001) );
  XNOR U18208 ( .A(y[7218]), .B(x[7218]), .Z(n9998) );
  XNOR U18209 ( .A(n9999), .B(n10000), .Z(n9997) );
  XNOR U18210 ( .A(y[7219]), .B(x[7219]), .Z(n10000) );
  XNOR U18211 ( .A(y[7220]), .B(x[7220]), .Z(n9999) );
  XNOR U18212 ( .A(n9991), .B(n9992), .Z(n10002) );
  XNOR U18213 ( .A(y[7215]), .B(x[7215]), .Z(n9992) );
  XNOR U18214 ( .A(n9993), .B(n9994), .Z(n9991) );
  XNOR U18215 ( .A(y[7216]), .B(x[7216]), .Z(n9994) );
  XNOR U18216 ( .A(y[7217]), .B(x[7217]), .Z(n9993) );
  NAND U18217 ( .A(n10058), .B(n10059), .Z(N64496) );
  NANDN U18218 ( .A(n10060), .B(n10061), .Z(n10059) );
  OR U18219 ( .A(n10062), .B(n10063), .Z(n10061) );
  NAND U18220 ( .A(n10062), .B(n10063), .Z(n10058) );
  XOR U18221 ( .A(n10062), .B(n10064), .Z(N64495) );
  XNOR U18222 ( .A(n10060), .B(n10063), .Z(n10064) );
  AND U18223 ( .A(n10065), .B(n10066), .Z(n10063) );
  NANDN U18224 ( .A(n10067), .B(n10068), .Z(n10066) );
  NANDN U18225 ( .A(n10069), .B(n10070), .Z(n10068) );
  NANDN U18226 ( .A(n10070), .B(n10069), .Z(n10065) );
  NAND U18227 ( .A(n10071), .B(n10072), .Z(n10060) );
  NANDN U18228 ( .A(n10073), .B(n10074), .Z(n10072) );
  OR U18229 ( .A(n10075), .B(n10076), .Z(n10074) );
  NAND U18230 ( .A(n10076), .B(n10075), .Z(n10071) );
  AND U18231 ( .A(n10077), .B(n10078), .Z(n10062) );
  NANDN U18232 ( .A(n10079), .B(n10080), .Z(n10078) );
  NANDN U18233 ( .A(n10081), .B(n10082), .Z(n10080) );
  NANDN U18234 ( .A(n10082), .B(n10081), .Z(n10077) );
  XOR U18235 ( .A(n10076), .B(n10083), .Z(N64494) );
  XOR U18236 ( .A(n10073), .B(n10075), .Z(n10083) );
  XNOR U18237 ( .A(n10069), .B(n10084), .Z(n10075) );
  XNOR U18238 ( .A(n10067), .B(n10070), .Z(n10084) );
  NAND U18239 ( .A(n10085), .B(n10086), .Z(n10070) );
  NAND U18240 ( .A(n10087), .B(n10088), .Z(n10086) );
  OR U18241 ( .A(n10089), .B(n10090), .Z(n10087) );
  NANDN U18242 ( .A(n10091), .B(n10089), .Z(n10085) );
  IV U18243 ( .A(n10090), .Z(n10091) );
  NAND U18244 ( .A(n10092), .B(n10093), .Z(n10067) );
  NAND U18245 ( .A(n10094), .B(n10095), .Z(n10093) );
  NANDN U18246 ( .A(n10096), .B(n10097), .Z(n10094) );
  NANDN U18247 ( .A(n10097), .B(n10096), .Z(n10092) );
  AND U18248 ( .A(n10098), .B(n10099), .Z(n10069) );
  NAND U18249 ( .A(n10100), .B(n10101), .Z(n10099) );
  OR U18250 ( .A(n10102), .B(n10103), .Z(n10100) );
  NANDN U18251 ( .A(n10104), .B(n10102), .Z(n10098) );
  NAND U18252 ( .A(n10105), .B(n10106), .Z(n10073) );
  NANDN U18253 ( .A(n10107), .B(n10108), .Z(n10106) );
  OR U18254 ( .A(n10109), .B(n10110), .Z(n10108) );
  NANDN U18255 ( .A(n10111), .B(n10109), .Z(n10105) );
  IV U18256 ( .A(n10110), .Z(n10111) );
  XNOR U18257 ( .A(n10081), .B(n10112), .Z(n10076) );
  XNOR U18258 ( .A(n10079), .B(n10082), .Z(n10112) );
  NAND U18259 ( .A(n10113), .B(n10114), .Z(n10082) );
  NAND U18260 ( .A(n10115), .B(n10116), .Z(n10114) );
  OR U18261 ( .A(n10117), .B(n10118), .Z(n10115) );
  NANDN U18262 ( .A(n10119), .B(n10117), .Z(n10113) );
  IV U18263 ( .A(n10118), .Z(n10119) );
  NAND U18264 ( .A(n10120), .B(n10121), .Z(n10079) );
  NAND U18265 ( .A(n10122), .B(n10123), .Z(n10121) );
  NANDN U18266 ( .A(n10124), .B(n10125), .Z(n10122) );
  NANDN U18267 ( .A(n10125), .B(n10124), .Z(n10120) );
  AND U18268 ( .A(n10126), .B(n10127), .Z(n10081) );
  NAND U18269 ( .A(n10128), .B(n10129), .Z(n10127) );
  OR U18270 ( .A(n10130), .B(n10131), .Z(n10128) );
  NANDN U18271 ( .A(n10132), .B(n10130), .Z(n10126) );
  XNOR U18272 ( .A(n10107), .B(n10133), .Z(N64493) );
  XOR U18273 ( .A(n10109), .B(n10110), .Z(n10133) );
  XNOR U18274 ( .A(n10123), .B(n10134), .Z(n10110) );
  XOR U18275 ( .A(n10124), .B(n10125), .Z(n10134) );
  XOR U18276 ( .A(n10130), .B(n10135), .Z(n10125) );
  XOR U18277 ( .A(n10129), .B(n10132), .Z(n10135) );
  IV U18278 ( .A(n10131), .Z(n10132) );
  NAND U18279 ( .A(n10136), .B(n10137), .Z(n10131) );
  OR U18280 ( .A(n10138), .B(n10139), .Z(n10137) );
  OR U18281 ( .A(n10140), .B(n10141), .Z(n10136) );
  NAND U18282 ( .A(n10142), .B(n10143), .Z(n10129) );
  OR U18283 ( .A(n10144), .B(n10145), .Z(n10143) );
  OR U18284 ( .A(n10146), .B(n10147), .Z(n10142) );
  NOR U18285 ( .A(n10148), .B(n10149), .Z(n10130) );
  ANDN U18286 ( .B(n10150), .A(n10151), .Z(n10124) );
  XNOR U18287 ( .A(n10117), .B(n10152), .Z(n10123) );
  XNOR U18288 ( .A(n10116), .B(n10118), .Z(n10152) );
  NAND U18289 ( .A(n10153), .B(n10154), .Z(n10118) );
  OR U18290 ( .A(n10155), .B(n10156), .Z(n10154) );
  OR U18291 ( .A(n10157), .B(n10158), .Z(n10153) );
  NAND U18292 ( .A(n10159), .B(n10160), .Z(n10116) );
  OR U18293 ( .A(n10161), .B(n10162), .Z(n10160) );
  OR U18294 ( .A(n10163), .B(n10164), .Z(n10159) );
  ANDN U18295 ( .B(n10165), .A(n10166), .Z(n10117) );
  IV U18296 ( .A(n10167), .Z(n10165) );
  ANDN U18297 ( .B(n10168), .A(n10169), .Z(n10109) );
  XOR U18298 ( .A(n10095), .B(n10170), .Z(n10107) );
  XOR U18299 ( .A(n10096), .B(n10097), .Z(n10170) );
  XOR U18300 ( .A(n10102), .B(n10171), .Z(n10097) );
  XOR U18301 ( .A(n10101), .B(n10104), .Z(n10171) );
  IV U18302 ( .A(n10103), .Z(n10104) );
  NAND U18303 ( .A(n10172), .B(n10173), .Z(n10103) );
  OR U18304 ( .A(n10174), .B(n10175), .Z(n10173) );
  OR U18305 ( .A(n10176), .B(n10177), .Z(n10172) );
  NAND U18306 ( .A(n10178), .B(n10179), .Z(n10101) );
  OR U18307 ( .A(n10180), .B(n10181), .Z(n10179) );
  OR U18308 ( .A(n10182), .B(n10183), .Z(n10178) );
  NOR U18309 ( .A(n10184), .B(n10185), .Z(n10102) );
  ANDN U18310 ( .B(n10186), .A(n10187), .Z(n10096) );
  IV U18311 ( .A(n10188), .Z(n10186) );
  XNOR U18312 ( .A(n10089), .B(n10189), .Z(n10095) );
  XNOR U18313 ( .A(n10088), .B(n10090), .Z(n10189) );
  NAND U18314 ( .A(n10190), .B(n10191), .Z(n10090) );
  OR U18315 ( .A(n10192), .B(n10193), .Z(n10191) );
  OR U18316 ( .A(n10194), .B(n10195), .Z(n10190) );
  NAND U18317 ( .A(n10196), .B(n10197), .Z(n10088) );
  OR U18318 ( .A(n10198), .B(n10199), .Z(n10197) );
  OR U18319 ( .A(n10200), .B(n10201), .Z(n10196) );
  ANDN U18320 ( .B(n10202), .A(n10203), .Z(n10089) );
  IV U18321 ( .A(n10204), .Z(n10202) );
  XNOR U18322 ( .A(n10169), .B(n10168), .Z(N64492) );
  XOR U18323 ( .A(n10188), .B(n10187), .Z(n10168) );
  XNOR U18324 ( .A(n10203), .B(n10204), .Z(n10187) );
  XNOR U18325 ( .A(n10198), .B(n10199), .Z(n10204) );
  XNOR U18326 ( .A(n10200), .B(n10201), .Z(n10199) );
  XNOR U18327 ( .A(y[7213]), .B(x[7213]), .Z(n10201) );
  XNOR U18328 ( .A(y[7214]), .B(x[7214]), .Z(n10200) );
  XNOR U18329 ( .A(y[7212]), .B(x[7212]), .Z(n10198) );
  XNOR U18330 ( .A(n10192), .B(n10193), .Z(n10203) );
  XNOR U18331 ( .A(y[7209]), .B(x[7209]), .Z(n10193) );
  XNOR U18332 ( .A(n10194), .B(n10195), .Z(n10192) );
  XNOR U18333 ( .A(y[7210]), .B(x[7210]), .Z(n10195) );
  XNOR U18334 ( .A(y[7211]), .B(x[7211]), .Z(n10194) );
  XNOR U18335 ( .A(n10185), .B(n10184), .Z(n10188) );
  XNOR U18336 ( .A(n10180), .B(n10181), .Z(n10184) );
  XNOR U18337 ( .A(y[7206]), .B(x[7206]), .Z(n10181) );
  XNOR U18338 ( .A(n10182), .B(n10183), .Z(n10180) );
  XNOR U18339 ( .A(y[7207]), .B(x[7207]), .Z(n10183) );
  XNOR U18340 ( .A(y[7208]), .B(x[7208]), .Z(n10182) );
  XNOR U18341 ( .A(n10174), .B(n10175), .Z(n10185) );
  XNOR U18342 ( .A(y[7203]), .B(x[7203]), .Z(n10175) );
  XNOR U18343 ( .A(n10176), .B(n10177), .Z(n10174) );
  XNOR U18344 ( .A(y[7204]), .B(x[7204]), .Z(n10177) );
  XNOR U18345 ( .A(y[7205]), .B(x[7205]), .Z(n10176) );
  XOR U18346 ( .A(n10150), .B(n10151), .Z(n10169) );
  XNOR U18347 ( .A(n10166), .B(n10167), .Z(n10151) );
  XNOR U18348 ( .A(n10161), .B(n10162), .Z(n10167) );
  XNOR U18349 ( .A(n10163), .B(n10164), .Z(n10162) );
  XNOR U18350 ( .A(y[7201]), .B(x[7201]), .Z(n10164) );
  XNOR U18351 ( .A(y[7202]), .B(x[7202]), .Z(n10163) );
  XNOR U18352 ( .A(y[7200]), .B(x[7200]), .Z(n10161) );
  XNOR U18353 ( .A(n10155), .B(n10156), .Z(n10166) );
  XNOR U18354 ( .A(y[7197]), .B(x[7197]), .Z(n10156) );
  XNOR U18355 ( .A(n10157), .B(n10158), .Z(n10155) );
  XNOR U18356 ( .A(y[7198]), .B(x[7198]), .Z(n10158) );
  XNOR U18357 ( .A(y[7199]), .B(x[7199]), .Z(n10157) );
  XOR U18358 ( .A(n10149), .B(n10148), .Z(n10150) );
  XNOR U18359 ( .A(n10144), .B(n10145), .Z(n10148) );
  XNOR U18360 ( .A(y[7194]), .B(x[7194]), .Z(n10145) );
  XNOR U18361 ( .A(n10146), .B(n10147), .Z(n10144) );
  XNOR U18362 ( .A(y[7195]), .B(x[7195]), .Z(n10147) );
  XNOR U18363 ( .A(y[7196]), .B(x[7196]), .Z(n10146) );
  XNOR U18364 ( .A(n10138), .B(n10139), .Z(n10149) );
  XNOR U18365 ( .A(y[7191]), .B(x[7191]), .Z(n10139) );
  XNOR U18366 ( .A(n10140), .B(n10141), .Z(n10138) );
  XNOR U18367 ( .A(y[7192]), .B(x[7192]), .Z(n10141) );
  XNOR U18368 ( .A(y[7193]), .B(x[7193]), .Z(n10140) );
  NAND U18369 ( .A(n10205), .B(n10206), .Z(N64483) );
  NANDN U18370 ( .A(n10207), .B(n10208), .Z(n10206) );
  OR U18371 ( .A(n10209), .B(n10210), .Z(n10208) );
  NAND U18372 ( .A(n10209), .B(n10210), .Z(n10205) );
  XOR U18373 ( .A(n10209), .B(n10211), .Z(N64482) );
  XNOR U18374 ( .A(n10207), .B(n10210), .Z(n10211) );
  AND U18375 ( .A(n10212), .B(n10213), .Z(n10210) );
  NANDN U18376 ( .A(n10214), .B(n10215), .Z(n10213) );
  NANDN U18377 ( .A(n10216), .B(n10217), .Z(n10215) );
  NANDN U18378 ( .A(n10217), .B(n10216), .Z(n10212) );
  NAND U18379 ( .A(n10218), .B(n10219), .Z(n10207) );
  NANDN U18380 ( .A(n10220), .B(n10221), .Z(n10219) );
  OR U18381 ( .A(n10222), .B(n10223), .Z(n10221) );
  NAND U18382 ( .A(n10223), .B(n10222), .Z(n10218) );
  AND U18383 ( .A(n10224), .B(n10225), .Z(n10209) );
  NANDN U18384 ( .A(n10226), .B(n10227), .Z(n10225) );
  NANDN U18385 ( .A(n10228), .B(n10229), .Z(n10227) );
  NANDN U18386 ( .A(n10229), .B(n10228), .Z(n10224) );
  XOR U18387 ( .A(n10223), .B(n10230), .Z(N64481) );
  XOR U18388 ( .A(n10220), .B(n10222), .Z(n10230) );
  XNOR U18389 ( .A(n10216), .B(n10231), .Z(n10222) );
  XNOR U18390 ( .A(n10214), .B(n10217), .Z(n10231) );
  NAND U18391 ( .A(n10232), .B(n10233), .Z(n10217) );
  NAND U18392 ( .A(n10234), .B(n10235), .Z(n10233) );
  OR U18393 ( .A(n10236), .B(n10237), .Z(n10234) );
  NANDN U18394 ( .A(n10238), .B(n10236), .Z(n10232) );
  IV U18395 ( .A(n10237), .Z(n10238) );
  NAND U18396 ( .A(n10239), .B(n10240), .Z(n10214) );
  NAND U18397 ( .A(n10241), .B(n10242), .Z(n10240) );
  NANDN U18398 ( .A(n10243), .B(n10244), .Z(n10241) );
  NANDN U18399 ( .A(n10244), .B(n10243), .Z(n10239) );
  AND U18400 ( .A(n10245), .B(n10246), .Z(n10216) );
  NAND U18401 ( .A(n10247), .B(n10248), .Z(n10246) );
  OR U18402 ( .A(n10249), .B(n10250), .Z(n10247) );
  NANDN U18403 ( .A(n10251), .B(n10249), .Z(n10245) );
  NAND U18404 ( .A(n10252), .B(n10253), .Z(n10220) );
  NANDN U18405 ( .A(n10254), .B(n10255), .Z(n10253) );
  OR U18406 ( .A(n10256), .B(n10257), .Z(n10255) );
  NANDN U18407 ( .A(n10258), .B(n10256), .Z(n10252) );
  IV U18408 ( .A(n10257), .Z(n10258) );
  XNOR U18409 ( .A(n10228), .B(n10259), .Z(n10223) );
  XNOR U18410 ( .A(n10226), .B(n10229), .Z(n10259) );
  NAND U18411 ( .A(n10260), .B(n10261), .Z(n10229) );
  NAND U18412 ( .A(n10262), .B(n10263), .Z(n10261) );
  OR U18413 ( .A(n10264), .B(n10265), .Z(n10262) );
  NANDN U18414 ( .A(n10266), .B(n10264), .Z(n10260) );
  IV U18415 ( .A(n10265), .Z(n10266) );
  NAND U18416 ( .A(n10267), .B(n10268), .Z(n10226) );
  NAND U18417 ( .A(n10269), .B(n10270), .Z(n10268) );
  NANDN U18418 ( .A(n10271), .B(n10272), .Z(n10269) );
  NANDN U18419 ( .A(n10272), .B(n10271), .Z(n10267) );
  AND U18420 ( .A(n10273), .B(n10274), .Z(n10228) );
  NAND U18421 ( .A(n10275), .B(n10276), .Z(n10274) );
  OR U18422 ( .A(n10277), .B(n10278), .Z(n10275) );
  NANDN U18423 ( .A(n10279), .B(n10277), .Z(n10273) );
  XNOR U18424 ( .A(n10254), .B(n10280), .Z(N64480) );
  XOR U18425 ( .A(n10256), .B(n10257), .Z(n10280) );
  XNOR U18426 ( .A(n10270), .B(n10281), .Z(n10257) );
  XOR U18427 ( .A(n10271), .B(n10272), .Z(n10281) );
  XOR U18428 ( .A(n10277), .B(n10282), .Z(n10272) );
  XOR U18429 ( .A(n10276), .B(n10279), .Z(n10282) );
  IV U18430 ( .A(n10278), .Z(n10279) );
  NAND U18431 ( .A(n10283), .B(n10284), .Z(n10278) );
  OR U18432 ( .A(n10285), .B(n10286), .Z(n10284) );
  OR U18433 ( .A(n10287), .B(n10288), .Z(n10283) );
  NAND U18434 ( .A(n10289), .B(n10290), .Z(n10276) );
  OR U18435 ( .A(n10291), .B(n10292), .Z(n10290) );
  OR U18436 ( .A(n10293), .B(n10294), .Z(n10289) );
  NOR U18437 ( .A(n10295), .B(n10296), .Z(n10277) );
  ANDN U18438 ( .B(n10297), .A(n10298), .Z(n10271) );
  XNOR U18439 ( .A(n10264), .B(n10299), .Z(n10270) );
  XNOR U18440 ( .A(n10263), .B(n10265), .Z(n10299) );
  NAND U18441 ( .A(n10300), .B(n10301), .Z(n10265) );
  OR U18442 ( .A(n10302), .B(n10303), .Z(n10301) );
  OR U18443 ( .A(n10304), .B(n10305), .Z(n10300) );
  NAND U18444 ( .A(n10306), .B(n10307), .Z(n10263) );
  OR U18445 ( .A(n10308), .B(n10309), .Z(n10307) );
  OR U18446 ( .A(n10310), .B(n10311), .Z(n10306) );
  ANDN U18447 ( .B(n10312), .A(n10313), .Z(n10264) );
  IV U18448 ( .A(n10314), .Z(n10312) );
  ANDN U18449 ( .B(n10315), .A(n10316), .Z(n10256) );
  XOR U18450 ( .A(n10242), .B(n10317), .Z(n10254) );
  XOR U18451 ( .A(n10243), .B(n10244), .Z(n10317) );
  XOR U18452 ( .A(n10249), .B(n10318), .Z(n10244) );
  XOR U18453 ( .A(n10248), .B(n10251), .Z(n10318) );
  IV U18454 ( .A(n10250), .Z(n10251) );
  NAND U18455 ( .A(n10319), .B(n10320), .Z(n10250) );
  OR U18456 ( .A(n10321), .B(n10322), .Z(n10320) );
  OR U18457 ( .A(n10323), .B(n10324), .Z(n10319) );
  NAND U18458 ( .A(n10325), .B(n10326), .Z(n10248) );
  OR U18459 ( .A(n10327), .B(n10328), .Z(n10326) );
  OR U18460 ( .A(n10329), .B(n10330), .Z(n10325) );
  NOR U18461 ( .A(n10331), .B(n10332), .Z(n10249) );
  ANDN U18462 ( .B(n10333), .A(n10334), .Z(n10243) );
  IV U18463 ( .A(n10335), .Z(n10333) );
  XNOR U18464 ( .A(n10236), .B(n10336), .Z(n10242) );
  XNOR U18465 ( .A(n10235), .B(n10237), .Z(n10336) );
  NAND U18466 ( .A(n10337), .B(n10338), .Z(n10237) );
  OR U18467 ( .A(n10339), .B(n10340), .Z(n10338) );
  OR U18468 ( .A(n10341), .B(n10342), .Z(n10337) );
  NAND U18469 ( .A(n10343), .B(n10344), .Z(n10235) );
  OR U18470 ( .A(n10345), .B(n10346), .Z(n10344) );
  OR U18471 ( .A(n10347), .B(n10348), .Z(n10343) );
  ANDN U18472 ( .B(n10349), .A(n10350), .Z(n10236) );
  IV U18473 ( .A(n10351), .Z(n10349) );
  XNOR U18474 ( .A(n10316), .B(n10315), .Z(N64479) );
  XOR U18475 ( .A(n10335), .B(n10334), .Z(n10315) );
  XNOR U18476 ( .A(n10350), .B(n10351), .Z(n10334) );
  XNOR U18477 ( .A(n10345), .B(n10346), .Z(n10351) );
  XNOR U18478 ( .A(n10347), .B(n10348), .Z(n10346) );
  XNOR U18479 ( .A(y[7189]), .B(x[7189]), .Z(n10348) );
  XNOR U18480 ( .A(y[7190]), .B(x[7190]), .Z(n10347) );
  XNOR U18481 ( .A(y[7188]), .B(x[7188]), .Z(n10345) );
  XNOR U18482 ( .A(n10339), .B(n10340), .Z(n10350) );
  XNOR U18483 ( .A(y[7185]), .B(x[7185]), .Z(n10340) );
  XNOR U18484 ( .A(n10341), .B(n10342), .Z(n10339) );
  XNOR U18485 ( .A(y[7186]), .B(x[7186]), .Z(n10342) );
  XNOR U18486 ( .A(y[7187]), .B(x[7187]), .Z(n10341) );
  XNOR U18487 ( .A(n10332), .B(n10331), .Z(n10335) );
  XNOR U18488 ( .A(n10327), .B(n10328), .Z(n10331) );
  XNOR U18489 ( .A(y[7182]), .B(x[7182]), .Z(n10328) );
  XNOR U18490 ( .A(n10329), .B(n10330), .Z(n10327) );
  XNOR U18491 ( .A(y[7183]), .B(x[7183]), .Z(n10330) );
  XNOR U18492 ( .A(y[7184]), .B(x[7184]), .Z(n10329) );
  XNOR U18493 ( .A(n10321), .B(n10322), .Z(n10332) );
  XNOR U18494 ( .A(y[7179]), .B(x[7179]), .Z(n10322) );
  XNOR U18495 ( .A(n10323), .B(n10324), .Z(n10321) );
  XNOR U18496 ( .A(y[7180]), .B(x[7180]), .Z(n10324) );
  XNOR U18497 ( .A(y[7181]), .B(x[7181]), .Z(n10323) );
  XOR U18498 ( .A(n10297), .B(n10298), .Z(n10316) );
  XNOR U18499 ( .A(n10313), .B(n10314), .Z(n10298) );
  XNOR U18500 ( .A(n10308), .B(n10309), .Z(n10314) );
  XNOR U18501 ( .A(n10310), .B(n10311), .Z(n10309) );
  XNOR U18502 ( .A(y[7177]), .B(x[7177]), .Z(n10311) );
  XNOR U18503 ( .A(y[7178]), .B(x[7178]), .Z(n10310) );
  XNOR U18504 ( .A(y[7176]), .B(x[7176]), .Z(n10308) );
  XNOR U18505 ( .A(n10302), .B(n10303), .Z(n10313) );
  XNOR U18506 ( .A(y[7173]), .B(x[7173]), .Z(n10303) );
  XNOR U18507 ( .A(n10304), .B(n10305), .Z(n10302) );
  XNOR U18508 ( .A(y[7174]), .B(x[7174]), .Z(n10305) );
  XNOR U18509 ( .A(y[7175]), .B(x[7175]), .Z(n10304) );
  XOR U18510 ( .A(n10296), .B(n10295), .Z(n10297) );
  XNOR U18511 ( .A(n10291), .B(n10292), .Z(n10295) );
  XNOR U18512 ( .A(y[7170]), .B(x[7170]), .Z(n10292) );
  XNOR U18513 ( .A(n10293), .B(n10294), .Z(n10291) );
  XNOR U18514 ( .A(y[7171]), .B(x[7171]), .Z(n10294) );
  XNOR U18515 ( .A(y[7172]), .B(x[7172]), .Z(n10293) );
  XNOR U18516 ( .A(n10285), .B(n10286), .Z(n10296) );
  XNOR U18517 ( .A(y[7167]), .B(x[7167]), .Z(n10286) );
  XNOR U18518 ( .A(n10287), .B(n10288), .Z(n10285) );
  XNOR U18519 ( .A(y[7168]), .B(x[7168]), .Z(n10288) );
  XNOR U18520 ( .A(y[7169]), .B(x[7169]), .Z(n10287) );
  NAND U18521 ( .A(n10352), .B(n10353), .Z(N64470) );
  NANDN U18522 ( .A(n10354), .B(n10355), .Z(n10353) );
  OR U18523 ( .A(n10356), .B(n10357), .Z(n10355) );
  NAND U18524 ( .A(n10356), .B(n10357), .Z(n10352) );
  XOR U18525 ( .A(n10356), .B(n10358), .Z(N64469) );
  XNOR U18526 ( .A(n10354), .B(n10357), .Z(n10358) );
  AND U18527 ( .A(n10359), .B(n10360), .Z(n10357) );
  NANDN U18528 ( .A(n10361), .B(n10362), .Z(n10360) );
  NANDN U18529 ( .A(n10363), .B(n10364), .Z(n10362) );
  NANDN U18530 ( .A(n10364), .B(n10363), .Z(n10359) );
  NAND U18531 ( .A(n10365), .B(n10366), .Z(n10354) );
  NANDN U18532 ( .A(n10367), .B(n10368), .Z(n10366) );
  OR U18533 ( .A(n10369), .B(n10370), .Z(n10368) );
  NAND U18534 ( .A(n10370), .B(n10369), .Z(n10365) );
  AND U18535 ( .A(n10371), .B(n10372), .Z(n10356) );
  NANDN U18536 ( .A(n10373), .B(n10374), .Z(n10372) );
  NANDN U18537 ( .A(n10375), .B(n10376), .Z(n10374) );
  NANDN U18538 ( .A(n10376), .B(n10375), .Z(n10371) );
  XOR U18539 ( .A(n10370), .B(n10377), .Z(N64468) );
  XOR U18540 ( .A(n10367), .B(n10369), .Z(n10377) );
  XNOR U18541 ( .A(n10363), .B(n10378), .Z(n10369) );
  XNOR U18542 ( .A(n10361), .B(n10364), .Z(n10378) );
  NAND U18543 ( .A(n10379), .B(n10380), .Z(n10364) );
  NAND U18544 ( .A(n10381), .B(n10382), .Z(n10380) );
  OR U18545 ( .A(n10383), .B(n10384), .Z(n10381) );
  NANDN U18546 ( .A(n10385), .B(n10383), .Z(n10379) );
  IV U18547 ( .A(n10384), .Z(n10385) );
  NAND U18548 ( .A(n10386), .B(n10387), .Z(n10361) );
  NAND U18549 ( .A(n10388), .B(n10389), .Z(n10387) );
  NANDN U18550 ( .A(n10390), .B(n10391), .Z(n10388) );
  NANDN U18551 ( .A(n10391), .B(n10390), .Z(n10386) );
  AND U18552 ( .A(n10392), .B(n10393), .Z(n10363) );
  NAND U18553 ( .A(n10394), .B(n10395), .Z(n10393) );
  OR U18554 ( .A(n10396), .B(n10397), .Z(n10394) );
  NANDN U18555 ( .A(n10398), .B(n10396), .Z(n10392) );
  NAND U18556 ( .A(n10399), .B(n10400), .Z(n10367) );
  NANDN U18557 ( .A(n10401), .B(n10402), .Z(n10400) );
  OR U18558 ( .A(n10403), .B(n10404), .Z(n10402) );
  NANDN U18559 ( .A(n10405), .B(n10403), .Z(n10399) );
  IV U18560 ( .A(n10404), .Z(n10405) );
  XNOR U18561 ( .A(n10375), .B(n10406), .Z(n10370) );
  XNOR U18562 ( .A(n10373), .B(n10376), .Z(n10406) );
  NAND U18563 ( .A(n10407), .B(n10408), .Z(n10376) );
  NAND U18564 ( .A(n10409), .B(n10410), .Z(n10408) );
  OR U18565 ( .A(n10411), .B(n10412), .Z(n10409) );
  NANDN U18566 ( .A(n10413), .B(n10411), .Z(n10407) );
  IV U18567 ( .A(n10412), .Z(n10413) );
  NAND U18568 ( .A(n10414), .B(n10415), .Z(n10373) );
  NAND U18569 ( .A(n10416), .B(n10417), .Z(n10415) );
  NANDN U18570 ( .A(n10418), .B(n10419), .Z(n10416) );
  NANDN U18571 ( .A(n10419), .B(n10418), .Z(n10414) );
  AND U18572 ( .A(n10420), .B(n10421), .Z(n10375) );
  NAND U18573 ( .A(n10422), .B(n10423), .Z(n10421) );
  OR U18574 ( .A(n10424), .B(n10425), .Z(n10422) );
  NANDN U18575 ( .A(n10426), .B(n10424), .Z(n10420) );
  XNOR U18576 ( .A(n10401), .B(n10427), .Z(N64467) );
  XOR U18577 ( .A(n10403), .B(n10404), .Z(n10427) );
  XNOR U18578 ( .A(n10417), .B(n10428), .Z(n10404) );
  XOR U18579 ( .A(n10418), .B(n10419), .Z(n10428) );
  XOR U18580 ( .A(n10424), .B(n10429), .Z(n10419) );
  XOR U18581 ( .A(n10423), .B(n10426), .Z(n10429) );
  IV U18582 ( .A(n10425), .Z(n10426) );
  NAND U18583 ( .A(n10430), .B(n10431), .Z(n10425) );
  OR U18584 ( .A(n10432), .B(n10433), .Z(n10431) );
  OR U18585 ( .A(n10434), .B(n10435), .Z(n10430) );
  NAND U18586 ( .A(n10436), .B(n10437), .Z(n10423) );
  OR U18587 ( .A(n10438), .B(n10439), .Z(n10437) );
  OR U18588 ( .A(n10440), .B(n10441), .Z(n10436) );
  NOR U18589 ( .A(n10442), .B(n10443), .Z(n10424) );
  ANDN U18590 ( .B(n10444), .A(n10445), .Z(n10418) );
  XNOR U18591 ( .A(n10411), .B(n10446), .Z(n10417) );
  XNOR U18592 ( .A(n10410), .B(n10412), .Z(n10446) );
  NAND U18593 ( .A(n10447), .B(n10448), .Z(n10412) );
  OR U18594 ( .A(n10449), .B(n10450), .Z(n10448) );
  OR U18595 ( .A(n10451), .B(n10452), .Z(n10447) );
  NAND U18596 ( .A(n10453), .B(n10454), .Z(n10410) );
  OR U18597 ( .A(n10455), .B(n10456), .Z(n10454) );
  OR U18598 ( .A(n10457), .B(n10458), .Z(n10453) );
  ANDN U18599 ( .B(n10459), .A(n10460), .Z(n10411) );
  IV U18600 ( .A(n10461), .Z(n10459) );
  ANDN U18601 ( .B(n10462), .A(n10463), .Z(n10403) );
  XOR U18602 ( .A(n10389), .B(n10464), .Z(n10401) );
  XOR U18603 ( .A(n10390), .B(n10391), .Z(n10464) );
  XOR U18604 ( .A(n10396), .B(n10465), .Z(n10391) );
  XOR U18605 ( .A(n10395), .B(n10398), .Z(n10465) );
  IV U18606 ( .A(n10397), .Z(n10398) );
  NAND U18607 ( .A(n10466), .B(n10467), .Z(n10397) );
  OR U18608 ( .A(n10468), .B(n10469), .Z(n10467) );
  OR U18609 ( .A(n10470), .B(n10471), .Z(n10466) );
  NAND U18610 ( .A(n10472), .B(n10473), .Z(n10395) );
  OR U18611 ( .A(n10474), .B(n10475), .Z(n10473) );
  OR U18612 ( .A(n10476), .B(n10477), .Z(n10472) );
  NOR U18613 ( .A(n10478), .B(n10479), .Z(n10396) );
  ANDN U18614 ( .B(n10480), .A(n10481), .Z(n10390) );
  IV U18615 ( .A(n10482), .Z(n10480) );
  XNOR U18616 ( .A(n10383), .B(n10483), .Z(n10389) );
  XNOR U18617 ( .A(n10382), .B(n10384), .Z(n10483) );
  NAND U18618 ( .A(n10484), .B(n10485), .Z(n10384) );
  OR U18619 ( .A(n10486), .B(n10487), .Z(n10485) );
  OR U18620 ( .A(n10488), .B(n10489), .Z(n10484) );
  NAND U18621 ( .A(n10490), .B(n10491), .Z(n10382) );
  OR U18622 ( .A(n10492), .B(n10493), .Z(n10491) );
  OR U18623 ( .A(n10494), .B(n10495), .Z(n10490) );
  ANDN U18624 ( .B(n10496), .A(n10497), .Z(n10383) );
  IV U18625 ( .A(n10498), .Z(n10496) );
  XNOR U18626 ( .A(n10463), .B(n10462), .Z(N64466) );
  XOR U18627 ( .A(n10482), .B(n10481), .Z(n10462) );
  XNOR U18628 ( .A(n10497), .B(n10498), .Z(n10481) );
  XNOR U18629 ( .A(n10492), .B(n10493), .Z(n10498) );
  XNOR U18630 ( .A(n10494), .B(n10495), .Z(n10493) );
  XNOR U18631 ( .A(y[7165]), .B(x[7165]), .Z(n10495) );
  XNOR U18632 ( .A(y[7166]), .B(x[7166]), .Z(n10494) );
  XNOR U18633 ( .A(y[7164]), .B(x[7164]), .Z(n10492) );
  XNOR U18634 ( .A(n10486), .B(n10487), .Z(n10497) );
  XNOR U18635 ( .A(y[7161]), .B(x[7161]), .Z(n10487) );
  XNOR U18636 ( .A(n10488), .B(n10489), .Z(n10486) );
  XNOR U18637 ( .A(y[7162]), .B(x[7162]), .Z(n10489) );
  XNOR U18638 ( .A(y[7163]), .B(x[7163]), .Z(n10488) );
  XNOR U18639 ( .A(n10479), .B(n10478), .Z(n10482) );
  XNOR U18640 ( .A(n10474), .B(n10475), .Z(n10478) );
  XNOR U18641 ( .A(y[7158]), .B(x[7158]), .Z(n10475) );
  XNOR U18642 ( .A(n10476), .B(n10477), .Z(n10474) );
  XNOR U18643 ( .A(y[7159]), .B(x[7159]), .Z(n10477) );
  XNOR U18644 ( .A(y[7160]), .B(x[7160]), .Z(n10476) );
  XNOR U18645 ( .A(n10468), .B(n10469), .Z(n10479) );
  XNOR U18646 ( .A(y[7155]), .B(x[7155]), .Z(n10469) );
  XNOR U18647 ( .A(n10470), .B(n10471), .Z(n10468) );
  XNOR U18648 ( .A(y[7156]), .B(x[7156]), .Z(n10471) );
  XNOR U18649 ( .A(y[7157]), .B(x[7157]), .Z(n10470) );
  XOR U18650 ( .A(n10444), .B(n10445), .Z(n10463) );
  XNOR U18651 ( .A(n10460), .B(n10461), .Z(n10445) );
  XNOR U18652 ( .A(n10455), .B(n10456), .Z(n10461) );
  XNOR U18653 ( .A(n10457), .B(n10458), .Z(n10456) );
  XNOR U18654 ( .A(y[7153]), .B(x[7153]), .Z(n10458) );
  XNOR U18655 ( .A(y[7154]), .B(x[7154]), .Z(n10457) );
  XNOR U18656 ( .A(y[7152]), .B(x[7152]), .Z(n10455) );
  XNOR U18657 ( .A(n10449), .B(n10450), .Z(n10460) );
  XNOR U18658 ( .A(y[7149]), .B(x[7149]), .Z(n10450) );
  XNOR U18659 ( .A(n10451), .B(n10452), .Z(n10449) );
  XNOR U18660 ( .A(y[7150]), .B(x[7150]), .Z(n10452) );
  XNOR U18661 ( .A(y[7151]), .B(x[7151]), .Z(n10451) );
  XOR U18662 ( .A(n10443), .B(n10442), .Z(n10444) );
  XNOR U18663 ( .A(n10438), .B(n10439), .Z(n10442) );
  XNOR U18664 ( .A(y[7146]), .B(x[7146]), .Z(n10439) );
  XNOR U18665 ( .A(n10440), .B(n10441), .Z(n10438) );
  XNOR U18666 ( .A(y[7147]), .B(x[7147]), .Z(n10441) );
  XNOR U18667 ( .A(y[7148]), .B(x[7148]), .Z(n10440) );
  XNOR U18668 ( .A(n10432), .B(n10433), .Z(n10443) );
  XNOR U18669 ( .A(y[7143]), .B(x[7143]), .Z(n10433) );
  XNOR U18670 ( .A(n10434), .B(n10435), .Z(n10432) );
  XNOR U18671 ( .A(y[7144]), .B(x[7144]), .Z(n10435) );
  XNOR U18672 ( .A(y[7145]), .B(x[7145]), .Z(n10434) );
  NAND U18673 ( .A(n10499), .B(n10500), .Z(N64457) );
  NANDN U18674 ( .A(n10501), .B(n10502), .Z(n10500) );
  OR U18675 ( .A(n10503), .B(n10504), .Z(n10502) );
  NAND U18676 ( .A(n10503), .B(n10504), .Z(n10499) );
  XOR U18677 ( .A(n10503), .B(n10505), .Z(N64456) );
  XNOR U18678 ( .A(n10501), .B(n10504), .Z(n10505) );
  AND U18679 ( .A(n10506), .B(n10507), .Z(n10504) );
  NANDN U18680 ( .A(n10508), .B(n10509), .Z(n10507) );
  NANDN U18681 ( .A(n10510), .B(n10511), .Z(n10509) );
  NANDN U18682 ( .A(n10511), .B(n10510), .Z(n10506) );
  NAND U18683 ( .A(n10512), .B(n10513), .Z(n10501) );
  NANDN U18684 ( .A(n10514), .B(n10515), .Z(n10513) );
  OR U18685 ( .A(n10516), .B(n10517), .Z(n10515) );
  NAND U18686 ( .A(n10517), .B(n10516), .Z(n10512) );
  AND U18687 ( .A(n10518), .B(n10519), .Z(n10503) );
  NANDN U18688 ( .A(n10520), .B(n10521), .Z(n10519) );
  NANDN U18689 ( .A(n10522), .B(n10523), .Z(n10521) );
  NANDN U18690 ( .A(n10523), .B(n10522), .Z(n10518) );
  XOR U18691 ( .A(n10517), .B(n10524), .Z(N64455) );
  XOR U18692 ( .A(n10514), .B(n10516), .Z(n10524) );
  XNOR U18693 ( .A(n10510), .B(n10525), .Z(n10516) );
  XNOR U18694 ( .A(n10508), .B(n10511), .Z(n10525) );
  NAND U18695 ( .A(n10526), .B(n10527), .Z(n10511) );
  NAND U18696 ( .A(n10528), .B(n10529), .Z(n10527) );
  OR U18697 ( .A(n10530), .B(n10531), .Z(n10528) );
  NANDN U18698 ( .A(n10532), .B(n10530), .Z(n10526) );
  IV U18699 ( .A(n10531), .Z(n10532) );
  NAND U18700 ( .A(n10533), .B(n10534), .Z(n10508) );
  NAND U18701 ( .A(n10535), .B(n10536), .Z(n10534) );
  NANDN U18702 ( .A(n10537), .B(n10538), .Z(n10535) );
  NANDN U18703 ( .A(n10538), .B(n10537), .Z(n10533) );
  AND U18704 ( .A(n10539), .B(n10540), .Z(n10510) );
  NAND U18705 ( .A(n10541), .B(n10542), .Z(n10540) );
  OR U18706 ( .A(n10543), .B(n10544), .Z(n10541) );
  NANDN U18707 ( .A(n10545), .B(n10543), .Z(n10539) );
  NAND U18708 ( .A(n10546), .B(n10547), .Z(n10514) );
  NANDN U18709 ( .A(n10548), .B(n10549), .Z(n10547) );
  OR U18710 ( .A(n10550), .B(n10551), .Z(n10549) );
  NANDN U18711 ( .A(n10552), .B(n10550), .Z(n10546) );
  IV U18712 ( .A(n10551), .Z(n10552) );
  XNOR U18713 ( .A(n10522), .B(n10553), .Z(n10517) );
  XNOR U18714 ( .A(n10520), .B(n10523), .Z(n10553) );
  NAND U18715 ( .A(n10554), .B(n10555), .Z(n10523) );
  NAND U18716 ( .A(n10556), .B(n10557), .Z(n10555) );
  OR U18717 ( .A(n10558), .B(n10559), .Z(n10556) );
  NANDN U18718 ( .A(n10560), .B(n10558), .Z(n10554) );
  IV U18719 ( .A(n10559), .Z(n10560) );
  NAND U18720 ( .A(n10561), .B(n10562), .Z(n10520) );
  NAND U18721 ( .A(n10563), .B(n10564), .Z(n10562) );
  NANDN U18722 ( .A(n10565), .B(n10566), .Z(n10563) );
  NANDN U18723 ( .A(n10566), .B(n10565), .Z(n10561) );
  AND U18724 ( .A(n10567), .B(n10568), .Z(n10522) );
  NAND U18725 ( .A(n10569), .B(n10570), .Z(n10568) );
  OR U18726 ( .A(n10571), .B(n10572), .Z(n10569) );
  NANDN U18727 ( .A(n10573), .B(n10571), .Z(n10567) );
  XNOR U18728 ( .A(n10548), .B(n10574), .Z(N64454) );
  XOR U18729 ( .A(n10550), .B(n10551), .Z(n10574) );
  XNOR U18730 ( .A(n10564), .B(n10575), .Z(n10551) );
  XOR U18731 ( .A(n10565), .B(n10566), .Z(n10575) );
  XOR U18732 ( .A(n10571), .B(n10576), .Z(n10566) );
  XOR U18733 ( .A(n10570), .B(n10573), .Z(n10576) );
  IV U18734 ( .A(n10572), .Z(n10573) );
  NAND U18735 ( .A(n10577), .B(n10578), .Z(n10572) );
  OR U18736 ( .A(n10579), .B(n10580), .Z(n10578) );
  OR U18737 ( .A(n10581), .B(n10582), .Z(n10577) );
  NAND U18738 ( .A(n10583), .B(n10584), .Z(n10570) );
  OR U18739 ( .A(n10585), .B(n10586), .Z(n10584) );
  OR U18740 ( .A(n10587), .B(n10588), .Z(n10583) );
  NOR U18741 ( .A(n10589), .B(n10590), .Z(n10571) );
  ANDN U18742 ( .B(n10591), .A(n10592), .Z(n10565) );
  XNOR U18743 ( .A(n10558), .B(n10593), .Z(n10564) );
  XNOR U18744 ( .A(n10557), .B(n10559), .Z(n10593) );
  NAND U18745 ( .A(n10594), .B(n10595), .Z(n10559) );
  OR U18746 ( .A(n10596), .B(n10597), .Z(n10595) );
  OR U18747 ( .A(n10598), .B(n10599), .Z(n10594) );
  NAND U18748 ( .A(n10600), .B(n10601), .Z(n10557) );
  OR U18749 ( .A(n10602), .B(n10603), .Z(n10601) );
  OR U18750 ( .A(n10604), .B(n10605), .Z(n10600) );
  ANDN U18751 ( .B(n10606), .A(n10607), .Z(n10558) );
  IV U18752 ( .A(n10608), .Z(n10606) );
  ANDN U18753 ( .B(n10609), .A(n10610), .Z(n10550) );
  XOR U18754 ( .A(n10536), .B(n10611), .Z(n10548) );
  XOR U18755 ( .A(n10537), .B(n10538), .Z(n10611) );
  XOR U18756 ( .A(n10543), .B(n10612), .Z(n10538) );
  XOR U18757 ( .A(n10542), .B(n10545), .Z(n10612) );
  IV U18758 ( .A(n10544), .Z(n10545) );
  NAND U18759 ( .A(n10613), .B(n10614), .Z(n10544) );
  OR U18760 ( .A(n10615), .B(n10616), .Z(n10614) );
  OR U18761 ( .A(n10617), .B(n10618), .Z(n10613) );
  NAND U18762 ( .A(n10619), .B(n10620), .Z(n10542) );
  OR U18763 ( .A(n10621), .B(n10622), .Z(n10620) );
  OR U18764 ( .A(n10623), .B(n10624), .Z(n10619) );
  NOR U18765 ( .A(n10625), .B(n10626), .Z(n10543) );
  ANDN U18766 ( .B(n10627), .A(n10628), .Z(n10537) );
  IV U18767 ( .A(n10629), .Z(n10627) );
  XNOR U18768 ( .A(n10530), .B(n10630), .Z(n10536) );
  XNOR U18769 ( .A(n10529), .B(n10531), .Z(n10630) );
  NAND U18770 ( .A(n10631), .B(n10632), .Z(n10531) );
  OR U18771 ( .A(n10633), .B(n10634), .Z(n10632) );
  OR U18772 ( .A(n10635), .B(n10636), .Z(n10631) );
  NAND U18773 ( .A(n10637), .B(n10638), .Z(n10529) );
  OR U18774 ( .A(n10639), .B(n10640), .Z(n10638) );
  OR U18775 ( .A(n10641), .B(n10642), .Z(n10637) );
  ANDN U18776 ( .B(n10643), .A(n10644), .Z(n10530) );
  IV U18777 ( .A(n10645), .Z(n10643) );
  XNOR U18778 ( .A(n10610), .B(n10609), .Z(N64453) );
  XOR U18779 ( .A(n10629), .B(n10628), .Z(n10609) );
  XNOR U18780 ( .A(n10644), .B(n10645), .Z(n10628) );
  XNOR U18781 ( .A(n10639), .B(n10640), .Z(n10645) );
  XNOR U18782 ( .A(n10641), .B(n10642), .Z(n10640) );
  XNOR U18783 ( .A(y[7141]), .B(x[7141]), .Z(n10642) );
  XNOR U18784 ( .A(y[7142]), .B(x[7142]), .Z(n10641) );
  XNOR U18785 ( .A(y[7140]), .B(x[7140]), .Z(n10639) );
  XNOR U18786 ( .A(n10633), .B(n10634), .Z(n10644) );
  XNOR U18787 ( .A(y[7137]), .B(x[7137]), .Z(n10634) );
  XNOR U18788 ( .A(n10635), .B(n10636), .Z(n10633) );
  XNOR U18789 ( .A(y[7138]), .B(x[7138]), .Z(n10636) );
  XNOR U18790 ( .A(y[7139]), .B(x[7139]), .Z(n10635) );
  XNOR U18791 ( .A(n10626), .B(n10625), .Z(n10629) );
  XNOR U18792 ( .A(n10621), .B(n10622), .Z(n10625) );
  XNOR U18793 ( .A(y[7134]), .B(x[7134]), .Z(n10622) );
  XNOR U18794 ( .A(n10623), .B(n10624), .Z(n10621) );
  XNOR U18795 ( .A(y[7135]), .B(x[7135]), .Z(n10624) );
  XNOR U18796 ( .A(y[7136]), .B(x[7136]), .Z(n10623) );
  XNOR U18797 ( .A(n10615), .B(n10616), .Z(n10626) );
  XNOR U18798 ( .A(y[7131]), .B(x[7131]), .Z(n10616) );
  XNOR U18799 ( .A(n10617), .B(n10618), .Z(n10615) );
  XNOR U18800 ( .A(y[7132]), .B(x[7132]), .Z(n10618) );
  XNOR U18801 ( .A(y[7133]), .B(x[7133]), .Z(n10617) );
  XOR U18802 ( .A(n10591), .B(n10592), .Z(n10610) );
  XNOR U18803 ( .A(n10607), .B(n10608), .Z(n10592) );
  XNOR U18804 ( .A(n10602), .B(n10603), .Z(n10608) );
  XNOR U18805 ( .A(n10604), .B(n10605), .Z(n10603) );
  XNOR U18806 ( .A(y[7129]), .B(x[7129]), .Z(n10605) );
  XNOR U18807 ( .A(y[7130]), .B(x[7130]), .Z(n10604) );
  XNOR U18808 ( .A(y[7128]), .B(x[7128]), .Z(n10602) );
  XNOR U18809 ( .A(n10596), .B(n10597), .Z(n10607) );
  XNOR U18810 ( .A(y[7125]), .B(x[7125]), .Z(n10597) );
  XNOR U18811 ( .A(n10598), .B(n10599), .Z(n10596) );
  XNOR U18812 ( .A(y[7126]), .B(x[7126]), .Z(n10599) );
  XNOR U18813 ( .A(y[7127]), .B(x[7127]), .Z(n10598) );
  XOR U18814 ( .A(n10590), .B(n10589), .Z(n10591) );
  XNOR U18815 ( .A(n10585), .B(n10586), .Z(n10589) );
  XNOR U18816 ( .A(y[7122]), .B(x[7122]), .Z(n10586) );
  XNOR U18817 ( .A(n10587), .B(n10588), .Z(n10585) );
  XNOR U18818 ( .A(y[7123]), .B(x[7123]), .Z(n10588) );
  XNOR U18819 ( .A(y[7124]), .B(x[7124]), .Z(n10587) );
  XNOR U18820 ( .A(n10579), .B(n10580), .Z(n10590) );
  XNOR U18821 ( .A(y[7119]), .B(x[7119]), .Z(n10580) );
  XNOR U18822 ( .A(n10581), .B(n10582), .Z(n10579) );
  XNOR U18823 ( .A(y[7120]), .B(x[7120]), .Z(n10582) );
  XNOR U18824 ( .A(y[7121]), .B(x[7121]), .Z(n10581) );
  NAND U18825 ( .A(n10646), .B(n10647), .Z(N64444) );
  NANDN U18826 ( .A(n10648), .B(n10649), .Z(n10647) );
  OR U18827 ( .A(n10650), .B(n10651), .Z(n10649) );
  NAND U18828 ( .A(n10650), .B(n10651), .Z(n10646) );
  XOR U18829 ( .A(n10650), .B(n10652), .Z(N64443) );
  XNOR U18830 ( .A(n10648), .B(n10651), .Z(n10652) );
  AND U18831 ( .A(n10653), .B(n10654), .Z(n10651) );
  NANDN U18832 ( .A(n10655), .B(n10656), .Z(n10654) );
  NANDN U18833 ( .A(n10657), .B(n10658), .Z(n10656) );
  NANDN U18834 ( .A(n10658), .B(n10657), .Z(n10653) );
  NAND U18835 ( .A(n10659), .B(n10660), .Z(n10648) );
  NANDN U18836 ( .A(n10661), .B(n10662), .Z(n10660) );
  OR U18837 ( .A(n10663), .B(n10664), .Z(n10662) );
  NAND U18838 ( .A(n10664), .B(n10663), .Z(n10659) );
  AND U18839 ( .A(n10665), .B(n10666), .Z(n10650) );
  NANDN U18840 ( .A(n10667), .B(n10668), .Z(n10666) );
  NANDN U18841 ( .A(n10669), .B(n10670), .Z(n10668) );
  NANDN U18842 ( .A(n10670), .B(n10669), .Z(n10665) );
  XOR U18843 ( .A(n10664), .B(n10671), .Z(N64442) );
  XOR U18844 ( .A(n10661), .B(n10663), .Z(n10671) );
  XNOR U18845 ( .A(n10657), .B(n10672), .Z(n10663) );
  XNOR U18846 ( .A(n10655), .B(n10658), .Z(n10672) );
  NAND U18847 ( .A(n10673), .B(n10674), .Z(n10658) );
  NAND U18848 ( .A(n10675), .B(n10676), .Z(n10674) );
  OR U18849 ( .A(n10677), .B(n10678), .Z(n10675) );
  NANDN U18850 ( .A(n10679), .B(n10677), .Z(n10673) );
  IV U18851 ( .A(n10678), .Z(n10679) );
  NAND U18852 ( .A(n10680), .B(n10681), .Z(n10655) );
  NAND U18853 ( .A(n10682), .B(n10683), .Z(n10681) );
  NANDN U18854 ( .A(n10684), .B(n10685), .Z(n10682) );
  NANDN U18855 ( .A(n10685), .B(n10684), .Z(n10680) );
  AND U18856 ( .A(n10686), .B(n10687), .Z(n10657) );
  NAND U18857 ( .A(n10688), .B(n10689), .Z(n10687) );
  OR U18858 ( .A(n10690), .B(n10691), .Z(n10688) );
  NANDN U18859 ( .A(n10692), .B(n10690), .Z(n10686) );
  NAND U18860 ( .A(n10693), .B(n10694), .Z(n10661) );
  NANDN U18861 ( .A(n10695), .B(n10696), .Z(n10694) );
  OR U18862 ( .A(n10697), .B(n10698), .Z(n10696) );
  NANDN U18863 ( .A(n10699), .B(n10697), .Z(n10693) );
  IV U18864 ( .A(n10698), .Z(n10699) );
  XNOR U18865 ( .A(n10669), .B(n10700), .Z(n10664) );
  XNOR U18866 ( .A(n10667), .B(n10670), .Z(n10700) );
  NAND U18867 ( .A(n10701), .B(n10702), .Z(n10670) );
  NAND U18868 ( .A(n10703), .B(n10704), .Z(n10702) );
  OR U18869 ( .A(n10705), .B(n10706), .Z(n10703) );
  NANDN U18870 ( .A(n10707), .B(n10705), .Z(n10701) );
  IV U18871 ( .A(n10706), .Z(n10707) );
  NAND U18872 ( .A(n10708), .B(n10709), .Z(n10667) );
  NAND U18873 ( .A(n10710), .B(n10711), .Z(n10709) );
  NANDN U18874 ( .A(n10712), .B(n10713), .Z(n10710) );
  NANDN U18875 ( .A(n10713), .B(n10712), .Z(n10708) );
  AND U18876 ( .A(n10714), .B(n10715), .Z(n10669) );
  NAND U18877 ( .A(n10716), .B(n10717), .Z(n10715) );
  OR U18878 ( .A(n10718), .B(n10719), .Z(n10716) );
  NANDN U18879 ( .A(n10720), .B(n10718), .Z(n10714) );
  XNOR U18880 ( .A(n10695), .B(n10721), .Z(N64441) );
  XOR U18881 ( .A(n10697), .B(n10698), .Z(n10721) );
  XNOR U18882 ( .A(n10711), .B(n10722), .Z(n10698) );
  XOR U18883 ( .A(n10712), .B(n10713), .Z(n10722) );
  XOR U18884 ( .A(n10718), .B(n10723), .Z(n10713) );
  XOR U18885 ( .A(n10717), .B(n10720), .Z(n10723) );
  IV U18886 ( .A(n10719), .Z(n10720) );
  NAND U18887 ( .A(n10724), .B(n10725), .Z(n10719) );
  OR U18888 ( .A(n10726), .B(n10727), .Z(n10725) );
  OR U18889 ( .A(n10728), .B(n10729), .Z(n10724) );
  NAND U18890 ( .A(n10730), .B(n10731), .Z(n10717) );
  OR U18891 ( .A(n10732), .B(n10733), .Z(n10731) );
  OR U18892 ( .A(n10734), .B(n10735), .Z(n10730) );
  NOR U18893 ( .A(n10736), .B(n10737), .Z(n10718) );
  ANDN U18894 ( .B(n10738), .A(n10739), .Z(n10712) );
  XNOR U18895 ( .A(n10705), .B(n10740), .Z(n10711) );
  XNOR U18896 ( .A(n10704), .B(n10706), .Z(n10740) );
  NAND U18897 ( .A(n10741), .B(n10742), .Z(n10706) );
  OR U18898 ( .A(n10743), .B(n10744), .Z(n10742) );
  OR U18899 ( .A(n10745), .B(n10746), .Z(n10741) );
  NAND U18900 ( .A(n10747), .B(n10748), .Z(n10704) );
  OR U18901 ( .A(n10749), .B(n10750), .Z(n10748) );
  OR U18902 ( .A(n10751), .B(n10752), .Z(n10747) );
  ANDN U18903 ( .B(n10753), .A(n10754), .Z(n10705) );
  IV U18904 ( .A(n10755), .Z(n10753) );
  ANDN U18905 ( .B(n10756), .A(n10757), .Z(n10697) );
  XOR U18906 ( .A(n10683), .B(n10758), .Z(n10695) );
  XOR U18907 ( .A(n10684), .B(n10685), .Z(n10758) );
  XOR U18908 ( .A(n10690), .B(n10759), .Z(n10685) );
  XOR U18909 ( .A(n10689), .B(n10692), .Z(n10759) );
  IV U18910 ( .A(n10691), .Z(n10692) );
  NAND U18911 ( .A(n10760), .B(n10761), .Z(n10691) );
  OR U18912 ( .A(n10762), .B(n10763), .Z(n10761) );
  OR U18913 ( .A(n10764), .B(n10765), .Z(n10760) );
  NAND U18914 ( .A(n10766), .B(n10767), .Z(n10689) );
  OR U18915 ( .A(n10768), .B(n10769), .Z(n10767) );
  OR U18916 ( .A(n10770), .B(n10771), .Z(n10766) );
  NOR U18917 ( .A(n10772), .B(n10773), .Z(n10690) );
  ANDN U18918 ( .B(n10774), .A(n10775), .Z(n10684) );
  IV U18919 ( .A(n10776), .Z(n10774) );
  XNOR U18920 ( .A(n10677), .B(n10777), .Z(n10683) );
  XNOR U18921 ( .A(n10676), .B(n10678), .Z(n10777) );
  NAND U18922 ( .A(n10778), .B(n10779), .Z(n10678) );
  OR U18923 ( .A(n10780), .B(n10781), .Z(n10779) );
  OR U18924 ( .A(n10782), .B(n10783), .Z(n10778) );
  NAND U18925 ( .A(n10784), .B(n10785), .Z(n10676) );
  OR U18926 ( .A(n10786), .B(n10787), .Z(n10785) );
  OR U18927 ( .A(n10788), .B(n10789), .Z(n10784) );
  ANDN U18928 ( .B(n10790), .A(n10791), .Z(n10677) );
  IV U18929 ( .A(n10792), .Z(n10790) );
  XNOR U18930 ( .A(n10757), .B(n10756), .Z(N64440) );
  XOR U18931 ( .A(n10776), .B(n10775), .Z(n10756) );
  XNOR U18932 ( .A(n10791), .B(n10792), .Z(n10775) );
  XNOR U18933 ( .A(n10786), .B(n10787), .Z(n10792) );
  XNOR U18934 ( .A(n10788), .B(n10789), .Z(n10787) );
  XNOR U18935 ( .A(y[7117]), .B(x[7117]), .Z(n10789) );
  XNOR U18936 ( .A(y[7118]), .B(x[7118]), .Z(n10788) );
  XNOR U18937 ( .A(y[7116]), .B(x[7116]), .Z(n10786) );
  XNOR U18938 ( .A(n10780), .B(n10781), .Z(n10791) );
  XNOR U18939 ( .A(y[7113]), .B(x[7113]), .Z(n10781) );
  XNOR U18940 ( .A(n10782), .B(n10783), .Z(n10780) );
  XNOR U18941 ( .A(y[7114]), .B(x[7114]), .Z(n10783) );
  XNOR U18942 ( .A(y[7115]), .B(x[7115]), .Z(n10782) );
  XNOR U18943 ( .A(n10773), .B(n10772), .Z(n10776) );
  XNOR U18944 ( .A(n10768), .B(n10769), .Z(n10772) );
  XNOR U18945 ( .A(y[7110]), .B(x[7110]), .Z(n10769) );
  XNOR U18946 ( .A(n10770), .B(n10771), .Z(n10768) );
  XNOR U18947 ( .A(y[7111]), .B(x[7111]), .Z(n10771) );
  XNOR U18948 ( .A(y[7112]), .B(x[7112]), .Z(n10770) );
  XNOR U18949 ( .A(n10762), .B(n10763), .Z(n10773) );
  XNOR U18950 ( .A(y[7107]), .B(x[7107]), .Z(n10763) );
  XNOR U18951 ( .A(n10764), .B(n10765), .Z(n10762) );
  XNOR U18952 ( .A(y[7108]), .B(x[7108]), .Z(n10765) );
  XNOR U18953 ( .A(y[7109]), .B(x[7109]), .Z(n10764) );
  XOR U18954 ( .A(n10738), .B(n10739), .Z(n10757) );
  XNOR U18955 ( .A(n10754), .B(n10755), .Z(n10739) );
  XNOR U18956 ( .A(n10749), .B(n10750), .Z(n10755) );
  XNOR U18957 ( .A(n10751), .B(n10752), .Z(n10750) );
  XNOR U18958 ( .A(y[7105]), .B(x[7105]), .Z(n10752) );
  XNOR U18959 ( .A(y[7106]), .B(x[7106]), .Z(n10751) );
  XNOR U18960 ( .A(y[7104]), .B(x[7104]), .Z(n10749) );
  XNOR U18961 ( .A(n10743), .B(n10744), .Z(n10754) );
  XNOR U18962 ( .A(y[7101]), .B(x[7101]), .Z(n10744) );
  XNOR U18963 ( .A(n10745), .B(n10746), .Z(n10743) );
  XNOR U18964 ( .A(y[7102]), .B(x[7102]), .Z(n10746) );
  XNOR U18965 ( .A(y[7103]), .B(x[7103]), .Z(n10745) );
  XOR U18966 ( .A(n10737), .B(n10736), .Z(n10738) );
  XNOR U18967 ( .A(n10732), .B(n10733), .Z(n10736) );
  XNOR U18968 ( .A(y[7098]), .B(x[7098]), .Z(n10733) );
  XNOR U18969 ( .A(n10734), .B(n10735), .Z(n10732) );
  XNOR U18970 ( .A(y[7099]), .B(x[7099]), .Z(n10735) );
  XNOR U18971 ( .A(y[7100]), .B(x[7100]), .Z(n10734) );
  XNOR U18972 ( .A(n10726), .B(n10727), .Z(n10737) );
  XNOR U18973 ( .A(y[7095]), .B(x[7095]), .Z(n10727) );
  XNOR U18974 ( .A(n10728), .B(n10729), .Z(n10726) );
  XNOR U18975 ( .A(y[7096]), .B(x[7096]), .Z(n10729) );
  XNOR U18976 ( .A(y[7097]), .B(x[7097]), .Z(n10728) );
  NAND U18977 ( .A(n10793), .B(n10794), .Z(N64431) );
  NANDN U18978 ( .A(n10795), .B(n10796), .Z(n10794) );
  OR U18979 ( .A(n10797), .B(n10798), .Z(n10796) );
  NAND U18980 ( .A(n10797), .B(n10798), .Z(n10793) );
  XOR U18981 ( .A(n10797), .B(n10799), .Z(N64430) );
  XNOR U18982 ( .A(n10795), .B(n10798), .Z(n10799) );
  AND U18983 ( .A(n10800), .B(n10801), .Z(n10798) );
  NANDN U18984 ( .A(n10802), .B(n10803), .Z(n10801) );
  NANDN U18985 ( .A(n10804), .B(n10805), .Z(n10803) );
  NANDN U18986 ( .A(n10805), .B(n10804), .Z(n10800) );
  NAND U18987 ( .A(n10806), .B(n10807), .Z(n10795) );
  NANDN U18988 ( .A(n10808), .B(n10809), .Z(n10807) );
  OR U18989 ( .A(n10810), .B(n10811), .Z(n10809) );
  NAND U18990 ( .A(n10811), .B(n10810), .Z(n10806) );
  AND U18991 ( .A(n10812), .B(n10813), .Z(n10797) );
  NANDN U18992 ( .A(n10814), .B(n10815), .Z(n10813) );
  NANDN U18993 ( .A(n10816), .B(n10817), .Z(n10815) );
  NANDN U18994 ( .A(n10817), .B(n10816), .Z(n10812) );
  XOR U18995 ( .A(n10811), .B(n10818), .Z(N64429) );
  XOR U18996 ( .A(n10808), .B(n10810), .Z(n10818) );
  XNOR U18997 ( .A(n10804), .B(n10819), .Z(n10810) );
  XNOR U18998 ( .A(n10802), .B(n10805), .Z(n10819) );
  NAND U18999 ( .A(n10820), .B(n10821), .Z(n10805) );
  NAND U19000 ( .A(n10822), .B(n10823), .Z(n10821) );
  OR U19001 ( .A(n10824), .B(n10825), .Z(n10822) );
  NANDN U19002 ( .A(n10826), .B(n10824), .Z(n10820) );
  IV U19003 ( .A(n10825), .Z(n10826) );
  NAND U19004 ( .A(n10827), .B(n10828), .Z(n10802) );
  NAND U19005 ( .A(n10829), .B(n10830), .Z(n10828) );
  NANDN U19006 ( .A(n10831), .B(n10832), .Z(n10829) );
  NANDN U19007 ( .A(n10832), .B(n10831), .Z(n10827) );
  AND U19008 ( .A(n10833), .B(n10834), .Z(n10804) );
  NAND U19009 ( .A(n10835), .B(n10836), .Z(n10834) );
  OR U19010 ( .A(n10837), .B(n10838), .Z(n10835) );
  NANDN U19011 ( .A(n10839), .B(n10837), .Z(n10833) );
  NAND U19012 ( .A(n10840), .B(n10841), .Z(n10808) );
  NANDN U19013 ( .A(n10842), .B(n10843), .Z(n10841) );
  OR U19014 ( .A(n10844), .B(n10845), .Z(n10843) );
  NANDN U19015 ( .A(n10846), .B(n10844), .Z(n10840) );
  IV U19016 ( .A(n10845), .Z(n10846) );
  XNOR U19017 ( .A(n10816), .B(n10847), .Z(n10811) );
  XNOR U19018 ( .A(n10814), .B(n10817), .Z(n10847) );
  NAND U19019 ( .A(n10848), .B(n10849), .Z(n10817) );
  NAND U19020 ( .A(n10850), .B(n10851), .Z(n10849) );
  OR U19021 ( .A(n10852), .B(n10853), .Z(n10850) );
  NANDN U19022 ( .A(n10854), .B(n10852), .Z(n10848) );
  IV U19023 ( .A(n10853), .Z(n10854) );
  NAND U19024 ( .A(n10855), .B(n10856), .Z(n10814) );
  NAND U19025 ( .A(n10857), .B(n10858), .Z(n10856) );
  NANDN U19026 ( .A(n10859), .B(n10860), .Z(n10857) );
  NANDN U19027 ( .A(n10860), .B(n10859), .Z(n10855) );
  AND U19028 ( .A(n10861), .B(n10862), .Z(n10816) );
  NAND U19029 ( .A(n10863), .B(n10864), .Z(n10862) );
  OR U19030 ( .A(n10865), .B(n10866), .Z(n10863) );
  NANDN U19031 ( .A(n10867), .B(n10865), .Z(n10861) );
  XNOR U19032 ( .A(n10842), .B(n10868), .Z(N64428) );
  XOR U19033 ( .A(n10844), .B(n10845), .Z(n10868) );
  XNOR U19034 ( .A(n10858), .B(n10869), .Z(n10845) );
  XOR U19035 ( .A(n10859), .B(n10860), .Z(n10869) );
  XOR U19036 ( .A(n10865), .B(n10870), .Z(n10860) );
  XOR U19037 ( .A(n10864), .B(n10867), .Z(n10870) );
  IV U19038 ( .A(n10866), .Z(n10867) );
  NAND U19039 ( .A(n10871), .B(n10872), .Z(n10866) );
  OR U19040 ( .A(n10873), .B(n10874), .Z(n10872) );
  OR U19041 ( .A(n10875), .B(n10876), .Z(n10871) );
  NAND U19042 ( .A(n10877), .B(n10878), .Z(n10864) );
  OR U19043 ( .A(n10879), .B(n10880), .Z(n10878) );
  OR U19044 ( .A(n10881), .B(n10882), .Z(n10877) );
  NOR U19045 ( .A(n10883), .B(n10884), .Z(n10865) );
  ANDN U19046 ( .B(n10885), .A(n10886), .Z(n10859) );
  XNOR U19047 ( .A(n10852), .B(n10887), .Z(n10858) );
  XNOR U19048 ( .A(n10851), .B(n10853), .Z(n10887) );
  NAND U19049 ( .A(n10888), .B(n10889), .Z(n10853) );
  OR U19050 ( .A(n10890), .B(n10891), .Z(n10889) );
  OR U19051 ( .A(n10892), .B(n10893), .Z(n10888) );
  NAND U19052 ( .A(n10894), .B(n10895), .Z(n10851) );
  OR U19053 ( .A(n10896), .B(n10897), .Z(n10895) );
  OR U19054 ( .A(n10898), .B(n10899), .Z(n10894) );
  ANDN U19055 ( .B(n10900), .A(n10901), .Z(n10852) );
  IV U19056 ( .A(n10902), .Z(n10900) );
  ANDN U19057 ( .B(n10903), .A(n10904), .Z(n10844) );
  XOR U19058 ( .A(n10830), .B(n10905), .Z(n10842) );
  XOR U19059 ( .A(n10831), .B(n10832), .Z(n10905) );
  XOR U19060 ( .A(n10837), .B(n10906), .Z(n10832) );
  XOR U19061 ( .A(n10836), .B(n10839), .Z(n10906) );
  IV U19062 ( .A(n10838), .Z(n10839) );
  NAND U19063 ( .A(n10907), .B(n10908), .Z(n10838) );
  OR U19064 ( .A(n10909), .B(n10910), .Z(n10908) );
  OR U19065 ( .A(n10911), .B(n10912), .Z(n10907) );
  NAND U19066 ( .A(n10913), .B(n10914), .Z(n10836) );
  OR U19067 ( .A(n10915), .B(n10916), .Z(n10914) );
  OR U19068 ( .A(n10917), .B(n10918), .Z(n10913) );
  NOR U19069 ( .A(n10919), .B(n10920), .Z(n10837) );
  ANDN U19070 ( .B(n10921), .A(n10922), .Z(n10831) );
  IV U19071 ( .A(n10923), .Z(n10921) );
  XNOR U19072 ( .A(n10824), .B(n10924), .Z(n10830) );
  XNOR U19073 ( .A(n10823), .B(n10825), .Z(n10924) );
  NAND U19074 ( .A(n10925), .B(n10926), .Z(n10825) );
  OR U19075 ( .A(n10927), .B(n10928), .Z(n10926) );
  OR U19076 ( .A(n10929), .B(n10930), .Z(n10925) );
  NAND U19077 ( .A(n10931), .B(n10932), .Z(n10823) );
  OR U19078 ( .A(n10933), .B(n10934), .Z(n10932) );
  OR U19079 ( .A(n10935), .B(n10936), .Z(n10931) );
  ANDN U19080 ( .B(n10937), .A(n10938), .Z(n10824) );
  IV U19081 ( .A(n10939), .Z(n10937) );
  XNOR U19082 ( .A(n10904), .B(n10903), .Z(N64427) );
  XOR U19083 ( .A(n10923), .B(n10922), .Z(n10903) );
  XNOR U19084 ( .A(n10938), .B(n10939), .Z(n10922) );
  XNOR U19085 ( .A(n10933), .B(n10934), .Z(n10939) );
  XNOR U19086 ( .A(n10935), .B(n10936), .Z(n10934) );
  XNOR U19087 ( .A(y[7093]), .B(x[7093]), .Z(n10936) );
  XNOR U19088 ( .A(y[7094]), .B(x[7094]), .Z(n10935) );
  XNOR U19089 ( .A(y[7092]), .B(x[7092]), .Z(n10933) );
  XNOR U19090 ( .A(n10927), .B(n10928), .Z(n10938) );
  XNOR U19091 ( .A(y[7089]), .B(x[7089]), .Z(n10928) );
  XNOR U19092 ( .A(n10929), .B(n10930), .Z(n10927) );
  XNOR U19093 ( .A(y[7090]), .B(x[7090]), .Z(n10930) );
  XNOR U19094 ( .A(y[7091]), .B(x[7091]), .Z(n10929) );
  XNOR U19095 ( .A(n10920), .B(n10919), .Z(n10923) );
  XNOR U19096 ( .A(n10915), .B(n10916), .Z(n10919) );
  XNOR U19097 ( .A(y[7086]), .B(x[7086]), .Z(n10916) );
  XNOR U19098 ( .A(n10917), .B(n10918), .Z(n10915) );
  XNOR U19099 ( .A(y[7087]), .B(x[7087]), .Z(n10918) );
  XNOR U19100 ( .A(y[7088]), .B(x[7088]), .Z(n10917) );
  XNOR U19101 ( .A(n10909), .B(n10910), .Z(n10920) );
  XNOR U19102 ( .A(y[7083]), .B(x[7083]), .Z(n10910) );
  XNOR U19103 ( .A(n10911), .B(n10912), .Z(n10909) );
  XNOR U19104 ( .A(y[7084]), .B(x[7084]), .Z(n10912) );
  XNOR U19105 ( .A(y[7085]), .B(x[7085]), .Z(n10911) );
  XOR U19106 ( .A(n10885), .B(n10886), .Z(n10904) );
  XNOR U19107 ( .A(n10901), .B(n10902), .Z(n10886) );
  XNOR U19108 ( .A(n10896), .B(n10897), .Z(n10902) );
  XNOR U19109 ( .A(n10898), .B(n10899), .Z(n10897) );
  XNOR U19110 ( .A(y[7081]), .B(x[7081]), .Z(n10899) );
  XNOR U19111 ( .A(y[7082]), .B(x[7082]), .Z(n10898) );
  XNOR U19112 ( .A(y[7080]), .B(x[7080]), .Z(n10896) );
  XNOR U19113 ( .A(n10890), .B(n10891), .Z(n10901) );
  XNOR U19114 ( .A(y[7077]), .B(x[7077]), .Z(n10891) );
  XNOR U19115 ( .A(n10892), .B(n10893), .Z(n10890) );
  XNOR U19116 ( .A(y[7078]), .B(x[7078]), .Z(n10893) );
  XNOR U19117 ( .A(y[7079]), .B(x[7079]), .Z(n10892) );
  XOR U19118 ( .A(n10884), .B(n10883), .Z(n10885) );
  XNOR U19119 ( .A(n10879), .B(n10880), .Z(n10883) );
  XNOR U19120 ( .A(y[7074]), .B(x[7074]), .Z(n10880) );
  XNOR U19121 ( .A(n10881), .B(n10882), .Z(n10879) );
  XNOR U19122 ( .A(y[7075]), .B(x[7075]), .Z(n10882) );
  XNOR U19123 ( .A(y[7076]), .B(x[7076]), .Z(n10881) );
  XNOR U19124 ( .A(n10873), .B(n10874), .Z(n10884) );
  XNOR U19125 ( .A(y[7071]), .B(x[7071]), .Z(n10874) );
  XNOR U19126 ( .A(n10875), .B(n10876), .Z(n10873) );
  XNOR U19127 ( .A(y[7072]), .B(x[7072]), .Z(n10876) );
  XNOR U19128 ( .A(y[7073]), .B(x[7073]), .Z(n10875) );
  NAND U19129 ( .A(n10940), .B(n10941), .Z(N64418) );
  NANDN U19130 ( .A(n10942), .B(n10943), .Z(n10941) );
  OR U19131 ( .A(n10944), .B(n10945), .Z(n10943) );
  NAND U19132 ( .A(n10944), .B(n10945), .Z(n10940) );
  XOR U19133 ( .A(n10944), .B(n10946), .Z(N64417) );
  XNOR U19134 ( .A(n10942), .B(n10945), .Z(n10946) );
  AND U19135 ( .A(n10947), .B(n10948), .Z(n10945) );
  NANDN U19136 ( .A(n10949), .B(n10950), .Z(n10948) );
  NANDN U19137 ( .A(n10951), .B(n10952), .Z(n10950) );
  NANDN U19138 ( .A(n10952), .B(n10951), .Z(n10947) );
  NAND U19139 ( .A(n10953), .B(n10954), .Z(n10942) );
  NANDN U19140 ( .A(n10955), .B(n10956), .Z(n10954) );
  OR U19141 ( .A(n10957), .B(n10958), .Z(n10956) );
  NAND U19142 ( .A(n10958), .B(n10957), .Z(n10953) );
  AND U19143 ( .A(n10959), .B(n10960), .Z(n10944) );
  NANDN U19144 ( .A(n10961), .B(n10962), .Z(n10960) );
  NANDN U19145 ( .A(n10963), .B(n10964), .Z(n10962) );
  NANDN U19146 ( .A(n10964), .B(n10963), .Z(n10959) );
  XOR U19147 ( .A(n10958), .B(n10965), .Z(N64416) );
  XOR U19148 ( .A(n10955), .B(n10957), .Z(n10965) );
  XNOR U19149 ( .A(n10951), .B(n10966), .Z(n10957) );
  XNOR U19150 ( .A(n10949), .B(n10952), .Z(n10966) );
  NAND U19151 ( .A(n10967), .B(n10968), .Z(n10952) );
  NAND U19152 ( .A(n10969), .B(n10970), .Z(n10968) );
  OR U19153 ( .A(n10971), .B(n10972), .Z(n10969) );
  NANDN U19154 ( .A(n10973), .B(n10971), .Z(n10967) );
  IV U19155 ( .A(n10972), .Z(n10973) );
  NAND U19156 ( .A(n10974), .B(n10975), .Z(n10949) );
  NAND U19157 ( .A(n10976), .B(n10977), .Z(n10975) );
  NANDN U19158 ( .A(n10978), .B(n10979), .Z(n10976) );
  NANDN U19159 ( .A(n10979), .B(n10978), .Z(n10974) );
  AND U19160 ( .A(n10980), .B(n10981), .Z(n10951) );
  NAND U19161 ( .A(n10982), .B(n10983), .Z(n10981) );
  OR U19162 ( .A(n10984), .B(n10985), .Z(n10982) );
  NANDN U19163 ( .A(n10986), .B(n10984), .Z(n10980) );
  NAND U19164 ( .A(n10987), .B(n10988), .Z(n10955) );
  NANDN U19165 ( .A(n10989), .B(n10990), .Z(n10988) );
  OR U19166 ( .A(n10991), .B(n10992), .Z(n10990) );
  NANDN U19167 ( .A(n10993), .B(n10991), .Z(n10987) );
  IV U19168 ( .A(n10992), .Z(n10993) );
  XNOR U19169 ( .A(n10963), .B(n10994), .Z(n10958) );
  XNOR U19170 ( .A(n10961), .B(n10964), .Z(n10994) );
  NAND U19171 ( .A(n10995), .B(n10996), .Z(n10964) );
  NAND U19172 ( .A(n10997), .B(n10998), .Z(n10996) );
  OR U19173 ( .A(n10999), .B(n11000), .Z(n10997) );
  NANDN U19174 ( .A(n11001), .B(n10999), .Z(n10995) );
  IV U19175 ( .A(n11000), .Z(n11001) );
  NAND U19176 ( .A(n11002), .B(n11003), .Z(n10961) );
  NAND U19177 ( .A(n11004), .B(n11005), .Z(n11003) );
  NANDN U19178 ( .A(n11006), .B(n11007), .Z(n11004) );
  NANDN U19179 ( .A(n11007), .B(n11006), .Z(n11002) );
  AND U19180 ( .A(n11008), .B(n11009), .Z(n10963) );
  NAND U19181 ( .A(n11010), .B(n11011), .Z(n11009) );
  OR U19182 ( .A(n11012), .B(n11013), .Z(n11010) );
  NANDN U19183 ( .A(n11014), .B(n11012), .Z(n11008) );
  XNOR U19184 ( .A(n10989), .B(n11015), .Z(N64415) );
  XOR U19185 ( .A(n10991), .B(n10992), .Z(n11015) );
  XNOR U19186 ( .A(n11005), .B(n11016), .Z(n10992) );
  XOR U19187 ( .A(n11006), .B(n11007), .Z(n11016) );
  XOR U19188 ( .A(n11012), .B(n11017), .Z(n11007) );
  XOR U19189 ( .A(n11011), .B(n11014), .Z(n11017) );
  IV U19190 ( .A(n11013), .Z(n11014) );
  NAND U19191 ( .A(n11018), .B(n11019), .Z(n11013) );
  OR U19192 ( .A(n11020), .B(n11021), .Z(n11019) );
  OR U19193 ( .A(n11022), .B(n11023), .Z(n11018) );
  NAND U19194 ( .A(n11024), .B(n11025), .Z(n11011) );
  OR U19195 ( .A(n11026), .B(n11027), .Z(n11025) );
  OR U19196 ( .A(n11028), .B(n11029), .Z(n11024) );
  NOR U19197 ( .A(n11030), .B(n11031), .Z(n11012) );
  ANDN U19198 ( .B(n11032), .A(n11033), .Z(n11006) );
  XNOR U19199 ( .A(n10999), .B(n11034), .Z(n11005) );
  XNOR U19200 ( .A(n10998), .B(n11000), .Z(n11034) );
  NAND U19201 ( .A(n11035), .B(n11036), .Z(n11000) );
  OR U19202 ( .A(n11037), .B(n11038), .Z(n11036) );
  OR U19203 ( .A(n11039), .B(n11040), .Z(n11035) );
  NAND U19204 ( .A(n11041), .B(n11042), .Z(n10998) );
  OR U19205 ( .A(n11043), .B(n11044), .Z(n11042) );
  OR U19206 ( .A(n11045), .B(n11046), .Z(n11041) );
  ANDN U19207 ( .B(n11047), .A(n11048), .Z(n10999) );
  IV U19208 ( .A(n11049), .Z(n11047) );
  ANDN U19209 ( .B(n11050), .A(n11051), .Z(n10991) );
  XOR U19210 ( .A(n10977), .B(n11052), .Z(n10989) );
  XOR U19211 ( .A(n10978), .B(n10979), .Z(n11052) );
  XOR U19212 ( .A(n10984), .B(n11053), .Z(n10979) );
  XOR U19213 ( .A(n10983), .B(n10986), .Z(n11053) );
  IV U19214 ( .A(n10985), .Z(n10986) );
  NAND U19215 ( .A(n11054), .B(n11055), .Z(n10985) );
  OR U19216 ( .A(n11056), .B(n11057), .Z(n11055) );
  OR U19217 ( .A(n11058), .B(n11059), .Z(n11054) );
  NAND U19218 ( .A(n11060), .B(n11061), .Z(n10983) );
  OR U19219 ( .A(n11062), .B(n11063), .Z(n11061) );
  OR U19220 ( .A(n11064), .B(n11065), .Z(n11060) );
  NOR U19221 ( .A(n11066), .B(n11067), .Z(n10984) );
  ANDN U19222 ( .B(n11068), .A(n11069), .Z(n10978) );
  IV U19223 ( .A(n11070), .Z(n11068) );
  XNOR U19224 ( .A(n10971), .B(n11071), .Z(n10977) );
  XNOR U19225 ( .A(n10970), .B(n10972), .Z(n11071) );
  NAND U19226 ( .A(n11072), .B(n11073), .Z(n10972) );
  OR U19227 ( .A(n11074), .B(n11075), .Z(n11073) );
  OR U19228 ( .A(n11076), .B(n11077), .Z(n11072) );
  NAND U19229 ( .A(n11078), .B(n11079), .Z(n10970) );
  OR U19230 ( .A(n11080), .B(n11081), .Z(n11079) );
  OR U19231 ( .A(n11082), .B(n11083), .Z(n11078) );
  ANDN U19232 ( .B(n11084), .A(n11085), .Z(n10971) );
  IV U19233 ( .A(n11086), .Z(n11084) );
  XNOR U19234 ( .A(n11051), .B(n11050), .Z(N64414) );
  XOR U19235 ( .A(n11070), .B(n11069), .Z(n11050) );
  XNOR U19236 ( .A(n11085), .B(n11086), .Z(n11069) );
  XNOR U19237 ( .A(n11080), .B(n11081), .Z(n11086) );
  XNOR U19238 ( .A(n11082), .B(n11083), .Z(n11081) );
  XNOR U19239 ( .A(y[7069]), .B(x[7069]), .Z(n11083) );
  XNOR U19240 ( .A(y[7070]), .B(x[7070]), .Z(n11082) );
  XNOR U19241 ( .A(y[7068]), .B(x[7068]), .Z(n11080) );
  XNOR U19242 ( .A(n11074), .B(n11075), .Z(n11085) );
  XNOR U19243 ( .A(y[7065]), .B(x[7065]), .Z(n11075) );
  XNOR U19244 ( .A(n11076), .B(n11077), .Z(n11074) );
  XNOR U19245 ( .A(y[7066]), .B(x[7066]), .Z(n11077) );
  XNOR U19246 ( .A(y[7067]), .B(x[7067]), .Z(n11076) );
  XNOR U19247 ( .A(n11067), .B(n11066), .Z(n11070) );
  XNOR U19248 ( .A(n11062), .B(n11063), .Z(n11066) );
  XNOR U19249 ( .A(y[7062]), .B(x[7062]), .Z(n11063) );
  XNOR U19250 ( .A(n11064), .B(n11065), .Z(n11062) );
  XNOR U19251 ( .A(y[7063]), .B(x[7063]), .Z(n11065) );
  XNOR U19252 ( .A(y[7064]), .B(x[7064]), .Z(n11064) );
  XNOR U19253 ( .A(n11056), .B(n11057), .Z(n11067) );
  XNOR U19254 ( .A(y[7059]), .B(x[7059]), .Z(n11057) );
  XNOR U19255 ( .A(n11058), .B(n11059), .Z(n11056) );
  XNOR U19256 ( .A(y[7060]), .B(x[7060]), .Z(n11059) );
  XNOR U19257 ( .A(y[7061]), .B(x[7061]), .Z(n11058) );
  XOR U19258 ( .A(n11032), .B(n11033), .Z(n11051) );
  XNOR U19259 ( .A(n11048), .B(n11049), .Z(n11033) );
  XNOR U19260 ( .A(n11043), .B(n11044), .Z(n11049) );
  XNOR U19261 ( .A(n11045), .B(n11046), .Z(n11044) );
  XNOR U19262 ( .A(y[7057]), .B(x[7057]), .Z(n11046) );
  XNOR U19263 ( .A(y[7058]), .B(x[7058]), .Z(n11045) );
  XNOR U19264 ( .A(y[7056]), .B(x[7056]), .Z(n11043) );
  XNOR U19265 ( .A(n11037), .B(n11038), .Z(n11048) );
  XNOR U19266 ( .A(y[7053]), .B(x[7053]), .Z(n11038) );
  XNOR U19267 ( .A(n11039), .B(n11040), .Z(n11037) );
  XNOR U19268 ( .A(y[7054]), .B(x[7054]), .Z(n11040) );
  XNOR U19269 ( .A(y[7055]), .B(x[7055]), .Z(n11039) );
  XOR U19270 ( .A(n11031), .B(n11030), .Z(n11032) );
  XNOR U19271 ( .A(n11026), .B(n11027), .Z(n11030) );
  XNOR U19272 ( .A(y[7050]), .B(x[7050]), .Z(n11027) );
  XNOR U19273 ( .A(n11028), .B(n11029), .Z(n11026) );
  XNOR U19274 ( .A(y[7051]), .B(x[7051]), .Z(n11029) );
  XNOR U19275 ( .A(y[7052]), .B(x[7052]), .Z(n11028) );
  XNOR U19276 ( .A(n11020), .B(n11021), .Z(n11031) );
  XNOR U19277 ( .A(y[7047]), .B(x[7047]), .Z(n11021) );
  XNOR U19278 ( .A(n11022), .B(n11023), .Z(n11020) );
  XNOR U19279 ( .A(y[7048]), .B(x[7048]), .Z(n11023) );
  XNOR U19280 ( .A(y[7049]), .B(x[7049]), .Z(n11022) );
  NAND U19281 ( .A(n11087), .B(n11088), .Z(N64405) );
  NANDN U19282 ( .A(n11089), .B(n11090), .Z(n11088) );
  OR U19283 ( .A(n11091), .B(n11092), .Z(n11090) );
  NAND U19284 ( .A(n11091), .B(n11092), .Z(n11087) );
  XOR U19285 ( .A(n11091), .B(n11093), .Z(N64404) );
  XNOR U19286 ( .A(n11089), .B(n11092), .Z(n11093) );
  AND U19287 ( .A(n11094), .B(n11095), .Z(n11092) );
  NANDN U19288 ( .A(n11096), .B(n11097), .Z(n11095) );
  NANDN U19289 ( .A(n11098), .B(n11099), .Z(n11097) );
  NANDN U19290 ( .A(n11099), .B(n11098), .Z(n11094) );
  NAND U19291 ( .A(n11100), .B(n11101), .Z(n11089) );
  NANDN U19292 ( .A(n11102), .B(n11103), .Z(n11101) );
  OR U19293 ( .A(n11104), .B(n11105), .Z(n11103) );
  NAND U19294 ( .A(n11105), .B(n11104), .Z(n11100) );
  AND U19295 ( .A(n11106), .B(n11107), .Z(n11091) );
  NANDN U19296 ( .A(n11108), .B(n11109), .Z(n11107) );
  NANDN U19297 ( .A(n11110), .B(n11111), .Z(n11109) );
  NANDN U19298 ( .A(n11111), .B(n11110), .Z(n11106) );
  XOR U19299 ( .A(n11105), .B(n11112), .Z(N64403) );
  XOR U19300 ( .A(n11102), .B(n11104), .Z(n11112) );
  XNOR U19301 ( .A(n11098), .B(n11113), .Z(n11104) );
  XNOR U19302 ( .A(n11096), .B(n11099), .Z(n11113) );
  NAND U19303 ( .A(n11114), .B(n11115), .Z(n11099) );
  NAND U19304 ( .A(n11116), .B(n11117), .Z(n11115) );
  OR U19305 ( .A(n11118), .B(n11119), .Z(n11116) );
  NANDN U19306 ( .A(n11120), .B(n11118), .Z(n11114) );
  IV U19307 ( .A(n11119), .Z(n11120) );
  NAND U19308 ( .A(n11121), .B(n11122), .Z(n11096) );
  NAND U19309 ( .A(n11123), .B(n11124), .Z(n11122) );
  NANDN U19310 ( .A(n11125), .B(n11126), .Z(n11123) );
  NANDN U19311 ( .A(n11126), .B(n11125), .Z(n11121) );
  AND U19312 ( .A(n11127), .B(n11128), .Z(n11098) );
  NAND U19313 ( .A(n11129), .B(n11130), .Z(n11128) );
  OR U19314 ( .A(n11131), .B(n11132), .Z(n11129) );
  NANDN U19315 ( .A(n11133), .B(n11131), .Z(n11127) );
  NAND U19316 ( .A(n11134), .B(n11135), .Z(n11102) );
  NANDN U19317 ( .A(n11136), .B(n11137), .Z(n11135) );
  OR U19318 ( .A(n11138), .B(n11139), .Z(n11137) );
  NANDN U19319 ( .A(n11140), .B(n11138), .Z(n11134) );
  IV U19320 ( .A(n11139), .Z(n11140) );
  XNOR U19321 ( .A(n11110), .B(n11141), .Z(n11105) );
  XNOR U19322 ( .A(n11108), .B(n11111), .Z(n11141) );
  NAND U19323 ( .A(n11142), .B(n11143), .Z(n11111) );
  NAND U19324 ( .A(n11144), .B(n11145), .Z(n11143) );
  OR U19325 ( .A(n11146), .B(n11147), .Z(n11144) );
  NANDN U19326 ( .A(n11148), .B(n11146), .Z(n11142) );
  IV U19327 ( .A(n11147), .Z(n11148) );
  NAND U19328 ( .A(n11149), .B(n11150), .Z(n11108) );
  NAND U19329 ( .A(n11151), .B(n11152), .Z(n11150) );
  NANDN U19330 ( .A(n11153), .B(n11154), .Z(n11151) );
  NANDN U19331 ( .A(n11154), .B(n11153), .Z(n11149) );
  AND U19332 ( .A(n11155), .B(n11156), .Z(n11110) );
  NAND U19333 ( .A(n11157), .B(n11158), .Z(n11156) );
  OR U19334 ( .A(n11159), .B(n11160), .Z(n11157) );
  NANDN U19335 ( .A(n11161), .B(n11159), .Z(n11155) );
  XNOR U19336 ( .A(n11136), .B(n11162), .Z(N64402) );
  XOR U19337 ( .A(n11138), .B(n11139), .Z(n11162) );
  XNOR U19338 ( .A(n11152), .B(n11163), .Z(n11139) );
  XOR U19339 ( .A(n11153), .B(n11154), .Z(n11163) );
  XOR U19340 ( .A(n11159), .B(n11164), .Z(n11154) );
  XOR U19341 ( .A(n11158), .B(n11161), .Z(n11164) );
  IV U19342 ( .A(n11160), .Z(n11161) );
  NAND U19343 ( .A(n11165), .B(n11166), .Z(n11160) );
  OR U19344 ( .A(n11167), .B(n11168), .Z(n11166) );
  OR U19345 ( .A(n11169), .B(n11170), .Z(n11165) );
  NAND U19346 ( .A(n11171), .B(n11172), .Z(n11158) );
  OR U19347 ( .A(n11173), .B(n11174), .Z(n11172) );
  OR U19348 ( .A(n11175), .B(n11176), .Z(n11171) );
  NOR U19349 ( .A(n11177), .B(n11178), .Z(n11159) );
  ANDN U19350 ( .B(n11179), .A(n11180), .Z(n11153) );
  XNOR U19351 ( .A(n11146), .B(n11181), .Z(n11152) );
  XNOR U19352 ( .A(n11145), .B(n11147), .Z(n11181) );
  NAND U19353 ( .A(n11182), .B(n11183), .Z(n11147) );
  OR U19354 ( .A(n11184), .B(n11185), .Z(n11183) );
  OR U19355 ( .A(n11186), .B(n11187), .Z(n11182) );
  NAND U19356 ( .A(n11188), .B(n11189), .Z(n11145) );
  OR U19357 ( .A(n11190), .B(n11191), .Z(n11189) );
  OR U19358 ( .A(n11192), .B(n11193), .Z(n11188) );
  ANDN U19359 ( .B(n11194), .A(n11195), .Z(n11146) );
  IV U19360 ( .A(n11196), .Z(n11194) );
  ANDN U19361 ( .B(n11197), .A(n11198), .Z(n11138) );
  XOR U19362 ( .A(n11124), .B(n11199), .Z(n11136) );
  XOR U19363 ( .A(n11125), .B(n11126), .Z(n11199) );
  XOR U19364 ( .A(n11131), .B(n11200), .Z(n11126) );
  XOR U19365 ( .A(n11130), .B(n11133), .Z(n11200) );
  IV U19366 ( .A(n11132), .Z(n11133) );
  NAND U19367 ( .A(n11201), .B(n11202), .Z(n11132) );
  OR U19368 ( .A(n11203), .B(n11204), .Z(n11202) );
  OR U19369 ( .A(n11205), .B(n11206), .Z(n11201) );
  NAND U19370 ( .A(n11207), .B(n11208), .Z(n11130) );
  OR U19371 ( .A(n11209), .B(n11210), .Z(n11208) );
  OR U19372 ( .A(n11211), .B(n11212), .Z(n11207) );
  NOR U19373 ( .A(n11213), .B(n11214), .Z(n11131) );
  ANDN U19374 ( .B(n11215), .A(n11216), .Z(n11125) );
  IV U19375 ( .A(n11217), .Z(n11215) );
  XNOR U19376 ( .A(n11118), .B(n11218), .Z(n11124) );
  XNOR U19377 ( .A(n11117), .B(n11119), .Z(n11218) );
  NAND U19378 ( .A(n11219), .B(n11220), .Z(n11119) );
  OR U19379 ( .A(n11221), .B(n11222), .Z(n11220) );
  OR U19380 ( .A(n11223), .B(n11224), .Z(n11219) );
  NAND U19381 ( .A(n11225), .B(n11226), .Z(n11117) );
  OR U19382 ( .A(n11227), .B(n11228), .Z(n11226) );
  OR U19383 ( .A(n11229), .B(n11230), .Z(n11225) );
  ANDN U19384 ( .B(n11231), .A(n11232), .Z(n11118) );
  IV U19385 ( .A(n11233), .Z(n11231) );
  XNOR U19386 ( .A(n11198), .B(n11197), .Z(N64401) );
  XOR U19387 ( .A(n11217), .B(n11216), .Z(n11197) );
  XNOR U19388 ( .A(n11232), .B(n11233), .Z(n11216) );
  XNOR U19389 ( .A(n11227), .B(n11228), .Z(n11233) );
  XNOR U19390 ( .A(n11229), .B(n11230), .Z(n11228) );
  XNOR U19391 ( .A(y[7045]), .B(x[7045]), .Z(n11230) );
  XNOR U19392 ( .A(y[7046]), .B(x[7046]), .Z(n11229) );
  XNOR U19393 ( .A(y[7044]), .B(x[7044]), .Z(n11227) );
  XNOR U19394 ( .A(n11221), .B(n11222), .Z(n11232) );
  XNOR U19395 ( .A(y[7041]), .B(x[7041]), .Z(n11222) );
  XNOR U19396 ( .A(n11223), .B(n11224), .Z(n11221) );
  XNOR U19397 ( .A(y[7042]), .B(x[7042]), .Z(n11224) );
  XNOR U19398 ( .A(y[7043]), .B(x[7043]), .Z(n11223) );
  XNOR U19399 ( .A(n11214), .B(n11213), .Z(n11217) );
  XNOR U19400 ( .A(n11209), .B(n11210), .Z(n11213) );
  XNOR U19401 ( .A(y[7038]), .B(x[7038]), .Z(n11210) );
  XNOR U19402 ( .A(n11211), .B(n11212), .Z(n11209) );
  XNOR U19403 ( .A(y[7039]), .B(x[7039]), .Z(n11212) );
  XNOR U19404 ( .A(y[7040]), .B(x[7040]), .Z(n11211) );
  XNOR U19405 ( .A(n11203), .B(n11204), .Z(n11214) );
  XNOR U19406 ( .A(y[7035]), .B(x[7035]), .Z(n11204) );
  XNOR U19407 ( .A(n11205), .B(n11206), .Z(n11203) );
  XNOR U19408 ( .A(y[7036]), .B(x[7036]), .Z(n11206) );
  XNOR U19409 ( .A(y[7037]), .B(x[7037]), .Z(n11205) );
  XOR U19410 ( .A(n11179), .B(n11180), .Z(n11198) );
  XNOR U19411 ( .A(n11195), .B(n11196), .Z(n11180) );
  XNOR U19412 ( .A(n11190), .B(n11191), .Z(n11196) );
  XNOR U19413 ( .A(n11192), .B(n11193), .Z(n11191) );
  XNOR U19414 ( .A(y[7033]), .B(x[7033]), .Z(n11193) );
  XNOR U19415 ( .A(y[7034]), .B(x[7034]), .Z(n11192) );
  XNOR U19416 ( .A(y[7032]), .B(x[7032]), .Z(n11190) );
  XNOR U19417 ( .A(n11184), .B(n11185), .Z(n11195) );
  XNOR U19418 ( .A(y[7029]), .B(x[7029]), .Z(n11185) );
  XNOR U19419 ( .A(n11186), .B(n11187), .Z(n11184) );
  XNOR U19420 ( .A(y[7030]), .B(x[7030]), .Z(n11187) );
  XNOR U19421 ( .A(y[7031]), .B(x[7031]), .Z(n11186) );
  XOR U19422 ( .A(n11178), .B(n11177), .Z(n11179) );
  XNOR U19423 ( .A(n11173), .B(n11174), .Z(n11177) );
  XNOR U19424 ( .A(y[7026]), .B(x[7026]), .Z(n11174) );
  XNOR U19425 ( .A(n11175), .B(n11176), .Z(n11173) );
  XNOR U19426 ( .A(y[7027]), .B(x[7027]), .Z(n11176) );
  XNOR U19427 ( .A(y[7028]), .B(x[7028]), .Z(n11175) );
  XNOR U19428 ( .A(n11167), .B(n11168), .Z(n11178) );
  XNOR U19429 ( .A(y[7023]), .B(x[7023]), .Z(n11168) );
  XNOR U19430 ( .A(n11169), .B(n11170), .Z(n11167) );
  XNOR U19431 ( .A(y[7024]), .B(x[7024]), .Z(n11170) );
  XNOR U19432 ( .A(y[7025]), .B(x[7025]), .Z(n11169) );
  NAND U19433 ( .A(n11234), .B(n11235), .Z(N64392) );
  NANDN U19434 ( .A(n11236), .B(n11237), .Z(n11235) );
  OR U19435 ( .A(n11238), .B(n11239), .Z(n11237) );
  NAND U19436 ( .A(n11238), .B(n11239), .Z(n11234) );
  XOR U19437 ( .A(n11238), .B(n11240), .Z(N64391) );
  XNOR U19438 ( .A(n11236), .B(n11239), .Z(n11240) );
  AND U19439 ( .A(n11241), .B(n11242), .Z(n11239) );
  NANDN U19440 ( .A(n11243), .B(n11244), .Z(n11242) );
  NANDN U19441 ( .A(n11245), .B(n11246), .Z(n11244) );
  NANDN U19442 ( .A(n11246), .B(n11245), .Z(n11241) );
  NAND U19443 ( .A(n11247), .B(n11248), .Z(n11236) );
  NANDN U19444 ( .A(n11249), .B(n11250), .Z(n11248) );
  OR U19445 ( .A(n11251), .B(n11252), .Z(n11250) );
  NAND U19446 ( .A(n11252), .B(n11251), .Z(n11247) );
  AND U19447 ( .A(n11253), .B(n11254), .Z(n11238) );
  NANDN U19448 ( .A(n11255), .B(n11256), .Z(n11254) );
  NANDN U19449 ( .A(n11257), .B(n11258), .Z(n11256) );
  NANDN U19450 ( .A(n11258), .B(n11257), .Z(n11253) );
  XOR U19451 ( .A(n11252), .B(n11259), .Z(N64390) );
  XOR U19452 ( .A(n11249), .B(n11251), .Z(n11259) );
  XNOR U19453 ( .A(n11245), .B(n11260), .Z(n11251) );
  XNOR U19454 ( .A(n11243), .B(n11246), .Z(n11260) );
  NAND U19455 ( .A(n11261), .B(n11262), .Z(n11246) );
  NAND U19456 ( .A(n11263), .B(n11264), .Z(n11262) );
  OR U19457 ( .A(n11265), .B(n11266), .Z(n11263) );
  NANDN U19458 ( .A(n11267), .B(n11265), .Z(n11261) );
  IV U19459 ( .A(n11266), .Z(n11267) );
  NAND U19460 ( .A(n11268), .B(n11269), .Z(n11243) );
  NAND U19461 ( .A(n11270), .B(n11271), .Z(n11269) );
  NANDN U19462 ( .A(n11272), .B(n11273), .Z(n11270) );
  NANDN U19463 ( .A(n11273), .B(n11272), .Z(n11268) );
  AND U19464 ( .A(n11274), .B(n11275), .Z(n11245) );
  NAND U19465 ( .A(n11276), .B(n11277), .Z(n11275) );
  OR U19466 ( .A(n11278), .B(n11279), .Z(n11276) );
  NANDN U19467 ( .A(n11280), .B(n11278), .Z(n11274) );
  NAND U19468 ( .A(n11281), .B(n11282), .Z(n11249) );
  NANDN U19469 ( .A(n11283), .B(n11284), .Z(n11282) );
  OR U19470 ( .A(n11285), .B(n11286), .Z(n11284) );
  NANDN U19471 ( .A(n11287), .B(n11285), .Z(n11281) );
  IV U19472 ( .A(n11286), .Z(n11287) );
  XNOR U19473 ( .A(n11257), .B(n11288), .Z(n11252) );
  XNOR U19474 ( .A(n11255), .B(n11258), .Z(n11288) );
  NAND U19475 ( .A(n11289), .B(n11290), .Z(n11258) );
  NAND U19476 ( .A(n11291), .B(n11292), .Z(n11290) );
  OR U19477 ( .A(n11293), .B(n11294), .Z(n11291) );
  NANDN U19478 ( .A(n11295), .B(n11293), .Z(n11289) );
  IV U19479 ( .A(n11294), .Z(n11295) );
  NAND U19480 ( .A(n11296), .B(n11297), .Z(n11255) );
  NAND U19481 ( .A(n11298), .B(n11299), .Z(n11297) );
  NANDN U19482 ( .A(n11300), .B(n11301), .Z(n11298) );
  NANDN U19483 ( .A(n11301), .B(n11300), .Z(n11296) );
  AND U19484 ( .A(n11302), .B(n11303), .Z(n11257) );
  NAND U19485 ( .A(n11304), .B(n11305), .Z(n11303) );
  OR U19486 ( .A(n11306), .B(n11307), .Z(n11304) );
  NANDN U19487 ( .A(n11308), .B(n11306), .Z(n11302) );
  XNOR U19488 ( .A(n11283), .B(n11309), .Z(N64389) );
  XOR U19489 ( .A(n11285), .B(n11286), .Z(n11309) );
  XNOR U19490 ( .A(n11299), .B(n11310), .Z(n11286) );
  XOR U19491 ( .A(n11300), .B(n11301), .Z(n11310) );
  XOR U19492 ( .A(n11306), .B(n11311), .Z(n11301) );
  XOR U19493 ( .A(n11305), .B(n11308), .Z(n11311) );
  IV U19494 ( .A(n11307), .Z(n11308) );
  NAND U19495 ( .A(n11312), .B(n11313), .Z(n11307) );
  OR U19496 ( .A(n11314), .B(n11315), .Z(n11313) );
  OR U19497 ( .A(n11316), .B(n11317), .Z(n11312) );
  NAND U19498 ( .A(n11318), .B(n11319), .Z(n11305) );
  OR U19499 ( .A(n11320), .B(n11321), .Z(n11319) );
  OR U19500 ( .A(n11322), .B(n11323), .Z(n11318) );
  NOR U19501 ( .A(n11324), .B(n11325), .Z(n11306) );
  ANDN U19502 ( .B(n11326), .A(n11327), .Z(n11300) );
  XNOR U19503 ( .A(n11293), .B(n11328), .Z(n11299) );
  XNOR U19504 ( .A(n11292), .B(n11294), .Z(n11328) );
  NAND U19505 ( .A(n11329), .B(n11330), .Z(n11294) );
  OR U19506 ( .A(n11331), .B(n11332), .Z(n11330) );
  OR U19507 ( .A(n11333), .B(n11334), .Z(n11329) );
  NAND U19508 ( .A(n11335), .B(n11336), .Z(n11292) );
  OR U19509 ( .A(n11337), .B(n11338), .Z(n11336) );
  OR U19510 ( .A(n11339), .B(n11340), .Z(n11335) );
  ANDN U19511 ( .B(n11341), .A(n11342), .Z(n11293) );
  IV U19512 ( .A(n11343), .Z(n11341) );
  ANDN U19513 ( .B(n11344), .A(n11345), .Z(n11285) );
  XOR U19514 ( .A(n11271), .B(n11346), .Z(n11283) );
  XOR U19515 ( .A(n11272), .B(n11273), .Z(n11346) );
  XOR U19516 ( .A(n11278), .B(n11347), .Z(n11273) );
  XOR U19517 ( .A(n11277), .B(n11280), .Z(n11347) );
  IV U19518 ( .A(n11279), .Z(n11280) );
  NAND U19519 ( .A(n11348), .B(n11349), .Z(n11279) );
  OR U19520 ( .A(n11350), .B(n11351), .Z(n11349) );
  OR U19521 ( .A(n11352), .B(n11353), .Z(n11348) );
  NAND U19522 ( .A(n11354), .B(n11355), .Z(n11277) );
  OR U19523 ( .A(n11356), .B(n11357), .Z(n11355) );
  OR U19524 ( .A(n11358), .B(n11359), .Z(n11354) );
  NOR U19525 ( .A(n11360), .B(n11361), .Z(n11278) );
  ANDN U19526 ( .B(n11362), .A(n11363), .Z(n11272) );
  IV U19527 ( .A(n11364), .Z(n11362) );
  XNOR U19528 ( .A(n11265), .B(n11365), .Z(n11271) );
  XNOR U19529 ( .A(n11264), .B(n11266), .Z(n11365) );
  NAND U19530 ( .A(n11366), .B(n11367), .Z(n11266) );
  OR U19531 ( .A(n11368), .B(n11369), .Z(n11367) );
  OR U19532 ( .A(n11370), .B(n11371), .Z(n11366) );
  NAND U19533 ( .A(n11372), .B(n11373), .Z(n11264) );
  OR U19534 ( .A(n11374), .B(n11375), .Z(n11373) );
  OR U19535 ( .A(n11376), .B(n11377), .Z(n11372) );
  ANDN U19536 ( .B(n11378), .A(n11379), .Z(n11265) );
  IV U19537 ( .A(n11380), .Z(n11378) );
  XNOR U19538 ( .A(n11345), .B(n11344), .Z(N64388) );
  XOR U19539 ( .A(n11364), .B(n11363), .Z(n11344) );
  XNOR U19540 ( .A(n11379), .B(n11380), .Z(n11363) );
  XNOR U19541 ( .A(n11374), .B(n11375), .Z(n11380) );
  XNOR U19542 ( .A(n11376), .B(n11377), .Z(n11375) );
  XNOR U19543 ( .A(y[7021]), .B(x[7021]), .Z(n11377) );
  XNOR U19544 ( .A(y[7022]), .B(x[7022]), .Z(n11376) );
  XNOR U19545 ( .A(y[7020]), .B(x[7020]), .Z(n11374) );
  XNOR U19546 ( .A(n11368), .B(n11369), .Z(n11379) );
  XNOR U19547 ( .A(y[7017]), .B(x[7017]), .Z(n11369) );
  XNOR U19548 ( .A(n11370), .B(n11371), .Z(n11368) );
  XNOR U19549 ( .A(y[7018]), .B(x[7018]), .Z(n11371) );
  XNOR U19550 ( .A(y[7019]), .B(x[7019]), .Z(n11370) );
  XNOR U19551 ( .A(n11361), .B(n11360), .Z(n11364) );
  XNOR U19552 ( .A(n11356), .B(n11357), .Z(n11360) );
  XNOR U19553 ( .A(y[7014]), .B(x[7014]), .Z(n11357) );
  XNOR U19554 ( .A(n11358), .B(n11359), .Z(n11356) );
  XNOR U19555 ( .A(y[7015]), .B(x[7015]), .Z(n11359) );
  XNOR U19556 ( .A(y[7016]), .B(x[7016]), .Z(n11358) );
  XNOR U19557 ( .A(n11350), .B(n11351), .Z(n11361) );
  XNOR U19558 ( .A(y[7011]), .B(x[7011]), .Z(n11351) );
  XNOR U19559 ( .A(n11352), .B(n11353), .Z(n11350) );
  XNOR U19560 ( .A(y[7012]), .B(x[7012]), .Z(n11353) );
  XNOR U19561 ( .A(y[7013]), .B(x[7013]), .Z(n11352) );
  XOR U19562 ( .A(n11326), .B(n11327), .Z(n11345) );
  XNOR U19563 ( .A(n11342), .B(n11343), .Z(n11327) );
  XNOR U19564 ( .A(n11337), .B(n11338), .Z(n11343) );
  XNOR U19565 ( .A(n11339), .B(n11340), .Z(n11338) );
  XNOR U19566 ( .A(y[7009]), .B(x[7009]), .Z(n11340) );
  XNOR U19567 ( .A(y[7010]), .B(x[7010]), .Z(n11339) );
  XNOR U19568 ( .A(y[7008]), .B(x[7008]), .Z(n11337) );
  XNOR U19569 ( .A(n11331), .B(n11332), .Z(n11342) );
  XNOR U19570 ( .A(y[7005]), .B(x[7005]), .Z(n11332) );
  XNOR U19571 ( .A(n11333), .B(n11334), .Z(n11331) );
  XNOR U19572 ( .A(y[7006]), .B(x[7006]), .Z(n11334) );
  XNOR U19573 ( .A(y[7007]), .B(x[7007]), .Z(n11333) );
  XOR U19574 ( .A(n11325), .B(n11324), .Z(n11326) );
  XNOR U19575 ( .A(n11320), .B(n11321), .Z(n11324) );
  XNOR U19576 ( .A(y[7002]), .B(x[7002]), .Z(n11321) );
  XNOR U19577 ( .A(n11322), .B(n11323), .Z(n11320) );
  XNOR U19578 ( .A(y[7003]), .B(x[7003]), .Z(n11323) );
  XNOR U19579 ( .A(y[7004]), .B(x[7004]), .Z(n11322) );
  XNOR U19580 ( .A(n11314), .B(n11315), .Z(n11325) );
  XNOR U19581 ( .A(y[6999]), .B(x[6999]), .Z(n11315) );
  XNOR U19582 ( .A(n11316), .B(n11317), .Z(n11314) );
  XNOR U19583 ( .A(y[7000]), .B(x[7000]), .Z(n11317) );
  XNOR U19584 ( .A(y[7001]), .B(x[7001]), .Z(n11316) );
  NAND U19585 ( .A(n11381), .B(n11382), .Z(N64379) );
  NANDN U19586 ( .A(n11383), .B(n11384), .Z(n11382) );
  OR U19587 ( .A(n11385), .B(n11386), .Z(n11384) );
  NAND U19588 ( .A(n11385), .B(n11386), .Z(n11381) );
  XOR U19589 ( .A(n11385), .B(n11387), .Z(N64378) );
  XNOR U19590 ( .A(n11383), .B(n11386), .Z(n11387) );
  AND U19591 ( .A(n11388), .B(n11389), .Z(n11386) );
  NANDN U19592 ( .A(n11390), .B(n11391), .Z(n11389) );
  NANDN U19593 ( .A(n11392), .B(n11393), .Z(n11391) );
  NANDN U19594 ( .A(n11393), .B(n11392), .Z(n11388) );
  NAND U19595 ( .A(n11394), .B(n11395), .Z(n11383) );
  NANDN U19596 ( .A(n11396), .B(n11397), .Z(n11395) );
  OR U19597 ( .A(n11398), .B(n11399), .Z(n11397) );
  NAND U19598 ( .A(n11399), .B(n11398), .Z(n11394) );
  AND U19599 ( .A(n11400), .B(n11401), .Z(n11385) );
  NANDN U19600 ( .A(n11402), .B(n11403), .Z(n11401) );
  NANDN U19601 ( .A(n11404), .B(n11405), .Z(n11403) );
  NANDN U19602 ( .A(n11405), .B(n11404), .Z(n11400) );
  XOR U19603 ( .A(n11399), .B(n11406), .Z(N64377) );
  XOR U19604 ( .A(n11396), .B(n11398), .Z(n11406) );
  XNOR U19605 ( .A(n11392), .B(n11407), .Z(n11398) );
  XNOR U19606 ( .A(n11390), .B(n11393), .Z(n11407) );
  NAND U19607 ( .A(n11408), .B(n11409), .Z(n11393) );
  NAND U19608 ( .A(n11410), .B(n11411), .Z(n11409) );
  OR U19609 ( .A(n11412), .B(n11413), .Z(n11410) );
  NANDN U19610 ( .A(n11414), .B(n11412), .Z(n11408) );
  IV U19611 ( .A(n11413), .Z(n11414) );
  NAND U19612 ( .A(n11415), .B(n11416), .Z(n11390) );
  NAND U19613 ( .A(n11417), .B(n11418), .Z(n11416) );
  NANDN U19614 ( .A(n11419), .B(n11420), .Z(n11417) );
  NANDN U19615 ( .A(n11420), .B(n11419), .Z(n11415) );
  AND U19616 ( .A(n11421), .B(n11422), .Z(n11392) );
  NAND U19617 ( .A(n11423), .B(n11424), .Z(n11422) );
  OR U19618 ( .A(n11425), .B(n11426), .Z(n11423) );
  NANDN U19619 ( .A(n11427), .B(n11425), .Z(n11421) );
  NAND U19620 ( .A(n11428), .B(n11429), .Z(n11396) );
  NANDN U19621 ( .A(n11430), .B(n11431), .Z(n11429) );
  OR U19622 ( .A(n11432), .B(n11433), .Z(n11431) );
  NANDN U19623 ( .A(n11434), .B(n11432), .Z(n11428) );
  IV U19624 ( .A(n11433), .Z(n11434) );
  XNOR U19625 ( .A(n11404), .B(n11435), .Z(n11399) );
  XNOR U19626 ( .A(n11402), .B(n11405), .Z(n11435) );
  NAND U19627 ( .A(n11436), .B(n11437), .Z(n11405) );
  NAND U19628 ( .A(n11438), .B(n11439), .Z(n11437) );
  OR U19629 ( .A(n11440), .B(n11441), .Z(n11438) );
  NANDN U19630 ( .A(n11442), .B(n11440), .Z(n11436) );
  IV U19631 ( .A(n11441), .Z(n11442) );
  NAND U19632 ( .A(n11443), .B(n11444), .Z(n11402) );
  NAND U19633 ( .A(n11445), .B(n11446), .Z(n11444) );
  NANDN U19634 ( .A(n11447), .B(n11448), .Z(n11445) );
  NANDN U19635 ( .A(n11448), .B(n11447), .Z(n11443) );
  AND U19636 ( .A(n11449), .B(n11450), .Z(n11404) );
  NAND U19637 ( .A(n11451), .B(n11452), .Z(n11450) );
  OR U19638 ( .A(n11453), .B(n11454), .Z(n11451) );
  NANDN U19639 ( .A(n11455), .B(n11453), .Z(n11449) );
  XNOR U19640 ( .A(n11430), .B(n11456), .Z(N64376) );
  XOR U19641 ( .A(n11432), .B(n11433), .Z(n11456) );
  XNOR U19642 ( .A(n11446), .B(n11457), .Z(n11433) );
  XOR U19643 ( .A(n11447), .B(n11448), .Z(n11457) );
  XOR U19644 ( .A(n11453), .B(n11458), .Z(n11448) );
  XOR U19645 ( .A(n11452), .B(n11455), .Z(n11458) );
  IV U19646 ( .A(n11454), .Z(n11455) );
  NAND U19647 ( .A(n11459), .B(n11460), .Z(n11454) );
  OR U19648 ( .A(n11461), .B(n11462), .Z(n11460) );
  OR U19649 ( .A(n11463), .B(n11464), .Z(n11459) );
  NAND U19650 ( .A(n11465), .B(n11466), .Z(n11452) );
  OR U19651 ( .A(n11467), .B(n11468), .Z(n11466) );
  OR U19652 ( .A(n11469), .B(n11470), .Z(n11465) );
  NOR U19653 ( .A(n11471), .B(n11472), .Z(n11453) );
  ANDN U19654 ( .B(n11473), .A(n11474), .Z(n11447) );
  XNOR U19655 ( .A(n11440), .B(n11475), .Z(n11446) );
  XNOR U19656 ( .A(n11439), .B(n11441), .Z(n11475) );
  NAND U19657 ( .A(n11476), .B(n11477), .Z(n11441) );
  OR U19658 ( .A(n11478), .B(n11479), .Z(n11477) );
  OR U19659 ( .A(n11480), .B(n11481), .Z(n11476) );
  NAND U19660 ( .A(n11482), .B(n11483), .Z(n11439) );
  OR U19661 ( .A(n11484), .B(n11485), .Z(n11483) );
  OR U19662 ( .A(n11486), .B(n11487), .Z(n11482) );
  ANDN U19663 ( .B(n11488), .A(n11489), .Z(n11440) );
  IV U19664 ( .A(n11490), .Z(n11488) );
  ANDN U19665 ( .B(n11491), .A(n11492), .Z(n11432) );
  XOR U19666 ( .A(n11418), .B(n11493), .Z(n11430) );
  XOR U19667 ( .A(n11419), .B(n11420), .Z(n11493) );
  XOR U19668 ( .A(n11425), .B(n11494), .Z(n11420) );
  XOR U19669 ( .A(n11424), .B(n11427), .Z(n11494) );
  IV U19670 ( .A(n11426), .Z(n11427) );
  NAND U19671 ( .A(n11495), .B(n11496), .Z(n11426) );
  OR U19672 ( .A(n11497), .B(n11498), .Z(n11496) );
  OR U19673 ( .A(n11499), .B(n11500), .Z(n11495) );
  NAND U19674 ( .A(n11501), .B(n11502), .Z(n11424) );
  OR U19675 ( .A(n11503), .B(n11504), .Z(n11502) );
  OR U19676 ( .A(n11505), .B(n11506), .Z(n11501) );
  NOR U19677 ( .A(n11507), .B(n11508), .Z(n11425) );
  ANDN U19678 ( .B(n11509), .A(n11510), .Z(n11419) );
  IV U19679 ( .A(n11511), .Z(n11509) );
  XNOR U19680 ( .A(n11412), .B(n11512), .Z(n11418) );
  XNOR U19681 ( .A(n11411), .B(n11413), .Z(n11512) );
  NAND U19682 ( .A(n11513), .B(n11514), .Z(n11413) );
  OR U19683 ( .A(n11515), .B(n11516), .Z(n11514) );
  OR U19684 ( .A(n11517), .B(n11518), .Z(n11513) );
  NAND U19685 ( .A(n11519), .B(n11520), .Z(n11411) );
  OR U19686 ( .A(n11521), .B(n11522), .Z(n11520) );
  OR U19687 ( .A(n11523), .B(n11524), .Z(n11519) );
  ANDN U19688 ( .B(n11525), .A(n11526), .Z(n11412) );
  IV U19689 ( .A(n11527), .Z(n11525) );
  XNOR U19690 ( .A(n11492), .B(n11491), .Z(N64375) );
  XOR U19691 ( .A(n11511), .B(n11510), .Z(n11491) );
  XNOR U19692 ( .A(n11526), .B(n11527), .Z(n11510) );
  XNOR U19693 ( .A(n11521), .B(n11522), .Z(n11527) );
  XNOR U19694 ( .A(n11523), .B(n11524), .Z(n11522) );
  XNOR U19695 ( .A(y[6997]), .B(x[6997]), .Z(n11524) );
  XNOR U19696 ( .A(y[6998]), .B(x[6998]), .Z(n11523) );
  XNOR U19697 ( .A(y[6996]), .B(x[6996]), .Z(n11521) );
  XNOR U19698 ( .A(n11515), .B(n11516), .Z(n11526) );
  XNOR U19699 ( .A(y[6993]), .B(x[6993]), .Z(n11516) );
  XNOR U19700 ( .A(n11517), .B(n11518), .Z(n11515) );
  XNOR U19701 ( .A(y[6994]), .B(x[6994]), .Z(n11518) );
  XNOR U19702 ( .A(y[6995]), .B(x[6995]), .Z(n11517) );
  XNOR U19703 ( .A(n11508), .B(n11507), .Z(n11511) );
  XNOR U19704 ( .A(n11503), .B(n11504), .Z(n11507) );
  XNOR U19705 ( .A(y[6990]), .B(x[6990]), .Z(n11504) );
  XNOR U19706 ( .A(n11505), .B(n11506), .Z(n11503) );
  XNOR U19707 ( .A(y[6991]), .B(x[6991]), .Z(n11506) );
  XNOR U19708 ( .A(y[6992]), .B(x[6992]), .Z(n11505) );
  XNOR U19709 ( .A(n11497), .B(n11498), .Z(n11508) );
  XNOR U19710 ( .A(y[6987]), .B(x[6987]), .Z(n11498) );
  XNOR U19711 ( .A(n11499), .B(n11500), .Z(n11497) );
  XNOR U19712 ( .A(y[6988]), .B(x[6988]), .Z(n11500) );
  XNOR U19713 ( .A(y[6989]), .B(x[6989]), .Z(n11499) );
  XOR U19714 ( .A(n11473), .B(n11474), .Z(n11492) );
  XNOR U19715 ( .A(n11489), .B(n11490), .Z(n11474) );
  XNOR U19716 ( .A(n11484), .B(n11485), .Z(n11490) );
  XNOR U19717 ( .A(n11486), .B(n11487), .Z(n11485) );
  XNOR U19718 ( .A(y[6985]), .B(x[6985]), .Z(n11487) );
  XNOR U19719 ( .A(y[6986]), .B(x[6986]), .Z(n11486) );
  XNOR U19720 ( .A(y[6984]), .B(x[6984]), .Z(n11484) );
  XNOR U19721 ( .A(n11478), .B(n11479), .Z(n11489) );
  XNOR U19722 ( .A(y[6981]), .B(x[6981]), .Z(n11479) );
  XNOR U19723 ( .A(n11480), .B(n11481), .Z(n11478) );
  XNOR U19724 ( .A(y[6982]), .B(x[6982]), .Z(n11481) );
  XNOR U19725 ( .A(y[6983]), .B(x[6983]), .Z(n11480) );
  XOR U19726 ( .A(n11472), .B(n11471), .Z(n11473) );
  XNOR U19727 ( .A(n11467), .B(n11468), .Z(n11471) );
  XNOR U19728 ( .A(y[6978]), .B(x[6978]), .Z(n11468) );
  XNOR U19729 ( .A(n11469), .B(n11470), .Z(n11467) );
  XNOR U19730 ( .A(y[6979]), .B(x[6979]), .Z(n11470) );
  XNOR U19731 ( .A(y[6980]), .B(x[6980]), .Z(n11469) );
  XNOR U19732 ( .A(n11461), .B(n11462), .Z(n11472) );
  XNOR U19733 ( .A(y[6975]), .B(x[6975]), .Z(n11462) );
  XNOR U19734 ( .A(n11463), .B(n11464), .Z(n11461) );
  XNOR U19735 ( .A(y[6976]), .B(x[6976]), .Z(n11464) );
  XNOR U19736 ( .A(y[6977]), .B(x[6977]), .Z(n11463) );
  NAND U19737 ( .A(n11528), .B(n11529), .Z(N64366) );
  NANDN U19738 ( .A(n11530), .B(n11531), .Z(n11529) );
  OR U19739 ( .A(n11532), .B(n11533), .Z(n11531) );
  NAND U19740 ( .A(n11532), .B(n11533), .Z(n11528) );
  XOR U19741 ( .A(n11532), .B(n11534), .Z(N64365) );
  XNOR U19742 ( .A(n11530), .B(n11533), .Z(n11534) );
  AND U19743 ( .A(n11535), .B(n11536), .Z(n11533) );
  NANDN U19744 ( .A(n11537), .B(n11538), .Z(n11536) );
  NANDN U19745 ( .A(n11539), .B(n11540), .Z(n11538) );
  NANDN U19746 ( .A(n11540), .B(n11539), .Z(n11535) );
  NAND U19747 ( .A(n11541), .B(n11542), .Z(n11530) );
  NANDN U19748 ( .A(n11543), .B(n11544), .Z(n11542) );
  OR U19749 ( .A(n11545), .B(n11546), .Z(n11544) );
  NAND U19750 ( .A(n11546), .B(n11545), .Z(n11541) );
  AND U19751 ( .A(n11547), .B(n11548), .Z(n11532) );
  NANDN U19752 ( .A(n11549), .B(n11550), .Z(n11548) );
  NANDN U19753 ( .A(n11551), .B(n11552), .Z(n11550) );
  NANDN U19754 ( .A(n11552), .B(n11551), .Z(n11547) );
  XOR U19755 ( .A(n11546), .B(n11553), .Z(N64364) );
  XOR U19756 ( .A(n11543), .B(n11545), .Z(n11553) );
  XNOR U19757 ( .A(n11539), .B(n11554), .Z(n11545) );
  XNOR U19758 ( .A(n11537), .B(n11540), .Z(n11554) );
  NAND U19759 ( .A(n11555), .B(n11556), .Z(n11540) );
  NAND U19760 ( .A(n11557), .B(n11558), .Z(n11556) );
  OR U19761 ( .A(n11559), .B(n11560), .Z(n11557) );
  NANDN U19762 ( .A(n11561), .B(n11559), .Z(n11555) );
  IV U19763 ( .A(n11560), .Z(n11561) );
  NAND U19764 ( .A(n11562), .B(n11563), .Z(n11537) );
  NAND U19765 ( .A(n11564), .B(n11565), .Z(n11563) );
  NANDN U19766 ( .A(n11566), .B(n11567), .Z(n11564) );
  NANDN U19767 ( .A(n11567), .B(n11566), .Z(n11562) );
  AND U19768 ( .A(n11568), .B(n11569), .Z(n11539) );
  NAND U19769 ( .A(n11570), .B(n11571), .Z(n11569) );
  OR U19770 ( .A(n11572), .B(n11573), .Z(n11570) );
  NANDN U19771 ( .A(n11574), .B(n11572), .Z(n11568) );
  NAND U19772 ( .A(n11575), .B(n11576), .Z(n11543) );
  NANDN U19773 ( .A(n11577), .B(n11578), .Z(n11576) );
  OR U19774 ( .A(n11579), .B(n11580), .Z(n11578) );
  NANDN U19775 ( .A(n11581), .B(n11579), .Z(n11575) );
  IV U19776 ( .A(n11580), .Z(n11581) );
  XNOR U19777 ( .A(n11551), .B(n11582), .Z(n11546) );
  XNOR U19778 ( .A(n11549), .B(n11552), .Z(n11582) );
  NAND U19779 ( .A(n11583), .B(n11584), .Z(n11552) );
  NAND U19780 ( .A(n11585), .B(n11586), .Z(n11584) );
  OR U19781 ( .A(n11587), .B(n11588), .Z(n11585) );
  NANDN U19782 ( .A(n11589), .B(n11587), .Z(n11583) );
  IV U19783 ( .A(n11588), .Z(n11589) );
  NAND U19784 ( .A(n11590), .B(n11591), .Z(n11549) );
  NAND U19785 ( .A(n11592), .B(n11593), .Z(n11591) );
  NANDN U19786 ( .A(n11594), .B(n11595), .Z(n11592) );
  NANDN U19787 ( .A(n11595), .B(n11594), .Z(n11590) );
  AND U19788 ( .A(n11596), .B(n11597), .Z(n11551) );
  NAND U19789 ( .A(n11598), .B(n11599), .Z(n11597) );
  OR U19790 ( .A(n11600), .B(n11601), .Z(n11598) );
  NANDN U19791 ( .A(n11602), .B(n11600), .Z(n11596) );
  XNOR U19792 ( .A(n11577), .B(n11603), .Z(N64363) );
  XOR U19793 ( .A(n11579), .B(n11580), .Z(n11603) );
  XNOR U19794 ( .A(n11593), .B(n11604), .Z(n11580) );
  XOR U19795 ( .A(n11594), .B(n11595), .Z(n11604) );
  XOR U19796 ( .A(n11600), .B(n11605), .Z(n11595) );
  XOR U19797 ( .A(n11599), .B(n11602), .Z(n11605) );
  IV U19798 ( .A(n11601), .Z(n11602) );
  NAND U19799 ( .A(n11606), .B(n11607), .Z(n11601) );
  OR U19800 ( .A(n11608), .B(n11609), .Z(n11607) );
  OR U19801 ( .A(n11610), .B(n11611), .Z(n11606) );
  NAND U19802 ( .A(n11612), .B(n11613), .Z(n11599) );
  OR U19803 ( .A(n11614), .B(n11615), .Z(n11613) );
  OR U19804 ( .A(n11616), .B(n11617), .Z(n11612) );
  NOR U19805 ( .A(n11618), .B(n11619), .Z(n11600) );
  ANDN U19806 ( .B(n11620), .A(n11621), .Z(n11594) );
  XNOR U19807 ( .A(n11587), .B(n11622), .Z(n11593) );
  XNOR U19808 ( .A(n11586), .B(n11588), .Z(n11622) );
  NAND U19809 ( .A(n11623), .B(n11624), .Z(n11588) );
  OR U19810 ( .A(n11625), .B(n11626), .Z(n11624) );
  OR U19811 ( .A(n11627), .B(n11628), .Z(n11623) );
  NAND U19812 ( .A(n11629), .B(n11630), .Z(n11586) );
  OR U19813 ( .A(n11631), .B(n11632), .Z(n11630) );
  OR U19814 ( .A(n11633), .B(n11634), .Z(n11629) );
  ANDN U19815 ( .B(n11635), .A(n11636), .Z(n11587) );
  IV U19816 ( .A(n11637), .Z(n11635) );
  ANDN U19817 ( .B(n11638), .A(n11639), .Z(n11579) );
  XOR U19818 ( .A(n11565), .B(n11640), .Z(n11577) );
  XOR U19819 ( .A(n11566), .B(n11567), .Z(n11640) );
  XOR U19820 ( .A(n11572), .B(n11641), .Z(n11567) );
  XOR U19821 ( .A(n11571), .B(n11574), .Z(n11641) );
  IV U19822 ( .A(n11573), .Z(n11574) );
  NAND U19823 ( .A(n11642), .B(n11643), .Z(n11573) );
  OR U19824 ( .A(n11644), .B(n11645), .Z(n11643) );
  OR U19825 ( .A(n11646), .B(n11647), .Z(n11642) );
  NAND U19826 ( .A(n11648), .B(n11649), .Z(n11571) );
  OR U19827 ( .A(n11650), .B(n11651), .Z(n11649) );
  OR U19828 ( .A(n11652), .B(n11653), .Z(n11648) );
  NOR U19829 ( .A(n11654), .B(n11655), .Z(n11572) );
  ANDN U19830 ( .B(n11656), .A(n11657), .Z(n11566) );
  IV U19831 ( .A(n11658), .Z(n11656) );
  XNOR U19832 ( .A(n11559), .B(n11659), .Z(n11565) );
  XNOR U19833 ( .A(n11558), .B(n11560), .Z(n11659) );
  NAND U19834 ( .A(n11660), .B(n11661), .Z(n11560) );
  OR U19835 ( .A(n11662), .B(n11663), .Z(n11661) );
  OR U19836 ( .A(n11664), .B(n11665), .Z(n11660) );
  NAND U19837 ( .A(n11666), .B(n11667), .Z(n11558) );
  OR U19838 ( .A(n11668), .B(n11669), .Z(n11667) );
  OR U19839 ( .A(n11670), .B(n11671), .Z(n11666) );
  ANDN U19840 ( .B(n11672), .A(n11673), .Z(n11559) );
  IV U19841 ( .A(n11674), .Z(n11672) );
  XNOR U19842 ( .A(n11639), .B(n11638), .Z(N64362) );
  XOR U19843 ( .A(n11658), .B(n11657), .Z(n11638) );
  XNOR U19844 ( .A(n11673), .B(n11674), .Z(n11657) );
  XNOR U19845 ( .A(n11668), .B(n11669), .Z(n11674) );
  XNOR U19846 ( .A(n11670), .B(n11671), .Z(n11669) );
  XNOR U19847 ( .A(y[6973]), .B(x[6973]), .Z(n11671) );
  XNOR U19848 ( .A(y[6974]), .B(x[6974]), .Z(n11670) );
  XNOR U19849 ( .A(y[6972]), .B(x[6972]), .Z(n11668) );
  XNOR U19850 ( .A(n11662), .B(n11663), .Z(n11673) );
  XNOR U19851 ( .A(y[6969]), .B(x[6969]), .Z(n11663) );
  XNOR U19852 ( .A(n11664), .B(n11665), .Z(n11662) );
  XNOR U19853 ( .A(y[6970]), .B(x[6970]), .Z(n11665) );
  XNOR U19854 ( .A(y[6971]), .B(x[6971]), .Z(n11664) );
  XNOR U19855 ( .A(n11655), .B(n11654), .Z(n11658) );
  XNOR U19856 ( .A(n11650), .B(n11651), .Z(n11654) );
  XNOR U19857 ( .A(y[6966]), .B(x[6966]), .Z(n11651) );
  XNOR U19858 ( .A(n11652), .B(n11653), .Z(n11650) );
  XNOR U19859 ( .A(y[6967]), .B(x[6967]), .Z(n11653) );
  XNOR U19860 ( .A(y[6968]), .B(x[6968]), .Z(n11652) );
  XNOR U19861 ( .A(n11644), .B(n11645), .Z(n11655) );
  XNOR U19862 ( .A(y[6963]), .B(x[6963]), .Z(n11645) );
  XNOR U19863 ( .A(n11646), .B(n11647), .Z(n11644) );
  XNOR U19864 ( .A(y[6964]), .B(x[6964]), .Z(n11647) );
  XNOR U19865 ( .A(y[6965]), .B(x[6965]), .Z(n11646) );
  XOR U19866 ( .A(n11620), .B(n11621), .Z(n11639) );
  XNOR U19867 ( .A(n11636), .B(n11637), .Z(n11621) );
  XNOR U19868 ( .A(n11631), .B(n11632), .Z(n11637) );
  XNOR U19869 ( .A(n11633), .B(n11634), .Z(n11632) );
  XNOR U19870 ( .A(y[6961]), .B(x[6961]), .Z(n11634) );
  XNOR U19871 ( .A(y[6962]), .B(x[6962]), .Z(n11633) );
  XNOR U19872 ( .A(y[6960]), .B(x[6960]), .Z(n11631) );
  XNOR U19873 ( .A(n11625), .B(n11626), .Z(n11636) );
  XNOR U19874 ( .A(y[6957]), .B(x[6957]), .Z(n11626) );
  XNOR U19875 ( .A(n11627), .B(n11628), .Z(n11625) );
  XNOR U19876 ( .A(y[6958]), .B(x[6958]), .Z(n11628) );
  XNOR U19877 ( .A(y[6959]), .B(x[6959]), .Z(n11627) );
  XOR U19878 ( .A(n11619), .B(n11618), .Z(n11620) );
  XNOR U19879 ( .A(n11614), .B(n11615), .Z(n11618) );
  XNOR U19880 ( .A(y[6954]), .B(x[6954]), .Z(n11615) );
  XNOR U19881 ( .A(n11616), .B(n11617), .Z(n11614) );
  XNOR U19882 ( .A(y[6955]), .B(x[6955]), .Z(n11617) );
  XNOR U19883 ( .A(y[6956]), .B(x[6956]), .Z(n11616) );
  XNOR U19884 ( .A(n11608), .B(n11609), .Z(n11619) );
  XNOR U19885 ( .A(y[6951]), .B(x[6951]), .Z(n11609) );
  XNOR U19886 ( .A(n11610), .B(n11611), .Z(n11608) );
  XNOR U19887 ( .A(y[6952]), .B(x[6952]), .Z(n11611) );
  XNOR U19888 ( .A(y[6953]), .B(x[6953]), .Z(n11610) );
  NAND U19889 ( .A(n11675), .B(n11676), .Z(N64353) );
  NANDN U19890 ( .A(n11677), .B(n11678), .Z(n11676) );
  OR U19891 ( .A(n11679), .B(n11680), .Z(n11678) );
  NAND U19892 ( .A(n11679), .B(n11680), .Z(n11675) );
  XOR U19893 ( .A(n11679), .B(n11681), .Z(N64352) );
  XNOR U19894 ( .A(n11677), .B(n11680), .Z(n11681) );
  AND U19895 ( .A(n11682), .B(n11683), .Z(n11680) );
  NANDN U19896 ( .A(n11684), .B(n11685), .Z(n11683) );
  NANDN U19897 ( .A(n11686), .B(n11687), .Z(n11685) );
  NANDN U19898 ( .A(n11687), .B(n11686), .Z(n11682) );
  NAND U19899 ( .A(n11688), .B(n11689), .Z(n11677) );
  NANDN U19900 ( .A(n11690), .B(n11691), .Z(n11689) );
  OR U19901 ( .A(n11692), .B(n11693), .Z(n11691) );
  NAND U19902 ( .A(n11693), .B(n11692), .Z(n11688) );
  AND U19903 ( .A(n11694), .B(n11695), .Z(n11679) );
  NANDN U19904 ( .A(n11696), .B(n11697), .Z(n11695) );
  NANDN U19905 ( .A(n11698), .B(n11699), .Z(n11697) );
  NANDN U19906 ( .A(n11699), .B(n11698), .Z(n11694) );
  XOR U19907 ( .A(n11693), .B(n11700), .Z(N64351) );
  XOR U19908 ( .A(n11690), .B(n11692), .Z(n11700) );
  XNOR U19909 ( .A(n11686), .B(n11701), .Z(n11692) );
  XNOR U19910 ( .A(n11684), .B(n11687), .Z(n11701) );
  NAND U19911 ( .A(n11702), .B(n11703), .Z(n11687) );
  NAND U19912 ( .A(n11704), .B(n11705), .Z(n11703) );
  OR U19913 ( .A(n11706), .B(n11707), .Z(n11704) );
  NANDN U19914 ( .A(n11708), .B(n11706), .Z(n11702) );
  IV U19915 ( .A(n11707), .Z(n11708) );
  NAND U19916 ( .A(n11709), .B(n11710), .Z(n11684) );
  NAND U19917 ( .A(n11711), .B(n11712), .Z(n11710) );
  NANDN U19918 ( .A(n11713), .B(n11714), .Z(n11711) );
  NANDN U19919 ( .A(n11714), .B(n11713), .Z(n11709) );
  AND U19920 ( .A(n11715), .B(n11716), .Z(n11686) );
  NAND U19921 ( .A(n11717), .B(n11718), .Z(n11716) );
  OR U19922 ( .A(n11719), .B(n11720), .Z(n11717) );
  NANDN U19923 ( .A(n11721), .B(n11719), .Z(n11715) );
  NAND U19924 ( .A(n11722), .B(n11723), .Z(n11690) );
  NANDN U19925 ( .A(n11724), .B(n11725), .Z(n11723) );
  OR U19926 ( .A(n11726), .B(n11727), .Z(n11725) );
  NANDN U19927 ( .A(n11728), .B(n11726), .Z(n11722) );
  IV U19928 ( .A(n11727), .Z(n11728) );
  XNOR U19929 ( .A(n11698), .B(n11729), .Z(n11693) );
  XNOR U19930 ( .A(n11696), .B(n11699), .Z(n11729) );
  NAND U19931 ( .A(n11730), .B(n11731), .Z(n11699) );
  NAND U19932 ( .A(n11732), .B(n11733), .Z(n11731) );
  OR U19933 ( .A(n11734), .B(n11735), .Z(n11732) );
  NANDN U19934 ( .A(n11736), .B(n11734), .Z(n11730) );
  IV U19935 ( .A(n11735), .Z(n11736) );
  NAND U19936 ( .A(n11737), .B(n11738), .Z(n11696) );
  NAND U19937 ( .A(n11739), .B(n11740), .Z(n11738) );
  NANDN U19938 ( .A(n11741), .B(n11742), .Z(n11739) );
  NANDN U19939 ( .A(n11742), .B(n11741), .Z(n11737) );
  AND U19940 ( .A(n11743), .B(n11744), .Z(n11698) );
  NAND U19941 ( .A(n11745), .B(n11746), .Z(n11744) );
  OR U19942 ( .A(n11747), .B(n11748), .Z(n11745) );
  NANDN U19943 ( .A(n11749), .B(n11747), .Z(n11743) );
  XNOR U19944 ( .A(n11724), .B(n11750), .Z(N64350) );
  XOR U19945 ( .A(n11726), .B(n11727), .Z(n11750) );
  XNOR U19946 ( .A(n11740), .B(n11751), .Z(n11727) );
  XOR U19947 ( .A(n11741), .B(n11742), .Z(n11751) );
  XOR U19948 ( .A(n11747), .B(n11752), .Z(n11742) );
  XOR U19949 ( .A(n11746), .B(n11749), .Z(n11752) );
  IV U19950 ( .A(n11748), .Z(n11749) );
  NAND U19951 ( .A(n11753), .B(n11754), .Z(n11748) );
  OR U19952 ( .A(n11755), .B(n11756), .Z(n11754) );
  OR U19953 ( .A(n11757), .B(n11758), .Z(n11753) );
  NAND U19954 ( .A(n11759), .B(n11760), .Z(n11746) );
  OR U19955 ( .A(n11761), .B(n11762), .Z(n11760) );
  OR U19956 ( .A(n11763), .B(n11764), .Z(n11759) );
  NOR U19957 ( .A(n11765), .B(n11766), .Z(n11747) );
  ANDN U19958 ( .B(n11767), .A(n11768), .Z(n11741) );
  XNOR U19959 ( .A(n11734), .B(n11769), .Z(n11740) );
  XNOR U19960 ( .A(n11733), .B(n11735), .Z(n11769) );
  NAND U19961 ( .A(n11770), .B(n11771), .Z(n11735) );
  OR U19962 ( .A(n11772), .B(n11773), .Z(n11771) );
  OR U19963 ( .A(n11774), .B(n11775), .Z(n11770) );
  NAND U19964 ( .A(n11776), .B(n11777), .Z(n11733) );
  OR U19965 ( .A(n11778), .B(n11779), .Z(n11777) );
  OR U19966 ( .A(n11780), .B(n11781), .Z(n11776) );
  ANDN U19967 ( .B(n11782), .A(n11783), .Z(n11734) );
  IV U19968 ( .A(n11784), .Z(n11782) );
  ANDN U19969 ( .B(n11785), .A(n11786), .Z(n11726) );
  XOR U19970 ( .A(n11712), .B(n11787), .Z(n11724) );
  XOR U19971 ( .A(n11713), .B(n11714), .Z(n11787) );
  XOR U19972 ( .A(n11719), .B(n11788), .Z(n11714) );
  XOR U19973 ( .A(n11718), .B(n11721), .Z(n11788) );
  IV U19974 ( .A(n11720), .Z(n11721) );
  NAND U19975 ( .A(n11789), .B(n11790), .Z(n11720) );
  OR U19976 ( .A(n11791), .B(n11792), .Z(n11790) );
  OR U19977 ( .A(n11793), .B(n11794), .Z(n11789) );
  NAND U19978 ( .A(n11795), .B(n11796), .Z(n11718) );
  OR U19979 ( .A(n11797), .B(n11798), .Z(n11796) );
  OR U19980 ( .A(n11799), .B(n11800), .Z(n11795) );
  NOR U19981 ( .A(n11801), .B(n11802), .Z(n11719) );
  ANDN U19982 ( .B(n11803), .A(n11804), .Z(n11713) );
  IV U19983 ( .A(n11805), .Z(n11803) );
  XNOR U19984 ( .A(n11706), .B(n11806), .Z(n11712) );
  XNOR U19985 ( .A(n11705), .B(n11707), .Z(n11806) );
  NAND U19986 ( .A(n11807), .B(n11808), .Z(n11707) );
  OR U19987 ( .A(n11809), .B(n11810), .Z(n11808) );
  OR U19988 ( .A(n11811), .B(n11812), .Z(n11807) );
  NAND U19989 ( .A(n11813), .B(n11814), .Z(n11705) );
  OR U19990 ( .A(n11815), .B(n11816), .Z(n11814) );
  OR U19991 ( .A(n11817), .B(n11818), .Z(n11813) );
  ANDN U19992 ( .B(n11819), .A(n11820), .Z(n11706) );
  IV U19993 ( .A(n11821), .Z(n11819) );
  XNOR U19994 ( .A(n11786), .B(n11785), .Z(N64349) );
  XOR U19995 ( .A(n11805), .B(n11804), .Z(n11785) );
  XNOR U19996 ( .A(n11820), .B(n11821), .Z(n11804) );
  XNOR U19997 ( .A(n11815), .B(n11816), .Z(n11821) );
  XNOR U19998 ( .A(n11817), .B(n11818), .Z(n11816) );
  XNOR U19999 ( .A(y[6949]), .B(x[6949]), .Z(n11818) );
  XNOR U20000 ( .A(y[6950]), .B(x[6950]), .Z(n11817) );
  XNOR U20001 ( .A(y[6948]), .B(x[6948]), .Z(n11815) );
  XNOR U20002 ( .A(n11809), .B(n11810), .Z(n11820) );
  XNOR U20003 ( .A(y[6945]), .B(x[6945]), .Z(n11810) );
  XNOR U20004 ( .A(n11811), .B(n11812), .Z(n11809) );
  XNOR U20005 ( .A(y[6946]), .B(x[6946]), .Z(n11812) );
  XNOR U20006 ( .A(y[6947]), .B(x[6947]), .Z(n11811) );
  XNOR U20007 ( .A(n11802), .B(n11801), .Z(n11805) );
  XNOR U20008 ( .A(n11797), .B(n11798), .Z(n11801) );
  XNOR U20009 ( .A(y[6942]), .B(x[6942]), .Z(n11798) );
  XNOR U20010 ( .A(n11799), .B(n11800), .Z(n11797) );
  XNOR U20011 ( .A(y[6943]), .B(x[6943]), .Z(n11800) );
  XNOR U20012 ( .A(y[6944]), .B(x[6944]), .Z(n11799) );
  XNOR U20013 ( .A(n11791), .B(n11792), .Z(n11802) );
  XNOR U20014 ( .A(y[6939]), .B(x[6939]), .Z(n11792) );
  XNOR U20015 ( .A(n11793), .B(n11794), .Z(n11791) );
  XNOR U20016 ( .A(y[6940]), .B(x[6940]), .Z(n11794) );
  XNOR U20017 ( .A(y[6941]), .B(x[6941]), .Z(n11793) );
  XOR U20018 ( .A(n11767), .B(n11768), .Z(n11786) );
  XNOR U20019 ( .A(n11783), .B(n11784), .Z(n11768) );
  XNOR U20020 ( .A(n11778), .B(n11779), .Z(n11784) );
  XNOR U20021 ( .A(n11780), .B(n11781), .Z(n11779) );
  XNOR U20022 ( .A(y[6937]), .B(x[6937]), .Z(n11781) );
  XNOR U20023 ( .A(y[6938]), .B(x[6938]), .Z(n11780) );
  XNOR U20024 ( .A(y[6936]), .B(x[6936]), .Z(n11778) );
  XNOR U20025 ( .A(n11772), .B(n11773), .Z(n11783) );
  XNOR U20026 ( .A(y[6933]), .B(x[6933]), .Z(n11773) );
  XNOR U20027 ( .A(n11774), .B(n11775), .Z(n11772) );
  XNOR U20028 ( .A(y[6934]), .B(x[6934]), .Z(n11775) );
  XNOR U20029 ( .A(y[6935]), .B(x[6935]), .Z(n11774) );
  XOR U20030 ( .A(n11766), .B(n11765), .Z(n11767) );
  XNOR U20031 ( .A(n11761), .B(n11762), .Z(n11765) );
  XNOR U20032 ( .A(y[6930]), .B(x[6930]), .Z(n11762) );
  XNOR U20033 ( .A(n11763), .B(n11764), .Z(n11761) );
  XNOR U20034 ( .A(y[6931]), .B(x[6931]), .Z(n11764) );
  XNOR U20035 ( .A(y[6932]), .B(x[6932]), .Z(n11763) );
  XNOR U20036 ( .A(n11755), .B(n11756), .Z(n11766) );
  XNOR U20037 ( .A(y[6927]), .B(x[6927]), .Z(n11756) );
  XNOR U20038 ( .A(n11757), .B(n11758), .Z(n11755) );
  XNOR U20039 ( .A(y[6928]), .B(x[6928]), .Z(n11758) );
  XNOR U20040 ( .A(y[6929]), .B(x[6929]), .Z(n11757) );
  NAND U20041 ( .A(n11822), .B(n11823), .Z(N64340) );
  NANDN U20042 ( .A(n11824), .B(n11825), .Z(n11823) );
  OR U20043 ( .A(n11826), .B(n11827), .Z(n11825) );
  NAND U20044 ( .A(n11826), .B(n11827), .Z(n11822) );
  XOR U20045 ( .A(n11826), .B(n11828), .Z(N64339) );
  XNOR U20046 ( .A(n11824), .B(n11827), .Z(n11828) );
  AND U20047 ( .A(n11829), .B(n11830), .Z(n11827) );
  NANDN U20048 ( .A(n11831), .B(n11832), .Z(n11830) );
  NANDN U20049 ( .A(n11833), .B(n11834), .Z(n11832) );
  NANDN U20050 ( .A(n11834), .B(n11833), .Z(n11829) );
  NAND U20051 ( .A(n11835), .B(n11836), .Z(n11824) );
  NANDN U20052 ( .A(n11837), .B(n11838), .Z(n11836) );
  OR U20053 ( .A(n11839), .B(n11840), .Z(n11838) );
  NAND U20054 ( .A(n11840), .B(n11839), .Z(n11835) );
  AND U20055 ( .A(n11841), .B(n11842), .Z(n11826) );
  NANDN U20056 ( .A(n11843), .B(n11844), .Z(n11842) );
  NANDN U20057 ( .A(n11845), .B(n11846), .Z(n11844) );
  NANDN U20058 ( .A(n11846), .B(n11845), .Z(n11841) );
  XOR U20059 ( .A(n11840), .B(n11847), .Z(N64338) );
  XOR U20060 ( .A(n11837), .B(n11839), .Z(n11847) );
  XNOR U20061 ( .A(n11833), .B(n11848), .Z(n11839) );
  XNOR U20062 ( .A(n11831), .B(n11834), .Z(n11848) );
  NAND U20063 ( .A(n11849), .B(n11850), .Z(n11834) );
  NAND U20064 ( .A(n11851), .B(n11852), .Z(n11850) );
  OR U20065 ( .A(n11853), .B(n11854), .Z(n11851) );
  NANDN U20066 ( .A(n11855), .B(n11853), .Z(n11849) );
  IV U20067 ( .A(n11854), .Z(n11855) );
  NAND U20068 ( .A(n11856), .B(n11857), .Z(n11831) );
  NAND U20069 ( .A(n11858), .B(n11859), .Z(n11857) );
  NANDN U20070 ( .A(n11860), .B(n11861), .Z(n11858) );
  NANDN U20071 ( .A(n11861), .B(n11860), .Z(n11856) );
  AND U20072 ( .A(n11862), .B(n11863), .Z(n11833) );
  NAND U20073 ( .A(n11864), .B(n11865), .Z(n11863) );
  OR U20074 ( .A(n11866), .B(n11867), .Z(n11864) );
  NANDN U20075 ( .A(n11868), .B(n11866), .Z(n11862) );
  NAND U20076 ( .A(n11869), .B(n11870), .Z(n11837) );
  NANDN U20077 ( .A(n11871), .B(n11872), .Z(n11870) );
  OR U20078 ( .A(n11873), .B(n11874), .Z(n11872) );
  NANDN U20079 ( .A(n11875), .B(n11873), .Z(n11869) );
  IV U20080 ( .A(n11874), .Z(n11875) );
  XNOR U20081 ( .A(n11845), .B(n11876), .Z(n11840) );
  XNOR U20082 ( .A(n11843), .B(n11846), .Z(n11876) );
  NAND U20083 ( .A(n11877), .B(n11878), .Z(n11846) );
  NAND U20084 ( .A(n11879), .B(n11880), .Z(n11878) );
  OR U20085 ( .A(n11881), .B(n11882), .Z(n11879) );
  NANDN U20086 ( .A(n11883), .B(n11881), .Z(n11877) );
  IV U20087 ( .A(n11882), .Z(n11883) );
  NAND U20088 ( .A(n11884), .B(n11885), .Z(n11843) );
  NAND U20089 ( .A(n11886), .B(n11887), .Z(n11885) );
  NANDN U20090 ( .A(n11888), .B(n11889), .Z(n11886) );
  NANDN U20091 ( .A(n11889), .B(n11888), .Z(n11884) );
  AND U20092 ( .A(n11890), .B(n11891), .Z(n11845) );
  NAND U20093 ( .A(n11892), .B(n11893), .Z(n11891) );
  OR U20094 ( .A(n11894), .B(n11895), .Z(n11892) );
  NANDN U20095 ( .A(n11896), .B(n11894), .Z(n11890) );
  XNOR U20096 ( .A(n11871), .B(n11897), .Z(N64337) );
  XOR U20097 ( .A(n11873), .B(n11874), .Z(n11897) );
  XNOR U20098 ( .A(n11887), .B(n11898), .Z(n11874) );
  XOR U20099 ( .A(n11888), .B(n11889), .Z(n11898) );
  XOR U20100 ( .A(n11894), .B(n11899), .Z(n11889) );
  XOR U20101 ( .A(n11893), .B(n11896), .Z(n11899) );
  IV U20102 ( .A(n11895), .Z(n11896) );
  NAND U20103 ( .A(n11900), .B(n11901), .Z(n11895) );
  OR U20104 ( .A(n11902), .B(n11903), .Z(n11901) );
  OR U20105 ( .A(n11904), .B(n11905), .Z(n11900) );
  NAND U20106 ( .A(n11906), .B(n11907), .Z(n11893) );
  OR U20107 ( .A(n11908), .B(n11909), .Z(n11907) );
  OR U20108 ( .A(n11910), .B(n11911), .Z(n11906) );
  NOR U20109 ( .A(n11912), .B(n11913), .Z(n11894) );
  ANDN U20110 ( .B(n11914), .A(n11915), .Z(n11888) );
  XNOR U20111 ( .A(n11881), .B(n11916), .Z(n11887) );
  XNOR U20112 ( .A(n11880), .B(n11882), .Z(n11916) );
  NAND U20113 ( .A(n11917), .B(n11918), .Z(n11882) );
  OR U20114 ( .A(n11919), .B(n11920), .Z(n11918) );
  OR U20115 ( .A(n11921), .B(n11922), .Z(n11917) );
  NAND U20116 ( .A(n11923), .B(n11924), .Z(n11880) );
  OR U20117 ( .A(n11925), .B(n11926), .Z(n11924) );
  OR U20118 ( .A(n11927), .B(n11928), .Z(n11923) );
  ANDN U20119 ( .B(n11929), .A(n11930), .Z(n11881) );
  IV U20120 ( .A(n11931), .Z(n11929) );
  ANDN U20121 ( .B(n11932), .A(n11933), .Z(n11873) );
  XOR U20122 ( .A(n11859), .B(n11934), .Z(n11871) );
  XOR U20123 ( .A(n11860), .B(n11861), .Z(n11934) );
  XOR U20124 ( .A(n11866), .B(n11935), .Z(n11861) );
  XOR U20125 ( .A(n11865), .B(n11868), .Z(n11935) );
  IV U20126 ( .A(n11867), .Z(n11868) );
  NAND U20127 ( .A(n11936), .B(n11937), .Z(n11867) );
  OR U20128 ( .A(n11938), .B(n11939), .Z(n11937) );
  OR U20129 ( .A(n11940), .B(n11941), .Z(n11936) );
  NAND U20130 ( .A(n11942), .B(n11943), .Z(n11865) );
  OR U20131 ( .A(n11944), .B(n11945), .Z(n11943) );
  OR U20132 ( .A(n11946), .B(n11947), .Z(n11942) );
  NOR U20133 ( .A(n11948), .B(n11949), .Z(n11866) );
  ANDN U20134 ( .B(n11950), .A(n11951), .Z(n11860) );
  IV U20135 ( .A(n11952), .Z(n11950) );
  XNOR U20136 ( .A(n11853), .B(n11953), .Z(n11859) );
  XNOR U20137 ( .A(n11852), .B(n11854), .Z(n11953) );
  NAND U20138 ( .A(n11954), .B(n11955), .Z(n11854) );
  OR U20139 ( .A(n11956), .B(n11957), .Z(n11955) );
  OR U20140 ( .A(n11958), .B(n11959), .Z(n11954) );
  NAND U20141 ( .A(n11960), .B(n11961), .Z(n11852) );
  OR U20142 ( .A(n11962), .B(n11963), .Z(n11961) );
  OR U20143 ( .A(n11964), .B(n11965), .Z(n11960) );
  ANDN U20144 ( .B(n11966), .A(n11967), .Z(n11853) );
  IV U20145 ( .A(n11968), .Z(n11966) );
  XNOR U20146 ( .A(n11933), .B(n11932), .Z(N64336) );
  XOR U20147 ( .A(n11952), .B(n11951), .Z(n11932) );
  XNOR U20148 ( .A(n11967), .B(n11968), .Z(n11951) );
  XNOR U20149 ( .A(n11962), .B(n11963), .Z(n11968) );
  XNOR U20150 ( .A(n11964), .B(n11965), .Z(n11963) );
  XNOR U20151 ( .A(y[6925]), .B(x[6925]), .Z(n11965) );
  XNOR U20152 ( .A(y[6926]), .B(x[6926]), .Z(n11964) );
  XNOR U20153 ( .A(y[6924]), .B(x[6924]), .Z(n11962) );
  XNOR U20154 ( .A(n11956), .B(n11957), .Z(n11967) );
  XNOR U20155 ( .A(y[6921]), .B(x[6921]), .Z(n11957) );
  XNOR U20156 ( .A(n11958), .B(n11959), .Z(n11956) );
  XNOR U20157 ( .A(y[6922]), .B(x[6922]), .Z(n11959) );
  XNOR U20158 ( .A(y[6923]), .B(x[6923]), .Z(n11958) );
  XNOR U20159 ( .A(n11949), .B(n11948), .Z(n11952) );
  XNOR U20160 ( .A(n11944), .B(n11945), .Z(n11948) );
  XNOR U20161 ( .A(y[6918]), .B(x[6918]), .Z(n11945) );
  XNOR U20162 ( .A(n11946), .B(n11947), .Z(n11944) );
  XNOR U20163 ( .A(y[6919]), .B(x[6919]), .Z(n11947) );
  XNOR U20164 ( .A(y[6920]), .B(x[6920]), .Z(n11946) );
  XNOR U20165 ( .A(n11938), .B(n11939), .Z(n11949) );
  XNOR U20166 ( .A(y[6915]), .B(x[6915]), .Z(n11939) );
  XNOR U20167 ( .A(n11940), .B(n11941), .Z(n11938) );
  XNOR U20168 ( .A(y[6916]), .B(x[6916]), .Z(n11941) );
  XNOR U20169 ( .A(y[6917]), .B(x[6917]), .Z(n11940) );
  XOR U20170 ( .A(n11914), .B(n11915), .Z(n11933) );
  XNOR U20171 ( .A(n11930), .B(n11931), .Z(n11915) );
  XNOR U20172 ( .A(n11925), .B(n11926), .Z(n11931) );
  XNOR U20173 ( .A(n11927), .B(n11928), .Z(n11926) );
  XNOR U20174 ( .A(y[6913]), .B(x[6913]), .Z(n11928) );
  XNOR U20175 ( .A(y[6914]), .B(x[6914]), .Z(n11927) );
  XNOR U20176 ( .A(y[6912]), .B(x[6912]), .Z(n11925) );
  XNOR U20177 ( .A(n11919), .B(n11920), .Z(n11930) );
  XNOR U20178 ( .A(y[6909]), .B(x[6909]), .Z(n11920) );
  XNOR U20179 ( .A(n11921), .B(n11922), .Z(n11919) );
  XNOR U20180 ( .A(y[6910]), .B(x[6910]), .Z(n11922) );
  XNOR U20181 ( .A(y[6911]), .B(x[6911]), .Z(n11921) );
  XOR U20182 ( .A(n11913), .B(n11912), .Z(n11914) );
  XNOR U20183 ( .A(n11908), .B(n11909), .Z(n11912) );
  XNOR U20184 ( .A(y[6906]), .B(x[6906]), .Z(n11909) );
  XNOR U20185 ( .A(n11910), .B(n11911), .Z(n11908) );
  XNOR U20186 ( .A(y[6907]), .B(x[6907]), .Z(n11911) );
  XNOR U20187 ( .A(y[6908]), .B(x[6908]), .Z(n11910) );
  XNOR U20188 ( .A(n11902), .B(n11903), .Z(n11913) );
  XNOR U20189 ( .A(y[6903]), .B(x[6903]), .Z(n11903) );
  XNOR U20190 ( .A(n11904), .B(n11905), .Z(n11902) );
  XNOR U20191 ( .A(y[6904]), .B(x[6904]), .Z(n11905) );
  XNOR U20192 ( .A(y[6905]), .B(x[6905]), .Z(n11904) );
  NAND U20193 ( .A(n11969), .B(n11970), .Z(N64327) );
  NANDN U20194 ( .A(n11971), .B(n11972), .Z(n11970) );
  OR U20195 ( .A(n11973), .B(n11974), .Z(n11972) );
  NAND U20196 ( .A(n11973), .B(n11974), .Z(n11969) );
  XOR U20197 ( .A(n11973), .B(n11975), .Z(N64326) );
  XNOR U20198 ( .A(n11971), .B(n11974), .Z(n11975) );
  AND U20199 ( .A(n11976), .B(n11977), .Z(n11974) );
  NANDN U20200 ( .A(n11978), .B(n11979), .Z(n11977) );
  NANDN U20201 ( .A(n11980), .B(n11981), .Z(n11979) );
  NANDN U20202 ( .A(n11981), .B(n11980), .Z(n11976) );
  NAND U20203 ( .A(n11982), .B(n11983), .Z(n11971) );
  NANDN U20204 ( .A(n11984), .B(n11985), .Z(n11983) );
  OR U20205 ( .A(n11986), .B(n11987), .Z(n11985) );
  NAND U20206 ( .A(n11987), .B(n11986), .Z(n11982) );
  AND U20207 ( .A(n11988), .B(n11989), .Z(n11973) );
  NANDN U20208 ( .A(n11990), .B(n11991), .Z(n11989) );
  NANDN U20209 ( .A(n11992), .B(n11993), .Z(n11991) );
  NANDN U20210 ( .A(n11993), .B(n11992), .Z(n11988) );
  XOR U20211 ( .A(n11987), .B(n11994), .Z(N64325) );
  XOR U20212 ( .A(n11984), .B(n11986), .Z(n11994) );
  XNOR U20213 ( .A(n11980), .B(n11995), .Z(n11986) );
  XNOR U20214 ( .A(n11978), .B(n11981), .Z(n11995) );
  NAND U20215 ( .A(n11996), .B(n11997), .Z(n11981) );
  NAND U20216 ( .A(n11998), .B(n11999), .Z(n11997) );
  OR U20217 ( .A(n12000), .B(n12001), .Z(n11998) );
  NANDN U20218 ( .A(n12002), .B(n12000), .Z(n11996) );
  IV U20219 ( .A(n12001), .Z(n12002) );
  NAND U20220 ( .A(n12003), .B(n12004), .Z(n11978) );
  NAND U20221 ( .A(n12005), .B(n12006), .Z(n12004) );
  NANDN U20222 ( .A(n12007), .B(n12008), .Z(n12005) );
  NANDN U20223 ( .A(n12008), .B(n12007), .Z(n12003) );
  AND U20224 ( .A(n12009), .B(n12010), .Z(n11980) );
  NAND U20225 ( .A(n12011), .B(n12012), .Z(n12010) );
  OR U20226 ( .A(n12013), .B(n12014), .Z(n12011) );
  NANDN U20227 ( .A(n12015), .B(n12013), .Z(n12009) );
  NAND U20228 ( .A(n12016), .B(n12017), .Z(n11984) );
  NANDN U20229 ( .A(n12018), .B(n12019), .Z(n12017) );
  OR U20230 ( .A(n12020), .B(n12021), .Z(n12019) );
  NANDN U20231 ( .A(n12022), .B(n12020), .Z(n12016) );
  IV U20232 ( .A(n12021), .Z(n12022) );
  XNOR U20233 ( .A(n11992), .B(n12023), .Z(n11987) );
  XNOR U20234 ( .A(n11990), .B(n11993), .Z(n12023) );
  NAND U20235 ( .A(n12024), .B(n12025), .Z(n11993) );
  NAND U20236 ( .A(n12026), .B(n12027), .Z(n12025) );
  OR U20237 ( .A(n12028), .B(n12029), .Z(n12026) );
  NANDN U20238 ( .A(n12030), .B(n12028), .Z(n12024) );
  IV U20239 ( .A(n12029), .Z(n12030) );
  NAND U20240 ( .A(n12031), .B(n12032), .Z(n11990) );
  NAND U20241 ( .A(n12033), .B(n12034), .Z(n12032) );
  NANDN U20242 ( .A(n12035), .B(n12036), .Z(n12033) );
  NANDN U20243 ( .A(n12036), .B(n12035), .Z(n12031) );
  AND U20244 ( .A(n12037), .B(n12038), .Z(n11992) );
  NAND U20245 ( .A(n12039), .B(n12040), .Z(n12038) );
  OR U20246 ( .A(n12041), .B(n12042), .Z(n12039) );
  NANDN U20247 ( .A(n12043), .B(n12041), .Z(n12037) );
  XNOR U20248 ( .A(n12018), .B(n12044), .Z(N64324) );
  XOR U20249 ( .A(n12020), .B(n12021), .Z(n12044) );
  XNOR U20250 ( .A(n12034), .B(n12045), .Z(n12021) );
  XOR U20251 ( .A(n12035), .B(n12036), .Z(n12045) );
  XOR U20252 ( .A(n12041), .B(n12046), .Z(n12036) );
  XOR U20253 ( .A(n12040), .B(n12043), .Z(n12046) );
  IV U20254 ( .A(n12042), .Z(n12043) );
  NAND U20255 ( .A(n12047), .B(n12048), .Z(n12042) );
  OR U20256 ( .A(n12049), .B(n12050), .Z(n12048) );
  OR U20257 ( .A(n12051), .B(n12052), .Z(n12047) );
  NAND U20258 ( .A(n12053), .B(n12054), .Z(n12040) );
  OR U20259 ( .A(n12055), .B(n12056), .Z(n12054) );
  OR U20260 ( .A(n12057), .B(n12058), .Z(n12053) );
  NOR U20261 ( .A(n12059), .B(n12060), .Z(n12041) );
  ANDN U20262 ( .B(n12061), .A(n12062), .Z(n12035) );
  XNOR U20263 ( .A(n12028), .B(n12063), .Z(n12034) );
  XNOR U20264 ( .A(n12027), .B(n12029), .Z(n12063) );
  NAND U20265 ( .A(n12064), .B(n12065), .Z(n12029) );
  OR U20266 ( .A(n12066), .B(n12067), .Z(n12065) );
  OR U20267 ( .A(n12068), .B(n12069), .Z(n12064) );
  NAND U20268 ( .A(n12070), .B(n12071), .Z(n12027) );
  OR U20269 ( .A(n12072), .B(n12073), .Z(n12071) );
  OR U20270 ( .A(n12074), .B(n12075), .Z(n12070) );
  ANDN U20271 ( .B(n12076), .A(n12077), .Z(n12028) );
  IV U20272 ( .A(n12078), .Z(n12076) );
  ANDN U20273 ( .B(n12079), .A(n12080), .Z(n12020) );
  XOR U20274 ( .A(n12006), .B(n12081), .Z(n12018) );
  XOR U20275 ( .A(n12007), .B(n12008), .Z(n12081) );
  XOR U20276 ( .A(n12013), .B(n12082), .Z(n12008) );
  XOR U20277 ( .A(n12012), .B(n12015), .Z(n12082) );
  IV U20278 ( .A(n12014), .Z(n12015) );
  NAND U20279 ( .A(n12083), .B(n12084), .Z(n12014) );
  OR U20280 ( .A(n12085), .B(n12086), .Z(n12084) );
  OR U20281 ( .A(n12087), .B(n12088), .Z(n12083) );
  NAND U20282 ( .A(n12089), .B(n12090), .Z(n12012) );
  OR U20283 ( .A(n12091), .B(n12092), .Z(n12090) );
  OR U20284 ( .A(n12093), .B(n12094), .Z(n12089) );
  NOR U20285 ( .A(n12095), .B(n12096), .Z(n12013) );
  ANDN U20286 ( .B(n12097), .A(n12098), .Z(n12007) );
  IV U20287 ( .A(n12099), .Z(n12097) );
  XNOR U20288 ( .A(n12000), .B(n12100), .Z(n12006) );
  XNOR U20289 ( .A(n11999), .B(n12001), .Z(n12100) );
  NAND U20290 ( .A(n12101), .B(n12102), .Z(n12001) );
  OR U20291 ( .A(n12103), .B(n12104), .Z(n12102) );
  OR U20292 ( .A(n12105), .B(n12106), .Z(n12101) );
  NAND U20293 ( .A(n12107), .B(n12108), .Z(n11999) );
  OR U20294 ( .A(n12109), .B(n12110), .Z(n12108) );
  OR U20295 ( .A(n12111), .B(n12112), .Z(n12107) );
  ANDN U20296 ( .B(n12113), .A(n12114), .Z(n12000) );
  IV U20297 ( .A(n12115), .Z(n12113) );
  XNOR U20298 ( .A(n12080), .B(n12079), .Z(N64323) );
  XOR U20299 ( .A(n12099), .B(n12098), .Z(n12079) );
  XNOR U20300 ( .A(n12114), .B(n12115), .Z(n12098) );
  XNOR U20301 ( .A(n12109), .B(n12110), .Z(n12115) );
  XNOR U20302 ( .A(n12111), .B(n12112), .Z(n12110) );
  XNOR U20303 ( .A(y[6901]), .B(x[6901]), .Z(n12112) );
  XNOR U20304 ( .A(y[6902]), .B(x[6902]), .Z(n12111) );
  XNOR U20305 ( .A(y[6900]), .B(x[6900]), .Z(n12109) );
  XNOR U20306 ( .A(n12103), .B(n12104), .Z(n12114) );
  XNOR U20307 ( .A(y[6897]), .B(x[6897]), .Z(n12104) );
  XNOR U20308 ( .A(n12105), .B(n12106), .Z(n12103) );
  XNOR U20309 ( .A(y[6898]), .B(x[6898]), .Z(n12106) );
  XNOR U20310 ( .A(y[6899]), .B(x[6899]), .Z(n12105) );
  XNOR U20311 ( .A(n12096), .B(n12095), .Z(n12099) );
  XNOR U20312 ( .A(n12091), .B(n12092), .Z(n12095) );
  XNOR U20313 ( .A(y[6894]), .B(x[6894]), .Z(n12092) );
  XNOR U20314 ( .A(n12093), .B(n12094), .Z(n12091) );
  XNOR U20315 ( .A(y[6895]), .B(x[6895]), .Z(n12094) );
  XNOR U20316 ( .A(y[6896]), .B(x[6896]), .Z(n12093) );
  XNOR U20317 ( .A(n12085), .B(n12086), .Z(n12096) );
  XNOR U20318 ( .A(y[6891]), .B(x[6891]), .Z(n12086) );
  XNOR U20319 ( .A(n12087), .B(n12088), .Z(n12085) );
  XNOR U20320 ( .A(y[6892]), .B(x[6892]), .Z(n12088) );
  XNOR U20321 ( .A(y[6893]), .B(x[6893]), .Z(n12087) );
  XOR U20322 ( .A(n12061), .B(n12062), .Z(n12080) );
  XNOR U20323 ( .A(n12077), .B(n12078), .Z(n12062) );
  XNOR U20324 ( .A(n12072), .B(n12073), .Z(n12078) );
  XNOR U20325 ( .A(n12074), .B(n12075), .Z(n12073) );
  XNOR U20326 ( .A(y[6889]), .B(x[6889]), .Z(n12075) );
  XNOR U20327 ( .A(y[6890]), .B(x[6890]), .Z(n12074) );
  XNOR U20328 ( .A(y[6888]), .B(x[6888]), .Z(n12072) );
  XNOR U20329 ( .A(n12066), .B(n12067), .Z(n12077) );
  XNOR U20330 ( .A(y[6885]), .B(x[6885]), .Z(n12067) );
  XNOR U20331 ( .A(n12068), .B(n12069), .Z(n12066) );
  XNOR U20332 ( .A(y[6886]), .B(x[6886]), .Z(n12069) );
  XNOR U20333 ( .A(y[6887]), .B(x[6887]), .Z(n12068) );
  XOR U20334 ( .A(n12060), .B(n12059), .Z(n12061) );
  XNOR U20335 ( .A(n12055), .B(n12056), .Z(n12059) );
  XNOR U20336 ( .A(y[6882]), .B(x[6882]), .Z(n12056) );
  XNOR U20337 ( .A(n12057), .B(n12058), .Z(n12055) );
  XNOR U20338 ( .A(y[6883]), .B(x[6883]), .Z(n12058) );
  XNOR U20339 ( .A(y[6884]), .B(x[6884]), .Z(n12057) );
  XNOR U20340 ( .A(n12049), .B(n12050), .Z(n12060) );
  XNOR U20341 ( .A(y[6879]), .B(x[6879]), .Z(n12050) );
  XNOR U20342 ( .A(n12051), .B(n12052), .Z(n12049) );
  XNOR U20343 ( .A(y[6880]), .B(x[6880]), .Z(n12052) );
  XNOR U20344 ( .A(y[6881]), .B(x[6881]), .Z(n12051) );
  NAND U20345 ( .A(n12116), .B(n12117), .Z(N64314) );
  NANDN U20346 ( .A(n12118), .B(n12119), .Z(n12117) );
  OR U20347 ( .A(n12120), .B(n12121), .Z(n12119) );
  NAND U20348 ( .A(n12120), .B(n12121), .Z(n12116) );
  XOR U20349 ( .A(n12120), .B(n12122), .Z(N64313) );
  XNOR U20350 ( .A(n12118), .B(n12121), .Z(n12122) );
  AND U20351 ( .A(n12123), .B(n12124), .Z(n12121) );
  NANDN U20352 ( .A(n12125), .B(n12126), .Z(n12124) );
  NANDN U20353 ( .A(n12127), .B(n12128), .Z(n12126) );
  NANDN U20354 ( .A(n12128), .B(n12127), .Z(n12123) );
  NAND U20355 ( .A(n12129), .B(n12130), .Z(n12118) );
  NANDN U20356 ( .A(n12131), .B(n12132), .Z(n12130) );
  OR U20357 ( .A(n12133), .B(n12134), .Z(n12132) );
  NAND U20358 ( .A(n12134), .B(n12133), .Z(n12129) );
  AND U20359 ( .A(n12135), .B(n12136), .Z(n12120) );
  NANDN U20360 ( .A(n12137), .B(n12138), .Z(n12136) );
  NANDN U20361 ( .A(n12139), .B(n12140), .Z(n12138) );
  NANDN U20362 ( .A(n12140), .B(n12139), .Z(n12135) );
  XOR U20363 ( .A(n12134), .B(n12141), .Z(N64312) );
  XOR U20364 ( .A(n12131), .B(n12133), .Z(n12141) );
  XNOR U20365 ( .A(n12127), .B(n12142), .Z(n12133) );
  XNOR U20366 ( .A(n12125), .B(n12128), .Z(n12142) );
  NAND U20367 ( .A(n12143), .B(n12144), .Z(n12128) );
  NAND U20368 ( .A(n12145), .B(n12146), .Z(n12144) );
  OR U20369 ( .A(n12147), .B(n12148), .Z(n12145) );
  NANDN U20370 ( .A(n12149), .B(n12147), .Z(n12143) );
  IV U20371 ( .A(n12148), .Z(n12149) );
  NAND U20372 ( .A(n12150), .B(n12151), .Z(n12125) );
  NAND U20373 ( .A(n12152), .B(n12153), .Z(n12151) );
  NANDN U20374 ( .A(n12154), .B(n12155), .Z(n12152) );
  NANDN U20375 ( .A(n12155), .B(n12154), .Z(n12150) );
  AND U20376 ( .A(n12156), .B(n12157), .Z(n12127) );
  NAND U20377 ( .A(n12158), .B(n12159), .Z(n12157) );
  OR U20378 ( .A(n12160), .B(n12161), .Z(n12158) );
  NANDN U20379 ( .A(n12162), .B(n12160), .Z(n12156) );
  NAND U20380 ( .A(n12163), .B(n12164), .Z(n12131) );
  NANDN U20381 ( .A(n12165), .B(n12166), .Z(n12164) );
  OR U20382 ( .A(n12167), .B(n12168), .Z(n12166) );
  NANDN U20383 ( .A(n12169), .B(n12167), .Z(n12163) );
  IV U20384 ( .A(n12168), .Z(n12169) );
  XNOR U20385 ( .A(n12139), .B(n12170), .Z(n12134) );
  XNOR U20386 ( .A(n12137), .B(n12140), .Z(n12170) );
  NAND U20387 ( .A(n12171), .B(n12172), .Z(n12140) );
  NAND U20388 ( .A(n12173), .B(n12174), .Z(n12172) );
  OR U20389 ( .A(n12175), .B(n12176), .Z(n12173) );
  NANDN U20390 ( .A(n12177), .B(n12175), .Z(n12171) );
  IV U20391 ( .A(n12176), .Z(n12177) );
  NAND U20392 ( .A(n12178), .B(n12179), .Z(n12137) );
  NAND U20393 ( .A(n12180), .B(n12181), .Z(n12179) );
  NANDN U20394 ( .A(n12182), .B(n12183), .Z(n12180) );
  NANDN U20395 ( .A(n12183), .B(n12182), .Z(n12178) );
  AND U20396 ( .A(n12184), .B(n12185), .Z(n12139) );
  NAND U20397 ( .A(n12186), .B(n12187), .Z(n12185) );
  OR U20398 ( .A(n12188), .B(n12189), .Z(n12186) );
  NANDN U20399 ( .A(n12190), .B(n12188), .Z(n12184) );
  XNOR U20400 ( .A(n12165), .B(n12191), .Z(N64311) );
  XOR U20401 ( .A(n12167), .B(n12168), .Z(n12191) );
  XNOR U20402 ( .A(n12181), .B(n12192), .Z(n12168) );
  XOR U20403 ( .A(n12182), .B(n12183), .Z(n12192) );
  XOR U20404 ( .A(n12188), .B(n12193), .Z(n12183) );
  XOR U20405 ( .A(n12187), .B(n12190), .Z(n12193) );
  IV U20406 ( .A(n12189), .Z(n12190) );
  NAND U20407 ( .A(n12194), .B(n12195), .Z(n12189) );
  OR U20408 ( .A(n12196), .B(n12197), .Z(n12195) );
  OR U20409 ( .A(n12198), .B(n12199), .Z(n12194) );
  NAND U20410 ( .A(n12200), .B(n12201), .Z(n12187) );
  OR U20411 ( .A(n12202), .B(n12203), .Z(n12201) );
  OR U20412 ( .A(n12204), .B(n12205), .Z(n12200) );
  NOR U20413 ( .A(n12206), .B(n12207), .Z(n12188) );
  ANDN U20414 ( .B(n12208), .A(n12209), .Z(n12182) );
  XNOR U20415 ( .A(n12175), .B(n12210), .Z(n12181) );
  XNOR U20416 ( .A(n12174), .B(n12176), .Z(n12210) );
  NAND U20417 ( .A(n12211), .B(n12212), .Z(n12176) );
  OR U20418 ( .A(n12213), .B(n12214), .Z(n12212) );
  OR U20419 ( .A(n12215), .B(n12216), .Z(n12211) );
  NAND U20420 ( .A(n12217), .B(n12218), .Z(n12174) );
  OR U20421 ( .A(n12219), .B(n12220), .Z(n12218) );
  OR U20422 ( .A(n12221), .B(n12222), .Z(n12217) );
  ANDN U20423 ( .B(n12223), .A(n12224), .Z(n12175) );
  IV U20424 ( .A(n12225), .Z(n12223) );
  ANDN U20425 ( .B(n12226), .A(n12227), .Z(n12167) );
  XOR U20426 ( .A(n12153), .B(n12228), .Z(n12165) );
  XOR U20427 ( .A(n12154), .B(n12155), .Z(n12228) );
  XOR U20428 ( .A(n12160), .B(n12229), .Z(n12155) );
  XOR U20429 ( .A(n12159), .B(n12162), .Z(n12229) );
  IV U20430 ( .A(n12161), .Z(n12162) );
  NAND U20431 ( .A(n12230), .B(n12231), .Z(n12161) );
  OR U20432 ( .A(n12232), .B(n12233), .Z(n12231) );
  OR U20433 ( .A(n12234), .B(n12235), .Z(n12230) );
  NAND U20434 ( .A(n12236), .B(n12237), .Z(n12159) );
  OR U20435 ( .A(n12238), .B(n12239), .Z(n12237) );
  OR U20436 ( .A(n12240), .B(n12241), .Z(n12236) );
  NOR U20437 ( .A(n12242), .B(n12243), .Z(n12160) );
  ANDN U20438 ( .B(n12244), .A(n12245), .Z(n12154) );
  IV U20439 ( .A(n12246), .Z(n12244) );
  XNOR U20440 ( .A(n12147), .B(n12247), .Z(n12153) );
  XNOR U20441 ( .A(n12146), .B(n12148), .Z(n12247) );
  NAND U20442 ( .A(n12248), .B(n12249), .Z(n12148) );
  OR U20443 ( .A(n12250), .B(n12251), .Z(n12249) );
  OR U20444 ( .A(n12252), .B(n12253), .Z(n12248) );
  NAND U20445 ( .A(n12254), .B(n12255), .Z(n12146) );
  OR U20446 ( .A(n12256), .B(n12257), .Z(n12255) );
  OR U20447 ( .A(n12258), .B(n12259), .Z(n12254) );
  ANDN U20448 ( .B(n12260), .A(n12261), .Z(n12147) );
  IV U20449 ( .A(n12262), .Z(n12260) );
  XNOR U20450 ( .A(n12227), .B(n12226), .Z(N64310) );
  XOR U20451 ( .A(n12246), .B(n12245), .Z(n12226) );
  XNOR U20452 ( .A(n12261), .B(n12262), .Z(n12245) );
  XNOR U20453 ( .A(n12256), .B(n12257), .Z(n12262) );
  XNOR U20454 ( .A(n12258), .B(n12259), .Z(n12257) );
  XNOR U20455 ( .A(y[6877]), .B(x[6877]), .Z(n12259) );
  XNOR U20456 ( .A(y[6878]), .B(x[6878]), .Z(n12258) );
  XNOR U20457 ( .A(y[6876]), .B(x[6876]), .Z(n12256) );
  XNOR U20458 ( .A(n12250), .B(n12251), .Z(n12261) );
  XNOR U20459 ( .A(y[6873]), .B(x[6873]), .Z(n12251) );
  XNOR U20460 ( .A(n12252), .B(n12253), .Z(n12250) );
  XNOR U20461 ( .A(y[6874]), .B(x[6874]), .Z(n12253) );
  XNOR U20462 ( .A(y[6875]), .B(x[6875]), .Z(n12252) );
  XNOR U20463 ( .A(n12243), .B(n12242), .Z(n12246) );
  XNOR U20464 ( .A(n12238), .B(n12239), .Z(n12242) );
  XNOR U20465 ( .A(y[6870]), .B(x[6870]), .Z(n12239) );
  XNOR U20466 ( .A(n12240), .B(n12241), .Z(n12238) );
  XNOR U20467 ( .A(y[6871]), .B(x[6871]), .Z(n12241) );
  XNOR U20468 ( .A(y[6872]), .B(x[6872]), .Z(n12240) );
  XNOR U20469 ( .A(n12232), .B(n12233), .Z(n12243) );
  XNOR U20470 ( .A(y[6867]), .B(x[6867]), .Z(n12233) );
  XNOR U20471 ( .A(n12234), .B(n12235), .Z(n12232) );
  XNOR U20472 ( .A(y[6868]), .B(x[6868]), .Z(n12235) );
  XNOR U20473 ( .A(y[6869]), .B(x[6869]), .Z(n12234) );
  XOR U20474 ( .A(n12208), .B(n12209), .Z(n12227) );
  XNOR U20475 ( .A(n12224), .B(n12225), .Z(n12209) );
  XNOR U20476 ( .A(n12219), .B(n12220), .Z(n12225) );
  XNOR U20477 ( .A(n12221), .B(n12222), .Z(n12220) );
  XNOR U20478 ( .A(y[6865]), .B(x[6865]), .Z(n12222) );
  XNOR U20479 ( .A(y[6866]), .B(x[6866]), .Z(n12221) );
  XNOR U20480 ( .A(y[6864]), .B(x[6864]), .Z(n12219) );
  XNOR U20481 ( .A(n12213), .B(n12214), .Z(n12224) );
  XNOR U20482 ( .A(y[6861]), .B(x[6861]), .Z(n12214) );
  XNOR U20483 ( .A(n12215), .B(n12216), .Z(n12213) );
  XNOR U20484 ( .A(y[6862]), .B(x[6862]), .Z(n12216) );
  XNOR U20485 ( .A(y[6863]), .B(x[6863]), .Z(n12215) );
  XOR U20486 ( .A(n12207), .B(n12206), .Z(n12208) );
  XNOR U20487 ( .A(n12202), .B(n12203), .Z(n12206) );
  XNOR U20488 ( .A(y[6858]), .B(x[6858]), .Z(n12203) );
  XNOR U20489 ( .A(n12204), .B(n12205), .Z(n12202) );
  XNOR U20490 ( .A(y[6859]), .B(x[6859]), .Z(n12205) );
  XNOR U20491 ( .A(y[6860]), .B(x[6860]), .Z(n12204) );
  XNOR U20492 ( .A(n12196), .B(n12197), .Z(n12207) );
  XNOR U20493 ( .A(y[6855]), .B(x[6855]), .Z(n12197) );
  XNOR U20494 ( .A(n12198), .B(n12199), .Z(n12196) );
  XNOR U20495 ( .A(y[6856]), .B(x[6856]), .Z(n12199) );
  XNOR U20496 ( .A(y[6857]), .B(x[6857]), .Z(n12198) );
  NAND U20497 ( .A(n12263), .B(n12264), .Z(N64301) );
  NANDN U20498 ( .A(n12265), .B(n12266), .Z(n12264) );
  OR U20499 ( .A(n12267), .B(n12268), .Z(n12266) );
  NAND U20500 ( .A(n12267), .B(n12268), .Z(n12263) );
  XOR U20501 ( .A(n12267), .B(n12269), .Z(N64300) );
  XNOR U20502 ( .A(n12265), .B(n12268), .Z(n12269) );
  AND U20503 ( .A(n12270), .B(n12271), .Z(n12268) );
  NANDN U20504 ( .A(n12272), .B(n12273), .Z(n12271) );
  NANDN U20505 ( .A(n12274), .B(n12275), .Z(n12273) );
  NANDN U20506 ( .A(n12275), .B(n12274), .Z(n12270) );
  NAND U20507 ( .A(n12276), .B(n12277), .Z(n12265) );
  NANDN U20508 ( .A(n12278), .B(n12279), .Z(n12277) );
  OR U20509 ( .A(n12280), .B(n12281), .Z(n12279) );
  NAND U20510 ( .A(n12281), .B(n12280), .Z(n12276) );
  AND U20511 ( .A(n12282), .B(n12283), .Z(n12267) );
  NANDN U20512 ( .A(n12284), .B(n12285), .Z(n12283) );
  NANDN U20513 ( .A(n12286), .B(n12287), .Z(n12285) );
  NANDN U20514 ( .A(n12287), .B(n12286), .Z(n12282) );
  XOR U20515 ( .A(n12281), .B(n12288), .Z(N64299) );
  XOR U20516 ( .A(n12278), .B(n12280), .Z(n12288) );
  XNOR U20517 ( .A(n12274), .B(n12289), .Z(n12280) );
  XNOR U20518 ( .A(n12272), .B(n12275), .Z(n12289) );
  NAND U20519 ( .A(n12290), .B(n12291), .Z(n12275) );
  NAND U20520 ( .A(n12292), .B(n12293), .Z(n12291) );
  OR U20521 ( .A(n12294), .B(n12295), .Z(n12292) );
  NANDN U20522 ( .A(n12296), .B(n12294), .Z(n12290) );
  IV U20523 ( .A(n12295), .Z(n12296) );
  NAND U20524 ( .A(n12297), .B(n12298), .Z(n12272) );
  NAND U20525 ( .A(n12299), .B(n12300), .Z(n12298) );
  NANDN U20526 ( .A(n12301), .B(n12302), .Z(n12299) );
  NANDN U20527 ( .A(n12302), .B(n12301), .Z(n12297) );
  AND U20528 ( .A(n12303), .B(n12304), .Z(n12274) );
  NAND U20529 ( .A(n12305), .B(n12306), .Z(n12304) );
  OR U20530 ( .A(n12307), .B(n12308), .Z(n12305) );
  NANDN U20531 ( .A(n12309), .B(n12307), .Z(n12303) );
  NAND U20532 ( .A(n12310), .B(n12311), .Z(n12278) );
  NANDN U20533 ( .A(n12312), .B(n12313), .Z(n12311) );
  OR U20534 ( .A(n12314), .B(n12315), .Z(n12313) );
  NANDN U20535 ( .A(n12316), .B(n12314), .Z(n12310) );
  IV U20536 ( .A(n12315), .Z(n12316) );
  XNOR U20537 ( .A(n12286), .B(n12317), .Z(n12281) );
  XNOR U20538 ( .A(n12284), .B(n12287), .Z(n12317) );
  NAND U20539 ( .A(n12318), .B(n12319), .Z(n12287) );
  NAND U20540 ( .A(n12320), .B(n12321), .Z(n12319) );
  OR U20541 ( .A(n12322), .B(n12323), .Z(n12320) );
  NANDN U20542 ( .A(n12324), .B(n12322), .Z(n12318) );
  IV U20543 ( .A(n12323), .Z(n12324) );
  NAND U20544 ( .A(n12325), .B(n12326), .Z(n12284) );
  NAND U20545 ( .A(n12327), .B(n12328), .Z(n12326) );
  NANDN U20546 ( .A(n12329), .B(n12330), .Z(n12327) );
  NANDN U20547 ( .A(n12330), .B(n12329), .Z(n12325) );
  AND U20548 ( .A(n12331), .B(n12332), .Z(n12286) );
  NAND U20549 ( .A(n12333), .B(n12334), .Z(n12332) );
  OR U20550 ( .A(n12335), .B(n12336), .Z(n12333) );
  NANDN U20551 ( .A(n12337), .B(n12335), .Z(n12331) );
  XNOR U20552 ( .A(n12312), .B(n12338), .Z(N64298) );
  XOR U20553 ( .A(n12314), .B(n12315), .Z(n12338) );
  XNOR U20554 ( .A(n12328), .B(n12339), .Z(n12315) );
  XOR U20555 ( .A(n12329), .B(n12330), .Z(n12339) );
  XOR U20556 ( .A(n12335), .B(n12340), .Z(n12330) );
  XOR U20557 ( .A(n12334), .B(n12337), .Z(n12340) );
  IV U20558 ( .A(n12336), .Z(n12337) );
  NAND U20559 ( .A(n12341), .B(n12342), .Z(n12336) );
  OR U20560 ( .A(n12343), .B(n12344), .Z(n12342) );
  OR U20561 ( .A(n12345), .B(n12346), .Z(n12341) );
  NAND U20562 ( .A(n12347), .B(n12348), .Z(n12334) );
  OR U20563 ( .A(n12349), .B(n12350), .Z(n12348) );
  OR U20564 ( .A(n12351), .B(n12352), .Z(n12347) );
  NOR U20565 ( .A(n12353), .B(n12354), .Z(n12335) );
  ANDN U20566 ( .B(n12355), .A(n12356), .Z(n12329) );
  XNOR U20567 ( .A(n12322), .B(n12357), .Z(n12328) );
  XNOR U20568 ( .A(n12321), .B(n12323), .Z(n12357) );
  NAND U20569 ( .A(n12358), .B(n12359), .Z(n12323) );
  OR U20570 ( .A(n12360), .B(n12361), .Z(n12359) );
  OR U20571 ( .A(n12362), .B(n12363), .Z(n12358) );
  NAND U20572 ( .A(n12364), .B(n12365), .Z(n12321) );
  OR U20573 ( .A(n12366), .B(n12367), .Z(n12365) );
  OR U20574 ( .A(n12368), .B(n12369), .Z(n12364) );
  ANDN U20575 ( .B(n12370), .A(n12371), .Z(n12322) );
  IV U20576 ( .A(n12372), .Z(n12370) );
  ANDN U20577 ( .B(n12373), .A(n12374), .Z(n12314) );
  XOR U20578 ( .A(n12300), .B(n12375), .Z(n12312) );
  XOR U20579 ( .A(n12301), .B(n12302), .Z(n12375) );
  XOR U20580 ( .A(n12307), .B(n12376), .Z(n12302) );
  XOR U20581 ( .A(n12306), .B(n12309), .Z(n12376) );
  IV U20582 ( .A(n12308), .Z(n12309) );
  NAND U20583 ( .A(n12377), .B(n12378), .Z(n12308) );
  OR U20584 ( .A(n12379), .B(n12380), .Z(n12378) );
  OR U20585 ( .A(n12381), .B(n12382), .Z(n12377) );
  NAND U20586 ( .A(n12383), .B(n12384), .Z(n12306) );
  OR U20587 ( .A(n12385), .B(n12386), .Z(n12384) );
  OR U20588 ( .A(n12387), .B(n12388), .Z(n12383) );
  NOR U20589 ( .A(n12389), .B(n12390), .Z(n12307) );
  ANDN U20590 ( .B(n12391), .A(n12392), .Z(n12301) );
  IV U20591 ( .A(n12393), .Z(n12391) );
  XNOR U20592 ( .A(n12294), .B(n12394), .Z(n12300) );
  XNOR U20593 ( .A(n12293), .B(n12295), .Z(n12394) );
  NAND U20594 ( .A(n12395), .B(n12396), .Z(n12295) );
  OR U20595 ( .A(n12397), .B(n12398), .Z(n12396) );
  OR U20596 ( .A(n12399), .B(n12400), .Z(n12395) );
  NAND U20597 ( .A(n12401), .B(n12402), .Z(n12293) );
  OR U20598 ( .A(n12403), .B(n12404), .Z(n12402) );
  OR U20599 ( .A(n12405), .B(n12406), .Z(n12401) );
  ANDN U20600 ( .B(n12407), .A(n12408), .Z(n12294) );
  IV U20601 ( .A(n12409), .Z(n12407) );
  XNOR U20602 ( .A(n12374), .B(n12373), .Z(N64297) );
  XOR U20603 ( .A(n12393), .B(n12392), .Z(n12373) );
  XNOR U20604 ( .A(n12408), .B(n12409), .Z(n12392) );
  XNOR U20605 ( .A(n12403), .B(n12404), .Z(n12409) );
  XNOR U20606 ( .A(n12405), .B(n12406), .Z(n12404) );
  XNOR U20607 ( .A(y[6853]), .B(x[6853]), .Z(n12406) );
  XNOR U20608 ( .A(y[6854]), .B(x[6854]), .Z(n12405) );
  XNOR U20609 ( .A(y[6852]), .B(x[6852]), .Z(n12403) );
  XNOR U20610 ( .A(n12397), .B(n12398), .Z(n12408) );
  XNOR U20611 ( .A(y[6849]), .B(x[6849]), .Z(n12398) );
  XNOR U20612 ( .A(n12399), .B(n12400), .Z(n12397) );
  XNOR U20613 ( .A(y[6850]), .B(x[6850]), .Z(n12400) );
  XNOR U20614 ( .A(y[6851]), .B(x[6851]), .Z(n12399) );
  XNOR U20615 ( .A(n12390), .B(n12389), .Z(n12393) );
  XNOR U20616 ( .A(n12385), .B(n12386), .Z(n12389) );
  XNOR U20617 ( .A(y[6846]), .B(x[6846]), .Z(n12386) );
  XNOR U20618 ( .A(n12387), .B(n12388), .Z(n12385) );
  XNOR U20619 ( .A(y[6847]), .B(x[6847]), .Z(n12388) );
  XNOR U20620 ( .A(y[6848]), .B(x[6848]), .Z(n12387) );
  XNOR U20621 ( .A(n12379), .B(n12380), .Z(n12390) );
  XNOR U20622 ( .A(y[6843]), .B(x[6843]), .Z(n12380) );
  XNOR U20623 ( .A(n12381), .B(n12382), .Z(n12379) );
  XNOR U20624 ( .A(y[6844]), .B(x[6844]), .Z(n12382) );
  XNOR U20625 ( .A(y[6845]), .B(x[6845]), .Z(n12381) );
  XOR U20626 ( .A(n12355), .B(n12356), .Z(n12374) );
  XNOR U20627 ( .A(n12371), .B(n12372), .Z(n12356) );
  XNOR U20628 ( .A(n12366), .B(n12367), .Z(n12372) );
  XNOR U20629 ( .A(n12368), .B(n12369), .Z(n12367) );
  XNOR U20630 ( .A(y[6841]), .B(x[6841]), .Z(n12369) );
  XNOR U20631 ( .A(y[6842]), .B(x[6842]), .Z(n12368) );
  XNOR U20632 ( .A(y[6840]), .B(x[6840]), .Z(n12366) );
  XNOR U20633 ( .A(n12360), .B(n12361), .Z(n12371) );
  XNOR U20634 ( .A(y[6837]), .B(x[6837]), .Z(n12361) );
  XNOR U20635 ( .A(n12362), .B(n12363), .Z(n12360) );
  XNOR U20636 ( .A(y[6838]), .B(x[6838]), .Z(n12363) );
  XNOR U20637 ( .A(y[6839]), .B(x[6839]), .Z(n12362) );
  XOR U20638 ( .A(n12354), .B(n12353), .Z(n12355) );
  XNOR U20639 ( .A(n12349), .B(n12350), .Z(n12353) );
  XNOR U20640 ( .A(y[6834]), .B(x[6834]), .Z(n12350) );
  XNOR U20641 ( .A(n12351), .B(n12352), .Z(n12349) );
  XNOR U20642 ( .A(y[6835]), .B(x[6835]), .Z(n12352) );
  XNOR U20643 ( .A(y[6836]), .B(x[6836]), .Z(n12351) );
  XNOR U20644 ( .A(n12343), .B(n12344), .Z(n12354) );
  XNOR U20645 ( .A(y[6831]), .B(x[6831]), .Z(n12344) );
  XNOR U20646 ( .A(n12345), .B(n12346), .Z(n12343) );
  XNOR U20647 ( .A(y[6832]), .B(x[6832]), .Z(n12346) );
  XNOR U20648 ( .A(y[6833]), .B(x[6833]), .Z(n12345) );
  NAND U20649 ( .A(n12410), .B(n12411), .Z(N64288) );
  NANDN U20650 ( .A(n12412), .B(n12413), .Z(n12411) );
  OR U20651 ( .A(n12414), .B(n12415), .Z(n12413) );
  NAND U20652 ( .A(n12414), .B(n12415), .Z(n12410) );
  XOR U20653 ( .A(n12414), .B(n12416), .Z(N64287) );
  XNOR U20654 ( .A(n12412), .B(n12415), .Z(n12416) );
  AND U20655 ( .A(n12417), .B(n12418), .Z(n12415) );
  NANDN U20656 ( .A(n12419), .B(n12420), .Z(n12418) );
  NANDN U20657 ( .A(n12421), .B(n12422), .Z(n12420) );
  NANDN U20658 ( .A(n12422), .B(n12421), .Z(n12417) );
  NAND U20659 ( .A(n12423), .B(n12424), .Z(n12412) );
  NANDN U20660 ( .A(n12425), .B(n12426), .Z(n12424) );
  OR U20661 ( .A(n12427), .B(n12428), .Z(n12426) );
  NAND U20662 ( .A(n12428), .B(n12427), .Z(n12423) );
  AND U20663 ( .A(n12429), .B(n12430), .Z(n12414) );
  NANDN U20664 ( .A(n12431), .B(n12432), .Z(n12430) );
  NANDN U20665 ( .A(n12433), .B(n12434), .Z(n12432) );
  NANDN U20666 ( .A(n12434), .B(n12433), .Z(n12429) );
  XOR U20667 ( .A(n12428), .B(n12435), .Z(N64286) );
  XOR U20668 ( .A(n12425), .B(n12427), .Z(n12435) );
  XNOR U20669 ( .A(n12421), .B(n12436), .Z(n12427) );
  XNOR U20670 ( .A(n12419), .B(n12422), .Z(n12436) );
  NAND U20671 ( .A(n12437), .B(n12438), .Z(n12422) );
  NAND U20672 ( .A(n12439), .B(n12440), .Z(n12438) );
  OR U20673 ( .A(n12441), .B(n12442), .Z(n12439) );
  NANDN U20674 ( .A(n12443), .B(n12441), .Z(n12437) );
  IV U20675 ( .A(n12442), .Z(n12443) );
  NAND U20676 ( .A(n12444), .B(n12445), .Z(n12419) );
  NAND U20677 ( .A(n12446), .B(n12447), .Z(n12445) );
  NANDN U20678 ( .A(n12448), .B(n12449), .Z(n12446) );
  NANDN U20679 ( .A(n12449), .B(n12448), .Z(n12444) );
  AND U20680 ( .A(n12450), .B(n12451), .Z(n12421) );
  NAND U20681 ( .A(n12452), .B(n12453), .Z(n12451) );
  OR U20682 ( .A(n12454), .B(n12455), .Z(n12452) );
  NANDN U20683 ( .A(n12456), .B(n12454), .Z(n12450) );
  NAND U20684 ( .A(n12457), .B(n12458), .Z(n12425) );
  NANDN U20685 ( .A(n12459), .B(n12460), .Z(n12458) );
  OR U20686 ( .A(n12461), .B(n12462), .Z(n12460) );
  NANDN U20687 ( .A(n12463), .B(n12461), .Z(n12457) );
  IV U20688 ( .A(n12462), .Z(n12463) );
  XNOR U20689 ( .A(n12433), .B(n12464), .Z(n12428) );
  XNOR U20690 ( .A(n12431), .B(n12434), .Z(n12464) );
  NAND U20691 ( .A(n12465), .B(n12466), .Z(n12434) );
  NAND U20692 ( .A(n12467), .B(n12468), .Z(n12466) );
  OR U20693 ( .A(n12469), .B(n12470), .Z(n12467) );
  NANDN U20694 ( .A(n12471), .B(n12469), .Z(n12465) );
  IV U20695 ( .A(n12470), .Z(n12471) );
  NAND U20696 ( .A(n12472), .B(n12473), .Z(n12431) );
  NAND U20697 ( .A(n12474), .B(n12475), .Z(n12473) );
  NANDN U20698 ( .A(n12476), .B(n12477), .Z(n12474) );
  NANDN U20699 ( .A(n12477), .B(n12476), .Z(n12472) );
  AND U20700 ( .A(n12478), .B(n12479), .Z(n12433) );
  NAND U20701 ( .A(n12480), .B(n12481), .Z(n12479) );
  OR U20702 ( .A(n12482), .B(n12483), .Z(n12480) );
  NANDN U20703 ( .A(n12484), .B(n12482), .Z(n12478) );
  XNOR U20704 ( .A(n12459), .B(n12485), .Z(N64285) );
  XOR U20705 ( .A(n12461), .B(n12462), .Z(n12485) );
  XNOR U20706 ( .A(n12475), .B(n12486), .Z(n12462) );
  XOR U20707 ( .A(n12476), .B(n12477), .Z(n12486) );
  XOR U20708 ( .A(n12482), .B(n12487), .Z(n12477) );
  XOR U20709 ( .A(n12481), .B(n12484), .Z(n12487) );
  IV U20710 ( .A(n12483), .Z(n12484) );
  NAND U20711 ( .A(n12488), .B(n12489), .Z(n12483) );
  OR U20712 ( .A(n12490), .B(n12491), .Z(n12489) );
  OR U20713 ( .A(n12492), .B(n12493), .Z(n12488) );
  NAND U20714 ( .A(n12494), .B(n12495), .Z(n12481) );
  OR U20715 ( .A(n12496), .B(n12497), .Z(n12495) );
  OR U20716 ( .A(n12498), .B(n12499), .Z(n12494) );
  NOR U20717 ( .A(n12500), .B(n12501), .Z(n12482) );
  ANDN U20718 ( .B(n12502), .A(n12503), .Z(n12476) );
  XNOR U20719 ( .A(n12469), .B(n12504), .Z(n12475) );
  XNOR U20720 ( .A(n12468), .B(n12470), .Z(n12504) );
  NAND U20721 ( .A(n12505), .B(n12506), .Z(n12470) );
  OR U20722 ( .A(n12507), .B(n12508), .Z(n12506) );
  OR U20723 ( .A(n12509), .B(n12510), .Z(n12505) );
  NAND U20724 ( .A(n12511), .B(n12512), .Z(n12468) );
  OR U20725 ( .A(n12513), .B(n12514), .Z(n12512) );
  OR U20726 ( .A(n12515), .B(n12516), .Z(n12511) );
  ANDN U20727 ( .B(n12517), .A(n12518), .Z(n12469) );
  IV U20728 ( .A(n12519), .Z(n12517) );
  ANDN U20729 ( .B(n12520), .A(n12521), .Z(n12461) );
  XOR U20730 ( .A(n12447), .B(n12522), .Z(n12459) );
  XOR U20731 ( .A(n12448), .B(n12449), .Z(n12522) );
  XOR U20732 ( .A(n12454), .B(n12523), .Z(n12449) );
  XOR U20733 ( .A(n12453), .B(n12456), .Z(n12523) );
  IV U20734 ( .A(n12455), .Z(n12456) );
  NAND U20735 ( .A(n12524), .B(n12525), .Z(n12455) );
  OR U20736 ( .A(n12526), .B(n12527), .Z(n12525) );
  OR U20737 ( .A(n12528), .B(n12529), .Z(n12524) );
  NAND U20738 ( .A(n12530), .B(n12531), .Z(n12453) );
  OR U20739 ( .A(n12532), .B(n12533), .Z(n12531) );
  OR U20740 ( .A(n12534), .B(n12535), .Z(n12530) );
  NOR U20741 ( .A(n12536), .B(n12537), .Z(n12454) );
  ANDN U20742 ( .B(n12538), .A(n12539), .Z(n12448) );
  IV U20743 ( .A(n12540), .Z(n12538) );
  XNOR U20744 ( .A(n12441), .B(n12541), .Z(n12447) );
  XNOR U20745 ( .A(n12440), .B(n12442), .Z(n12541) );
  NAND U20746 ( .A(n12542), .B(n12543), .Z(n12442) );
  OR U20747 ( .A(n12544), .B(n12545), .Z(n12543) );
  OR U20748 ( .A(n12546), .B(n12547), .Z(n12542) );
  NAND U20749 ( .A(n12548), .B(n12549), .Z(n12440) );
  OR U20750 ( .A(n12550), .B(n12551), .Z(n12549) );
  OR U20751 ( .A(n12552), .B(n12553), .Z(n12548) );
  ANDN U20752 ( .B(n12554), .A(n12555), .Z(n12441) );
  IV U20753 ( .A(n12556), .Z(n12554) );
  XNOR U20754 ( .A(n12521), .B(n12520), .Z(N64284) );
  XOR U20755 ( .A(n12540), .B(n12539), .Z(n12520) );
  XNOR U20756 ( .A(n12555), .B(n12556), .Z(n12539) );
  XNOR U20757 ( .A(n12550), .B(n12551), .Z(n12556) );
  XNOR U20758 ( .A(n12552), .B(n12553), .Z(n12551) );
  XNOR U20759 ( .A(y[6829]), .B(x[6829]), .Z(n12553) );
  XNOR U20760 ( .A(y[6830]), .B(x[6830]), .Z(n12552) );
  XNOR U20761 ( .A(y[6828]), .B(x[6828]), .Z(n12550) );
  XNOR U20762 ( .A(n12544), .B(n12545), .Z(n12555) );
  XNOR U20763 ( .A(y[6825]), .B(x[6825]), .Z(n12545) );
  XNOR U20764 ( .A(n12546), .B(n12547), .Z(n12544) );
  XNOR U20765 ( .A(y[6826]), .B(x[6826]), .Z(n12547) );
  XNOR U20766 ( .A(y[6827]), .B(x[6827]), .Z(n12546) );
  XNOR U20767 ( .A(n12537), .B(n12536), .Z(n12540) );
  XNOR U20768 ( .A(n12532), .B(n12533), .Z(n12536) );
  XNOR U20769 ( .A(y[6822]), .B(x[6822]), .Z(n12533) );
  XNOR U20770 ( .A(n12534), .B(n12535), .Z(n12532) );
  XNOR U20771 ( .A(y[6823]), .B(x[6823]), .Z(n12535) );
  XNOR U20772 ( .A(y[6824]), .B(x[6824]), .Z(n12534) );
  XNOR U20773 ( .A(n12526), .B(n12527), .Z(n12537) );
  XNOR U20774 ( .A(y[6819]), .B(x[6819]), .Z(n12527) );
  XNOR U20775 ( .A(n12528), .B(n12529), .Z(n12526) );
  XNOR U20776 ( .A(y[6820]), .B(x[6820]), .Z(n12529) );
  XNOR U20777 ( .A(y[6821]), .B(x[6821]), .Z(n12528) );
  XOR U20778 ( .A(n12502), .B(n12503), .Z(n12521) );
  XNOR U20779 ( .A(n12518), .B(n12519), .Z(n12503) );
  XNOR U20780 ( .A(n12513), .B(n12514), .Z(n12519) );
  XNOR U20781 ( .A(n12515), .B(n12516), .Z(n12514) );
  XNOR U20782 ( .A(y[6817]), .B(x[6817]), .Z(n12516) );
  XNOR U20783 ( .A(y[6818]), .B(x[6818]), .Z(n12515) );
  XNOR U20784 ( .A(y[6816]), .B(x[6816]), .Z(n12513) );
  XNOR U20785 ( .A(n12507), .B(n12508), .Z(n12518) );
  XNOR U20786 ( .A(y[6813]), .B(x[6813]), .Z(n12508) );
  XNOR U20787 ( .A(n12509), .B(n12510), .Z(n12507) );
  XNOR U20788 ( .A(y[6814]), .B(x[6814]), .Z(n12510) );
  XNOR U20789 ( .A(y[6815]), .B(x[6815]), .Z(n12509) );
  XOR U20790 ( .A(n12501), .B(n12500), .Z(n12502) );
  XNOR U20791 ( .A(n12496), .B(n12497), .Z(n12500) );
  XNOR U20792 ( .A(y[6810]), .B(x[6810]), .Z(n12497) );
  XNOR U20793 ( .A(n12498), .B(n12499), .Z(n12496) );
  XNOR U20794 ( .A(y[6811]), .B(x[6811]), .Z(n12499) );
  XNOR U20795 ( .A(y[6812]), .B(x[6812]), .Z(n12498) );
  XNOR U20796 ( .A(n12490), .B(n12491), .Z(n12501) );
  XNOR U20797 ( .A(y[6807]), .B(x[6807]), .Z(n12491) );
  XNOR U20798 ( .A(n12492), .B(n12493), .Z(n12490) );
  XNOR U20799 ( .A(y[6808]), .B(x[6808]), .Z(n12493) );
  XNOR U20800 ( .A(y[6809]), .B(x[6809]), .Z(n12492) );
  NAND U20801 ( .A(n12557), .B(n12558), .Z(N64275) );
  NANDN U20802 ( .A(n12559), .B(n12560), .Z(n12558) );
  OR U20803 ( .A(n12561), .B(n12562), .Z(n12560) );
  NAND U20804 ( .A(n12561), .B(n12562), .Z(n12557) );
  XOR U20805 ( .A(n12561), .B(n12563), .Z(N64274) );
  XNOR U20806 ( .A(n12559), .B(n12562), .Z(n12563) );
  AND U20807 ( .A(n12564), .B(n12565), .Z(n12562) );
  NANDN U20808 ( .A(n12566), .B(n12567), .Z(n12565) );
  NANDN U20809 ( .A(n12568), .B(n12569), .Z(n12567) );
  NANDN U20810 ( .A(n12569), .B(n12568), .Z(n12564) );
  NAND U20811 ( .A(n12570), .B(n12571), .Z(n12559) );
  NANDN U20812 ( .A(n12572), .B(n12573), .Z(n12571) );
  OR U20813 ( .A(n12574), .B(n12575), .Z(n12573) );
  NAND U20814 ( .A(n12575), .B(n12574), .Z(n12570) );
  AND U20815 ( .A(n12576), .B(n12577), .Z(n12561) );
  NANDN U20816 ( .A(n12578), .B(n12579), .Z(n12577) );
  NANDN U20817 ( .A(n12580), .B(n12581), .Z(n12579) );
  NANDN U20818 ( .A(n12581), .B(n12580), .Z(n12576) );
  XOR U20819 ( .A(n12575), .B(n12582), .Z(N64273) );
  XOR U20820 ( .A(n12572), .B(n12574), .Z(n12582) );
  XNOR U20821 ( .A(n12568), .B(n12583), .Z(n12574) );
  XNOR U20822 ( .A(n12566), .B(n12569), .Z(n12583) );
  NAND U20823 ( .A(n12584), .B(n12585), .Z(n12569) );
  NAND U20824 ( .A(n12586), .B(n12587), .Z(n12585) );
  OR U20825 ( .A(n12588), .B(n12589), .Z(n12586) );
  NANDN U20826 ( .A(n12590), .B(n12588), .Z(n12584) );
  IV U20827 ( .A(n12589), .Z(n12590) );
  NAND U20828 ( .A(n12591), .B(n12592), .Z(n12566) );
  NAND U20829 ( .A(n12593), .B(n12594), .Z(n12592) );
  NANDN U20830 ( .A(n12595), .B(n12596), .Z(n12593) );
  NANDN U20831 ( .A(n12596), .B(n12595), .Z(n12591) );
  AND U20832 ( .A(n12597), .B(n12598), .Z(n12568) );
  NAND U20833 ( .A(n12599), .B(n12600), .Z(n12598) );
  OR U20834 ( .A(n12601), .B(n12602), .Z(n12599) );
  NANDN U20835 ( .A(n12603), .B(n12601), .Z(n12597) );
  NAND U20836 ( .A(n12604), .B(n12605), .Z(n12572) );
  NANDN U20837 ( .A(n12606), .B(n12607), .Z(n12605) );
  OR U20838 ( .A(n12608), .B(n12609), .Z(n12607) );
  NANDN U20839 ( .A(n12610), .B(n12608), .Z(n12604) );
  IV U20840 ( .A(n12609), .Z(n12610) );
  XNOR U20841 ( .A(n12580), .B(n12611), .Z(n12575) );
  XNOR U20842 ( .A(n12578), .B(n12581), .Z(n12611) );
  NAND U20843 ( .A(n12612), .B(n12613), .Z(n12581) );
  NAND U20844 ( .A(n12614), .B(n12615), .Z(n12613) );
  OR U20845 ( .A(n12616), .B(n12617), .Z(n12614) );
  NANDN U20846 ( .A(n12618), .B(n12616), .Z(n12612) );
  IV U20847 ( .A(n12617), .Z(n12618) );
  NAND U20848 ( .A(n12619), .B(n12620), .Z(n12578) );
  NAND U20849 ( .A(n12621), .B(n12622), .Z(n12620) );
  NANDN U20850 ( .A(n12623), .B(n12624), .Z(n12621) );
  NANDN U20851 ( .A(n12624), .B(n12623), .Z(n12619) );
  AND U20852 ( .A(n12625), .B(n12626), .Z(n12580) );
  NAND U20853 ( .A(n12627), .B(n12628), .Z(n12626) );
  OR U20854 ( .A(n12629), .B(n12630), .Z(n12627) );
  NANDN U20855 ( .A(n12631), .B(n12629), .Z(n12625) );
  XNOR U20856 ( .A(n12606), .B(n12632), .Z(N64272) );
  XOR U20857 ( .A(n12608), .B(n12609), .Z(n12632) );
  XNOR U20858 ( .A(n12622), .B(n12633), .Z(n12609) );
  XOR U20859 ( .A(n12623), .B(n12624), .Z(n12633) );
  XOR U20860 ( .A(n12629), .B(n12634), .Z(n12624) );
  XOR U20861 ( .A(n12628), .B(n12631), .Z(n12634) );
  IV U20862 ( .A(n12630), .Z(n12631) );
  NAND U20863 ( .A(n12635), .B(n12636), .Z(n12630) );
  OR U20864 ( .A(n12637), .B(n12638), .Z(n12636) );
  OR U20865 ( .A(n12639), .B(n12640), .Z(n12635) );
  NAND U20866 ( .A(n12641), .B(n12642), .Z(n12628) );
  OR U20867 ( .A(n12643), .B(n12644), .Z(n12642) );
  OR U20868 ( .A(n12645), .B(n12646), .Z(n12641) );
  NOR U20869 ( .A(n12647), .B(n12648), .Z(n12629) );
  ANDN U20870 ( .B(n12649), .A(n12650), .Z(n12623) );
  XNOR U20871 ( .A(n12616), .B(n12651), .Z(n12622) );
  XNOR U20872 ( .A(n12615), .B(n12617), .Z(n12651) );
  NAND U20873 ( .A(n12652), .B(n12653), .Z(n12617) );
  OR U20874 ( .A(n12654), .B(n12655), .Z(n12653) );
  OR U20875 ( .A(n12656), .B(n12657), .Z(n12652) );
  NAND U20876 ( .A(n12658), .B(n12659), .Z(n12615) );
  OR U20877 ( .A(n12660), .B(n12661), .Z(n12659) );
  OR U20878 ( .A(n12662), .B(n12663), .Z(n12658) );
  ANDN U20879 ( .B(n12664), .A(n12665), .Z(n12616) );
  IV U20880 ( .A(n12666), .Z(n12664) );
  ANDN U20881 ( .B(n12667), .A(n12668), .Z(n12608) );
  XOR U20882 ( .A(n12594), .B(n12669), .Z(n12606) );
  XOR U20883 ( .A(n12595), .B(n12596), .Z(n12669) );
  XOR U20884 ( .A(n12601), .B(n12670), .Z(n12596) );
  XOR U20885 ( .A(n12600), .B(n12603), .Z(n12670) );
  IV U20886 ( .A(n12602), .Z(n12603) );
  NAND U20887 ( .A(n12671), .B(n12672), .Z(n12602) );
  OR U20888 ( .A(n12673), .B(n12674), .Z(n12672) );
  OR U20889 ( .A(n12675), .B(n12676), .Z(n12671) );
  NAND U20890 ( .A(n12677), .B(n12678), .Z(n12600) );
  OR U20891 ( .A(n12679), .B(n12680), .Z(n12678) );
  OR U20892 ( .A(n12681), .B(n12682), .Z(n12677) );
  NOR U20893 ( .A(n12683), .B(n12684), .Z(n12601) );
  ANDN U20894 ( .B(n12685), .A(n12686), .Z(n12595) );
  IV U20895 ( .A(n12687), .Z(n12685) );
  XNOR U20896 ( .A(n12588), .B(n12688), .Z(n12594) );
  XNOR U20897 ( .A(n12587), .B(n12589), .Z(n12688) );
  NAND U20898 ( .A(n12689), .B(n12690), .Z(n12589) );
  OR U20899 ( .A(n12691), .B(n12692), .Z(n12690) );
  OR U20900 ( .A(n12693), .B(n12694), .Z(n12689) );
  NAND U20901 ( .A(n12695), .B(n12696), .Z(n12587) );
  OR U20902 ( .A(n12697), .B(n12698), .Z(n12696) );
  OR U20903 ( .A(n12699), .B(n12700), .Z(n12695) );
  ANDN U20904 ( .B(n12701), .A(n12702), .Z(n12588) );
  IV U20905 ( .A(n12703), .Z(n12701) );
  XNOR U20906 ( .A(n12668), .B(n12667), .Z(N64271) );
  XOR U20907 ( .A(n12687), .B(n12686), .Z(n12667) );
  XNOR U20908 ( .A(n12702), .B(n12703), .Z(n12686) );
  XNOR U20909 ( .A(n12697), .B(n12698), .Z(n12703) );
  XNOR U20910 ( .A(n12699), .B(n12700), .Z(n12698) );
  XNOR U20911 ( .A(y[6805]), .B(x[6805]), .Z(n12700) );
  XNOR U20912 ( .A(y[6806]), .B(x[6806]), .Z(n12699) );
  XNOR U20913 ( .A(y[6804]), .B(x[6804]), .Z(n12697) );
  XNOR U20914 ( .A(n12691), .B(n12692), .Z(n12702) );
  XNOR U20915 ( .A(y[6801]), .B(x[6801]), .Z(n12692) );
  XNOR U20916 ( .A(n12693), .B(n12694), .Z(n12691) );
  XNOR U20917 ( .A(y[6802]), .B(x[6802]), .Z(n12694) );
  XNOR U20918 ( .A(y[6803]), .B(x[6803]), .Z(n12693) );
  XNOR U20919 ( .A(n12684), .B(n12683), .Z(n12687) );
  XNOR U20920 ( .A(n12679), .B(n12680), .Z(n12683) );
  XNOR U20921 ( .A(y[6798]), .B(x[6798]), .Z(n12680) );
  XNOR U20922 ( .A(n12681), .B(n12682), .Z(n12679) );
  XNOR U20923 ( .A(y[6799]), .B(x[6799]), .Z(n12682) );
  XNOR U20924 ( .A(y[6800]), .B(x[6800]), .Z(n12681) );
  XNOR U20925 ( .A(n12673), .B(n12674), .Z(n12684) );
  XNOR U20926 ( .A(y[6795]), .B(x[6795]), .Z(n12674) );
  XNOR U20927 ( .A(n12675), .B(n12676), .Z(n12673) );
  XNOR U20928 ( .A(y[6796]), .B(x[6796]), .Z(n12676) );
  XNOR U20929 ( .A(y[6797]), .B(x[6797]), .Z(n12675) );
  XOR U20930 ( .A(n12649), .B(n12650), .Z(n12668) );
  XNOR U20931 ( .A(n12665), .B(n12666), .Z(n12650) );
  XNOR U20932 ( .A(n12660), .B(n12661), .Z(n12666) );
  XNOR U20933 ( .A(n12662), .B(n12663), .Z(n12661) );
  XNOR U20934 ( .A(y[6793]), .B(x[6793]), .Z(n12663) );
  XNOR U20935 ( .A(y[6794]), .B(x[6794]), .Z(n12662) );
  XNOR U20936 ( .A(y[6792]), .B(x[6792]), .Z(n12660) );
  XNOR U20937 ( .A(n12654), .B(n12655), .Z(n12665) );
  XNOR U20938 ( .A(y[6789]), .B(x[6789]), .Z(n12655) );
  XNOR U20939 ( .A(n12656), .B(n12657), .Z(n12654) );
  XNOR U20940 ( .A(y[6790]), .B(x[6790]), .Z(n12657) );
  XNOR U20941 ( .A(y[6791]), .B(x[6791]), .Z(n12656) );
  XOR U20942 ( .A(n12648), .B(n12647), .Z(n12649) );
  XNOR U20943 ( .A(n12643), .B(n12644), .Z(n12647) );
  XNOR U20944 ( .A(y[6786]), .B(x[6786]), .Z(n12644) );
  XNOR U20945 ( .A(n12645), .B(n12646), .Z(n12643) );
  XNOR U20946 ( .A(y[6787]), .B(x[6787]), .Z(n12646) );
  XNOR U20947 ( .A(y[6788]), .B(x[6788]), .Z(n12645) );
  XNOR U20948 ( .A(n12637), .B(n12638), .Z(n12648) );
  XNOR U20949 ( .A(y[6783]), .B(x[6783]), .Z(n12638) );
  XNOR U20950 ( .A(n12639), .B(n12640), .Z(n12637) );
  XNOR U20951 ( .A(y[6784]), .B(x[6784]), .Z(n12640) );
  XNOR U20952 ( .A(y[6785]), .B(x[6785]), .Z(n12639) );
  NAND U20953 ( .A(n12704), .B(n12705), .Z(N64262) );
  NANDN U20954 ( .A(n12706), .B(n12707), .Z(n12705) );
  OR U20955 ( .A(n12708), .B(n12709), .Z(n12707) );
  NAND U20956 ( .A(n12708), .B(n12709), .Z(n12704) );
  XOR U20957 ( .A(n12708), .B(n12710), .Z(N64261) );
  XNOR U20958 ( .A(n12706), .B(n12709), .Z(n12710) );
  AND U20959 ( .A(n12711), .B(n12712), .Z(n12709) );
  NANDN U20960 ( .A(n12713), .B(n12714), .Z(n12712) );
  NANDN U20961 ( .A(n12715), .B(n12716), .Z(n12714) );
  NANDN U20962 ( .A(n12716), .B(n12715), .Z(n12711) );
  NAND U20963 ( .A(n12717), .B(n12718), .Z(n12706) );
  NANDN U20964 ( .A(n12719), .B(n12720), .Z(n12718) );
  OR U20965 ( .A(n12721), .B(n12722), .Z(n12720) );
  NAND U20966 ( .A(n12722), .B(n12721), .Z(n12717) );
  AND U20967 ( .A(n12723), .B(n12724), .Z(n12708) );
  NANDN U20968 ( .A(n12725), .B(n12726), .Z(n12724) );
  NANDN U20969 ( .A(n12727), .B(n12728), .Z(n12726) );
  NANDN U20970 ( .A(n12728), .B(n12727), .Z(n12723) );
  XOR U20971 ( .A(n12722), .B(n12729), .Z(N64260) );
  XOR U20972 ( .A(n12719), .B(n12721), .Z(n12729) );
  XNOR U20973 ( .A(n12715), .B(n12730), .Z(n12721) );
  XNOR U20974 ( .A(n12713), .B(n12716), .Z(n12730) );
  NAND U20975 ( .A(n12731), .B(n12732), .Z(n12716) );
  NAND U20976 ( .A(n12733), .B(n12734), .Z(n12732) );
  OR U20977 ( .A(n12735), .B(n12736), .Z(n12733) );
  NANDN U20978 ( .A(n12737), .B(n12735), .Z(n12731) );
  IV U20979 ( .A(n12736), .Z(n12737) );
  NAND U20980 ( .A(n12738), .B(n12739), .Z(n12713) );
  NAND U20981 ( .A(n12740), .B(n12741), .Z(n12739) );
  NANDN U20982 ( .A(n12742), .B(n12743), .Z(n12740) );
  NANDN U20983 ( .A(n12743), .B(n12742), .Z(n12738) );
  AND U20984 ( .A(n12744), .B(n12745), .Z(n12715) );
  NAND U20985 ( .A(n12746), .B(n12747), .Z(n12745) );
  OR U20986 ( .A(n12748), .B(n12749), .Z(n12746) );
  NANDN U20987 ( .A(n12750), .B(n12748), .Z(n12744) );
  NAND U20988 ( .A(n12751), .B(n12752), .Z(n12719) );
  NANDN U20989 ( .A(n12753), .B(n12754), .Z(n12752) );
  OR U20990 ( .A(n12755), .B(n12756), .Z(n12754) );
  NANDN U20991 ( .A(n12757), .B(n12755), .Z(n12751) );
  IV U20992 ( .A(n12756), .Z(n12757) );
  XNOR U20993 ( .A(n12727), .B(n12758), .Z(n12722) );
  XNOR U20994 ( .A(n12725), .B(n12728), .Z(n12758) );
  NAND U20995 ( .A(n12759), .B(n12760), .Z(n12728) );
  NAND U20996 ( .A(n12761), .B(n12762), .Z(n12760) );
  OR U20997 ( .A(n12763), .B(n12764), .Z(n12761) );
  NANDN U20998 ( .A(n12765), .B(n12763), .Z(n12759) );
  IV U20999 ( .A(n12764), .Z(n12765) );
  NAND U21000 ( .A(n12766), .B(n12767), .Z(n12725) );
  NAND U21001 ( .A(n12768), .B(n12769), .Z(n12767) );
  NANDN U21002 ( .A(n12770), .B(n12771), .Z(n12768) );
  NANDN U21003 ( .A(n12771), .B(n12770), .Z(n12766) );
  AND U21004 ( .A(n12772), .B(n12773), .Z(n12727) );
  NAND U21005 ( .A(n12774), .B(n12775), .Z(n12773) );
  OR U21006 ( .A(n12776), .B(n12777), .Z(n12774) );
  NANDN U21007 ( .A(n12778), .B(n12776), .Z(n12772) );
  XNOR U21008 ( .A(n12753), .B(n12779), .Z(N64259) );
  XOR U21009 ( .A(n12755), .B(n12756), .Z(n12779) );
  XNOR U21010 ( .A(n12769), .B(n12780), .Z(n12756) );
  XOR U21011 ( .A(n12770), .B(n12771), .Z(n12780) );
  XOR U21012 ( .A(n12776), .B(n12781), .Z(n12771) );
  XOR U21013 ( .A(n12775), .B(n12778), .Z(n12781) );
  IV U21014 ( .A(n12777), .Z(n12778) );
  NAND U21015 ( .A(n12782), .B(n12783), .Z(n12777) );
  OR U21016 ( .A(n12784), .B(n12785), .Z(n12783) );
  OR U21017 ( .A(n12786), .B(n12787), .Z(n12782) );
  NAND U21018 ( .A(n12788), .B(n12789), .Z(n12775) );
  OR U21019 ( .A(n12790), .B(n12791), .Z(n12789) );
  OR U21020 ( .A(n12792), .B(n12793), .Z(n12788) );
  NOR U21021 ( .A(n12794), .B(n12795), .Z(n12776) );
  ANDN U21022 ( .B(n12796), .A(n12797), .Z(n12770) );
  XNOR U21023 ( .A(n12763), .B(n12798), .Z(n12769) );
  XNOR U21024 ( .A(n12762), .B(n12764), .Z(n12798) );
  NAND U21025 ( .A(n12799), .B(n12800), .Z(n12764) );
  OR U21026 ( .A(n12801), .B(n12802), .Z(n12800) );
  OR U21027 ( .A(n12803), .B(n12804), .Z(n12799) );
  NAND U21028 ( .A(n12805), .B(n12806), .Z(n12762) );
  OR U21029 ( .A(n12807), .B(n12808), .Z(n12806) );
  OR U21030 ( .A(n12809), .B(n12810), .Z(n12805) );
  ANDN U21031 ( .B(n12811), .A(n12812), .Z(n12763) );
  IV U21032 ( .A(n12813), .Z(n12811) );
  ANDN U21033 ( .B(n12814), .A(n12815), .Z(n12755) );
  XOR U21034 ( .A(n12741), .B(n12816), .Z(n12753) );
  XOR U21035 ( .A(n12742), .B(n12743), .Z(n12816) );
  XOR U21036 ( .A(n12748), .B(n12817), .Z(n12743) );
  XOR U21037 ( .A(n12747), .B(n12750), .Z(n12817) );
  IV U21038 ( .A(n12749), .Z(n12750) );
  NAND U21039 ( .A(n12818), .B(n12819), .Z(n12749) );
  OR U21040 ( .A(n12820), .B(n12821), .Z(n12819) );
  OR U21041 ( .A(n12822), .B(n12823), .Z(n12818) );
  NAND U21042 ( .A(n12824), .B(n12825), .Z(n12747) );
  OR U21043 ( .A(n12826), .B(n12827), .Z(n12825) );
  OR U21044 ( .A(n12828), .B(n12829), .Z(n12824) );
  NOR U21045 ( .A(n12830), .B(n12831), .Z(n12748) );
  ANDN U21046 ( .B(n12832), .A(n12833), .Z(n12742) );
  IV U21047 ( .A(n12834), .Z(n12832) );
  XNOR U21048 ( .A(n12735), .B(n12835), .Z(n12741) );
  XNOR U21049 ( .A(n12734), .B(n12736), .Z(n12835) );
  NAND U21050 ( .A(n12836), .B(n12837), .Z(n12736) );
  OR U21051 ( .A(n12838), .B(n12839), .Z(n12837) );
  OR U21052 ( .A(n12840), .B(n12841), .Z(n12836) );
  NAND U21053 ( .A(n12842), .B(n12843), .Z(n12734) );
  OR U21054 ( .A(n12844), .B(n12845), .Z(n12843) );
  OR U21055 ( .A(n12846), .B(n12847), .Z(n12842) );
  ANDN U21056 ( .B(n12848), .A(n12849), .Z(n12735) );
  IV U21057 ( .A(n12850), .Z(n12848) );
  XNOR U21058 ( .A(n12815), .B(n12814), .Z(N64258) );
  XOR U21059 ( .A(n12834), .B(n12833), .Z(n12814) );
  XNOR U21060 ( .A(n12849), .B(n12850), .Z(n12833) );
  XNOR U21061 ( .A(n12844), .B(n12845), .Z(n12850) );
  XNOR U21062 ( .A(n12846), .B(n12847), .Z(n12845) );
  XNOR U21063 ( .A(y[6781]), .B(x[6781]), .Z(n12847) );
  XNOR U21064 ( .A(y[6782]), .B(x[6782]), .Z(n12846) );
  XNOR U21065 ( .A(y[6780]), .B(x[6780]), .Z(n12844) );
  XNOR U21066 ( .A(n12838), .B(n12839), .Z(n12849) );
  XNOR U21067 ( .A(y[6777]), .B(x[6777]), .Z(n12839) );
  XNOR U21068 ( .A(n12840), .B(n12841), .Z(n12838) );
  XNOR U21069 ( .A(y[6778]), .B(x[6778]), .Z(n12841) );
  XNOR U21070 ( .A(y[6779]), .B(x[6779]), .Z(n12840) );
  XNOR U21071 ( .A(n12831), .B(n12830), .Z(n12834) );
  XNOR U21072 ( .A(n12826), .B(n12827), .Z(n12830) );
  XNOR U21073 ( .A(y[6774]), .B(x[6774]), .Z(n12827) );
  XNOR U21074 ( .A(n12828), .B(n12829), .Z(n12826) );
  XNOR U21075 ( .A(y[6775]), .B(x[6775]), .Z(n12829) );
  XNOR U21076 ( .A(y[6776]), .B(x[6776]), .Z(n12828) );
  XNOR U21077 ( .A(n12820), .B(n12821), .Z(n12831) );
  XNOR U21078 ( .A(y[6771]), .B(x[6771]), .Z(n12821) );
  XNOR U21079 ( .A(n12822), .B(n12823), .Z(n12820) );
  XNOR U21080 ( .A(y[6772]), .B(x[6772]), .Z(n12823) );
  XNOR U21081 ( .A(y[6773]), .B(x[6773]), .Z(n12822) );
  XOR U21082 ( .A(n12796), .B(n12797), .Z(n12815) );
  XNOR U21083 ( .A(n12812), .B(n12813), .Z(n12797) );
  XNOR U21084 ( .A(n12807), .B(n12808), .Z(n12813) );
  XNOR U21085 ( .A(n12809), .B(n12810), .Z(n12808) );
  XNOR U21086 ( .A(y[6769]), .B(x[6769]), .Z(n12810) );
  XNOR U21087 ( .A(y[6770]), .B(x[6770]), .Z(n12809) );
  XNOR U21088 ( .A(y[6768]), .B(x[6768]), .Z(n12807) );
  XNOR U21089 ( .A(n12801), .B(n12802), .Z(n12812) );
  XNOR U21090 ( .A(y[6765]), .B(x[6765]), .Z(n12802) );
  XNOR U21091 ( .A(n12803), .B(n12804), .Z(n12801) );
  XNOR U21092 ( .A(y[6766]), .B(x[6766]), .Z(n12804) );
  XNOR U21093 ( .A(y[6767]), .B(x[6767]), .Z(n12803) );
  XOR U21094 ( .A(n12795), .B(n12794), .Z(n12796) );
  XNOR U21095 ( .A(n12790), .B(n12791), .Z(n12794) );
  XNOR U21096 ( .A(y[6762]), .B(x[6762]), .Z(n12791) );
  XNOR U21097 ( .A(n12792), .B(n12793), .Z(n12790) );
  XNOR U21098 ( .A(y[6763]), .B(x[6763]), .Z(n12793) );
  XNOR U21099 ( .A(y[6764]), .B(x[6764]), .Z(n12792) );
  XNOR U21100 ( .A(n12784), .B(n12785), .Z(n12795) );
  XNOR U21101 ( .A(y[6759]), .B(x[6759]), .Z(n12785) );
  XNOR U21102 ( .A(n12786), .B(n12787), .Z(n12784) );
  XNOR U21103 ( .A(y[6760]), .B(x[6760]), .Z(n12787) );
  XNOR U21104 ( .A(y[6761]), .B(x[6761]), .Z(n12786) );
  NAND U21105 ( .A(n12851), .B(n12852), .Z(N64249) );
  NANDN U21106 ( .A(n12853), .B(n12854), .Z(n12852) );
  OR U21107 ( .A(n12855), .B(n12856), .Z(n12854) );
  NAND U21108 ( .A(n12855), .B(n12856), .Z(n12851) );
  XOR U21109 ( .A(n12855), .B(n12857), .Z(N64248) );
  XNOR U21110 ( .A(n12853), .B(n12856), .Z(n12857) );
  AND U21111 ( .A(n12858), .B(n12859), .Z(n12856) );
  NANDN U21112 ( .A(n12860), .B(n12861), .Z(n12859) );
  NANDN U21113 ( .A(n12862), .B(n12863), .Z(n12861) );
  NANDN U21114 ( .A(n12863), .B(n12862), .Z(n12858) );
  NAND U21115 ( .A(n12864), .B(n12865), .Z(n12853) );
  NANDN U21116 ( .A(n12866), .B(n12867), .Z(n12865) );
  OR U21117 ( .A(n12868), .B(n12869), .Z(n12867) );
  NAND U21118 ( .A(n12869), .B(n12868), .Z(n12864) );
  AND U21119 ( .A(n12870), .B(n12871), .Z(n12855) );
  NANDN U21120 ( .A(n12872), .B(n12873), .Z(n12871) );
  NANDN U21121 ( .A(n12874), .B(n12875), .Z(n12873) );
  NANDN U21122 ( .A(n12875), .B(n12874), .Z(n12870) );
  XOR U21123 ( .A(n12869), .B(n12876), .Z(N64247) );
  XOR U21124 ( .A(n12866), .B(n12868), .Z(n12876) );
  XNOR U21125 ( .A(n12862), .B(n12877), .Z(n12868) );
  XNOR U21126 ( .A(n12860), .B(n12863), .Z(n12877) );
  NAND U21127 ( .A(n12878), .B(n12879), .Z(n12863) );
  NAND U21128 ( .A(n12880), .B(n12881), .Z(n12879) );
  OR U21129 ( .A(n12882), .B(n12883), .Z(n12880) );
  NANDN U21130 ( .A(n12884), .B(n12882), .Z(n12878) );
  IV U21131 ( .A(n12883), .Z(n12884) );
  NAND U21132 ( .A(n12885), .B(n12886), .Z(n12860) );
  NAND U21133 ( .A(n12887), .B(n12888), .Z(n12886) );
  NANDN U21134 ( .A(n12889), .B(n12890), .Z(n12887) );
  NANDN U21135 ( .A(n12890), .B(n12889), .Z(n12885) );
  AND U21136 ( .A(n12891), .B(n12892), .Z(n12862) );
  NAND U21137 ( .A(n12893), .B(n12894), .Z(n12892) );
  OR U21138 ( .A(n12895), .B(n12896), .Z(n12893) );
  NANDN U21139 ( .A(n12897), .B(n12895), .Z(n12891) );
  NAND U21140 ( .A(n12898), .B(n12899), .Z(n12866) );
  NANDN U21141 ( .A(n12900), .B(n12901), .Z(n12899) );
  OR U21142 ( .A(n12902), .B(n12903), .Z(n12901) );
  NANDN U21143 ( .A(n12904), .B(n12902), .Z(n12898) );
  IV U21144 ( .A(n12903), .Z(n12904) );
  XNOR U21145 ( .A(n12874), .B(n12905), .Z(n12869) );
  XNOR U21146 ( .A(n12872), .B(n12875), .Z(n12905) );
  NAND U21147 ( .A(n12906), .B(n12907), .Z(n12875) );
  NAND U21148 ( .A(n12908), .B(n12909), .Z(n12907) );
  OR U21149 ( .A(n12910), .B(n12911), .Z(n12908) );
  NANDN U21150 ( .A(n12912), .B(n12910), .Z(n12906) );
  IV U21151 ( .A(n12911), .Z(n12912) );
  NAND U21152 ( .A(n12913), .B(n12914), .Z(n12872) );
  NAND U21153 ( .A(n12915), .B(n12916), .Z(n12914) );
  NANDN U21154 ( .A(n12917), .B(n12918), .Z(n12915) );
  NANDN U21155 ( .A(n12918), .B(n12917), .Z(n12913) );
  AND U21156 ( .A(n12919), .B(n12920), .Z(n12874) );
  NAND U21157 ( .A(n12921), .B(n12922), .Z(n12920) );
  OR U21158 ( .A(n12923), .B(n12924), .Z(n12921) );
  NANDN U21159 ( .A(n12925), .B(n12923), .Z(n12919) );
  XNOR U21160 ( .A(n12900), .B(n12926), .Z(N64246) );
  XOR U21161 ( .A(n12902), .B(n12903), .Z(n12926) );
  XNOR U21162 ( .A(n12916), .B(n12927), .Z(n12903) );
  XOR U21163 ( .A(n12917), .B(n12918), .Z(n12927) );
  XOR U21164 ( .A(n12923), .B(n12928), .Z(n12918) );
  XOR U21165 ( .A(n12922), .B(n12925), .Z(n12928) );
  IV U21166 ( .A(n12924), .Z(n12925) );
  NAND U21167 ( .A(n12929), .B(n12930), .Z(n12924) );
  OR U21168 ( .A(n12931), .B(n12932), .Z(n12930) );
  OR U21169 ( .A(n12933), .B(n12934), .Z(n12929) );
  NAND U21170 ( .A(n12935), .B(n12936), .Z(n12922) );
  OR U21171 ( .A(n12937), .B(n12938), .Z(n12936) );
  OR U21172 ( .A(n12939), .B(n12940), .Z(n12935) );
  NOR U21173 ( .A(n12941), .B(n12942), .Z(n12923) );
  ANDN U21174 ( .B(n12943), .A(n12944), .Z(n12917) );
  XNOR U21175 ( .A(n12910), .B(n12945), .Z(n12916) );
  XNOR U21176 ( .A(n12909), .B(n12911), .Z(n12945) );
  NAND U21177 ( .A(n12946), .B(n12947), .Z(n12911) );
  OR U21178 ( .A(n12948), .B(n12949), .Z(n12947) );
  OR U21179 ( .A(n12950), .B(n12951), .Z(n12946) );
  NAND U21180 ( .A(n12952), .B(n12953), .Z(n12909) );
  OR U21181 ( .A(n12954), .B(n12955), .Z(n12953) );
  OR U21182 ( .A(n12956), .B(n12957), .Z(n12952) );
  ANDN U21183 ( .B(n12958), .A(n12959), .Z(n12910) );
  IV U21184 ( .A(n12960), .Z(n12958) );
  ANDN U21185 ( .B(n12961), .A(n12962), .Z(n12902) );
  XOR U21186 ( .A(n12888), .B(n12963), .Z(n12900) );
  XOR U21187 ( .A(n12889), .B(n12890), .Z(n12963) );
  XOR U21188 ( .A(n12895), .B(n12964), .Z(n12890) );
  XOR U21189 ( .A(n12894), .B(n12897), .Z(n12964) );
  IV U21190 ( .A(n12896), .Z(n12897) );
  NAND U21191 ( .A(n12965), .B(n12966), .Z(n12896) );
  OR U21192 ( .A(n12967), .B(n12968), .Z(n12966) );
  OR U21193 ( .A(n12969), .B(n12970), .Z(n12965) );
  NAND U21194 ( .A(n12971), .B(n12972), .Z(n12894) );
  OR U21195 ( .A(n12973), .B(n12974), .Z(n12972) );
  OR U21196 ( .A(n12975), .B(n12976), .Z(n12971) );
  NOR U21197 ( .A(n12977), .B(n12978), .Z(n12895) );
  ANDN U21198 ( .B(n12979), .A(n12980), .Z(n12889) );
  IV U21199 ( .A(n12981), .Z(n12979) );
  XNOR U21200 ( .A(n12882), .B(n12982), .Z(n12888) );
  XNOR U21201 ( .A(n12881), .B(n12883), .Z(n12982) );
  NAND U21202 ( .A(n12983), .B(n12984), .Z(n12883) );
  OR U21203 ( .A(n12985), .B(n12986), .Z(n12984) );
  OR U21204 ( .A(n12987), .B(n12988), .Z(n12983) );
  NAND U21205 ( .A(n12989), .B(n12990), .Z(n12881) );
  OR U21206 ( .A(n12991), .B(n12992), .Z(n12990) );
  OR U21207 ( .A(n12993), .B(n12994), .Z(n12989) );
  ANDN U21208 ( .B(n12995), .A(n12996), .Z(n12882) );
  IV U21209 ( .A(n12997), .Z(n12995) );
  XNOR U21210 ( .A(n12962), .B(n12961), .Z(N64245) );
  XOR U21211 ( .A(n12981), .B(n12980), .Z(n12961) );
  XNOR U21212 ( .A(n12996), .B(n12997), .Z(n12980) );
  XNOR U21213 ( .A(n12991), .B(n12992), .Z(n12997) );
  XNOR U21214 ( .A(n12993), .B(n12994), .Z(n12992) );
  XNOR U21215 ( .A(y[6757]), .B(x[6757]), .Z(n12994) );
  XNOR U21216 ( .A(y[6758]), .B(x[6758]), .Z(n12993) );
  XNOR U21217 ( .A(y[6756]), .B(x[6756]), .Z(n12991) );
  XNOR U21218 ( .A(n12985), .B(n12986), .Z(n12996) );
  XNOR U21219 ( .A(y[6753]), .B(x[6753]), .Z(n12986) );
  XNOR U21220 ( .A(n12987), .B(n12988), .Z(n12985) );
  XNOR U21221 ( .A(y[6754]), .B(x[6754]), .Z(n12988) );
  XNOR U21222 ( .A(y[6755]), .B(x[6755]), .Z(n12987) );
  XNOR U21223 ( .A(n12978), .B(n12977), .Z(n12981) );
  XNOR U21224 ( .A(n12973), .B(n12974), .Z(n12977) );
  XNOR U21225 ( .A(y[6750]), .B(x[6750]), .Z(n12974) );
  XNOR U21226 ( .A(n12975), .B(n12976), .Z(n12973) );
  XNOR U21227 ( .A(y[6751]), .B(x[6751]), .Z(n12976) );
  XNOR U21228 ( .A(y[6752]), .B(x[6752]), .Z(n12975) );
  XNOR U21229 ( .A(n12967), .B(n12968), .Z(n12978) );
  XNOR U21230 ( .A(y[6747]), .B(x[6747]), .Z(n12968) );
  XNOR U21231 ( .A(n12969), .B(n12970), .Z(n12967) );
  XNOR U21232 ( .A(y[6748]), .B(x[6748]), .Z(n12970) );
  XNOR U21233 ( .A(y[6749]), .B(x[6749]), .Z(n12969) );
  XOR U21234 ( .A(n12943), .B(n12944), .Z(n12962) );
  XNOR U21235 ( .A(n12959), .B(n12960), .Z(n12944) );
  XNOR U21236 ( .A(n12954), .B(n12955), .Z(n12960) );
  XNOR U21237 ( .A(n12956), .B(n12957), .Z(n12955) );
  XNOR U21238 ( .A(y[6745]), .B(x[6745]), .Z(n12957) );
  XNOR U21239 ( .A(y[6746]), .B(x[6746]), .Z(n12956) );
  XNOR U21240 ( .A(y[6744]), .B(x[6744]), .Z(n12954) );
  XNOR U21241 ( .A(n12948), .B(n12949), .Z(n12959) );
  XNOR U21242 ( .A(y[6741]), .B(x[6741]), .Z(n12949) );
  XNOR U21243 ( .A(n12950), .B(n12951), .Z(n12948) );
  XNOR U21244 ( .A(y[6742]), .B(x[6742]), .Z(n12951) );
  XNOR U21245 ( .A(y[6743]), .B(x[6743]), .Z(n12950) );
  XOR U21246 ( .A(n12942), .B(n12941), .Z(n12943) );
  XNOR U21247 ( .A(n12937), .B(n12938), .Z(n12941) );
  XNOR U21248 ( .A(y[6738]), .B(x[6738]), .Z(n12938) );
  XNOR U21249 ( .A(n12939), .B(n12940), .Z(n12937) );
  XNOR U21250 ( .A(y[6739]), .B(x[6739]), .Z(n12940) );
  XNOR U21251 ( .A(y[6740]), .B(x[6740]), .Z(n12939) );
  XNOR U21252 ( .A(n12931), .B(n12932), .Z(n12942) );
  XNOR U21253 ( .A(y[6735]), .B(x[6735]), .Z(n12932) );
  XNOR U21254 ( .A(n12933), .B(n12934), .Z(n12931) );
  XNOR U21255 ( .A(y[6736]), .B(x[6736]), .Z(n12934) );
  XNOR U21256 ( .A(y[6737]), .B(x[6737]), .Z(n12933) );
  NAND U21257 ( .A(n12998), .B(n12999), .Z(N64236) );
  NANDN U21258 ( .A(n13000), .B(n13001), .Z(n12999) );
  OR U21259 ( .A(n13002), .B(n13003), .Z(n13001) );
  NAND U21260 ( .A(n13002), .B(n13003), .Z(n12998) );
  XOR U21261 ( .A(n13002), .B(n13004), .Z(N64235) );
  XNOR U21262 ( .A(n13000), .B(n13003), .Z(n13004) );
  AND U21263 ( .A(n13005), .B(n13006), .Z(n13003) );
  NANDN U21264 ( .A(n13007), .B(n13008), .Z(n13006) );
  NANDN U21265 ( .A(n13009), .B(n13010), .Z(n13008) );
  NANDN U21266 ( .A(n13010), .B(n13009), .Z(n13005) );
  NAND U21267 ( .A(n13011), .B(n13012), .Z(n13000) );
  NANDN U21268 ( .A(n13013), .B(n13014), .Z(n13012) );
  OR U21269 ( .A(n13015), .B(n13016), .Z(n13014) );
  NAND U21270 ( .A(n13016), .B(n13015), .Z(n13011) );
  AND U21271 ( .A(n13017), .B(n13018), .Z(n13002) );
  NANDN U21272 ( .A(n13019), .B(n13020), .Z(n13018) );
  NANDN U21273 ( .A(n13021), .B(n13022), .Z(n13020) );
  NANDN U21274 ( .A(n13022), .B(n13021), .Z(n13017) );
  XOR U21275 ( .A(n13016), .B(n13023), .Z(N64234) );
  XOR U21276 ( .A(n13013), .B(n13015), .Z(n13023) );
  XNOR U21277 ( .A(n13009), .B(n13024), .Z(n13015) );
  XNOR U21278 ( .A(n13007), .B(n13010), .Z(n13024) );
  NAND U21279 ( .A(n13025), .B(n13026), .Z(n13010) );
  NAND U21280 ( .A(n13027), .B(n13028), .Z(n13026) );
  OR U21281 ( .A(n13029), .B(n13030), .Z(n13027) );
  NANDN U21282 ( .A(n13031), .B(n13029), .Z(n13025) );
  IV U21283 ( .A(n13030), .Z(n13031) );
  NAND U21284 ( .A(n13032), .B(n13033), .Z(n13007) );
  NAND U21285 ( .A(n13034), .B(n13035), .Z(n13033) );
  NANDN U21286 ( .A(n13036), .B(n13037), .Z(n13034) );
  NANDN U21287 ( .A(n13037), .B(n13036), .Z(n13032) );
  AND U21288 ( .A(n13038), .B(n13039), .Z(n13009) );
  NAND U21289 ( .A(n13040), .B(n13041), .Z(n13039) );
  OR U21290 ( .A(n13042), .B(n13043), .Z(n13040) );
  NANDN U21291 ( .A(n13044), .B(n13042), .Z(n13038) );
  NAND U21292 ( .A(n13045), .B(n13046), .Z(n13013) );
  NANDN U21293 ( .A(n13047), .B(n13048), .Z(n13046) );
  OR U21294 ( .A(n13049), .B(n13050), .Z(n13048) );
  NANDN U21295 ( .A(n13051), .B(n13049), .Z(n13045) );
  IV U21296 ( .A(n13050), .Z(n13051) );
  XNOR U21297 ( .A(n13021), .B(n13052), .Z(n13016) );
  XNOR U21298 ( .A(n13019), .B(n13022), .Z(n13052) );
  NAND U21299 ( .A(n13053), .B(n13054), .Z(n13022) );
  NAND U21300 ( .A(n13055), .B(n13056), .Z(n13054) );
  OR U21301 ( .A(n13057), .B(n13058), .Z(n13055) );
  NANDN U21302 ( .A(n13059), .B(n13057), .Z(n13053) );
  IV U21303 ( .A(n13058), .Z(n13059) );
  NAND U21304 ( .A(n13060), .B(n13061), .Z(n13019) );
  NAND U21305 ( .A(n13062), .B(n13063), .Z(n13061) );
  NANDN U21306 ( .A(n13064), .B(n13065), .Z(n13062) );
  NANDN U21307 ( .A(n13065), .B(n13064), .Z(n13060) );
  AND U21308 ( .A(n13066), .B(n13067), .Z(n13021) );
  NAND U21309 ( .A(n13068), .B(n13069), .Z(n13067) );
  OR U21310 ( .A(n13070), .B(n13071), .Z(n13068) );
  NANDN U21311 ( .A(n13072), .B(n13070), .Z(n13066) );
  XNOR U21312 ( .A(n13047), .B(n13073), .Z(N64233) );
  XOR U21313 ( .A(n13049), .B(n13050), .Z(n13073) );
  XNOR U21314 ( .A(n13063), .B(n13074), .Z(n13050) );
  XOR U21315 ( .A(n13064), .B(n13065), .Z(n13074) );
  XOR U21316 ( .A(n13070), .B(n13075), .Z(n13065) );
  XOR U21317 ( .A(n13069), .B(n13072), .Z(n13075) );
  IV U21318 ( .A(n13071), .Z(n13072) );
  NAND U21319 ( .A(n13076), .B(n13077), .Z(n13071) );
  OR U21320 ( .A(n13078), .B(n13079), .Z(n13077) );
  OR U21321 ( .A(n13080), .B(n13081), .Z(n13076) );
  NAND U21322 ( .A(n13082), .B(n13083), .Z(n13069) );
  OR U21323 ( .A(n13084), .B(n13085), .Z(n13083) );
  OR U21324 ( .A(n13086), .B(n13087), .Z(n13082) );
  NOR U21325 ( .A(n13088), .B(n13089), .Z(n13070) );
  ANDN U21326 ( .B(n13090), .A(n13091), .Z(n13064) );
  XNOR U21327 ( .A(n13057), .B(n13092), .Z(n13063) );
  XNOR U21328 ( .A(n13056), .B(n13058), .Z(n13092) );
  NAND U21329 ( .A(n13093), .B(n13094), .Z(n13058) );
  OR U21330 ( .A(n13095), .B(n13096), .Z(n13094) );
  OR U21331 ( .A(n13097), .B(n13098), .Z(n13093) );
  NAND U21332 ( .A(n13099), .B(n13100), .Z(n13056) );
  OR U21333 ( .A(n13101), .B(n13102), .Z(n13100) );
  OR U21334 ( .A(n13103), .B(n13104), .Z(n13099) );
  ANDN U21335 ( .B(n13105), .A(n13106), .Z(n13057) );
  IV U21336 ( .A(n13107), .Z(n13105) );
  ANDN U21337 ( .B(n13108), .A(n13109), .Z(n13049) );
  XOR U21338 ( .A(n13035), .B(n13110), .Z(n13047) );
  XOR U21339 ( .A(n13036), .B(n13037), .Z(n13110) );
  XOR U21340 ( .A(n13042), .B(n13111), .Z(n13037) );
  XOR U21341 ( .A(n13041), .B(n13044), .Z(n13111) );
  IV U21342 ( .A(n13043), .Z(n13044) );
  NAND U21343 ( .A(n13112), .B(n13113), .Z(n13043) );
  OR U21344 ( .A(n13114), .B(n13115), .Z(n13113) );
  OR U21345 ( .A(n13116), .B(n13117), .Z(n13112) );
  NAND U21346 ( .A(n13118), .B(n13119), .Z(n13041) );
  OR U21347 ( .A(n13120), .B(n13121), .Z(n13119) );
  OR U21348 ( .A(n13122), .B(n13123), .Z(n13118) );
  NOR U21349 ( .A(n13124), .B(n13125), .Z(n13042) );
  ANDN U21350 ( .B(n13126), .A(n13127), .Z(n13036) );
  IV U21351 ( .A(n13128), .Z(n13126) );
  XNOR U21352 ( .A(n13029), .B(n13129), .Z(n13035) );
  XNOR U21353 ( .A(n13028), .B(n13030), .Z(n13129) );
  NAND U21354 ( .A(n13130), .B(n13131), .Z(n13030) );
  OR U21355 ( .A(n13132), .B(n13133), .Z(n13131) );
  OR U21356 ( .A(n13134), .B(n13135), .Z(n13130) );
  NAND U21357 ( .A(n13136), .B(n13137), .Z(n13028) );
  OR U21358 ( .A(n13138), .B(n13139), .Z(n13137) );
  OR U21359 ( .A(n13140), .B(n13141), .Z(n13136) );
  ANDN U21360 ( .B(n13142), .A(n13143), .Z(n13029) );
  IV U21361 ( .A(n13144), .Z(n13142) );
  XNOR U21362 ( .A(n13109), .B(n13108), .Z(N64232) );
  XOR U21363 ( .A(n13128), .B(n13127), .Z(n13108) );
  XNOR U21364 ( .A(n13143), .B(n13144), .Z(n13127) );
  XNOR U21365 ( .A(n13138), .B(n13139), .Z(n13144) );
  XNOR U21366 ( .A(n13140), .B(n13141), .Z(n13139) );
  XNOR U21367 ( .A(y[6733]), .B(x[6733]), .Z(n13141) );
  XNOR U21368 ( .A(y[6734]), .B(x[6734]), .Z(n13140) );
  XNOR U21369 ( .A(y[6732]), .B(x[6732]), .Z(n13138) );
  XNOR U21370 ( .A(n13132), .B(n13133), .Z(n13143) );
  XNOR U21371 ( .A(y[6729]), .B(x[6729]), .Z(n13133) );
  XNOR U21372 ( .A(n13134), .B(n13135), .Z(n13132) );
  XNOR U21373 ( .A(y[6730]), .B(x[6730]), .Z(n13135) );
  XNOR U21374 ( .A(y[6731]), .B(x[6731]), .Z(n13134) );
  XNOR U21375 ( .A(n13125), .B(n13124), .Z(n13128) );
  XNOR U21376 ( .A(n13120), .B(n13121), .Z(n13124) );
  XNOR U21377 ( .A(y[6726]), .B(x[6726]), .Z(n13121) );
  XNOR U21378 ( .A(n13122), .B(n13123), .Z(n13120) );
  XNOR U21379 ( .A(y[6727]), .B(x[6727]), .Z(n13123) );
  XNOR U21380 ( .A(y[6728]), .B(x[6728]), .Z(n13122) );
  XNOR U21381 ( .A(n13114), .B(n13115), .Z(n13125) );
  XNOR U21382 ( .A(y[6723]), .B(x[6723]), .Z(n13115) );
  XNOR U21383 ( .A(n13116), .B(n13117), .Z(n13114) );
  XNOR U21384 ( .A(y[6724]), .B(x[6724]), .Z(n13117) );
  XNOR U21385 ( .A(y[6725]), .B(x[6725]), .Z(n13116) );
  XOR U21386 ( .A(n13090), .B(n13091), .Z(n13109) );
  XNOR U21387 ( .A(n13106), .B(n13107), .Z(n13091) );
  XNOR U21388 ( .A(n13101), .B(n13102), .Z(n13107) );
  XNOR U21389 ( .A(n13103), .B(n13104), .Z(n13102) );
  XNOR U21390 ( .A(y[6721]), .B(x[6721]), .Z(n13104) );
  XNOR U21391 ( .A(y[6722]), .B(x[6722]), .Z(n13103) );
  XNOR U21392 ( .A(y[6720]), .B(x[6720]), .Z(n13101) );
  XNOR U21393 ( .A(n13095), .B(n13096), .Z(n13106) );
  XNOR U21394 ( .A(y[6717]), .B(x[6717]), .Z(n13096) );
  XNOR U21395 ( .A(n13097), .B(n13098), .Z(n13095) );
  XNOR U21396 ( .A(y[6718]), .B(x[6718]), .Z(n13098) );
  XNOR U21397 ( .A(y[6719]), .B(x[6719]), .Z(n13097) );
  XOR U21398 ( .A(n13089), .B(n13088), .Z(n13090) );
  XNOR U21399 ( .A(n13084), .B(n13085), .Z(n13088) );
  XNOR U21400 ( .A(y[6714]), .B(x[6714]), .Z(n13085) );
  XNOR U21401 ( .A(n13086), .B(n13087), .Z(n13084) );
  XNOR U21402 ( .A(y[6715]), .B(x[6715]), .Z(n13087) );
  XNOR U21403 ( .A(y[6716]), .B(x[6716]), .Z(n13086) );
  XNOR U21404 ( .A(n13078), .B(n13079), .Z(n13089) );
  XNOR U21405 ( .A(y[6711]), .B(x[6711]), .Z(n13079) );
  XNOR U21406 ( .A(n13080), .B(n13081), .Z(n13078) );
  XNOR U21407 ( .A(y[6712]), .B(x[6712]), .Z(n13081) );
  XNOR U21408 ( .A(y[6713]), .B(x[6713]), .Z(n13080) );
  NAND U21409 ( .A(n13145), .B(n13146), .Z(N64223) );
  NANDN U21410 ( .A(n13147), .B(n13148), .Z(n13146) );
  OR U21411 ( .A(n13149), .B(n13150), .Z(n13148) );
  NAND U21412 ( .A(n13149), .B(n13150), .Z(n13145) );
  XOR U21413 ( .A(n13149), .B(n13151), .Z(N64222) );
  XNOR U21414 ( .A(n13147), .B(n13150), .Z(n13151) );
  AND U21415 ( .A(n13152), .B(n13153), .Z(n13150) );
  NANDN U21416 ( .A(n13154), .B(n13155), .Z(n13153) );
  NANDN U21417 ( .A(n13156), .B(n13157), .Z(n13155) );
  NANDN U21418 ( .A(n13157), .B(n13156), .Z(n13152) );
  NAND U21419 ( .A(n13158), .B(n13159), .Z(n13147) );
  NANDN U21420 ( .A(n13160), .B(n13161), .Z(n13159) );
  OR U21421 ( .A(n13162), .B(n13163), .Z(n13161) );
  NAND U21422 ( .A(n13163), .B(n13162), .Z(n13158) );
  AND U21423 ( .A(n13164), .B(n13165), .Z(n13149) );
  NANDN U21424 ( .A(n13166), .B(n13167), .Z(n13165) );
  NANDN U21425 ( .A(n13168), .B(n13169), .Z(n13167) );
  NANDN U21426 ( .A(n13169), .B(n13168), .Z(n13164) );
  XOR U21427 ( .A(n13163), .B(n13170), .Z(N64221) );
  XOR U21428 ( .A(n13160), .B(n13162), .Z(n13170) );
  XNOR U21429 ( .A(n13156), .B(n13171), .Z(n13162) );
  XNOR U21430 ( .A(n13154), .B(n13157), .Z(n13171) );
  NAND U21431 ( .A(n13172), .B(n13173), .Z(n13157) );
  NAND U21432 ( .A(n13174), .B(n13175), .Z(n13173) );
  OR U21433 ( .A(n13176), .B(n13177), .Z(n13174) );
  NANDN U21434 ( .A(n13178), .B(n13176), .Z(n13172) );
  IV U21435 ( .A(n13177), .Z(n13178) );
  NAND U21436 ( .A(n13179), .B(n13180), .Z(n13154) );
  NAND U21437 ( .A(n13181), .B(n13182), .Z(n13180) );
  NANDN U21438 ( .A(n13183), .B(n13184), .Z(n13181) );
  NANDN U21439 ( .A(n13184), .B(n13183), .Z(n13179) );
  AND U21440 ( .A(n13185), .B(n13186), .Z(n13156) );
  NAND U21441 ( .A(n13187), .B(n13188), .Z(n13186) );
  OR U21442 ( .A(n13189), .B(n13190), .Z(n13187) );
  NANDN U21443 ( .A(n13191), .B(n13189), .Z(n13185) );
  NAND U21444 ( .A(n13192), .B(n13193), .Z(n13160) );
  NANDN U21445 ( .A(n13194), .B(n13195), .Z(n13193) );
  OR U21446 ( .A(n13196), .B(n13197), .Z(n13195) );
  NANDN U21447 ( .A(n13198), .B(n13196), .Z(n13192) );
  IV U21448 ( .A(n13197), .Z(n13198) );
  XNOR U21449 ( .A(n13168), .B(n13199), .Z(n13163) );
  XNOR U21450 ( .A(n13166), .B(n13169), .Z(n13199) );
  NAND U21451 ( .A(n13200), .B(n13201), .Z(n13169) );
  NAND U21452 ( .A(n13202), .B(n13203), .Z(n13201) );
  OR U21453 ( .A(n13204), .B(n13205), .Z(n13202) );
  NANDN U21454 ( .A(n13206), .B(n13204), .Z(n13200) );
  IV U21455 ( .A(n13205), .Z(n13206) );
  NAND U21456 ( .A(n13207), .B(n13208), .Z(n13166) );
  NAND U21457 ( .A(n13209), .B(n13210), .Z(n13208) );
  NANDN U21458 ( .A(n13211), .B(n13212), .Z(n13209) );
  NANDN U21459 ( .A(n13212), .B(n13211), .Z(n13207) );
  AND U21460 ( .A(n13213), .B(n13214), .Z(n13168) );
  NAND U21461 ( .A(n13215), .B(n13216), .Z(n13214) );
  OR U21462 ( .A(n13217), .B(n13218), .Z(n13215) );
  NANDN U21463 ( .A(n13219), .B(n13217), .Z(n13213) );
  XNOR U21464 ( .A(n13194), .B(n13220), .Z(N64220) );
  XOR U21465 ( .A(n13196), .B(n13197), .Z(n13220) );
  XNOR U21466 ( .A(n13210), .B(n13221), .Z(n13197) );
  XOR U21467 ( .A(n13211), .B(n13212), .Z(n13221) );
  XOR U21468 ( .A(n13217), .B(n13222), .Z(n13212) );
  XOR U21469 ( .A(n13216), .B(n13219), .Z(n13222) );
  IV U21470 ( .A(n13218), .Z(n13219) );
  NAND U21471 ( .A(n13223), .B(n13224), .Z(n13218) );
  OR U21472 ( .A(n13225), .B(n13226), .Z(n13224) );
  OR U21473 ( .A(n13227), .B(n13228), .Z(n13223) );
  NAND U21474 ( .A(n13229), .B(n13230), .Z(n13216) );
  OR U21475 ( .A(n13231), .B(n13232), .Z(n13230) );
  OR U21476 ( .A(n13233), .B(n13234), .Z(n13229) );
  NOR U21477 ( .A(n13235), .B(n13236), .Z(n13217) );
  ANDN U21478 ( .B(n13237), .A(n13238), .Z(n13211) );
  XNOR U21479 ( .A(n13204), .B(n13239), .Z(n13210) );
  XNOR U21480 ( .A(n13203), .B(n13205), .Z(n13239) );
  NAND U21481 ( .A(n13240), .B(n13241), .Z(n13205) );
  OR U21482 ( .A(n13242), .B(n13243), .Z(n13241) );
  OR U21483 ( .A(n13244), .B(n13245), .Z(n13240) );
  NAND U21484 ( .A(n13246), .B(n13247), .Z(n13203) );
  OR U21485 ( .A(n13248), .B(n13249), .Z(n13247) );
  OR U21486 ( .A(n13250), .B(n13251), .Z(n13246) );
  ANDN U21487 ( .B(n13252), .A(n13253), .Z(n13204) );
  IV U21488 ( .A(n13254), .Z(n13252) );
  ANDN U21489 ( .B(n13255), .A(n13256), .Z(n13196) );
  XOR U21490 ( .A(n13182), .B(n13257), .Z(n13194) );
  XOR U21491 ( .A(n13183), .B(n13184), .Z(n13257) );
  XOR U21492 ( .A(n13189), .B(n13258), .Z(n13184) );
  XOR U21493 ( .A(n13188), .B(n13191), .Z(n13258) );
  IV U21494 ( .A(n13190), .Z(n13191) );
  NAND U21495 ( .A(n13259), .B(n13260), .Z(n13190) );
  OR U21496 ( .A(n13261), .B(n13262), .Z(n13260) );
  OR U21497 ( .A(n13263), .B(n13264), .Z(n13259) );
  NAND U21498 ( .A(n13265), .B(n13266), .Z(n13188) );
  OR U21499 ( .A(n13267), .B(n13268), .Z(n13266) );
  OR U21500 ( .A(n13269), .B(n13270), .Z(n13265) );
  NOR U21501 ( .A(n13271), .B(n13272), .Z(n13189) );
  ANDN U21502 ( .B(n13273), .A(n13274), .Z(n13183) );
  IV U21503 ( .A(n13275), .Z(n13273) );
  XNOR U21504 ( .A(n13176), .B(n13276), .Z(n13182) );
  XNOR U21505 ( .A(n13175), .B(n13177), .Z(n13276) );
  NAND U21506 ( .A(n13277), .B(n13278), .Z(n13177) );
  OR U21507 ( .A(n13279), .B(n13280), .Z(n13278) );
  OR U21508 ( .A(n13281), .B(n13282), .Z(n13277) );
  NAND U21509 ( .A(n13283), .B(n13284), .Z(n13175) );
  OR U21510 ( .A(n13285), .B(n13286), .Z(n13284) );
  OR U21511 ( .A(n13287), .B(n13288), .Z(n13283) );
  ANDN U21512 ( .B(n13289), .A(n13290), .Z(n13176) );
  IV U21513 ( .A(n13291), .Z(n13289) );
  XNOR U21514 ( .A(n13256), .B(n13255), .Z(N64219) );
  XOR U21515 ( .A(n13275), .B(n13274), .Z(n13255) );
  XNOR U21516 ( .A(n13290), .B(n13291), .Z(n13274) );
  XNOR U21517 ( .A(n13285), .B(n13286), .Z(n13291) );
  XNOR U21518 ( .A(n13287), .B(n13288), .Z(n13286) );
  XNOR U21519 ( .A(y[6709]), .B(x[6709]), .Z(n13288) );
  XNOR U21520 ( .A(y[6710]), .B(x[6710]), .Z(n13287) );
  XNOR U21521 ( .A(y[6708]), .B(x[6708]), .Z(n13285) );
  XNOR U21522 ( .A(n13279), .B(n13280), .Z(n13290) );
  XNOR U21523 ( .A(y[6705]), .B(x[6705]), .Z(n13280) );
  XNOR U21524 ( .A(n13281), .B(n13282), .Z(n13279) );
  XNOR U21525 ( .A(y[6706]), .B(x[6706]), .Z(n13282) );
  XNOR U21526 ( .A(y[6707]), .B(x[6707]), .Z(n13281) );
  XNOR U21527 ( .A(n13272), .B(n13271), .Z(n13275) );
  XNOR U21528 ( .A(n13267), .B(n13268), .Z(n13271) );
  XNOR U21529 ( .A(y[6702]), .B(x[6702]), .Z(n13268) );
  XNOR U21530 ( .A(n13269), .B(n13270), .Z(n13267) );
  XNOR U21531 ( .A(y[6703]), .B(x[6703]), .Z(n13270) );
  XNOR U21532 ( .A(y[6704]), .B(x[6704]), .Z(n13269) );
  XNOR U21533 ( .A(n13261), .B(n13262), .Z(n13272) );
  XNOR U21534 ( .A(y[6699]), .B(x[6699]), .Z(n13262) );
  XNOR U21535 ( .A(n13263), .B(n13264), .Z(n13261) );
  XNOR U21536 ( .A(y[6700]), .B(x[6700]), .Z(n13264) );
  XNOR U21537 ( .A(y[6701]), .B(x[6701]), .Z(n13263) );
  XOR U21538 ( .A(n13237), .B(n13238), .Z(n13256) );
  XNOR U21539 ( .A(n13253), .B(n13254), .Z(n13238) );
  XNOR U21540 ( .A(n13248), .B(n13249), .Z(n13254) );
  XNOR U21541 ( .A(n13250), .B(n13251), .Z(n13249) );
  XNOR U21542 ( .A(y[6697]), .B(x[6697]), .Z(n13251) );
  XNOR U21543 ( .A(y[6698]), .B(x[6698]), .Z(n13250) );
  XNOR U21544 ( .A(y[6696]), .B(x[6696]), .Z(n13248) );
  XNOR U21545 ( .A(n13242), .B(n13243), .Z(n13253) );
  XNOR U21546 ( .A(y[6693]), .B(x[6693]), .Z(n13243) );
  XNOR U21547 ( .A(n13244), .B(n13245), .Z(n13242) );
  XNOR U21548 ( .A(y[6694]), .B(x[6694]), .Z(n13245) );
  XNOR U21549 ( .A(y[6695]), .B(x[6695]), .Z(n13244) );
  XOR U21550 ( .A(n13236), .B(n13235), .Z(n13237) );
  XNOR U21551 ( .A(n13231), .B(n13232), .Z(n13235) );
  XNOR U21552 ( .A(y[6690]), .B(x[6690]), .Z(n13232) );
  XNOR U21553 ( .A(n13233), .B(n13234), .Z(n13231) );
  XNOR U21554 ( .A(y[6691]), .B(x[6691]), .Z(n13234) );
  XNOR U21555 ( .A(y[6692]), .B(x[6692]), .Z(n13233) );
  XNOR U21556 ( .A(n13225), .B(n13226), .Z(n13236) );
  XNOR U21557 ( .A(y[6687]), .B(x[6687]), .Z(n13226) );
  XNOR U21558 ( .A(n13227), .B(n13228), .Z(n13225) );
  XNOR U21559 ( .A(y[6688]), .B(x[6688]), .Z(n13228) );
  XNOR U21560 ( .A(y[6689]), .B(x[6689]), .Z(n13227) );
  NAND U21561 ( .A(n13292), .B(n13293), .Z(N64210) );
  NANDN U21562 ( .A(n13294), .B(n13295), .Z(n13293) );
  OR U21563 ( .A(n13296), .B(n13297), .Z(n13295) );
  NAND U21564 ( .A(n13296), .B(n13297), .Z(n13292) );
  XOR U21565 ( .A(n13296), .B(n13298), .Z(N64209) );
  XNOR U21566 ( .A(n13294), .B(n13297), .Z(n13298) );
  AND U21567 ( .A(n13299), .B(n13300), .Z(n13297) );
  NANDN U21568 ( .A(n13301), .B(n13302), .Z(n13300) );
  NANDN U21569 ( .A(n13303), .B(n13304), .Z(n13302) );
  NANDN U21570 ( .A(n13304), .B(n13303), .Z(n13299) );
  NAND U21571 ( .A(n13305), .B(n13306), .Z(n13294) );
  NANDN U21572 ( .A(n13307), .B(n13308), .Z(n13306) );
  OR U21573 ( .A(n13309), .B(n13310), .Z(n13308) );
  NAND U21574 ( .A(n13310), .B(n13309), .Z(n13305) );
  AND U21575 ( .A(n13311), .B(n13312), .Z(n13296) );
  NANDN U21576 ( .A(n13313), .B(n13314), .Z(n13312) );
  NANDN U21577 ( .A(n13315), .B(n13316), .Z(n13314) );
  NANDN U21578 ( .A(n13316), .B(n13315), .Z(n13311) );
  XOR U21579 ( .A(n13310), .B(n13317), .Z(N64208) );
  XOR U21580 ( .A(n13307), .B(n13309), .Z(n13317) );
  XNOR U21581 ( .A(n13303), .B(n13318), .Z(n13309) );
  XNOR U21582 ( .A(n13301), .B(n13304), .Z(n13318) );
  NAND U21583 ( .A(n13319), .B(n13320), .Z(n13304) );
  NAND U21584 ( .A(n13321), .B(n13322), .Z(n13320) );
  OR U21585 ( .A(n13323), .B(n13324), .Z(n13321) );
  NANDN U21586 ( .A(n13325), .B(n13323), .Z(n13319) );
  IV U21587 ( .A(n13324), .Z(n13325) );
  NAND U21588 ( .A(n13326), .B(n13327), .Z(n13301) );
  NAND U21589 ( .A(n13328), .B(n13329), .Z(n13327) );
  NANDN U21590 ( .A(n13330), .B(n13331), .Z(n13328) );
  NANDN U21591 ( .A(n13331), .B(n13330), .Z(n13326) );
  AND U21592 ( .A(n13332), .B(n13333), .Z(n13303) );
  NAND U21593 ( .A(n13334), .B(n13335), .Z(n13333) );
  OR U21594 ( .A(n13336), .B(n13337), .Z(n13334) );
  NANDN U21595 ( .A(n13338), .B(n13336), .Z(n13332) );
  NAND U21596 ( .A(n13339), .B(n13340), .Z(n13307) );
  NANDN U21597 ( .A(n13341), .B(n13342), .Z(n13340) );
  OR U21598 ( .A(n13343), .B(n13344), .Z(n13342) );
  NANDN U21599 ( .A(n13345), .B(n13343), .Z(n13339) );
  IV U21600 ( .A(n13344), .Z(n13345) );
  XNOR U21601 ( .A(n13315), .B(n13346), .Z(n13310) );
  XNOR U21602 ( .A(n13313), .B(n13316), .Z(n13346) );
  NAND U21603 ( .A(n13347), .B(n13348), .Z(n13316) );
  NAND U21604 ( .A(n13349), .B(n13350), .Z(n13348) );
  OR U21605 ( .A(n13351), .B(n13352), .Z(n13349) );
  NANDN U21606 ( .A(n13353), .B(n13351), .Z(n13347) );
  IV U21607 ( .A(n13352), .Z(n13353) );
  NAND U21608 ( .A(n13354), .B(n13355), .Z(n13313) );
  NAND U21609 ( .A(n13356), .B(n13357), .Z(n13355) );
  NANDN U21610 ( .A(n13358), .B(n13359), .Z(n13356) );
  NANDN U21611 ( .A(n13359), .B(n13358), .Z(n13354) );
  AND U21612 ( .A(n13360), .B(n13361), .Z(n13315) );
  NAND U21613 ( .A(n13362), .B(n13363), .Z(n13361) );
  OR U21614 ( .A(n13364), .B(n13365), .Z(n13362) );
  NANDN U21615 ( .A(n13366), .B(n13364), .Z(n13360) );
  XNOR U21616 ( .A(n13341), .B(n13367), .Z(N64207) );
  XOR U21617 ( .A(n13343), .B(n13344), .Z(n13367) );
  XNOR U21618 ( .A(n13357), .B(n13368), .Z(n13344) );
  XOR U21619 ( .A(n13358), .B(n13359), .Z(n13368) );
  XOR U21620 ( .A(n13364), .B(n13369), .Z(n13359) );
  XOR U21621 ( .A(n13363), .B(n13366), .Z(n13369) );
  IV U21622 ( .A(n13365), .Z(n13366) );
  NAND U21623 ( .A(n13370), .B(n13371), .Z(n13365) );
  OR U21624 ( .A(n13372), .B(n13373), .Z(n13371) );
  OR U21625 ( .A(n13374), .B(n13375), .Z(n13370) );
  NAND U21626 ( .A(n13376), .B(n13377), .Z(n13363) );
  OR U21627 ( .A(n13378), .B(n13379), .Z(n13377) );
  OR U21628 ( .A(n13380), .B(n13381), .Z(n13376) );
  NOR U21629 ( .A(n13382), .B(n13383), .Z(n13364) );
  ANDN U21630 ( .B(n13384), .A(n13385), .Z(n13358) );
  XNOR U21631 ( .A(n13351), .B(n13386), .Z(n13357) );
  XNOR U21632 ( .A(n13350), .B(n13352), .Z(n13386) );
  NAND U21633 ( .A(n13387), .B(n13388), .Z(n13352) );
  OR U21634 ( .A(n13389), .B(n13390), .Z(n13388) );
  OR U21635 ( .A(n13391), .B(n13392), .Z(n13387) );
  NAND U21636 ( .A(n13393), .B(n13394), .Z(n13350) );
  OR U21637 ( .A(n13395), .B(n13396), .Z(n13394) );
  OR U21638 ( .A(n13397), .B(n13398), .Z(n13393) );
  ANDN U21639 ( .B(n13399), .A(n13400), .Z(n13351) );
  IV U21640 ( .A(n13401), .Z(n13399) );
  ANDN U21641 ( .B(n13402), .A(n13403), .Z(n13343) );
  XOR U21642 ( .A(n13329), .B(n13404), .Z(n13341) );
  XOR U21643 ( .A(n13330), .B(n13331), .Z(n13404) );
  XOR U21644 ( .A(n13336), .B(n13405), .Z(n13331) );
  XOR U21645 ( .A(n13335), .B(n13338), .Z(n13405) );
  IV U21646 ( .A(n13337), .Z(n13338) );
  NAND U21647 ( .A(n13406), .B(n13407), .Z(n13337) );
  OR U21648 ( .A(n13408), .B(n13409), .Z(n13407) );
  OR U21649 ( .A(n13410), .B(n13411), .Z(n13406) );
  NAND U21650 ( .A(n13412), .B(n13413), .Z(n13335) );
  OR U21651 ( .A(n13414), .B(n13415), .Z(n13413) );
  OR U21652 ( .A(n13416), .B(n13417), .Z(n13412) );
  NOR U21653 ( .A(n13418), .B(n13419), .Z(n13336) );
  ANDN U21654 ( .B(n13420), .A(n13421), .Z(n13330) );
  IV U21655 ( .A(n13422), .Z(n13420) );
  XNOR U21656 ( .A(n13323), .B(n13423), .Z(n13329) );
  XNOR U21657 ( .A(n13322), .B(n13324), .Z(n13423) );
  NAND U21658 ( .A(n13424), .B(n13425), .Z(n13324) );
  OR U21659 ( .A(n13426), .B(n13427), .Z(n13425) );
  OR U21660 ( .A(n13428), .B(n13429), .Z(n13424) );
  NAND U21661 ( .A(n13430), .B(n13431), .Z(n13322) );
  OR U21662 ( .A(n13432), .B(n13433), .Z(n13431) );
  OR U21663 ( .A(n13434), .B(n13435), .Z(n13430) );
  ANDN U21664 ( .B(n13436), .A(n13437), .Z(n13323) );
  IV U21665 ( .A(n13438), .Z(n13436) );
  XNOR U21666 ( .A(n13403), .B(n13402), .Z(N64206) );
  XOR U21667 ( .A(n13422), .B(n13421), .Z(n13402) );
  XNOR U21668 ( .A(n13437), .B(n13438), .Z(n13421) );
  XNOR U21669 ( .A(n13432), .B(n13433), .Z(n13438) );
  XNOR U21670 ( .A(n13434), .B(n13435), .Z(n13433) );
  XNOR U21671 ( .A(y[6685]), .B(x[6685]), .Z(n13435) );
  XNOR U21672 ( .A(y[6686]), .B(x[6686]), .Z(n13434) );
  XNOR U21673 ( .A(y[6684]), .B(x[6684]), .Z(n13432) );
  XNOR U21674 ( .A(n13426), .B(n13427), .Z(n13437) );
  XNOR U21675 ( .A(y[6681]), .B(x[6681]), .Z(n13427) );
  XNOR U21676 ( .A(n13428), .B(n13429), .Z(n13426) );
  XNOR U21677 ( .A(y[6682]), .B(x[6682]), .Z(n13429) );
  XNOR U21678 ( .A(y[6683]), .B(x[6683]), .Z(n13428) );
  XNOR U21679 ( .A(n13419), .B(n13418), .Z(n13422) );
  XNOR U21680 ( .A(n13414), .B(n13415), .Z(n13418) );
  XNOR U21681 ( .A(y[6678]), .B(x[6678]), .Z(n13415) );
  XNOR U21682 ( .A(n13416), .B(n13417), .Z(n13414) );
  XNOR U21683 ( .A(y[6679]), .B(x[6679]), .Z(n13417) );
  XNOR U21684 ( .A(y[6680]), .B(x[6680]), .Z(n13416) );
  XNOR U21685 ( .A(n13408), .B(n13409), .Z(n13419) );
  XNOR U21686 ( .A(y[6675]), .B(x[6675]), .Z(n13409) );
  XNOR U21687 ( .A(n13410), .B(n13411), .Z(n13408) );
  XNOR U21688 ( .A(y[6676]), .B(x[6676]), .Z(n13411) );
  XNOR U21689 ( .A(y[6677]), .B(x[6677]), .Z(n13410) );
  XOR U21690 ( .A(n13384), .B(n13385), .Z(n13403) );
  XNOR U21691 ( .A(n13400), .B(n13401), .Z(n13385) );
  XNOR U21692 ( .A(n13395), .B(n13396), .Z(n13401) );
  XNOR U21693 ( .A(n13397), .B(n13398), .Z(n13396) );
  XNOR U21694 ( .A(y[6673]), .B(x[6673]), .Z(n13398) );
  XNOR U21695 ( .A(y[6674]), .B(x[6674]), .Z(n13397) );
  XNOR U21696 ( .A(y[6672]), .B(x[6672]), .Z(n13395) );
  XNOR U21697 ( .A(n13389), .B(n13390), .Z(n13400) );
  XNOR U21698 ( .A(y[6669]), .B(x[6669]), .Z(n13390) );
  XNOR U21699 ( .A(n13391), .B(n13392), .Z(n13389) );
  XNOR U21700 ( .A(y[6670]), .B(x[6670]), .Z(n13392) );
  XNOR U21701 ( .A(y[6671]), .B(x[6671]), .Z(n13391) );
  XOR U21702 ( .A(n13383), .B(n13382), .Z(n13384) );
  XNOR U21703 ( .A(n13378), .B(n13379), .Z(n13382) );
  XNOR U21704 ( .A(y[6666]), .B(x[6666]), .Z(n13379) );
  XNOR U21705 ( .A(n13380), .B(n13381), .Z(n13378) );
  XNOR U21706 ( .A(y[6667]), .B(x[6667]), .Z(n13381) );
  XNOR U21707 ( .A(y[6668]), .B(x[6668]), .Z(n13380) );
  XNOR U21708 ( .A(n13372), .B(n13373), .Z(n13383) );
  XNOR U21709 ( .A(y[6663]), .B(x[6663]), .Z(n13373) );
  XNOR U21710 ( .A(n13374), .B(n13375), .Z(n13372) );
  XNOR U21711 ( .A(y[6664]), .B(x[6664]), .Z(n13375) );
  XNOR U21712 ( .A(y[6665]), .B(x[6665]), .Z(n13374) );
  NAND U21713 ( .A(n13439), .B(n13440), .Z(N64197) );
  NANDN U21714 ( .A(n13441), .B(n13442), .Z(n13440) );
  OR U21715 ( .A(n13443), .B(n13444), .Z(n13442) );
  NAND U21716 ( .A(n13443), .B(n13444), .Z(n13439) );
  XOR U21717 ( .A(n13443), .B(n13445), .Z(N64196) );
  XNOR U21718 ( .A(n13441), .B(n13444), .Z(n13445) );
  AND U21719 ( .A(n13446), .B(n13447), .Z(n13444) );
  NANDN U21720 ( .A(n13448), .B(n13449), .Z(n13447) );
  NANDN U21721 ( .A(n13450), .B(n13451), .Z(n13449) );
  NANDN U21722 ( .A(n13451), .B(n13450), .Z(n13446) );
  NAND U21723 ( .A(n13452), .B(n13453), .Z(n13441) );
  NANDN U21724 ( .A(n13454), .B(n13455), .Z(n13453) );
  OR U21725 ( .A(n13456), .B(n13457), .Z(n13455) );
  NAND U21726 ( .A(n13457), .B(n13456), .Z(n13452) );
  AND U21727 ( .A(n13458), .B(n13459), .Z(n13443) );
  NANDN U21728 ( .A(n13460), .B(n13461), .Z(n13459) );
  NANDN U21729 ( .A(n13462), .B(n13463), .Z(n13461) );
  NANDN U21730 ( .A(n13463), .B(n13462), .Z(n13458) );
  XOR U21731 ( .A(n13457), .B(n13464), .Z(N64195) );
  XOR U21732 ( .A(n13454), .B(n13456), .Z(n13464) );
  XNOR U21733 ( .A(n13450), .B(n13465), .Z(n13456) );
  XNOR U21734 ( .A(n13448), .B(n13451), .Z(n13465) );
  NAND U21735 ( .A(n13466), .B(n13467), .Z(n13451) );
  NAND U21736 ( .A(n13468), .B(n13469), .Z(n13467) );
  OR U21737 ( .A(n13470), .B(n13471), .Z(n13468) );
  NANDN U21738 ( .A(n13472), .B(n13470), .Z(n13466) );
  IV U21739 ( .A(n13471), .Z(n13472) );
  NAND U21740 ( .A(n13473), .B(n13474), .Z(n13448) );
  NAND U21741 ( .A(n13475), .B(n13476), .Z(n13474) );
  NANDN U21742 ( .A(n13477), .B(n13478), .Z(n13475) );
  NANDN U21743 ( .A(n13478), .B(n13477), .Z(n13473) );
  AND U21744 ( .A(n13479), .B(n13480), .Z(n13450) );
  NAND U21745 ( .A(n13481), .B(n13482), .Z(n13480) );
  OR U21746 ( .A(n13483), .B(n13484), .Z(n13481) );
  NANDN U21747 ( .A(n13485), .B(n13483), .Z(n13479) );
  NAND U21748 ( .A(n13486), .B(n13487), .Z(n13454) );
  NANDN U21749 ( .A(n13488), .B(n13489), .Z(n13487) );
  OR U21750 ( .A(n13490), .B(n13491), .Z(n13489) );
  NANDN U21751 ( .A(n13492), .B(n13490), .Z(n13486) );
  IV U21752 ( .A(n13491), .Z(n13492) );
  XNOR U21753 ( .A(n13462), .B(n13493), .Z(n13457) );
  XNOR U21754 ( .A(n13460), .B(n13463), .Z(n13493) );
  NAND U21755 ( .A(n13494), .B(n13495), .Z(n13463) );
  NAND U21756 ( .A(n13496), .B(n13497), .Z(n13495) );
  OR U21757 ( .A(n13498), .B(n13499), .Z(n13496) );
  NANDN U21758 ( .A(n13500), .B(n13498), .Z(n13494) );
  IV U21759 ( .A(n13499), .Z(n13500) );
  NAND U21760 ( .A(n13501), .B(n13502), .Z(n13460) );
  NAND U21761 ( .A(n13503), .B(n13504), .Z(n13502) );
  NANDN U21762 ( .A(n13505), .B(n13506), .Z(n13503) );
  NANDN U21763 ( .A(n13506), .B(n13505), .Z(n13501) );
  AND U21764 ( .A(n13507), .B(n13508), .Z(n13462) );
  NAND U21765 ( .A(n13509), .B(n13510), .Z(n13508) );
  OR U21766 ( .A(n13511), .B(n13512), .Z(n13509) );
  NANDN U21767 ( .A(n13513), .B(n13511), .Z(n13507) );
  XNOR U21768 ( .A(n13488), .B(n13514), .Z(N64194) );
  XOR U21769 ( .A(n13490), .B(n13491), .Z(n13514) );
  XNOR U21770 ( .A(n13504), .B(n13515), .Z(n13491) );
  XOR U21771 ( .A(n13505), .B(n13506), .Z(n13515) );
  XOR U21772 ( .A(n13511), .B(n13516), .Z(n13506) );
  XOR U21773 ( .A(n13510), .B(n13513), .Z(n13516) );
  IV U21774 ( .A(n13512), .Z(n13513) );
  NAND U21775 ( .A(n13517), .B(n13518), .Z(n13512) );
  OR U21776 ( .A(n13519), .B(n13520), .Z(n13518) );
  OR U21777 ( .A(n13521), .B(n13522), .Z(n13517) );
  NAND U21778 ( .A(n13523), .B(n13524), .Z(n13510) );
  OR U21779 ( .A(n13525), .B(n13526), .Z(n13524) );
  OR U21780 ( .A(n13527), .B(n13528), .Z(n13523) );
  NOR U21781 ( .A(n13529), .B(n13530), .Z(n13511) );
  ANDN U21782 ( .B(n13531), .A(n13532), .Z(n13505) );
  XNOR U21783 ( .A(n13498), .B(n13533), .Z(n13504) );
  XNOR U21784 ( .A(n13497), .B(n13499), .Z(n13533) );
  NAND U21785 ( .A(n13534), .B(n13535), .Z(n13499) );
  OR U21786 ( .A(n13536), .B(n13537), .Z(n13535) );
  OR U21787 ( .A(n13538), .B(n13539), .Z(n13534) );
  NAND U21788 ( .A(n13540), .B(n13541), .Z(n13497) );
  OR U21789 ( .A(n13542), .B(n13543), .Z(n13541) );
  OR U21790 ( .A(n13544), .B(n13545), .Z(n13540) );
  ANDN U21791 ( .B(n13546), .A(n13547), .Z(n13498) );
  IV U21792 ( .A(n13548), .Z(n13546) );
  ANDN U21793 ( .B(n13549), .A(n13550), .Z(n13490) );
  XOR U21794 ( .A(n13476), .B(n13551), .Z(n13488) );
  XOR U21795 ( .A(n13477), .B(n13478), .Z(n13551) );
  XOR U21796 ( .A(n13483), .B(n13552), .Z(n13478) );
  XOR U21797 ( .A(n13482), .B(n13485), .Z(n13552) );
  IV U21798 ( .A(n13484), .Z(n13485) );
  NAND U21799 ( .A(n13553), .B(n13554), .Z(n13484) );
  OR U21800 ( .A(n13555), .B(n13556), .Z(n13554) );
  OR U21801 ( .A(n13557), .B(n13558), .Z(n13553) );
  NAND U21802 ( .A(n13559), .B(n13560), .Z(n13482) );
  OR U21803 ( .A(n13561), .B(n13562), .Z(n13560) );
  OR U21804 ( .A(n13563), .B(n13564), .Z(n13559) );
  NOR U21805 ( .A(n13565), .B(n13566), .Z(n13483) );
  ANDN U21806 ( .B(n13567), .A(n13568), .Z(n13477) );
  IV U21807 ( .A(n13569), .Z(n13567) );
  XNOR U21808 ( .A(n13470), .B(n13570), .Z(n13476) );
  XNOR U21809 ( .A(n13469), .B(n13471), .Z(n13570) );
  NAND U21810 ( .A(n13571), .B(n13572), .Z(n13471) );
  OR U21811 ( .A(n13573), .B(n13574), .Z(n13572) );
  OR U21812 ( .A(n13575), .B(n13576), .Z(n13571) );
  NAND U21813 ( .A(n13577), .B(n13578), .Z(n13469) );
  OR U21814 ( .A(n13579), .B(n13580), .Z(n13578) );
  OR U21815 ( .A(n13581), .B(n13582), .Z(n13577) );
  ANDN U21816 ( .B(n13583), .A(n13584), .Z(n13470) );
  IV U21817 ( .A(n13585), .Z(n13583) );
  XNOR U21818 ( .A(n13550), .B(n13549), .Z(N64193) );
  XOR U21819 ( .A(n13569), .B(n13568), .Z(n13549) );
  XNOR U21820 ( .A(n13584), .B(n13585), .Z(n13568) );
  XNOR U21821 ( .A(n13579), .B(n13580), .Z(n13585) );
  XNOR U21822 ( .A(n13581), .B(n13582), .Z(n13580) );
  XNOR U21823 ( .A(y[6661]), .B(x[6661]), .Z(n13582) );
  XNOR U21824 ( .A(y[6662]), .B(x[6662]), .Z(n13581) );
  XNOR U21825 ( .A(y[6660]), .B(x[6660]), .Z(n13579) );
  XNOR U21826 ( .A(n13573), .B(n13574), .Z(n13584) );
  XNOR U21827 ( .A(y[6657]), .B(x[6657]), .Z(n13574) );
  XNOR U21828 ( .A(n13575), .B(n13576), .Z(n13573) );
  XNOR U21829 ( .A(y[6658]), .B(x[6658]), .Z(n13576) );
  XNOR U21830 ( .A(y[6659]), .B(x[6659]), .Z(n13575) );
  XNOR U21831 ( .A(n13566), .B(n13565), .Z(n13569) );
  XNOR U21832 ( .A(n13561), .B(n13562), .Z(n13565) );
  XNOR U21833 ( .A(y[6654]), .B(x[6654]), .Z(n13562) );
  XNOR U21834 ( .A(n13563), .B(n13564), .Z(n13561) );
  XNOR U21835 ( .A(y[6655]), .B(x[6655]), .Z(n13564) );
  XNOR U21836 ( .A(y[6656]), .B(x[6656]), .Z(n13563) );
  XNOR U21837 ( .A(n13555), .B(n13556), .Z(n13566) );
  XNOR U21838 ( .A(y[6651]), .B(x[6651]), .Z(n13556) );
  XNOR U21839 ( .A(n13557), .B(n13558), .Z(n13555) );
  XNOR U21840 ( .A(y[6652]), .B(x[6652]), .Z(n13558) );
  XNOR U21841 ( .A(y[6653]), .B(x[6653]), .Z(n13557) );
  XOR U21842 ( .A(n13531), .B(n13532), .Z(n13550) );
  XNOR U21843 ( .A(n13547), .B(n13548), .Z(n13532) );
  XNOR U21844 ( .A(n13542), .B(n13543), .Z(n13548) );
  XNOR U21845 ( .A(n13544), .B(n13545), .Z(n13543) );
  XNOR U21846 ( .A(y[6649]), .B(x[6649]), .Z(n13545) );
  XNOR U21847 ( .A(y[6650]), .B(x[6650]), .Z(n13544) );
  XNOR U21848 ( .A(y[6648]), .B(x[6648]), .Z(n13542) );
  XNOR U21849 ( .A(n13536), .B(n13537), .Z(n13547) );
  XNOR U21850 ( .A(y[6645]), .B(x[6645]), .Z(n13537) );
  XNOR U21851 ( .A(n13538), .B(n13539), .Z(n13536) );
  XNOR U21852 ( .A(y[6646]), .B(x[6646]), .Z(n13539) );
  XNOR U21853 ( .A(y[6647]), .B(x[6647]), .Z(n13538) );
  XOR U21854 ( .A(n13530), .B(n13529), .Z(n13531) );
  XNOR U21855 ( .A(n13525), .B(n13526), .Z(n13529) );
  XNOR U21856 ( .A(y[6642]), .B(x[6642]), .Z(n13526) );
  XNOR U21857 ( .A(n13527), .B(n13528), .Z(n13525) );
  XNOR U21858 ( .A(y[6643]), .B(x[6643]), .Z(n13528) );
  XNOR U21859 ( .A(y[6644]), .B(x[6644]), .Z(n13527) );
  XNOR U21860 ( .A(n13519), .B(n13520), .Z(n13530) );
  XNOR U21861 ( .A(y[6639]), .B(x[6639]), .Z(n13520) );
  XNOR U21862 ( .A(n13521), .B(n13522), .Z(n13519) );
  XNOR U21863 ( .A(y[6640]), .B(x[6640]), .Z(n13522) );
  XNOR U21864 ( .A(y[6641]), .B(x[6641]), .Z(n13521) );
  NAND U21865 ( .A(n13586), .B(n13587), .Z(N64184) );
  NANDN U21866 ( .A(n13588), .B(n13589), .Z(n13587) );
  OR U21867 ( .A(n13590), .B(n13591), .Z(n13589) );
  NAND U21868 ( .A(n13590), .B(n13591), .Z(n13586) );
  XOR U21869 ( .A(n13590), .B(n13592), .Z(N64183) );
  XNOR U21870 ( .A(n13588), .B(n13591), .Z(n13592) );
  AND U21871 ( .A(n13593), .B(n13594), .Z(n13591) );
  NANDN U21872 ( .A(n13595), .B(n13596), .Z(n13594) );
  NANDN U21873 ( .A(n13597), .B(n13598), .Z(n13596) );
  NANDN U21874 ( .A(n13598), .B(n13597), .Z(n13593) );
  NAND U21875 ( .A(n13599), .B(n13600), .Z(n13588) );
  NANDN U21876 ( .A(n13601), .B(n13602), .Z(n13600) );
  OR U21877 ( .A(n13603), .B(n13604), .Z(n13602) );
  NAND U21878 ( .A(n13604), .B(n13603), .Z(n13599) );
  AND U21879 ( .A(n13605), .B(n13606), .Z(n13590) );
  NANDN U21880 ( .A(n13607), .B(n13608), .Z(n13606) );
  NANDN U21881 ( .A(n13609), .B(n13610), .Z(n13608) );
  NANDN U21882 ( .A(n13610), .B(n13609), .Z(n13605) );
  XOR U21883 ( .A(n13604), .B(n13611), .Z(N64182) );
  XOR U21884 ( .A(n13601), .B(n13603), .Z(n13611) );
  XNOR U21885 ( .A(n13597), .B(n13612), .Z(n13603) );
  XNOR U21886 ( .A(n13595), .B(n13598), .Z(n13612) );
  NAND U21887 ( .A(n13613), .B(n13614), .Z(n13598) );
  NAND U21888 ( .A(n13615), .B(n13616), .Z(n13614) );
  OR U21889 ( .A(n13617), .B(n13618), .Z(n13615) );
  NANDN U21890 ( .A(n13619), .B(n13617), .Z(n13613) );
  IV U21891 ( .A(n13618), .Z(n13619) );
  NAND U21892 ( .A(n13620), .B(n13621), .Z(n13595) );
  NAND U21893 ( .A(n13622), .B(n13623), .Z(n13621) );
  NANDN U21894 ( .A(n13624), .B(n13625), .Z(n13622) );
  NANDN U21895 ( .A(n13625), .B(n13624), .Z(n13620) );
  AND U21896 ( .A(n13626), .B(n13627), .Z(n13597) );
  NAND U21897 ( .A(n13628), .B(n13629), .Z(n13627) );
  OR U21898 ( .A(n13630), .B(n13631), .Z(n13628) );
  NANDN U21899 ( .A(n13632), .B(n13630), .Z(n13626) );
  NAND U21900 ( .A(n13633), .B(n13634), .Z(n13601) );
  NANDN U21901 ( .A(n13635), .B(n13636), .Z(n13634) );
  OR U21902 ( .A(n13637), .B(n13638), .Z(n13636) );
  NANDN U21903 ( .A(n13639), .B(n13637), .Z(n13633) );
  IV U21904 ( .A(n13638), .Z(n13639) );
  XNOR U21905 ( .A(n13609), .B(n13640), .Z(n13604) );
  XNOR U21906 ( .A(n13607), .B(n13610), .Z(n13640) );
  NAND U21907 ( .A(n13641), .B(n13642), .Z(n13610) );
  NAND U21908 ( .A(n13643), .B(n13644), .Z(n13642) );
  OR U21909 ( .A(n13645), .B(n13646), .Z(n13643) );
  NANDN U21910 ( .A(n13647), .B(n13645), .Z(n13641) );
  IV U21911 ( .A(n13646), .Z(n13647) );
  NAND U21912 ( .A(n13648), .B(n13649), .Z(n13607) );
  NAND U21913 ( .A(n13650), .B(n13651), .Z(n13649) );
  NANDN U21914 ( .A(n13652), .B(n13653), .Z(n13650) );
  NANDN U21915 ( .A(n13653), .B(n13652), .Z(n13648) );
  AND U21916 ( .A(n13654), .B(n13655), .Z(n13609) );
  NAND U21917 ( .A(n13656), .B(n13657), .Z(n13655) );
  OR U21918 ( .A(n13658), .B(n13659), .Z(n13656) );
  NANDN U21919 ( .A(n13660), .B(n13658), .Z(n13654) );
  XNOR U21920 ( .A(n13635), .B(n13661), .Z(N64181) );
  XOR U21921 ( .A(n13637), .B(n13638), .Z(n13661) );
  XNOR U21922 ( .A(n13651), .B(n13662), .Z(n13638) );
  XOR U21923 ( .A(n13652), .B(n13653), .Z(n13662) );
  XOR U21924 ( .A(n13658), .B(n13663), .Z(n13653) );
  XOR U21925 ( .A(n13657), .B(n13660), .Z(n13663) );
  IV U21926 ( .A(n13659), .Z(n13660) );
  NAND U21927 ( .A(n13664), .B(n13665), .Z(n13659) );
  OR U21928 ( .A(n13666), .B(n13667), .Z(n13665) );
  OR U21929 ( .A(n13668), .B(n13669), .Z(n13664) );
  NAND U21930 ( .A(n13670), .B(n13671), .Z(n13657) );
  OR U21931 ( .A(n13672), .B(n13673), .Z(n13671) );
  OR U21932 ( .A(n13674), .B(n13675), .Z(n13670) );
  NOR U21933 ( .A(n13676), .B(n13677), .Z(n13658) );
  ANDN U21934 ( .B(n13678), .A(n13679), .Z(n13652) );
  XNOR U21935 ( .A(n13645), .B(n13680), .Z(n13651) );
  XNOR U21936 ( .A(n13644), .B(n13646), .Z(n13680) );
  NAND U21937 ( .A(n13681), .B(n13682), .Z(n13646) );
  OR U21938 ( .A(n13683), .B(n13684), .Z(n13682) );
  OR U21939 ( .A(n13685), .B(n13686), .Z(n13681) );
  NAND U21940 ( .A(n13687), .B(n13688), .Z(n13644) );
  OR U21941 ( .A(n13689), .B(n13690), .Z(n13688) );
  OR U21942 ( .A(n13691), .B(n13692), .Z(n13687) );
  ANDN U21943 ( .B(n13693), .A(n13694), .Z(n13645) );
  IV U21944 ( .A(n13695), .Z(n13693) );
  ANDN U21945 ( .B(n13696), .A(n13697), .Z(n13637) );
  XOR U21946 ( .A(n13623), .B(n13698), .Z(n13635) );
  XOR U21947 ( .A(n13624), .B(n13625), .Z(n13698) );
  XOR U21948 ( .A(n13630), .B(n13699), .Z(n13625) );
  XOR U21949 ( .A(n13629), .B(n13632), .Z(n13699) );
  IV U21950 ( .A(n13631), .Z(n13632) );
  NAND U21951 ( .A(n13700), .B(n13701), .Z(n13631) );
  OR U21952 ( .A(n13702), .B(n13703), .Z(n13701) );
  OR U21953 ( .A(n13704), .B(n13705), .Z(n13700) );
  NAND U21954 ( .A(n13706), .B(n13707), .Z(n13629) );
  OR U21955 ( .A(n13708), .B(n13709), .Z(n13707) );
  OR U21956 ( .A(n13710), .B(n13711), .Z(n13706) );
  NOR U21957 ( .A(n13712), .B(n13713), .Z(n13630) );
  ANDN U21958 ( .B(n13714), .A(n13715), .Z(n13624) );
  IV U21959 ( .A(n13716), .Z(n13714) );
  XNOR U21960 ( .A(n13617), .B(n13717), .Z(n13623) );
  XNOR U21961 ( .A(n13616), .B(n13618), .Z(n13717) );
  NAND U21962 ( .A(n13718), .B(n13719), .Z(n13618) );
  OR U21963 ( .A(n13720), .B(n13721), .Z(n13719) );
  OR U21964 ( .A(n13722), .B(n13723), .Z(n13718) );
  NAND U21965 ( .A(n13724), .B(n13725), .Z(n13616) );
  OR U21966 ( .A(n13726), .B(n13727), .Z(n13725) );
  OR U21967 ( .A(n13728), .B(n13729), .Z(n13724) );
  ANDN U21968 ( .B(n13730), .A(n13731), .Z(n13617) );
  IV U21969 ( .A(n13732), .Z(n13730) );
  XNOR U21970 ( .A(n13697), .B(n13696), .Z(N64180) );
  XOR U21971 ( .A(n13716), .B(n13715), .Z(n13696) );
  XNOR U21972 ( .A(n13731), .B(n13732), .Z(n13715) );
  XNOR U21973 ( .A(n13726), .B(n13727), .Z(n13732) );
  XNOR U21974 ( .A(n13728), .B(n13729), .Z(n13727) );
  XNOR U21975 ( .A(y[6637]), .B(x[6637]), .Z(n13729) );
  XNOR U21976 ( .A(y[6638]), .B(x[6638]), .Z(n13728) );
  XNOR U21977 ( .A(y[6636]), .B(x[6636]), .Z(n13726) );
  XNOR U21978 ( .A(n13720), .B(n13721), .Z(n13731) );
  XNOR U21979 ( .A(y[6633]), .B(x[6633]), .Z(n13721) );
  XNOR U21980 ( .A(n13722), .B(n13723), .Z(n13720) );
  XNOR U21981 ( .A(y[6634]), .B(x[6634]), .Z(n13723) );
  XNOR U21982 ( .A(y[6635]), .B(x[6635]), .Z(n13722) );
  XNOR U21983 ( .A(n13713), .B(n13712), .Z(n13716) );
  XNOR U21984 ( .A(n13708), .B(n13709), .Z(n13712) );
  XNOR U21985 ( .A(y[6630]), .B(x[6630]), .Z(n13709) );
  XNOR U21986 ( .A(n13710), .B(n13711), .Z(n13708) );
  XNOR U21987 ( .A(y[6631]), .B(x[6631]), .Z(n13711) );
  XNOR U21988 ( .A(y[6632]), .B(x[6632]), .Z(n13710) );
  XNOR U21989 ( .A(n13702), .B(n13703), .Z(n13713) );
  XNOR U21990 ( .A(y[6627]), .B(x[6627]), .Z(n13703) );
  XNOR U21991 ( .A(n13704), .B(n13705), .Z(n13702) );
  XNOR U21992 ( .A(y[6628]), .B(x[6628]), .Z(n13705) );
  XNOR U21993 ( .A(y[6629]), .B(x[6629]), .Z(n13704) );
  XOR U21994 ( .A(n13678), .B(n13679), .Z(n13697) );
  XNOR U21995 ( .A(n13694), .B(n13695), .Z(n13679) );
  XNOR U21996 ( .A(n13689), .B(n13690), .Z(n13695) );
  XNOR U21997 ( .A(n13691), .B(n13692), .Z(n13690) );
  XNOR U21998 ( .A(y[6625]), .B(x[6625]), .Z(n13692) );
  XNOR U21999 ( .A(y[6626]), .B(x[6626]), .Z(n13691) );
  XNOR U22000 ( .A(y[6624]), .B(x[6624]), .Z(n13689) );
  XNOR U22001 ( .A(n13683), .B(n13684), .Z(n13694) );
  XNOR U22002 ( .A(y[6621]), .B(x[6621]), .Z(n13684) );
  XNOR U22003 ( .A(n13685), .B(n13686), .Z(n13683) );
  XNOR U22004 ( .A(y[6622]), .B(x[6622]), .Z(n13686) );
  XNOR U22005 ( .A(y[6623]), .B(x[6623]), .Z(n13685) );
  XOR U22006 ( .A(n13677), .B(n13676), .Z(n13678) );
  XNOR U22007 ( .A(n13672), .B(n13673), .Z(n13676) );
  XNOR U22008 ( .A(y[6618]), .B(x[6618]), .Z(n13673) );
  XNOR U22009 ( .A(n13674), .B(n13675), .Z(n13672) );
  XNOR U22010 ( .A(y[6619]), .B(x[6619]), .Z(n13675) );
  XNOR U22011 ( .A(y[6620]), .B(x[6620]), .Z(n13674) );
  XNOR U22012 ( .A(n13666), .B(n13667), .Z(n13677) );
  XNOR U22013 ( .A(y[6615]), .B(x[6615]), .Z(n13667) );
  XNOR U22014 ( .A(n13668), .B(n13669), .Z(n13666) );
  XNOR U22015 ( .A(y[6616]), .B(x[6616]), .Z(n13669) );
  XNOR U22016 ( .A(y[6617]), .B(x[6617]), .Z(n13668) );
  NAND U22017 ( .A(n13733), .B(n13734), .Z(N64171) );
  NANDN U22018 ( .A(n13735), .B(n13736), .Z(n13734) );
  OR U22019 ( .A(n13737), .B(n13738), .Z(n13736) );
  NAND U22020 ( .A(n13737), .B(n13738), .Z(n13733) );
  XOR U22021 ( .A(n13737), .B(n13739), .Z(N64170) );
  XNOR U22022 ( .A(n13735), .B(n13738), .Z(n13739) );
  AND U22023 ( .A(n13740), .B(n13741), .Z(n13738) );
  NANDN U22024 ( .A(n13742), .B(n13743), .Z(n13741) );
  NANDN U22025 ( .A(n13744), .B(n13745), .Z(n13743) );
  NANDN U22026 ( .A(n13745), .B(n13744), .Z(n13740) );
  NAND U22027 ( .A(n13746), .B(n13747), .Z(n13735) );
  NANDN U22028 ( .A(n13748), .B(n13749), .Z(n13747) );
  OR U22029 ( .A(n13750), .B(n13751), .Z(n13749) );
  NAND U22030 ( .A(n13751), .B(n13750), .Z(n13746) );
  AND U22031 ( .A(n13752), .B(n13753), .Z(n13737) );
  NANDN U22032 ( .A(n13754), .B(n13755), .Z(n13753) );
  NANDN U22033 ( .A(n13756), .B(n13757), .Z(n13755) );
  NANDN U22034 ( .A(n13757), .B(n13756), .Z(n13752) );
  XOR U22035 ( .A(n13751), .B(n13758), .Z(N64169) );
  XOR U22036 ( .A(n13748), .B(n13750), .Z(n13758) );
  XNOR U22037 ( .A(n13744), .B(n13759), .Z(n13750) );
  XNOR U22038 ( .A(n13742), .B(n13745), .Z(n13759) );
  NAND U22039 ( .A(n13760), .B(n13761), .Z(n13745) );
  NAND U22040 ( .A(n13762), .B(n13763), .Z(n13761) );
  OR U22041 ( .A(n13764), .B(n13765), .Z(n13762) );
  NANDN U22042 ( .A(n13766), .B(n13764), .Z(n13760) );
  IV U22043 ( .A(n13765), .Z(n13766) );
  NAND U22044 ( .A(n13767), .B(n13768), .Z(n13742) );
  NAND U22045 ( .A(n13769), .B(n13770), .Z(n13768) );
  NANDN U22046 ( .A(n13771), .B(n13772), .Z(n13769) );
  NANDN U22047 ( .A(n13772), .B(n13771), .Z(n13767) );
  AND U22048 ( .A(n13773), .B(n13774), .Z(n13744) );
  NAND U22049 ( .A(n13775), .B(n13776), .Z(n13774) );
  OR U22050 ( .A(n13777), .B(n13778), .Z(n13775) );
  NANDN U22051 ( .A(n13779), .B(n13777), .Z(n13773) );
  NAND U22052 ( .A(n13780), .B(n13781), .Z(n13748) );
  NANDN U22053 ( .A(n13782), .B(n13783), .Z(n13781) );
  OR U22054 ( .A(n13784), .B(n13785), .Z(n13783) );
  NANDN U22055 ( .A(n13786), .B(n13784), .Z(n13780) );
  IV U22056 ( .A(n13785), .Z(n13786) );
  XNOR U22057 ( .A(n13756), .B(n13787), .Z(n13751) );
  XNOR U22058 ( .A(n13754), .B(n13757), .Z(n13787) );
  NAND U22059 ( .A(n13788), .B(n13789), .Z(n13757) );
  NAND U22060 ( .A(n13790), .B(n13791), .Z(n13789) );
  OR U22061 ( .A(n13792), .B(n13793), .Z(n13790) );
  NANDN U22062 ( .A(n13794), .B(n13792), .Z(n13788) );
  IV U22063 ( .A(n13793), .Z(n13794) );
  NAND U22064 ( .A(n13795), .B(n13796), .Z(n13754) );
  NAND U22065 ( .A(n13797), .B(n13798), .Z(n13796) );
  NANDN U22066 ( .A(n13799), .B(n13800), .Z(n13797) );
  NANDN U22067 ( .A(n13800), .B(n13799), .Z(n13795) );
  AND U22068 ( .A(n13801), .B(n13802), .Z(n13756) );
  NAND U22069 ( .A(n13803), .B(n13804), .Z(n13802) );
  OR U22070 ( .A(n13805), .B(n13806), .Z(n13803) );
  NANDN U22071 ( .A(n13807), .B(n13805), .Z(n13801) );
  XNOR U22072 ( .A(n13782), .B(n13808), .Z(N64168) );
  XOR U22073 ( .A(n13784), .B(n13785), .Z(n13808) );
  XNOR U22074 ( .A(n13798), .B(n13809), .Z(n13785) );
  XOR U22075 ( .A(n13799), .B(n13800), .Z(n13809) );
  XOR U22076 ( .A(n13805), .B(n13810), .Z(n13800) );
  XOR U22077 ( .A(n13804), .B(n13807), .Z(n13810) );
  IV U22078 ( .A(n13806), .Z(n13807) );
  NAND U22079 ( .A(n13811), .B(n13812), .Z(n13806) );
  OR U22080 ( .A(n13813), .B(n13814), .Z(n13812) );
  OR U22081 ( .A(n13815), .B(n13816), .Z(n13811) );
  NAND U22082 ( .A(n13817), .B(n13818), .Z(n13804) );
  OR U22083 ( .A(n13819), .B(n13820), .Z(n13818) );
  OR U22084 ( .A(n13821), .B(n13822), .Z(n13817) );
  NOR U22085 ( .A(n13823), .B(n13824), .Z(n13805) );
  ANDN U22086 ( .B(n13825), .A(n13826), .Z(n13799) );
  XNOR U22087 ( .A(n13792), .B(n13827), .Z(n13798) );
  XNOR U22088 ( .A(n13791), .B(n13793), .Z(n13827) );
  NAND U22089 ( .A(n13828), .B(n13829), .Z(n13793) );
  OR U22090 ( .A(n13830), .B(n13831), .Z(n13829) );
  OR U22091 ( .A(n13832), .B(n13833), .Z(n13828) );
  NAND U22092 ( .A(n13834), .B(n13835), .Z(n13791) );
  OR U22093 ( .A(n13836), .B(n13837), .Z(n13835) );
  OR U22094 ( .A(n13838), .B(n13839), .Z(n13834) );
  ANDN U22095 ( .B(n13840), .A(n13841), .Z(n13792) );
  IV U22096 ( .A(n13842), .Z(n13840) );
  ANDN U22097 ( .B(n13843), .A(n13844), .Z(n13784) );
  XOR U22098 ( .A(n13770), .B(n13845), .Z(n13782) );
  XOR U22099 ( .A(n13771), .B(n13772), .Z(n13845) );
  XOR U22100 ( .A(n13777), .B(n13846), .Z(n13772) );
  XOR U22101 ( .A(n13776), .B(n13779), .Z(n13846) );
  IV U22102 ( .A(n13778), .Z(n13779) );
  NAND U22103 ( .A(n13847), .B(n13848), .Z(n13778) );
  OR U22104 ( .A(n13849), .B(n13850), .Z(n13848) );
  OR U22105 ( .A(n13851), .B(n13852), .Z(n13847) );
  NAND U22106 ( .A(n13853), .B(n13854), .Z(n13776) );
  OR U22107 ( .A(n13855), .B(n13856), .Z(n13854) );
  OR U22108 ( .A(n13857), .B(n13858), .Z(n13853) );
  NOR U22109 ( .A(n13859), .B(n13860), .Z(n13777) );
  ANDN U22110 ( .B(n13861), .A(n13862), .Z(n13771) );
  IV U22111 ( .A(n13863), .Z(n13861) );
  XNOR U22112 ( .A(n13764), .B(n13864), .Z(n13770) );
  XNOR U22113 ( .A(n13763), .B(n13765), .Z(n13864) );
  NAND U22114 ( .A(n13865), .B(n13866), .Z(n13765) );
  OR U22115 ( .A(n13867), .B(n13868), .Z(n13866) );
  OR U22116 ( .A(n13869), .B(n13870), .Z(n13865) );
  NAND U22117 ( .A(n13871), .B(n13872), .Z(n13763) );
  OR U22118 ( .A(n13873), .B(n13874), .Z(n13872) );
  OR U22119 ( .A(n13875), .B(n13876), .Z(n13871) );
  ANDN U22120 ( .B(n13877), .A(n13878), .Z(n13764) );
  IV U22121 ( .A(n13879), .Z(n13877) );
  XNOR U22122 ( .A(n13844), .B(n13843), .Z(N64167) );
  XOR U22123 ( .A(n13863), .B(n13862), .Z(n13843) );
  XNOR U22124 ( .A(n13878), .B(n13879), .Z(n13862) );
  XNOR U22125 ( .A(n13873), .B(n13874), .Z(n13879) );
  XNOR U22126 ( .A(n13875), .B(n13876), .Z(n13874) );
  XNOR U22127 ( .A(y[6613]), .B(x[6613]), .Z(n13876) );
  XNOR U22128 ( .A(y[6614]), .B(x[6614]), .Z(n13875) );
  XNOR U22129 ( .A(y[6612]), .B(x[6612]), .Z(n13873) );
  XNOR U22130 ( .A(n13867), .B(n13868), .Z(n13878) );
  XNOR U22131 ( .A(y[6609]), .B(x[6609]), .Z(n13868) );
  XNOR U22132 ( .A(n13869), .B(n13870), .Z(n13867) );
  XNOR U22133 ( .A(y[6610]), .B(x[6610]), .Z(n13870) );
  XNOR U22134 ( .A(y[6611]), .B(x[6611]), .Z(n13869) );
  XNOR U22135 ( .A(n13860), .B(n13859), .Z(n13863) );
  XNOR U22136 ( .A(n13855), .B(n13856), .Z(n13859) );
  XNOR U22137 ( .A(y[6606]), .B(x[6606]), .Z(n13856) );
  XNOR U22138 ( .A(n13857), .B(n13858), .Z(n13855) );
  XNOR U22139 ( .A(y[6607]), .B(x[6607]), .Z(n13858) );
  XNOR U22140 ( .A(y[6608]), .B(x[6608]), .Z(n13857) );
  XNOR U22141 ( .A(n13849), .B(n13850), .Z(n13860) );
  XNOR U22142 ( .A(y[6603]), .B(x[6603]), .Z(n13850) );
  XNOR U22143 ( .A(n13851), .B(n13852), .Z(n13849) );
  XNOR U22144 ( .A(y[6604]), .B(x[6604]), .Z(n13852) );
  XNOR U22145 ( .A(y[6605]), .B(x[6605]), .Z(n13851) );
  XOR U22146 ( .A(n13825), .B(n13826), .Z(n13844) );
  XNOR U22147 ( .A(n13841), .B(n13842), .Z(n13826) );
  XNOR U22148 ( .A(n13836), .B(n13837), .Z(n13842) );
  XNOR U22149 ( .A(n13838), .B(n13839), .Z(n13837) );
  XNOR U22150 ( .A(y[6601]), .B(x[6601]), .Z(n13839) );
  XNOR U22151 ( .A(y[6602]), .B(x[6602]), .Z(n13838) );
  XNOR U22152 ( .A(y[6600]), .B(x[6600]), .Z(n13836) );
  XNOR U22153 ( .A(n13830), .B(n13831), .Z(n13841) );
  XNOR U22154 ( .A(y[6597]), .B(x[6597]), .Z(n13831) );
  XNOR U22155 ( .A(n13832), .B(n13833), .Z(n13830) );
  XNOR U22156 ( .A(y[6598]), .B(x[6598]), .Z(n13833) );
  XNOR U22157 ( .A(y[6599]), .B(x[6599]), .Z(n13832) );
  XOR U22158 ( .A(n13824), .B(n13823), .Z(n13825) );
  XNOR U22159 ( .A(n13819), .B(n13820), .Z(n13823) );
  XNOR U22160 ( .A(y[6594]), .B(x[6594]), .Z(n13820) );
  XNOR U22161 ( .A(n13821), .B(n13822), .Z(n13819) );
  XNOR U22162 ( .A(y[6595]), .B(x[6595]), .Z(n13822) );
  XNOR U22163 ( .A(y[6596]), .B(x[6596]), .Z(n13821) );
  XNOR U22164 ( .A(n13813), .B(n13814), .Z(n13824) );
  XNOR U22165 ( .A(y[6591]), .B(x[6591]), .Z(n13814) );
  XNOR U22166 ( .A(n13815), .B(n13816), .Z(n13813) );
  XNOR U22167 ( .A(y[6592]), .B(x[6592]), .Z(n13816) );
  XNOR U22168 ( .A(y[6593]), .B(x[6593]), .Z(n13815) );
  NAND U22169 ( .A(n13880), .B(n13881), .Z(N64158) );
  NANDN U22170 ( .A(n13882), .B(n13883), .Z(n13881) );
  OR U22171 ( .A(n13884), .B(n13885), .Z(n13883) );
  NAND U22172 ( .A(n13884), .B(n13885), .Z(n13880) );
  XOR U22173 ( .A(n13884), .B(n13886), .Z(N64157) );
  XNOR U22174 ( .A(n13882), .B(n13885), .Z(n13886) );
  AND U22175 ( .A(n13887), .B(n13888), .Z(n13885) );
  NANDN U22176 ( .A(n13889), .B(n13890), .Z(n13888) );
  NANDN U22177 ( .A(n13891), .B(n13892), .Z(n13890) );
  NANDN U22178 ( .A(n13892), .B(n13891), .Z(n13887) );
  NAND U22179 ( .A(n13893), .B(n13894), .Z(n13882) );
  NANDN U22180 ( .A(n13895), .B(n13896), .Z(n13894) );
  OR U22181 ( .A(n13897), .B(n13898), .Z(n13896) );
  NAND U22182 ( .A(n13898), .B(n13897), .Z(n13893) );
  AND U22183 ( .A(n13899), .B(n13900), .Z(n13884) );
  NANDN U22184 ( .A(n13901), .B(n13902), .Z(n13900) );
  NANDN U22185 ( .A(n13903), .B(n13904), .Z(n13902) );
  NANDN U22186 ( .A(n13904), .B(n13903), .Z(n13899) );
  XOR U22187 ( .A(n13898), .B(n13905), .Z(N64156) );
  XOR U22188 ( .A(n13895), .B(n13897), .Z(n13905) );
  XNOR U22189 ( .A(n13891), .B(n13906), .Z(n13897) );
  XNOR U22190 ( .A(n13889), .B(n13892), .Z(n13906) );
  NAND U22191 ( .A(n13907), .B(n13908), .Z(n13892) );
  NAND U22192 ( .A(n13909), .B(n13910), .Z(n13908) );
  OR U22193 ( .A(n13911), .B(n13912), .Z(n13909) );
  NANDN U22194 ( .A(n13913), .B(n13911), .Z(n13907) );
  IV U22195 ( .A(n13912), .Z(n13913) );
  NAND U22196 ( .A(n13914), .B(n13915), .Z(n13889) );
  NAND U22197 ( .A(n13916), .B(n13917), .Z(n13915) );
  NANDN U22198 ( .A(n13918), .B(n13919), .Z(n13916) );
  NANDN U22199 ( .A(n13919), .B(n13918), .Z(n13914) );
  AND U22200 ( .A(n13920), .B(n13921), .Z(n13891) );
  NAND U22201 ( .A(n13922), .B(n13923), .Z(n13921) );
  OR U22202 ( .A(n13924), .B(n13925), .Z(n13922) );
  NANDN U22203 ( .A(n13926), .B(n13924), .Z(n13920) );
  NAND U22204 ( .A(n13927), .B(n13928), .Z(n13895) );
  NANDN U22205 ( .A(n13929), .B(n13930), .Z(n13928) );
  OR U22206 ( .A(n13931), .B(n13932), .Z(n13930) );
  NANDN U22207 ( .A(n13933), .B(n13931), .Z(n13927) );
  IV U22208 ( .A(n13932), .Z(n13933) );
  XNOR U22209 ( .A(n13903), .B(n13934), .Z(n13898) );
  XNOR U22210 ( .A(n13901), .B(n13904), .Z(n13934) );
  NAND U22211 ( .A(n13935), .B(n13936), .Z(n13904) );
  NAND U22212 ( .A(n13937), .B(n13938), .Z(n13936) );
  OR U22213 ( .A(n13939), .B(n13940), .Z(n13937) );
  NANDN U22214 ( .A(n13941), .B(n13939), .Z(n13935) );
  IV U22215 ( .A(n13940), .Z(n13941) );
  NAND U22216 ( .A(n13942), .B(n13943), .Z(n13901) );
  NAND U22217 ( .A(n13944), .B(n13945), .Z(n13943) );
  NANDN U22218 ( .A(n13946), .B(n13947), .Z(n13944) );
  NANDN U22219 ( .A(n13947), .B(n13946), .Z(n13942) );
  AND U22220 ( .A(n13948), .B(n13949), .Z(n13903) );
  NAND U22221 ( .A(n13950), .B(n13951), .Z(n13949) );
  OR U22222 ( .A(n13952), .B(n13953), .Z(n13950) );
  NANDN U22223 ( .A(n13954), .B(n13952), .Z(n13948) );
  XNOR U22224 ( .A(n13929), .B(n13955), .Z(N64155) );
  XOR U22225 ( .A(n13931), .B(n13932), .Z(n13955) );
  XNOR U22226 ( .A(n13945), .B(n13956), .Z(n13932) );
  XOR U22227 ( .A(n13946), .B(n13947), .Z(n13956) );
  XOR U22228 ( .A(n13952), .B(n13957), .Z(n13947) );
  XOR U22229 ( .A(n13951), .B(n13954), .Z(n13957) );
  IV U22230 ( .A(n13953), .Z(n13954) );
  NAND U22231 ( .A(n13958), .B(n13959), .Z(n13953) );
  OR U22232 ( .A(n13960), .B(n13961), .Z(n13959) );
  OR U22233 ( .A(n13962), .B(n13963), .Z(n13958) );
  NAND U22234 ( .A(n13964), .B(n13965), .Z(n13951) );
  OR U22235 ( .A(n13966), .B(n13967), .Z(n13965) );
  OR U22236 ( .A(n13968), .B(n13969), .Z(n13964) );
  NOR U22237 ( .A(n13970), .B(n13971), .Z(n13952) );
  ANDN U22238 ( .B(n13972), .A(n13973), .Z(n13946) );
  XNOR U22239 ( .A(n13939), .B(n13974), .Z(n13945) );
  XNOR U22240 ( .A(n13938), .B(n13940), .Z(n13974) );
  NAND U22241 ( .A(n13975), .B(n13976), .Z(n13940) );
  OR U22242 ( .A(n13977), .B(n13978), .Z(n13976) );
  OR U22243 ( .A(n13979), .B(n13980), .Z(n13975) );
  NAND U22244 ( .A(n13981), .B(n13982), .Z(n13938) );
  OR U22245 ( .A(n13983), .B(n13984), .Z(n13982) );
  OR U22246 ( .A(n13985), .B(n13986), .Z(n13981) );
  ANDN U22247 ( .B(n13987), .A(n13988), .Z(n13939) );
  IV U22248 ( .A(n13989), .Z(n13987) );
  ANDN U22249 ( .B(n13990), .A(n13991), .Z(n13931) );
  XOR U22250 ( .A(n13917), .B(n13992), .Z(n13929) );
  XOR U22251 ( .A(n13918), .B(n13919), .Z(n13992) );
  XOR U22252 ( .A(n13924), .B(n13993), .Z(n13919) );
  XOR U22253 ( .A(n13923), .B(n13926), .Z(n13993) );
  IV U22254 ( .A(n13925), .Z(n13926) );
  NAND U22255 ( .A(n13994), .B(n13995), .Z(n13925) );
  OR U22256 ( .A(n13996), .B(n13997), .Z(n13995) );
  OR U22257 ( .A(n13998), .B(n13999), .Z(n13994) );
  NAND U22258 ( .A(n14000), .B(n14001), .Z(n13923) );
  OR U22259 ( .A(n14002), .B(n14003), .Z(n14001) );
  OR U22260 ( .A(n14004), .B(n14005), .Z(n14000) );
  NOR U22261 ( .A(n14006), .B(n14007), .Z(n13924) );
  ANDN U22262 ( .B(n14008), .A(n14009), .Z(n13918) );
  IV U22263 ( .A(n14010), .Z(n14008) );
  XNOR U22264 ( .A(n13911), .B(n14011), .Z(n13917) );
  XNOR U22265 ( .A(n13910), .B(n13912), .Z(n14011) );
  NAND U22266 ( .A(n14012), .B(n14013), .Z(n13912) );
  OR U22267 ( .A(n14014), .B(n14015), .Z(n14013) );
  OR U22268 ( .A(n14016), .B(n14017), .Z(n14012) );
  NAND U22269 ( .A(n14018), .B(n14019), .Z(n13910) );
  OR U22270 ( .A(n14020), .B(n14021), .Z(n14019) );
  OR U22271 ( .A(n14022), .B(n14023), .Z(n14018) );
  ANDN U22272 ( .B(n14024), .A(n14025), .Z(n13911) );
  IV U22273 ( .A(n14026), .Z(n14024) );
  XNOR U22274 ( .A(n13991), .B(n13990), .Z(N64154) );
  XOR U22275 ( .A(n14010), .B(n14009), .Z(n13990) );
  XNOR U22276 ( .A(n14025), .B(n14026), .Z(n14009) );
  XNOR U22277 ( .A(n14020), .B(n14021), .Z(n14026) );
  XNOR U22278 ( .A(n14022), .B(n14023), .Z(n14021) );
  XNOR U22279 ( .A(y[6589]), .B(x[6589]), .Z(n14023) );
  XNOR U22280 ( .A(y[6590]), .B(x[6590]), .Z(n14022) );
  XNOR U22281 ( .A(y[6588]), .B(x[6588]), .Z(n14020) );
  XNOR U22282 ( .A(n14014), .B(n14015), .Z(n14025) );
  XNOR U22283 ( .A(y[6585]), .B(x[6585]), .Z(n14015) );
  XNOR U22284 ( .A(n14016), .B(n14017), .Z(n14014) );
  XNOR U22285 ( .A(y[6586]), .B(x[6586]), .Z(n14017) );
  XNOR U22286 ( .A(y[6587]), .B(x[6587]), .Z(n14016) );
  XNOR U22287 ( .A(n14007), .B(n14006), .Z(n14010) );
  XNOR U22288 ( .A(n14002), .B(n14003), .Z(n14006) );
  XNOR U22289 ( .A(y[6582]), .B(x[6582]), .Z(n14003) );
  XNOR U22290 ( .A(n14004), .B(n14005), .Z(n14002) );
  XNOR U22291 ( .A(y[6583]), .B(x[6583]), .Z(n14005) );
  XNOR U22292 ( .A(y[6584]), .B(x[6584]), .Z(n14004) );
  XNOR U22293 ( .A(n13996), .B(n13997), .Z(n14007) );
  XNOR U22294 ( .A(y[6579]), .B(x[6579]), .Z(n13997) );
  XNOR U22295 ( .A(n13998), .B(n13999), .Z(n13996) );
  XNOR U22296 ( .A(y[6580]), .B(x[6580]), .Z(n13999) );
  XNOR U22297 ( .A(y[6581]), .B(x[6581]), .Z(n13998) );
  XOR U22298 ( .A(n13972), .B(n13973), .Z(n13991) );
  XNOR U22299 ( .A(n13988), .B(n13989), .Z(n13973) );
  XNOR U22300 ( .A(n13983), .B(n13984), .Z(n13989) );
  XNOR U22301 ( .A(n13985), .B(n13986), .Z(n13984) );
  XNOR U22302 ( .A(y[6577]), .B(x[6577]), .Z(n13986) );
  XNOR U22303 ( .A(y[6578]), .B(x[6578]), .Z(n13985) );
  XNOR U22304 ( .A(y[6576]), .B(x[6576]), .Z(n13983) );
  XNOR U22305 ( .A(n13977), .B(n13978), .Z(n13988) );
  XNOR U22306 ( .A(y[6573]), .B(x[6573]), .Z(n13978) );
  XNOR U22307 ( .A(n13979), .B(n13980), .Z(n13977) );
  XNOR U22308 ( .A(y[6574]), .B(x[6574]), .Z(n13980) );
  XNOR U22309 ( .A(y[6575]), .B(x[6575]), .Z(n13979) );
  XOR U22310 ( .A(n13971), .B(n13970), .Z(n13972) );
  XNOR U22311 ( .A(n13966), .B(n13967), .Z(n13970) );
  XNOR U22312 ( .A(y[6570]), .B(x[6570]), .Z(n13967) );
  XNOR U22313 ( .A(n13968), .B(n13969), .Z(n13966) );
  XNOR U22314 ( .A(y[6571]), .B(x[6571]), .Z(n13969) );
  XNOR U22315 ( .A(y[6572]), .B(x[6572]), .Z(n13968) );
  XNOR U22316 ( .A(n13960), .B(n13961), .Z(n13971) );
  XNOR U22317 ( .A(y[6567]), .B(x[6567]), .Z(n13961) );
  XNOR U22318 ( .A(n13962), .B(n13963), .Z(n13960) );
  XNOR U22319 ( .A(y[6568]), .B(x[6568]), .Z(n13963) );
  XNOR U22320 ( .A(y[6569]), .B(x[6569]), .Z(n13962) );
  NAND U22321 ( .A(n14027), .B(n14028), .Z(N64145) );
  NANDN U22322 ( .A(n14029), .B(n14030), .Z(n14028) );
  OR U22323 ( .A(n14031), .B(n14032), .Z(n14030) );
  NAND U22324 ( .A(n14031), .B(n14032), .Z(n14027) );
  XOR U22325 ( .A(n14031), .B(n14033), .Z(N64144) );
  XNOR U22326 ( .A(n14029), .B(n14032), .Z(n14033) );
  AND U22327 ( .A(n14034), .B(n14035), .Z(n14032) );
  NANDN U22328 ( .A(n14036), .B(n14037), .Z(n14035) );
  NANDN U22329 ( .A(n14038), .B(n14039), .Z(n14037) );
  NANDN U22330 ( .A(n14039), .B(n14038), .Z(n14034) );
  NAND U22331 ( .A(n14040), .B(n14041), .Z(n14029) );
  NANDN U22332 ( .A(n14042), .B(n14043), .Z(n14041) );
  OR U22333 ( .A(n14044), .B(n14045), .Z(n14043) );
  NAND U22334 ( .A(n14045), .B(n14044), .Z(n14040) );
  AND U22335 ( .A(n14046), .B(n14047), .Z(n14031) );
  NANDN U22336 ( .A(n14048), .B(n14049), .Z(n14047) );
  NANDN U22337 ( .A(n14050), .B(n14051), .Z(n14049) );
  NANDN U22338 ( .A(n14051), .B(n14050), .Z(n14046) );
  XOR U22339 ( .A(n14045), .B(n14052), .Z(N64143) );
  XOR U22340 ( .A(n14042), .B(n14044), .Z(n14052) );
  XNOR U22341 ( .A(n14038), .B(n14053), .Z(n14044) );
  XNOR U22342 ( .A(n14036), .B(n14039), .Z(n14053) );
  NAND U22343 ( .A(n14054), .B(n14055), .Z(n14039) );
  NAND U22344 ( .A(n14056), .B(n14057), .Z(n14055) );
  OR U22345 ( .A(n14058), .B(n14059), .Z(n14056) );
  NANDN U22346 ( .A(n14060), .B(n14058), .Z(n14054) );
  IV U22347 ( .A(n14059), .Z(n14060) );
  NAND U22348 ( .A(n14061), .B(n14062), .Z(n14036) );
  NAND U22349 ( .A(n14063), .B(n14064), .Z(n14062) );
  NANDN U22350 ( .A(n14065), .B(n14066), .Z(n14063) );
  NANDN U22351 ( .A(n14066), .B(n14065), .Z(n14061) );
  AND U22352 ( .A(n14067), .B(n14068), .Z(n14038) );
  NAND U22353 ( .A(n14069), .B(n14070), .Z(n14068) );
  OR U22354 ( .A(n14071), .B(n14072), .Z(n14069) );
  NANDN U22355 ( .A(n14073), .B(n14071), .Z(n14067) );
  NAND U22356 ( .A(n14074), .B(n14075), .Z(n14042) );
  NANDN U22357 ( .A(n14076), .B(n14077), .Z(n14075) );
  OR U22358 ( .A(n14078), .B(n14079), .Z(n14077) );
  NANDN U22359 ( .A(n14080), .B(n14078), .Z(n14074) );
  IV U22360 ( .A(n14079), .Z(n14080) );
  XNOR U22361 ( .A(n14050), .B(n14081), .Z(n14045) );
  XNOR U22362 ( .A(n14048), .B(n14051), .Z(n14081) );
  NAND U22363 ( .A(n14082), .B(n14083), .Z(n14051) );
  NAND U22364 ( .A(n14084), .B(n14085), .Z(n14083) );
  OR U22365 ( .A(n14086), .B(n14087), .Z(n14084) );
  NANDN U22366 ( .A(n14088), .B(n14086), .Z(n14082) );
  IV U22367 ( .A(n14087), .Z(n14088) );
  NAND U22368 ( .A(n14089), .B(n14090), .Z(n14048) );
  NAND U22369 ( .A(n14091), .B(n14092), .Z(n14090) );
  NANDN U22370 ( .A(n14093), .B(n14094), .Z(n14091) );
  NANDN U22371 ( .A(n14094), .B(n14093), .Z(n14089) );
  AND U22372 ( .A(n14095), .B(n14096), .Z(n14050) );
  NAND U22373 ( .A(n14097), .B(n14098), .Z(n14096) );
  OR U22374 ( .A(n14099), .B(n14100), .Z(n14097) );
  NANDN U22375 ( .A(n14101), .B(n14099), .Z(n14095) );
  XNOR U22376 ( .A(n14076), .B(n14102), .Z(N64142) );
  XOR U22377 ( .A(n14078), .B(n14079), .Z(n14102) );
  XNOR U22378 ( .A(n14092), .B(n14103), .Z(n14079) );
  XOR U22379 ( .A(n14093), .B(n14094), .Z(n14103) );
  XOR U22380 ( .A(n14099), .B(n14104), .Z(n14094) );
  XOR U22381 ( .A(n14098), .B(n14101), .Z(n14104) );
  IV U22382 ( .A(n14100), .Z(n14101) );
  NAND U22383 ( .A(n14105), .B(n14106), .Z(n14100) );
  OR U22384 ( .A(n14107), .B(n14108), .Z(n14106) );
  OR U22385 ( .A(n14109), .B(n14110), .Z(n14105) );
  NAND U22386 ( .A(n14111), .B(n14112), .Z(n14098) );
  OR U22387 ( .A(n14113), .B(n14114), .Z(n14112) );
  OR U22388 ( .A(n14115), .B(n14116), .Z(n14111) );
  NOR U22389 ( .A(n14117), .B(n14118), .Z(n14099) );
  ANDN U22390 ( .B(n14119), .A(n14120), .Z(n14093) );
  XNOR U22391 ( .A(n14086), .B(n14121), .Z(n14092) );
  XNOR U22392 ( .A(n14085), .B(n14087), .Z(n14121) );
  NAND U22393 ( .A(n14122), .B(n14123), .Z(n14087) );
  OR U22394 ( .A(n14124), .B(n14125), .Z(n14123) );
  OR U22395 ( .A(n14126), .B(n14127), .Z(n14122) );
  NAND U22396 ( .A(n14128), .B(n14129), .Z(n14085) );
  OR U22397 ( .A(n14130), .B(n14131), .Z(n14129) );
  OR U22398 ( .A(n14132), .B(n14133), .Z(n14128) );
  ANDN U22399 ( .B(n14134), .A(n14135), .Z(n14086) );
  IV U22400 ( .A(n14136), .Z(n14134) );
  ANDN U22401 ( .B(n14137), .A(n14138), .Z(n14078) );
  XOR U22402 ( .A(n14064), .B(n14139), .Z(n14076) );
  XOR U22403 ( .A(n14065), .B(n14066), .Z(n14139) );
  XOR U22404 ( .A(n14071), .B(n14140), .Z(n14066) );
  XOR U22405 ( .A(n14070), .B(n14073), .Z(n14140) );
  IV U22406 ( .A(n14072), .Z(n14073) );
  NAND U22407 ( .A(n14141), .B(n14142), .Z(n14072) );
  OR U22408 ( .A(n14143), .B(n14144), .Z(n14142) );
  OR U22409 ( .A(n14145), .B(n14146), .Z(n14141) );
  NAND U22410 ( .A(n14147), .B(n14148), .Z(n14070) );
  OR U22411 ( .A(n14149), .B(n14150), .Z(n14148) );
  OR U22412 ( .A(n14151), .B(n14152), .Z(n14147) );
  NOR U22413 ( .A(n14153), .B(n14154), .Z(n14071) );
  ANDN U22414 ( .B(n14155), .A(n14156), .Z(n14065) );
  IV U22415 ( .A(n14157), .Z(n14155) );
  XNOR U22416 ( .A(n14058), .B(n14158), .Z(n14064) );
  XNOR U22417 ( .A(n14057), .B(n14059), .Z(n14158) );
  NAND U22418 ( .A(n14159), .B(n14160), .Z(n14059) );
  OR U22419 ( .A(n14161), .B(n14162), .Z(n14160) );
  OR U22420 ( .A(n14163), .B(n14164), .Z(n14159) );
  NAND U22421 ( .A(n14165), .B(n14166), .Z(n14057) );
  OR U22422 ( .A(n14167), .B(n14168), .Z(n14166) );
  OR U22423 ( .A(n14169), .B(n14170), .Z(n14165) );
  ANDN U22424 ( .B(n14171), .A(n14172), .Z(n14058) );
  IV U22425 ( .A(n14173), .Z(n14171) );
  XNOR U22426 ( .A(n14138), .B(n14137), .Z(N64141) );
  XOR U22427 ( .A(n14157), .B(n14156), .Z(n14137) );
  XNOR U22428 ( .A(n14172), .B(n14173), .Z(n14156) );
  XNOR U22429 ( .A(n14167), .B(n14168), .Z(n14173) );
  XNOR U22430 ( .A(n14169), .B(n14170), .Z(n14168) );
  XNOR U22431 ( .A(y[6565]), .B(x[6565]), .Z(n14170) );
  XNOR U22432 ( .A(y[6566]), .B(x[6566]), .Z(n14169) );
  XNOR U22433 ( .A(y[6564]), .B(x[6564]), .Z(n14167) );
  XNOR U22434 ( .A(n14161), .B(n14162), .Z(n14172) );
  XNOR U22435 ( .A(y[6561]), .B(x[6561]), .Z(n14162) );
  XNOR U22436 ( .A(n14163), .B(n14164), .Z(n14161) );
  XNOR U22437 ( .A(y[6562]), .B(x[6562]), .Z(n14164) );
  XNOR U22438 ( .A(y[6563]), .B(x[6563]), .Z(n14163) );
  XNOR U22439 ( .A(n14154), .B(n14153), .Z(n14157) );
  XNOR U22440 ( .A(n14149), .B(n14150), .Z(n14153) );
  XNOR U22441 ( .A(y[6558]), .B(x[6558]), .Z(n14150) );
  XNOR U22442 ( .A(n14151), .B(n14152), .Z(n14149) );
  XNOR U22443 ( .A(y[6559]), .B(x[6559]), .Z(n14152) );
  XNOR U22444 ( .A(y[6560]), .B(x[6560]), .Z(n14151) );
  XNOR U22445 ( .A(n14143), .B(n14144), .Z(n14154) );
  XNOR U22446 ( .A(y[6555]), .B(x[6555]), .Z(n14144) );
  XNOR U22447 ( .A(n14145), .B(n14146), .Z(n14143) );
  XNOR U22448 ( .A(y[6556]), .B(x[6556]), .Z(n14146) );
  XNOR U22449 ( .A(y[6557]), .B(x[6557]), .Z(n14145) );
  XOR U22450 ( .A(n14119), .B(n14120), .Z(n14138) );
  XNOR U22451 ( .A(n14135), .B(n14136), .Z(n14120) );
  XNOR U22452 ( .A(n14130), .B(n14131), .Z(n14136) );
  XNOR U22453 ( .A(n14132), .B(n14133), .Z(n14131) );
  XNOR U22454 ( .A(y[6553]), .B(x[6553]), .Z(n14133) );
  XNOR U22455 ( .A(y[6554]), .B(x[6554]), .Z(n14132) );
  XNOR U22456 ( .A(y[6552]), .B(x[6552]), .Z(n14130) );
  XNOR U22457 ( .A(n14124), .B(n14125), .Z(n14135) );
  XNOR U22458 ( .A(y[6549]), .B(x[6549]), .Z(n14125) );
  XNOR U22459 ( .A(n14126), .B(n14127), .Z(n14124) );
  XNOR U22460 ( .A(y[6550]), .B(x[6550]), .Z(n14127) );
  XNOR U22461 ( .A(y[6551]), .B(x[6551]), .Z(n14126) );
  XOR U22462 ( .A(n14118), .B(n14117), .Z(n14119) );
  XNOR U22463 ( .A(n14113), .B(n14114), .Z(n14117) );
  XNOR U22464 ( .A(y[6546]), .B(x[6546]), .Z(n14114) );
  XNOR U22465 ( .A(n14115), .B(n14116), .Z(n14113) );
  XNOR U22466 ( .A(y[6547]), .B(x[6547]), .Z(n14116) );
  XNOR U22467 ( .A(y[6548]), .B(x[6548]), .Z(n14115) );
  XNOR U22468 ( .A(n14107), .B(n14108), .Z(n14118) );
  XNOR U22469 ( .A(y[6543]), .B(x[6543]), .Z(n14108) );
  XNOR U22470 ( .A(n14109), .B(n14110), .Z(n14107) );
  XNOR U22471 ( .A(y[6544]), .B(x[6544]), .Z(n14110) );
  XNOR U22472 ( .A(y[6545]), .B(x[6545]), .Z(n14109) );
  NAND U22473 ( .A(n14174), .B(n14175), .Z(N64132) );
  NANDN U22474 ( .A(n14176), .B(n14177), .Z(n14175) );
  OR U22475 ( .A(n14178), .B(n14179), .Z(n14177) );
  NAND U22476 ( .A(n14178), .B(n14179), .Z(n14174) );
  XOR U22477 ( .A(n14178), .B(n14180), .Z(N64131) );
  XNOR U22478 ( .A(n14176), .B(n14179), .Z(n14180) );
  AND U22479 ( .A(n14181), .B(n14182), .Z(n14179) );
  NANDN U22480 ( .A(n14183), .B(n14184), .Z(n14182) );
  NANDN U22481 ( .A(n14185), .B(n14186), .Z(n14184) );
  NANDN U22482 ( .A(n14186), .B(n14185), .Z(n14181) );
  NAND U22483 ( .A(n14187), .B(n14188), .Z(n14176) );
  NANDN U22484 ( .A(n14189), .B(n14190), .Z(n14188) );
  OR U22485 ( .A(n14191), .B(n14192), .Z(n14190) );
  NAND U22486 ( .A(n14192), .B(n14191), .Z(n14187) );
  AND U22487 ( .A(n14193), .B(n14194), .Z(n14178) );
  NANDN U22488 ( .A(n14195), .B(n14196), .Z(n14194) );
  NANDN U22489 ( .A(n14197), .B(n14198), .Z(n14196) );
  NANDN U22490 ( .A(n14198), .B(n14197), .Z(n14193) );
  XOR U22491 ( .A(n14192), .B(n14199), .Z(N64130) );
  XOR U22492 ( .A(n14189), .B(n14191), .Z(n14199) );
  XNOR U22493 ( .A(n14185), .B(n14200), .Z(n14191) );
  XNOR U22494 ( .A(n14183), .B(n14186), .Z(n14200) );
  NAND U22495 ( .A(n14201), .B(n14202), .Z(n14186) );
  NAND U22496 ( .A(n14203), .B(n14204), .Z(n14202) );
  OR U22497 ( .A(n14205), .B(n14206), .Z(n14203) );
  NANDN U22498 ( .A(n14207), .B(n14205), .Z(n14201) );
  IV U22499 ( .A(n14206), .Z(n14207) );
  NAND U22500 ( .A(n14208), .B(n14209), .Z(n14183) );
  NAND U22501 ( .A(n14210), .B(n14211), .Z(n14209) );
  NANDN U22502 ( .A(n14212), .B(n14213), .Z(n14210) );
  NANDN U22503 ( .A(n14213), .B(n14212), .Z(n14208) );
  AND U22504 ( .A(n14214), .B(n14215), .Z(n14185) );
  NAND U22505 ( .A(n14216), .B(n14217), .Z(n14215) );
  OR U22506 ( .A(n14218), .B(n14219), .Z(n14216) );
  NANDN U22507 ( .A(n14220), .B(n14218), .Z(n14214) );
  NAND U22508 ( .A(n14221), .B(n14222), .Z(n14189) );
  NANDN U22509 ( .A(n14223), .B(n14224), .Z(n14222) );
  OR U22510 ( .A(n14225), .B(n14226), .Z(n14224) );
  NANDN U22511 ( .A(n14227), .B(n14225), .Z(n14221) );
  IV U22512 ( .A(n14226), .Z(n14227) );
  XNOR U22513 ( .A(n14197), .B(n14228), .Z(n14192) );
  XNOR U22514 ( .A(n14195), .B(n14198), .Z(n14228) );
  NAND U22515 ( .A(n14229), .B(n14230), .Z(n14198) );
  NAND U22516 ( .A(n14231), .B(n14232), .Z(n14230) );
  OR U22517 ( .A(n14233), .B(n14234), .Z(n14231) );
  NANDN U22518 ( .A(n14235), .B(n14233), .Z(n14229) );
  IV U22519 ( .A(n14234), .Z(n14235) );
  NAND U22520 ( .A(n14236), .B(n14237), .Z(n14195) );
  NAND U22521 ( .A(n14238), .B(n14239), .Z(n14237) );
  NANDN U22522 ( .A(n14240), .B(n14241), .Z(n14238) );
  NANDN U22523 ( .A(n14241), .B(n14240), .Z(n14236) );
  AND U22524 ( .A(n14242), .B(n14243), .Z(n14197) );
  NAND U22525 ( .A(n14244), .B(n14245), .Z(n14243) );
  OR U22526 ( .A(n14246), .B(n14247), .Z(n14244) );
  NANDN U22527 ( .A(n14248), .B(n14246), .Z(n14242) );
  XNOR U22528 ( .A(n14223), .B(n14249), .Z(N64129) );
  XOR U22529 ( .A(n14225), .B(n14226), .Z(n14249) );
  XNOR U22530 ( .A(n14239), .B(n14250), .Z(n14226) );
  XOR U22531 ( .A(n14240), .B(n14241), .Z(n14250) );
  XOR U22532 ( .A(n14246), .B(n14251), .Z(n14241) );
  XOR U22533 ( .A(n14245), .B(n14248), .Z(n14251) );
  IV U22534 ( .A(n14247), .Z(n14248) );
  NAND U22535 ( .A(n14252), .B(n14253), .Z(n14247) );
  OR U22536 ( .A(n14254), .B(n14255), .Z(n14253) );
  OR U22537 ( .A(n14256), .B(n14257), .Z(n14252) );
  NAND U22538 ( .A(n14258), .B(n14259), .Z(n14245) );
  OR U22539 ( .A(n14260), .B(n14261), .Z(n14259) );
  OR U22540 ( .A(n14262), .B(n14263), .Z(n14258) );
  NOR U22541 ( .A(n14264), .B(n14265), .Z(n14246) );
  ANDN U22542 ( .B(n14266), .A(n14267), .Z(n14240) );
  XNOR U22543 ( .A(n14233), .B(n14268), .Z(n14239) );
  XNOR U22544 ( .A(n14232), .B(n14234), .Z(n14268) );
  NAND U22545 ( .A(n14269), .B(n14270), .Z(n14234) );
  OR U22546 ( .A(n14271), .B(n14272), .Z(n14270) );
  OR U22547 ( .A(n14273), .B(n14274), .Z(n14269) );
  NAND U22548 ( .A(n14275), .B(n14276), .Z(n14232) );
  OR U22549 ( .A(n14277), .B(n14278), .Z(n14276) );
  OR U22550 ( .A(n14279), .B(n14280), .Z(n14275) );
  ANDN U22551 ( .B(n14281), .A(n14282), .Z(n14233) );
  IV U22552 ( .A(n14283), .Z(n14281) );
  ANDN U22553 ( .B(n14284), .A(n14285), .Z(n14225) );
  XOR U22554 ( .A(n14211), .B(n14286), .Z(n14223) );
  XOR U22555 ( .A(n14212), .B(n14213), .Z(n14286) );
  XOR U22556 ( .A(n14218), .B(n14287), .Z(n14213) );
  XOR U22557 ( .A(n14217), .B(n14220), .Z(n14287) );
  IV U22558 ( .A(n14219), .Z(n14220) );
  NAND U22559 ( .A(n14288), .B(n14289), .Z(n14219) );
  OR U22560 ( .A(n14290), .B(n14291), .Z(n14289) );
  OR U22561 ( .A(n14292), .B(n14293), .Z(n14288) );
  NAND U22562 ( .A(n14294), .B(n14295), .Z(n14217) );
  OR U22563 ( .A(n14296), .B(n14297), .Z(n14295) );
  OR U22564 ( .A(n14298), .B(n14299), .Z(n14294) );
  NOR U22565 ( .A(n14300), .B(n14301), .Z(n14218) );
  ANDN U22566 ( .B(n14302), .A(n14303), .Z(n14212) );
  IV U22567 ( .A(n14304), .Z(n14302) );
  XNOR U22568 ( .A(n14205), .B(n14305), .Z(n14211) );
  XNOR U22569 ( .A(n14204), .B(n14206), .Z(n14305) );
  NAND U22570 ( .A(n14306), .B(n14307), .Z(n14206) );
  OR U22571 ( .A(n14308), .B(n14309), .Z(n14307) );
  OR U22572 ( .A(n14310), .B(n14311), .Z(n14306) );
  NAND U22573 ( .A(n14312), .B(n14313), .Z(n14204) );
  OR U22574 ( .A(n14314), .B(n14315), .Z(n14313) );
  OR U22575 ( .A(n14316), .B(n14317), .Z(n14312) );
  ANDN U22576 ( .B(n14318), .A(n14319), .Z(n14205) );
  IV U22577 ( .A(n14320), .Z(n14318) );
  XNOR U22578 ( .A(n14285), .B(n14284), .Z(N64128) );
  XOR U22579 ( .A(n14304), .B(n14303), .Z(n14284) );
  XNOR U22580 ( .A(n14319), .B(n14320), .Z(n14303) );
  XNOR U22581 ( .A(n14314), .B(n14315), .Z(n14320) );
  XNOR U22582 ( .A(n14316), .B(n14317), .Z(n14315) );
  XNOR U22583 ( .A(y[6541]), .B(x[6541]), .Z(n14317) );
  XNOR U22584 ( .A(y[6542]), .B(x[6542]), .Z(n14316) );
  XNOR U22585 ( .A(y[6540]), .B(x[6540]), .Z(n14314) );
  XNOR U22586 ( .A(n14308), .B(n14309), .Z(n14319) );
  XNOR U22587 ( .A(y[6537]), .B(x[6537]), .Z(n14309) );
  XNOR U22588 ( .A(n14310), .B(n14311), .Z(n14308) );
  XNOR U22589 ( .A(y[6538]), .B(x[6538]), .Z(n14311) );
  XNOR U22590 ( .A(y[6539]), .B(x[6539]), .Z(n14310) );
  XNOR U22591 ( .A(n14301), .B(n14300), .Z(n14304) );
  XNOR U22592 ( .A(n14296), .B(n14297), .Z(n14300) );
  XNOR U22593 ( .A(y[6534]), .B(x[6534]), .Z(n14297) );
  XNOR U22594 ( .A(n14298), .B(n14299), .Z(n14296) );
  XNOR U22595 ( .A(y[6535]), .B(x[6535]), .Z(n14299) );
  XNOR U22596 ( .A(y[6536]), .B(x[6536]), .Z(n14298) );
  XNOR U22597 ( .A(n14290), .B(n14291), .Z(n14301) );
  XNOR U22598 ( .A(y[6531]), .B(x[6531]), .Z(n14291) );
  XNOR U22599 ( .A(n14292), .B(n14293), .Z(n14290) );
  XNOR U22600 ( .A(y[6532]), .B(x[6532]), .Z(n14293) );
  XNOR U22601 ( .A(y[6533]), .B(x[6533]), .Z(n14292) );
  XOR U22602 ( .A(n14266), .B(n14267), .Z(n14285) );
  XNOR U22603 ( .A(n14282), .B(n14283), .Z(n14267) );
  XNOR U22604 ( .A(n14277), .B(n14278), .Z(n14283) );
  XNOR U22605 ( .A(n14279), .B(n14280), .Z(n14278) );
  XNOR U22606 ( .A(y[6529]), .B(x[6529]), .Z(n14280) );
  XNOR U22607 ( .A(y[6530]), .B(x[6530]), .Z(n14279) );
  XNOR U22608 ( .A(y[6528]), .B(x[6528]), .Z(n14277) );
  XNOR U22609 ( .A(n14271), .B(n14272), .Z(n14282) );
  XNOR U22610 ( .A(y[6525]), .B(x[6525]), .Z(n14272) );
  XNOR U22611 ( .A(n14273), .B(n14274), .Z(n14271) );
  XNOR U22612 ( .A(y[6526]), .B(x[6526]), .Z(n14274) );
  XNOR U22613 ( .A(y[6527]), .B(x[6527]), .Z(n14273) );
  XOR U22614 ( .A(n14265), .B(n14264), .Z(n14266) );
  XNOR U22615 ( .A(n14260), .B(n14261), .Z(n14264) );
  XNOR U22616 ( .A(y[6522]), .B(x[6522]), .Z(n14261) );
  XNOR U22617 ( .A(n14262), .B(n14263), .Z(n14260) );
  XNOR U22618 ( .A(y[6523]), .B(x[6523]), .Z(n14263) );
  XNOR U22619 ( .A(y[6524]), .B(x[6524]), .Z(n14262) );
  XNOR U22620 ( .A(n14254), .B(n14255), .Z(n14265) );
  XNOR U22621 ( .A(y[6519]), .B(x[6519]), .Z(n14255) );
  XNOR U22622 ( .A(n14256), .B(n14257), .Z(n14254) );
  XNOR U22623 ( .A(y[6520]), .B(x[6520]), .Z(n14257) );
  XNOR U22624 ( .A(y[6521]), .B(x[6521]), .Z(n14256) );
  NAND U22625 ( .A(n14321), .B(n14322), .Z(N64119) );
  NANDN U22626 ( .A(n14323), .B(n14324), .Z(n14322) );
  OR U22627 ( .A(n14325), .B(n14326), .Z(n14324) );
  NAND U22628 ( .A(n14325), .B(n14326), .Z(n14321) );
  XOR U22629 ( .A(n14325), .B(n14327), .Z(N64118) );
  XNOR U22630 ( .A(n14323), .B(n14326), .Z(n14327) );
  AND U22631 ( .A(n14328), .B(n14329), .Z(n14326) );
  NANDN U22632 ( .A(n14330), .B(n14331), .Z(n14329) );
  NANDN U22633 ( .A(n14332), .B(n14333), .Z(n14331) );
  NANDN U22634 ( .A(n14333), .B(n14332), .Z(n14328) );
  NAND U22635 ( .A(n14334), .B(n14335), .Z(n14323) );
  NANDN U22636 ( .A(n14336), .B(n14337), .Z(n14335) );
  OR U22637 ( .A(n14338), .B(n14339), .Z(n14337) );
  NAND U22638 ( .A(n14339), .B(n14338), .Z(n14334) );
  AND U22639 ( .A(n14340), .B(n14341), .Z(n14325) );
  NANDN U22640 ( .A(n14342), .B(n14343), .Z(n14341) );
  NANDN U22641 ( .A(n14344), .B(n14345), .Z(n14343) );
  NANDN U22642 ( .A(n14345), .B(n14344), .Z(n14340) );
  XOR U22643 ( .A(n14339), .B(n14346), .Z(N64117) );
  XOR U22644 ( .A(n14336), .B(n14338), .Z(n14346) );
  XNOR U22645 ( .A(n14332), .B(n14347), .Z(n14338) );
  XNOR U22646 ( .A(n14330), .B(n14333), .Z(n14347) );
  NAND U22647 ( .A(n14348), .B(n14349), .Z(n14333) );
  NAND U22648 ( .A(n14350), .B(n14351), .Z(n14349) );
  OR U22649 ( .A(n14352), .B(n14353), .Z(n14350) );
  NANDN U22650 ( .A(n14354), .B(n14352), .Z(n14348) );
  IV U22651 ( .A(n14353), .Z(n14354) );
  NAND U22652 ( .A(n14355), .B(n14356), .Z(n14330) );
  NAND U22653 ( .A(n14357), .B(n14358), .Z(n14356) );
  NANDN U22654 ( .A(n14359), .B(n14360), .Z(n14357) );
  NANDN U22655 ( .A(n14360), .B(n14359), .Z(n14355) );
  AND U22656 ( .A(n14361), .B(n14362), .Z(n14332) );
  NAND U22657 ( .A(n14363), .B(n14364), .Z(n14362) );
  OR U22658 ( .A(n14365), .B(n14366), .Z(n14363) );
  NANDN U22659 ( .A(n14367), .B(n14365), .Z(n14361) );
  NAND U22660 ( .A(n14368), .B(n14369), .Z(n14336) );
  NANDN U22661 ( .A(n14370), .B(n14371), .Z(n14369) );
  OR U22662 ( .A(n14372), .B(n14373), .Z(n14371) );
  NANDN U22663 ( .A(n14374), .B(n14372), .Z(n14368) );
  IV U22664 ( .A(n14373), .Z(n14374) );
  XNOR U22665 ( .A(n14344), .B(n14375), .Z(n14339) );
  XNOR U22666 ( .A(n14342), .B(n14345), .Z(n14375) );
  NAND U22667 ( .A(n14376), .B(n14377), .Z(n14345) );
  NAND U22668 ( .A(n14378), .B(n14379), .Z(n14377) );
  OR U22669 ( .A(n14380), .B(n14381), .Z(n14378) );
  NANDN U22670 ( .A(n14382), .B(n14380), .Z(n14376) );
  IV U22671 ( .A(n14381), .Z(n14382) );
  NAND U22672 ( .A(n14383), .B(n14384), .Z(n14342) );
  NAND U22673 ( .A(n14385), .B(n14386), .Z(n14384) );
  NANDN U22674 ( .A(n14387), .B(n14388), .Z(n14385) );
  NANDN U22675 ( .A(n14388), .B(n14387), .Z(n14383) );
  AND U22676 ( .A(n14389), .B(n14390), .Z(n14344) );
  NAND U22677 ( .A(n14391), .B(n14392), .Z(n14390) );
  OR U22678 ( .A(n14393), .B(n14394), .Z(n14391) );
  NANDN U22679 ( .A(n14395), .B(n14393), .Z(n14389) );
  XNOR U22680 ( .A(n14370), .B(n14396), .Z(N64116) );
  XOR U22681 ( .A(n14372), .B(n14373), .Z(n14396) );
  XNOR U22682 ( .A(n14386), .B(n14397), .Z(n14373) );
  XOR U22683 ( .A(n14387), .B(n14388), .Z(n14397) );
  XOR U22684 ( .A(n14393), .B(n14398), .Z(n14388) );
  XOR U22685 ( .A(n14392), .B(n14395), .Z(n14398) );
  IV U22686 ( .A(n14394), .Z(n14395) );
  NAND U22687 ( .A(n14399), .B(n14400), .Z(n14394) );
  OR U22688 ( .A(n14401), .B(n14402), .Z(n14400) );
  OR U22689 ( .A(n14403), .B(n14404), .Z(n14399) );
  NAND U22690 ( .A(n14405), .B(n14406), .Z(n14392) );
  OR U22691 ( .A(n14407), .B(n14408), .Z(n14406) );
  OR U22692 ( .A(n14409), .B(n14410), .Z(n14405) );
  NOR U22693 ( .A(n14411), .B(n14412), .Z(n14393) );
  ANDN U22694 ( .B(n14413), .A(n14414), .Z(n14387) );
  XNOR U22695 ( .A(n14380), .B(n14415), .Z(n14386) );
  XNOR U22696 ( .A(n14379), .B(n14381), .Z(n14415) );
  NAND U22697 ( .A(n14416), .B(n14417), .Z(n14381) );
  OR U22698 ( .A(n14418), .B(n14419), .Z(n14417) );
  OR U22699 ( .A(n14420), .B(n14421), .Z(n14416) );
  NAND U22700 ( .A(n14422), .B(n14423), .Z(n14379) );
  OR U22701 ( .A(n14424), .B(n14425), .Z(n14423) );
  OR U22702 ( .A(n14426), .B(n14427), .Z(n14422) );
  ANDN U22703 ( .B(n14428), .A(n14429), .Z(n14380) );
  IV U22704 ( .A(n14430), .Z(n14428) );
  ANDN U22705 ( .B(n14431), .A(n14432), .Z(n14372) );
  XOR U22706 ( .A(n14358), .B(n14433), .Z(n14370) );
  XOR U22707 ( .A(n14359), .B(n14360), .Z(n14433) );
  XOR U22708 ( .A(n14365), .B(n14434), .Z(n14360) );
  XOR U22709 ( .A(n14364), .B(n14367), .Z(n14434) );
  IV U22710 ( .A(n14366), .Z(n14367) );
  NAND U22711 ( .A(n14435), .B(n14436), .Z(n14366) );
  OR U22712 ( .A(n14437), .B(n14438), .Z(n14436) );
  OR U22713 ( .A(n14439), .B(n14440), .Z(n14435) );
  NAND U22714 ( .A(n14441), .B(n14442), .Z(n14364) );
  OR U22715 ( .A(n14443), .B(n14444), .Z(n14442) );
  OR U22716 ( .A(n14445), .B(n14446), .Z(n14441) );
  NOR U22717 ( .A(n14447), .B(n14448), .Z(n14365) );
  ANDN U22718 ( .B(n14449), .A(n14450), .Z(n14359) );
  IV U22719 ( .A(n14451), .Z(n14449) );
  XNOR U22720 ( .A(n14352), .B(n14452), .Z(n14358) );
  XNOR U22721 ( .A(n14351), .B(n14353), .Z(n14452) );
  NAND U22722 ( .A(n14453), .B(n14454), .Z(n14353) );
  OR U22723 ( .A(n14455), .B(n14456), .Z(n14454) );
  OR U22724 ( .A(n14457), .B(n14458), .Z(n14453) );
  NAND U22725 ( .A(n14459), .B(n14460), .Z(n14351) );
  OR U22726 ( .A(n14461), .B(n14462), .Z(n14460) );
  OR U22727 ( .A(n14463), .B(n14464), .Z(n14459) );
  ANDN U22728 ( .B(n14465), .A(n14466), .Z(n14352) );
  IV U22729 ( .A(n14467), .Z(n14465) );
  XNOR U22730 ( .A(n14432), .B(n14431), .Z(N64115) );
  XOR U22731 ( .A(n14451), .B(n14450), .Z(n14431) );
  XNOR U22732 ( .A(n14466), .B(n14467), .Z(n14450) );
  XNOR U22733 ( .A(n14461), .B(n14462), .Z(n14467) );
  XNOR U22734 ( .A(n14463), .B(n14464), .Z(n14462) );
  XNOR U22735 ( .A(y[6517]), .B(x[6517]), .Z(n14464) );
  XNOR U22736 ( .A(y[6518]), .B(x[6518]), .Z(n14463) );
  XNOR U22737 ( .A(y[6516]), .B(x[6516]), .Z(n14461) );
  XNOR U22738 ( .A(n14455), .B(n14456), .Z(n14466) );
  XNOR U22739 ( .A(y[6513]), .B(x[6513]), .Z(n14456) );
  XNOR U22740 ( .A(n14457), .B(n14458), .Z(n14455) );
  XNOR U22741 ( .A(y[6514]), .B(x[6514]), .Z(n14458) );
  XNOR U22742 ( .A(y[6515]), .B(x[6515]), .Z(n14457) );
  XNOR U22743 ( .A(n14448), .B(n14447), .Z(n14451) );
  XNOR U22744 ( .A(n14443), .B(n14444), .Z(n14447) );
  XNOR U22745 ( .A(y[6510]), .B(x[6510]), .Z(n14444) );
  XNOR U22746 ( .A(n14445), .B(n14446), .Z(n14443) );
  XNOR U22747 ( .A(y[6511]), .B(x[6511]), .Z(n14446) );
  XNOR U22748 ( .A(y[6512]), .B(x[6512]), .Z(n14445) );
  XNOR U22749 ( .A(n14437), .B(n14438), .Z(n14448) );
  XNOR U22750 ( .A(y[6507]), .B(x[6507]), .Z(n14438) );
  XNOR U22751 ( .A(n14439), .B(n14440), .Z(n14437) );
  XNOR U22752 ( .A(y[6508]), .B(x[6508]), .Z(n14440) );
  XNOR U22753 ( .A(y[6509]), .B(x[6509]), .Z(n14439) );
  XOR U22754 ( .A(n14413), .B(n14414), .Z(n14432) );
  XNOR U22755 ( .A(n14429), .B(n14430), .Z(n14414) );
  XNOR U22756 ( .A(n14424), .B(n14425), .Z(n14430) );
  XNOR U22757 ( .A(n14426), .B(n14427), .Z(n14425) );
  XNOR U22758 ( .A(y[6505]), .B(x[6505]), .Z(n14427) );
  XNOR U22759 ( .A(y[6506]), .B(x[6506]), .Z(n14426) );
  XNOR U22760 ( .A(y[6504]), .B(x[6504]), .Z(n14424) );
  XNOR U22761 ( .A(n14418), .B(n14419), .Z(n14429) );
  XNOR U22762 ( .A(y[6501]), .B(x[6501]), .Z(n14419) );
  XNOR U22763 ( .A(n14420), .B(n14421), .Z(n14418) );
  XNOR U22764 ( .A(y[6502]), .B(x[6502]), .Z(n14421) );
  XNOR U22765 ( .A(y[6503]), .B(x[6503]), .Z(n14420) );
  XOR U22766 ( .A(n14412), .B(n14411), .Z(n14413) );
  XNOR U22767 ( .A(n14407), .B(n14408), .Z(n14411) );
  XNOR U22768 ( .A(y[6498]), .B(x[6498]), .Z(n14408) );
  XNOR U22769 ( .A(n14409), .B(n14410), .Z(n14407) );
  XNOR U22770 ( .A(y[6499]), .B(x[6499]), .Z(n14410) );
  XNOR U22771 ( .A(y[6500]), .B(x[6500]), .Z(n14409) );
  XNOR U22772 ( .A(n14401), .B(n14402), .Z(n14412) );
  XNOR U22773 ( .A(y[6495]), .B(x[6495]), .Z(n14402) );
  XNOR U22774 ( .A(n14403), .B(n14404), .Z(n14401) );
  XNOR U22775 ( .A(y[6496]), .B(x[6496]), .Z(n14404) );
  XNOR U22776 ( .A(y[6497]), .B(x[6497]), .Z(n14403) );
  NAND U22777 ( .A(n14468), .B(n14469), .Z(N64106) );
  NANDN U22778 ( .A(n14470), .B(n14471), .Z(n14469) );
  OR U22779 ( .A(n14472), .B(n14473), .Z(n14471) );
  NAND U22780 ( .A(n14472), .B(n14473), .Z(n14468) );
  XOR U22781 ( .A(n14472), .B(n14474), .Z(N64105) );
  XNOR U22782 ( .A(n14470), .B(n14473), .Z(n14474) );
  AND U22783 ( .A(n14475), .B(n14476), .Z(n14473) );
  NANDN U22784 ( .A(n14477), .B(n14478), .Z(n14476) );
  NANDN U22785 ( .A(n14479), .B(n14480), .Z(n14478) );
  NANDN U22786 ( .A(n14480), .B(n14479), .Z(n14475) );
  NAND U22787 ( .A(n14481), .B(n14482), .Z(n14470) );
  NANDN U22788 ( .A(n14483), .B(n14484), .Z(n14482) );
  OR U22789 ( .A(n14485), .B(n14486), .Z(n14484) );
  NAND U22790 ( .A(n14486), .B(n14485), .Z(n14481) );
  AND U22791 ( .A(n14487), .B(n14488), .Z(n14472) );
  NANDN U22792 ( .A(n14489), .B(n14490), .Z(n14488) );
  NANDN U22793 ( .A(n14491), .B(n14492), .Z(n14490) );
  NANDN U22794 ( .A(n14492), .B(n14491), .Z(n14487) );
  XOR U22795 ( .A(n14486), .B(n14493), .Z(N64104) );
  XOR U22796 ( .A(n14483), .B(n14485), .Z(n14493) );
  XNOR U22797 ( .A(n14479), .B(n14494), .Z(n14485) );
  XNOR U22798 ( .A(n14477), .B(n14480), .Z(n14494) );
  NAND U22799 ( .A(n14495), .B(n14496), .Z(n14480) );
  NAND U22800 ( .A(n14497), .B(n14498), .Z(n14496) );
  OR U22801 ( .A(n14499), .B(n14500), .Z(n14497) );
  NANDN U22802 ( .A(n14501), .B(n14499), .Z(n14495) );
  IV U22803 ( .A(n14500), .Z(n14501) );
  NAND U22804 ( .A(n14502), .B(n14503), .Z(n14477) );
  NAND U22805 ( .A(n14504), .B(n14505), .Z(n14503) );
  NANDN U22806 ( .A(n14506), .B(n14507), .Z(n14504) );
  NANDN U22807 ( .A(n14507), .B(n14506), .Z(n14502) );
  AND U22808 ( .A(n14508), .B(n14509), .Z(n14479) );
  NAND U22809 ( .A(n14510), .B(n14511), .Z(n14509) );
  OR U22810 ( .A(n14512), .B(n14513), .Z(n14510) );
  NANDN U22811 ( .A(n14514), .B(n14512), .Z(n14508) );
  NAND U22812 ( .A(n14515), .B(n14516), .Z(n14483) );
  NANDN U22813 ( .A(n14517), .B(n14518), .Z(n14516) );
  OR U22814 ( .A(n14519), .B(n14520), .Z(n14518) );
  NANDN U22815 ( .A(n14521), .B(n14519), .Z(n14515) );
  IV U22816 ( .A(n14520), .Z(n14521) );
  XNOR U22817 ( .A(n14491), .B(n14522), .Z(n14486) );
  XNOR U22818 ( .A(n14489), .B(n14492), .Z(n14522) );
  NAND U22819 ( .A(n14523), .B(n14524), .Z(n14492) );
  NAND U22820 ( .A(n14525), .B(n14526), .Z(n14524) );
  OR U22821 ( .A(n14527), .B(n14528), .Z(n14525) );
  NANDN U22822 ( .A(n14529), .B(n14527), .Z(n14523) );
  IV U22823 ( .A(n14528), .Z(n14529) );
  NAND U22824 ( .A(n14530), .B(n14531), .Z(n14489) );
  NAND U22825 ( .A(n14532), .B(n14533), .Z(n14531) );
  NANDN U22826 ( .A(n14534), .B(n14535), .Z(n14532) );
  NANDN U22827 ( .A(n14535), .B(n14534), .Z(n14530) );
  AND U22828 ( .A(n14536), .B(n14537), .Z(n14491) );
  NAND U22829 ( .A(n14538), .B(n14539), .Z(n14537) );
  OR U22830 ( .A(n14540), .B(n14541), .Z(n14538) );
  NANDN U22831 ( .A(n14542), .B(n14540), .Z(n14536) );
  XNOR U22832 ( .A(n14517), .B(n14543), .Z(N64103) );
  XOR U22833 ( .A(n14519), .B(n14520), .Z(n14543) );
  XNOR U22834 ( .A(n14533), .B(n14544), .Z(n14520) );
  XOR U22835 ( .A(n14534), .B(n14535), .Z(n14544) );
  XOR U22836 ( .A(n14540), .B(n14545), .Z(n14535) );
  XOR U22837 ( .A(n14539), .B(n14542), .Z(n14545) );
  IV U22838 ( .A(n14541), .Z(n14542) );
  NAND U22839 ( .A(n14546), .B(n14547), .Z(n14541) );
  OR U22840 ( .A(n14548), .B(n14549), .Z(n14547) );
  OR U22841 ( .A(n14550), .B(n14551), .Z(n14546) );
  NAND U22842 ( .A(n14552), .B(n14553), .Z(n14539) );
  OR U22843 ( .A(n14554), .B(n14555), .Z(n14553) );
  OR U22844 ( .A(n14556), .B(n14557), .Z(n14552) );
  NOR U22845 ( .A(n14558), .B(n14559), .Z(n14540) );
  ANDN U22846 ( .B(n14560), .A(n14561), .Z(n14534) );
  XNOR U22847 ( .A(n14527), .B(n14562), .Z(n14533) );
  XNOR U22848 ( .A(n14526), .B(n14528), .Z(n14562) );
  NAND U22849 ( .A(n14563), .B(n14564), .Z(n14528) );
  OR U22850 ( .A(n14565), .B(n14566), .Z(n14564) );
  OR U22851 ( .A(n14567), .B(n14568), .Z(n14563) );
  NAND U22852 ( .A(n14569), .B(n14570), .Z(n14526) );
  OR U22853 ( .A(n14571), .B(n14572), .Z(n14570) );
  OR U22854 ( .A(n14573), .B(n14574), .Z(n14569) );
  ANDN U22855 ( .B(n14575), .A(n14576), .Z(n14527) );
  IV U22856 ( .A(n14577), .Z(n14575) );
  ANDN U22857 ( .B(n14578), .A(n14579), .Z(n14519) );
  XOR U22858 ( .A(n14505), .B(n14580), .Z(n14517) );
  XOR U22859 ( .A(n14506), .B(n14507), .Z(n14580) );
  XOR U22860 ( .A(n14512), .B(n14581), .Z(n14507) );
  XOR U22861 ( .A(n14511), .B(n14514), .Z(n14581) );
  IV U22862 ( .A(n14513), .Z(n14514) );
  NAND U22863 ( .A(n14582), .B(n14583), .Z(n14513) );
  OR U22864 ( .A(n14584), .B(n14585), .Z(n14583) );
  OR U22865 ( .A(n14586), .B(n14587), .Z(n14582) );
  NAND U22866 ( .A(n14588), .B(n14589), .Z(n14511) );
  OR U22867 ( .A(n14590), .B(n14591), .Z(n14589) );
  OR U22868 ( .A(n14592), .B(n14593), .Z(n14588) );
  NOR U22869 ( .A(n14594), .B(n14595), .Z(n14512) );
  ANDN U22870 ( .B(n14596), .A(n14597), .Z(n14506) );
  IV U22871 ( .A(n14598), .Z(n14596) );
  XNOR U22872 ( .A(n14499), .B(n14599), .Z(n14505) );
  XNOR U22873 ( .A(n14498), .B(n14500), .Z(n14599) );
  NAND U22874 ( .A(n14600), .B(n14601), .Z(n14500) );
  OR U22875 ( .A(n14602), .B(n14603), .Z(n14601) );
  OR U22876 ( .A(n14604), .B(n14605), .Z(n14600) );
  NAND U22877 ( .A(n14606), .B(n14607), .Z(n14498) );
  OR U22878 ( .A(n14608), .B(n14609), .Z(n14607) );
  OR U22879 ( .A(n14610), .B(n14611), .Z(n14606) );
  ANDN U22880 ( .B(n14612), .A(n14613), .Z(n14499) );
  IV U22881 ( .A(n14614), .Z(n14612) );
  XNOR U22882 ( .A(n14579), .B(n14578), .Z(N64102) );
  XOR U22883 ( .A(n14598), .B(n14597), .Z(n14578) );
  XNOR U22884 ( .A(n14613), .B(n14614), .Z(n14597) );
  XNOR U22885 ( .A(n14608), .B(n14609), .Z(n14614) );
  XNOR U22886 ( .A(n14610), .B(n14611), .Z(n14609) );
  XNOR U22887 ( .A(y[6493]), .B(x[6493]), .Z(n14611) );
  XNOR U22888 ( .A(y[6494]), .B(x[6494]), .Z(n14610) );
  XNOR U22889 ( .A(y[6492]), .B(x[6492]), .Z(n14608) );
  XNOR U22890 ( .A(n14602), .B(n14603), .Z(n14613) );
  XNOR U22891 ( .A(y[6489]), .B(x[6489]), .Z(n14603) );
  XNOR U22892 ( .A(n14604), .B(n14605), .Z(n14602) );
  XNOR U22893 ( .A(y[6490]), .B(x[6490]), .Z(n14605) );
  XNOR U22894 ( .A(y[6491]), .B(x[6491]), .Z(n14604) );
  XNOR U22895 ( .A(n14595), .B(n14594), .Z(n14598) );
  XNOR U22896 ( .A(n14590), .B(n14591), .Z(n14594) );
  XNOR U22897 ( .A(y[6486]), .B(x[6486]), .Z(n14591) );
  XNOR U22898 ( .A(n14592), .B(n14593), .Z(n14590) );
  XNOR U22899 ( .A(y[6487]), .B(x[6487]), .Z(n14593) );
  XNOR U22900 ( .A(y[6488]), .B(x[6488]), .Z(n14592) );
  XNOR U22901 ( .A(n14584), .B(n14585), .Z(n14595) );
  XNOR U22902 ( .A(y[6483]), .B(x[6483]), .Z(n14585) );
  XNOR U22903 ( .A(n14586), .B(n14587), .Z(n14584) );
  XNOR U22904 ( .A(y[6484]), .B(x[6484]), .Z(n14587) );
  XNOR U22905 ( .A(y[6485]), .B(x[6485]), .Z(n14586) );
  XOR U22906 ( .A(n14560), .B(n14561), .Z(n14579) );
  XNOR U22907 ( .A(n14576), .B(n14577), .Z(n14561) );
  XNOR U22908 ( .A(n14571), .B(n14572), .Z(n14577) );
  XNOR U22909 ( .A(n14573), .B(n14574), .Z(n14572) );
  XNOR U22910 ( .A(y[6481]), .B(x[6481]), .Z(n14574) );
  XNOR U22911 ( .A(y[6482]), .B(x[6482]), .Z(n14573) );
  XNOR U22912 ( .A(y[6480]), .B(x[6480]), .Z(n14571) );
  XNOR U22913 ( .A(n14565), .B(n14566), .Z(n14576) );
  XNOR U22914 ( .A(y[6477]), .B(x[6477]), .Z(n14566) );
  XNOR U22915 ( .A(n14567), .B(n14568), .Z(n14565) );
  XNOR U22916 ( .A(y[6478]), .B(x[6478]), .Z(n14568) );
  XNOR U22917 ( .A(y[6479]), .B(x[6479]), .Z(n14567) );
  XOR U22918 ( .A(n14559), .B(n14558), .Z(n14560) );
  XNOR U22919 ( .A(n14554), .B(n14555), .Z(n14558) );
  XNOR U22920 ( .A(y[6474]), .B(x[6474]), .Z(n14555) );
  XNOR U22921 ( .A(n14556), .B(n14557), .Z(n14554) );
  XNOR U22922 ( .A(y[6475]), .B(x[6475]), .Z(n14557) );
  XNOR U22923 ( .A(y[6476]), .B(x[6476]), .Z(n14556) );
  XNOR U22924 ( .A(n14548), .B(n14549), .Z(n14559) );
  XNOR U22925 ( .A(y[6471]), .B(x[6471]), .Z(n14549) );
  XNOR U22926 ( .A(n14550), .B(n14551), .Z(n14548) );
  XNOR U22927 ( .A(y[6472]), .B(x[6472]), .Z(n14551) );
  XNOR U22928 ( .A(y[6473]), .B(x[6473]), .Z(n14550) );
  NAND U22929 ( .A(n14615), .B(n14616), .Z(N64093) );
  NANDN U22930 ( .A(n14617), .B(n14618), .Z(n14616) );
  OR U22931 ( .A(n14619), .B(n14620), .Z(n14618) );
  NAND U22932 ( .A(n14619), .B(n14620), .Z(n14615) );
  XOR U22933 ( .A(n14619), .B(n14621), .Z(N64092) );
  XNOR U22934 ( .A(n14617), .B(n14620), .Z(n14621) );
  AND U22935 ( .A(n14622), .B(n14623), .Z(n14620) );
  NANDN U22936 ( .A(n14624), .B(n14625), .Z(n14623) );
  NANDN U22937 ( .A(n14626), .B(n14627), .Z(n14625) );
  NANDN U22938 ( .A(n14627), .B(n14626), .Z(n14622) );
  NAND U22939 ( .A(n14628), .B(n14629), .Z(n14617) );
  NANDN U22940 ( .A(n14630), .B(n14631), .Z(n14629) );
  OR U22941 ( .A(n14632), .B(n14633), .Z(n14631) );
  NAND U22942 ( .A(n14633), .B(n14632), .Z(n14628) );
  AND U22943 ( .A(n14634), .B(n14635), .Z(n14619) );
  NANDN U22944 ( .A(n14636), .B(n14637), .Z(n14635) );
  NANDN U22945 ( .A(n14638), .B(n14639), .Z(n14637) );
  NANDN U22946 ( .A(n14639), .B(n14638), .Z(n14634) );
  XOR U22947 ( .A(n14633), .B(n14640), .Z(N64091) );
  XOR U22948 ( .A(n14630), .B(n14632), .Z(n14640) );
  XNOR U22949 ( .A(n14626), .B(n14641), .Z(n14632) );
  XNOR U22950 ( .A(n14624), .B(n14627), .Z(n14641) );
  NAND U22951 ( .A(n14642), .B(n14643), .Z(n14627) );
  NAND U22952 ( .A(n14644), .B(n14645), .Z(n14643) );
  OR U22953 ( .A(n14646), .B(n14647), .Z(n14644) );
  NANDN U22954 ( .A(n14648), .B(n14646), .Z(n14642) );
  IV U22955 ( .A(n14647), .Z(n14648) );
  NAND U22956 ( .A(n14649), .B(n14650), .Z(n14624) );
  NAND U22957 ( .A(n14651), .B(n14652), .Z(n14650) );
  NANDN U22958 ( .A(n14653), .B(n14654), .Z(n14651) );
  NANDN U22959 ( .A(n14654), .B(n14653), .Z(n14649) );
  AND U22960 ( .A(n14655), .B(n14656), .Z(n14626) );
  NAND U22961 ( .A(n14657), .B(n14658), .Z(n14656) );
  OR U22962 ( .A(n14659), .B(n14660), .Z(n14657) );
  NANDN U22963 ( .A(n14661), .B(n14659), .Z(n14655) );
  NAND U22964 ( .A(n14662), .B(n14663), .Z(n14630) );
  NANDN U22965 ( .A(n14664), .B(n14665), .Z(n14663) );
  OR U22966 ( .A(n14666), .B(n14667), .Z(n14665) );
  NANDN U22967 ( .A(n14668), .B(n14666), .Z(n14662) );
  IV U22968 ( .A(n14667), .Z(n14668) );
  XNOR U22969 ( .A(n14638), .B(n14669), .Z(n14633) );
  XNOR U22970 ( .A(n14636), .B(n14639), .Z(n14669) );
  NAND U22971 ( .A(n14670), .B(n14671), .Z(n14639) );
  NAND U22972 ( .A(n14672), .B(n14673), .Z(n14671) );
  OR U22973 ( .A(n14674), .B(n14675), .Z(n14672) );
  NANDN U22974 ( .A(n14676), .B(n14674), .Z(n14670) );
  IV U22975 ( .A(n14675), .Z(n14676) );
  NAND U22976 ( .A(n14677), .B(n14678), .Z(n14636) );
  NAND U22977 ( .A(n14679), .B(n14680), .Z(n14678) );
  NANDN U22978 ( .A(n14681), .B(n14682), .Z(n14679) );
  NANDN U22979 ( .A(n14682), .B(n14681), .Z(n14677) );
  AND U22980 ( .A(n14683), .B(n14684), .Z(n14638) );
  NAND U22981 ( .A(n14685), .B(n14686), .Z(n14684) );
  OR U22982 ( .A(n14687), .B(n14688), .Z(n14685) );
  NANDN U22983 ( .A(n14689), .B(n14687), .Z(n14683) );
  XNOR U22984 ( .A(n14664), .B(n14690), .Z(N64090) );
  XOR U22985 ( .A(n14666), .B(n14667), .Z(n14690) );
  XNOR U22986 ( .A(n14680), .B(n14691), .Z(n14667) );
  XOR U22987 ( .A(n14681), .B(n14682), .Z(n14691) );
  XOR U22988 ( .A(n14687), .B(n14692), .Z(n14682) );
  XOR U22989 ( .A(n14686), .B(n14689), .Z(n14692) );
  IV U22990 ( .A(n14688), .Z(n14689) );
  NAND U22991 ( .A(n14693), .B(n14694), .Z(n14688) );
  OR U22992 ( .A(n14695), .B(n14696), .Z(n14694) );
  OR U22993 ( .A(n14697), .B(n14698), .Z(n14693) );
  NAND U22994 ( .A(n14699), .B(n14700), .Z(n14686) );
  OR U22995 ( .A(n14701), .B(n14702), .Z(n14700) );
  OR U22996 ( .A(n14703), .B(n14704), .Z(n14699) );
  NOR U22997 ( .A(n14705), .B(n14706), .Z(n14687) );
  ANDN U22998 ( .B(n14707), .A(n14708), .Z(n14681) );
  XNOR U22999 ( .A(n14674), .B(n14709), .Z(n14680) );
  XNOR U23000 ( .A(n14673), .B(n14675), .Z(n14709) );
  NAND U23001 ( .A(n14710), .B(n14711), .Z(n14675) );
  OR U23002 ( .A(n14712), .B(n14713), .Z(n14711) );
  OR U23003 ( .A(n14714), .B(n14715), .Z(n14710) );
  NAND U23004 ( .A(n14716), .B(n14717), .Z(n14673) );
  OR U23005 ( .A(n14718), .B(n14719), .Z(n14717) );
  OR U23006 ( .A(n14720), .B(n14721), .Z(n14716) );
  ANDN U23007 ( .B(n14722), .A(n14723), .Z(n14674) );
  IV U23008 ( .A(n14724), .Z(n14722) );
  ANDN U23009 ( .B(n14725), .A(n14726), .Z(n14666) );
  XOR U23010 ( .A(n14652), .B(n14727), .Z(n14664) );
  XOR U23011 ( .A(n14653), .B(n14654), .Z(n14727) );
  XOR U23012 ( .A(n14659), .B(n14728), .Z(n14654) );
  XOR U23013 ( .A(n14658), .B(n14661), .Z(n14728) );
  IV U23014 ( .A(n14660), .Z(n14661) );
  NAND U23015 ( .A(n14729), .B(n14730), .Z(n14660) );
  OR U23016 ( .A(n14731), .B(n14732), .Z(n14730) );
  OR U23017 ( .A(n14733), .B(n14734), .Z(n14729) );
  NAND U23018 ( .A(n14735), .B(n14736), .Z(n14658) );
  OR U23019 ( .A(n14737), .B(n14738), .Z(n14736) );
  OR U23020 ( .A(n14739), .B(n14740), .Z(n14735) );
  NOR U23021 ( .A(n14741), .B(n14742), .Z(n14659) );
  ANDN U23022 ( .B(n14743), .A(n14744), .Z(n14653) );
  IV U23023 ( .A(n14745), .Z(n14743) );
  XNOR U23024 ( .A(n14646), .B(n14746), .Z(n14652) );
  XNOR U23025 ( .A(n14645), .B(n14647), .Z(n14746) );
  NAND U23026 ( .A(n14747), .B(n14748), .Z(n14647) );
  OR U23027 ( .A(n14749), .B(n14750), .Z(n14748) );
  OR U23028 ( .A(n14751), .B(n14752), .Z(n14747) );
  NAND U23029 ( .A(n14753), .B(n14754), .Z(n14645) );
  OR U23030 ( .A(n14755), .B(n14756), .Z(n14754) );
  OR U23031 ( .A(n14757), .B(n14758), .Z(n14753) );
  ANDN U23032 ( .B(n14759), .A(n14760), .Z(n14646) );
  IV U23033 ( .A(n14761), .Z(n14759) );
  XNOR U23034 ( .A(n14726), .B(n14725), .Z(N64089) );
  XOR U23035 ( .A(n14745), .B(n14744), .Z(n14725) );
  XNOR U23036 ( .A(n14760), .B(n14761), .Z(n14744) );
  XNOR U23037 ( .A(n14755), .B(n14756), .Z(n14761) );
  XNOR U23038 ( .A(n14757), .B(n14758), .Z(n14756) );
  XNOR U23039 ( .A(y[6469]), .B(x[6469]), .Z(n14758) );
  XNOR U23040 ( .A(y[6470]), .B(x[6470]), .Z(n14757) );
  XNOR U23041 ( .A(y[6468]), .B(x[6468]), .Z(n14755) );
  XNOR U23042 ( .A(n14749), .B(n14750), .Z(n14760) );
  XNOR U23043 ( .A(y[6465]), .B(x[6465]), .Z(n14750) );
  XNOR U23044 ( .A(n14751), .B(n14752), .Z(n14749) );
  XNOR U23045 ( .A(y[6466]), .B(x[6466]), .Z(n14752) );
  XNOR U23046 ( .A(y[6467]), .B(x[6467]), .Z(n14751) );
  XNOR U23047 ( .A(n14742), .B(n14741), .Z(n14745) );
  XNOR U23048 ( .A(n14737), .B(n14738), .Z(n14741) );
  XNOR U23049 ( .A(y[6462]), .B(x[6462]), .Z(n14738) );
  XNOR U23050 ( .A(n14739), .B(n14740), .Z(n14737) );
  XNOR U23051 ( .A(y[6463]), .B(x[6463]), .Z(n14740) );
  XNOR U23052 ( .A(y[6464]), .B(x[6464]), .Z(n14739) );
  XNOR U23053 ( .A(n14731), .B(n14732), .Z(n14742) );
  XNOR U23054 ( .A(y[6459]), .B(x[6459]), .Z(n14732) );
  XNOR U23055 ( .A(n14733), .B(n14734), .Z(n14731) );
  XNOR U23056 ( .A(y[6460]), .B(x[6460]), .Z(n14734) );
  XNOR U23057 ( .A(y[6461]), .B(x[6461]), .Z(n14733) );
  XOR U23058 ( .A(n14707), .B(n14708), .Z(n14726) );
  XNOR U23059 ( .A(n14723), .B(n14724), .Z(n14708) );
  XNOR U23060 ( .A(n14718), .B(n14719), .Z(n14724) );
  XNOR U23061 ( .A(n14720), .B(n14721), .Z(n14719) );
  XNOR U23062 ( .A(y[6457]), .B(x[6457]), .Z(n14721) );
  XNOR U23063 ( .A(y[6458]), .B(x[6458]), .Z(n14720) );
  XNOR U23064 ( .A(y[6456]), .B(x[6456]), .Z(n14718) );
  XNOR U23065 ( .A(n14712), .B(n14713), .Z(n14723) );
  XNOR U23066 ( .A(y[6453]), .B(x[6453]), .Z(n14713) );
  XNOR U23067 ( .A(n14714), .B(n14715), .Z(n14712) );
  XNOR U23068 ( .A(y[6454]), .B(x[6454]), .Z(n14715) );
  XNOR U23069 ( .A(y[6455]), .B(x[6455]), .Z(n14714) );
  XOR U23070 ( .A(n14706), .B(n14705), .Z(n14707) );
  XNOR U23071 ( .A(n14701), .B(n14702), .Z(n14705) );
  XNOR U23072 ( .A(y[6450]), .B(x[6450]), .Z(n14702) );
  XNOR U23073 ( .A(n14703), .B(n14704), .Z(n14701) );
  XNOR U23074 ( .A(y[6451]), .B(x[6451]), .Z(n14704) );
  XNOR U23075 ( .A(y[6452]), .B(x[6452]), .Z(n14703) );
  XNOR U23076 ( .A(n14695), .B(n14696), .Z(n14706) );
  XNOR U23077 ( .A(y[6447]), .B(x[6447]), .Z(n14696) );
  XNOR U23078 ( .A(n14697), .B(n14698), .Z(n14695) );
  XNOR U23079 ( .A(y[6448]), .B(x[6448]), .Z(n14698) );
  XNOR U23080 ( .A(y[6449]), .B(x[6449]), .Z(n14697) );
  NAND U23081 ( .A(n14762), .B(n14763), .Z(N64080) );
  NANDN U23082 ( .A(n14764), .B(n14765), .Z(n14763) );
  OR U23083 ( .A(n14766), .B(n14767), .Z(n14765) );
  NAND U23084 ( .A(n14766), .B(n14767), .Z(n14762) );
  XOR U23085 ( .A(n14766), .B(n14768), .Z(N64079) );
  XNOR U23086 ( .A(n14764), .B(n14767), .Z(n14768) );
  AND U23087 ( .A(n14769), .B(n14770), .Z(n14767) );
  NANDN U23088 ( .A(n14771), .B(n14772), .Z(n14770) );
  NANDN U23089 ( .A(n14773), .B(n14774), .Z(n14772) );
  NANDN U23090 ( .A(n14774), .B(n14773), .Z(n14769) );
  NAND U23091 ( .A(n14775), .B(n14776), .Z(n14764) );
  NANDN U23092 ( .A(n14777), .B(n14778), .Z(n14776) );
  OR U23093 ( .A(n14779), .B(n14780), .Z(n14778) );
  NAND U23094 ( .A(n14780), .B(n14779), .Z(n14775) );
  AND U23095 ( .A(n14781), .B(n14782), .Z(n14766) );
  NANDN U23096 ( .A(n14783), .B(n14784), .Z(n14782) );
  NANDN U23097 ( .A(n14785), .B(n14786), .Z(n14784) );
  NANDN U23098 ( .A(n14786), .B(n14785), .Z(n14781) );
  XOR U23099 ( .A(n14780), .B(n14787), .Z(N64078) );
  XOR U23100 ( .A(n14777), .B(n14779), .Z(n14787) );
  XNOR U23101 ( .A(n14773), .B(n14788), .Z(n14779) );
  XNOR U23102 ( .A(n14771), .B(n14774), .Z(n14788) );
  NAND U23103 ( .A(n14789), .B(n14790), .Z(n14774) );
  NAND U23104 ( .A(n14791), .B(n14792), .Z(n14790) );
  OR U23105 ( .A(n14793), .B(n14794), .Z(n14791) );
  NANDN U23106 ( .A(n14795), .B(n14793), .Z(n14789) );
  IV U23107 ( .A(n14794), .Z(n14795) );
  NAND U23108 ( .A(n14796), .B(n14797), .Z(n14771) );
  NAND U23109 ( .A(n14798), .B(n14799), .Z(n14797) );
  NANDN U23110 ( .A(n14800), .B(n14801), .Z(n14798) );
  NANDN U23111 ( .A(n14801), .B(n14800), .Z(n14796) );
  AND U23112 ( .A(n14802), .B(n14803), .Z(n14773) );
  NAND U23113 ( .A(n14804), .B(n14805), .Z(n14803) );
  OR U23114 ( .A(n14806), .B(n14807), .Z(n14804) );
  NANDN U23115 ( .A(n14808), .B(n14806), .Z(n14802) );
  NAND U23116 ( .A(n14809), .B(n14810), .Z(n14777) );
  NANDN U23117 ( .A(n14811), .B(n14812), .Z(n14810) );
  OR U23118 ( .A(n14813), .B(n14814), .Z(n14812) );
  NANDN U23119 ( .A(n14815), .B(n14813), .Z(n14809) );
  IV U23120 ( .A(n14814), .Z(n14815) );
  XNOR U23121 ( .A(n14785), .B(n14816), .Z(n14780) );
  XNOR U23122 ( .A(n14783), .B(n14786), .Z(n14816) );
  NAND U23123 ( .A(n14817), .B(n14818), .Z(n14786) );
  NAND U23124 ( .A(n14819), .B(n14820), .Z(n14818) );
  OR U23125 ( .A(n14821), .B(n14822), .Z(n14819) );
  NANDN U23126 ( .A(n14823), .B(n14821), .Z(n14817) );
  IV U23127 ( .A(n14822), .Z(n14823) );
  NAND U23128 ( .A(n14824), .B(n14825), .Z(n14783) );
  NAND U23129 ( .A(n14826), .B(n14827), .Z(n14825) );
  NANDN U23130 ( .A(n14828), .B(n14829), .Z(n14826) );
  NANDN U23131 ( .A(n14829), .B(n14828), .Z(n14824) );
  AND U23132 ( .A(n14830), .B(n14831), .Z(n14785) );
  NAND U23133 ( .A(n14832), .B(n14833), .Z(n14831) );
  OR U23134 ( .A(n14834), .B(n14835), .Z(n14832) );
  NANDN U23135 ( .A(n14836), .B(n14834), .Z(n14830) );
  XNOR U23136 ( .A(n14811), .B(n14837), .Z(N64077) );
  XOR U23137 ( .A(n14813), .B(n14814), .Z(n14837) );
  XNOR U23138 ( .A(n14827), .B(n14838), .Z(n14814) );
  XOR U23139 ( .A(n14828), .B(n14829), .Z(n14838) );
  XOR U23140 ( .A(n14834), .B(n14839), .Z(n14829) );
  XOR U23141 ( .A(n14833), .B(n14836), .Z(n14839) );
  IV U23142 ( .A(n14835), .Z(n14836) );
  NAND U23143 ( .A(n14840), .B(n14841), .Z(n14835) );
  OR U23144 ( .A(n14842), .B(n14843), .Z(n14841) );
  OR U23145 ( .A(n14844), .B(n14845), .Z(n14840) );
  NAND U23146 ( .A(n14846), .B(n14847), .Z(n14833) );
  OR U23147 ( .A(n14848), .B(n14849), .Z(n14847) );
  OR U23148 ( .A(n14850), .B(n14851), .Z(n14846) );
  NOR U23149 ( .A(n14852), .B(n14853), .Z(n14834) );
  ANDN U23150 ( .B(n14854), .A(n14855), .Z(n14828) );
  XNOR U23151 ( .A(n14821), .B(n14856), .Z(n14827) );
  XNOR U23152 ( .A(n14820), .B(n14822), .Z(n14856) );
  NAND U23153 ( .A(n14857), .B(n14858), .Z(n14822) );
  OR U23154 ( .A(n14859), .B(n14860), .Z(n14858) );
  OR U23155 ( .A(n14861), .B(n14862), .Z(n14857) );
  NAND U23156 ( .A(n14863), .B(n14864), .Z(n14820) );
  OR U23157 ( .A(n14865), .B(n14866), .Z(n14864) );
  OR U23158 ( .A(n14867), .B(n14868), .Z(n14863) );
  ANDN U23159 ( .B(n14869), .A(n14870), .Z(n14821) );
  IV U23160 ( .A(n14871), .Z(n14869) );
  ANDN U23161 ( .B(n14872), .A(n14873), .Z(n14813) );
  XOR U23162 ( .A(n14799), .B(n14874), .Z(n14811) );
  XOR U23163 ( .A(n14800), .B(n14801), .Z(n14874) );
  XOR U23164 ( .A(n14806), .B(n14875), .Z(n14801) );
  XOR U23165 ( .A(n14805), .B(n14808), .Z(n14875) );
  IV U23166 ( .A(n14807), .Z(n14808) );
  NAND U23167 ( .A(n14876), .B(n14877), .Z(n14807) );
  OR U23168 ( .A(n14878), .B(n14879), .Z(n14877) );
  OR U23169 ( .A(n14880), .B(n14881), .Z(n14876) );
  NAND U23170 ( .A(n14882), .B(n14883), .Z(n14805) );
  OR U23171 ( .A(n14884), .B(n14885), .Z(n14883) );
  OR U23172 ( .A(n14886), .B(n14887), .Z(n14882) );
  NOR U23173 ( .A(n14888), .B(n14889), .Z(n14806) );
  ANDN U23174 ( .B(n14890), .A(n14891), .Z(n14800) );
  IV U23175 ( .A(n14892), .Z(n14890) );
  XNOR U23176 ( .A(n14793), .B(n14893), .Z(n14799) );
  XNOR U23177 ( .A(n14792), .B(n14794), .Z(n14893) );
  NAND U23178 ( .A(n14894), .B(n14895), .Z(n14794) );
  OR U23179 ( .A(n14896), .B(n14897), .Z(n14895) );
  OR U23180 ( .A(n14898), .B(n14899), .Z(n14894) );
  NAND U23181 ( .A(n14900), .B(n14901), .Z(n14792) );
  OR U23182 ( .A(n14902), .B(n14903), .Z(n14901) );
  OR U23183 ( .A(n14904), .B(n14905), .Z(n14900) );
  ANDN U23184 ( .B(n14906), .A(n14907), .Z(n14793) );
  IV U23185 ( .A(n14908), .Z(n14906) );
  XNOR U23186 ( .A(n14873), .B(n14872), .Z(N64076) );
  XOR U23187 ( .A(n14892), .B(n14891), .Z(n14872) );
  XNOR U23188 ( .A(n14907), .B(n14908), .Z(n14891) );
  XNOR U23189 ( .A(n14902), .B(n14903), .Z(n14908) );
  XNOR U23190 ( .A(n14904), .B(n14905), .Z(n14903) );
  XNOR U23191 ( .A(y[6445]), .B(x[6445]), .Z(n14905) );
  XNOR U23192 ( .A(y[6446]), .B(x[6446]), .Z(n14904) );
  XNOR U23193 ( .A(y[6444]), .B(x[6444]), .Z(n14902) );
  XNOR U23194 ( .A(n14896), .B(n14897), .Z(n14907) );
  XNOR U23195 ( .A(y[6441]), .B(x[6441]), .Z(n14897) );
  XNOR U23196 ( .A(n14898), .B(n14899), .Z(n14896) );
  XNOR U23197 ( .A(y[6442]), .B(x[6442]), .Z(n14899) );
  XNOR U23198 ( .A(y[6443]), .B(x[6443]), .Z(n14898) );
  XNOR U23199 ( .A(n14889), .B(n14888), .Z(n14892) );
  XNOR U23200 ( .A(n14884), .B(n14885), .Z(n14888) );
  XNOR U23201 ( .A(y[6438]), .B(x[6438]), .Z(n14885) );
  XNOR U23202 ( .A(n14886), .B(n14887), .Z(n14884) );
  XNOR U23203 ( .A(y[6439]), .B(x[6439]), .Z(n14887) );
  XNOR U23204 ( .A(y[6440]), .B(x[6440]), .Z(n14886) );
  XNOR U23205 ( .A(n14878), .B(n14879), .Z(n14889) );
  XNOR U23206 ( .A(y[6435]), .B(x[6435]), .Z(n14879) );
  XNOR U23207 ( .A(n14880), .B(n14881), .Z(n14878) );
  XNOR U23208 ( .A(y[6436]), .B(x[6436]), .Z(n14881) );
  XNOR U23209 ( .A(y[6437]), .B(x[6437]), .Z(n14880) );
  XOR U23210 ( .A(n14854), .B(n14855), .Z(n14873) );
  XNOR U23211 ( .A(n14870), .B(n14871), .Z(n14855) );
  XNOR U23212 ( .A(n14865), .B(n14866), .Z(n14871) );
  XNOR U23213 ( .A(n14867), .B(n14868), .Z(n14866) );
  XNOR U23214 ( .A(y[6433]), .B(x[6433]), .Z(n14868) );
  XNOR U23215 ( .A(y[6434]), .B(x[6434]), .Z(n14867) );
  XNOR U23216 ( .A(y[6432]), .B(x[6432]), .Z(n14865) );
  XNOR U23217 ( .A(n14859), .B(n14860), .Z(n14870) );
  XNOR U23218 ( .A(y[6429]), .B(x[6429]), .Z(n14860) );
  XNOR U23219 ( .A(n14861), .B(n14862), .Z(n14859) );
  XNOR U23220 ( .A(y[6430]), .B(x[6430]), .Z(n14862) );
  XNOR U23221 ( .A(y[6431]), .B(x[6431]), .Z(n14861) );
  XOR U23222 ( .A(n14853), .B(n14852), .Z(n14854) );
  XNOR U23223 ( .A(n14848), .B(n14849), .Z(n14852) );
  XNOR U23224 ( .A(y[6426]), .B(x[6426]), .Z(n14849) );
  XNOR U23225 ( .A(n14850), .B(n14851), .Z(n14848) );
  XNOR U23226 ( .A(y[6427]), .B(x[6427]), .Z(n14851) );
  XNOR U23227 ( .A(y[6428]), .B(x[6428]), .Z(n14850) );
  XNOR U23228 ( .A(n14842), .B(n14843), .Z(n14853) );
  XNOR U23229 ( .A(y[6423]), .B(x[6423]), .Z(n14843) );
  XNOR U23230 ( .A(n14844), .B(n14845), .Z(n14842) );
  XNOR U23231 ( .A(y[6424]), .B(x[6424]), .Z(n14845) );
  XNOR U23232 ( .A(y[6425]), .B(x[6425]), .Z(n14844) );
  NAND U23233 ( .A(n14909), .B(n14910), .Z(N64067) );
  NANDN U23234 ( .A(n14911), .B(n14912), .Z(n14910) );
  OR U23235 ( .A(n14913), .B(n14914), .Z(n14912) );
  NAND U23236 ( .A(n14913), .B(n14914), .Z(n14909) );
  XOR U23237 ( .A(n14913), .B(n14915), .Z(N64066) );
  XNOR U23238 ( .A(n14911), .B(n14914), .Z(n14915) );
  AND U23239 ( .A(n14916), .B(n14917), .Z(n14914) );
  NANDN U23240 ( .A(n14918), .B(n14919), .Z(n14917) );
  NANDN U23241 ( .A(n14920), .B(n14921), .Z(n14919) );
  NANDN U23242 ( .A(n14921), .B(n14920), .Z(n14916) );
  NAND U23243 ( .A(n14922), .B(n14923), .Z(n14911) );
  NANDN U23244 ( .A(n14924), .B(n14925), .Z(n14923) );
  OR U23245 ( .A(n14926), .B(n14927), .Z(n14925) );
  NAND U23246 ( .A(n14927), .B(n14926), .Z(n14922) );
  AND U23247 ( .A(n14928), .B(n14929), .Z(n14913) );
  NANDN U23248 ( .A(n14930), .B(n14931), .Z(n14929) );
  NANDN U23249 ( .A(n14932), .B(n14933), .Z(n14931) );
  NANDN U23250 ( .A(n14933), .B(n14932), .Z(n14928) );
  XOR U23251 ( .A(n14927), .B(n14934), .Z(N64065) );
  XOR U23252 ( .A(n14924), .B(n14926), .Z(n14934) );
  XNOR U23253 ( .A(n14920), .B(n14935), .Z(n14926) );
  XNOR U23254 ( .A(n14918), .B(n14921), .Z(n14935) );
  NAND U23255 ( .A(n14936), .B(n14937), .Z(n14921) );
  NAND U23256 ( .A(n14938), .B(n14939), .Z(n14937) );
  OR U23257 ( .A(n14940), .B(n14941), .Z(n14938) );
  NANDN U23258 ( .A(n14942), .B(n14940), .Z(n14936) );
  IV U23259 ( .A(n14941), .Z(n14942) );
  NAND U23260 ( .A(n14943), .B(n14944), .Z(n14918) );
  NAND U23261 ( .A(n14945), .B(n14946), .Z(n14944) );
  NANDN U23262 ( .A(n14947), .B(n14948), .Z(n14945) );
  NANDN U23263 ( .A(n14948), .B(n14947), .Z(n14943) );
  AND U23264 ( .A(n14949), .B(n14950), .Z(n14920) );
  NAND U23265 ( .A(n14951), .B(n14952), .Z(n14950) );
  OR U23266 ( .A(n14953), .B(n14954), .Z(n14951) );
  NANDN U23267 ( .A(n14955), .B(n14953), .Z(n14949) );
  NAND U23268 ( .A(n14956), .B(n14957), .Z(n14924) );
  NANDN U23269 ( .A(n14958), .B(n14959), .Z(n14957) );
  OR U23270 ( .A(n14960), .B(n14961), .Z(n14959) );
  NANDN U23271 ( .A(n14962), .B(n14960), .Z(n14956) );
  IV U23272 ( .A(n14961), .Z(n14962) );
  XNOR U23273 ( .A(n14932), .B(n14963), .Z(n14927) );
  XNOR U23274 ( .A(n14930), .B(n14933), .Z(n14963) );
  NAND U23275 ( .A(n14964), .B(n14965), .Z(n14933) );
  NAND U23276 ( .A(n14966), .B(n14967), .Z(n14965) );
  OR U23277 ( .A(n14968), .B(n14969), .Z(n14966) );
  NANDN U23278 ( .A(n14970), .B(n14968), .Z(n14964) );
  IV U23279 ( .A(n14969), .Z(n14970) );
  NAND U23280 ( .A(n14971), .B(n14972), .Z(n14930) );
  NAND U23281 ( .A(n14973), .B(n14974), .Z(n14972) );
  NANDN U23282 ( .A(n14975), .B(n14976), .Z(n14973) );
  NANDN U23283 ( .A(n14976), .B(n14975), .Z(n14971) );
  AND U23284 ( .A(n14977), .B(n14978), .Z(n14932) );
  NAND U23285 ( .A(n14979), .B(n14980), .Z(n14978) );
  OR U23286 ( .A(n14981), .B(n14982), .Z(n14979) );
  NANDN U23287 ( .A(n14983), .B(n14981), .Z(n14977) );
  XNOR U23288 ( .A(n14958), .B(n14984), .Z(N64064) );
  XOR U23289 ( .A(n14960), .B(n14961), .Z(n14984) );
  XNOR U23290 ( .A(n14974), .B(n14985), .Z(n14961) );
  XOR U23291 ( .A(n14975), .B(n14976), .Z(n14985) );
  XOR U23292 ( .A(n14981), .B(n14986), .Z(n14976) );
  XOR U23293 ( .A(n14980), .B(n14983), .Z(n14986) );
  IV U23294 ( .A(n14982), .Z(n14983) );
  NAND U23295 ( .A(n14987), .B(n14988), .Z(n14982) );
  OR U23296 ( .A(n14989), .B(n14990), .Z(n14988) );
  OR U23297 ( .A(n14991), .B(n14992), .Z(n14987) );
  NAND U23298 ( .A(n14993), .B(n14994), .Z(n14980) );
  OR U23299 ( .A(n14995), .B(n14996), .Z(n14994) );
  OR U23300 ( .A(n14997), .B(n14998), .Z(n14993) );
  NOR U23301 ( .A(n14999), .B(n15000), .Z(n14981) );
  ANDN U23302 ( .B(n15001), .A(n15002), .Z(n14975) );
  XNOR U23303 ( .A(n14968), .B(n15003), .Z(n14974) );
  XNOR U23304 ( .A(n14967), .B(n14969), .Z(n15003) );
  NAND U23305 ( .A(n15004), .B(n15005), .Z(n14969) );
  OR U23306 ( .A(n15006), .B(n15007), .Z(n15005) );
  OR U23307 ( .A(n15008), .B(n15009), .Z(n15004) );
  NAND U23308 ( .A(n15010), .B(n15011), .Z(n14967) );
  OR U23309 ( .A(n15012), .B(n15013), .Z(n15011) );
  OR U23310 ( .A(n15014), .B(n15015), .Z(n15010) );
  ANDN U23311 ( .B(n15016), .A(n15017), .Z(n14968) );
  IV U23312 ( .A(n15018), .Z(n15016) );
  ANDN U23313 ( .B(n15019), .A(n15020), .Z(n14960) );
  XOR U23314 ( .A(n14946), .B(n15021), .Z(n14958) );
  XOR U23315 ( .A(n14947), .B(n14948), .Z(n15021) );
  XOR U23316 ( .A(n14953), .B(n15022), .Z(n14948) );
  XOR U23317 ( .A(n14952), .B(n14955), .Z(n15022) );
  IV U23318 ( .A(n14954), .Z(n14955) );
  NAND U23319 ( .A(n15023), .B(n15024), .Z(n14954) );
  OR U23320 ( .A(n15025), .B(n15026), .Z(n15024) );
  OR U23321 ( .A(n15027), .B(n15028), .Z(n15023) );
  NAND U23322 ( .A(n15029), .B(n15030), .Z(n14952) );
  OR U23323 ( .A(n15031), .B(n15032), .Z(n15030) );
  OR U23324 ( .A(n15033), .B(n15034), .Z(n15029) );
  NOR U23325 ( .A(n15035), .B(n15036), .Z(n14953) );
  ANDN U23326 ( .B(n15037), .A(n15038), .Z(n14947) );
  IV U23327 ( .A(n15039), .Z(n15037) );
  XNOR U23328 ( .A(n14940), .B(n15040), .Z(n14946) );
  XNOR U23329 ( .A(n14939), .B(n14941), .Z(n15040) );
  NAND U23330 ( .A(n15041), .B(n15042), .Z(n14941) );
  OR U23331 ( .A(n15043), .B(n15044), .Z(n15042) );
  OR U23332 ( .A(n15045), .B(n15046), .Z(n15041) );
  NAND U23333 ( .A(n15047), .B(n15048), .Z(n14939) );
  OR U23334 ( .A(n15049), .B(n15050), .Z(n15048) );
  OR U23335 ( .A(n15051), .B(n15052), .Z(n15047) );
  ANDN U23336 ( .B(n15053), .A(n15054), .Z(n14940) );
  IV U23337 ( .A(n15055), .Z(n15053) );
  XNOR U23338 ( .A(n15020), .B(n15019), .Z(N64063) );
  XOR U23339 ( .A(n15039), .B(n15038), .Z(n15019) );
  XNOR U23340 ( .A(n15054), .B(n15055), .Z(n15038) );
  XNOR U23341 ( .A(n15049), .B(n15050), .Z(n15055) );
  XNOR U23342 ( .A(n15051), .B(n15052), .Z(n15050) );
  XNOR U23343 ( .A(y[6421]), .B(x[6421]), .Z(n15052) );
  XNOR U23344 ( .A(y[6422]), .B(x[6422]), .Z(n15051) );
  XNOR U23345 ( .A(y[6420]), .B(x[6420]), .Z(n15049) );
  XNOR U23346 ( .A(n15043), .B(n15044), .Z(n15054) );
  XNOR U23347 ( .A(y[6417]), .B(x[6417]), .Z(n15044) );
  XNOR U23348 ( .A(n15045), .B(n15046), .Z(n15043) );
  XNOR U23349 ( .A(y[6418]), .B(x[6418]), .Z(n15046) );
  XNOR U23350 ( .A(y[6419]), .B(x[6419]), .Z(n15045) );
  XNOR U23351 ( .A(n15036), .B(n15035), .Z(n15039) );
  XNOR U23352 ( .A(n15031), .B(n15032), .Z(n15035) );
  XNOR U23353 ( .A(y[6414]), .B(x[6414]), .Z(n15032) );
  XNOR U23354 ( .A(n15033), .B(n15034), .Z(n15031) );
  XNOR U23355 ( .A(y[6415]), .B(x[6415]), .Z(n15034) );
  XNOR U23356 ( .A(y[6416]), .B(x[6416]), .Z(n15033) );
  XNOR U23357 ( .A(n15025), .B(n15026), .Z(n15036) );
  XNOR U23358 ( .A(y[6411]), .B(x[6411]), .Z(n15026) );
  XNOR U23359 ( .A(n15027), .B(n15028), .Z(n15025) );
  XNOR U23360 ( .A(y[6412]), .B(x[6412]), .Z(n15028) );
  XNOR U23361 ( .A(y[6413]), .B(x[6413]), .Z(n15027) );
  XOR U23362 ( .A(n15001), .B(n15002), .Z(n15020) );
  XNOR U23363 ( .A(n15017), .B(n15018), .Z(n15002) );
  XNOR U23364 ( .A(n15012), .B(n15013), .Z(n15018) );
  XNOR U23365 ( .A(n15014), .B(n15015), .Z(n15013) );
  XNOR U23366 ( .A(y[6409]), .B(x[6409]), .Z(n15015) );
  XNOR U23367 ( .A(y[6410]), .B(x[6410]), .Z(n15014) );
  XNOR U23368 ( .A(y[6408]), .B(x[6408]), .Z(n15012) );
  XNOR U23369 ( .A(n15006), .B(n15007), .Z(n15017) );
  XNOR U23370 ( .A(y[6405]), .B(x[6405]), .Z(n15007) );
  XNOR U23371 ( .A(n15008), .B(n15009), .Z(n15006) );
  XNOR U23372 ( .A(y[6406]), .B(x[6406]), .Z(n15009) );
  XNOR U23373 ( .A(y[6407]), .B(x[6407]), .Z(n15008) );
  XOR U23374 ( .A(n15000), .B(n14999), .Z(n15001) );
  XNOR U23375 ( .A(n14995), .B(n14996), .Z(n14999) );
  XNOR U23376 ( .A(y[6402]), .B(x[6402]), .Z(n14996) );
  XNOR U23377 ( .A(n14997), .B(n14998), .Z(n14995) );
  XNOR U23378 ( .A(y[6403]), .B(x[6403]), .Z(n14998) );
  XNOR U23379 ( .A(y[6404]), .B(x[6404]), .Z(n14997) );
  XNOR U23380 ( .A(n14989), .B(n14990), .Z(n15000) );
  XNOR U23381 ( .A(y[6399]), .B(x[6399]), .Z(n14990) );
  XNOR U23382 ( .A(n14991), .B(n14992), .Z(n14989) );
  XNOR U23383 ( .A(y[6400]), .B(x[6400]), .Z(n14992) );
  XNOR U23384 ( .A(y[6401]), .B(x[6401]), .Z(n14991) );
  NAND U23385 ( .A(n15056), .B(n15057), .Z(N64054) );
  NANDN U23386 ( .A(n15058), .B(n15059), .Z(n15057) );
  OR U23387 ( .A(n15060), .B(n15061), .Z(n15059) );
  NAND U23388 ( .A(n15060), .B(n15061), .Z(n15056) );
  XOR U23389 ( .A(n15060), .B(n15062), .Z(N64053) );
  XNOR U23390 ( .A(n15058), .B(n15061), .Z(n15062) );
  AND U23391 ( .A(n15063), .B(n15064), .Z(n15061) );
  NANDN U23392 ( .A(n15065), .B(n15066), .Z(n15064) );
  NANDN U23393 ( .A(n15067), .B(n15068), .Z(n15066) );
  NANDN U23394 ( .A(n15068), .B(n15067), .Z(n15063) );
  NAND U23395 ( .A(n15069), .B(n15070), .Z(n15058) );
  NANDN U23396 ( .A(n15071), .B(n15072), .Z(n15070) );
  OR U23397 ( .A(n15073), .B(n15074), .Z(n15072) );
  NAND U23398 ( .A(n15074), .B(n15073), .Z(n15069) );
  AND U23399 ( .A(n15075), .B(n15076), .Z(n15060) );
  NANDN U23400 ( .A(n15077), .B(n15078), .Z(n15076) );
  NANDN U23401 ( .A(n15079), .B(n15080), .Z(n15078) );
  NANDN U23402 ( .A(n15080), .B(n15079), .Z(n15075) );
  XOR U23403 ( .A(n15074), .B(n15081), .Z(N64052) );
  XOR U23404 ( .A(n15071), .B(n15073), .Z(n15081) );
  XNOR U23405 ( .A(n15067), .B(n15082), .Z(n15073) );
  XNOR U23406 ( .A(n15065), .B(n15068), .Z(n15082) );
  NAND U23407 ( .A(n15083), .B(n15084), .Z(n15068) );
  NAND U23408 ( .A(n15085), .B(n15086), .Z(n15084) );
  OR U23409 ( .A(n15087), .B(n15088), .Z(n15085) );
  NANDN U23410 ( .A(n15089), .B(n15087), .Z(n15083) );
  IV U23411 ( .A(n15088), .Z(n15089) );
  NAND U23412 ( .A(n15090), .B(n15091), .Z(n15065) );
  NAND U23413 ( .A(n15092), .B(n15093), .Z(n15091) );
  NANDN U23414 ( .A(n15094), .B(n15095), .Z(n15092) );
  NANDN U23415 ( .A(n15095), .B(n15094), .Z(n15090) );
  AND U23416 ( .A(n15096), .B(n15097), .Z(n15067) );
  NAND U23417 ( .A(n15098), .B(n15099), .Z(n15097) );
  OR U23418 ( .A(n15100), .B(n15101), .Z(n15098) );
  NANDN U23419 ( .A(n15102), .B(n15100), .Z(n15096) );
  NAND U23420 ( .A(n15103), .B(n15104), .Z(n15071) );
  NANDN U23421 ( .A(n15105), .B(n15106), .Z(n15104) );
  OR U23422 ( .A(n15107), .B(n15108), .Z(n15106) );
  NANDN U23423 ( .A(n15109), .B(n15107), .Z(n15103) );
  IV U23424 ( .A(n15108), .Z(n15109) );
  XNOR U23425 ( .A(n15079), .B(n15110), .Z(n15074) );
  XNOR U23426 ( .A(n15077), .B(n15080), .Z(n15110) );
  NAND U23427 ( .A(n15111), .B(n15112), .Z(n15080) );
  NAND U23428 ( .A(n15113), .B(n15114), .Z(n15112) );
  OR U23429 ( .A(n15115), .B(n15116), .Z(n15113) );
  NANDN U23430 ( .A(n15117), .B(n15115), .Z(n15111) );
  IV U23431 ( .A(n15116), .Z(n15117) );
  NAND U23432 ( .A(n15118), .B(n15119), .Z(n15077) );
  NAND U23433 ( .A(n15120), .B(n15121), .Z(n15119) );
  NANDN U23434 ( .A(n15122), .B(n15123), .Z(n15120) );
  NANDN U23435 ( .A(n15123), .B(n15122), .Z(n15118) );
  AND U23436 ( .A(n15124), .B(n15125), .Z(n15079) );
  NAND U23437 ( .A(n15126), .B(n15127), .Z(n15125) );
  OR U23438 ( .A(n15128), .B(n15129), .Z(n15126) );
  NANDN U23439 ( .A(n15130), .B(n15128), .Z(n15124) );
  XNOR U23440 ( .A(n15105), .B(n15131), .Z(N64051) );
  XOR U23441 ( .A(n15107), .B(n15108), .Z(n15131) );
  XNOR U23442 ( .A(n15121), .B(n15132), .Z(n15108) );
  XOR U23443 ( .A(n15122), .B(n15123), .Z(n15132) );
  XOR U23444 ( .A(n15128), .B(n15133), .Z(n15123) );
  XOR U23445 ( .A(n15127), .B(n15130), .Z(n15133) );
  IV U23446 ( .A(n15129), .Z(n15130) );
  NAND U23447 ( .A(n15134), .B(n15135), .Z(n15129) );
  OR U23448 ( .A(n15136), .B(n15137), .Z(n15135) );
  OR U23449 ( .A(n15138), .B(n15139), .Z(n15134) );
  NAND U23450 ( .A(n15140), .B(n15141), .Z(n15127) );
  OR U23451 ( .A(n15142), .B(n15143), .Z(n15141) );
  OR U23452 ( .A(n15144), .B(n15145), .Z(n15140) );
  NOR U23453 ( .A(n15146), .B(n15147), .Z(n15128) );
  ANDN U23454 ( .B(n15148), .A(n15149), .Z(n15122) );
  XNOR U23455 ( .A(n15115), .B(n15150), .Z(n15121) );
  XNOR U23456 ( .A(n15114), .B(n15116), .Z(n15150) );
  NAND U23457 ( .A(n15151), .B(n15152), .Z(n15116) );
  OR U23458 ( .A(n15153), .B(n15154), .Z(n15152) );
  OR U23459 ( .A(n15155), .B(n15156), .Z(n15151) );
  NAND U23460 ( .A(n15157), .B(n15158), .Z(n15114) );
  OR U23461 ( .A(n15159), .B(n15160), .Z(n15158) );
  OR U23462 ( .A(n15161), .B(n15162), .Z(n15157) );
  ANDN U23463 ( .B(n15163), .A(n15164), .Z(n15115) );
  IV U23464 ( .A(n15165), .Z(n15163) );
  ANDN U23465 ( .B(n15166), .A(n15167), .Z(n15107) );
  XOR U23466 ( .A(n15093), .B(n15168), .Z(n15105) );
  XOR U23467 ( .A(n15094), .B(n15095), .Z(n15168) );
  XOR U23468 ( .A(n15100), .B(n15169), .Z(n15095) );
  XOR U23469 ( .A(n15099), .B(n15102), .Z(n15169) );
  IV U23470 ( .A(n15101), .Z(n15102) );
  NAND U23471 ( .A(n15170), .B(n15171), .Z(n15101) );
  OR U23472 ( .A(n15172), .B(n15173), .Z(n15171) );
  OR U23473 ( .A(n15174), .B(n15175), .Z(n15170) );
  NAND U23474 ( .A(n15176), .B(n15177), .Z(n15099) );
  OR U23475 ( .A(n15178), .B(n15179), .Z(n15177) );
  OR U23476 ( .A(n15180), .B(n15181), .Z(n15176) );
  NOR U23477 ( .A(n15182), .B(n15183), .Z(n15100) );
  ANDN U23478 ( .B(n15184), .A(n15185), .Z(n15094) );
  IV U23479 ( .A(n15186), .Z(n15184) );
  XNOR U23480 ( .A(n15087), .B(n15187), .Z(n15093) );
  XNOR U23481 ( .A(n15086), .B(n15088), .Z(n15187) );
  NAND U23482 ( .A(n15188), .B(n15189), .Z(n15088) );
  OR U23483 ( .A(n15190), .B(n15191), .Z(n15189) );
  OR U23484 ( .A(n15192), .B(n15193), .Z(n15188) );
  NAND U23485 ( .A(n15194), .B(n15195), .Z(n15086) );
  OR U23486 ( .A(n15196), .B(n15197), .Z(n15195) );
  OR U23487 ( .A(n15198), .B(n15199), .Z(n15194) );
  ANDN U23488 ( .B(n15200), .A(n15201), .Z(n15087) );
  IV U23489 ( .A(n15202), .Z(n15200) );
  XNOR U23490 ( .A(n15167), .B(n15166), .Z(N64050) );
  XOR U23491 ( .A(n15186), .B(n15185), .Z(n15166) );
  XNOR U23492 ( .A(n15201), .B(n15202), .Z(n15185) );
  XNOR U23493 ( .A(n15196), .B(n15197), .Z(n15202) );
  XNOR U23494 ( .A(n15198), .B(n15199), .Z(n15197) );
  XNOR U23495 ( .A(y[6397]), .B(x[6397]), .Z(n15199) );
  XNOR U23496 ( .A(y[6398]), .B(x[6398]), .Z(n15198) );
  XNOR U23497 ( .A(y[6396]), .B(x[6396]), .Z(n15196) );
  XNOR U23498 ( .A(n15190), .B(n15191), .Z(n15201) );
  XNOR U23499 ( .A(y[6393]), .B(x[6393]), .Z(n15191) );
  XNOR U23500 ( .A(n15192), .B(n15193), .Z(n15190) );
  XNOR U23501 ( .A(y[6394]), .B(x[6394]), .Z(n15193) );
  XNOR U23502 ( .A(y[6395]), .B(x[6395]), .Z(n15192) );
  XNOR U23503 ( .A(n15183), .B(n15182), .Z(n15186) );
  XNOR U23504 ( .A(n15178), .B(n15179), .Z(n15182) );
  XNOR U23505 ( .A(y[6390]), .B(x[6390]), .Z(n15179) );
  XNOR U23506 ( .A(n15180), .B(n15181), .Z(n15178) );
  XNOR U23507 ( .A(y[6391]), .B(x[6391]), .Z(n15181) );
  XNOR U23508 ( .A(y[6392]), .B(x[6392]), .Z(n15180) );
  XNOR U23509 ( .A(n15172), .B(n15173), .Z(n15183) );
  XNOR U23510 ( .A(y[6387]), .B(x[6387]), .Z(n15173) );
  XNOR U23511 ( .A(n15174), .B(n15175), .Z(n15172) );
  XNOR U23512 ( .A(y[6388]), .B(x[6388]), .Z(n15175) );
  XNOR U23513 ( .A(y[6389]), .B(x[6389]), .Z(n15174) );
  XOR U23514 ( .A(n15148), .B(n15149), .Z(n15167) );
  XNOR U23515 ( .A(n15164), .B(n15165), .Z(n15149) );
  XNOR U23516 ( .A(n15159), .B(n15160), .Z(n15165) );
  XNOR U23517 ( .A(n15161), .B(n15162), .Z(n15160) );
  XNOR U23518 ( .A(y[6385]), .B(x[6385]), .Z(n15162) );
  XNOR U23519 ( .A(y[6386]), .B(x[6386]), .Z(n15161) );
  XNOR U23520 ( .A(y[6384]), .B(x[6384]), .Z(n15159) );
  XNOR U23521 ( .A(n15153), .B(n15154), .Z(n15164) );
  XNOR U23522 ( .A(y[6381]), .B(x[6381]), .Z(n15154) );
  XNOR U23523 ( .A(n15155), .B(n15156), .Z(n15153) );
  XNOR U23524 ( .A(y[6382]), .B(x[6382]), .Z(n15156) );
  XNOR U23525 ( .A(y[6383]), .B(x[6383]), .Z(n15155) );
  XOR U23526 ( .A(n15147), .B(n15146), .Z(n15148) );
  XNOR U23527 ( .A(n15142), .B(n15143), .Z(n15146) );
  XNOR U23528 ( .A(y[6378]), .B(x[6378]), .Z(n15143) );
  XNOR U23529 ( .A(n15144), .B(n15145), .Z(n15142) );
  XNOR U23530 ( .A(y[6379]), .B(x[6379]), .Z(n15145) );
  XNOR U23531 ( .A(y[6380]), .B(x[6380]), .Z(n15144) );
  XNOR U23532 ( .A(n15136), .B(n15137), .Z(n15147) );
  XNOR U23533 ( .A(y[6375]), .B(x[6375]), .Z(n15137) );
  XNOR U23534 ( .A(n15138), .B(n15139), .Z(n15136) );
  XNOR U23535 ( .A(y[6376]), .B(x[6376]), .Z(n15139) );
  XNOR U23536 ( .A(y[6377]), .B(x[6377]), .Z(n15138) );
  NAND U23537 ( .A(n15203), .B(n15204), .Z(N64041) );
  NANDN U23538 ( .A(n15205), .B(n15206), .Z(n15204) );
  OR U23539 ( .A(n15207), .B(n15208), .Z(n15206) );
  NAND U23540 ( .A(n15207), .B(n15208), .Z(n15203) );
  XOR U23541 ( .A(n15207), .B(n15209), .Z(N64040) );
  XNOR U23542 ( .A(n15205), .B(n15208), .Z(n15209) );
  AND U23543 ( .A(n15210), .B(n15211), .Z(n15208) );
  NANDN U23544 ( .A(n15212), .B(n15213), .Z(n15211) );
  NANDN U23545 ( .A(n15214), .B(n15215), .Z(n15213) );
  NANDN U23546 ( .A(n15215), .B(n15214), .Z(n15210) );
  NAND U23547 ( .A(n15216), .B(n15217), .Z(n15205) );
  NANDN U23548 ( .A(n15218), .B(n15219), .Z(n15217) );
  OR U23549 ( .A(n15220), .B(n15221), .Z(n15219) );
  NAND U23550 ( .A(n15221), .B(n15220), .Z(n15216) );
  AND U23551 ( .A(n15222), .B(n15223), .Z(n15207) );
  NANDN U23552 ( .A(n15224), .B(n15225), .Z(n15223) );
  NANDN U23553 ( .A(n15226), .B(n15227), .Z(n15225) );
  NANDN U23554 ( .A(n15227), .B(n15226), .Z(n15222) );
  XOR U23555 ( .A(n15221), .B(n15228), .Z(N64039) );
  XOR U23556 ( .A(n15218), .B(n15220), .Z(n15228) );
  XNOR U23557 ( .A(n15214), .B(n15229), .Z(n15220) );
  XNOR U23558 ( .A(n15212), .B(n15215), .Z(n15229) );
  NAND U23559 ( .A(n15230), .B(n15231), .Z(n15215) );
  NAND U23560 ( .A(n15232), .B(n15233), .Z(n15231) );
  OR U23561 ( .A(n15234), .B(n15235), .Z(n15232) );
  NANDN U23562 ( .A(n15236), .B(n15234), .Z(n15230) );
  IV U23563 ( .A(n15235), .Z(n15236) );
  NAND U23564 ( .A(n15237), .B(n15238), .Z(n15212) );
  NAND U23565 ( .A(n15239), .B(n15240), .Z(n15238) );
  NANDN U23566 ( .A(n15241), .B(n15242), .Z(n15239) );
  NANDN U23567 ( .A(n15242), .B(n15241), .Z(n15237) );
  AND U23568 ( .A(n15243), .B(n15244), .Z(n15214) );
  NAND U23569 ( .A(n15245), .B(n15246), .Z(n15244) );
  OR U23570 ( .A(n15247), .B(n15248), .Z(n15245) );
  NANDN U23571 ( .A(n15249), .B(n15247), .Z(n15243) );
  NAND U23572 ( .A(n15250), .B(n15251), .Z(n15218) );
  NANDN U23573 ( .A(n15252), .B(n15253), .Z(n15251) );
  OR U23574 ( .A(n15254), .B(n15255), .Z(n15253) );
  NANDN U23575 ( .A(n15256), .B(n15254), .Z(n15250) );
  IV U23576 ( .A(n15255), .Z(n15256) );
  XNOR U23577 ( .A(n15226), .B(n15257), .Z(n15221) );
  XNOR U23578 ( .A(n15224), .B(n15227), .Z(n15257) );
  NAND U23579 ( .A(n15258), .B(n15259), .Z(n15227) );
  NAND U23580 ( .A(n15260), .B(n15261), .Z(n15259) );
  OR U23581 ( .A(n15262), .B(n15263), .Z(n15260) );
  NANDN U23582 ( .A(n15264), .B(n15262), .Z(n15258) );
  IV U23583 ( .A(n15263), .Z(n15264) );
  NAND U23584 ( .A(n15265), .B(n15266), .Z(n15224) );
  NAND U23585 ( .A(n15267), .B(n15268), .Z(n15266) );
  NANDN U23586 ( .A(n15269), .B(n15270), .Z(n15267) );
  NANDN U23587 ( .A(n15270), .B(n15269), .Z(n15265) );
  AND U23588 ( .A(n15271), .B(n15272), .Z(n15226) );
  NAND U23589 ( .A(n15273), .B(n15274), .Z(n15272) );
  OR U23590 ( .A(n15275), .B(n15276), .Z(n15273) );
  NANDN U23591 ( .A(n15277), .B(n15275), .Z(n15271) );
  XNOR U23592 ( .A(n15252), .B(n15278), .Z(N64038) );
  XOR U23593 ( .A(n15254), .B(n15255), .Z(n15278) );
  XNOR U23594 ( .A(n15268), .B(n15279), .Z(n15255) );
  XOR U23595 ( .A(n15269), .B(n15270), .Z(n15279) );
  XOR U23596 ( .A(n15275), .B(n15280), .Z(n15270) );
  XOR U23597 ( .A(n15274), .B(n15277), .Z(n15280) );
  IV U23598 ( .A(n15276), .Z(n15277) );
  NAND U23599 ( .A(n15281), .B(n15282), .Z(n15276) );
  OR U23600 ( .A(n15283), .B(n15284), .Z(n15282) );
  OR U23601 ( .A(n15285), .B(n15286), .Z(n15281) );
  NAND U23602 ( .A(n15287), .B(n15288), .Z(n15274) );
  OR U23603 ( .A(n15289), .B(n15290), .Z(n15288) );
  OR U23604 ( .A(n15291), .B(n15292), .Z(n15287) );
  NOR U23605 ( .A(n15293), .B(n15294), .Z(n15275) );
  ANDN U23606 ( .B(n15295), .A(n15296), .Z(n15269) );
  XNOR U23607 ( .A(n15262), .B(n15297), .Z(n15268) );
  XNOR U23608 ( .A(n15261), .B(n15263), .Z(n15297) );
  NAND U23609 ( .A(n15298), .B(n15299), .Z(n15263) );
  OR U23610 ( .A(n15300), .B(n15301), .Z(n15299) );
  OR U23611 ( .A(n15302), .B(n15303), .Z(n15298) );
  NAND U23612 ( .A(n15304), .B(n15305), .Z(n15261) );
  OR U23613 ( .A(n15306), .B(n15307), .Z(n15305) );
  OR U23614 ( .A(n15308), .B(n15309), .Z(n15304) );
  ANDN U23615 ( .B(n15310), .A(n15311), .Z(n15262) );
  IV U23616 ( .A(n15312), .Z(n15310) );
  ANDN U23617 ( .B(n15313), .A(n15314), .Z(n15254) );
  XOR U23618 ( .A(n15240), .B(n15315), .Z(n15252) );
  XOR U23619 ( .A(n15241), .B(n15242), .Z(n15315) );
  XOR U23620 ( .A(n15247), .B(n15316), .Z(n15242) );
  XOR U23621 ( .A(n15246), .B(n15249), .Z(n15316) );
  IV U23622 ( .A(n15248), .Z(n15249) );
  NAND U23623 ( .A(n15317), .B(n15318), .Z(n15248) );
  OR U23624 ( .A(n15319), .B(n15320), .Z(n15318) );
  OR U23625 ( .A(n15321), .B(n15322), .Z(n15317) );
  NAND U23626 ( .A(n15323), .B(n15324), .Z(n15246) );
  OR U23627 ( .A(n15325), .B(n15326), .Z(n15324) );
  OR U23628 ( .A(n15327), .B(n15328), .Z(n15323) );
  NOR U23629 ( .A(n15329), .B(n15330), .Z(n15247) );
  ANDN U23630 ( .B(n15331), .A(n15332), .Z(n15241) );
  IV U23631 ( .A(n15333), .Z(n15331) );
  XNOR U23632 ( .A(n15234), .B(n15334), .Z(n15240) );
  XNOR U23633 ( .A(n15233), .B(n15235), .Z(n15334) );
  NAND U23634 ( .A(n15335), .B(n15336), .Z(n15235) );
  OR U23635 ( .A(n15337), .B(n15338), .Z(n15336) );
  OR U23636 ( .A(n15339), .B(n15340), .Z(n15335) );
  NAND U23637 ( .A(n15341), .B(n15342), .Z(n15233) );
  OR U23638 ( .A(n15343), .B(n15344), .Z(n15342) );
  OR U23639 ( .A(n15345), .B(n15346), .Z(n15341) );
  ANDN U23640 ( .B(n15347), .A(n15348), .Z(n15234) );
  IV U23641 ( .A(n15349), .Z(n15347) );
  XNOR U23642 ( .A(n15314), .B(n15313), .Z(N64037) );
  XOR U23643 ( .A(n15333), .B(n15332), .Z(n15313) );
  XNOR U23644 ( .A(n15348), .B(n15349), .Z(n15332) );
  XNOR U23645 ( .A(n15343), .B(n15344), .Z(n15349) );
  XNOR U23646 ( .A(n15345), .B(n15346), .Z(n15344) );
  XNOR U23647 ( .A(y[6373]), .B(x[6373]), .Z(n15346) );
  XNOR U23648 ( .A(y[6374]), .B(x[6374]), .Z(n15345) );
  XNOR U23649 ( .A(y[6372]), .B(x[6372]), .Z(n15343) );
  XNOR U23650 ( .A(n15337), .B(n15338), .Z(n15348) );
  XNOR U23651 ( .A(y[6369]), .B(x[6369]), .Z(n15338) );
  XNOR U23652 ( .A(n15339), .B(n15340), .Z(n15337) );
  XNOR U23653 ( .A(y[6370]), .B(x[6370]), .Z(n15340) );
  XNOR U23654 ( .A(y[6371]), .B(x[6371]), .Z(n15339) );
  XNOR U23655 ( .A(n15330), .B(n15329), .Z(n15333) );
  XNOR U23656 ( .A(n15325), .B(n15326), .Z(n15329) );
  XNOR U23657 ( .A(y[6366]), .B(x[6366]), .Z(n15326) );
  XNOR U23658 ( .A(n15327), .B(n15328), .Z(n15325) );
  XNOR U23659 ( .A(y[6367]), .B(x[6367]), .Z(n15328) );
  XNOR U23660 ( .A(y[6368]), .B(x[6368]), .Z(n15327) );
  XNOR U23661 ( .A(n15319), .B(n15320), .Z(n15330) );
  XNOR U23662 ( .A(y[6363]), .B(x[6363]), .Z(n15320) );
  XNOR U23663 ( .A(n15321), .B(n15322), .Z(n15319) );
  XNOR U23664 ( .A(y[6364]), .B(x[6364]), .Z(n15322) );
  XNOR U23665 ( .A(y[6365]), .B(x[6365]), .Z(n15321) );
  XOR U23666 ( .A(n15295), .B(n15296), .Z(n15314) );
  XNOR U23667 ( .A(n15311), .B(n15312), .Z(n15296) );
  XNOR U23668 ( .A(n15306), .B(n15307), .Z(n15312) );
  XNOR U23669 ( .A(n15308), .B(n15309), .Z(n15307) );
  XNOR U23670 ( .A(y[6361]), .B(x[6361]), .Z(n15309) );
  XNOR U23671 ( .A(y[6362]), .B(x[6362]), .Z(n15308) );
  XNOR U23672 ( .A(y[6360]), .B(x[6360]), .Z(n15306) );
  XNOR U23673 ( .A(n15300), .B(n15301), .Z(n15311) );
  XNOR U23674 ( .A(y[6357]), .B(x[6357]), .Z(n15301) );
  XNOR U23675 ( .A(n15302), .B(n15303), .Z(n15300) );
  XNOR U23676 ( .A(y[6358]), .B(x[6358]), .Z(n15303) );
  XNOR U23677 ( .A(y[6359]), .B(x[6359]), .Z(n15302) );
  XOR U23678 ( .A(n15294), .B(n15293), .Z(n15295) );
  XNOR U23679 ( .A(n15289), .B(n15290), .Z(n15293) );
  XNOR U23680 ( .A(y[6354]), .B(x[6354]), .Z(n15290) );
  XNOR U23681 ( .A(n15291), .B(n15292), .Z(n15289) );
  XNOR U23682 ( .A(y[6355]), .B(x[6355]), .Z(n15292) );
  XNOR U23683 ( .A(y[6356]), .B(x[6356]), .Z(n15291) );
  XNOR U23684 ( .A(n15283), .B(n15284), .Z(n15294) );
  XNOR U23685 ( .A(y[6351]), .B(x[6351]), .Z(n15284) );
  XNOR U23686 ( .A(n15285), .B(n15286), .Z(n15283) );
  XNOR U23687 ( .A(y[6352]), .B(x[6352]), .Z(n15286) );
  XNOR U23688 ( .A(y[6353]), .B(x[6353]), .Z(n15285) );
  NAND U23689 ( .A(n15350), .B(n15351), .Z(N64028) );
  NANDN U23690 ( .A(n15352), .B(n15353), .Z(n15351) );
  OR U23691 ( .A(n15354), .B(n15355), .Z(n15353) );
  NAND U23692 ( .A(n15354), .B(n15355), .Z(n15350) );
  XOR U23693 ( .A(n15354), .B(n15356), .Z(N64027) );
  XNOR U23694 ( .A(n15352), .B(n15355), .Z(n15356) );
  AND U23695 ( .A(n15357), .B(n15358), .Z(n15355) );
  NANDN U23696 ( .A(n15359), .B(n15360), .Z(n15358) );
  NANDN U23697 ( .A(n15361), .B(n15362), .Z(n15360) );
  NANDN U23698 ( .A(n15362), .B(n15361), .Z(n15357) );
  NAND U23699 ( .A(n15363), .B(n15364), .Z(n15352) );
  NANDN U23700 ( .A(n15365), .B(n15366), .Z(n15364) );
  OR U23701 ( .A(n15367), .B(n15368), .Z(n15366) );
  NAND U23702 ( .A(n15368), .B(n15367), .Z(n15363) );
  AND U23703 ( .A(n15369), .B(n15370), .Z(n15354) );
  NANDN U23704 ( .A(n15371), .B(n15372), .Z(n15370) );
  NANDN U23705 ( .A(n15373), .B(n15374), .Z(n15372) );
  NANDN U23706 ( .A(n15374), .B(n15373), .Z(n15369) );
  XOR U23707 ( .A(n15368), .B(n15375), .Z(N64026) );
  XOR U23708 ( .A(n15365), .B(n15367), .Z(n15375) );
  XNOR U23709 ( .A(n15361), .B(n15376), .Z(n15367) );
  XNOR U23710 ( .A(n15359), .B(n15362), .Z(n15376) );
  NAND U23711 ( .A(n15377), .B(n15378), .Z(n15362) );
  NAND U23712 ( .A(n15379), .B(n15380), .Z(n15378) );
  OR U23713 ( .A(n15381), .B(n15382), .Z(n15379) );
  NANDN U23714 ( .A(n15383), .B(n15381), .Z(n15377) );
  IV U23715 ( .A(n15382), .Z(n15383) );
  NAND U23716 ( .A(n15384), .B(n15385), .Z(n15359) );
  NAND U23717 ( .A(n15386), .B(n15387), .Z(n15385) );
  NANDN U23718 ( .A(n15388), .B(n15389), .Z(n15386) );
  NANDN U23719 ( .A(n15389), .B(n15388), .Z(n15384) );
  AND U23720 ( .A(n15390), .B(n15391), .Z(n15361) );
  NAND U23721 ( .A(n15392), .B(n15393), .Z(n15391) );
  OR U23722 ( .A(n15394), .B(n15395), .Z(n15392) );
  NANDN U23723 ( .A(n15396), .B(n15394), .Z(n15390) );
  NAND U23724 ( .A(n15397), .B(n15398), .Z(n15365) );
  NANDN U23725 ( .A(n15399), .B(n15400), .Z(n15398) );
  OR U23726 ( .A(n15401), .B(n15402), .Z(n15400) );
  NANDN U23727 ( .A(n15403), .B(n15401), .Z(n15397) );
  IV U23728 ( .A(n15402), .Z(n15403) );
  XNOR U23729 ( .A(n15373), .B(n15404), .Z(n15368) );
  XNOR U23730 ( .A(n15371), .B(n15374), .Z(n15404) );
  NAND U23731 ( .A(n15405), .B(n15406), .Z(n15374) );
  NAND U23732 ( .A(n15407), .B(n15408), .Z(n15406) );
  OR U23733 ( .A(n15409), .B(n15410), .Z(n15407) );
  NANDN U23734 ( .A(n15411), .B(n15409), .Z(n15405) );
  IV U23735 ( .A(n15410), .Z(n15411) );
  NAND U23736 ( .A(n15412), .B(n15413), .Z(n15371) );
  NAND U23737 ( .A(n15414), .B(n15415), .Z(n15413) );
  NANDN U23738 ( .A(n15416), .B(n15417), .Z(n15414) );
  NANDN U23739 ( .A(n15417), .B(n15416), .Z(n15412) );
  AND U23740 ( .A(n15418), .B(n15419), .Z(n15373) );
  NAND U23741 ( .A(n15420), .B(n15421), .Z(n15419) );
  OR U23742 ( .A(n15422), .B(n15423), .Z(n15420) );
  NANDN U23743 ( .A(n15424), .B(n15422), .Z(n15418) );
  XNOR U23744 ( .A(n15399), .B(n15425), .Z(N64025) );
  XOR U23745 ( .A(n15401), .B(n15402), .Z(n15425) );
  XNOR U23746 ( .A(n15415), .B(n15426), .Z(n15402) );
  XOR U23747 ( .A(n15416), .B(n15417), .Z(n15426) );
  XOR U23748 ( .A(n15422), .B(n15427), .Z(n15417) );
  XOR U23749 ( .A(n15421), .B(n15424), .Z(n15427) );
  IV U23750 ( .A(n15423), .Z(n15424) );
  NAND U23751 ( .A(n15428), .B(n15429), .Z(n15423) );
  OR U23752 ( .A(n15430), .B(n15431), .Z(n15429) );
  OR U23753 ( .A(n15432), .B(n15433), .Z(n15428) );
  NAND U23754 ( .A(n15434), .B(n15435), .Z(n15421) );
  OR U23755 ( .A(n15436), .B(n15437), .Z(n15435) );
  OR U23756 ( .A(n15438), .B(n15439), .Z(n15434) );
  NOR U23757 ( .A(n15440), .B(n15441), .Z(n15422) );
  ANDN U23758 ( .B(n15442), .A(n15443), .Z(n15416) );
  XNOR U23759 ( .A(n15409), .B(n15444), .Z(n15415) );
  XNOR U23760 ( .A(n15408), .B(n15410), .Z(n15444) );
  NAND U23761 ( .A(n15445), .B(n15446), .Z(n15410) );
  OR U23762 ( .A(n15447), .B(n15448), .Z(n15446) );
  OR U23763 ( .A(n15449), .B(n15450), .Z(n15445) );
  NAND U23764 ( .A(n15451), .B(n15452), .Z(n15408) );
  OR U23765 ( .A(n15453), .B(n15454), .Z(n15452) );
  OR U23766 ( .A(n15455), .B(n15456), .Z(n15451) );
  ANDN U23767 ( .B(n15457), .A(n15458), .Z(n15409) );
  IV U23768 ( .A(n15459), .Z(n15457) );
  ANDN U23769 ( .B(n15460), .A(n15461), .Z(n15401) );
  XOR U23770 ( .A(n15387), .B(n15462), .Z(n15399) );
  XOR U23771 ( .A(n15388), .B(n15389), .Z(n15462) );
  XOR U23772 ( .A(n15394), .B(n15463), .Z(n15389) );
  XOR U23773 ( .A(n15393), .B(n15396), .Z(n15463) );
  IV U23774 ( .A(n15395), .Z(n15396) );
  NAND U23775 ( .A(n15464), .B(n15465), .Z(n15395) );
  OR U23776 ( .A(n15466), .B(n15467), .Z(n15465) );
  OR U23777 ( .A(n15468), .B(n15469), .Z(n15464) );
  NAND U23778 ( .A(n15470), .B(n15471), .Z(n15393) );
  OR U23779 ( .A(n15472), .B(n15473), .Z(n15471) );
  OR U23780 ( .A(n15474), .B(n15475), .Z(n15470) );
  NOR U23781 ( .A(n15476), .B(n15477), .Z(n15394) );
  ANDN U23782 ( .B(n15478), .A(n15479), .Z(n15388) );
  IV U23783 ( .A(n15480), .Z(n15478) );
  XNOR U23784 ( .A(n15381), .B(n15481), .Z(n15387) );
  XNOR U23785 ( .A(n15380), .B(n15382), .Z(n15481) );
  NAND U23786 ( .A(n15482), .B(n15483), .Z(n15382) );
  OR U23787 ( .A(n15484), .B(n15485), .Z(n15483) );
  OR U23788 ( .A(n15486), .B(n15487), .Z(n15482) );
  NAND U23789 ( .A(n15488), .B(n15489), .Z(n15380) );
  OR U23790 ( .A(n15490), .B(n15491), .Z(n15489) );
  OR U23791 ( .A(n15492), .B(n15493), .Z(n15488) );
  ANDN U23792 ( .B(n15494), .A(n15495), .Z(n15381) );
  IV U23793 ( .A(n15496), .Z(n15494) );
  XNOR U23794 ( .A(n15461), .B(n15460), .Z(N64024) );
  XOR U23795 ( .A(n15480), .B(n15479), .Z(n15460) );
  XNOR U23796 ( .A(n15495), .B(n15496), .Z(n15479) );
  XNOR U23797 ( .A(n15490), .B(n15491), .Z(n15496) );
  XNOR U23798 ( .A(n15492), .B(n15493), .Z(n15491) );
  XNOR U23799 ( .A(y[6349]), .B(x[6349]), .Z(n15493) );
  XNOR U23800 ( .A(y[6350]), .B(x[6350]), .Z(n15492) );
  XNOR U23801 ( .A(y[6348]), .B(x[6348]), .Z(n15490) );
  XNOR U23802 ( .A(n15484), .B(n15485), .Z(n15495) );
  XNOR U23803 ( .A(y[6345]), .B(x[6345]), .Z(n15485) );
  XNOR U23804 ( .A(n15486), .B(n15487), .Z(n15484) );
  XNOR U23805 ( .A(y[6346]), .B(x[6346]), .Z(n15487) );
  XNOR U23806 ( .A(y[6347]), .B(x[6347]), .Z(n15486) );
  XNOR U23807 ( .A(n15477), .B(n15476), .Z(n15480) );
  XNOR U23808 ( .A(n15472), .B(n15473), .Z(n15476) );
  XNOR U23809 ( .A(y[6342]), .B(x[6342]), .Z(n15473) );
  XNOR U23810 ( .A(n15474), .B(n15475), .Z(n15472) );
  XNOR U23811 ( .A(y[6343]), .B(x[6343]), .Z(n15475) );
  XNOR U23812 ( .A(y[6344]), .B(x[6344]), .Z(n15474) );
  XNOR U23813 ( .A(n15466), .B(n15467), .Z(n15477) );
  XNOR U23814 ( .A(y[6339]), .B(x[6339]), .Z(n15467) );
  XNOR U23815 ( .A(n15468), .B(n15469), .Z(n15466) );
  XNOR U23816 ( .A(y[6340]), .B(x[6340]), .Z(n15469) );
  XNOR U23817 ( .A(y[6341]), .B(x[6341]), .Z(n15468) );
  XOR U23818 ( .A(n15442), .B(n15443), .Z(n15461) );
  XNOR U23819 ( .A(n15458), .B(n15459), .Z(n15443) );
  XNOR U23820 ( .A(n15453), .B(n15454), .Z(n15459) );
  XNOR U23821 ( .A(n15455), .B(n15456), .Z(n15454) );
  XNOR U23822 ( .A(y[6337]), .B(x[6337]), .Z(n15456) );
  XNOR U23823 ( .A(y[6338]), .B(x[6338]), .Z(n15455) );
  XNOR U23824 ( .A(y[6336]), .B(x[6336]), .Z(n15453) );
  XNOR U23825 ( .A(n15447), .B(n15448), .Z(n15458) );
  XNOR U23826 ( .A(y[6333]), .B(x[6333]), .Z(n15448) );
  XNOR U23827 ( .A(n15449), .B(n15450), .Z(n15447) );
  XNOR U23828 ( .A(y[6334]), .B(x[6334]), .Z(n15450) );
  XNOR U23829 ( .A(y[6335]), .B(x[6335]), .Z(n15449) );
  XOR U23830 ( .A(n15441), .B(n15440), .Z(n15442) );
  XNOR U23831 ( .A(n15436), .B(n15437), .Z(n15440) );
  XNOR U23832 ( .A(y[6330]), .B(x[6330]), .Z(n15437) );
  XNOR U23833 ( .A(n15438), .B(n15439), .Z(n15436) );
  XNOR U23834 ( .A(y[6331]), .B(x[6331]), .Z(n15439) );
  XNOR U23835 ( .A(y[6332]), .B(x[6332]), .Z(n15438) );
  XNOR U23836 ( .A(n15430), .B(n15431), .Z(n15441) );
  XNOR U23837 ( .A(y[6327]), .B(x[6327]), .Z(n15431) );
  XNOR U23838 ( .A(n15432), .B(n15433), .Z(n15430) );
  XNOR U23839 ( .A(y[6328]), .B(x[6328]), .Z(n15433) );
  XNOR U23840 ( .A(y[6329]), .B(x[6329]), .Z(n15432) );
  NAND U23841 ( .A(n15497), .B(n15498), .Z(N64015) );
  NANDN U23842 ( .A(n15499), .B(n15500), .Z(n15498) );
  OR U23843 ( .A(n15501), .B(n15502), .Z(n15500) );
  NAND U23844 ( .A(n15501), .B(n15502), .Z(n15497) );
  XOR U23845 ( .A(n15501), .B(n15503), .Z(N64014) );
  XNOR U23846 ( .A(n15499), .B(n15502), .Z(n15503) );
  AND U23847 ( .A(n15504), .B(n15505), .Z(n15502) );
  NANDN U23848 ( .A(n15506), .B(n15507), .Z(n15505) );
  NANDN U23849 ( .A(n15508), .B(n15509), .Z(n15507) );
  NANDN U23850 ( .A(n15509), .B(n15508), .Z(n15504) );
  NAND U23851 ( .A(n15510), .B(n15511), .Z(n15499) );
  NANDN U23852 ( .A(n15512), .B(n15513), .Z(n15511) );
  OR U23853 ( .A(n15514), .B(n15515), .Z(n15513) );
  NAND U23854 ( .A(n15515), .B(n15514), .Z(n15510) );
  AND U23855 ( .A(n15516), .B(n15517), .Z(n15501) );
  NANDN U23856 ( .A(n15518), .B(n15519), .Z(n15517) );
  NANDN U23857 ( .A(n15520), .B(n15521), .Z(n15519) );
  NANDN U23858 ( .A(n15521), .B(n15520), .Z(n15516) );
  XOR U23859 ( .A(n15515), .B(n15522), .Z(N64013) );
  XOR U23860 ( .A(n15512), .B(n15514), .Z(n15522) );
  XNOR U23861 ( .A(n15508), .B(n15523), .Z(n15514) );
  XNOR U23862 ( .A(n15506), .B(n15509), .Z(n15523) );
  NAND U23863 ( .A(n15524), .B(n15525), .Z(n15509) );
  NAND U23864 ( .A(n15526), .B(n15527), .Z(n15525) );
  OR U23865 ( .A(n15528), .B(n15529), .Z(n15526) );
  NANDN U23866 ( .A(n15530), .B(n15528), .Z(n15524) );
  IV U23867 ( .A(n15529), .Z(n15530) );
  NAND U23868 ( .A(n15531), .B(n15532), .Z(n15506) );
  NAND U23869 ( .A(n15533), .B(n15534), .Z(n15532) );
  NANDN U23870 ( .A(n15535), .B(n15536), .Z(n15533) );
  NANDN U23871 ( .A(n15536), .B(n15535), .Z(n15531) );
  AND U23872 ( .A(n15537), .B(n15538), .Z(n15508) );
  NAND U23873 ( .A(n15539), .B(n15540), .Z(n15538) );
  OR U23874 ( .A(n15541), .B(n15542), .Z(n15539) );
  NANDN U23875 ( .A(n15543), .B(n15541), .Z(n15537) );
  NAND U23876 ( .A(n15544), .B(n15545), .Z(n15512) );
  NANDN U23877 ( .A(n15546), .B(n15547), .Z(n15545) );
  OR U23878 ( .A(n15548), .B(n15549), .Z(n15547) );
  NANDN U23879 ( .A(n15550), .B(n15548), .Z(n15544) );
  IV U23880 ( .A(n15549), .Z(n15550) );
  XNOR U23881 ( .A(n15520), .B(n15551), .Z(n15515) );
  XNOR U23882 ( .A(n15518), .B(n15521), .Z(n15551) );
  NAND U23883 ( .A(n15552), .B(n15553), .Z(n15521) );
  NAND U23884 ( .A(n15554), .B(n15555), .Z(n15553) );
  OR U23885 ( .A(n15556), .B(n15557), .Z(n15554) );
  NANDN U23886 ( .A(n15558), .B(n15556), .Z(n15552) );
  IV U23887 ( .A(n15557), .Z(n15558) );
  NAND U23888 ( .A(n15559), .B(n15560), .Z(n15518) );
  NAND U23889 ( .A(n15561), .B(n15562), .Z(n15560) );
  NANDN U23890 ( .A(n15563), .B(n15564), .Z(n15561) );
  NANDN U23891 ( .A(n15564), .B(n15563), .Z(n15559) );
  AND U23892 ( .A(n15565), .B(n15566), .Z(n15520) );
  NAND U23893 ( .A(n15567), .B(n15568), .Z(n15566) );
  OR U23894 ( .A(n15569), .B(n15570), .Z(n15567) );
  NANDN U23895 ( .A(n15571), .B(n15569), .Z(n15565) );
  XNOR U23896 ( .A(n15546), .B(n15572), .Z(N64012) );
  XOR U23897 ( .A(n15548), .B(n15549), .Z(n15572) );
  XNOR U23898 ( .A(n15562), .B(n15573), .Z(n15549) );
  XOR U23899 ( .A(n15563), .B(n15564), .Z(n15573) );
  XOR U23900 ( .A(n15569), .B(n15574), .Z(n15564) );
  XOR U23901 ( .A(n15568), .B(n15571), .Z(n15574) );
  IV U23902 ( .A(n15570), .Z(n15571) );
  NAND U23903 ( .A(n15575), .B(n15576), .Z(n15570) );
  OR U23904 ( .A(n15577), .B(n15578), .Z(n15576) );
  OR U23905 ( .A(n15579), .B(n15580), .Z(n15575) );
  NAND U23906 ( .A(n15581), .B(n15582), .Z(n15568) );
  OR U23907 ( .A(n15583), .B(n15584), .Z(n15582) );
  OR U23908 ( .A(n15585), .B(n15586), .Z(n15581) );
  NOR U23909 ( .A(n15587), .B(n15588), .Z(n15569) );
  ANDN U23910 ( .B(n15589), .A(n15590), .Z(n15563) );
  XNOR U23911 ( .A(n15556), .B(n15591), .Z(n15562) );
  XNOR U23912 ( .A(n15555), .B(n15557), .Z(n15591) );
  NAND U23913 ( .A(n15592), .B(n15593), .Z(n15557) );
  OR U23914 ( .A(n15594), .B(n15595), .Z(n15593) );
  OR U23915 ( .A(n15596), .B(n15597), .Z(n15592) );
  NAND U23916 ( .A(n15598), .B(n15599), .Z(n15555) );
  OR U23917 ( .A(n15600), .B(n15601), .Z(n15599) );
  OR U23918 ( .A(n15602), .B(n15603), .Z(n15598) );
  ANDN U23919 ( .B(n15604), .A(n15605), .Z(n15556) );
  IV U23920 ( .A(n15606), .Z(n15604) );
  ANDN U23921 ( .B(n15607), .A(n15608), .Z(n15548) );
  XOR U23922 ( .A(n15534), .B(n15609), .Z(n15546) );
  XOR U23923 ( .A(n15535), .B(n15536), .Z(n15609) );
  XOR U23924 ( .A(n15541), .B(n15610), .Z(n15536) );
  XOR U23925 ( .A(n15540), .B(n15543), .Z(n15610) );
  IV U23926 ( .A(n15542), .Z(n15543) );
  NAND U23927 ( .A(n15611), .B(n15612), .Z(n15542) );
  OR U23928 ( .A(n15613), .B(n15614), .Z(n15612) );
  OR U23929 ( .A(n15615), .B(n15616), .Z(n15611) );
  NAND U23930 ( .A(n15617), .B(n15618), .Z(n15540) );
  OR U23931 ( .A(n15619), .B(n15620), .Z(n15618) );
  OR U23932 ( .A(n15621), .B(n15622), .Z(n15617) );
  NOR U23933 ( .A(n15623), .B(n15624), .Z(n15541) );
  ANDN U23934 ( .B(n15625), .A(n15626), .Z(n15535) );
  IV U23935 ( .A(n15627), .Z(n15625) );
  XNOR U23936 ( .A(n15528), .B(n15628), .Z(n15534) );
  XNOR U23937 ( .A(n15527), .B(n15529), .Z(n15628) );
  NAND U23938 ( .A(n15629), .B(n15630), .Z(n15529) );
  OR U23939 ( .A(n15631), .B(n15632), .Z(n15630) );
  OR U23940 ( .A(n15633), .B(n15634), .Z(n15629) );
  NAND U23941 ( .A(n15635), .B(n15636), .Z(n15527) );
  OR U23942 ( .A(n15637), .B(n15638), .Z(n15636) );
  OR U23943 ( .A(n15639), .B(n15640), .Z(n15635) );
  ANDN U23944 ( .B(n15641), .A(n15642), .Z(n15528) );
  IV U23945 ( .A(n15643), .Z(n15641) );
  XNOR U23946 ( .A(n15608), .B(n15607), .Z(N64011) );
  XOR U23947 ( .A(n15627), .B(n15626), .Z(n15607) );
  XNOR U23948 ( .A(n15642), .B(n15643), .Z(n15626) );
  XNOR U23949 ( .A(n15637), .B(n15638), .Z(n15643) );
  XNOR U23950 ( .A(n15639), .B(n15640), .Z(n15638) );
  XNOR U23951 ( .A(y[6325]), .B(x[6325]), .Z(n15640) );
  XNOR U23952 ( .A(y[6326]), .B(x[6326]), .Z(n15639) );
  XNOR U23953 ( .A(y[6324]), .B(x[6324]), .Z(n15637) );
  XNOR U23954 ( .A(n15631), .B(n15632), .Z(n15642) );
  XNOR U23955 ( .A(y[6321]), .B(x[6321]), .Z(n15632) );
  XNOR U23956 ( .A(n15633), .B(n15634), .Z(n15631) );
  XNOR U23957 ( .A(y[6322]), .B(x[6322]), .Z(n15634) );
  XNOR U23958 ( .A(y[6323]), .B(x[6323]), .Z(n15633) );
  XNOR U23959 ( .A(n15624), .B(n15623), .Z(n15627) );
  XNOR U23960 ( .A(n15619), .B(n15620), .Z(n15623) );
  XNOR U23961 ( .A(y[6318]), .B(x[6318]), .Z(n15620) );
  XNOR U23962 ( .A(n15621), .B(n15622), .Z(n15619) );
  XNOR U23963 ( .A(y[6319]), .B(x[6319]), .Z(n15622) );
  XNOR U23964 ( .A(y[6320]), .B(x[6320]), .Z(n15621) );
  XNOR U23965 ( .A(n15613), .B(n15614), .Z(n15624) );
  XNOR U23966 ( .A(y[6315]), .B(x[6315]), .Z(n15614) );
  XNOR U23967 ( .A(n15615), .B(n15616), .Z(n15613) );
  XNOR U23968 ( .A(y[6316]), .B(x[6316]), .Z(n15616) );
  XNOR U23969 ( .A(y[6317]), .B(x[6317]), .Z(n15615) );
  XOR U23970 ( .A(n15589), .B(n15590), .Z(n15608) );
  XNOR U23971 ( .A(n15605), .B(n15606), .Z(n15590) );
  XNOR U23972 ( .A(n15600), .B(n15601), .Z(n15606) );
  XNOR U23973 ( .A(n15602), .B(n15603), .Z(n15601) );
  XNOR U23974 ( .A(y[6313]), .B(x[6313]), .Z(n15603) );
  XNOR U23975 ( .A(y[6314]), .B(x[6314]), .Z(n15602) );
  XNOR U23976 ( .A(y[6312]), .B(x[6312]), .Z(n15600) );
  XNOR U23977 ( .A(n15594), .B(n15595), .Z(n15605) );
  XNOR U23978 ( .A(y[6309]), .B(x[6309]), .Z(n15595) );
  XNOR U23979 ( .A(n15596), .B(n15597), .Z(n15594) );
  XNOR U23980 ( .A(y[6310]), .B(x[6310]), .Z(n15597) );
  XNOR U23981 ( .A(y[6311]), .B(x[6311]), .Z(n15596) );
  XOR U23982 ( .A(n15588), .B(n15587), .Z(n15589) );
  XNOR U23983 ( .A(n15583), .B(n15584), .Z(n15587) );
  XNOR U23984 ( .A(y[6306]), .B(x[6306]), .Z(n15584) );
  XNOR U23985 ( .A(n15585), .B(n15586), .Z(n15583) );
  XNOR U23986 ( .A(y[6307]), .B(x[6307]), .Z(n15586) );
  XNOR U23987 ( .A(y[6308]), .B(x[6308]), .Z(n15585) );
  XNOR U23988 ( .A(n15577), .B(n15578), .Z(n15588) );
  XNOR U23989 ( .A(y[6303]), .B(x[6303]), .Z(n15578) );
  XNOR U23990 ( .A(n15579), .B(n15580), .Z(n15577) );
  XNOR U23991 ( .A(y[6304]), .B(x[6304]), .Z(n15580) );
  XNOR U23992 ( .A(y[6305]), .B(x[6305]), .Z(n15579) );
  NAND U23993 ( .A(n15644), .B(n15645), .Z(N64002) );
  NANDN U23994 ( .A(n15646), .B(n15647), .Z(n15645) );
  OR U23995 ( .A(n15648), .B(n15649), .Z(n15647) );
  NAND U23996 ( .A(n15648), .B(n15649), .Z(n15644) );
  XOR U23997 ( .A(n15648), .B(n15650), .Z(N64001) );
  XNOR U23998 ( .A(n15646), .B(n15649), .Z(n15650) );
  AND U23999 ( .A(n15651), .B(n15652), .Z(n15649) );
  NANDN U24000 ( .A(n15653), .B(n15654), .Z(n15652) );
  NANDN U24001 ( .A(n15655), .B(n15656), .Z(n15654) );
  NANDN U24002 ( .A(n15656), .B(n15655), .Z(n15651) );
  NAND U24003 ( .A(n15657), .B(n15658), .Z(n15646) );
  NANDN U24004 ( .A(n15659), .B(n15660), .Z(n15658) );
  OR U24005 ( .A(n15661), .B(n15662), .Z(n15660) );
  NAND U24006 ( .A(n15662), .B(n15661), .Z(n15657) );
  AND U24007 ( .A(n15663), .B(n15664), .Z(n15648) );
  NANDN U24008 ( .A(n15665), .B(n15666), .Z(n15664) );
  NANDN U24009 ( .A(n15667), .B(n15668), .Z(n15666) );
  NANDN U24010 ( .A(n15668), .B(n15667), .Z(n15663) );
  XOR U24011 ( .A(n15662), .B(n15669), .Z(N64000) );
  XOR U24012 ( .A(n15659), .B(n15661), .Z(n15669) );
  XNOR U24013 ( .A(n15655), .B(n15670), .Z(n15661) );
  XNOR U24014 ( .A(n15653), .B(n15656), .Z(n15670) );
  NAND U24015 ( .A(n15671), .B(n15672), .Z(n15656) );
  NAND U24016 ( .A(n15673), .B(n15674), .Z(n15672) );
  OR U24017 ( .A(n15675), .B(n15676), .Z(n15673) );
  NANDN U24018 ( .A(n15677), .B(n15675), .Z(n15671) );
  IV U24019 ( .A(n15676), .Z(n15677) );
  NAND U24020 ( .A(n15678), .B(n15679), .Z(n15653) );
  NAND U24021 ( .A(n15680), .B(n15681), .Z(n15679) );
  NANDN U24022 ( .A(n15682), .B(n15683), .Z(n15680) );
  NANDN U24023 ( .A(n15683), .B(n15682), .Z(n15678) );
  AND U24024 ( .A(n15684), .B(n15685), .Z(n15655) );
  NAND U24025 ( .A(n15686), .B(n15687), .Z(n15685) );
  OR U24026 ( .A(n15688), .B(n15689), .Z(n15686) );
  NANDN U24027 ( .A(n15690), .B(n15688), .Z(n15684) );
  NAND U24028 ( .A(n15691), .B(n15692), .Z(n15659) );
  NANDN U24029 ( .A(n15693), .B(n15694), .Z(n15692) );
  OR U24030 ( .A(n15695), .B(n15696), .Z(n15694) );
  NANDN U24031 ( .A(n15697), .B(n15695), .Z(n15691) );
  IV U24032 ( .A(n15696), .Z(n15697) );
  XNOR U24033 ( .A(n15667), .B(n15698), .Z(n15662) );
  XNOR U24034 ( .A(n15665), .B(n15668), .Z(n15698) );
  NAND U24035 ( .A(n15699), .B(n15700), .Z(n15668) );
  NAND U24036 ( .A(n15701), .B(n15702), .Z(n15700) );
  OR U24037 ( .A(n15703), .B(n15704), .Z(n15701) );
  NANDN U24038 ( .A(n15705), .B(n15703), .Z(n15699) );
  IV U24039 ( .A(n15704), .Z(n15705) );
  NAND U24040 ( .A(n15706), .B(n15707), .Z(n15665) );
  NAND U24041 ( .A(n15708), .B(n15709), .Z(n15707) );
  NANDN U24042 ( .A(n15710), .B(n15711), .Z(n15708) );
  NANDN U24043 ( .A(n15711), .B(n15710), .Z(n15706) );
  AND U24044 ( .A(n15712), .B(n15713), .Z(n15667) );
  NAND U24045 ( .A(n15714), .B(n15715), .Z(n15713) );
  OR U24046 ( .A(n15716), .B(n15717), .Z(n15714) );
  NANDN U24047 ( .A(n15718), .B(n15716), .Z(n15712) );
  XNOR U24048 ( .A(n15693), .B(n15719), .Z(N63999) );
  XOR U24049 ( .A(n15695), .B(n15696), .Z(n15719) );
  XNOR U24050 ( .A(n15709), .B(n15720), .Z(n15696) );
  XOR U24051 ( .A(n15710), .B(n15711), .Z(n15720) );
  XOR U24052 ( .A(n15716), .B(n15721), .Z(n15711) );
  XOR U24053 ( .A(n15715), .B(n15718), .Z(n15721) );
  IV U24054 ( .A(n15717), .Z(n15718) );
  NAND U24055 ( .A(n15722), .B(n15723), .Z(n15717) );
  OR U24056 ( .A(n15724), .B(n15725), .Z(n15723) );
  OR U24057 ( .A(n15726), .B(n15727), .Z(n15722) );
  NAND U24058 ( .A(n15728), .B(n15729), .Z(n15715) );
  OR U24059 ( .A(n15730), .B(n15731), .Z(n15729) );
  OR U24060 ( .A(n15732), .B(n15733), .Z(n15728) );
  NOR U24061 ( .A(n15734), .B(n15735), .Z(n15716) );
  ANDN U24062 ( .B(n15736), .A(n15737), .Z(n15710) );
  XNOR U24063 ( .A(n15703), .B(n15738), .Z(n15709) );
  XNOR U24064 ( .A(n15702), .B(n15704), .Z(n15738) );
  NAND U24065 ( .A(n15739), .B(n15740), .Z(n15704) );
  OR U24066 ( .A(n15741), .B(n15742), .Z(n15740) );
  OR U24067 ( .A(n15743), .B(n15744), .Z(n15739) );
  NAND U24068 ( .A(n15745), .B(n15746), .Z(n15702) );
  OR U24069 ( .A(n15747), .B(n15748), .Z(n15746) );
  OR U24070 ( .A(n15749), .B(n15750), .Z(n15745) );
  ANDN U24071 ( .B(n15751), .A(n15752), .Z(n15703) );
  IV U24072 ( .A(n15753), .Z(n15751) );
  ANDN U24073 ( .B(n15754), .A(n15755), .Z(n15695) );
  XOR U24074 ( .A(n15681), .B(n15756), .Z(n15693) );
  XOR U24075 ( .A(n15682), .B(n15683), .Z(n15756) );
  XOR U24076 ( .A(n15688), .B(n15757), .Z(n15683) );
  XOR U24077 ( .A(n15687), .B(n15690), .Z(n15757) );
  IV U24078 ( .A(n15689), .Z(n15690) );
  NAND U24079 ( .A(n15758), .B(n15759), .Z(n15689) );
  OR U24080 ( .A(n15760), .B(n15761), .Z(n15759) );
  OR U24081 ( .A(n15762), .B(n15763), .Z(n15758) );
  NAND U24082 ( .A(n15764), .B(n15765), .Z(n15687) );
  OR U24083 ( .A(n15766), .B(n15767), .Z(n15765) );
  OR U24084 ( .A(n15768), .B(n15769), .Z(n15764) );
  NOR U24085 ( .A(n15770), .B(n15771), .Z(n15688) );
  ANDN U24086 ( .B(n15772), .A(n15773), .Z(n15682) );
  IV U24087 ( .A(n15774), .Z(n15772) );
  XNOR U24088 ( .A(n15675), .B(n15775), .Z(n15681) );
  XNOR U24089 ( .A(n15674), .B(n15676), .Z(n15775) );
  NAND U24090 ( .A(n15776), .B(n15777), .Z(n15676) );
  OR U24091 ( .A(n15778), .B(n15779), .Z(n15777) );
  OR U24092 ( .A(n15780), .B(n15781), .Z(n15776) );
  NAND U24093 ( .A(n15782), .B(n15783), .Z(n15674) );
  OR U24094 ( .A(n15784), .B(n15785), .Z(n15783) );
  OR U24095 ( .A(n15786), .B(n15787), .Z(n15782) );
  ANDN U24096 ( .B(n15788), .A(n15789), .Z(n15675) );
  IV U24097 ( .A(n15790), .Z(n15788) );
  XNOR U24098 ( .A(n15755), .B(n15754), .Z(N63998) );
  XOR U24099 ( .A(n15774), .B(n15773), .Z(n15754) );
  XNOR U24100 ( .A(n15789), .B(n15790), .Z(n15773) );
  XNOR U24101 ( .A(n15784), .B(n15785), .Z(n15790) );
  XNOR U24102 ( .A(n15786), .B(n15787), .Z(n15785) );
  XNOR U24103 ( .A(y[6301]), .B(x[6301]), .Z(n15787) );
  XNOR U24104 ( .A(y[6302]), .B(x[6302]), .Z(n15786) );
  XNOR U24105 ( .A(y[6300]), .B(x[6300]), .Z(n15784) );
  XNOR U24106 ( .A(n15778), .B(n15779), .Z(n15789) );
  XNOR U24107 ( .A(y[6297]), .B(x[6297]), .Z(n15779) );
  XNOR U24108 ( .A(n15780), .B(n15781), .Z(n15778) );
  XNOR U24109 ( .A(y[6298]), .B(x[6298]), .Z(n15781) );
  XNOR U24110 ( .A(y[6299]), .B(x[6299]), .Z(n15780) );
  XNOR U24111 ( .A(n15771), .B(n15770), .Z(n15774) );
  XNOR U24112 ( .A(n15766), .B(n15767), .Z(n15770) );
  XNOR U24113 ( .A(y[6294]), .B(x[6294]), .Z(n15767) );
  XNOR U24114 ( .A(n15768), .B(n15769), .Z(n15766) );
  XNOR U24115 ( .A(y[6295]), .B(x[6295]), .Z(n15769) );
  XNOR U24116 ( .A(y[6296]), .B(x[6296]), .Z(n15768) );
  XNOR U24117 ( .A(n15760), .B(n15761), .Z(n15771) );
  XNOR U24118 ( .A(y[6291]), .B(x[6291]), .Z(n15761) );
  XNOR U24119 ( .A(n15762), .B(n15763), .Z(n15760) );
  XNOR U24120 ( .A(y[6292]), .B(x[6292]), .Z(n15763) );
  XNOR U24121 ( .A(y[6293]), .B(x[6293]), .Z(n15762) );
  XOR U24122 ( .A(n15736), .B(n15737), .Z(n15755) );
  XNOR U24123 ( .A(n15752), .B(n15753), .Z(n15737) );
  XNOR U24124 ( .A(n15747), .B(n15748), .Z(n15753) );
  XNOR U24125 ( .A(n15749), .B(n15750), .Z(n15748) );
  XNOR U24126 ( .A(y[6289]), .B(x[6289]), .Z(n15750) );
  XNOR U24127 ( .A(y[6290]), .B(x[6290]), .Z(n15749) );
  XNOR U24128 ( .A(y[6288]), .B(x[6288]), .Z(n15747) );
  XNOR U24129 ( .A(n15741), .B(n15742), .Z(n15752) );
  XNOR U24130 ( .A(y[6285]), .B(x[6285]), .Z(n15742) );
  XNOR U24131 ( .A(n15743), .B(n15744), .Z(n15741) );
  XNOR U24132 ( .A(y[6286]), .B(x[6286]), .Z(n15744) );
  XNOR U24133 ( .A(y[6287]), .B(x[6287]), .Z(n15743) );
  XOR U24134 ( .A(n15735), .B(n15734), .Z(n15736) );
  XNOR U24135 ( .A(n15730), .B(n15731), .Z(n15734) );
  XNOR U24136 ( .A(y[6282]), .B(x[6282]), .Z(n15731) );
  XNOR U24137 ( .A(n15732), .B(n15733), .Z(n15730) );
  XNOR U24138 ( .A(y[6283]), .B(x[6283]), .Z(n15733) );
  XNOR U24139 ( .A(y[6284]), .B(x[6284]), .Z(n15732) );
  XNOR U24140 ( .A(n15724), .B(n15725), .Z(n15735) );
  XNOR U24141 ( .A(y[6279]), .B(x[6279]), .Z(n15725) );
  XNOR U24142 ( .A(n15726), .B(n15727), .Z(n15724) );
  XNOR U24143 ( .A(y[6280]), .B(x[6280]), .Z(n15727) );
  XNOR U24144 ( .A(y[6281]), .B(x[6281]), .Z(n15726) );
  NAND U24145 ( .A(n15791), .B(n15792), .Z(N63989) );
  NANDN U24146 ( .A(n15793), .B(n15794), .Z(n15792) );
  OR U24147 ( .A(n15795), .B(n15796), .Z(n15794) );
  NAND U24148 ( .A(n15795), .B(n15796), .Z(n15791) );
  XOR U24149 ( .A(n15795), .B(n15797), .Z(N63988) );
  XNOR U24150 ( .A(n15793), .B(n15796), .Z(n15797) );
  AND U24151 ( .A(n15798), .B(n15799), .Z(n15796) );
  NANDN U24152 ( .A(n15800), .B(n15801), .Z(n15799) );
  NANDN U24153 ( .A(n15802), .B(n15803), .Z(n15801) );
  NANDN U24154 ( .A(n15803), .B(n15802), .Z(n15798) );
  NAND U24155 ( .A(n15804), .B(n15805), .Z(n15793) );
  NANDN U24156 ( .A(n15806), .B(n15807), .Z(n15805) );
  OR U24157 ( .A(n15808), .B(n15809), .Z(n15807) );
  NAND U24158 ( .A(n15809), .B(n15808), .Z(n15804) );
  AND U24159 ( .A(n15810), .B(n15811), .Z(n15795) );
  NANDN U24160 ( .A(n15812), .B(n15813), .Z(n15811) );
  NANDN U24161 ( .A(n15814), .B(n15815), .Z(n15813) );
  NANDN U24162 ( .A(n15815), .B(n15814), .Z(n15810) );
  XOR U24163 ( .A(n15809), .B(n15816), .Z(N63987) );
  XOR U24164 ( .A(n15806), .B(n15808), .Z(n15816) );
  XNOR U24165 ( .A(n15802), .B(n15817), .Z(n15808) );
  XNOR U24166 ( .A(n15800), .B(n15803), .Z(n15817) );
  NAND U24167 ( .A(n15818), .B(n15819), .Z(n15803) );
  NAND U24168 ( .A(n15820), .B(n15821), .Z(n15819) );
  OR U24169 ( .A(n15822), .B(n15823), .Z(n15820) );
  NANDN U24170 ( .A(n15824), .B(n15822), .Z(n15818) );
  IV U24171 ( .A(n15823), .Z(n15824) );
  NAND U24172 ( .A(n15825), .B(n15826), .Z(n15800) );
  NAND U24173 ( .A(n15827), .B(n15828), .Z(n15826) );
  NANDN U24174 ( .A(n15829), .B(n15830), .Z(n15827) );
  NANDN U24175 ( .A(n15830), .B(n15829), .Z(n15825) );
  AND U24176 ( .A(n15831), .B(n15832), .Z(n15802) );
  NAND U24177 ( .A(n15833), .B(n15834), .Z(n15832) );
  OR U24178 ( .A(n15835), .B(n15836), .Z(n15833) );
  NANDN U24179 ( .A(n15837), .B(n15835), .Z(n15831) );
  NAND U24180 ( .A(n15838), .B(n15839), .Z(n15806) );
  NANDN U24181 ( .A(n15840), .B(n15841), .Z(n15839) );
  OR U24182 ( .A(n15842), .B(n15843), .Z(n15841) );
  NANDN U24183 ( .A(n15844), .B(n15842), .Z(n15838) );
  IV U24184 ( .A(n15843), .Z(n15844) );
  XNOR U24185 ( .A(n15814), .B(n15845), .Z(n15809) );
  XNOR U24186 ( .A(n15812), .B(n15815), .Z(n15845) );
  NAND U24187 ( .A(n15846), .B(n15847), .Z(n15815) );
  NAND U24188 ( .A(n15848), .B(n15849), .Z(n15847) );
  OR U24189 ( .A(n15850), .B(n15851), .Z(n15848) );
  NANDN U24190 ( .A(n15852), .B(n15850), .Z(n15846) );
  IV U24191 ( .A(n15851), .Z(n15852) );
  NAND U24192 ( .A(n15853), .B(n15854), .Z(n15812) );
  NAND U24193 ( .A(n15855), .B(n15856), .Z(n15854) );
  NANDN U24194 ( .A(n15857), .B(n15858), .Z(n15855) );
  NANDN U24195 ( .A(n15858), .B(n15857), .Z(n15853) );
  AND U24196 ( .A(n15859), .B(n15860), .Z(n15814) );
  NAND U24197 ( .A(n15861), .B(n15862), .Z(n15860) );
  OR U24198 ( .A(n15863), .B(n15864), .Z(n15861) );
  NANDN U24199 ( .A(n15865), .B(n15863), .Z(n15859) );
  XNOR U24200 ( .A(n15840), .B(n15866), .Z(N63986) );
  XOR U24201 ( .A(n15842), .B(n15843), .Z(n15866) );
  XNOR U24202 ( .A(n15856), .B(n15867), .Z(n15843) );
  XOR U24203 ( .A(n15857), .B(n15858), .Z(n15867) );
  XOR U24204 ( .A(n15863), .B(n15868), .Z(n15858) );
  XOR U24205 ( .A(n15862), .B(n15865), .Z(n15868) );
  IV U24206 ( .A(n15864), .Z(n15865) );
  NAND U24207 ( .A(n15869), .B(n15870), .Z(n15864) );
  OR U24208 ( .A(n15871), .B(n15872), .Z(n15870) );
  OR U24209 ( .A(n15873), .B(n15874), .Z(n15869) );
  NAND U24210 ( .A(n15875), .B(n15876), .Z(n15862) );
  OR U24211 ( .A(n15877), .B(n15878), .Z(n15876) );
  OR U24212 ( .A(n15879), .B(n15880), .Z(n15875) );
  NOR U24213 ( .A(n15881), .B(n15882), .Z(n15863) );
  ANDN U24214 ( .B(n15883), .A(n15884), .Z(n15857) );
  XNOR U24215 ( .A(n15850), .B(n15885), .Z(n15856) );
  XNOR U24216 ( .A(n15849), .B(n15851), .Z(n15885) );
  NAND U24217 ( .A(n15886), .B(n15887), .Z(n15851) );
  OR U24218 ( .A(n15888), .B(n15889), .Z(n15887) );
  OR U24219 ( .A(n15890), .B(n15891), .Z(n15886) );
  NAND U24220 ( .A(n15892), .B(n15893), .Z(n15849) );
  OR U24221 ( .A(n15894), .B(n15895), .Z(n15893) );
  OR U24222 ( .A(n15896), .B(n15897), .Z(n15892) );
  ANDN U24223 ( .B(n15898), .A(n15899), .Z(n15850) );
  IV U24224 ( .A(n15900), .Z(n15898) );
  ANDN U24225 ( .B(n15901), .A(n15902), .Z(n15842) );
  XOR U24226 ( .A(n15828), .B(n15903), .Z(n15840) );
  XOR U24227 ( .A(n15829), .B(n15830), .Z(n15903) );
  XOR U24228 ( .A(n15835), .B(n15904), .Z(n15830) );
  XOR U24229 ( .A(n15834), .B(n15837), .Z(n15904) );
  IV U24230 ( .A(n15836), .Z(n15837) );
  NAND U24231 ( .A(n15905), .B(n15906), .Z(n15836) );
  OR U24232 ( .A(n15907), .B(n15908), .Z(n15906) );
  OR U24233 ( .A(n15909), .B(n15910), .Z(n15905) );
  NAND U24234 ( .A(n15911), .B(n15912), .Z(n15834) );
  OR U24235 ( .A(n15913), .B(n15914), .Z(n15912) );
  OR U24236 ( .A(n15915), .B(n15916), .Z(n15911) );
  NOR U24237 ( .A(n15917), .B(n15918), .Z(n15835) );
  ANDN U24238 ( .B(n15919), .A(n15920), .Z(n15829) );
  IV U24239 ( .A(n15921), .Z(n15919) );
  XNOR U24240 ( .A(n15822), .B(n15922), .Z(n15828) );
  XNOR U24241 ( .A(n15821), .B(n15823), .Z(n15922) );
  NAND U24242 ( .A(n15923), .B(n15924), .Z(n15823) );
  OR U24243 ( .A(n15925), .B(n15926), .Z(n15924) );
  OR U24244 ( .A(n15927), .B(n15928), .Z(n15923) );
  NAND U24245 ( .A(n15929), .B(n15930), .Z(n15821) );
  OR U24246 ( .A(n15931), .B(n15932), .Z(n15930) );
  OR U24247 ( .A(n15933), .B(n15934), .Z(n15929) );
  ANDN U24248 ( .B(n15935), .A(n15936), .Z(n15822) );
  IV U24249 ( .A(n15937), .Z(n15935) );
  XNOR U24250 ( .A(n15902), .B(n15901), .Z(N63985) );
  XOR U24251 ( .A(n15921), .B(n15920), .Z(n15901) );
  XNOR U24252 ( .A(n15936), .B(n15937), .Z(n15920) );
  XNOR U24253 ( .A(n15931), .B(n15932), .Z(n15937) );
  XNOR U24254 ( .A(n15933), .B(n15934), .Z(n15932) );
  XNOR U24255 ( .A(y[6277]), .B(x[6277]), .Z(n15934) );
  XNOR U24256 ( .A(y[6278]), .B(x[6278]), .Z(n15933) );
  XNOR U24257 ( .A(y[6276]), .B(x[6276]), .Z(n15931) );
  XNOR U24258 ( .A(n15925), .B(n15926), .Z(n15936) );
  XNOR U24259 ( .A(y[6273]), .B(x[6273]), .Z(n15926) );
  XNOR U24260 ( .A(n15927), .B(n15928), .Z(n15925) );
  XNOR U24261 ( .A(y[6274]), .B(x[6274]), .Z(n15928) );
  XNOR U24262 ( .A(y[6275]), .B(x[6275]), .Z(n15927) );
  XNOR U24263 ( .A(n15918), .B(n15917), .Z(n15921) );
  XNOR U24264 ( .A(n15913), .B(n15914), .Z(n15917) );
  XNOR U24265 ( .A(y[6270]), .B(x[6270]), .Z(n15914) );
  XNOR U24266 ( .A(n15915), .B(n15916), .Z(n15913) );
  XNOR U24267 ( .A(y[6271]), .B(x[6271]), .Z(n15916) );
  XNOR U24268 ( .A(y[6272]), .B(x[6272]), .Z(n15915) );
  XNOR U24269 ( .A(n15907), .B(n15908), .Z(n15918) );
  XNOR U24270 ( .A(y[6267]), .B(x[6267]), .Z(n15908) );
  XNOR U24271 ( .A(n15909), .B(n15910), .Z(n15907) );
  XNOR U24272 ( .A(y[6268]), .B(x[6268]), .Z(n15910) );
  XNOR U24273 ( .A(y[6269]), .B(x[6269]), .Z(n15909) );
  XOR U24274 ( .A(n15883), .B(n15884), .Z(n15902) );
  XNOR U24275 ( .A(n15899), .B(n15900), .Z(n15884) );
  XNOR U24276 ( .A(n15894), .B(n15895), .Z(n15900) );
  XNOR U24277 ( .A(n15896), .B(n15897), .Z(n15895) );
  XNOR U24278 ( .A(y[6265]), .B(x[6265]), .Z(n15897) );
  XNOR U24279 ( .A(y[6266]), .B(x[6266]), .Z(n15896) );
  XNOR U24280 ( .A(y[6264]), .B(x[6264]), .Z(n15894) );
  XNOR U24281 ( .A(n15888), .B(n15889), .Z(n15899) );
  XNOR U24282 ( .A(y[6261]), .B(x[6261]), .Z(n15889) );
  XNOR U24283 ( .A(n15890), .B(n15891), .Z(n15888) );
  XNOR U24284 ( .A(y[6262]), .B(x[6262]), .Z(n15891) );
  XNOR U24285 ( .A(y[6263]), .B(x[6263]), .Z(n15890) );
  XOR U24286 ( .A(n15882), .B(n15881), .Z(n15883) );
  XNOR U24287 ( .A(n15877), .B(n15878), .Z(n15881) );
  XNOR U24288 ( .A(y[6258]), .B(x[6258]), .Z(n15878) );
  XNOR U24289 ( .A(n15879), .B(n15880), .Z(n15877) );
  XNOR U24290 ( .A(y[6259]), .B(x[6259]), .Z(n15880) );
  XNOR U24291 ( .A(y[6260]), .B(x[6260]), .Z(n15879) );
  XNOR U24292 ( .A(n15871), .B(n15872), .Z(n15882) );
  XNOR U24293 ( .A(y[6255]), .B(x[6255]), .Z(n15872) );
  XNOR U24294 ( .A(n15873), .B(n15874), .Z(n15871) );
  XNOR U24295 ( .A(y[6256]), .B(x[6256]), .Z(n15874) );
  XNOR U24296 ( .A(y[6257]), .B(x[6257]), .Z(n15873) );
  NAND U24297 ( .A(n15938), .B(n15939), .Z(N63976) );
  NANDN U24298 ( .A(n15940), .B(n15941), .Z(n15939) );
  OR U24299 ( .A(n15942), .B(n15943), .Z(n15941) );
  NAND U24300 ( .A(n15942), .B(n15943), .Z(n15938) );
  XOR U24301 ( .A(n15942), .B(n15944), .Z(N63975) );
  XNOR U24302 ( .A(n15940), .B(n15943), .Z(n15944) );
  AND U24303 ( .A(n15945), .B(n15946), .Z(n15943) );
  NANDN U24304 ( .A(n15947), .B(n15948), .Z(n15946) );
  NANDN U24305 ( .A(n15949), .B(n15950), .Z(n15948) );
  NANDN U24306 ( .A(n15950), .B(n15949), .Z(n15945) );
  NAND U24307 ( .A(n15951), .B(n15952), .Z(n15940) );
  NANDN U24308 ( .A(n15953), .B(n15954), .Z(n15952) );
  OR U24309 ( .A(n15955), .B(n15956), .Z(n15954) );
  NAND U24310 ( .A(n15956), .B(n15955), .Z(n15951) );
  AND U24311 ( .A(n15957), .B(n15958), .Z(n15942) );
  NANDN U24312 ( .A(n15959), .B(n15960), .Z(n15958) );
  NANDN U24313 ( .A(n15961), .B(n15962), .Z(n15960) );
  NANDN U24314 ( .A(n15962), .B(n15961), .Z(n15957) );
  XOR U24315 ( .A(n15956), .B(n15963), .Z(N63974) );
  XOR U24316 ( .A(n15953), .B(n15955), .Z(n15963) );
  XNOR U24317 ( .A(n15949), .B(n15964), .Z(n15955) );
  XNOR U24318 ( .A(n15947), .B(n15950), .Z(n15964) );
  NAND U24319 ( .A(n15965), .B(n15966), .Z(n15950) );
  NAND U24320 ( .A(n15967), .B(n15968), .Z(n15966) );
  OR U24321 ( .A(n15969), .B(n15970), .Z(n15967) );
  NANDN U24322 ( .A(n15971), .B(n15969), .Z(n15965) );
  IV U24323 ( .A(n15970), .Z(n15971) );
  NAND U24324 ( .A(n15972), .B(n15973), .Z(n15947) );
  NAND U24325 ( .A(n15974), .B(n15975), .Z(n15973) );
  NANDN U24326 ( .A(n15976), .B(n15977), .Z(n15974) );
  NANDN U24327 ( .A(n15977), .B(n15976), .Z(n15972) );
  AND U24328 ( .A(n15978), .B(n15979), .Z(n15949) );
  NAND U24329 ( .A(n15980), .B(n15981), .Z(n15979) );
  OR U24330 ( .A(n15982), .B(n15983), .Z(n15980) );
  NANDN U24331 ( .A(n15984), .B(n15982), .Z(n15978) );
  NAND U24332 ( .A(n15985), .B(n15986), .Z(n15953) );
  NANDN U24333 ( .A(n15987), .B(n15988), .Z(n15986) );
  OR U24334 ( .A(n15989), .B(n15990), .Z(n15988) );
  NANDN U24335 ( .A(n15991), .B(n15989), .Z(n15985) );
  IV U24336 ( .A(n15990), .Z(n15991) );
  XNOR U24337 ( .A(n15961), .B(n15992), .Z(n15956) );
  XNOR U24338 ( .A(n15959), .B(n15962), .Z(n15992) );
  NAND U24339 ( .A(n15993), .B(n15994), .Z(n15962) );
  NAND U24340 ( .A(n15995), .B(n15996), .Z(n15994) );
  OR U24341 ( .A(n15997), .B(n15998), .Z(n15995) );
  NANDN U24342 ( .A(n15999), .B(n15997), .Z(n15993) );
  IV U24343 ( .A(n15998), .Z(n15999) );
  NAND U24344 ( .A(n16000), .B(n16001), .Z(n15959) );
  NAND U24345 ( .A(n16002), .B(n16003), .Z(n16001) );
  NANDN U24346 ( .A(n16004), .B(n16005), .Z(n16002) );
  NANDN U24347 ( .A(n16005), .B(n16004), .Z(n16000) );
  AND U24348 ( .A(n16006), .B(n16007), .Z(n15961) );
  NAND U24349 ( .A(n16008), .B(n16009), .Z(n16007) );
  OR U24350 ( .A(n16010), .B(n16011), .Z(n16008) );
  NANDN U24351 ( .A(n16012), .B(n16010), .Z(n16006) );
  XNOR U24352 ( .A(n15987), .B(n16013), .Z(N63973) );
  XOR U24353 ( .A(n15989), .B(n15990), .Z(n16013) );
  XNOR U24354 ( .A(n16003), .B(n16014), .Z(n15990) );
  XOR U24355 ( .A(n16004), .B(n16005), .Z(n16014) );
  XOR U24356 ( .A(n16010), .B(n16015), .Z(n16005) );
  XOR U24357 ( .A(n16009), .B(n16012), .Z(n16015) );
  IV U24358 ( .A(n16011), .Z(n16012) );
  NAND U24359 ( .A(n16016), .B(n16017), .Z(n16011) );
  OR U24360 ( .A(n16018), .B(n16019), .Z(n16017) );
  OR U24361 ( .A(n16020), .B(n16021), .Z(n16016) );
  NAND U24362 ( .A(n16022), .B(n16023), .Z(n16009) );
  OR U24363 ( .A(n16024), .B(n16025), .Z(n16023) );
  OR U24364 ( .A(n16026), .B(n16027), .Z(n16022) );
  NOR U24365 ( .A(n16028), .B(n16029), .Z(n16010) );
  ANDN U24366 ( .B(n16030), .A(n16031), .Z(n16004) );
  XNOR U24367 ( .A(n15997), .B(n16032), .Z(n16003) );
  XNOR U24368 ( .A(n15996), .B(n15998), .Z(n16032) );
  NAND U24369 ( .A(n16033), .B(n16034), .Z(n15998) );
  OR U24370 ( .A(n16035), .B(n16036), .Z(n16034) );
  OR U24371 ( .A(n16037), .B(n16038), .Z(n16033) );
  NAND U24372 ( .A(n16039), .B(n16040), .Z(n15996) );
  OR U24373 ( .A(n16041), .B(n16042), .Z(n16040) );
  OR U24374 ( .A(n16043), .B(n16044), .Z(n16039) );
  ANDN U24375 ( .B(n16045), .A(n16046), .Z(n15997) );
  IV U24376 ( .A(n16047), .Z(n16045) );
  ANDN U24377 ( .B(n16048), .A(n16049), .Z(n15989) );
  XOR U24378 ( .A(n15975), .B(n16050), .Z(n15987) );
  XOR U24379 ( .A(n15976), .B(n15977), .Z(n16050) );
  XOR U24380 ( .A(n15982), .B(n16051), .Z(n15977) );
  XOR U24381 ( .A(n15981), .B(n15984), .Z(n16051) );
  IV U24382 ( .A(n15983), .Z(n15984) );
  NAND U24383 ( .A(n16052), .B(n16053), .Z(n15983) );
  OR U24384 ( .A(n16054), .B(n16055), .Z(n16053) );
  OR U24385 ( .A(n16056), .B(n16057), .Z(n16052) );
  NAND U24386 ( .A(n16058), .B(n16059), .Z(n15981) );
  OR U24387 ( .A(n16060), .B(n16061), .Z(n16059) );
  OR U24388 ( .A(n16062), .B(n16063), .Z(n16058) );
  NOR U24389 ( .A(n16064), .B(n16065), .Z(n15982) );
  ANDN U24390 ( .B(n16066), .A(n16067), .Z(n15976) );
  IV U24391 ( .A(n16068), .Z(n16066) );
  XNOR U24392 ( .A(n15969), .B(n16069), .Z(n15975) );
  XNOR U24393 ( .A(n15968), .B(n15970), .Z(n16069) );
  NAND U24394 ( .A(n16070), .B(n16071), .Z(n15970) );
  OR U24395 ( .A(n16072), .B(n16073), .Z(n16071) );
  OR U24396 ( .A(n16074), .B(n16075), .Z(n16070) );
  NAND U24397 ( .A(n16076), .B(n16077), .Z(n15968) );
  OR U24398 ( .A(n16078), .B(n16079), .Z(n16077) );
  OR U24399 ( .A(n16080), .B(n16081), .Z(n16076) );
  ANDN U24400 ( .B(n16082), .A(n16083), .Z(n15969) );
  IV U24401 ( .A(n16084), .Z(n16082) );
  XNOR U24402 ( .A(n16049), .B(n16048), .Z(N63972) );
  XOR U24403 ( .A(n16068), .B(n16067), .Z(n16048) );
  XNOR U24404 ( .A(n16083), .B(n16084), .Z(n16067) );
  XNOR U24405 ( .A(n16078), .B(n16079), .Z(n16084) );
  XNOR U24406 ( .A(n16080), .B(n16081), .Z(n16079) );
  XNOR U24407 ( .A(y[6253]), .B(x[6253]), .Z(n16081) );
  XNOR U24408 ( .A(y[6254]), .B(x[6254]), .Z(n16080) );
  XNOR U24409 ( .A(y[6252]), .B(x[6252]), .Z(n16078) );
  XNOR U24410 ( .A(n16072), .B(n16073), .Z(n16083) );
  XNOR U24411 ( .A(y[6249]), .B(x[6249]), .Z(n16073) );
  XNOR U24412 ( .A(n16074), .B(n16075), .Z(n16072) );
  XNOR U24413 ( .A(y[6250]), .B(x[6250]), .Z(n16075) );
  XNOR U24414 ( .A(y[6251]), .B(x[6251]), .Z(n16074) );
  XNOR U24415 ( .A(n16065), .B(n16064), .Z(n16068) );
  XNOR U24416 ( .A(n16060), .B(n16061), .Z(n16064) );
  XNOR U24417 ( .A(y[6246]), .B(x[6246]), .Z(n16061) );
  XNOR U24418 ( .A(n16062), .B(n16063), .Z(n16060) );
  XNOR U24419 ( .A(y[6247]), .B(x[6247]), .Z(n16063) );
  XNOR U24420 ( .A(y[6248]), .B(x[6248]), .Z(n16062) );
  XNOR U24421 ( .A(n16054), .B(n16055), .Z(n16065) );
  XNOR U24422 ( .A(y[6243]), .B(x[6243]), .Z(n16055) );
  XNOR U24423 ( .A(n16056), .B(n16057), .Z(n16054) );
  XNOR U24424 ( .A(y[6244]), .B(x[6244]), .Z(n16057) );
  XNOR U24425 ( .A(y[6245]), .B(x[6245]), .Z(n16056) );
  XOR U24426 ( .A(n16030), .B(n16031), .Z(n16049) );
  XNOR U24427 ( .A(n16046), .B(n16047), .Z(n16031) );
  XNOR U24428 ( .A(n16041), .B(n16042), .Z(n16047) );
  XNOR U24429 ( .A(n16043), .B(n16044), .Z(n16042) );
  XNOR U24430 ( .A(y[6241]), .B(x[6241]), .Z(n16044) );
  XNOR U24431 ( .A(y[6242]), .B(x[6242]), .Z(n16043) );
  XNOR U24432 ( .A(y[6240]), .B(x[6240]), .Z(n16041) );
  XNOR U24433 ( .A(n16035), .B(n16036), .Z(n16046) );
  XNOR U24434 ( .A(y[6237]), .B(x[6237]), .Z(n16036) );
  XNOR U24435 ( .A(n16037), .B(n16038), .Z(n16035) );
  XNOR U24436 ( .A(y[6238]), .B(x[6238]), .Z(n16038) );
  XNOR U24437 ( .A(y[6239]), .B(x[6239]), .Z(n16037) );
  XOR U24438 ( .A(n16029), .B(n16028), .Z(n16030) );
  XNOR U24439 ( .A(n16024), .B(n16025), .Z(n16028) );
  XNOR U24440 ( .A(y[6234]), .B(x[6234]), .Z(n16025) );
  XNOR U24441 ( .A(n16026), .B(n16027), .Z(n16024) );
  XNOR U24442 ( .A(y[6235]), .B(x[6235]), .Z(n16027) );
  XNOR U24443 ( .A(y[6236]), .B(x[6236]), .Z(n16026) );
  XNOR U24444 ( .A(n16018), .B(n16019), .Z(n16029) );
  XNOR U24445 ( .A(y[6231]), .B(x[6231]), .Z(n16019) );
  XNOR U24446 ( .A(n16020), .B(n16021), .Z(n16018) );
  XNOR U24447 ( .A(y[6232]), .B(x[6232]), .Z(n16021) );
  XNOR U24448 ( .A(y[6233]), .B(x[6233]), .Z(n16020) );
  NAND U24449 ( .A(n16085), .B(n16086), .Z(N63963) );
  NANDN U24450 ( .A(n16087), .B(n16088), .Z(n16086) );
  OR U24451 ( .A(n16089), .B(n16090), .Z(n16088) );
  NAND U24452 ( .A(n16089), .B(n16090), .Z(n16085) );
  XOR U24453 ( .A(n16089), .B(n16091), .Z(N63962) );
  XNOR U24454 ( .A(n16087), .B(n16090), .Z(n16091) );
  AND U24455 ( .A(n16092), .B(n16093), .Z(n16090) );
  NANDN U24456 ( .A(n16094), .B(n16095), .Z(n16093) );
  NANDN U24457 ( .A(n16096), .B(n16097), .Z(n16095) );
  NANDN U24458 ( .A(n16097), .B(n16096), .Z(n16092) );
  NAND U24459 ( .A(n16098), .B(n16099), .Z(n16087) );
  NANDN U24460 ( .A(n16100), .B(n16101), .Z(n16099) );
  OR U24461 ( .A(n16102), .B(n16103), .Z(n16101) );
  NAND U24462 ( .A(n16103), .B(n16102), .Z(n16098) );
  AND U24463 ( .A(n16104), .B(n16105), .Z(n16089) );
  NANDN U24464 ( .A(n16106), .B(n16107), .Z(n16105) );
  NANDN U24465 ( .A(n16108), .B(n16109), .Z(n16107) );
  NANDN U24466 ( .A(n16109), .B(n16108), .Z(n16104) );
  XOR U24467 ( .A(n16103), .B(n16110), .Z(N63961) );
  XOR U24468 ( .A(n16100), .B(n16102), .Z(n16110) );
  XNOR U24469 ( .A(n16096), .B(n16111), .Z(n16102) );
  XNOR U24470 ( .A(n16094), .B(n16097), .Z(n16111) );
  NAND U24471 ( .A(n16112), .B(n16113), .Z(n16097) );
  NAND U24472 ( .A(n16114), .B(n16115), .Z(n16113) );
  OR U24473 ( .A(n16116), .B(n16117), .Z(n16114) );
  NANDN U24474 ( .A(n16118), .B(n16116), .Z(n16112) );
  IV U24475 ( .A(n16117), .Z(n16118) );
  NAND U24476 ( .A(n16119), .B(n16120), .Z(n16094) );
  NAND U24477 ( .A(n16121), .B(n16122), .Z(n16120) );
  NANDN U24478 ( .A(n16123), .B(n16124), .Z(n16121) );
  NANDN U24479 ( .A(n16124), .B(n16123), .Z(n16119) );
  AND U24480 ( .A(n16125), .B(n16126), .Z(n16096) );
  NAND U24481 ( .A(n16127), .B(n16128), .Z(n16126) );
  OR U24482 ( .A(n16129), .B(n16130), .Z(n16127) );
  NANDN U24483 ( .A(n16131), .B(n16129), .Z(n16125) );
  NAND U24484 ( .A(n16132), .B(n16133), .Z(n16100) );
  NANDN U24485 ( .A(n16134), .B(n16135), .Z(n16133) );
  OR U24486 ( .A(n16136), .B(n16137), .Z(n16135) );
  NANDN U24487 ( .A(n16138), .B(n16136), .Z(n16132) );
  IV U24488 ( .A(n16137), .Z(n16138) );
  XNOR U24489 ( .A(n16108), .B(n16139), .Z(n16103) );
  XNOR U24490 ( .A(n16106), .B(n16109), .Z(n16139) );
  NAND U24491 ( .A(n16140), .B(n16141), .Z(n16109) );
  NAND U24492 ( .A(n16142), .B(n16143), .Z(n16141) );
  OR U24493 ( .A(n16144), .B(n16145), .Z(n16142) );
  NANDN U24494 ( .A(n16146), .B(n16144), .Z(n16140) );
  IV U24495 ( .A(n16145), .Z(n16146) );
  NAND U24496 ( .A(n16147), .B(n16148), .Z(n16106) );
  NAND U24497 ( .A(n16149), .B(n16150), .Z(n16148) );
  NANDN U24498 ( .A(n16151), .B(n16152), .Z(n16149) );
  NANDN U24499 ( .A(n16152), .B(n16151), .Z(n16147) );
  AND U24500 ( .A(n16153), .B(n16154), .Z(n16108) );
  NAND U24501 ( .A(n16155), .B(n16156), .Z(n16154) );
  OR U24502 ( .A(n16157), .B(n16158), .Z(n16155) );
  NANDN U24503 ( .A(n16159), .B(n16157), .Z(n16153) );
  XNOR U24504 ( .A(n16134), .B(n16160), .Z(N63960) );
  XOR U24505 ( .A(n16136), .B(n16137), .Z(n16160) );
  XNOR U24506 ( .A(n16150), .B(n16161), .Z(n16137) );
  XOR U24507 ( .A(n16151), .B(n16152), .Z(n16161) );
  XOR U24508 ( .A(n16157), .B(n16162), .Z(n16152) );
  XOR U24509 ( .A(n16156), .B(n16159), .Z(n16162) );
  IV U24510 ( .A(n16158), .Z(n16159) );
  NAND U24511 ( .A(n16163), .B(n16164), .Z(n16158) );
  OR U24512 ( .A(n16165), .B(n16166), .Z(n16164) );
  OR U24513 ( .A(n16167), .B(n16168), .Z(n16163) );
  NAND U24514 ( .A(n16169), .B(n16170), .Z(n16156) );
  OR U24515 ( .A(n16171), .B(n16172), .Z(n16170) );
  OR U24516 ( .A(n16173), .B(n16174), .Z(n16169) );
  NOR U24517 ( .A(n16175), .B(n16176), .Z(n16157) );
  ANDN U24518 ( .B(n16177), .A(n16178), .Z(n16151) );
  XNOR U24519 ( .A(n16144), .B(n16179), .Z(n16150) );
  XNOR U24520 ( .A(n16143), .B(n16145), .Z(n16179) );
  NAND U24521 ( .A(n16180), .B(n16181), .Z(n16145) );
  OR U24522 ( .A(n16182), .B(n16183), .Z(n16181) );
  OR U24523 ( .A(n16184), .B(n16185), .Z(n16180) );
  NAND U24524 ( .A(n16186), .B(n16187), .Z(n16143) );
  OR U24525 ( .A(n16188), .B(n16189), .Z(n16187) );
  OR U24526 ( .A(n16190), .B(n16191), .Z(n16186) );
  ANDN U24527 ( .B(n16192), .A(n16193), .Z(n16144) );
  IV U24528 ( .A(n16194), .Z(n16192) );
  ANDN U24529 ( .B(n16195), .A(n16196), .Z(n16136) );
  XOR U24530 ( .A(n16122), .B(n16197), .Z(n16134) );
  XOR U24531 ( .A(n16123), .B(n16124), .Z(n16197) );
  XOR U24532 ( .A(n16129), .B(n16198), .Z(n16124) );
  XOR U24533 ( .A(n16128), .B(n16131), .Z(n16198) );
  IV U24534 ( .A(n16130), .Z(n16131) );
  NAND U24535 ( .A(n16199), .B(n16200), .Z(n16130) );
  OR U24536 ( .A(n16201), .B(n16202), .Z(n16200) );
  OR U24537 ( .A(n16203), .B(n16204), .Z(n16199) );
  NAND U24538 ( .A(n16205), .B(n16206), .Z(n16128) );
  OR U24539 ( .A(n16207), .B(n16208), .Z(n16206) );
  OR U24540 ( .A(n16209), .B(n16210), .Z(n16205) );
  NOR U24541 ( .A(n16211), .B(n16212), .Z(n16129) );
  ANDN U24542 ( .B(n16213), .A(n16214), .Z(n16123) );
  IV U24543 ( .A(n16215), .Z(n16213) );
  XNOR U24544 ( .A(n16116), .B(n16216), .Z(n16122) );
  XNOR U24545 ( .A(n16115), .B(n16117), .Z(n16216) );
  NAND U24546 ( .A(n16217), .B(n16218), .Z(n16117) );
  OR U24547 ( .A(n16219), .B(n16220), .Z(n16218) );
  OR U24548 ( .A(n16221), .B(n16222), .Z(n16217) );
  NAND U24549 ( .A(n16223), .B(n16224), .Z(n16115) );
  OR U24550 ( .A(n16225), .B(n16226), .Z(n16224) );
  OR U24551 ( .A(n16227), .B(n16228), .Z(n16223) );
  ANDN U24552 ( .B(n16229), .A(n16230), .Z(n16116) );
  IV U24553 ( .A(n16231), .Z(n16229) );
  XNOR U24554 ( .A(n16196), .B(n16195), .Z(N63959) );
  XOR U24555 ( .A(n16215), .B(n16214), .Z(n16195) );
  XNOR U24556 ( .A(n16230), .B(n16231), .Z(n16214) );
  XNOR U24557 ( .A(n16225), .B(n16226), .Z(n16231) );
  XNOR U24558 ( .A(n16227), .B(n16228), .Z(n16226) );
  XNOR U24559 ( .A(y[6229]), .B(x[6229]), .Z(n16228) );
  XNOR U24560 ( .A(y[6230]), .B(x[6230]), .Z(n16227) );
  XNOR U24561 ( .A(y[6228]), .B(x[6228]), .Z(n16225) );
  XNOR U24562 ( .A(n16219), .B(n16220), .Z(n16230) );
  XNOR U24563 ( .A(y[6225]), .B(x[6225]), .Z(n16220) );
  XNOR U24564 ( .A(n16221), .B(n16222), .Z(n16219) );
  XNOR U24565 ( .A(y[6226]), .B(x[6226]), .Z(n16222) );
  XNOR U24566 ( .A(y[6227]), .B(x[6227]), .Z(n16221) );
  XNOR U24567 ( .A(n16212), .B(n16211), .Z(n16215) );
  XNOR U24568 ( .A(n16207), .B(n16208), .Z(n16211) );
  XNOR U24569 ( .A(y[6222]), .B(x[6222]), .Z(n16208) );
  XNOR U24570 ( .A(n16209), .B(n16210), .Z(n16207) );
  XNOR U24571 ( .A(y[6223]), .B(x[6223]), .Z(n16210) );
  XNOR U24572 ( .A(y[6224]), .B(x[6224]), .Z(n16209) );
  XNOR U24573 ( .A(n16201), .B(n16202), .Z(n16212) );
  XNOR U24574 ( .A(y[6219]), .B(x[6219]), .Z(n16202) );
  XNOR U24575 ( .A(n16203), .B(n16204), .Z(n16201) );
  XNOR U24576 ( .A(y[6220]), .B(x[6220]), .Z(n16204) );
  XNOR U24577 ( .A(y[6221]), .B(x[6221]), .Z(n16203) );
  XOR U24578 ( .A(n16177), .B(n16178), .Z(n16196) );
  XNOR U24579 ( .A(n16193), .B(n16194), .Z(n16178) );
  XNOR U24580 ( .A(n16188), .B(n16189), .Z(n16194) );
  XNOR U24581 ( .A(n16190), .B(n16191), .Z(n16189) );
  XNOR U24582 ( .A(y[6217]), .B(x[6217]), .Z(n16191) );
  XNOR U24583 ( .A(y[6218]), .B(x[6218]), .Z(n16190) );
  XNOR U24584 ( .A(y[6216]), .B(x[6216]), .Z(n16188) );
  XNOR U24585 ( .A(n16182), .B(n16183), .Z(n16193) );
  XNOR U24586 ( .A(y[6213]), .B(x[6213]), .Z(n16183) );
  XNOR U24587 ( .A(n16184), .B(n16185), .Z(n16182) );
  XNOR U24588 ( .A(y[6214]), .B(x[6214]), .Z(n16185) );
  XNOR U24589 ( .A(y[6215]), .B(x[6215]), .Z(n16184) );
  XOR U24590 ( .A(n16176), .B(n16175), .Z(n16177) );
  XNOR U24591 ( .A(n16171), .B(n16172), .Z(n16175) );
  XNOR U24592 ( .A(y[6210]), .B(x[6210]), .Z(n16172) );
  XNOR U24593 ( .A(n16173), .B(n16174), .Z(n16171) );
  XNOR U24594 ( .A(y[6211]), .B(x[6211]), .Z(n16174) );
  XNOR U24595 ( .A(y[6212]), .B(x[6212]), .Z(n16173) );
  XNOR U24596 ( .A(n16165), .B(n16166), .Z(n16176) );
  XNOR U24597 ( .A(y[6207]), .B(x[6207]), .Z(n16166) );
  XNOR U24598 ( .A(n16167), .B(n16168), .Z(n16165) );
  XNOR U24599 ( .A(y[6208]), .B(x[6208]), .Z(n16168) );
  XNOR U24600 ( .A(y[6209]), .B(x[6209]), .Z(n16167) );
  NAND U24601 ( .A(n16232), .B(n16233), .Z(N63950) );
  NANDN U24602 ( .A(n16234), .B(n16235), .Z(n16233) );
  OR U24603 ( .A(n16236), .B(n16237), .Z(n16235) );
  NAND U24604 ( .A(n16236), .B(n16237), .Z(n16232) );
  XOR U24605 ( .A(n16236), .B(n16238), .Z(N63949) );
  XNOR U24606 ( .A(n16234), .B(n16237), .Z(n16238) );
  AND U24607 ( .A(n16239), .B(n16240), .Z(n16237) );
  NANDN U24608 ( .A(n16241), .B(n16242), .Z(n16240) );
  NANDN U24609 ( .A(n16243), .B(n16244), .Z(n16242) );
  NANDN U24610 ( .A(n16244), .B(n16243), .Z(n16239) );
  NAND U24611 ( .A(n16245), .B(n16246), .Z(n16234) );
  NANDN U24612 ( .A(n16247), .B(n16248), .Z(n16246) );
  OR U24613 ( .A(n16249), .B(n16250), .Z(n16248) );
  NAND U24614 ( .A(n16250), .B(n16249), .Z(n16245) );
  AND U24615 ( .A(n16251), .B(n16252), .Z(n16236) );
  NANDN U24616 ( .A(n16253), .B(n16254), .Z(n16252) );
  NANDN U24617 ( .A(n16255), .B(n16256), .Z(n16254) );
  NANDN U24618 ( .A(n16256), .B(n16255), .Z(n16251) );
  XOR U24619 ( .A(n16250), .B(n16257), .Z(N63948) );
  XOR U24620 ( .A(n16247), .B(n16249), .Z(n16257) );
  XNOR U24621 ( .A(n16243), .B(n16258), .Z(n16249) );
  XNOR U24622 ( .A(n16241), .B(n16244), .Z(n16258) );
  NAND U24623 ( .A(n16259), .B(n16260), .Z(n16244) );
  NAND U24624 ( .A(n16261), .B(n16262), .Z(n16260) );
  OR U24625 ( .A(n16263), .B(n16264), .Z(n16261) );
  NANDN U24626 ( .A(n16265), .B(n16263), .Z(n16259) );
  IV U24627 ( .A(n16264), .Z(n16265) );
  NAND U24628 ( .A(n16266), .B(n16267), .Z(n16241) );
  NAND U24629 ( .A(n16268), .B(n16269), .Z(n16267) );
  NANDN U24630 ( .A(n16270), .B(n16271), .Z(n16268) );
  NANDN U24631 ( .A(n16271), .B(n16270), .Z(n16266) );
  AND U24632 ( .A(n16272), .B(n16273), .Z(n16243) );
  NAND U24633 ( .A(n16274), .B(n16275), .Z(n16273) );
  OR U24634 ( .A(n16276), .B(n16277), .Z(n16274) );
  NANDN U24635 ( .A(n16278), .B(n16276), .Z(n16272) );
  NAND U24636 ( .A(n16279), .B(n16280), .Z(n16247) );
  NANDN U24637 ( .A(n16281), .B(n16282), .Z(n16280) );
  OR U24638 ( .A(n16283), .B(n16284), .Z(n16282) );
  NANDN U24639 ( .A(n16285), .B(n16283), .Z(n16279) );
  IV U24640 ( .A(n16284), .Z(n16285) );
  XNOR U24641 ( .A(n16255), .B(n16286), .Z(n16250) );
  XNOR U24642 ( .A(n16253), .B(n16256), .Z(n16286) );
  NAND U24643 ( .A(n16287), .B(n16288), .Z(n16256) );
  NAND U24644 ( .A(n16289), .B(n16290), .Z(n16288) );
  OR U24645 ( .A(n16291), .B(n16292), .Z(n16289) );
  NANDN U24646 ( .A(n16293), .B(n16291), .Z(n16287) );
  IV U24647 ( .A(n16292), .Z(n16293) );
  NAND U24648 ( .A(n16294), .B(n16295), .Z(n16253) );
  NAND U24649 ( .A(n16296), .B(n16297), .Z(n16295) );
  NANDN U24650 ( .A(n16298), .B(n16299), .Z(n16296) );
  NANDN U24651 ( .A(n16299), .B(n16298), .Z(n16294) );
  AND U24652 ( .A(n16300), .B(n16301), .Z(n16255) );
  NAND U24653 ( .A(n16302), .B(n16303), .Z(n16301) );
  OR U24654 ( .A(n16304), .B(n16305), .Z(n16302) );
  NANDN U24655 ( .A(n16306), .B(n16304), .Z(n16300) );
  XNOR U24656 ( .A(n16281), .B(n16307), .Z(N63947) );
  XOR U24657 ( .A(n16283), .B(n16284), .Z(n16307) );
  XNOR U24658 ( .A(n16297), .B(n16308), .Z(n16284) );
  XOR U24659 ( .A(n16298), .B(n16299), .Z(n16308) );
  XOR U24660 ( .A(n16304), .B(n16309), .Z(n16299) );
  XOR U24661 ( .A(n16303), .B(n16306), .Z(n16309) );
  IV U24662 ( .A(n16305), .Z(n16306) );
  NAND U24663 ( .A(n16310), .B(n16311), .Z(n16305) );
  OR U24664 ( .A(n16312), .B(n16313), .Z(n16311) );
  OR U24665 ( .A(n16314), .B(n16315), .Z(n16310) );
  NAND U24666 ( .A(n16316), .B(n16317), .Z(n16303) );
  OR U24667 ( .A(n16318), .B(n16319), .Z(n16317) );
  OR U24668 ( .A(n16320), .B(n16321), .Z(n16316) );
  NOR U24669 ( .A(n16322), .B(n16323), .Z(n16304) );
  ANDN U24670 ( .B(n16324), .A(n16325), .Z(n16298) );
  XNOR U24671 ( .A(n16291), .B(n16326), .Z(n16297) );
  XNOR U24672 ( .A(n16290), .B(n16292), .Z(n16326) );
  NAND U24673 ( .A(n16327), .B(n16328), .Z(n16292) );
  OR U24674 ( .A(n16329), .B(n16330), .Z(n16328) );
  OR U24675 ( .A(n16331), .B(n16332), .Z(n16327) );
  NAND U24676 ( .A(n16333), .B(n16334), .Z(n16290) );
  OR U24677 ( .A(n16335), .B(n16336), .Z(n16334) );
  OR U24678 ( .A(n16337), .B(n16338), .Z(n16333) );
  ANDN U24679 ( .B(n16339), .A(n16340), .Z(n16291) );
  IV U24680 ( .A(n16341), .Z(n16339) );
  ANDN U24681 ( .B(n16342), .A(n16343), .Z(n16283) );
  XOR U24682 ( .A(n16269), .B(n16344), .Z(n16281) );
  XOR U24683 ( .A(n16270), .B(n16271), .Z(n16344) );
  XOR U24684 ( .A(n16276), .B(n16345), .Z(n16271) );
  XOR U24685 ( .A(n16275), .B(n16278), .Z(n16345) );
  IV U24686 ( .A(n16277), .Z(n16278) );
  NAND U24687 ( .A(n16346), .B(n16347), .Z(n16277) );
  OR U24688 ( .A(n16348), .B(n16349), .Z(n16347) );
  OR U24689 ( .A(n16350), .B(n16351), .Z(n16346) );
  NAND U24690 ( .A(n16352), .B(n16353), .Z(n16275) );
  OR U24691 ( .A(n16354), .B(n16355), .Z(n16353) );
  OR U24692 ( .A(n16356), .B(n16357), .Z(n16352) );
  NOR U24693 ( .A(n16358), .B(n16359), .Z(n16276) );
  ANDN U24694 ( .B(n16360), .A(n16361), .Z(n16270) );
  IV U24695 ( .A(n16362), .Z(n16360) );
  XNOR U24696 ( .A(n16263), .B(n16363), .Z(n16269) );
  XNOR U24697 ( .A(n16262), .B(n16264), .Z(n16363) );
  NAND U24698 ( .A(n16364), .B(n16365), .Z(n16264) );
  OR U24699 ( .A(n16366), .B(n16367), .Z(n16365) );
  OR U24700 ( .A(n16368), .B(n16369), .Z(n16364) );
  NAND U24701 ( .A(n16370), .B(n16371), .Z(n16262) );
  OR U24702 ( .A(n16372), .B(n16373), .Z(n16371) );
  OR U24703 ( .A(n16374), .B(n16375), .Z(n16370) );
  ANDN U24704 ( .B(n16376), .A(n16377), .Z(n16263) );
  IV U24705 ( .A(n16378), .Z(n16376) );
  XNOR U24706 ( .A(n16343), .B(n16342), .Z(N63946) );
  XOR U24707 ( .A(n16362), .B(n16361), .Z(n16342) );
  XNOR U24708 ( .A(n16377), .B(n16378), .Z(n16361) );
  XNOR U24709 ( .A(n16372), .B(n16373), .Z(n16378) );
  XNOR U24710 ( .A(n16374), .B(n16375), .Z(n16373) );
  XNOR U24711 ( .A(y[6205]), .B(x[6205]), .Z(n16375) );
  XNOR U24712 ( .A(y[6206]), .B(x[6206]), .Z(n16374) );
  XNOR U24713 ( .A(y[6204]), .B(x[6204]), .Z(n16372) );
  XNOR U24714 ( .A(n16366), .B(n16367), .Z(n16377) );
  XNOR U24715 ( .A(y[6201]), .B(x[6201]), .Z(n16367) );
  XNOR U24716 ( .A(n16368), .B(n16369), .Z(n16366) );
  XNOR U24717 ( .A(y[6202]), .B(x[6202]), .Z(n16369) );
  XNOR U24718 ( .A(y[6203]), .B(x[6203]), .Z(n16368) );
  XNOR U24719 ( .A(n16359), .B(n16358), .Z(n16362) );
  XNOR U24720 ( .A(n16354), .B(n16355), .Z(n16358) );
  XNOR U24721 ( .A(y[6198]), .B(x[6198]), .Z(n16355) );
  XNOR U24722 ( .A(n16356), .B(n16357), .Z(n16354) );
  XNOR U24723 ( .A(y[6199]), .B(x[6199]), .Z(n16357) );
  XNOR U24724 ( .A(y[6200]), .B(x[6200]), .Z(n16356) );
  XNOR U24725 ( .A(n16348), .B(n16349), .Z(n16359) );
  XNOR U24726 ( .A(y[6195]), .B(x[6195]), .Z(n16349) );
  XNOR U24727 ( .A(n16350), .B(n16351), .Z(n16348) );
  XNOR U24728 ( .A(y[6196]), .B(x[6196]), .Z(n16351) );
  XNOR U24729 ( .A(y[6197]), .B(x[6197]), .Z(n16350) );
  XOR U24730 ( .A(n16324), .B(n16325), .Z(n16343) );
  XNOR U24731 ( .A(n16340), .B(n16341), .Z(n16325) );
  XNOR U24732 ( .A(n16335), .B(n16336), .Z(n16341) );
  XNOR U24733 ( .A(n16337), .B(n16338), .Z(n16336) );
  XNOR U24734 ( .A(y[6193]), .B(x[6193]), .Z(n16338) );
  XNOR U24735 ( .A(y[6194]), .B(x[6194]), .Z(n16337) );
  XNOR U24736 ( .A(y[6192]), .B(x[6192]), .Z(n16335) );
  XNOR U24737 ( .A(n16329), .B(n16330), .Z(n16340) );
  XNOR U24738 ( .A(y[6189]), .B(x[6189]), .Z(n16330) );
  XNOR U24739 ( .A(n16331), .B(n16332), .Z(n16329) );
  XNOR U24740 ( .A(y[6190]), .B(x[6190]), .Z(n16332) );
  XNOR U24741 ( .A(y[6191]), .B(x[6191]), .Z(n16331) );
  XOR U24742 ( .A(n16323), .B(n16322), .Z(n16324) );
  XNOR U24743 ( .A(n16318), .B(n16319), .Z(n16322) );
  XNOR U24744 ( .A(y[6186]), .B(x[6186]), .Z(n16319) );
  XNOR U24745 ( .A(n16320), .B(n16321), .Z(n16318) );
  XNOR U24746 ( .A(y[6187]), .B(x[6187]), .Z(n16321) );
  XNOR U24747 ( .A(y[6188]), .B(x[6188]), .Z(n16320) );
  XNOR U24748 ( .A(n16312), .B(n16313), .Z(n16323) );
  XNOR U24749 ( .A(y[6183]), .B(x[6183]), .Z(n16313) );
  XNOR U24750 ( .A(n16314), .B(n16315), .Z(n16312) );
  XNOR U24751 ( .A(y[6184]), .B(x[6184]), .Z(n16315) );
  XNOR U24752 ( .A(y[6185]), .B(x[6185]), .Z(n16314) );
  NAND U24753 ( .A(n16379), .B(n16380), .Z(N63937) );
  NANDN U24754 ( .A(n16381), .B(n16382), .Z(n16380) );
  OR U24755 ( .A(n16383), .B(n16384), .Z(n16382) );
  NAND U24756 ( .A(n16383), .B(n16384), .Z(n16379) );
  XOR U24757 ( .A(n16383), .B(n16385), .Z(N63936) );
  XNOR U24758 ( .A(n16381), .B(n16384), .Z(n16385) );
  AND U24759 ( .A(n16386), .B(n16387), .Z(n16384) );
  NANDN U24760 ( .A(n16388), .B(n16389), .Z(n16387) );
  NANDN U24761 ( .A(n16390), .B(n16391), .Z(n16389) );
  NANDN U24762 ( .A(n16391), .B(n16390), .Z(n16386) );
  NAND U24763 ( .A(n16392), .B(n16393), .Z(n16381) );
  NANDN U24764 ( .A(n16394), .B(n16395), .Z(n16393) );
  OR U24765 ( .A(n16396), .B(n16397), .Z(n16395) );
  NAND U24766 ( .A(n16397), .B(n16396), .Z(n16392) );
  AND U24767 ( .A(n16398), .B(n16399), .Z(n16383) );
  NANDN U24768 ( .A(n16400), .B(n16401), .Z(n16399) );
  NANDN U24769 ( .A(n16402), .B(n16403), .Z(n16401) );
  NANDN U24770 ( .A(n16403), .B(n16402), .Z(n16398) );
  XOR U24771 ( .A(n16397), .B(n16404), .Z(N63935) );
  XOR U24772 ( .A(n16394), .B(n16396), .Z(n16404) );
  XNOR U24773 ( .A(n16390), .B(n16405), .Z(n16396) );
  XNOR U24774 ( .A(n16388), .B(n16391), .Z(n16405) );
  NAND U24775 ( .A(n16406), .B(n16407), .Z(n16391) );
  NAND U24776 ( .A(n16408), .B(n16409), .Z(n16407) );
  OR U24777 ( .A(n16410), .B(n16411), .Z(n16408) );
  NANDN U24778 ( .A(n16412), .B(n16410), .Z(n16406) );
  IV U24779 ( .A(n16411), .Z(n16412) );
  NAND U24780 ( .A(n16413), .B(n16414), .Z(n16388) );
  NAND U24781 ( .A(n16415), .B(n16416), .Z(n16414) );
  NANDN U24782 ( .A(n16417), .B(n16418), .Z(n16415) );
  NANDN U24783 ( .A(n16418), .B(n16417), .Z(n16413) );
  AND U24784 ( .A(n16419), .B(n16420), .Z(n16390) );
  NAND U24785 ( .A(n16421), .B(n16422), .Z(n16420) );
  OR U24786 ( .A(n16423), .B(n16424), .Z(n16421) );
  NANDN U24787 ( .A(n16425), .B(n16423), .Z(n16419) );
  NAND U24788 ( .A(n16426), .B(n16427), .Z(n16394) );
  NANDN U24789 ( .A(n16428), .B(n16429), .Z(n16427) );
  OR U24790 ( .A(n16430), .B(n16431), .Z(n16429) );
  NANDN U24791 ( .A(n16432), .B(n16430), .Z(n16426) );
  IV U24792 ( .A(n16431), .Z(n16432) );
  XNOR U24793 ( .A(n16402), .B(n16433), .Z(n16397) );
  XNOR U24794 ( .A(n16400), .B(n16403), .Z(n16433) );
  NAND U24795 ( .A(n16434), .B(n16435), .Z(n16403) );
  NAND U24796 ( .A(n16436), .B(n16437), .Z(n16435) );
  OR U24797 ( .A(n16438), .B(n16439), .Z(n16436) );
  NANDN U24798 ( .A(n16440), .B(n16438), .Z(n16434) );
  IV U24799 ( .A(n16439), .Z(n16440) );
  NAND U24800 ( .A(n16441), .B(n16442), .Z(n16400) );
  NAND U24801 ( .A(n16443), .B(n16444), .Z(n16442) );
  NANDN U24802 ( .A(n16445), .B(n16446), .Z(n16443) );
  NANDN U24803 ( .A(n16446), .B(n16445), .Z(n16441) );
  AND U24804 ( .A(n16447), .B(n16448), .Z(n16402) );
  NAND U24805 ( .A(n16449), .B(n16450), .Z(n16448) );
  OR U24806 ( .A(n16451), .B(n16452), .Z(n16449) );
  NANDN U24807 ( .A(n16453), .B(n16451), .Z(n16447) );
  XNOR U24808 ( .A(n16428), .B(n16454), .Z(N63934) );
  XOR U24809 ( .A(n16430), .B(n16431), .Z(n16454) );
  XNOR U24810 ( .A(n16444), .B(n16455), .Z(n16431) );
  XOR U24811 ( .A(n16445), .B(n16446), .Z(n16455) );
  XOR U24812 ( .A(n16451), .B(n16456), .Z(n16446) );
  XOR U24813 ( .A(n16450), .B(n16453), .Z(n16456) );
  IV U24814 ( .A(n16452), .Z(n16453) );
  NAND U24815 ( .A(n16457), .B(n16458), .Z(n16452) );
  OR U24816 ( .A(n16459), .B(n16460), .Z(n16458) );
  OR U24817 ( .A(n16461), .B(n16462), .Z(n16457) );
  NAND U24818 ( .A(n16463), .B(n16464), .Z(n16450) );
  OR U24819 ( .A(n16465), .B(n16466), .Z(n16464) );
  OR U24820 ( .A(n16467), .B(n16468), .Z(n16463) );
  NOR U24821 ( .A(n16469), .B(n16470), .Z(n16451) );
  ANDN U24822 ( .B(n16471), .A(n16472), .Z(n16445) );
  XNOR U24823 ( .A(n16438), .B(n16473), .Z(n16444) );
  XNOR U24824 ( .A(n16437), .B(n16439), .Z(n16473) );
  NAND U24825 ( .A(n16474), .B(n16475), .Z(n16439) );
  OR U24826 ( .A(n16476), .B(n16477), .Z(n16475) );
  OR U24827 ( .A(n16478), .B(n16479), .Z(n16474) );
  NAND U24828 ( .A(n16480), .B(n16481), .Z(n16437) );
  OR U24829 ( .A(n16482), .B(n16483), .Z(n16481) );
  OR U24830 ( .A(n16484), .B(n16485), .Z(n16480) );
  ANDN U24831 ( .B(n16486), .A(n16487), .Z(n16438) );
  IV U24832 ( .A(n16488), .Z(n16486) );
  ANDN U24833 ( .B(n16489), .A(n16490), .Z(n16430) );
  XOR U24834 ( .A(n16416), .B(n16491), .Z(n16428) );
  XOR U24835 ( .A(n16417), .B(n16418), .Z(n16491) );
  XOR U24836 ( .A(n16423), .B(n16492), .Z(n16418) );
  XOR U24837 ( .A(n16422), .B(n16425), .Z(n16492) );
  IV U24838 ( .A(n16424), .Z(n16425) );
  NAND U24839 ( .A(n16493), .B(n16494), .Z(n16424) );
  OR U24840 ( .A(n16495), .B(n16496), .Z(n16494) );
  OR U24841 ( .A(n16497), .B(n16498), .Z(n16493) );
  NAND U24842 ( .A(n16499), .B(n16500), .Z(n16422) );
  OR U24843 ( .A(n16501), .B(n16502), .Z(n16500) );
  OR U24844 ( .A(n16503), .B(n16504), .Z(n16499) );
  NOR U24845 ( .A(n16505), .B(n16506), .Z(n16423) );
  ANDN U24846 ( .B(n16507), .A(n16508), .Z(n16417) );
  IV U24847 ( .A(n16509), .Z(n16507) );
  XNOR U24848 ( .A(n16410), .B(n16510), .Z(n16416) );
  XNOR U24849 ( .A(n16409), .B(n16411), .Z(n16510) );
  NAND U24850 ( .A(n16511), .B(n16512), .Z(n16411) );
  OR U24851 ( .A(n16513), .B(n16514), .Z(n16512) );
  OR U24852 ( .A(n16515), .B(n16516), .Z(n16511) );
  NAND U24853 ( .A(n16517), .B(n16518), .Z(n16409) );
  OR U24854 ( .A(n16519), .B(n16520), .Z(n16518) );
  OR U24855 ( .A(n16521), .B(n16522), .Z(n16517) );
  ANDN U24856 ( .B(n16523), .A(n16524), .Z(n16410) );
  IV U24857 ( .A(n16525), .Z(n16523) );
  XNOR U24858 ( .A(n16490), .B(n16489), .Z(N63933) );
  XOR U24859 ( .A(n16509), .B(n16508), .Z(n16489) );
  XNOR U24860 ( .A(n16524), .B(n16525), .Z(n16508) );
  XNOR U24861 ( .A(n16519), .B(n16520), .Z(n16525) );
  XNOR U24862 ( .A(n16521), .B(n16522), .Z(n16520) );
  XNOR U24863 ( .A(y[6181]), .B(x[6181]), .Z(n16522) );
  XNOR U24864 ( .A(y[6182]), .B(x[6182]), .Z(n16521) );
  XNOR U24865 ( .A(y[6180]), .B(x[6180]), .Z(n16519) );
  XNOR U24866 ( .A(n16513), .B(n16514), .Z(n16524) );
  XNOR U24867 ( .A(y[6177]), .B(x[6177]), .Z(n16514) );
  XNOR U24868 ( .A(n16515), .B(n16516), .Z(n16513) );
  XNOR U24869 ( .A(y[6178]), .B(x[6178]), .Z(n16516) );
  XNOR U24870 ( .A(y[6179]), .B(x[6179]), .Z(n16515) );
  XNOR U24871 ( .A(n16506), .B(n16505), .Z(n16509) );
  XNOR U24872 ( .A(n16501), .B(n16502), .Z(n16505) );
  XNOR U24873 ( .A(y[6174]), .B(x[6174]), .Z(n16502) );
  XNOR U24874 ( .A(n16503), .B(n16504), .Z(n16501) );
  XNOR U24875 ( .A(y[6175]), .B(x[6175]), .Z(n16504) );
  XNOR U24876 ( .A(y[6176]), .B(x[6176]), .Z(n16503) );
  XNOR U24877 ( .A(n16495), .B(n16496), .Z(n16506) );
  XNOR U24878 ( .A(y[6171]), .B(x[6171]), .Z(n16496) );
  XNOR U24879 ( .A(n16497), .B(n16498), .Z(n16495) );
  XNOR U24880 ( .A(y[6172]), .B(x[6172]), .Z(n16498) );
  XNOR U24881 ( .A(y[6173]), .B(x[6173]), .Z(n16497) );
  XOR U24882 ( .A(n16471), .B(n16472), .Z(n16490) );
  XNOR U24883 ( .A(n16487), .B(n16488), .Z(n16472) );
  XNOR U24884 ( .A(n16482), .B(n16483), .Z(n16488) );
  XNOR U24885 ( .A(n16484), .B(n16485), .Z(n16483) );
  XNOR U24886 ( .A(y[6169]), .B(x[6169]), .Z(n16485) );
  XNOR U24887 ( .A(y[6170]), .B(x[6170]), .Z(n16484) );
  XNOR U24888 ( .A(y[6168]), .B(x[6168]), .Z(n16482) );
  XNOR U24889 ( .A(n16476), .B(n16477), .Z(n16487) );
  XNOR U24890 ( .A(y[6165]), .B(x[6165]), .Z(n16477) );
  XNOR U24891 ( .A(n16478), .B(n16479), .Z(n16476) );
  XNOR U24892 ( .A(y[6166]), .B(x[6166]), .Z(n16479) );
  XNOR U24893 ( .A(y[6167]), .B(x[6167]), .Z(n16478) );
  XOR U24894 ( .A(n16470), .B(n16469), .Z(n16471) );
  XNOR U24895 ( .A(n16465), .B(n16466), .Z(n16469) );
  XNOR U24896 ( .A(y[6162]), .B(x[6162]), .Z(n16466) );
  XNOR U24897 ( .A(n16467), .B(n16468), .Z(n16465) );
  XNOR U24898 ( .A(y[6163]), .B(x[6163]), .Z(n16468) );
  XNOR U24899 ( .A(y[6164]), .B(x[6164]), .Z(n16467) );
  XNOR U24900 ( .A(n16459), .B(n16460), .Z(n16470) );
  XNOR U24901 ( .A(y[6159]), .B(x[6159]), .Z(n16460) );
  XNOR U24902 ( .A(n16461), .B(n16462), .Z(n16459) );
  XNOR U24903 ( .A(y[6160]), .B(x[6160]), .Z(n16462) );
  XNOR U24904 ( .A(y[6161]), .B(x[6161]), .Z(n16461) );
  NAND U24905 ( .A(n16526), .B(n16527), .Z(N63924) );
  NANDN U24906 ( .A(n16528), .B(n16529), .Z(n16527) );
  OR U24907 ( .A(n16530), .B(n16531), .Z(n16529) );
  NAND U24908 ( .A(n16530), .B(n16531), .Z(n16526) );
  XOR U24909 ( .A(n16530), .B(n16532), .Z(N63923) );
  XNOR U24910 ( .A(n16528), .B(n16531), .Z(n16532) );
  AND U24911 ( .A(n16533), .B(n16534), .Z(n16531) );
  NANDN U24912 ( .A(n16535), .B(n16536), .Z(n16534) );
  NANDN U24913 ( .A(n16537), .B(n16538), .Z(n16536) );
  NANDN U24914 ( .A(n16538), .B(n16537), .Z(n16533) );
  NAND U24915 ( .A(n16539), .B(n16540), .Z(n16528) );
  NANDN U24916 ( .A(n16541), .B(n16542), .Z(n16540) );
  OR U24917 ( .A(n16543), .B(n16544), .Z(n16542) );
  NAND U24918 ( .A(n16544), .B(n16543), .Z(n16539) );
  AND U24919 ( .A(n16545), .B(n16546), .Z(n16530) );
  NANDN U24920 ( .A(n16547), .B(n16548), .Z(n16546) );
  NANDN U24921 ( .A(n16549), .B(n16550), .Z(n16548) );
  NANDN U24922 ( .A(n16550), .B(n16549), .Z(n16545) );
  XOR U24923 ( .A(n16544), .B(n16551), .Z(N63922) );
  XOR U24924 ( .A(n16541), .B(n16543), .Z(n16551) );
  XNOR U24925 ( .A(n16537), .B(n16552), .Z(n16543) );
  XNOR U24926 ( .A(n16535), .B(n16538), .Z(n16552) );
  NAND U24927 ( .A(n16553), .B(n16554), .Z(n16538) );
  NAND U24928 ( .A(n16555), .B(n16556), .Z(n16554) );
  OR U24929 ( .A(n16557), .B(n16558), .Z(n16555) );
  NANDN U24930 ( .A(n16559), .B(n16557), .Z(n16553) );
  IV U24931 ( .A(n16558), .Z(n16559) );
  NAND U24932 ( .A(n16560), .B(n16561), .Z(n16535) );
  NAND U24933 ( .A(n16562), .B(n16563), .Z(n16561) );
  NANDN U24934 ( .A(n16564), .B(n16565), .Z(n16562) );
  NANDN U24935 ( .A(n16565), .B(n16564), .Z(n16560) );
  AND U24936 ( .A(n16566), .B(n16567), .Z(n16537) );
  NAND U24937 ( .A(n16568), .B(n16569), .Z(n16567) );
  OR U24938 ( .A(n16570), .B(n16571), .Z(n16568) );
  NANDN U24939 ( .A(n16572), .B(n16570), .Z(n16566) );
  NAND U24940 ( .A(n16573), .B(n16574), .Z(n16541) );
  NANDN U24941 ( .A(n16575), .B(n16576), .Z(n16574) );
  OR U24942 ( .A(n16577), .B(n16578), .Z(n16576) );
  NANDN U24943 ( .A(n16579), .B(n16577), .Z(n16573) );
  IV U24944 ( .A(n16578), .Z(n16579) );
  XNOR U24945 ( .A(n16549), .B(n16580), .Z(n16544) );
  XNOR U24946 ( .A(n16547), .B(n16550), .Z(n16580) );
  NAND U24947 ( .A(n16581), .B(n16582), .Z(n16550) );
  NAND U24948 ( .A(n16583), .B(n16584), .Z(n16582) );
  OR U24949 ( .A(n16585), .B(n16586), .Z(n16583) );
  NANDN U24950 ( .A(n16587), .B(n16585), .Z(n16581) );
  IV U24951 ( .A(n16586), .Z(n16587) );
  NAND U24952 ( .A(n16588), .B(n16589), .Z(n16547) );
  NAND U24953 ( .A(n16590), .B(n16591), .Z(n16589) );
  NANDN U24954 ( .A(n16592), .B(n16593), .Z(n16590) );
  NANDN U24955 ( .A(n16593), .B(n16592), .Z(n16588) );
  AND U24956 ( .A(n16594), .B(n16595), .Z(n16549) );
  NAND U24957 ( .A(n16596), .B(n16597), .Z(n16595) );
  OR U24958 ( .A(n16598), .B(n16599), .Z(n16596) );
  NANDN U24959 ( .A(n16600), .B(n16598), .Z(n16594) );
  XNOR U24960 ( .A(n16575), .B(n16601), .Z(N63921) );
  XOR U24961 ( .A(n16577), .B(n16578), .Z(n16601) );
  XNOR U24962 ( .A(n16591), .B(n16602), .Z(n16578) );
  XOR U24963 ( .A(n16592), .B(n16593), .Z(n16602) );
  XOR U24964 ( .A(n16598), .B(n16603), .Z(n16593) );
  XOR U24965 ( .A(n16597), .B(n16600), .Z(n16603) );
  IV U24966 ( .A(n16599), .Z(n16600) );
  NAND U24967 ( .A(n16604), .B(n16605), .Z(n16599) );
  OR U24968 ( .A(n16606), .B(n16607), .Z(n16605) );
  OR U24969 ( .A(n16608), .B(n16609), .Z(n16604) );
  NAND U24970 ( .A(n16610), .B(n16611), .Z(n16597) );
  OR U24971 ( .A(n16612), .B(n16613), .Z(n16611) );
  OR U24972 ( .A(n16614), .B(n16615), .Z(n16610) );
  NOR U24973 ( .A(n16616), .B(n16617), .Z(n16598) );
  ANDN U24974 ( .B(n16618), .A(n16619), .Z(n16592) );
  XNOR U24975 ( .A(n16585), .B(n16620), .Z(n16591) );
  XNOR U24976 ( .A(n16584), .B(n16586), .Z(n16620) );
  NAND U24977 ( .A(n16621), .B(n16622), .Z(n16586) );
  OR U24978 ( .A(n16623), .B(n16624), .Z(n16622) );
  OR U24979 ( .A(n16625), .B(n16626), .Z(n16621) );
  NAND U24980 ( .A(n16627), .B(n16628), .Z(n16584) );
  OR U24981 ( .A(n16629), .B(n16630), .Z(n16628) );
  OR U24982 ( .A(n16631), .B(n16632), .Z(n16627) );
  ANDN U24983 ( .B(n16633), .A(n16634), .Z(n16585) );
  IV U24984 ( .A(n16635), .Z(n16633) );
  ANDN U24985 ( .B(n16636), .A(n16637), .Z(n16577) );
  XOR U24986 ( .A(n16563), .B(n16638), .Z(n16575) );
  XOR U24987 ( .A(n16564), .B(n16565), .Z(n16638) );
  XOR U24988 ( .A(n16570), .B(n16639), .Z(n16565) );
  XOR U24989 ( .A(n16569), .B(n16572), .Z(n16639) );
  IV U24990 ( .A(n16571), .Z(n16572) );
  NAND U24991 ( .A(n16640), .B(n16641), .Z(n16571) );
  OR U24992 ( .A(n16642), .B(n16643), .Z(n16641) );
  OR U24993 ( .A(n16644), .B(n16645), .Z(n16640) );
  NAND U24994 ( .A(n16646), .B(n16647), .Z(n16569) );
  OR U24995 ( .A(n16648), .B(n16649), .Z(n16647) );
  OR U24996 ( .A(n16650), .B(n16651), .Z(n16646) );
  NOR U24997 ( .A(n16652), .B(n16653), .Z(n16570) );
  ANDN U24998 ( .B(n16654), .A(n16655), .Z(n16564) );
  IV U24999 ( .A(n16656), .Z(n16654) );
  XNOR U25000 ( .A(n16557), .B(n16657), .Z(n16563) );
  XNOR U25001 ( .A(n16556), .B(n16558), .Z(n16657) );
  NAND U25002 ( .A(n16658), .B(n16659), .Z(n16558) );
  OR U25003 ( .A(n16660), .B(n16661), .Z(n16659) );
  OR U25004 ( .A(n16662), .B(n16663), .Z(n16658) );
  NAND U25005 ( .A(n16664), .B(n16665), .Z(n16556) );
  OR U25006 ( .A(n16666), .B(n16667), .Z(n16665) );
  OR U25007 ( .A(n16668), .B(n16669), .Z(n16664) );
  ANDN U25008 ( .B(n16670), .A(n16671), .Z(n16557) );
  IV U25009 ( .A(n16672), .Z(n16670) );
  XNOR U25010 ( .A(n16637), .B(n16636), .Z(N63920) );
  XOR U25011 ( .A(n16656), .B(n16655), .Z(n16636) );
  XNOR U25012 ( .A(n16671), .B(n16672), .Z(n16655) );
  XNOR U25013 ( .A(n16666), .B(n16667), .Z(n16672) );
  XNOR U25014 ( .A(n16668), .B(n16669), .Z(n16667) );
  XNOR U25015 ( .A(y[6157]), .B(x[6157]), .Z(n16669) );
  XNOR U25016 ( .A(y[6158]), .B(x[6158]), .Z(n16668) );
  XNOR U25017 ( .A(y[6156]), .B(x[6156]), .Z(n16666) );
  XNOR U25018 ( .A(n16660), .B(n16661), .Z(n16671) );
  XNOR U25019 ( .A(y[6153]), .B(x[6153]), .Z(n16661) );
  XNOR U25020 ( .A(n16662), .B(n16663), .Z(n16660) );
  XNOR U25021 ( .A(y[6154]), .B(x[6154]), .Z(n16663) );
  XNOR U25022 ( .A(y[6155]), .B(x[6155]), .Z(n16662) );
  XNOR U25023 ( .A(n16653), .B(n16652), .Z(n16656) );
  XNOR U25024 ( .A(n16648), .B(n16649), .Z(n16652) );
  XNOR U25025 ( .A(y[6150]), .B(x[6150]), .Z(n16649) );
  XNOR U25026 ( .A(n16650), .B(n16651), .Z(n16648) );
  XNOR U25027 ( .A(y[6151]), .B(x[6151]), .Z(n16651) );
  XNOR U25028 ( .A(y[6152]), .B(x[6152]), .Z(n16650) );
  XNOR U25029 ( .A(n16642), .B(n16643), .Z(n16653) );
  XNOR U25030 ( .A(y[6147]), .B(x[6147]), .Z(n16643) );
  XNOR U25031 ( .A(n16644), .B(n16645), .Z(n16642) );
  XNOR U25032 ( .A(y[6148]), .B(x[6148]), .Z(n16645) );
  XNOR U25033 ( .A(y[6149]), .B(x[6149]), .Z(n16644) );
  XOR U25034 ( .A(n16618), .B(n16619), .Z(n16637) );
  XNOR U25035 ( .A(n16634), .B(n16635), .Z(n16619) );
  XNOR U25036 ( .A(n16629), .B(n16630), .Z(n16635) );
  XNOR U25037 ( .A(n16631), .B(n16632), .Z(n16630) );
  XNOR U25038 ( .A(y[6145]), .B(x[6145]), .Z(n16632) );
  XNOR U25039 ( .A(y[6146]), .B(x[6146]), .Z(n16631) );
  XNOR U25040 ( .A(y[6144]), .B(x[6144]), .Z(n16629) );
  XNOR U25041 ( .A(n16623), .B(n16624), .Z(n16634) );
  XNOR U25042 ( .A(y[6141]), .B(x[6141]), .Z(n16624) );
  XNOR U25043 ( .A(n16625), .B(n16626), .Z(n16623) );
  XNOR U25044 ( .A(y[6142]), .B(x[6142]), .Z(n16626) );
  XNOR U25045 ( .A(y[6143]), .B(x[6143]), .Z(n16625) );
  XOR U25046 ( .A(n16617), .B(n16616), .Z(n16618) );
  XNOR U25047 ( .A(n16612), .B(n16613), .Z(n16616) );
  XNOR U25048 ( .A(y[6138]), .B(x[6138]), .Z(n16613) );
  XNOR U25049 ( .A(n16614), .B(n16615), .Z(n16612) );
  XNOR U25050 ( .A(y[6139]), .B(x[6139]), .Z(n16615) );
  XNOR U25051 ( .A(y[6140]), .B(x[6140]), .Z(n16614) );
  XNOR U25052 ( .A(n16606), .B(n16607), .Z(n16617) );
  XNOR U25053 ( .A(y[6135]), .B(x[6135]), .Z(n16607) );
  XNOR U25054 ( .A(n16608), .B(n16609), .Z(n16606) );
  XNOR U25055 ( .A(y[6136]), .B(x[6136]), .Z(n16609) );
  XNOR U25056 ( .A(y[6137]), .B(x[6137]), .Z(n16608) );
  NAND U25057 ( .A(n16673), .B(n16674), .Z(N63911) );
  NANDN U25058 ( .A(n16675), .B(n16676), .Z(n16674) );
  OR U25059 ( .A(n16677), .B(n16678), .Z(n16676) );
  NAND U25060 ( .A(n16677), .B(n16678), .Z(n16673) );
  XOR U25061 ( .A(n16677), .B(n16679), .Z(N63910) );
  XNOR U25062 ( .A(n16675), .B(n16678), .Z(n16679) );
  AND U25063 ( .A(n16680), .B(n16681), .Z(n16678) );
  NANDN U25064 ( .A(n16682), .B(n16683), .Z(n16681) );
  NANDN U25065 ( .A(n16684), .B(n16685), .Z(n16683) );
  NANDN U25066 ( .A(n16685), .B(n16684), .Z(n16680) );
  NAND U25067 ( .A(n16686), .B(n16687), .Z(n16675) );
  NANDN U25068 ( .A(n16688), .B(n16689), .Z(n16687) );
  OR U25069 ( .A(n16690), .B(n16691), .Z(n16689) );
  NAND U25070 ( .A(n16691), .B(n16690), .Z(n16686) );
  AND U25071 ( .A(n16692), .B(n16693), .Z(n16677) );
  NANDN U25072 ( .A(n16694), .B(n16695), .Z(n16693) );
  NANDN U25073 ( .A(n16696), .B(n16697), .Z(n16695) );
  NANDN U25074 ( .A(n16697), .B(n16696), .Z(n16692) );
  XOR U25075 ( .A(n16691), .B(n16698), .Z(N63909) );
  XOR U25076 ( .A(n16688), .B(n16690), .Z(n16698) );
  XNOR U25077 ( .A(n16684), .B(n16699), .Z(n16690) );
  XNOR U25078 ( .A(n16682), .B(n16685), .Z(n16699) );
  NAND U25079 ( .A(n16700), .B(n16701), .Z(n16685) );
  NAND U25080 ( .A(n16702), .B(n16703), .Z(n16701) );
  OR U25081 ( .A(n16704), .B(n16705), .Z(n16702) );
  NANDN U25082 ( .A(n16706), .B(n16704), .Z(n16700) );
  IV U25083 ( .A(n16705), .Z(n16706) );
  NAND U25084 ( .A(n16707), .B(n16708), .Z(n16682) );
  NAND U25085 ( .A(n16709), .B(n16710), .Z(n16708) );
  NANDN U25086 ( .A(n16711), .B(n16712), .Z(n16709) );
  NANDN U25087 ( .A(n16712), .B(n16711), .Z(n16707) );
  AND U25088 ( .A(n16713), .B(n16714), .Z(n16684) );
  NAND U25089 ( .A(n16715), .B(n16716), .Z(n16714) );
  OR U25090 ( .A(n16717), .B(n16718), .Z(n16715) );
  NANDN U25091 ( .A(n16719), .B(n16717), .Z(n16713) );
  NAND U25092 ( .A(n16720), .B(n16721), .Z(n16688) );
  NANDN U25093 ( .A(n16722), .B(n16723), .Z(n16721) );
  OR U25094 ( .A(n16724), .B(n16725), .Z(n16723) );
  NANDN U25095 ( .A(n16726), .B(n16724), .Z(n16720) );
  IV U25096 ( .A(n16725), .Z(n16726) );
  XNOR U25097 ( .A(n16696), .B(n16727), .Z(n16691) );
  XNOR U25098 ( .A(n16694), .B(n16697), .Z(n16727) );
  NAND U25099 ( .A(n16728), .B(n16729), .Z(n16697) );
  NAND U25100 ( .A(n16730), .B(n16731), .Z(n16729) );
  OR U25101 ( .A(n16732), .B(n16733), .Z(n16730) );
  NANDN U25102 ( .A(n16734), .B(n16732), .Z(n16728) );
  IV U25103 ( .A(n16733), .Z(n16734) );
  NAND U25104 ( .A(n16735), .B(n16736), .Z(n16694) );
  NAND U25105 ( .A(n16737), .B(n16738), .Z(n16736) );
  NANDN U25106 ( .A(n16739), .B(n16740), .Z(n16737) );
  NANDN U25107 ( .A(n16740), .B(n16739), .Z(n16735) );
  AND U25108 ( .A(n16741), .B(n16742), .Z(n16696) );
  NAND U25109 ( .A(n16743), .B(n16744), .Z(n16742) );
  OR U25110 ( .A(n16745), .B(n16746), .Z(n16743) );
  NANDN U25111 ( .A(n16747), .B(n16745), .Z(n16741) );
  XNOR U25112 ( .A(n16722), .B(n16748), .Z(N63908) );
  XOR U25113 ( .A(n16724), .B(n16725), .Z(n16748) );
  XNOR U25114 ( .A(n16738), .B(n16749), .Z(n16725) );
  XOR U25115 ( .A(n16739), .B(n16740), .Z(n16749) );
  XOR U25116 ( .A(n16745), .B(n16750), .Z(n16740) );
  XOR U25117 ( .A(n16744), .B(n16747), .Z(n16750) );
  IV U25118 ( .A(n16746), .Z(n16747) );
  NAND U25119 ( .A(n16751), .B(n16752), .Z(n16746) );
  OR U25120 ( .A(n16753), .B(n16754), .Z(n16752) );
  OR U25121 ( .A(n16755), .B(n16756), .Z(n16751) );
  NAND U25122 ( .A(n16757), .B(n16758), .Z(n16744) );
  OR U25123 ( .A(n16759), .B(n16760), .Z(n16758) );
  OR U25124 ( .A(n16761), .B(n16762), .Z(n16757) );
  NOR U25125 ( .A(n16763), .B(n16764), .Z(n16745) );
  ANDN U25126 ( .B(n16765), .A(n16766), .Z(n16739) );
  XNOR U25127 ( .A(n16732), .B(n16767), .Z(n16738) );
  XNOR U25128 ( .A(n16731), .B(n16733), .Z(n16767) );
  NAND U25129 ( .A(n16768), .B(n16769), .Z(n16733) );
  OR U25130 ( .A(n16770), .B(n16771), .Z(n16769) );
  OR U25131 ( .A(n16772), .B(n16773), .Z(n16768) );
  NAND U25132 ( .A(n16774), .B(n16775), .Z(n16731) );
  OR U25133 ( .A(n16776), .B(n16777), .Z(n16775) );
  OR U25134 ( .A(n16778), .B(n16779), .Z(n16774) );
  ANDN U25135 ( .B(n16780), .A(n16781), .Z(n16732) );
  IV U25136 ( .A(n16782), .Z(n16780) );
  ANDN U25137 ( .B(n16783), .A(n16784), .Z(n16724) );
  XOR U25138 ( .A(n16710), .B(n16785), .Z(n16722) );
  XOR U25139 ( .A(n16711), .B(n16712), .Z(n16785) );
  XOR U25140 ( .A(n16717), .B(n16786), .Z(n16712) );
  XOR U25141 ( .A(n16716), .B(n16719), .Z(n16786) );
  IV U25142 ( .A(n16718), .Z(n16719) );
  NAND U25143 ( .A(n16787), .B(n16788), .Z(n16718) );
  OR U25144 ( .A(n16789), .B(n16790), .Z(n16788) );
  OR U25145 ( .A(n16791), .B(n16792), .Z(n16787) );
  NAND U25146 ( .A(n16793), .B(n16794), .Z(n16716) );
  OR U25147 ( .A(n16795), .B(n16796), .Z(n16794) );
  OR U25148 ( .A(n16797), .B(n16798), .Z(n16793) );
  NOR U25149 ( .A(n16799), .B(n16800), .Z(n16717) );
  ANDN U25150 ( .B(n16801), .A(n16802), .Z(n16711) );
  IV U25151 ( .A(n16803), .Z(n16801) );
  XNOR U25152 ( .A(n16704), .B(n16804), .Z(n16710) );
  XNOR U25153 ( .A(n16703), .B(n16705), .Z(n16804) );
  NAND U25154 ( .A(n16805), .B(n16806), .Z(n16705) );
  OR U25155 ( .A(n16807), .B(n16808), .Z(n16806) );
  OR U25156 ( .A(n16809), .B(n16810), .Z(n16805) );
  NAND U25157 ( .A(n16811), .B(n16812), .Z(n16703) );
  OR U25158 ( .A(n16813), .B(n16814), .Z(n16812) );
  OR U25159 ( .A(n16815), .B(n16816), .Z(n16811) );
  ANDN U25160 ( .B(n16817), .A(n16818), .Z(n16704) );
  IV U25161 ( .A(n16819), .Z(n16817) );
  XNOR U25162 ( .A(n16784), .B(n16783), .Z(N63907) );
  XOR U25163 ( .A(n16803), .B(n16802), .Z(n16783) );
  XNOR U25164 ( .A(n16818), .B(n16819), .Z(n16802) );
  XNOR U25165 ( .A(n16813), .B(n16814), .Z(n16819) );
  XNOR U25166 ( .A(n16815), .B(n16816), .Z(n16814) );
  XNOR U25167 ( .A(y[6133]), .B(x[6133]), .Z(n16816) );
  XNOR U25168 ( .A(y[6134]), .B(x[6134]), .Z(n16815) );
  XNOR U25169 ( .A(y[6132]), .B(x[6132]), .Z(n16813) );
  XNOR U25170 ( .A(n16807), .B(n16808), .Z(n16818) );
  XNOR U25171 ( .A(y[6129]), .B(x[6129]), .Z(n16808) );
  XNOR U25172 ( .A(n16809), .B(n16810), .Z(n16807) );
  XNOR U25173 ( .A(y[6130]), .B(x[6130]), .Z(n16810) );
  XNOR U25174 ( .A(y[6131]), .B(x[6131]), .Z(n16809) );
  XNOR U25175 ( .A(n16800), .B(n16799), .Z(n16803) );
  XNOR U25176 ( .A(n16795), .B(n16796), .Z(n16799) );
  XNOR U25177 ( .A(y[6126]), .B(x[6126]), .Z(n16796) );
  XNOR U25178 ( .A(n16797), .B(n16798), .Z(n16795) );
  XNOR U25179 ( .A(y[6127]), .B(x[6127]), .Z(n16798) );
  XNOR U25180 ( .A(y[6128]), .B(x[6128]), .Z(n16797) );
  XNOR U25181 ( .A(n16789), .B(n16790), .Z(n16800) );
  XNOR U25182 ( .A(y[6123]), .B(x[6123]), .Z(n16790) );
  XNOR U25183 ( .A(n16791), .B(n16792), .Z(n16789) );
  XNOR U25184 ( .A(y[6124]), .B(x[6124]), .Z(n16792) );
  XNOR U25185 ( .A(y[6125]), .B(x[6125]), .Z(n16791) );
  XOR U25186 ( .A(n16765), .B(n16766), .Z(n16784) );
  XNOR U25187 ( .A(n16781), .B(n16782), .Z(n16766) );
  XNOR U25188 ( .A(n16776), .B(n16777), .Z(n16782) );
  XNOR U25189 ( .A(n16778), .B(n16779), .Z(n16777) );
  XNOR U25190 ( .A(y[6121]), .B(x[6121]), .Z(n16779) );
  XNOR U25191 ( .A(y[6122]), .B(x[6122]), .Z(n16778) );
  XNOR U25192 ( .A(y[6120]), .B(x[6120]), .Z(n16776) );
  XNOR U25193 ( .A(n16770), .B(n16771), .Z(n16781) );
  XNOR U25194 ( .A(y[6117]), .B(x[6117]), .Z(n16771) );
  XNOR U25195 ( .A(n16772), .B(n16773), .Z(n16770) );
  XNOR U25196 ( .A(y[6118]), .B(x[6118]), .Z(n16773) );
  XNOR U25197 ( .A(y[6119]), .B(x[6119]), .Z(n16772) );
  XOR U25198 ( .A(n16764), .B(n16763), .Z(n16765) );
  XNOR U25199 ( .A(n16759), .B(n16760), .Z(n16763) );
  XNOR U25200 ( .A(y[6114]), .B(x[6114]), .Z(n16760) );
  XNOR U25201 ( .A(n16761), .B(n16762), .Z(n16759) );
  XNOR U25202 ( .A(y[6115]), .B(x[6115]), .Z(n16762) );
  XNOR U25203 ( .A(y[6116]), .B(x[6116]), .Z(n16761) );
  XNOR U25204 ( .A(n16753), .B(n16754), .Z(n16764) );
  XNOR U25205 ( .A(y[6111]), .B(x[6111]), .Z(n16754) );
  XNOR U25206 ( .A(n16755), .B(n16756), .Z(n16753) );
  XNOR U25207 ( .A(y[6112]), .B(x[6112]), .Z(n16756) );
  XNOR U25208 ( .A(y[6113]), .B(x[6113]), .Z(n16755) );
  NAND U25209 ( .A(n16820), .B(n16821), .Z(N63898) );
  NANDN U25210 ( .A(n16822), .B(n16823), .Z(n16821) );
  OR U25211 ( .A(n16824), .B(n16825), .Z(n16823) );
  NAND U25212 ( .A(n16824), .B(n16825), .Z(n16820) );
  XOR U25213 ( .A(n16824), .B(n16826), .Z(N63897) );
  XNOR U25214 ( .A(n16822), .B(n16825), .Z(n16826) );
  AND U25215 ( .A(n16827), .B(n16828), .Z(n16825) );
  NANDN U25216 ( .A(n16829), .B(n16830), .Z(n16828) );
  NANDN U25217 ( .A(n16831), .B(n16832), .Z(n16830) );
  NANDN U25218 ( .A(n16832), .B(n16831), .Z(n16827) );
  NAND U25219 ( .A(n16833), .B(n16834), .Z(n16822) );
  NANDN U25220 ( .A(n16835), .B(n16836), .Z(n16834) );
  OR U25221 ( .A(n16837), .B(n16838), .Z(n16836) );
  NAND U25222 ( .A(n16838), .B(n16837), .Z(n16833) );
  AND U25223 ( .A(n16839), .B(n16840), .Z(n16824) );
  NANDN U25224 ( .A(n16841), .B(n16842), .Z(n16840) );
  NANDN U25225 ( .A(n16843), .B(n16844), .Z(n16842) );
  NANDN U25226 ( .A(n16844), .B(n16843), .Z(n16839) );
  XOR U25227 ( .A(n16838), .B(n16845), .Z(N63896) );
  XOR U25228 ( .A(n16835), .B(n16837), .Z(n16845) );
  XNOR U25229 ( .A(n16831), .B(n16846), .Z(n16837) );
  XNOR U25230 ( .A(n16829), .B(n16832), .Z(n16846) );
  NAND U25231 ( .A(n16847), .B(n16848), .Z(n16832) );
  NAND U25232 ( .A(n16849), .B(n16850), .Z(n16848) );
  OR U25233 ( .A(n16851), .B(n16852), .Z(n16849) );
  NANDN U25234 ( .A(n16853), .B(n16851), .Z(n16847) );
  IV U25235 ( .A(n16852), .Z(n16853) );
  NAND U25236 ( .A(n16854), .B(n16855), .Z(n16829) );
  NAND U25237 ( .A(n16856), .B(n16857), .Z(n16855) );
  NANDN U25238 ( .A(n16858), .B(n16859), .Z(n16856) );
  NANDN U25239 ( .A(n16859), .B(n16858), .Z(n16854) );
  AND U25240 ( .A(n16860), .B(n16861), .Z(n16831) );
  NAND U25241 ( .A(n16862), .B(n16863), .Z(n16861) );
  OR U25242 ( .A(n16864), .B(n16865), .Z(n16862) );
  NANDN U25243 ( .A(n16866), .B(n16864), .Z(n16860) );
  NAND U25244 ( .A(n16867), .B(n16868), .Z(n16835) );
  NANDN U25245 ( .A(n16869), .B(n16870), .Z(n16868) );
  OR U25246 ( .A(n16871), .B(n16872), .Z(n16870) );
  NANDN U25247 ( .A(n16873), .B(n16871), .Z(n16867) );
  IV U25248 ( .A(n16872), .Z(n16873) );
  XNOR U25249 ( .A(n16843), .B(n16874), .Z(n16838) );
  XNOR U25250 ( .A(n16841), .B(n16844), .Z(n16874) );
  NAND U25251 ( .A(n16875), .B(n16876), .Z(n16844) );
  NAND U25252 ( .A(n16877), .B(n16878), .Z(n16876) );
  OR U25253 ( .A(n16879), .B(n16880), .Z(n16877) );
  NANDN U25254 ( .A(n16881), .B(n16879), .Z(n16875) );
  IV U25255 ( .A(n16880), .Z(n16881) );
  NAND U25256 ( .A(n16882), .B(n16883), .Z(n16841) );
  NAND U25257 ( .A(n16884), .B(n16885), .Z(n16883) );
  NANDN U25258 ( .A(n16886), .B(n16887), .Z(n16884) );
  NANDN U25259 ( .A(n16887), .B(n16886), .Z(n16882) );
  AND U25260 ( .A(n16888), .B(n16889), .Z(n16843) );
  NAND U25261 ( .A(n16890), .B(n16891), .Z(n16889) );
  OR U25262 ( .A(n16892), .B(n16893), .Z(n16890) );
  NANDN U25263 ( .A(n16894), .B(n16892), .Z(n16888) );
  XNOR U25264 ( .A(n16869), .B(n16895), .Z(N63895) );
  XOR U25265 ( .A(n16871), .B(n16872), .Z(n16895) );
  XNOR U25266 ( .A(n16885), .B(n16896), .Z(n16872) );
  XOR U25267 ( .A(n16886), .B(n16887), .Z(n16896) );
  XOR U25268 ( .A(n16892), .B(n16897), .Z(n16887) );
  XOR U25269 ( .A(n16891), .B(n16894), .Z(n16897) );
  IV U25270 ( .A(n16893), .Z(n16894) );
  NAND U25271 ( .A(n16898), .B(n16899), .Z(n16893) );
  OR U25272 ( .A(n16900), .B(n16901), .Z(n16899) );
  OR U25273 ( .A(n16902), .B(n16903), .Z(n16898) );
  NAND U25274 ( .A(n16904), .B(n16905), .Z(n16891) );
  OR U25275 ( .A(n16906), .B(n16907), .Z(n16905) );
  OR U25276 ( .A(n16908), .B(n16909), .Z(n16904) );
  NOR U25277 ( .A(n16910), .B(n16911), .Z(n16892) );
  ANDN U25278 ( .B(n16912), .A(n16913), .Z(n16886) );
  XNOR U25279 ( .A(n16879), .B(n16914), .Z(n16885) );
  XNOR U25280 ( .A(n16878), .B(n16880), .Z(n16914) );
  NAND U25281 ( .A(n16915), .B(n16916), .Z(n16880) );
  OR U25282 ( .A(n16917), .B(n16918), .Z(n16916) );
  OR U25283 ( .A(n16919), .B(n16920), .Z(n16915) );
  NAND U25284 ( .A(n16921), .B(n16922), .Z(n16878) );
  OR U25285 ( .A(n16923), .B(n16924), .Z(n16922) );
  OR U25286 ( .A(n16925), .B(n16926), .Z(n16921) );
  ANDN U25287 ( .B(n16927), .A(n16928), .Z(n16879) );
  IV U25288 ( .A(n16929), .Z(n16927) );
  ANDN U25289 ( .B(n16930), .A(n16931), .Z(n16871) );
  XOR U25290 ( .A(n16857), .B(n16932), .Z(n16869) );
  XOR U25291 ( .A(n16858), .B(n16859), .Z(n16932) );
  XOR U25292 ( .A(n16864), .B(n16933), .Z(n16859) );
  XOR U25293 ( .A(n16863), .B(n16866), .Z(n16933) );
  IV U25294 ( .A(n16865), .Z(n16866) );
  NAND U25295 ( .A(n16934), .B(n16935), .Z(n16865) );
  OR U25296 ( .A(n16936), .B(n16937), .Z(n16935) );
  OR U25297 ( .A(n16938), .B(n16939), .Z(n16934) );
  NAND U25298 ( .A(n16940), .B(n16941), .Z(n16863) );
  OR U25299 ( .A(n16942), .B(n16943), .Z(n16941) );
  OR U25300 ( .A(n16944), .B(n16945), .Z(n16940) );
  NOR U25301 ( .A(n16946), .B(n16947), .Z(n16864) );
  ANDN U25302 ( .B(n16948), .A(n16949), .Z(n16858) );
  IV U25303 ( .A(n16950), .Z(n16948) );
  XNOR U25304 ( .A(n16851), .B(n16951), .Z(n16857) );
  XNOR U25305 ( .A(n16850), .B(n16852), .Z(n16951) );
  NAND U25306 ( .A(n16952), .B(n16953), .Z(n16852) );
  OR U25307 ( .A(n16954), .B(n16955), .Z(n16953) );
  OR U25308 ( .A(n16956), .B(n16957), .Z(n16952) );
  NAND U25309 ( .A(n16958), .B(n16959), .Z(n16850) );
  OR U25310 ( .A(n16960), .B(n16961), .Z(n16959) );
  OR U25311 ( .A(n16962), .B(n16963), .Z(n16958) );
  ANDN U25312 ( .B(n16964), .A(n16965), .Z(n16851) );
  IV U25313 ( .A(n16966), .Z(n16964) );
  XNOR U25314 ( .A(n16931), .B(n16930), .Z(N63894) );
  XOR U25315 ( .A(n16950), .B(n16949), .Z(n16930) );
  XNOR U25316 ( .A(n16965), .B(n16966), .Z(n16949) );
  XNOR U25317 ( .A(n16960), .B(n16961), .Z(n16966) );
  XNOR U25318 ( .A(n16962), .B(n16963), .Z(n16961) );
  XNOR U25319 ( .A(y[6109]), .B(x[6109]), .Z(n16963) );
  XNOR U25320 ( .A(y[6110]), .B(x[6110]), .Z(n16962) );
  XNOR U25321 ( .A(y[6108]), .B(x[6108]), .Z(n16960) );
  XNOR U25322 ( .A(n16954), .B(n16955), .Z(n16965) );
  XNOR U25323 ( .A(y[6105]), .B(x[6105]), .Z(n16955) );
  XNOR U25324 ( .A(n16956), .B(n16957), .Z(n16954) );
  XNOR U25325 ( .A(y[6106]), .B(x[6106]), .Z(n16957) );
  XNOR U25326 ( .A(y[6107]), .B(x[6107]), .Z(n16956) );
  XNOR U25327 ( .A(n16947), .B(n16946), .Z(n16950) );
  XNOR U25328 ( .A(n16942), .B(n16943), .Z(n16946) );
  XNOR U25329 ( .A(y[6102]), .B(x[6102]), .Z(n16943) );
  XNOR U25330 ( .A(n16944), .B(n16945), .Z(n16942) );
  XNOR U25331 ( .A(y[6103]), .B(x[6103]), .Z(n16945) );
  XNOR U25332 ( .A(y[6104]), .B(x[6104]), .Z(n16944) );
  XNOR U25333 ( .A(n16936), .B(n16937), .Z(n16947) );
  XNOR U25334 ( .A(y[6099]), .B(x[6099]), .Z(n16937) );
  XNOR U25335 ( .A(n16938), .B(n16939), .Z(n16936) );
  XNOR U25336 ( .A(y[6100]), .B(x[6100]), .Z(n16939) );
  XNOR U25337 ( .A(y[6101]), .B(x[6101]), .Z(n16938) );
  XOR U25338 ( .A(n16912), .B(n16913), .Z(n16931) );
  XNOR U25339 ( .A(n16928), .B(n16929), .Z(n16913) );
  XNOR U25340 ( .A(n16923), .B(n16924), .Z(n16929) );
  XNOR U25341 ( .A(n16925), .B(n16926), .Z(n16924) );
  XNOR U25342 ( .A(y[6097]), .B(x[6097]), .Z(n16926) );
  XNOR U25343 ( .A(y[6098]), .B(x[6098]), .Z(n16925) );
  XNOR U25344 ( .A(y[6096]), .B(x[6096]), .Z(n16923) );
  XNOR U25345 ( .A(n16917), .B(n16918), .Z(n16928) );
  XNOR U25346 ( .A(y[6093]), .B(x[6093]), .Z(n16918) );
  XNOR U25347 ( .A(n16919), .B(n16920), .Z(n16917) );
  XNOR U25348 ( .A(y[6094]), .B(x[6094]), .Z(n16920) );
  XNOR U25349 ( .A(y[6095]), .B(x[6095]), .Z(n16919) );
  XOR U25350 ( .A(n16911), .B(n16910), .Z(n16912) );
  XNOR U25351 ( .A(n16906), .B(n16907), .Z(n16910) );
  XNOR U25352 ( .A(y[6090]), .B(x[6090]), .Z(n16907) );
  XNOR U25353 ( .A(n16908), .B(n16909), .Z(n16906) );
  XNOR U25354 ( .A(y[6091]), .B(x[6091]), .Z(n16909) );
  XNOR U25355 ( .A(y[6092]), .B(x[6092]), .Z(n16908) );
  XNOR U25356 ( .A(n16900), .B(n16901), .Z(n16911) );
  XNOR U25357 ( .A(y[6087]), .B(x[6087]), .Z(n16901) );
  XNOR U25358 ( .A(n16902), .B(n16903), .Z(n16900) );
  XNOR U25359 ( .A(y[6088]), .B(x[6088]), .Z(n16903) );
  XNOR U25360 ( .A(y[6089]), .B(x[6089]), .Z(n16902) );
  NAND U25361 ( .A(n16967), .B(n16968), .Z(N63885) );
  NANDN U25362 ( .A(n16969), .B(n16970), .Z(n16968) );
  OR U25363 ( .A(n16971), .B(n16972), .Z(n16970) );
  NAND U25364 ( .A(n16971), .B(n16972), .Z(n16967) );
  XOR U25365 ( .A(n16971), .B(n16973), .Z(N63884) );
  XNOR U25366 ( .A(n16969), .B(n16972), .Z(n16973) );
  AND U25367 ( .A(n16974), .B(n16975), .Z(n16972) );
  NANDN U25368 ( .A(n16976), .B(n16977), .Z(n16975) );
  NANDN U25369 ( .A(n16978), .B(n16979), .Z(n16977) );
  NANDN U25370 ( .A(n16979), .B(n16978), .Z(n16974) );
  NAND U25371 ( .A(n16980), .B(n16981), .Z(n16969) );
  NANDN U25372 ( .A(n16982), .B(n16983), .Z(n16981) );
  OR U25373 ( .A(n16984), .B(n16985), .Z(n16983) );
  NAND U25374 ( .A(n16985), .B(n16984), .Z(n16980) );
  AND U25375 ( .A(n16986), .B(n16987), .Z(n16971) );
  NANDN U25376 ( .A(n16988), .B(n16989), .Z(n16987) );
  NANDN U25377 ( .A(n16990), .B(n16991), .Z(n16989) );
  NANDN U25378 ( .A(n16991), .B(n16990), .Z(n16986) );
  XOR U25379 ( .A(n16985), .B(n16992), .Z(N63883) );
  XOR U25380 ( .A(n16982), .B(n16984), .Z(n16992) );
  XNOR U25381 ( .A(n16978), .B(n16993), .Z(n16984) );
  XNOR U25382 ( .A(n16976), .B(n16979), .Z(n16993) );
  NAND U25383 ( .A(n16994), .B(n16995), .Z(n16979) );
  NAND U25384 ( .A(n16996), .B(n16997), .Z(n16995) );
  OR U25385 ( .A(n16998), .B(n16999), .Z(n16996) );
  NANDN U25386 ( .A(n17000), .B(n16998), .Z(n16994) );
  IV U25387 ( .A(n16999), .Z(n17000) );
  NAND U25388 ( .A(n17001), .B(n17002), .Z(n16976) );
  NAND U25389 ( .A(n17003), .B(n17004), .Z(n17002) );
  NANDN U25390 ( .A(n17005), .B(n17006), .Z(n17003) );
  NANDN U25391 ( .A(n17006), .B(n17005), .Z(n17001) );
  AND U25392 ( .A(n17007), .B(n17008), .Z(n16978) );
  NAND U25393 ( .A(n17009), .B(n17010), .Z(n17008) );
  OR U25394 ( .A(n17011), .B(n17012), .Z(n17009) );
  NANDN U25395 ( .A(n17013), .B(n17011), .Z(n17007) );
  NAND U25396 ( .A(n17014), .B(n17015), .Z(n16982) );
  NANDN U25397 ( .A(n17016), .B(n17017), .Z(n17015) );
  OR U25398 ( .A(n17018), .B(n17019), .Z(n17017) );
  NANDN U25399 ( .A(n17020), .B(n17018), .Z(n17014) );
  IV U25400 ( .A(n17019), .Z(n17020) );
  XNOR U25401 ( .A(n16990), .B(n17021), .Z(n16985) );
  XNOR U25402 ( .A(n16988), .B(n16991), .Z(n17021) );
  NAND U25403 ( .A(n17022), .B(n17023), .Z(n16991) );
  NAND U25404 ( .A(n17024), .B(n17025), .Z(n17023) );
  OR U25405 ( .A(n17026), .B(n17027), .Z(n17024) );
  NANDN U25406 ( .A(n17028), .B(n17026), .Z(n17022) );
  IV U25407 ( .A(n17027), .Z(n17028) );
  NAND U25408 ( .A(n17029), .B(n17030), .Z(n16988) );
  NAND U25409 ( .A(n17031), .B(n17032), .Z(n17030) );
  NANDN U25410 ( .A(n17033), .B(n17034), .Z(n17031) );
  NANDN U25411 ( .A(n17034), .B(n17033), .Z(n17029) );
  AND U25412 ( .A(n17035), .B(n17036), .Z(n16990) );
  NAND U25413 ( .A(n17037), .B(n17038), .Z(n17036) );
  OR U25414 ( .A(n17039), .B(n17040), .Z(n17037) );
  NANDN U25415 ( .A(n17041), .B(n17039), .Z(n17035) );
  XNOR U25416 ( .A(n17016), .B(n17042), .Z(N63882) );
  XOR U25417 ( .A(n17018), .B(n17019), .Z(n17042) );
  XNOR U25418 ( .A(n17032), .B(n17043), .Z(n17019) );
  XOR U25419 ( .A(n17033), .B(n17034), .Z(n17043) );
  XOR U25420 ( .A(n17039), .B(n17044), .Z(n17034) );
  XOR U25421 ( .A(n17038), .B(n17041), .Z(n17044) );
  IV U25422 ( .A(n17040), .Z(n17041) );
  NAND U25423 ( .A(n17045), .B(n17046), .Z(n17040) );
  OR U25424 ( .A(n17047), .B(n17048), .Z(n17046) );
  OR U25425 ( .A(n17049), .B(n17050), .Z(n17045) );
  NAND U25426 ( .A(n17051), .B(n17052), .Z(n17038) );
  OR U25427 ( .A(n17053), .B(n17054), .Z(n17052) );
  OR U25428 ( .A(n17055), .B(n17056), .Z(n17051) );
  NOR U25429 ( .A(n17057), .B(n17058), .Z(n17039) );
  ANDN U25430 ( .B(n17059), .A(n17060), .Z(n17033) );
  XNOR U25431 ( .A(n17026), .B(n17061), .Z(n17032) );
  XNOR U25432 ( .A(n17025), .B(n17027), .Z(n17061) );
  NAND U25433 ( .A(n17062), .B(n17063), .Z(n17027) );
  OR U25434 ( .A(n17064), .B(n17065), .Z(n17063) );
  OR U25435 ( .A(n17066), .B(n17067), .Z(n17062) );
  NAND U25436 ( .A(n17068), .B(n17069), .Z(n17025) );
  OR U25437 ( .A(n17070), .B(n17071), .Z(n17069) );
  OR U25438 ( .A(n17072), .B(n17073), .Z(n17068) );
  ANDN U25439 ( .B(n17074), .A(n17075), .Z(n17026) );
  IV U25440 ( .A(n17076), .Z(n17074) );
  ANDN U25441 ( .B(n17077), .A(n17078), .Z(n17018) );
  XOR U25442 ( .A(n17004), .B(n17079), .Z(n17016) );
  XOR U25443 ( .A(n17005), .B(n17006), .Z(n17079) );
  XOR U25444 ( .A(n17011), .B(n17080), .Z(n17006) );
  XOR U25445 ( .A(n17010), .B(n17013), .Z(n17080) );
  IV U25446 ( .A(n17012), .Z(n17013) );
  NAND U25447 ( .A(n17081), .B(n17082), .Z(n17012) );
  OR U25448 ( .A(n17083), .B(n17084), .Z(n17082) );
  OR U25449 ( .A(n17085), .B(n17086), .Z(n17081) );
  NAND U25450 ( .A(n17087), .B(n17088), .Z(n17010) );
  OR U25451 ( .A(n17089), .B(n17090), .Z(n17088) );
  OR U25452 ( .A(n17091), .B(n17092), .Z(n17087) );
  NOR U25453 ( .A(n17093), .B(n17094), .Z(n17011) );
  ANDN U25454 ( .B(n17095), .A(n17096), .Z(n17005) );
  IV U25455 ( .A(n17097), .Z(n17095) );
  XNOR U25456 ( .A(n16998), .B(n17098), .Z(n17004) );
  XNOR U25457 ( .A(n16997), .B(n16999), .Z(n17098) );
  NAND U25458 ( .A(n17099), .B(n17100), .Z(n16999) );
  OR U25459 ( .A(n17101), .B(n17102), .Z(n17100) );
  OR U25460 ( .A(n17103), .B(n17104), .Z(n17099) );
  NAND U25461 ( .A(n17105), .B(n17106), .Z(n16997) );
  OR U25462 ( .A(n17107), .B(n17108), .Z(n17106) );
  OR U25463 ( .A(n17109), .B(n17110), .Z(n17105) );
  ANDN U25464 ( .B(n17111), .A(n17112), .Z(n16998) );
  IV U25465 ( .A(n17113), .Z(n17111) );
  XNOR U25466 ( .A(n17078), .B(n17077), .Z(N63881) );
  XOR U25467 ( .A(n17097), .B(n17096), .Z(n17077) );
  XNOR U25468 ( .A(n17112), .B(n17113), .Z(n17096) );
  XNOR U25469 ( .A(n17107), .B(n17108), .Z(n17113) );
  XNOR U25470 ( .A(n17109), .B(n17110), .Z(n17108) );
  XNOR U25471 ( .A(y[6085]), .B(x[6085]), .Z(n17110) );
  XNOR U25472 ( .A(y[6086]), .B(x[6086]), .Z(n17109) );
  XNOR U25473 ( .A(y[6084]), .B(x[6084]), .Z(n17107) );
  XNOR U25474 ( .A(n17101), .B(n17102), .Z(n17112) );
  XNOR U25475 ( .A(y[6081]), .B(x[6081]), .Z(n17102) );
  XNOR U25476 ( .A(n17103), .B(n17104), .Z(n17101) );
  XNOR U25477 ( .A(y[6082]), .B(x[6082]), .Z(n17104) );
  XNOR U25478 ( .A(y[6083]), .B(x[6083]), .Z(n17103) );
  XNOR U25479 ( .A(n17094), .B(n17093), .Z(n17097) );
  XNOR U25480 ( .A(n17089), .B(n17090), .Z(n17093) );
  XNOR U25481 ( .A(y[6078]), .B(x[6078]), .Z(n17090) );
  XNOR U25482 ( .A(n17091), .B(n17092), .Z(n17089) );
  XNOR U25483 ( .A(y[6079]), .B(x[6079]), .Z(n17092) );
  XNOR U25484 ( .A(y[6080]), .B(x[6080]), .Z(n17091) );
  XNOR U25485 ( .A(n17083), .B(n17084), .Z(n17094) );
  XNOR U25486 ( .A(y[6075]), .B(x[6075]), .Z(n17084) );
  XNOR U25487 ( .A(n17085), .B(n17086), .Z(n17083) );
  XNOR U25488 ( .A(y[6076]), .B(x[6076]), .Z(n17086) );
  XNOR U25489 ( .A(y[6077]), .B(x[6077]), .Z(n17085) );
  XOR U25490 ( .A(n17059), .B(n17060), .Z(n17078) );
  XNOR U25491 ( .A(n17075), .B(n17076), .Z(n17060) );
  XNOR U25492 ( .A(n17070), .B(n17071), .Z(n17076) );
  XNOR U25493 ( .A(n17072), .B(n17073), .Z(n17071) );
  XNOR U25494 ( .A(y[6073]), .B(x[6073]), .Z(n17073) );
  XNOR U25495 ( .A(y[6074]), .B(x[6074]), .Z(n17072) );
  XNOR U25496 ( .A(y[6072]), .B(x[6072]), .Z(n17070) );
  XNOR U25497 ( .A(n17064), .B(n17065), .Z(n17075) );
  XNOR U25498 ( .A(y[6069]), .B(x[6069]), .Z(n17065) );
  XNOR U25499 ( .A(n17066), .B(n17067), .Z(n17064) );
  XNOR U25500 ( .A(y[6070]), .B(x[6070]), .Z(n17067) );
  XNOR U25501 ( .A(y[6071]), .B(x[6071]), .Z(n17066) );
  XOR U25502 ( .A(n17058), .B(n17057), .Z(n17059) );
  XNOR U25503 ( .A(n17053), .B(n17054), .Z(n17057) );
  XNOR U25504 ( .A(y[6066]), .B(x[6066]), .Z(n17054) );
  XNOR U25505 ( .A(n17055), .B(n17056), .Z(n17053) );
  XNOR U25506 ( .A(y[6067]), .B(x[6067]), .Z(n17056) );
  XNOR U25507 ( .A(y[6068]), .B(x[6068]), .Z(n17055) );
  XNOR U25508 ( .A(n17047), .B(n17048), .Z(n17058) );
  XNOR U25509 ( .A(y[6063]), .B(x[6063]), .Z(n17048) );
  XNOR U25510 ( .A(n17049), .B(n17050), .Z(n17047) );
  XNOR U25511 ( .A(y[6064]), .B(x[6064]), .Z(n17050) );
  XNOR U25512 ( .A(y[6065]), .B(x[6065]), .Z(n17049) );
  NAND U25513 ( .A(n17114), .B(n17115), .Z(N63872) );
  NANDN U25514 ( .A(n17116), .B(n17117), .Z(n17115) );
  OR U25515 ( .A(n17118), .B(n17119), .Z(n17117) );
  NAND U25516 ( .A(n17118), .B(n17119), .Z(n17114) );
  XOR U25517 ( .A(n17118), .B(n17120), .Z(N63871) );
  XNOR U25518 ( .A(n17116), .B(n17119), .Z(n17120) );
  AND U25519 ( .A(n17121), .B(n17122), .Z(n17119) );
  NANDN U25520 ( .A(n17123), .B(n17124), .Z(n17122) );
  NANDN U25521 ( .A(n17125), .B(n17126), .Z(n17124) );
  NANDN U25522 ( .A(n17126), .B(n17125), .Z(n17121) );
  NAND U25523 ( .A(n17127), .B(n17128), .Z(n17116) );
  NANDN U25524 ( .A(n17129), .B(n17130), .Z(n17128) );
  OR U25525 ( .A(n17131), .B(n17132), .Z(n17130) );
  NAND U25526 ( .A(n17132), .B(n17131), .Z(n17127) );
  AND U25527 ( .A(n17133), .B(n17134), .Z(n17118) );
  NANDN U25528 ( .A(n17135), .B(n17136), .Z(n17134) );
  NANDN U25529 ( .A(n17137), .B(n17138), .Z(n17136) );
  NANDN U25530 ( .A(n17138), .B(n17137), .Z(n17133) );
  XOR U25531 ( .A(n17132), .B(n17139), .Z(N63870) );
  XOR U25532 ( .A(n17129), .B(n17131), .Z(n17139) );
  XNOR U25533 ( .A(n17125), .B(n17140), .Z(n17131) );
  XNOR U25534 ( .A(n17123), .B(n17126), .Z(n17140) );
  NAND U25535 ( .A(n17141), .B(n17142), .Z(n17126) );
  NAND U25536 ( .A(n17143), .B(n17144), .Z(n17142) );
  OR U25537 ( .A(n17145), .B(n17146), .Z(n17143) );
  NANDN U25538 ( .A(n17147), .B(n17145), .Z(n17141) );
  IV U25539 ( .A(n17146), .Z(n17147) );
  NAND U25540 ( .A(n17148), .B(n17149), .Z(n17123) );
  NAND U25541 ( .A(n17150), .B(n17151), .Z(n17149) );
  NANDN U25542 ( .A(n17152), .B(n17153), .Z(n17150) );
  NANDN U25543 ( .A(n17153), .B(n17152), .Z(n17148) );
  AND U25544 ( .A(n17154), .B(n17155), .Z(n17125) );
  NAND U25545 ( .A(n17156), .B(n17157), .Z(n17155) );
  OR U25546 ( .A(n17158), .B(n17159), .Z(n17156) );
  NANDN U25547 ( .A(n17160), .B(n17158), .Z(n17154) );
  NAND U25548 ( .A(n17161), .B(n17162), .Z(n17129) );
  NANDN U25549 ( .A(n17163), .B(n17164), .Z(n17162) );
  OR U25550 ( .A(n17165), .B(n17166), .Z(n17164) );
  NANDN U25551 ( .A(n17167), .B(n17165), .Z(n17161) );
  IV U25552 ( .A(n17166), .Z(n17167) );
  XNOR U25553 ( .A(n17137), .B(n17168), .Z(n17132) );
  XNOR U25554 ( .A(n17135), .B(n17138), .Z(n17168) );
  NAND U25555 ( .A(n17169), .B(n17170), .Z(n17138) );
  NAND U25556 ( .A(n17171), .B(n17172), .Z(n17170) );
  OR U25557 ( .A(n17173), .B(n17174), .Z(n17171) );
  NANDN U25558 ( .A(n17175), .B(n17173), .Z(n17169) );
  IV U25559 ( .A(n17174), .Z(n17175) );
  NAND U25560 ( .A(n17176), .B(n17177), .Z(n17135) );
  NAND U25561 ( .A(n17178), .B(n17179), .Z(n17177) );
  NANDN U25562 ( .A(n17180), .B(n17181), .Z(n17178) );
  NANDN U25563 ( .A(n17181), .B(n17180), .Z(n17176) );
  AND U25564 ( .A(n17182), .B(n17183), .Z(n17137) );
  NAND U25565 ( .A(n17184), .B(n17185), .Z(n17183) );
  OR U25566 ( .A(n17186), .B(n17187), .Z(n17184) );
  NANDN U25567 ( .A(n17188), .B(n17186), .Z(n17182) );
  XNOR U25568 ( .A(n17163), .B(n17189), .Z(N63869) );
  XOR U25569 ( .A(n17165), .B(n17166), .Z(n17189) );
  XNOR U25570 ( .A(n17179), .B(n17190), .Z(n17166) );
  XOR U25571 ( .A(n17180), .B(n17181), .Z(n17190) );
  XOR U25572 ( .A(n17186), .B(n17191), .Z(n17181) );
  XOR U25573 ( .A(n17185), .B(n17188), .Z(n17191) );
  IV U25574 ( .A(n17187), .Z(n17188) );
  NAND U25575 ( .A(n17192), .B(n17193), .Z(n17187) );
  OR U25576 ( .A(n17194), .B(n17195), .Z(n17193) );
  OR U25577 ( .A(n17196), .B(n17197), .Z(n17192) );
  NAND U25578 ( .A(n17198), .B(n17199), .Z(n17185) );
  OR U25579 ( .A(n17200), .B(n17201), .Z(n17199) );
  OR U25580 ( .A(n17202), .B(n17203), .Z(n17198) );
  NOR U25581 ( .A(n17204), .B(n17205), .Z(n17186) );
  ANDN U25582 ( .B(n17206), .A(n17207), .Z(n17180) );
  XNOR U25583 ( .A(n17173), .B(n17208), .Z(n17179) );
  XNOR U25584 ( .A(n17172), .B(n17174), .Z(n17208) );
  NAND U25585 ( .A(n17209), .B(n17210), .Z(n17174) );
  OR U25586 ( .A(n17211), .B(n17212), .Z(n17210) );
  OR U25587 ( .A(n17213), .B(n17214), .Z(n17209) );
  NAND U25588 ( .A(n17215), .B(n17216), .Z(n17172) );
  OR U25589 ( .A(n17217), .B(n17218), .Z(n17216) );
  OR U25590 ( .A(n17219), .B(n17220), .Z(n17215) );
  ANDN U25591 ( .B(n17221), .A(n17222), .Z(n17173) );
  IV U25592 ( .A(n17223), .Z(n17221) );
  ANDN U25593 ( .B(n17224), .A(n17225), .Z(n17165) );
  XOR U25594 ( .A(n17151), .B(n17226), .Z(n17163) );
  XOR U25595 ( .A(n17152), .B(n17153), .Z(n17226) );
  XOR U25596 ( .A(n17158), .B(n17227), .Z(n17153) );
  XOR U25597 ( .A(n17157), .B(n17160), .Z(n17227) );
  IV U25598 ( .A(n17159), .Z(n17160) );
  NAND U25599 ( .A(n17228), .B(n17229), .Z(n17159) );
  OR U25600 ( .A(n17230), .B(n17231), .Z(n17229) );
  OR U25601 ( .A(n17232), .B(n17233), .Z(n17228) );
  NAND U25602 ( .A(n17234), .B(n17235), .Z(n17157) );
  OR U25603 ( .A(n17236), .B(n17237), .Z(n17235) );
  OR U25604 ( .A(n17238), .B(n17239), .Z(n17234) );
  NOR U25605 ( .A(n17240), .B(n17241), .Z(n17158) );
  ANDN U25606 ( .B(n17242), .A(n17243), .Z(n17152) );
  IV U25607 ( .A(n17244), .Z(n17242) );
  XNOR U25608 ( .A(n17145), .B(n17245), .Z(n17151) );
  XNOR U25609 ( .A(n17144), .B(n17146), .Z(n17245) );
  NAND U25610 ( .A(n17246), .B(n17247), .Z(n17146) );
  OR U25611 ( .A(n17248), .B(n17249), .Z(n17247) );
  OR U25612 ( .A(n17250), .B(n17251), .Z(n17246) );
  NAND U25613 ( .A(n17252), .B(n17253), .Z(n17144) );
  OR U25614 ( .A(n17254), .B(n17255), .Z(n17253) );
  OR U25615 ( .A(n17256), .B(n17257), .Z(n17252) );
  ANDN U25616 ( .B(n17258), .A(n17259), .Z(n17145) );
  IV U25617 ( .A(n17260), .Z(n17258) );
  XNOR U25618 ( .A(n17225), .B(n17224), .Z(N63868) );
  XOR U25619 ( .A(n17244), .B(n17243), .Z(n17224) );
  XNOR U25620 ( .A(n17259), .B(n17260), .Z(n17243) );
  XNOR U25621 ( .A(n17254), .B(n17255), .Z(n17260) );
  XNOR U25622 ( .A(n17256), .B(n17257), .Z(n17255) );
  XNOR U25623 ( .A(y[6061]), .B(x[6061]), .Z(n17257) );
  XNOR U25624 ( .A(y[6062]), .B(x[6062]), .Z(n17256) );
  XNOR U25625 ( .A(y[6060]), .B(x[6060]), .Z(n17254) );
  XNOR U25626 ( .A(n17248), .B(n17249), .Z(n17259) );
  XNOR U25627 ( .A(y[6057]), .B(x[6057]), .Z(n17249) );
  XNOR U25628 ( .A(n17250), .B(n17251), .Z(n17248) );
  XNOR U25629 ( .A(y[6058]), .B(x[6058]), .Z(n17251) );
  XNOR U25630 ( .A(y[6059]), .B(x[6059]), .Z(n17250) );
  XNOR U25631 ( .A(n17241), .B(n17240), .Z(n17244) );
  XNOR U25632 ( .A(n17236), .B(n17237), .Z(n17240) );
  XNOR U25633 ( .A(y[6054]), .B(x[6054]), .Z(n17237) );
  XNOR U25634 ( .A(n17238), .B(n17239), .Z(n17236) );
  XNOR U25635 ( .A(y[6055]), .B(x[6055]), .Z(n17239) );
  XNOR U25636 ( .A(y[6056]), .B(x[6056]), .Z(n17238) );
  XNOR U25637 ( .A(n17230), .B(n17231), .Z(n17241) );
  XNOR U25638 ( .A(y[6051]), .B(x[6051]), .Z(n17231) );
  XNOR U25639 ( .A(n17232), .B(n17233), .Z(n17230) );
  XNOR U25640 ( .A(y[6052]), .B(x[6052]), .Z(n17233) );
  XNOR U25641 ( .A(y[6053]), .B(x[6053]), .Z(n17232) );
  XOR U25642 ( .A(n17206), .B(n17207), .Z(n17225) );
  XNOR U25643 ( .A(n17222), .B(n17223), .Z(n17207) );
  XNOR U25644 ( .A(n17217), .B(n17218), .Z(n17223) );
  XNOR U25645 ( .A(n17219), .B(n17220), .Z(n17218) );
  XNOR U25646 ( .A(y[6049]), .B(x[6049]), .Z(n17220) );
  XNOR U25647 ( .A(y[6050]), .B(x[6050]), .Z(n17219) );
  XNOR U25648 ( .A(y[6048]), .B(x[6048]), .Z(n17217) );
  XNOR U25649 ( .A(n17211), .B(n17212), .Z(n17222) );
  XNOR U25650 ( .A(y[6045]), .B(x[6045]), .Z(n17212) );
  XNOR U25651 ( .A(n17213), .B(n17214), .Z(n17211) );
  XNOR U25652 ( .A(y[6046]), .B(x[6046]), .Z(n17214) );
  XNOR U25653 ( .A(y[6047]), .B(x[6047]), .Z(n17213) );
  XOR U25654 ( .A(n17205), .B(n17204), .Z(n17206) );
  XNOR U25655 ( .A(n17200), .B(n17201), .Z(n17204) );
  XNOR U25656 ( .A(y[6042]), .B(x[6042]), .Z(n17201) );
  XNOR U25657 ( .A(n17202), .B(n17203), .Z(n17200) );
  XNOR U25658 ( .A(y[6043]), .B(x[6043]), .Z(n17203) );
  XNOR U25659 ( .A(y[6044]), .B(x[6044]), .Z(n17202) );
  XNOR U25660 ( .A(n17194), .B(n17195), .Z(n17205) );
  XNOR U25661 ( .A(y[6039]), .B(x[6039]), .Z(n17195) );
  XNOR U25662 ( .A(n17196), .B(n17197), .Z(n17194) );
  XNOR U25663 ( .A(y[6040]), .B(x[6040]), .Z(n17197) );
  XNOR U25664 ( .A(y[6041]), .B(x[6041]), .Z(n17196) );
  NAND U25665 ( .A(n17261), .B(n17262), .Z(N63859) );
  NANDN U25666 ( .A(n17263), .B(n17264), .Z(n17262) );
  OR U25667 ( .A(n17265), .B(n17266), .Z(n17264) );
  NAND U25668 ( .A(n17265), .B(n17266), .Z(n17261) );
  XOR U25669 ( .A(n17265), .B(n17267), .Z(N63858) );
  XNOR U25670 ( .A(n17263), .B(n17266), .Z(n17267) );
  AND U25671 ( .A(n17268), .B(n17269), .Z(n17266) );
  NANDN U25672 ( .A(n17270), .B(n17271), .Z(n17269) );
  NANDN U25673 ( .A(n17272), .B(n17273), .Z(n17271) );
  NANDN U25674 ( .A(n17273), .B(n17272), .Z(n17268) );
  NAND U25675 ( .A(n17274), .B(n17275), .Z(n17263) );
  NANDN U25676 ( .A(n17276), .B(n17277), .Z(n17275) );
  OR U25677 ( .A(n17278), .B(n17279), .Z(n17277) );
  NAND U25678 ( .A(n17279), .B(n17278), .Z(n17274) );
  AND U25679 ( .A(n17280), .B(n17281), .Z(n17265) );
  NANDN U25680 ( .A(n17282), .B(n17283), .Z(n17281) );
  NANDN U25681 ( .A(n17284), .B(n17285), .Z(n17283) );
  NANDN U25682 ( .A(n17285), .B(n17284), .Z(n17280) );
  XOR U25683 ( .A(n17279), .B(n17286), .Z(N63857) );
  XOR U25684 ( .A(n17276), .B(n17278), .Z(n17286) );
  XNOR U25685 ( .A(n17272), .B(n17287), .Z(n17278) );
  XNOR U25686 ( .A(n17270), .B(n17273), .Z(n17287) );
  NAND U25687 ( .A(n17288), .B(n17289), .Z(n17273) );
  NAND U25688 ( .A(n17290), .B(n17291), .Z(n17289) );
  OR U25689 ( .A(n17292), .B(n17293), .Z(n17290) );
  NANDN U25690 ( .A(n17294), .B(n17292), .Z(n17288) );
  IV U25691 ( .A(n17293), .Z(n17294) );
  NAND U25692 ( .A(n17295), .B(n17296), .Z(n17270) );
  NAND U25693 ( .A(n17297), .B(n17298), .Z(n17296) );
  NANDN U25694 ( .A(n17299), .B(n17300), .Z(n17297) );
  NANDN U25695 ( .A(n17300), .B(n17299), .Z(n17295) );
  AND U25696 ( .A(n17301), .B(n17302), .Z(n17272) );
  NAND U25697 ( .A(n17303), .B(n17304), .Z(n17302) );
  OR U25698 ( .A(n17305), .B(n17306), .Z(n17303) );
  NANDN U25699 ( .A(n17307), .B(n17305), .Z(n17301) );
  NAND U25700 ( .A(n17308), .B(n17309), .Z(n17276) );
  NANDN U25701 ( .A(n17310), .B(n17311), .Z(n17309) );
  OR U25702 ( .A(n17312), .B(n17313), .Z(n17311) );
  NANDN U25703 ( .A(n17314), .B(n17312), .Z(n17308) );
  IV U25704 ( .A(n17313), .Z(n17314) );
  XNOR U25705 ( .A(n17284), .B(n17315), .Z(n17279) );
  XNOR U25706 ( .A(n17282), .B(n17285), .Z(n17315) );
  NAND U25707 ( .A(n17316), .B(n17317), .Z(n17285) );
  NAND U25708 ( .A(n17318), .B(n17319), .Z(n17317) );
  OR U25709 ( .A(n17320), .B(n17321), .Z(n17318) );
  NANDN U25710 ( .A(n17322), .B(n17320), .Z(n17316) );
  IV U25711 ( .A(n17321), .Z(n17322) );
  NAND U25712 ( .A(n17323), .B(n17324), .Z(n17282) );
  NAND U25713 ( .A(n17325), .B(n17326), .Z(n17324) );
  NANDN U25714 ( .A(n17327), .B(n17328), .Z(n17325) );
  NANDN U25715 ( .A(n17328), .B(n17327), .Z(n17323) );
  AND U25716 ( .A(n17329), .B(n17330), .Z(n17284) );
  NAND U25717 ( .A(n17331), .B(n17332), .Z(n17330) );
  OR U25718 ( .A(n17333), .B(n17334), .Z(n17331) );
  NANDN U25719 ( .A(n17335), .B(n17333), .Z(n17329) );
  XNOR U25720 ( .A(n17310), .B(n17336), .Z(N63856) );
  XOR U25721 ( .A(n17312), .B(n17313), .Z(n17336) );
  XNOR U25722 ( .A(n17326), .B(n17337), .Z(n17313) );
  XOR U25723 ( .A(n17327), .B(n17328), .Z(n17337) );
  XOR U25724 ( .A(n17333), .B(n17338), .Z(n17328) );
  XOR U25725 ( .A(n17332), .B(n17335), .Z(n17338) );
  IV U25726 ( .A(n17334), .Z(n17335) );
  NAND U25727 ( .A(n17339), .B(n17340), .Z(n17334) );
  OR U25728 ( .A(n17341), .B(n17342), .Z(n17340) );
  OR U25729 ( .A(n17343), .B(n17344), .Z(n17339) );
  NAND U25730 ( .A(n17345), .B(n17346), .Z(n17332) );
  OR U25731 ( .A(n17347), .B(n17348), .Z(n17346) );
  OR U25732 ( .A(n17349), .B(n17350), .Z(n17345) );
  NOR U25733 ( .A(n17351), .B(n17352), .Z(n17333) );
  ANDN U25734 ( .B(n17353), .A(n17354), .Z(n17327) );
  XNOR U25735 ( .A(n17320), .B(n17355), .Z(n17326) );
  XNOR U25736 ( .A(n17319), .B(n17321), .Z(n17355) );
  NAND U25737 ( .A(n17356), .B(n17357), .Z(n17321) );
  OR U25738 ( .A(n17358), .B(n17359), .Z(n17357) );
  OR U25739 ( .A(n17360), .B(n17361), .Z(n17356) );
  NAND U25740 ( .A(n17362), .B(n17363), .Z(n17319) );
  OR U25741 ( .A(n17364), .B(n17365), .Z(n17363) );
  OR U25742 ( .A(n17366), .B(n17367), .Z(n17362) );
  ANDN U25743 ( .B(n17368), .A(n17369), .Z(n17320) );
  IV U25744 ( .A(n17370), .Z(n17368) );
  ANDN U25745 ( .B(n17371), .A(n17372), .Z(n17312) );
  XOR U25746 ( .A(n17298), .B(n17373), .Z(n17310) );
  XOR U25747 ( .A(n17299), .B(n17300), .Z(n17373) );
  XOR U25748 ( .A(n17305), .B(n17374), .Z(n17300) );
  XOR U25749 ( .A(n17304), .B(n17307), .Z(n17374) );
  IV U25750 ( .A(n17306), .Z(n17307) );
  NAND U25751 ( .A(n17375), .B(n17376), .Z(n17306) );
  OR U25752 ( .A(n17377), .B(n17378), .Z(n17376) );
  OR U25753 ( .A(n17379), .B(n17380), .Z(n17375) );
  NAND U25754 ( .A(n17381), .B(n17382), .Z(n17304) );
  OR U25755 ( .A(n17383), .B(n17384), .Z(n17382) );
  OR U25756 ( .A(n17385), .B(n17386), .Z(n17381) );
  NOR U25757 ( .A(n17387), .B(n17388), .Z(n17305) );
  ANDN U25758 ( .B(n17389), .A(n17390), .Z(n17299) );
  IV U25759 ( .A(n17391), .Z(n17389) );
  XNOR U25760 ( .A(n17292), .B(n17392), .Z(n17298) );
  XNOR U25761 ( .A(n17291), .B(n17293), .Z(n17392) );
  NAND U25762 ( .A(n17393), .B(n17394), .Z(n17293) );
  OR U25763 ( .A(n17395), .B(n17396), .Z(n17394) );
  OR U25764 ( .A(n17397), .B(n17398), .Z(n17393) );
  NAND U25765 ( .A(n17399), .B(n17400), .Z(n17291) );
  OR U25766 ( .A(n17401), .B(n17402), .Z(n17400) );
  OR U25767 ( .A(n17403), .B(n17404), .Z(n17399) );
  ANDN U25768 ( .B(n17405), .A(n17406), .Z(n17292) );
  IV U25769 ( .A(n17407), .Z(n17405) );
  XNOR U25770 ( .A(n17372), .B(n17371), .Z(N63855) );
  XOR U25771 ( .A(n17391), .B(n17390), .Z(n17371) );
  XNOR U25772 ( .A(n17406), .B(n17407), .Z(n17390) );
  XNOR U25773 ( .A(n17401), .B(n17402), .Z(n17407) );
  XNOR U25774 ( .A(n17403), .B(n17404), .Z(n17402) );
  XNOR U25775 ( .A(y[6037]), .B(x[6037]), .Z(n17404) );
  XNOR U25776 ( .A(y[6038]), .B(x[6038]), .Z(n17403) );
  XNOR U25777 ( .A(y[6036]), .B(x[6036]), .Z(n17401) );
  XNOR U25778 ( .A(n17395), .B(n17396), .Z(n17406) );
  XNOR U25779 ( .A(y[6033]), .B(x[6033]), .Z(n17396) );
  XNOR U25780 ( .A(n17397), .B(n17398), .Z(n17395) );
  XNOR U25781 ( .A(y[6034]), .B(x[6034]), .Z(n17398) );
  XNOR U25782 ( .A(y[6035]), .B(x[6035]), .Z(n17397) );
  XNOR U25783 ( .A(n17388), .B(n17387), .Z(n17391) );
  XNOR U25784 ( .A(n17383), .B(n17384), .Z(n17387) );
  XNOR U25785 ( .A(y[6030]), .B(x[6030]), .Z(n17384) );
  XNOR U25786 ( .A(n17385), .B(n17386), .Z(n17383) );
  XNOR U25787 ( .A(y[6031]), .B(x[6031]), .Z(n17386) );
  XNOR U25788 ( .A(y[6032]), .B(x[6032]), .Z(n17385) );
  XNOR U25789 ( .A(n17377), .B(n17378), .Z(n17388) );
  XNOR U25790 ( .A(y[6027]), .B(x[6027]), .Z(n17378) );
  XNOR U25791 ( .A(n17379), .B(n17380), .Z(n17377) );
  XNOR U25792 ( .A(y[6028]), .B(x[6028]), .Z(n17380) );
  XNOR U25793 ( .A(y[6029]), .B(x[6029]), .Z(n17379) );
  XOR U25794 ( .A(n17353), .B(n17354), .Z(n17372) );
  XNOR U25795 ( .A(n17369), .B(n17370), .Z(n17354) );
  XNOR U25796 ( .A(n17364), .B(n17365), .Z(n17370) );
  XNOR U25797 ( .A(n17366), .B(n17367), .Z(n17365) );
  XNOR U25798 ( .A(y[6025]), .B(x[6025]), .Z(n17367) );
  XNOR U25799 ( .A(y[6026]), .B(x[6026]), .Z(n17366) );
  XNOR U25800 ( .A(y[6024]), .B(x[6024]), .Z(n17364) );
  XNOR U25801 ( .A(n17358), .B(n17359), .Z(n17369) );
  XNOR U25802 ( .A(y[6021]), .B(x[6021]), .Z(n17359) );
  XNOR U25803 ( .A(n17360), .B(n17361), .Z(n17358) );
  XNOR U25804 ( .A(y[6022]), .B(x[6022]), .Z(n17361) );
  XNOR U25805 ( .A(y[6023]), .B(x[6023]), .Z(n17360) );
  XOR U25806 ( .A(n17352), .B(n17351), .Z(n17353) );
  XNOR U25807 ( .A(n17347), .B(n17348), .Z(n17351) );
  XNOR U25808 ( .A(y[6018]), .B(x[6018]), .Z(n17348) );
  XNOR U25809 ( .A(n17349), .B(n17350), .Z(n17347) );
  XNOR U25810 ( .A(y[6019]), .B(x[6019]), .Z(n17350) );
  XNOR U25811 ( .A(y[6020]), .B(x[6020]), .Z(n17349) );
  XNOR U25812 ( .A(n17341), .B(n17342), .Z(n17352) );
  XNOR U25813 ( .A(y[6015]), .B(x[6015]), .Z(n17342) );
  XNOR U25814 ( .A(n17343), .B(n17344), .Z(n17341) );
  XNOR U25815 ( .A(y[6016]), .B(x[6016]), .Z(n17344) );
  XNOR U25816 ( .A(y[6017]), .B(x[6017]), .Z(n17343) );
  NAND U25817 ( .A(n17408), .B(n17409), .Z(N63846) );
  NANDN U25818 ( .A(n17410), .B(n17411), .Z(n17409) );
  OR U25819 ( .A(n17412), .B(n17413), .Z(n17411) );
  NAND U25820 ( .A(n17412), .B(n17413), .Z(n17408) );
  XOR U25821 ( .A(n17412), .B(n17414), .Z(N63845) );
  XNOR U25822 ( .A(n17410), .B(n17413), .Z(n17414) );
  AND U25823 ( .A(n17415), .B(n17416), .Z(n17413) );
  NANDN U25824 ( .A(n17417), .B(n17418), .Z(n17416) );
  NANDN U25825 ( .A(n17419), .B(n17420), .Z(n17418) );
  NANDN U25826 ( .A(n17420), .B(n17419), .Z(n17415) );
  NAND U25827 ( .A(n17421), .B(n17422), .Z(n17410) );
  NANDN U25828 ( .A(n17423), .B(n17424), .Z(n17422) );
  OR U25829 ( .A(n17425), .B(n17426), .Z(n17424) );
  NAND U25830 ( .A(n17426), .B(n17425), .Z(n17421) );
  AND U25831 ( .A(n17427), .B(n17428), .Z(n17412) );
  NANDN U25832 ( .A(n17429), .B(n17430), .Z(n17428) );
  NANDN U25833 ( .A(n17431), .B(n17432), .Z(n17430) );
  NANDN U25834 ( .A(n17432), .B(n17431), .Z(n17427) );
  XOR U25835 ( .A(n17426), .B(n17433), .Z(N63844) );
  XOR U25836 ( .A(n17423), .B(n17425), .Z(n17433) );
  XNOR U25837 ( .A(n17419), .B(n17434), .Z(n17425) );
  XNOR U25838 ( .A(n17417), .B(n17420), .Z(n17434) );
  NAND U25839 ( .A(n17435), .B(n17436), .Z(n17420) );
  NAND U25840 ( .A(n17437), .B(n17438), .Z(n17436) );
  OR U25841 ( .A(n17439), .B(n17440), .Z(n17437) );
  NANDN U25842 ( .A(n17441), .B(n17439), .Z(n17435) );
  IV U25843 ( .A(n17440), .Z(n17441) );
  NAND U25844 ( .A(n17442), .B(n17443), .Z(n17417) );
  NAND U25845 ( .A(n17444), .B(n17445), .Z(n17443) );
  NANDN U25846 ( .A(n17446), .B(n17447), .Z(n17444) );
  NANDN U25847 ( .A(n17447), .B(n17446), .Z(n17442) );
  AND U25848 ( .A(n17448), .B(n17449), .Z(n17419) );
  NAND U25849 ( .A(n17450), .B(n17451), .Z(n17449) );
  OR U25850 ( .A(n17452), .B(n17453), .Z(n17450) );
  NANDN U25851 ( .A(n17454), .B(n17452), .Z(n17448) );
  NAND U25852 ( .A(n17455), .B(n17456), .Z(n17423) );
  NANDN U25853 ( .A(n17457), .B(n17458), .Z(n17456) );
  OR U25854 ( .A(n17459), .B(n17460), .Z(n17458) );
  NANDN U25855 ( .A(n17461), .B(n17459), .Z(n17455) );
  IV U25856 ( .A(n17460), .Z(n17461) );
  XNOR U25857 ( .A(n17431), .B(n17462), .Z(n17426) );
  XNOR U25858 ( .A(n17429), .B(n17432), .Z(n17462) );
  NAND U25859 ( .A(n17463), .B(n17464), .Z(n17432) );
  NAND U25860 ( .A(n17465), .B(n17466), .Z(n17464) );
  OR U25861 ( .A(n17467), .B(n17468), .Z(n17465) );
  NANDN U25862 ( .A(n17469), .B(n17467), .Z(n17463) );
  IV U25863 ( .A(n17468), .Z(n17469) );
  NAND U25864 ( .A(n17470), .B(n17471), .Z(n17429) );
  NAND U25865 ( .A(n17472), .B(n17473), .Z(n17471) );
  NANDN U25866 ( .A(n17474), .B(n17475), .Z(n17472) );
  NANDN U25867 ( .A(n17475), .B(n17474), .Z(n17470) );
  AND U25868 ( .A(n17476), .B(n17477), .Z(n17431) );
  NAND U25869 ( .A(n17478), .B(n17479), .Z(n17477) );
  OR U25870 ( .A(n17480), .B(n17481), .Z(n17478) );
  NANDN U25871 ( .A(n17482), .B(n17480), .Z(n17476) );
  XNOR U25872 ( .A(n17457), .B(n17483), .Z(N63843) );
  XOR U25873 ( .A(n17459), .B(n17460), .Z(n17483) );
  XNOR U25874 ( .A(n17473), .B(n17484), .Z(n17460) );
  XOR U25875 ( .A(n17474), .B(n17475), .Z(n17484) );
  XOR U25876 ( .A(n17480), .B(n17485), .Z(n17475) );
  XOR U25877 ( .A(n17479), .B(n17482), .Z(n17485) );
  IV U25878 ( .A(n17481), .Z(n17482) );
  NAND U25879 ( .A(n17486), .B(n17487), .Z(n17481) );
  OR U25880 ( .A(n17488), .B(n17489), .Z(n17487) );
  OR U25881 ( .A(n17490), .B(n17491), .Z(n17486) );
  NAND U25882 ( .A(n17492), .B(n17493), .Z(n17479) );
  OR U25883 ( .A(n17494), .B(n17495), .Z(n17493) );
  OR U25884 ( .A(n17496), .B(n17497), .Z(n17492) );
  NOR U25885 ( .A(n17498), .B(n17499), .Z(n17480) );
  ANDN U25886 ( .B(n17500), .A(n17501), .Z(n17474) );
  XNOR U25887 ( .A(n17467), .B(n17502), .Z(n17473) );
  XNOR U25888 ( .A(n17466), .B(n17468), .Z(n17502) );
  NAND U25889 ( .A(n17503), .B(n17504), .Z(n17468) );
  OR U25890 ( .A(n17505), .B(n17506), .Z(n17504) );
  OR U25891 ( .A(n17507), .B(n17508), .Z(n17503) );
  NAND U25892 ( .A(n17509), .B(n17510), .Z(n17466) );
  OR U25893 ( .A(n17511), .B(n17512), .Z(n17510) );
  OR U25894 ( .A(n17513), .B(n17514), .Z(n17509) );
  ANDN U25895 ( .B(n17515), .A(n17516), .Z(n17467) );
  IV U25896 ( .A(n17517), .Z(n17515) );
  ANDN U25897 ( .B(n17518), .A(n17519), .Z(n17459) );
  XOR U25898 ( .A(n17445), .B(n17520), .Z(n17457) );
  XOR U25899 ( .A(n17446), .B(n17447), .Z(n17520) );
  XOR U25900 ( .A(n17452), .B(n17521), .Z(n17447) );
  XOR U25901 ( .A(n17451), .B(n17454), .Z(n17521) );
  IV U25902 ( .A(n17453), .Z(n17454) );
  NAND U25903 ( .A(n17522), .B(n17523), .Z(n17453) );
  OR U25904 ( .A(n17524), .B(n17525), .Z(n17523) );
  OR U25905 ( .A(n17526), .B(n17527), .Z(n17522) );
  NAND U25906 ( .A(n17528), .B(n17529), .Z(n17451) );
  OR U25907 ( .A(n17530), .B(n17531), .Z(n17529) );
  OR U25908 ( .A(n17532), .B(n17533), .Z(n17528) );
  NOR U25909 ( .A(n17534), .B(n17535), .Z(n17452) );
  ANDN U25910 ( .B(n17536), .A(n17537), .Z(n17446) );
  IV U25911 ( .A(n17538), .Z(n17536) );
  XNOR U25912 ( .A(n17439), .B(n17539), .Z(n17445) );
  XNOR U25913 ( .A(n17438), .B(n17440), .Z(n17539) );
  NAND U25914 ( .A(n17540), .B(n17541), .Z(n17440) );
  OR U25915 ( .A(n17542), .B(n17543), .Z(n17541) );
  OR U25916 ( .A(n17544), .B(n17545), .Z(n17540) );
  NAND U25917 ( .A(n17546), .B(n17547), .Z(n17438) );
  OR U25918 ( .A(n17548), .B(n17549), .Z(n17547) );
  OR U25919 ( .A(n17550), .B(n17551), .Z(n17546) );
  ANDN U25920 ( .B(n17552), .A(n17553), .Z(n17439) );
  IV U25921 ( .A(n17554), .Z(n17552) );
  XNOR U25922 ( .A(n17519), .B(n17518), .Z(N63842) );
  XOR U25923 ( .A(n17538), .B(n17537), .Z(n17518) );
  XNOR U25924 ( .A(n17553), .B(n17554), .Z(n17537) );
  XNOR U25925 ( .A(n17548), .B(n17549), .Z(n17554) );
  XNOR U25926 ( .A(n17550), .B(n17551), .Z(n17549) );
  XNOR U25927 ( .A(y[6013]), .B(x[6013]), .Z(n17551) );
  XNOR U25928 ( .A(y[6014]), .B(x[6014]), .Z(n17550) );
  XNOR U25929 ( .A(y[6012]), .B(x[6012]), .Z(n17548) );
  XNOR U25930 ( .A(n17542), .B(n17543), .Z(n17553) );
  XNOR U25931 ( .A(y[6009]), .B(x[6009]), .Z(n17543) );
  XNOR U25932 ( .A(n17544), .B(n17545), .Z(n17542) );
  XNOR U25933 ( .A(y[6010]), .B(x[6010]), .Z(n17545) );
  XNOR U25934 ( .A(y[6011]), .B(x[6011]), .Z(n17544) );
  XNOR U25935 ( .A(n17535), .B(n17534), .Z(n17538) );
  XNOR U25936 ( .A(n17530), .B(n17531), .Z(n17534) );
  XNOR U25937 ( .A(y[6006]), .B(x[6006]), .Z(n17531) );
  XNOR U25938 ( .A(n17532), .B(n17533), .Z(n17530) );
  XNOR U25939 ( .A(y[6007]), .B(x[6007]), .Z(n17533) );
  XNOR U25940 ( .A(y[6008]), .B(x[6008]), .Z(n17532) );
  XNOR U25941 ( .A(n17524), .B(n17525), .Z(n17535) );
  XNOR U25942 ( .A(y[6003]), .B(x[6003]), .Z(n17525) );
  XNOR U25943 ( .A(n17526), .B(n17527), .Z(n17524) );
  XNOR U25944 ( .A(y[6004]), .B(x[6004]), .Z(n17527) );
  XNOR U25945 ( .A(y[6005]), .B(x[6005]), .Z(n17526) );
  XOR U25946 ( .A(n17500), .B(n17501), .Z(n17519) );
  XNOR U25947 ( .A(n17516), .B(n17517), .Z(n17501) );
  XNOR U25948 ( .A(n17511), .B(n17512), .Z(n17517) );
  XNOR U25949 ( .A(n17513), .B(n17514), .Z(n17512) );
  XNOR U25950 ( .A(y[6001]), .B(x[6001]), .Z(n17514) );
  XNOR U25951 ( .A(y[6002]), .B(x[6002]), .Z(n17513) );
  XNOR U25952 ( .A(y[6000]), .B(x[6000]), .Z(n17511) );
  XNOR U25953 ( .A(n17505), .B(n17506), .Z(n17516) );
  XNOR U25954 ( .A(y[5997]), .B(x[5997]), .Z(n17506) );
  XNOR U25955 ( .A(n17507), .B(n17508), .Z(n17505) );
  XNOR U25956 ( .A(y[5998]), .B(x[5998]), .Z(n17508) );
  XNOR U25957 ( .A(y[5999]), .B(x[5999]), .Z(n17507) );
  XOR U25958 ( .A(n17499), .B(n17498), .Z(n17500) );
  XNOR U25959 ( .A(n17494), .B(n17495), .Z(n17498) );
  XNOR U25960 ( .A(y[5994]), .B(x[5994]), .Z(n17495) );
  XNOR U25961 ( .A(n17496), .B(n17497), .Z(n17494) );
  XNOR U25962 ( .A(y[5995]), .B(x[5995]), .Z(n17497) );
  XNOR U25963 ( .A(y[5996]), .B(x[5996]), .Z(n17496) );
  XNOR U25964 ( .A(n17488), .B(n17489), .Z(n17499) );
  XNOR U25965 ( .A(y[5991]), .B(x[5991]), .Z(n17489) );
  XNOR U25966 ( .A(n17490), .B(n17491), .Z(n17488) );
  XNOR U25967 ( .A(y[5992]), .B(x[5992]), .Z(n17491) );
  XNOR U25968 ( .A(y[5993]), .B(x[5993]), .Z(n17490) );
  NAND U25969 ( .A(n17555), .B(n17556), .Z(N63833) );
  NANDN U25970 ( .A(n17557), .B(n17558), .Z(n17556) );
  OR U25971 ( .A(n17559), .B(n17560), .Z(n17558) );
  NAND U25972 ( .A(n17559), .B(n17560), .Z(n17555) );
  XOR U25973 ( .A(n17559), .B(n17561), .Z(N63832) );
  XNOR U25974 ( .A(n17557), .B(n17560), .Z(n17561) );
  AND U25975 ( .A(n17562), .B(n17563), .Z(n17560) );
  NANDN U25976 ( .A(n17564), .B(n17565), .Z(n17563) );
  NANDN U25977 ( .A(n17566), .B(n17567), .Z(n17565) );
  NANDN U25978 ( .A(n17567), .B(n17566), .Z(n17562) );
  NAND U25979 ( .A(n17568), .B(n17569), .Z(n17557) );
  NANDN U25980 ( .A(n17570), .B(n17571), .Z(n17569) );
  OR U25981 ( .A(n17572), .B(n17573), .Z(n17571) );
  NAND U25982 ( .A(n17573), .B(n17572), .Z(n17568) );
  AND U25983 ( .A(n17574), .B(n17575), .Z(n17559) );
  NANDN U25984 ( .A(n17576), .B(n17577), .Z(n17575) );
  NANDN U25985 ( .A(n17578), .B(n17579), .Z(n17577) );
  NANDN U25986 ( .A(n17579), .B(n17578), .Z(n17574) );
  XOR U25987 ( .A(n17573), .B(n17580), .Z(N63831) );
  XOR U25988 ( .A(n17570), .B(n17572), .Z(n17580) );
  XNOR U25989 ( .A(n17566), .B(n17581), .Z(n17572) );
  XNOR U25990 ( .A(n17564), .B(n17567), .Z(n17581) );
  NAND U25991 ( .A(n17582), .B(n17583), .Z(n17567) );
  NAND U25992 ( .A(n17584), .B(n17585), .Z(n17583) );
  OR U25993 ( .A(n17586), .B(n17587), .Z(n17584) );
  NANDN U25994 ( .A(n17588), .B(n17586), .Z(n17582) );
  IV U25995 ( .A(n17587), .Z(n17588) );
  NAND U25996 ( .A(n17589), .B(n17590), .Z(n17564) );
  NAND U25997 ( .A(n17591), .B(n17592), .Z(n17590) );
  NANDN U25998 ( .A(n17593), .B(n17594), .Z(n17591) );
  NANDN U25999 ( .A(n17594), .B(n17593), .Z(n17589) );
  AND U26000 ( .A(n17595), .B(n17596), .Z(n17566) );
  NAND U26001 ( .A(n17597), .B(n17598), .Z(n17596) );
  OR U26002 ( .A(n17599), .B(n17600), .Z(n17597) );
  NANDN U26003 ( .A(n17601), .B(n17599), .Z(n17595) );
  NAND U26004 ( .A(n17602), .B(n17603), .Z(n17570) );
  NANDN U26005 ( .A(n17604), .B(n17605), .Z(n17603) );
  OR U26006 ( .A(n17606), .B(n17607), .Z(n17605) );
  NANDN U26007 ( .A(n17608), .B(n17606), .Z(n17602) );
  IV U26008 ( .A(n17607), .Z(n17608) );
  XNOR U26009 ( .A(n17578), .B(n17609), .Z(n17573) );
  XNOR U26010 ( .A(n17576), .B(n17579), .Z(n17609) );
  NAND U26011 ( .A(n17610), .B(n17611), .Z(n17579) );
  NAND U26012 ( .A(n17612), .B(n17613), .Z(n17611) );
  OR U26013 ( .A(n17614), .B(n17615), .Z(n17612) );
  NANDN U26014 ( .A(n17616), .B(n17614), .Z(n17610) );
  IV U26015 ( .A(n17615), .Z(n17616) );
  NAND U26016 ( .A(n17617), .B(n17618), .Z(n17576) );
  NAND U26017 ( .A(n17619), .B(n17620), .Z(n17618) );
  NANDN U26018 ( .A(n17621), .B(n17622), .Z(n17619) );
  NANDN U26019 ( .A(n17622), .B(n17621), .Z(n17617) );
  AND U26020 ( .A(n17623), .B(n17624), .Z(n17578) );
  NAND U26021 ( .A(n17625), .B(n17626), .Z(n17624) );
  OR U26022 ( .A(n17627), .B(n17628), .Z(n17625) );
  NANDN U26023 ( .A(n17629), .B(n17627), .Z(n17623) );
  XNOR U26024 ( .A(n17604), .B(n17630), .Z(N63830) );
  XOR U26025 ( .A(n17606), .B(n17607), .Z(n17630) );
  XNOR U26026 ( .A(n17620), .B(n17631), .Z(n17607) );
  XOR U26027 ( .A(n17621), .B(n17622), .Z(n17631) );
  XOR U26028 ( .A(n17627), .B(n17632), .Z(n17622) );
  XOR U26029 ( .A(n17626), .B(n17629), .Z(n17632) );
  IV U26030 ( .A(n17628), .Z(n17629) );
  NAND U26031 ( .A(n17633), .B(n17634), .Z(n17628) );
  OR U26032 ( .A(n17635), .B(n17636), .Z(n17634) );
  OR U26033 ( .A(n17637), .B(n17638), .Z(n17633) );
  NAND U26034 ( .A(n17639), .B(n17640), .Z(n17626) );
  OR U26035 ( .A(n17641), .B(n17642), .Z(n17640) );
  OR U26036 ( .A(n17643), .B(n17644), .Z(n17639) );
  NOR U26037 ( .A(n17645), .B(n17646), .Z(n17627) );
  ANDN U26038 ( .B(n17647), .A(n17648), .Z(n17621) );
  XNOR U26039 ( .A(n17614), .B(n17649), .Z(n17620) );
  XNOR U26040 ( .A(n17613), .B(n17615), .Z(n17649) );
  NAND U26041 ( .A(n17650), .B(n17651), .Z(n17615) );
  OR U26042 ( .A(n17652), .B(n17653), .Z(n17651) );
  OR U26043 ( .A(n17654), .B(n17655), .Z(n17650) );
  NAND U26044 ( .A(n17656), .B(n17657), .Z(n17613) );
  OR U26045 ( .A(n17658), .B(n17659), .Z(n17657) );
  OR U26046 ( .A(n17660), .B(n17661), .Z(n17656) );
  ANDN U26047 ( .B(n17662), .A(n17663), .Z(n17614) );
  IV U26048 ( .A(n17664), .Z(n17662) );
  ANDN U26049 ( .B(n17665), .A(n17666), .Z(n17606) );
  XOR U26050 ( .A(n17592), .B(n17667), .Z(n17604) );
  XOR U26051 ( .A(n17593), .B(n17594), .Z(n17667) );
  XOR U26052 ( .A(n17599), .B(n17668), .Z(n17594) );
  XOR U26053 ( .A(n17598), .B(n17601), .Z(n17668) );
  IV U26054 ( .A(n17600), .Z(n17601) );
  NAND U26055 ( .A(n17669), .B(n17670), .Z(n17600) );
  OR U26056 ( .A(n17671), .B(n17672), .Z(n17670) );
  OR U26057 ( .A(n17673), .B(n17674), .Z(n17669) );
  NAND U26058 ( .A(n17675), .B(n17676), .Z(n17598) );
  OR U26059 ( .A(n17677), .B(n17678), .Z(n17676) );
  OR U26060 ( .A(n17679), .B(n17680), .Z(n17675) );
  NOR U26061 ( .A(n17681), .B(n17682), .Z(n17599) );
  ANDN U26062 ( .B(n17683), .A(n17684), .Z(n17593) );
  IV U26063 ( .A(n17685), .Z(n17683) );
  XNOR U26064 ( .A(n17586), .B(n17686), .Z(n17592) );
  XNOR U26065 ( .A(n17585), .B(n17587), .Z(n17686) );
  NAND U26066 ( .A(n17687), .B(n17688), .Z(n17587) );
  OR U26067 ( .A(n17689), .B(n17690), .Z(n17688) );
  OR U26068 ( .A(n17691), .B(n17692), .Z(n17687) );
  NAND U26069 ( .A(n17693), .B(n17694), .Z(n17585) );
  OR U26070 ( .A(n17695), .B(n17696), .Z(n17694) );
  OR U26071 ( .A(n17697), .B(n17698), .Z(n17693) );
  ANDN U26072 ( .B(n17699), .A(n17700), .Z(n17586) );
  IV U26073 ( .A(n17701), .Z(n17699) );
  XNOR U26074 ( .A(n17666), .B(n17665), .Z(N63829) );
  XOR U26075 ( .A(n17685), .B(n17684), .Z(n17665) );
  XNOR U26076 ( .A(n17700), .B(n17701), .Z(n17684) );
  XNOR U26077 ( .A(n17695), .B(n17696), .Z(n17701) );
  XNOR U26078 ( .A(n17697), .B(n17698), .Z(n17696) );
  XNOR U26079 ( .A(y[5989]), .B(x[5989]), .Z(n17698) );
  XNOR U26080 ( .A(y[5990]), .B(x[5990]), .Z(n17697) );
  XNOR U26081 ( .A(y[5988]), .B(x[5988]), .Z(n17695) );
  XNOR U26082 ( .A(n17689), .B(n17690), .Z(n17700) );
  XNOR U26083 ( .A(y[5985]), .B(x[5985]), .Z(n17690) );
  XNOR U26084 ( .A(n17691), .B(n17692), .Z(n17689) );
  XNOR U26085 ( .A(y[5986]), .B(x[5986]), .Z(n17692) );
  XNOR U26086 ( .A(y[5987]), .B(x[5987]), .Z(n17691) );
  XNOR U26087 ( .A(n17682), .B(n17681), .Z(n17685) );
  XNOR U26088 ( .A(n17677), .B(n17678), .Z(n17681) );
  XNOR U26089 ( .A(y[5982]), .B(x[5982]), .Z(n17678) );
  XNOR U26090 ( .A(n17679), .B(n17680), .Z(n17677) );
  XNOR U26091 ( .A(y[5983]), .B(x[5983]), .Z(n17680) );
  XNOR U26092 ( .A(y[5984]), .B(x[5984]), .Z(n17679) );
  XNOR U26093 ( .A(n17671), .B(n17672), .Z(n17682) );
  XNOR U26094 ( .A(y[5979]), .B(x[5979]), .Z(n17672) );
  XNOR U26095 ( .A(n17673), .B(n17674), .Z(n17671) );
  XNOR U26096 ( .A(y[5980]), .B(x[5980]), .Z(n17674) );
  XNOR U26097 ( .A(y[5981]), .B(x[5981]), .Z(n17673) );
  XOR U26098 ( .A(n17647), .B(n17648), .Z(n17666) );
  XNOR U26099 ( .A(n17663), .B(n17664), .Z(n17648) );
  XNOR U26100 ( .A(n17658), .B(n17659), .Z(n17664) );
  XNOR U26101 ( .A(n17660), .B(n17661), .Z(n17659) );
  XNOR U26102 ( .A(y[5977]), .B(x[5977]), .Z(n17661) );
  XNOR U26103 ( .A(y[5978]), .B(x[5978]), .Z(n17660) );
  XNOR U26104 ( .A(y[5976]), .B(x[5976]), .Z(n17658) );
  XNOR U26105 ( .A(n17652), .B(n17653), .Z(n17663) );
  XNOR U26106 ( .A(y[5973]), .B(x[5973]), .Z(n17653) );
  XNOR U26107 ( .A(n17654), .B(n17655), .Z(n17652) );
  XNOR U26108 ( .A(y[5974]), .B(x[5974]), .Z(n17655) );
  XNOR U26109 ( .A(y[5975]), .B(x[5975]), .Z(n17654) );
  XOR U26110 ( .A(n17646), .B(n17645), .Z(n17647) );
  XNOR U26111 ( .A(n17641), .B(n17642), .Z(n17645) );
  XNOR U26112 ( .A(y[5970]), .B(x[5970]), .Z(n17642) );
  XNOR U26113 ( .A(n17643), .B(n17644), .Z(n17641) );
  XNOR U26114 ( .A(y[5971]), .B(x[5971]), .Z(n17644) );
  XNOR U26115 ( .A(y[5972]), .B(x[5972]), .Z(n17643) );
  XNOR U26116 ( .A(n17635), .B(n17636), .Z(n17646) );
  XNOR U26117 ( .A(y[5967]), .B(x[5967]), .Z(n17636) );
  XNOR U26118 ( .A(n17637), .B(n17638), .Z(n17635) );
  XNOR U26119 ( .A(y[5968]), .B(x[5968]), .Z(n17638) );
  XNOR U26120 ( .A(y[5969]), .B(x[5969]), .Z(n17637) );
  NAND U26121 ( .A(n17702), .B(n17703), .Z(N63820) );
  NANDN U26122 ( .A(n17704), .B(n17705), .Z(n17703) );
  OR U26123 ( .A(n17706), .B(n17707), .Z(n17705) );
  NAND U26124 ( .A(n17706), .B(n17707), .Z(n17702) );
  XOR U26125 ( .A(n17706), .B(n17708), .Z(N63819) );
  XNOR U26126 ( .A(n17704), .B(n17707), .Z(n17708) );
  AND U26127 ( .A(n17709), .B(n17710), .Z(n17707) );
  NANDN U26128 ( .A(n17711), .B(n17712), .Z(n17710) );
  NANDN U26129 ( .A(n17713), .B(n17714), .Z(n17712) );
  NANDN U26130 ( .A(n17714), .B(n17713), .Z(n17709) );
  NAND U26131 ( .A(n17715), .B(n17716), .Z(n17704) );
  NANDN U26132 ( .A(n17717), .B(n17718), .Z(n17716) );
  OR U26133 ( .A(n17719), .B(n17720), .Z(n17718) );
  NAND U26134 ( .A(n17720), .B(n17719), .Z(n17715) );
  AND U26135 ( .A(n17721), .B(n17722), .Z(n17706) );
  NANDN U26136 ( .A(n17723), .B(n17724), .Z(n17722) );
  NANDN U26137 ( .A(n17725), .B(n17726), .Z(n17724) );
  NANDN U26138 ( .A(n17726), .B(n17725), .Z(n17721) );
  XOR U26139 ( .A(n17720), .B(n17727), .Z(N63818) );
  XOR U26140 ( .A(n17717), .B(n17719), .Z(n17727) );
  XNOR U26141 ( .A(n17713), .B(n17728), .Z(n17719) );
  XNOR U26142 ( .A(n17711), .B(n17714), .Z(n17728) );
  NAND U26143 ( .A(n17729), .B(n17730), .Z(n17714) );
  NAND U26144 ( .A(n17731), .B(n17732), .Z(n17730) );
  OR U26145 ( .A(n17733), .B(n17734), .Z(n17731) );
  NANDN U26146 ( .A(n17735), .B(n17733), .Z(n17729) );
  IV U26147 ( .A(n17734), .Z(n17735) );
  NAND U26148 ( .A(n17736), .B(n17737), .Z(n17711) );
  NAND U26149 ( .A(n17738), .B(n17739), .Z(n17737) );
  NANDN U26150 ( .A(n17740), .B(n17741), .Z(n17738) );
  NANDN U26151 ( .A(n17741), .B(n17740), .Z(n17736) );
  AND U26152 ( .A(n17742), .B(n17743), .Z(n17713) );
  NAND U26153 ( .A(n17744), .B(n17745), .Z(n17743) );
  OR U26154 ( .A(n17746), .B(n17747), .Z(n17744) );
  NANDN U26155 ( .A(n17748), .B(n17746), .Z(n17742) );
  NAND U26156 ( .A(n17749), .B(n17750), .Z(n17717) );
  NANDN U26157 ( .A(n17751), .B(n17752), .Z(n17750) );
  OR U26158 ( .A(n17753), .B(n17754), .Z(n17752) );
  NANDN U26159 ( .A(n17755), .B(n17753), .Z(n17749) );
  IV U26160 ( .A(n17754), .Z(n17755) );
  XNOR U26161 ( .A(n17725), .B(n17756), .Z(n17720) );
  XNOR U26162 ( .A(n17723), .B(n17726), .Z(n17756) );
  NAND U26163 ( .A(n17757), .B(n17758), .Z(n17726) );
  NAND U26164 ( .A(n17759), .B(n17760), .Z(n17758) );
  OR U26165 ( .A(n17761), .B(n17762), .Z(n17759) );
  NANDN U26166 ( .A(n17763), .B(n17761), .Z(n17757) );
  IV U26167 ( .A(n17762), .Z(n17763) );
  NAND U26168 ( .A(n17764), .B(n17765), .Z(n17723) );
  NAND U26169 ( .A(n17766), .B(n17767), .Z(n17765) );
  NANDN U26170 ( .A(n17768), .B(n17769), .Z(n17766) );
  NANDN U26171 ( .A(n17769), .B(n17768), .Z(n17764) );
  AND U26172 ( .A(n17770), .B(n17771), .Z(n17725) );
  NAND U26173 ( .A(n17772), .B(n17773), .Z(n17771) );
  OR U26174 ( .A(n17774), .B(n17775), .Z(n17772) );
  NANDN U26175 ( .A(n17776), .B(n17774), .Z(n17770) );
  XNOR U26176 ( .A(n17751), .B(n17777), .Z(N63817) );
  XOR U26177 ( .A(n17753), .B(n17754), .Z(n17777) );
  XNOR U26178 ( .A(n17767), .B(n17778), .Z(n17754) );
  XOR U26179 ( .A(n17768), .B(n17769), .Z(n17778) );
  XOR U26180 ( .A(n17774), .B(n17779), .Z(n17769) );
  XOR U26181 ( .A(n17773), .B(n17776), .Z(n17779) );
  IV U26182 ( .A(n17775), .Z(n17776) );
  NAND U26183 ( .A(n17780), .B(n17781), .Z(n17775) );
  OR U26184 ( .A(n17782), .B(n17783), .Z(n17781) );
  OR U26185 ( .A(n17784), .B(n17785), .Z(n17780) );
  NAND U26186 ( .A(n17786), .B(n17787), .Z(n17773) );
  OR U26187 ( .A(n17788), .B(n17789), .Z(n17787) );
  OR U26188 ( .A(n17790), .B(n17791), .Z(n17786) );
  NOR U26189 ( .A(n17792), .B(n17793), .Z(n17774) );
  ANDN U26190 ( .B(n17794), .A(n17795), .Z(n17768) );
  XNOR U26191 ( .A(n17761), .B(n17796), .Z(n17767) );
  XNOR U26192 ( .A(n17760), .B(n17762), .Z(n17796) );
  NAND U26193 ( .A(n17797), .B(n17798), .Z(n17762) );
  OR U26194 ( .A(n17799), .B(n17800), .Z(n17798) );
  OR U26195 ( .A(n17801), .B(n17802), .Z(n17797) );
  NAND U26196 ( .A(n17803), .B(n17804), .Z(n17760) );
  OR U26197 ( .A(n17805), .B(n17806), .Z(n17804) );
  OR U26198 ( .A(n17807), .B(n17808), .Z(n17803) );
  ANDN U26199 ( .B(n17809), .A(n17810), .Z(n17761) );
  IV U26200 ( .A(n17811), .Z(n17809) );
  ANDN U26201 ( .B(n17812), .A(n17813), .Z(n17753) );
  XOR U26202 ( .A(n17739), .B(n17814), .Z(n17751) );
  XOR U26203 ( .A(n17740), .B(n17741), .Z(n17814) );
  XOR U26204 ( .A(n17746), .B(n17815), .Z(n17741) );
  XOR U26205 ( .A(n17745), .B(n17748), .Z(n17815) );
  IV U26206 ( .A(n17747), .Z(n17748) );
  NAND U26207 ( .A(n17816), .B(n17817), .Z(n17747) );
  OR U26208 ( .A(n17818), .B(n17819), .Z(n17817) );
  OR U26209 ( .A(n17820), .B(n17821), .Z(n17816) );
  NAND U26210 ( .A(n17822), .B(n17823), .Z(n17745) );
  OR U26211 ( .A(n17824), .B(n17825), .Z(n17823) );
  OR U26212 ( .A(n17826), .B(n17827), .Z(n17822) );
  NOR U26213 ( .A(n17828), .B(n17829), .Z(n17746) );
  ANDN U26214 ( .B(n17830), .A(n17831), .Z(n17740) );
  IV U26215 ( .A(n17832), .Z(n17830) );
  XNOR U26216 ( .A(n17733), .B(n17833), .Z(n17739) );
  XNOR U26217 ( .A(n17732), .B(n17734), .Z(n17833) );
  NAND U26218 ( .A(n17834), .B(n17835), .Z(n17734) );
  OR U26219 ( .A(n17836), .B(n17837), .Z(n17835) );
  OR U26220 ( .A(n17838), .B(n17839), .Z(n17834) );
  NAND U26221 ( .A(n17840), .B(n17841), .Z(n17732) );
  OR U26222 ( .A(n17842), .B(n17843), .Z(n17841) );
  OR U26223 ( .A(n17844), .B(n17845), .Z(n17840) );
  ANDN U26224 ( .B(n17846), .A(n17847), .Z(n17733) );
  IV U26225 ( .A(n17848), .Z(n17846) );
  XNOR U26226 ( .A(n17813), .B(n17812), .Z(N63816) );
  XOR U26227 ( .A(n17832), .B(n17831), .Z(n17812) );
  XNOR U26228 ( .A(n17847), .B(n17848), .Z(n17831) );
  XNOR U26229 ( .A(n17842), .B(n17843), .Z(n17848) );
  XNOR U26230 ( .A(n17844), .B(n17845), .Z(n17843) );
  XNOR U26231 ( .A(y[5965]), .B(x[5965]), .Z(n17845) );
  XNOR U26232 ( .A(y[5966]), .B(x[5966]), .Z(n17844) );
  XNOR U26233 ( .A(y[5964]), .B(x[5964]), .Z(n17842) );
  XNOR U26234 ( .A(n17836), .B(n17837), .Z(n17847) );
  XNOR U26235 ( .A(y[5961]), .B(x[5961]), .Z(n17837) );
  XNOR U26236 ( .A(n17838), .B(n17839), .Z(n17836) );
  XNOR U26237 ( .A(y[5962]), .B(x[5962]), .Z(n17839) );
  XNOR U26238 ( .A(y[5963]), .B(x[5963]), .Z(n17838) );
  XNOR U26239 ( .A(n17829), .B(n17828), .Z(n17832) );
  XNOR U26240 ( .A(n17824), .B(n17825), .Z(n17828) );
  XNOR U26241 ( .A(y[5958]), .B(x[5958]), .Z(n17825) );
  XNOR U26242 ( .A(n17826), .B(n17827), .Z(n17824) );
  XNOR U26243 ( .A(y[5959]), .B(x[5959]), .Z(n17827) );
  XNOR U26244 ( .A(y[5960]), .B(x[5960]), .Z(n17826) );
  XNOR U26245 ( .A(n17818), .B(n17819), .Z(n17829) );
  XNOR U26246 ( .A(y[5955]), .B(x[5955]), .Z(n17819) );
  XNOR U26247 ( .A(n17820), .B(n17821), .Z(n17818) );
  XNOR U26248 ( .A(y[5956]), .B(x[5956]), .Z(n17821) );
  XNOR U26249 ( .A(y[5957]), .B(x[5957]), .Z(n17820) );
  XOR U26250 ( .A(n17794), .B(n17795), .Z(n17813) );
  XNOR U26251 ( .A(n17810), .B(n17811), .Z(n17795) );
  XNOR U26252 ( .A(n17805), .B(n17806), .Z(n17811) );
  XNOR U26253 ( .A(n17807), .B(n17808), .Z(n17806) );
  XNOR U26254 ( .A(y[5953]), .B(x[5953]), .Z(n17808) );
  XNOR U26255 ( .A(y[5954]), .B(x[5954]), .Z(n17807) );
  XNOR U26256 ( .A(y[5952]), .B(x[5952]), .Z(n17805) );
  XNOR U26257 ( .A(n17799), .B(n17800), .Z(n17810) );
  XNOR U26258 ( .A(y[5949]), .B(x[5949]), .Z(n17800) );
  XNOR U26259 ( .A(n17801), .B(n17802), .Z(n17799) );
  XNOR U26260 ( .A(y[5950]), .B(x[5950]), .Z(n17802) );
  XNOR U26261 ( .A(y[5951]), .B(x[5951]), .Z(n17801) );
  XOR U26262 ( .A(n17793), .B(n17792), .Z(n17794) );
  XNOR U26263 ( .A(n17788), .B(n17789), .Z(n17792) );
  XNOR U26264 ( .A(y[5946]), .B(x[5946]), .Z(n17789) );
  XNOR U26265 ( .A(n17790), .B(n17791), .Z(n17788) );
  XNOR U26266 ( .A(y[5947]), .B(x[5947]), .Z(n17791) );
  XNOR U26267 ( .A(y[5948]), .B(x[5948]), .Z(n17790) );
  XNOR U26268 ( .A(n17782), .B(n17783), .Z(n17793) );
  XNOR U26269 ( .A(y[5943]), .B(x[5943]), .Z(n17783) );
  XNOR U26270 ( .A(n17784), .B(n17785), .Z(n17782) );
  XNOR U26271 ( .A(y[5944]), .B(x[5944]), .Z(n17785) );
  XNOR U26272 ( .A(y[5945]), .B(x[5945]), .Z(n17784) );
  NAND U26273 ( .A(n17849), .B(n17850), .Z(N63807) );
  NANDN U26274 ( .A(n17851), .B(n17852), .Z(n17850) );
  OR U26275 ( .A(n17853), .B(n17854), .Z(n17852) );
  NAND U26276 ( .A(n17853), .B(n17854), .Z(n17849) );
  XOR U26277 ( .A(n17853), .B(n17855), .Z(N63806) );
  XNOR U26278 ( .A(n17851), .B(n17854), .Z(n17855) );
  AND U26279 ( .A(n17856), .B(n17857), .Z(n17854) );
  NANDN U26280 ( .A(n17858), .B(n17859), .Z(n17857) );
  NANDN U26281 ( .A(n17860), .B(n17861), .Z(n17859) );
  NANDN U26282 ( .A(n17861), .B(n17860), .Z(n17856) );
  NAND U26283 ( .A(n17862), .B(n17863), .Z(n17851) );
  NANDN U26284 ( .A(n17864), .B(n17865), .Z(n17863) );
  OR U26285 ( .A(n17866), .B(n17867), .Z(n17865) );
  NAND U26286 ( .A(n17867), .B(n17866), .Z(n17862) );
  AND U26287 ( .A(n17868), .B(n17869), .Z(n17853) );
  NANDN U26288 ( .A(n17870), .B(n17871), .Z(n17869) );
  NANDN U26289 ( .A(n17872), .B(n17873), .Z(n17871) );
  NANDN U26290 ( .A(n17873), .B(n17872), .Z(n17868) );
  XOR U26291 ( .A(n17867), .B(n17874), .Z(N63805) );
  XOR U26292 ( .A(n17864), .B(n17866), .Z(n17874) );
  XNOR U26293 ( .A(n17860), .B(n17875), .Z(n17866) );
  XNOR U26294 ( .A(n17858), .B(n17861), .Z(n17875) );
  NAND U26295 ( .A(n17876), .B(n17877), .Z(n17861) );
  NAND U26296 ( .A(n17878), .B(n17879), .Z(n17877) );
  OR U26297 ( .A(n17880), .B(n17881), .Z(n17878) );
  NANDN U26298 ( .A(n17882), .B(n17880), .Z(n17876) );
  IV U26299 ( .A(n17881), .Z(n17882) );
  NAND U26300 ( .A(n17883), .B(n17884), .Z(n17858) );
  NAND U26301 ( .A(n17885), .B(n17886), .Z(n17884) );
  NANDN U26302 ( .A(n17887), .B(n17888), .Z(n17885) );
  NANDN U26303 ( .A(n17888), .B(n17887), .Z(n17883) );
  AND U26304 ( .A(n17889), .B(n17890), .Z(n17860) );
  NAND U26305 ( .A(n17891), .B(n17892), .Z(n17890) );
  OR U26306 ( .A(n17893), .B(n17894), .Z(n17891) );
  NANDN U26307 ( .A(n17895), .B(n17893), .Z(n17889) );
  NAND U26308 ( .A(n17896), .B(n17897), .Z(n17864) );
  NANDN U26309 ( .A(n17898), .B(n17899), .Z(n17897) );
  OR U26310 ( .A(n17900), .B(n17901), .Z(n17899) );
  NANDN U26311 ( .A(n17902), .B(n17900), .Z(n17896) );
  IV U26312 ( .A(n17901), .Z(n17902) );
  XNOR U26313 ( .A(n17872), .B(n17903), .Z(n17867) );
  XNOR U26314 ( .A(n17870), .B(n17873), .Z(n17903) );
  NAND U26315 ( .A(n17904), .B(n17905), .Z(n17873) );
  NAND U26316 ( .A(n17906), .B(n17907), .Z(n17905) );
  OR U26317 ( .A(n17908), .B(n17909), .Z(n17906) );
  NANDN U26318 ( .A(n17910), .B(n17908), .Z(n17904) );
  IV U26319 ( .A(n17909), .Z(n17910) );
  NAND U26320 ( .A(n17911), .B(n17912), .Z(n17870) );
  NAND U26321 ( .A(n17913), .B(n17914), .Z(n17912) );
  NANDN U26322 ( .A(n17915), .B(n17916), .Z(n17913) );
  NANDN U26323 ( .A(n17916), .B(n17915), .Z(n17911) );
  AND U26324 ( .A(n17917), .B(n17918), .Z(n17872) );
  NAND U26325 ( .A(n17919), .B(n17920), .Z(n17918) );
  OR U26326 ( .A(n17921), .B(n17922), .Z(n17919) );
  NANDN U26327 ( .A(n17923), .B(n17921), .Z(n17917) );
  XNOR U26328 ( .A(n17898), .B(n17924), .Z(N63804) );
  XOR U26329 ( .A(n17900), .B(n17901), .Z(n17924) );
  XNOR U26330 ( .A(n17914), .B(n17925), .Z(n17901) );
  XOR U26331 ( .A(n17915), .B(n17916), .Z(n17925) );
  XOR U26332 ( .A(n17921), .B(n17926), .Z(n17916) );
  XOR U26333 ( .A(n17920), .B(n17923), .Z(n17926) );
  IV U26334 ( .A(n17922), .Z(n17923) );
  NAND U26335 ( .A(n17927), .B(n17928), .Z(n17922) );
  OR U26336 ( .A(n17929), .B(n17930), .Z(n17928) );
  OR U26337 ( .A(n17931), .B(n17932), .Z(n17927) );
  NAND U26338 ( .A(n17933), .B(n17934), .Z(n17920) );
  OR U26339 ( .A(n17935), .B(n17936), .Z(n17934) );
  OR U26340 ( .A(n17937), .B(n17938), .Z(n17933) );
  NOR U26341 ( .A(n17939), .B(n17940), .Z(n17921) );
  ANDN U26342 ( .B(n17941), .A(n17942), .Z(n17915) );
  XNOR U26343 ( .A(n17908), .B(n17943), .Z(n17914) );
  XNOR U26344 ( .A(n17907), .B(n17909), .Z(n17943) );
  NAND U26345 ( .A(n17944), .B(n17945), .Z(n17909) );
  OR U26346 ( .A(n17946), .B(n17947), .Z(n17945) );
  OR U26347 ( .A(n17948), .B(n17949), .Z(n17944) );
  NAND U26348 ( .A(n17950), .B(n17951), .Z(n17907) );
  OR U26349 ( .A(n17952), .B(n17953), .Z(n17951) );
  OR U26350 ( .A(n17954), .B(n17955), .Z(n17950) );
  ANDN U26351 ( .B(n17956), .A(n17957), .Z(n17908) );
  IV U26352 ( .A(n17958), .Z(n17956) );
  ANDN U26353 ( .B(n17959), .A(n17960), .Z(n17900) );
  XOR U26354 ( .A(n17886), .B(n17961), .Z(n17898) );
  XOR U26355 ( .A(n17887), .B(n17888), .Z(n17961) );
  XOR U26356 ( .A(n17893), .B(n17962), .Z(n17888) );
  XOR U26357 ( .A(n17892), .B(n17895), .Z(n17962) );
  IV U26358 ( .A(n17894), .Z(n17895) );
  NAND U26359 ( .A(n17963), .B(n17964), .Z(n17894) );
  OR U26360 ( .A(n17965), .B(n17966), .Z(n17964) );
  OR U26361 ( .A(n17967), .B(n17968), .Z(n17963) );
  NAND U26362 ( .A(n17969), .B(n17970), .Z(n17892) );
  OR U26363 ( .A(n17971), .B(n17972), .Z(n17970) );
  OR U26364 ( .A(n17973), .B(n17974), .Z(n17969) );
  NOR U26365 ( .A(n17975), .B(n17976), .Z(n17893) );
  ANDN U26366 ( .B(n17977), .A(n17978), .Z(n17887) );
  IV U26367 ( .A(n17979), .Z(n17977) );
  XNOR U26368 ( .A(n17880), .B(n17980), .Z(n17886) );
  XNOR U26369 ( .A(n17879), .B(n17881), .Z(n17980) );
  NAND U26370 ( .A(n17981), .B(n17982), .Z(n17881) );
  OR U26371 ( .A(n17983), .B(n17984), .Z(n17982) );
  OR U26372 ( .A(n17985), .B(n17986), .Z(n17981) );
  NAND U26373 ( .A(n17987), .B(n17988), .Z(n17879) );
  OR U26374 ( .A(n17989), .B(n17990), .Z(n17988) );
  OR U26375 ( .A(n17991), .B(n17992), .Z(n17987) );
  ANDN U26376 ( .B(n17993), .A(n17994), .Z(n17880) );
  IV U26377 ( .A(n17995), .Z(n17993) );
  XNOR U26378 ( .A(n17960), .B(n17959), .Z(N63803) );
  XOR U26379 ( .A(n17979), .B(n17978), .Z(n17959) );
  XNOR U26380 ( .A(n17994), .B(n17995), .Z(n17978) );
  XNOR U26381 ( .A(n17989), .B(n17990), .Z(n17995) );
  XNOR U26382 ( .A(n17991), .B(n17992), .Z(n17990) );
  XNOR U26383 ( .A(y[5941]), .B(x[5941]), .Z(n17992) );
  XNOR U26384 ( .A(y[5942]), .B(x[5942]), .Z(n17991) );
  XNOR U26385 ( .A(y[5940]), .B(x[5940]), .Z(n17989) );
  XNOR U26386 ( .A(n17983), .B(n17984), .Z(n17994) );
  XNOR U26387 ( .A(y[5937]), .B(x[5937]), .Z(n17984) );
  XNOR U26388 ( .A(n17985), .B(n17986), .Z(n17983) );
  XNOR U26389 ( .A(y[5938]), .B(x[5938]), .Z(n17986) );
  XNOR U26390 ( .A(y[5939]), .B(x[5939]), .Z(n17985) );
  XNOR U26391 ( .A(n17976), .B(n17975), .Z(n17979) );
  XNOR U26392 ( .A(n17971), .B(n17972), .Z(n17975) );
  XNOR U26393 ( .A(y[5934]), .B(x[5934]), .Z(n17972) );
  XNOR U26394 ( .A(n17973), .B(n17974), .Z(n17971) );
  XNOR U26395 ( .A(y[5935]), .B(x[5935]), .Z(n17974) );
  XNOR U26396 ( .A(y[5936]), .B(x[5936]), .Z(n17973) );
  XNOR U26397 ( .A(n17965), .B(n17966), .Z(n17976) );
  XNOR U26398 ( .A(y[5931]), .B(x[5931]), .Z(n17966) );
  XNOR U26399 ( .A(n17967), .B(n17968), .Z(n17965) );
  XNOR U26400 ( .A(y[5932]), .B(x[5932]), .Z(n17968) );
  XNOR U26401 ( .A(y[5933]), .B(x[5933]), .Z(n17967) );
  XOR U26402 ( .A(n17941), .B(n17942), .Z(n17960) );
  XNOR U26403 ( .A(n17957), .B(n17958), .Z(n17942) );
  XNOR U26404 ( .A(n17952), .B(n17953), .Z(n17958) );
  XNOR U26405 ( .A(n17954), .B(n17955), .Z(n17953) );
  XNOR U26406 ( .A(y[5929]), .B(x[5929]), .Z(n17955) );
  XNOR U26407 ( .A(y[5930]), .B(x[5930]), .Z(n17954) );
  XNOR U26408 ( .A(y[5928]), .B(x[5928]), .Z(n17952) );
  XNOR U26409 ( .A(n17946), .B(n17947), .Z(n17957) );
  XNOR U26410 ( .A(y[5925]), .B(x[5925]), .Z(n17947) );
  XNOR U26411 ( .A(n17948), .B(n17949), .Z(n17946) );
  XNOR U26412 ( .A(y[5926]), .B(x[5926]), .Z(n17949) );
  XNOR U26413 ( .A(y[5927]), .B(x[5927]), .Z(n17948) );
  XOR U26414 ( .A(n17940), .B(n17939), .Z(n17941) );
  XNOR U26415 ( .A(n17935), .B(n17936), .Z(n17939) );
  XNOR U26416 ( .A(y[5922]), .B(x[5922]), .Z(n17936) );
  XNOR U26417 ( .A(n17937), .B(n17938), .Z(n17935) );
  XNOR U26418 ( .A(y[5923]), .B(x[5923]), .Z(n17938) );
  XNOR U26419 ( .A(y[5924]), .B(x[5924]), .Z(n17937) );
  XNOR U26420 ( .A(n17929), .B(n17930), .Z(n17940) );
  XNOR U26421 ( .A(y[5919]), .B(x[5919]), .Z(n17930) );
  XNOR U26422 ( .A(n17931), .B(n17932), .Z(n17929) );
  XNOR U26423 ( .A(y[5920]), .B(x[5920]), .Z(n17932) );
  XNOR U26424 ( .A(y[5921]), .B(x[5921]), .Z(n17931) );
  NAND U26425 ( .A(n17996), .B(n17997), .Z(N63794) );
  NANDN U26426 ( .A(n17998), .B(n17999), .Z(n17997) );
  OR U26427 ( .A(n18000), .B(n18001), .Z(n17999) );
  NAND U26428 ( .A(n18000), .B(n18001), .Z(n17996) );
  XOR U26429 ( .A(n18000), .B(n18002), .Z(N63793) );
  XNOR U26430 ( .A(n17998), .B(n18001), .Z(n18002) );
  AND U26431 ( .A(n18003), .B(n18004), .Z(n18001) );
  NANDN U26432 ( .A(n18005), .B(n18006), .Z(n18004) );
  NANDN U26433 ( .A(n18007), .B(n18008), .Z(n18006) );
  NANDN U26434 ( .A(n18008), .B(n18007), .Z(n18003) );
  NAND U26435 ( .A(n18009), .B(n18010), .Z(n17998) );
  NANDN U26436 ( .A(n18011), .B(n18012), .Z(n18010) );
  OR U26437 ( .A(n18013), .B(n18014), .Z(n18012) );
  NAND U26438 ( .A(n18014), .B(n18013), .Z(n18009) );
  AND U26439 ( .A(n18015), .B(n18016), .Z(n18000) );
  NANDN U26440 ( .A(n18017), .B(n18018), .Z(n18016) );
  NANDN U26441 ( .A(n18019), .B(n18020), .Z(n18018) );
  NANDN U26442 ( .A(n18020), .B(n18019), .Z(n18015) );
  XOR U26443 ( .A(n18014), .B(n18021), .Z(N63792) );
  XOR U26444 ( .A(n18011), .B(n18013), .Z(n18021) );
  XNOR U26445 ( .A(n18007), .B(n18022), .Z(n18013) );
  XNOR U26446 ( .A(n18005), .B(n18008), .Z(n18022) );
  NAND U26447 ( .A(n18023), .B(n18024), .Z(n18008) );
  NAND U26448 ( .A(n18025), .B(n18026), .Z(n18024) );
  OR U26449 ( .A(n18027), .B(n18028), .Z(n18025) );
  NANDN U26450 ( .A(n18029), .B(n18027), .Z(n18023) );
  IV U26451 ( .A(n18028), .Z(n18029) );
  NAND U26452 ( .A(n18030), .B(n18031), .Z(n18005) );
  NAND U26453 ( .A(n18032), .B(n18033), .Z(n18031) );
  NANDN U26454 ( .A(n18034), .B(n18035), .Z(n18032) );
  NANDN U26455 ( .A(n18035), .B(n18034), .Z(n18030) );
  AND U26456 ( .A(n18036), .B(n18037), .Z(n18007) );
  NAND U26457 ( .A(n18038), .B(n18039), .Z(n18037) );
  OR U26458 ( .A(n18040), .B(n18041), .Z(n18038) );
  NANDN U26459 ( .A(n18042), .B(n18040), .Z(n18036) );
  NAND U26460 ( .A(n18043), .B(n18044), .Z(n18011) );
  NANDN U26461 ( .A(n18045), .B(n18046), .Z(n18044) );
  OR U26462 ( .A(n18047), .B(n18048), .Z(n18046) );
  NANDN U26463 ( .A(n18049), .B(n18047), .Z(n18043) );
  IV U26464 ( .A(n18048), .Z(n18049) );
  XNOR U26465 ( .A(n18019), .B(n18050), .Z(n18014) );
  XNOR U26466 ( .A(n18017), .B(n18020), .Z(n18050) );
  NAND U26467 ( .A(n18051), .B(n18052), .Z(n18020) );
  NAND U26468 ( .A(n18053), .B(n18054), .Z(n18052) );
  OR U26469 ( .A(n18055), .B(n18056), .Z(n18053) );
  NANDN U26470 ( .A(n18057), .B(n18055), .Z(n18051) );
  IV U26471 ( .A(n18056), .Z(n18057) );
  NAND U26472 ( .A(n18058), .B(n18059), .Z(n18017) );
  NAND U26473 ( .A(n18060), .B(n18061), .Z(n18059) );
  NANDN U26474 ( .A(n18062), .B(n18063), .Z(n18060) );
  NANDN U26475 ( .A(n18063), .B(n18062), .Z(n18058) );
  AND U26476 ( .A(n18064), .B(n18065), .Z(n18019) );
  NAND U26477 ( .A(n18066), .B(n18067), .Z(n18065) );
  OR U26478 ( .A(n18068), .B(n18069), .Z(n18066) );
  NANDN U26479 ( .A(n18070), .B(n18068), .Z(n18064) );
  XNOR U26480 ( .A(n18045), .B(n18071), .Z(N63791) );
  XOR U26481 ( .A(n18047), .B(n18048), .Z(n18071) );
  XNOR U26482 ( .A(n18061), .B(n18072), .Z(n18048) );
  XOR U26483 ( .A(n18062), .B(n18063), .Z(n18072) );
  XOR U26484 ( .A(n18068), .B(n18073), .Z(n18063) );
  XOR U26485 ( .A(n18067), .B(n18070), .Z(n18073) );
  IV U26486 ( .A(n18069), .Z(n18070) );
  NAND U26487 ( .A(n18074), .B(n18075), .Z(n18069) );
  OR U26488 ( .A(n18076), .B(n18077), .Z(n18075) );
  OR U26489 ( .A(n18078), .B(n18079), .Z(n18074) );
  NAND U26490 ( .A(n18080), .B(n18081), .Z(n18067) );
  OR U26491 ( .A(n18082), .B(n18083), .Z(n18081) );
  OR U26492 ( .A(n18084), .B(n18085), .Z(n18080) );
  NOR U26493 ( .A(n18086), .B(n18087), .Z(n18068) );
  ANDN U26494 ( .B(n18088), .A(n18089), .Z(n18062) );
  XNOR U26495 ( .A(n18055), .B(n18090), .Z(n18061) );
  XNOR U26496 ( .A(n18054), .B(n18056), .Z(n18090) );
  NAND U26497 ( .A(n18091), .B(n18092), .Z(n18056) );
  OR U26498 ( .A(n18093), .B(n18094), .Z(n18092) );
  OR U26499 ( .A(n18095), .B(n18096), .Z(n18091) );
  NAND U26500 ( .A(n18097), .B(n18098), .Z(n18054) );
  OR U26501 ( .A(n18099), .B(n18100), .Z(n18098) );
  OR U26502 ( .A(n18101), .B(n18102), .Z(n18097) );
  ANDN U26503 ( .B(n18103), .A(n18104), .Z(n18055) );
  IV U26504 ( .A(n18105), .Z(n18103) );
  ANDN U26505 ( .B(n18106), .A(n18107), .Z(n18047) );
  XOR U26506 ( .A(n18033), .B(n18108), .Z(n18045) );
  XOR U26507 ( .A(n18034), .B(n18035), .Z(n18108) );
  XOR U26508 ( .A(n18040), .B(n18109), .Z(n18035) );
  XOR U26509 ( .A(n18039), .B(n18042), .Z(n18109) );
  IV U26510 ( .A(n18041), .Z(n18042) );
  NAND U26511 ( .A(n18110), .B(n18111), .Z(n18041) );
  OR U26512 ( .A(n18112), .B(n18113), .Z(n18111) );
  OR U26513 ( .A(n18114), .B(n18115), .Z(n18110) );
  NAND U26514 ( .A(n18116), .B(n18117), .Z(n18039) );
  OR U26515 ( .A(n18118), .B(n18119), .Z(n18117) );
  OR U26516 ( .A(n18120), .B(n18121), .Z(n18116) );
  NOR U26517 ( .A(n18122), .B(n18123), .Z(n18040) );
  ANDN U26518 ( .B(n18124), .A(n18125), .Z(n18034) );
  IV U26519 ( .A(n18126), .Z(n18124) );
  XNOR U26520 ( .A(n18027), .B(n18127), .Z(n18033) );
  XNOR U26521 ( .A(n18026), .B(n18028), .Z(n18127) );
  NAND U26522 ( .A(n18128), .B(n18129), .Z(n18028) );
  OR U26523 ( .A(n18130), .B(n18131), .Z(n18129) );
  OR U26524 ( .A(n18132), .B(n18133), .Z(n18128) );
  NAND U26525 ( .A(n18134), .B(n18135), .Z(n18026) );
  OR U26526 ( .A(n18136), .B(n18137), .Z(n18135) );
  OR U26527 ( .A(n18138), .B(n18139), .Z(n18134) );
  ANDN U26528 ( .B(n18140), .A(n18141), .Z(n18027) );
  IV U26529 ( .A(n18142), .Z(n18140) );
  XNOR U26530 ( .A(n18107), .B(n18106), .Z(N63790) );
  XOR U26531 ( .A(n18126), .B(n18125), .Z(n18106) );
  XNOR U26532 ( .A(n18141), .B(n18142), .Z(n18125) );
  XNOR U26533 ( .A(n18136), .B(n18137), .Z(n18142) );
  XNOR U26534 ( .A(n18138), .B(n18139), .Z(n18137) );
  XNOR U26535 ( .A(y[5917]), .B(x[5917]), .Z(n18139) );
  XNOR U26536 ( .A(y[5918]), .B(x[5918]), .Z(n18138) );
  XNOR U26537 ( .A(y[5916]), .B(x[5916]), .Z(n18136) );
  XNOR U26538 ( .A(n18130), .B(n18131), .Z(n18141) );
  XNOR U26539 ( .A(y[5913]), .B(x[5913]), .Z(n18131) );
  XNOR U26540 ( .A(n18132), .B(n18133), .Z(n18130) );
  XNOR U26541 ( .A(y[5914]), .B(x[5914]), .Z(n18133) );
  XNOR U26542 ( .A(y[5915]), .B(x[5915]), .Z(n18132) );
  XNOR U26543 ( .A(n18123), .B(n18122), .Z(n18126) );
  XNOR U26544 ( .A(n18118), .B(n18119), .Z(n18122) );
  XNOR U26545 ( .A(y[5910]), .B(x[5910]), .Z(n18119) );
  XNOR U26546 ( .A(n18120), .B(n18121), .Z(n18118) );
  XNOR U26547 ( .A(y[5911]), .B(x[5911]), .Z(n18121) );
  XNOR U26548 ( .A(y[5912]), .B(x[5912]), .Z(n18120) );
  XNOR U26549 ( .A(n18112), .B(n18113), .Z(n18123) );
  XNOR U26550 ( .A(y[5907]), .B(x[5907]), .Z(n18113) );
  XNOR U26551 ( .A(n18114), .B(n18115), .Z(n18112) );
  XNOR U26552 ( .A(y[5908]), .B(x[5908]), .Z(n18115) );
  XNOR U26553 ( .A(y[5909]), .B(x[5909]), .Z(n18114) );
  XOR U26554 ( .A(n18088), .B(n18089), .Z(n18107) );
  XNOR U26555 ( .A(n18104), .B(n18105), .Z(n18089) );
  XNOR U26556 ( .A(n18099), .B(n18100), .Z(n18105) );
  XNOR U26557 ( .A(n18101), .B(n18102), .Z(n18100) );
  XNOR U26558 ( .A(y[5905]), .B(x[5905]), .Z(n18102) );
  XNOR U26559 ( .A(y[5906]), .B(x[5906]), .Z(n18101) );
  XNOR U26560 ( .A(y[5904]), .B(x[5904]), .Z(n18099) );
  XNOR U26561 ( .A(n18093), .B(n18094), .Z(n18104) );
  XNOR U26562 ( .A(y[5901]), .B(x[5901]), .Z(n18094) );
  XNOR U26563 ( .A(n18095), .B(n18096), .Z(n18093) );
  XNOR U26564 ( .A(y[5902]), .B(x[5902]), .Z(n18096) );
  XNOR U26565 ( .A(y[5903]), .B(x[5903]), .Z(n18095) );
  XOR U26566 ( .A(n18087), .B(n18086), .Z(n18088) );
  XNOR U26567 ( .A(n18082), .B(n18083), .Z(n18086) );
  XNOR U26568 ( .A(y[5898]), .B(x[5898]), .Z(n18083) );
  XNOR U26569 ( .A(n18084), .B(n18085), .Z(n18082) );
  XNOR U26570 ( .A(y[5899]), .B(x[5899]), .Z(n18085) );
  XNOR U26571 ( .A(y[5900]), .B(x[5900]), .Z(n18084) );
  XNOR U26572 ( .A(n18076), .B(n18077), .Z(n18087) );
  XNOR U26573 ( .A(y[5895]), .B(x[5895]), .Z(n18077) );
  XNOR U26574 ( .A(n18078), .B(n18079), .Z(n18076) );
  XNOR U26575 ( .A(y[5896]), .B(x[5896]), .Z(n18079) );
  XNOR U26576 ( .A(y[5897]), .B(x[5897]), .Z(n18078) );
  NAND U26577 ( .A(n18143), .B(n18144), .Z(N63781) );
  NANDN U26578 ( .A(n18145), .B(n18146), .Z(n18144) );
  OR U26579 ( .A(n18147), .B(n18148), .Z(n18146) );
  NAND U26580 ( .A(n18147), .B(n18148), .Z(n18143) );
  XOR U26581 ( .A(n18147), .B(n18149), .Z(N63780) );
  XNOR U26582 ( .A(n18145), .B(n18148), .Z(n18149) );
  AND U26583 ( .A(n18150), .B(n18151), .Z(n18148) );
  NANDN U26584 ( .A(n18152), .B(n18153), .Z(n18151) );
  NANDN U26585 ( .A(n18154), .B(n18155), .Z(n18153) );
  NANDN U26586 ( .A(n18155), .B(n18154), .Z(n18150) );
  NAND U26587 ( .A(n18156), .B(n18157), .Z(n18145) );
  NANDN U26588 ( .A(n18158), .B(n18159), .Z(n18157) );
  OR U26589 ( .A(n18160), .B(n18161), .Z(n18159) );
  NAND U26590 ( .A(n18161), .B(n18160), .Z(n18156) );
  AND U26591 ( .A(n18162), .B(n18163), .Z(n18147) );
  NANDN U26592 ( .A(n18164), .B(n18165), .Z(n18163) );
  NANDN U26593 ( .A(n18166), .B(n18167), .Z(n18165) );
  NANDN U26594 ( .A(n18167), .B(n18166), .Z(n18162) );
  XOR U26595 ( .A(n18161), .B(n18168), .Z(N63779) );
  XOR U26596 ( .A(n18158), .B(n18160), .Z(n18168) );
  XNOR U26597 ( .A(n18154), .B(n18169), .Z(n18160) );
  XNOR U26598 ( .A(n18152), .B(n18155), .Z(n18169) );
  NAND U26599 ( .A(n18170), .B(n18171), .Z(n18155) );
  NAND U26600 ( .A(n18172), .B(n18173), .Z(n18171) );
  OR U26601 ( .A(n18174), .B(n18175), .Z(n18172) );
  NANDN U26602 ( .A(n18176), .B(n18174), .Z(n18170) );
  IV U26603 ( .A(n18175), .Z(n18176) );
  NAND U26604 ( .A(n18177), .B(n18178), .Z(n18152) );
  NAND U26605 ( .A(n18179), .B(n18180), .Z(n18178) );
  NANDN U26606 ( .A(n18181), .B(n18182), .Z(n18179) );
  NANDN U26607 ( .A(n18182), .B(n18181), .Z(n18177) );
  AND U26608 ( .A(n18183), .B(n18184), .Z(n18154) );
  NAND U26609 ( .A(n18185), .B(n18186), .Z(n18184) );
  OR U26610 ( .A(n18187), .B(n18188), .Z(n18185) );
  NANDN U26611 ( .A(n18189), .B(n18187), .Z(n18183) );
  NAND U26612 ( .A(n18190), .B(n18191), .Z(n18158) );
  NANDN U26613 ( .A(n18192), .B(n18193), .Z(n18191) );
  OR U26614 ( .A(n18194), .B(n18195), .Z(n18193) );
  NANDN U26615 ( .A(n18196), .B(n18194), .Z(n18190) );
  IV U26616 ( .A(n18195), .Z(n18196) );
  XNOR U26617 ( .A(n18166), .B(n18197), .Z(n18161) );
  XNOR U26618 ( .A(n18164), .B(n18167), .Z(n18197) );
  NAND U26619 ( .A(n18198), .B(n18199), .Z(n18167) );
  NAND U26620 ( .A(n18200), .B(n18201), .Z(n18199) );
  OR U26621 ( .A(n18202), .B(n18203), .Z(n18200) );
  NANDN U26622 ( .A(n18204), .B(n18202), .Z(n18198) );
  IV U26623 ( .A(n18203), .Z(n18204) );
  NAND U26624 ( .A(n18205), .B(n18206), .Z(n18164) );
  NAND U26625 ( .A(n18207), .B(n18208), .Z(n18206) );
  NANDN U26626 ( .A(n18209), .B(n18210), .Z(n18207) );
  NANDN U26627 ( .A(n18210), .B(n18209), .Z(n18205) );
  AND U26628 ( .A(n18211), .B(n18212), .Z(n18166) );
  NAND U26629 ( .A(n18213), .B(n18214), .Z(n18212) );
  OR U26630 ( .A(n18215), .B(n18216), .Z(n18213) );
  NANDN U26631 ( .A(n18217), .B(n18215), .Z(n18211) );
  XNOR U26632 ( .A(n18192), .B(n18218), .Z(N63778) );
  XOR U26633 ( .A(n18194), .B(n18195), .Z(n18218) );
  XNOR U26634 ( .A(n18208), .B(n18219), .Z(n18195) );
  XOR U26635 ( .A(n18209), .B(n18210), .Z(n18219) );
  XOR U26636 ( .A(n18215), .B(n18220), .Z(n18210) );
  XOR U26637 ( .A(n18214), .B(n18217), .Z(n18220) );
  IV U26638 ( .A(n18216), .Z(n18217) );
  NAND U26639 ( .A(n18221), .B(n18222), .Z(n18216) );
  OR U26640 ( .A(n18223), .B(n18224), .Z(n18222) );
  OR U26641 ( .A(n18225), .B(n18226), .Z(n18221) );
  NAND U26642 ( .A(n18227), .B(n18228), .Z(n18214) );
  OR U26643 ( .A(n18229), .B(n18230), .Z(n18228) );
  OR U26644 ( .A(n18231), .B(n18232), .Z(n18227) );
  NOR U26645 ( .A(n18233), .B(n18234), .Z(n18215) );
  ANDN U26646 ( .B(n18235), .A(n18236), .Z(n18209) );
  XNOR U26647 ( .A(n18202), .B(n18237), .Z(n18208) );
  XNOR U26648 ( .A(n18201), .B(n18203), .Z(n18237) );
  NAND U26649 ( .A(n18238), .B(n18239), .Z(n18203) );
  OR U26650 ( .A(n18240), .B(n18241), .Z(n18239) );
  OR U26651 ( .A(n18242), .B(n18243), .Z(n18238) );
  NAND U26652 ( .A(n18244), .B(n18245), .Z(n18201) );
  OR U26653 ( .A(n18246), .B(n18247), .Z(n18245) );
  OR U26654 ( .A(n18248), .B(n18249), .Z(n18244) );
  ANDN U26655 ( .B(n18250), .A(n18251), .Z(n18202) );
  IV U26656 ( .A(n18252), .Z(n18250) );
  ANDN U26657 ( .B(n18253), .A(n18254), .Z(n18194) );
  XOR U26658 ( .A(n18180), .B(n18255), .Z(n18192) );
  XOR U26659 ( .A(n18181), .B(n18182), .Z(n18255) );
  XOR U26660 ( .A(n18187), .B(n18256), .Z(n18182) );
  XOR U26661 ( .A(n18186), .B(n18189), .Z(n18256) );
  IV U26662 ( .A(n18188), .Z(n18189) );
  NAND U26663 ( .A(n18257), .B(n18258), .Z(n18188) );
  OR U26664 ( .A(n18259), .B(n18260), .Z(n18258) );
  OR U26665 ( .A(n18261), .B(n18262), .Z(n18257) );
  NAND U26666 ( .A(n18263), .B(n18264), .Z(n18186) );
  OR U26667 ( .A(n18265), .B(n18266), .Z(n18264) );
  OR U26668 ( .A(n18267), .B(n18268), .Z(n18263) );
  NOR U26669 ( .A(n18269), .B(n18270), .Z(n18187) );
  ANDN U26670 ( .B(n18271), .A(n18272), .Z(n18181) );
  IV U26671 ( .A(n18273), .Z(n18271) );
  XNOR U26672 ( .A(n18174), .B(n18274), .Z(n18180) );
  XNOR U26673 ( .A(n18173), .B(n18175), .Z(n18274) );
  NAND U26674 ( .A(n18275), .B(n18276), .Z(n18175) );
  OR U26675 ( .A(n18277), .B(n18278), .Z(n18276) );
  OR U26676 ( .A(n18279), .B(n18280), .Z(n18275) );
  NAND U26677 ( .A(n18281), .B(n18282), .Z(n18173) );
  OR U26678 ( .A(n18283), .B(n18284), .Z(n18282) );
  OR U26679 ( .A(n18285), .B(n18286), .Z(n18281) );
  ANDN U26680 ( .B(n18287), .A(n18288), .Z(n18174) );
  IV U26681 ( .A(n18289), .Z(n18287) );
  XNOR U26682 ( .A(n18254), .B(n18253), .Z(N63777) );
  XOR U26683 ( .A(n18273), .B(n18272), .Z(n18253) );
  XNOR U26684 ( .A(n18288), .B(n18289), .Z(n18272) );
  XNOR U26685 ( .A(n18283), .B(n18284), .Z(n18289) );
  XNOR U26686 ( .A(n18285), .B(n18286), .Z(n18284) );
  XNOR U26687 ( .A(y[5893]), .B(x[5893]), .Z(n18286) );
  XNOR U26688 ( .A(y[5894]), .B(x[5894]), .Z(n18285) );
  XNOR U26689 ( .A(y[5892]), .B(x[5892]), .Z(n18283) );
  XNOR U26690 ( .A(n18277), .B(n18278), .Z(n18288) );
  XNOR U26691 ( .A(y[5889]), .B(x[5889]), .Z(n18278) );
  XNOR U26692 ( .A(n18279), .B(n18280), .Z(n18277) );
  XNOR U26693 ( .A(y[5890]), .B(x[5890]), .Z(n18280) );
  XNOR U26694 ( .A(y[5891]), .B(x[5891]), .Z(n18279) );
  XNOR U26695 ( .A(n18270), .B(n18269), .Z(n18273) );
  XNOR U26696 ( .A(n18265), .B(n18266), .Z(n18269) );
  XNOR U26697 ( .A(y[5886]), .B(x[5886]), .Z(n18266) );
  XNOR U26698 ( .A(n18267), .B(n18268), .Z(n18265) );
  XNOR U26699 ( .A(y[5887]), .B(x[5887]), .Z(n18268) );
  XNOR U26700 ( .A(y[5888]), .B(x[5888]), .Z(n18267) );
  XNOR U26701 ( .A(n18259), .B(n18260), .Z(n18270) );
  XNOR U26702 ( .A(y[5883]), .B(x[5883]), .Z(n18260) );
  XNOR U26703 ( .A(n18261), .B(n18262), .Z(n18259) );
  XNOR U26704 ( .A(y[5884]), .B(x[5884]), .Z(n18262) );
  XNOR U26705 ( .A(y[5885]), .B(x[5885]), .Z(n18261) );
  XOR U26706 ( .A(n18235), .B(n18236), .Z(n18254) );
  XNOR U26707 ( .A(n18251), .B(n18252), .Z(n18236) );
  XNOR U26708 ( .A(n18246), .B(n18247), .Z(n18252) );
  XNOR U26709 ( .A(n18248), .B(n18249), .Z(n18247) );
  XNOR U26710 ( .A(y[5881]), .B(x[5881]), .Z(n18249) );
  XNOR U26711 ( .A(y[5882]), .B(x[5882]), .Z(n18248) );
  XNOR U26712 ( .A(y[5880]), .B(x[5880]), .Z(n18246) );
  XNOR U26713 ( .A(n18240), .B(n18241), .Z(n18251) );
  XNOR U26714 ( .A(y[5877]), .B(x[5877]), .Z(n18241) );
  XNOR U26715 ( .A(n18242), .B(n18243), .Z(n18240) );
  XNOR U26716 ( .A(y[5878]), .B(x[5878]), .Z(n18243) );
  XNOR U26717 ( .A(y[5879]), .B(x[5879]), .Z(n18242) );
  XOR U26718 ( .A(n18234), .B(n18233), .Z(n18235) );
  XNOR U26719 ( .A(n18229), .B(n18230), .Z(n18233) );
  XNOR U26720 ( .A(y[5874]), .B(x[5874]), .Z(n18230) );
  XNOR U26721 ( .A(n18231), .B(n18232), .Z(n18229) );
  XNOR U26722 ( .A(y[5875]), .B(x[5875]), .Z(n18232) );
  XNOR U26723 ( .A(y[5876]), .B(x[5876]), .Z(n18231) );
  XNOR U26724 ( .A(n18223), .B(n18224), .Z(n18234) );
  XNOR U26725 ( .A(y[5871]), .B(x[5871]), .Z(n18224) );
  XNOR U26726 ( .A(n18225), .B(n18226), .Z(n18223) );
  XNOR U26727 ( .A(y[5872]), .B(x[5872]), .Z(n18226) );
  XNOR U26728 ( .A(y[5873]), .B(x[5873]), .Z(n18225) );
  NAND U26729 ( .A(n18290), .B(n18291), .Z(N63768) );
  NANDN U26730 ( .A(n18292), .B(n18293), .Z(n18291) );
  OR U26731 ( .A(n18294), .B(n18295), .Z(n18293) );
  NAND U26732 ( .A(n18294), .B(n18295), .Z(n18290) );
  XOR U26733 ( .A(n18294), .B(n18296), .Z(N63767) );
  XNOR U26734 ( .A(n18292), .B(n18295), .Z(n18296) );
  AND U26735 ( .A(n18297), .B(n18298), .Z(n18295) );
  NANDN U26736 ( .A(n18299), .B(n18300), .Z(n18298) );
  NANDN U26737 ( .A(n18301), .B(n18302), .Z(n18300) );
  NANDN U26738 ( .A(n18302), .B(n18301), .Z(n18297) );
  NAND U26739 ( .A(n18303), .B(n18304), .Z(n18292) );
  NANDN U26740 ( .A(n18305), .B(n18306), .Z(n18304) );
  OR U26741 ( .A(n18307), .B(n18308), .Z(n18306) );
  NAND U26742 ( .A(n18308), .B(n18307), .Z(n18303) );
  AND U26743 ( .A(n18309), .B(n18310), .Z(n18294) );
  NANDN U26744 ( .A(n18311), .B(n18312), .Z(n18310) );
  NANDN U26745 ( .A(n18313), .B(n18314), .Z(n18312) );
  NANDN U26746 ( .A(n18314), .B(n18313), .Z(n18309) );
  XOR U26747 ( .A(n18308), .B(n18315), .Z(N63766) );
  XOR U26748 ( .A(n18305), .B(n18307), .Z(n18315) );
  XNOR U26749 ( .A(n18301), .B(n18316), .Z(n18307) );
  XNOR U26750 ( .A(n18299), .B(n18302), .Z(n18316) );
  NAND U26751 ( .A(n18317), .B(n18318), .Z(n18302) );
  NAND U26752 ( .A(n18319), .B(n18320), .Z(n18318) );
  OR U26753 ( .A(n18321), .B(n18322), .Z(n18319) );
  NANDN U26754 ( .A(n18323), .B(n18321), .Z(n18317) );
  IV U26755 ( .A(n18322), .Z(n18323) );
  NAND U26756 ( .A(n18324), .B(n18325), .Z(n18299) );
  NAND U26757 ( .A(n18326), .B(n18327), .Z(n18325) );
  NANDN U26758 ( .A(n18328), .B(n18329), .Z(n18326) );
  NANDN U26759 ( .A(n18329), .B(n18328), .Z(n18324) );
  AND U26760 ( .A(n18330), .B(n18331), .Z(n18301) );
  NAND U26761 ( .A(n18332), .B(n18333), .Z(n18331) );
  OR U26762 ( .A(n18334), .B(n18335), .Z(n18332) );
  NANDN U26763 ( .A(n18336), .B(n18334), .Z(n18330) );
  NAND U26764 ( .A(n18337), .B(n18338), .Z(n18305) );
  NANDN U26765 ( .A(n18339), .B(n18340), .Z(n18338) );
  OR U26766 ( .A(n18341), .B(n18342), .Z(n18340) );
  NANDN U26767 ( .A(n18343), .B(n18341), .Z(n18337) );
  IV U26768 ( .A(n18342), .Z(n18343) );
  XNOR U26769 ( .A(n18313), .B(n18344), .Z(n18308) );
  XNOR U26770 ( .A(n18311), .B(n18314), .Z(n18344) );
  NAND U26771 ( .A(n18345), .B(n18346), .Z(n18314) );
  NAND U26772 ( .A(n18347), .B(n18348), .Z(n18346) );
  OR U26773 ( .A(n18349), .B(n18350), .Z(n18347) );
  NANDN U26774 ( .A(n18351), .B(n18349), .Z(n18345) );
  IV U26775 ( .A(n18350), .Z(n18351) );
  NAND U26776 ( .A(n18352), .B(n18353), .Z(n18311) );
  NAND U26777 ( .A(n18354), .B(n18355), .Z(n18353) );
  NANDN U26778 ( .A(n18356), .B(n18357), .Z(n18354) );
  NANDN U26779 ( .A(n18357), .B(n18356), .Z(n18352) );
  AND U26780 ( .A(n18358), .B(n18359), .Z(n18313) );
  NAND U26781 ( .A(n18360), .B(n18361), .Z(n18359) );
  OR U26782 ( .A(n18362), .B(n18363), .Z(n18360) );
  NANDN U26783 ( .A(n18364), .B(n18362), .Z(n18358) );
  XNOR U26784 ( .A(n18339), .B(n18365), .Z(N63765) );
  XOR U26785 ( .A(n18341), .B(n18342), .Z(n18365) );
  XNOR U26786 ( .A(n18355), .B(n18366), .Z(n18342) );
  XOR U26787 ( .A(n18356), .B(n18357), .Z(n18366) );
  XOR U26788 ( .A(n18362), .B(n18367), .Z(n18357) );
  XOR U26789 ( .A(n18361), .B(n18364), .Z(n18367) );
  IV U26790 ( .A(n18363), .Z(n18364) );
  NAND U26791 ( .A(n18368), .B(n18369), .Z(n18363) );
  OR U26792 ( .A(n18370), .B(n18371), .Z(n18369) );
  OR U26793 ( .A(n18372), .B(n18373), .Z(n18368) );
  NAND U26794 ( .A(n18374), .B(n18375), .Z(n18361) );
  OR U26795 ( .A(n18376), .B(n18377), .Z(n18375) );
  OR U26796 ( .A(n18378), .B(n18379), .Z(n18374) );
  NOR U26797 ( .A(n18380), .B(n18381), .Z(n18362) );
  ANDN U26798 ( .B(n18382), .A(n18383), .Z(n18356) );
  XNOR U26799 ( .A(n18349), .B(n18384), .Z(n18355) );
  XNOR U26800 ( .A(n18348), .B(n18350), .Z(n18384) );
  NAND U26801 ( .A(n18385), .B(n18386), .Z(n18350) );
  OR U26802 ( .A(n18387), .B(n18388), .Z(n18386) );
  OR U26803 ( .A(n18389), .B(n18390), .Z(n18385) );
  NAND U26804 ( .A(n18391), .B(n18392), .Z(n18348) );
  OR U26805 ( .A(n18393), .B(n18394), .Z(n18392) );
  OR U26806 ( .A(n18395), .B(n18396), .Z(n18391) );
  ANDN U26807 ( .B(n18397), .A(n18398), .Z(n18349) );
  IV U26808 ( .A(n18399), .Z(n18397) );
  ANDN U26809 ( .B(n18400), .A(n18401), .Z(n18341) );
  XOR U26810 ( .A(n18327), .B(n18402), .Z(n18339) );
  XOR U26811 ( .A(n18328), .B(n18329), .Z(n18402) );
  XOR U26812 ( .A(n18334), .B(n18403), .Z(n18329) );
  XOR U26813 ( .A(n18333), .B(n18336), .Z(n18403) );
  IV U26814 ( .A(n18335), .Z(n18336) );
  NAND U26815 ( .A(n18404), .B(n18405), .Z(n18335) );
  OR U26816 ( .A(n18406), .B(n18407), .Z(n18405) );
  OR U26817 ( .A(n18408), .B(n18409), .Z(n18404) );
  NAND U26818 ( .A(n18410), .B(n18411), .Z(n18333) );
  OR U26819 ( .A(n18412), .B(n18413), .Z(n18411) );
  OR U26820 ( .A(n18414), .B(n18415), .Z(n18410) );
  NOR U26821 ( .A(n18416), .B(n18417), .Z(n18334) );
  ANDN U26822 ( .B(n18418), .A(n18419), .Z(n18328) );
  IV U26823 ( .A(n18420), .Z(n18418) );
  XNOR U26824 ( .A(n18321), .B(n18421), .Z(n18327) );
  XNOR U26825 ( .A(n18320), .B(n18322), .Z(n18421) );
  NAND U26826 ( .A(n18422), .B(n18423), .Z(n18322) );
  OR U26827 ( .A(n18424), .B(n18425), .Z(n18423) );
  OR U26828 ( .A(n18426), .B(n18427), .Z(n18422) );
  NAND U26829 ( .A(n18428), .B(n18429), .Z(n18320) );
  OR U26830 ( .A(n18430), .B(n18431), .Z(n18429) );
  OR U26831 ( .A(n18432), .B(n18433), .Z(n18428) );
  ANDN U26832 ( .B(n18434), .A(n18435), .Z(n18321) );
  IV U26833 ( .A(n18436), .Z(n18434) );
  XNOR U26834 ( .A(n18401), .B(n18400), .Z(N63764) );
  XOR U26835 ( .A(n18420), .B(n18419), .Z(n18400) );
  XNOR U26836 ( .A(n18435), .B(n18436), .Z(n18419) );
  XNOR U26837 ( .A(n18430), .B(n18431), .Z(n18436) );
  XNOR U26838 ( .A(n18432), .B(n18433), .Z(n18431) );
  XNOR U26839 ( .A(y[5869]), .B(x[5869]), .Z(n18433) );
  XNOR U26840 ( .A(y[5870]), .B(x[5870]), .Z(n18432) );
  XNOR U26841 ( .A(y[5868]), .B(x[5868]), .Z(n18430) );
  XNOR U26842 ( .A(n18424), .B(n18425), .Z(n18435) );
  XNOR U26843 ( .A(y[5865]), .B(x[5865]), .Z(n18425) );
  XNOR U26844 ( .A(n18426), .B(n18427), .Z(n18424) );
  XNOR U26845 ( .A(y[5866]), .B(x[5866]), .Z(n18427) );
  XNOR U26846 ( .A(y[5867]), .B(x[5867]), .Z(n18426) );
  XNOR U26847 ( .A(n18417), .B(n18416), .Z(n18420) );
  XNOR U26848 ( .A(n18412), .B(n18413), .Z(n18416) );
  XNOR U26849 ( .A(y[5862]), .B(x[5862]), .Z(n18413) );
  XNOR U26850 ( .A(n18414), .B(n18415), .Z(n18412) );
  XNOR U26851 ( .A(y[5863]), .B(x[5863]), .Z(n18415) );
  XNOR U26852 ( .A(y[5864]), .B(x[5864]), .Z(n18414) );
  XNOR U26853 ( .A(n18406), .B(n18407), .Z(n18417) );
  XNOR U26854 ( .A(y[5859]), .B(x[5859]), .Z(n18407) );
  XNOR U26855 ( .A(n18408), .B(n18409), .Z(n18406) );
  XNOR U26856 ( .A(y[5860]), .B(x[5860]), .Z(n18409) );
  XNOR U26857 ( .A(y[5861]), .B(x[5861]), .Z(n18408) );
  XOR U26858 ( .A(n18382), .B(n18383), .Z(n18401) );
  XNOR U26859 ( .A(n18398), .B(n18399), .Z(n18383) );
  XNOR U26860 ( .A(n18393), .B(n18394), .Z(n18399) );
  XNOR U26861 ( .A(n18395), .B(n18396), .Z(n18394) );
  XNOR U26862 ( .A(y[5857]), .B(x[5857]), .Z(n18396) );
  XNOR U26863 ( .A(y[5858]), .B(x[5858]), .Z(n18395) );
  XNOR U26864 ( .A(y[5856]), .B(x[5856]), .Z(n18393) );
  XNOR U26865 ( .A(n18387), .B(n18388), .Z(n18398) );
  XNOR U26866 ( .A(y[5853]), .B(x[5853]), .Z(n18388) );
  XNOR U26867 ( .A(n18389), .B(n18390), .Z(n18387) );
  XNOR U26868 ( .A(y[5854]), .B(x[5854]), .Z(n18390) );
  XNOR U26869 ( .A(y[5855]), .B(x[5855]), .Z(n18389) );
  XOR U26870 ( .A(n18381), .B(n18380), .Z(n18382) );
  XNOR U26871 ( .A(n18376), .B(n18377), .Z(n18380) );
  XNOR U26872 ( .A(y[5850]), .B(x[5850]), .Z(n18377) );
  XNOR U26873 ( .A(n18378), .B(n18379), .Z(n18376) );
  XNOR U26874 ( .A(y[5851]), .B(x[5851]), .Z(n18379) );
  XNOR U26875 ( .A(y[5852]), .B(x[5852]), .Z(n18378) );
  XNOR U26876 ( .A(n18370), .B(n18371), .Z(n18381) );
  XNOR U26877 ( .A(y[5847]), .B(x[5847]), .Z(n18371) );
  XNOR U26878 ( .A(n18372), .B(n18373), .Z(n18370) );
  XNOR U26879 ( .A(y[5848]), .B(x[5848]), .Z(n18373) );
  XNOR U26880 ( .A(y[5849]), .B(x[5849]), .Z(n18372) );
  NAND U26881 ( .A(n18437), .B(n18438), .Z(N63755) );
  NANDN U26882 ( .A(n18439), .B(n18440), .Z(n18438) );
  OR U26883 ( .A(n18441), .B(n18442), .Z(n18440) );
  NAND U26884 ( .A(n18441), .B(n18442), .Z(n18437) );
  XOR U26885 ( .A(n18441), .B(n18443), .Z(N63754) );
  XNOR U26886 ( .A(n18439), .B(n18442), .Z(n18443) );
  AND U26887 ( .A(n18444), .B(n18445), .Z(n18442) );
  NANDN U26888 ( .A(n18446), .B(n18447), .Z(n18445) );
  NANDN U26889 ( .A(n18448), .B(n18449), .Z(n18447) );
  NANDN U26890 ( .A(n18449), .B(n18448), .Z(n18444) );
  NAND U26891 ( .A(n18450), .B(n18451), .Z(n18439) );
  NANDN U26892 ( .A(n18452), .B(n18453), .Z(n18451) );
  OR U26893 ( .A(n18454), .B(n18455), .Z(n18453) );
  NAND U26894 ( .A(n18455), .B(n18454), .Z(n18450) );
  AND U26895 ( .A(n18456), .B(n18457), .Z(n18441) );
  NANDN U26896 ( .A(n18458), .B(n18459), .Z(n18457) );
  NANDN U26897 ( .A(n18460), .B(n18461), .Z(n18459) );
  NANDN U26898 ( .A(n18461), .B(n18460), .Z(n18456) );
  XOR U26899 ( .A(n18455), .B(n18462), .Z(N63753) );
  XOR U26900 ( .A(n18452), .B(n18454), .Z(n18462) );
  XNOR U26901 ( .A(n18448), .B(n18463), .Z(n18454) );
  XNOR U26902 ( .A(n18446), .B(n18449), .Z(n18463) );
  NAND U26903 ( .A(n18464), .B(n18465), .Z(n18449) );
  NAND U26904 ( .A(n18466), .B(n18467), .Z(n18465) );
  OR U26905 ( .A(n18468), .B(n18469), .Z(n18466) );
  NANDN U26906 ( .A(n18470), .B(n18468), .Z(n18464) );
  IV U26907 ( .A(n18469), .Z(n18470) );
  NAND U26908 ( .A(n18471), .B(n18472), .Z(n18446) );
  NAND U26909 ( .A(n18473), .B(n18474), .Z(n18472) );
  NANDN U26910 ( .A(n18475), .B(n18476), .Z(n18473) );
  NANDN U26911 ( .A(n18476), .B(n18475), .Z(n18471) );
  AND U26912 ( .A(n18477), .B(n18478), .Z(n18448) );
  NAND U26913 ( .A(n18479), .B(n18480), .Z(n18478) );
  OR U26914 ( .A(n18481), .B(n18482), .Z(n18479) );
  NANDN U26915 ( .A(n18483), .B(n18481), .Z(n18477) );
  NAND U26916 ( .A(n18484), .B(n18485), .Z(n18452) );
  NANDN U26917 ( .A(n18486), .B(n18487), .Z(n18485) );
  OR U26918 ( .A(n18488), .B(n18489), .Z(n18487) );
  NANDN U26919 ( .A(n18490), .B(n18488), .Z(n18484) );
  IV U26920 ( .A(n18489), .Z(n18490) );
  XNOR U26921 ( .A(n18460), .B(n18491), .Z(n18455) );
  XNOR U26922 ( .A(n18458), .B(n18461), .Z(n18491) );
  NAND U26923 ( .A(n18492), .B(n18493), .Z(n18461) );
  NAND U26924 ( .A(n18494), .B(n18495), .Z(n18493) );
  OR U26925 ( .A(n18496), .B(n18497), .Z(n18494) );
  NANDN U26926 ( .A(n18498), .B(n18496), .Z(n18492) );
  IV U26927 ( .A(n18497), .Z(n18498) );
  NAND U26928 ( .A(n18499), .B(n18500), .Z(n18458) );
  NAND U26929 ( .A(n18501), .B(n18502), .Z(n18500) );
  NANDN U26930 ( .A(n18503), .B(n18504), .Z(n18501) );
  NANDN U26931 ( .A(n18504), .B(n18503), .Z(n18499) );
  AND U26932 ( .A(n18505), .B(n18506), .Z(n18460) );
  NAND U26933 ( .A(n18507), .B(n18508), .Z(n18506) );
  OR U26934 ( .A(n18509), .B(n18510), .Z(n18507) );
  NANDN U26935 ( .A(n18511), .B(n18509), .Z(n18505) );
  XNOR U26936 ( .A(n18486), .B(n18512), .Z(N63752) );
  XOR U26937 ( .A(n18488), .B(n18489), .Z(n18512) );
  XNOR U26938 ( .A(n18502), .B(n18513), .Z(n18489) );
  XOR U26939 ( .A(n18503), .B(n18504), .Z(n18513) );
  XOR U26940 ( .A(n18509), .B(n18514), .Z(n18504) );
  XOR U26941 ( .A(n18508), .B(n18511), .Z(n18514) );
  IV U26942 ( .A(n18510), .Z(n18511) );
  NAND U26943 ( .A(n18515), .B(n18516), .Z(n18510) );
  OR U26944 ( .A(n18517), .B(n18518), .Z(n18516) );
  OR U26945 ( .A(n18519), .B(n18520), .Z(n18515) );
  NAND U26946 ( .A(n18521), .B(n18522), .Z(n18508) );
  OR U26947 ( .A(n18523), .B(n18524), .Z(n18522) );
  OR U26948 ( .A(n18525), .B(n18526), .Z(n18521) );
  NOR U26949 ( .A(n18527), .B(n18528), .Z(n18509) );
  ANDN U26950 ( .B(n18529), .A(n18530), .Z(n18503) );
  XNOR U26951 ( .A(n18496), .B(n18531), .Z(n18502) );
  XNOR U26952 ( .A(n18495), .B(n18497), .Z(n18531) );
  NAND U26953 ( .A(n18532), .B(n18533), .Z(n18497) );
  OR U26954 ( .A(n18534), .B(n18535), .Z(n18533) );
  OR U26955 ( .A(n18536), .B(n18537), .Z(n18532) );
  NAND U26956 ( .A(n18538), .B(n18539), .Z(n18495) );
  OR U26957 ( .A(n18540), .B(n18541), .Z(n18539) );
  OR U26958 ( .A(n18542), .B(n18543), .Z(n18538) );
  ANDN U26959 ( .B(n18544), .A(n18545), .Z(n18496) );
  IV U26960 ( .A(n18546), .Z(n18544) );
  ANDN U26961 ( .B(n18547), .A(n18548), .Z(n18488) );
  XOR U26962 ( .A(n18474), .B(n18549), .Z(n18486) );
  XOR U26963 ( .A(n18475), .B(n18476), .Z(n18549) );
  XOR U26964 ( .A(n18481), .B(n18550), .Z(n18476) );
  XOR U26965 ( .A(n18480), .B(n18483), .Z(n18550) );
  IV U26966 ( .A(n18482), .Z(n18483) );
  NAND U26967 ( .A(n18551), .B(n18552), .Z(n18482) );
  OR U26968 ( .A(n18553), .B(n18554), .Z(n18552) );
  OR U26969 ( .A(n18555), .B(n18556), .Z(n18551) );
  NAND U26970 ( .A(n18557), .B(n18558), .Z(n18480) );
  OR U26971 ( .A(n18559), .B(n18560), .Z(n18558) );
  OR U26972 ( .A(n18561), .B(n18562), .Z(n18557) );
  NOR U26973 ( .A(n18563), .B(n18564), .Z(n18481) );
  ANDN U26974 ( .B(n18565), .A(n18566), .Z(n18475) );
  IV U26975 ( .A(n18567), .Z(n18565) );
  XNOR U26976 ( .A(n18468), .B(n18568), .Z(n18474) );
  XNOR U26977 ( .A(n18467), .B(n18469), .Z(n18568) );
  NAND U26978 ( .A(n18569), .B(n18570), .Z(n18469) );
  OR U26979 ( .A(n18571), .B(n18572), .Z(n18570) );
  OR U26980 ( .A(n18573), .B(n18574), .Z(n18569) );
  NAND U26981 ( .A(n18575), .B(n18576), .Z(n18467) );
  OR U26982 ( .A(n18577), .B(n18578), .Z(n18576) );
  OR U26983 ( .A(n18579), .B(n18580), .Z(n18575) );
  ANDN U26984 ( .B(n18581), .A(n18582), .Z(n18468) );
  IV U26985 ( .A(n18583), .Z(n18581) );
  XNOR U26986 ( .A(n18548), .B(n18547), .Z(N63751) );
  XOR U26987 ( .A(n18567), .B(n18566), .Z(n18547) );
  XNOR U26988 ( .A(n18582), .B(n18583), .Z(n18566) );
  XNOR U26989 ( .A(n18577), .B(n18578), .Z(n18583) );
  XNOR U26990 ( .A(n18579), .B(n18580), .Z(n18578) );
  XNOR U26991 ( .A(y[5845]), .B(x[5845]), .Z(n18580) );
  XNOR U26992 ( .A(y[5846]), .B(x[5846]), .Z(n18579) );
  XNOR U26993 ( .A(y[5844]), .B(x[5844]), .Z(n18577) );
  XNOR U26994 ( .A(n18571), .B(n18572), .Z(n18582) );
  XNOR U26995 ( .A(y[5841]), .B(x[5841]), .Z(n18572) );
  XNOR U26996 ( .A(n18573), .B(n18574), .Z(n18571) );
  XNOR U26997 ( .A(y[5842]), .B(x[5842]), .Z(n18574) );
  XNOR U26998 ( .A(y[5843]), .B(x[5843]), .Z(n18573) );
  XNOR U26999 ( .A(n18564), .B(n18563), .Z(n18567) );
  XNOR U27000 ( .A(n18559), .B(n18560), .Z(n18563) );
  XNOR U27001 ( .A(y[5838]), .B(x[5838]), .Z(n18560) );
  XNOR U27002 ( .A(n18561), .B(n18562), .Z(n18559) );
  XNOR U27003 ( .A(y[5839]), .B(x[5839]), .Z(n18562) );
  XNOR U27004 ( .A(y[5840]), .B(x[5840]), .Z(n18561) );
  XNOR U27005 ( .A(n18553), .B(n18554), .Z(n18564) );
  XNOR U27006 ( .A(y[5835]), .B(x[5835]), .Z(n18554) );
  XNOR U27007 ( .A(n18555), .B(n18556), .Z(n18553) );
  XNOR U27008 ( .A(y[5836]), .B(x[5836]), .Z(n18556) );
  XNOR U27009 ( .A(y[5837]), .B(x[5837]), .Z(n18555) );
  XOR U27010 ( .A(n18529), .B(n18530), .Z(n18548) );
  XNOR U27011 ( .A(n18545), .B(n18546), .Z(n18530) );
  XNOR U27012 ( .A(n18540), .B(n18541), .Z(n18546) );
  XNOR U27013 ( .A(n18542), .B(n18543), .Z(n18541) );
  XNOR U27014 ( .A(y[5833]), .B(x[5833]), .Z(n18543) );
  XNOR U27015 ( .A(y[5834]), .B(x[5834]), .Z(n18542) );
  XNOR U27016 ( .A(y[5832]), .B(x[5832]), .Z(n18540) );
  XNOR U27017 ( .A(n18534), .B(n18535), .Z(n18545) );
  XNOR U27018 ( .A(y[5829]), .B(x[5829]), .Z(n18535) );
  XNOR U27019 ( .A(n18536), .B(n18537), .Z(n18534) );
  XNOR U27020 ( .A(y[5830]), .B(x[5830]), .Z(n18537) );
  XNOR U27021 ( .A(y[5831]), .B(x[5831]), .Z(n18536) );
  XOR U27022 ( .A(n18528), .B(n18527), .Z(n18529) );
  XNOR U27023 ( .A(n18523), .B(n18524), .Z(n18527) );
  XNOR U27024 ( .A(y[5826]), .B(x[5826]), .Z(n18524) );
  XNOR U27025 ( .A(n18525), .B(n18526), .Z(n18523) );
  XNOR U27026 ( .A(y[5827]), .B(x[5827]), .Z(n18526) );
  XNOR U27027 ( .A(y[5828]), .B(x[5828]), .Z(n18525) );
  XNOR U27028 ( .A(n18517), .B(n18518), .Z(n18528) );
  XNOR U27029 ( .A(y[5823]), .B(x[5823]), .Z(n18518) );
  XNOR U27030 ( .A(n18519), .B(n18520), .Z(n18517) );
  XNOR U27031 ( .A(y[5824]), .B(x[5824]), .Z(n18520) );
  XNOR U27032 ( .A(y[5825]), .B(x[5825]), .Z(n18519) );
  NAND U27033 ( .A(n18584), .B(n18585), .Z(N63742) );
  NANDN U27034 ( .A(n18586), .B(n18587), .Z(n18585) );
  OR U27035 ( .A(n18588), .B(n18589), .Z(n18587) );
  NAND U27036 ( .A(n18588), .B(n18589), .Z(n18584) );
  XOR U27037 ( .A(n18588), .B(n18590), .Z(N63741) );
  XNOR U27038 ( .A(n18586), .B(n18589), .Z(n18590) );
  AND U27039 ( .A(n18591), .B(n18592), .Z(n18589) );
  NANDN U27040 ( .A(n18593), .B(n18594), .Z(n18592) );
  NANDN U27041 ( .A(n18595), .B(n18596), .Z(n18594) );
  NANDN U27042 ( .A(n18596), .B(n18595), .Z(n18591) );
  NAND U27043 ( .A(n18597), .B(n18598), .Z(n18586) );
  NANDN U27044 ( .A(n18599), .B(n18600), .Z(n18598) );
  OR U27045 ( .A(n18601), .B(n18602), .Z(n18600) );
  NAND U27046 ( .A(n18602), .B(n18601), .Z(n18597) );
  AND U27047 ( .A(n18603), .B(n18604), .Z(n18588) );
  NANDN U27048 ( .A(n18605), .B(n18606), .Z(n18604) );
  NANDN U27049 ( .A(n18607), .B(n18608), .Z(n18606) );
  NANDN U27050 ( .A(n18608), .B(n18607), .Z(n18603) );
  XOR U27051 ( .A(n18602), .B(n18609), .Z(N63740) );
  XOR U27052 ( .A(n18599), .B(n18601), .Z(n18609) );
  XNOR U27053 ( .A(n18595), .B(n18610), .Z(n18601) );
  XNOR U27054 ( .A(n18593), .B(n18596), .Z(n18610) );
  NAND U27055 ( .A(n18611), .B(n18612), .Z(n18596) );
  NAND U27056 ( .A(n18613), .B(n18614), .Z(n18612) );
  OR U27057 ( .A(n18615), .B(n18616), .Z(n18613) );
  NANDN U27058 ( .A(n18617), .B(n18615), .Z(n18611) );
  IV U27059 ( .A(n18616), .Z(n18617) );
  NAND U27060 ( .A(n18618), .B(n18619), .Z(n18593) );
  NAND U27061 ( .A(n18620), .B(n18621), .Z(n18619) );
  NANDN U27062 ( .A(n18622), .B(n18623), .Z(n18620) );
  NANDN U27063 ( .A(n18623), .B(n18622), .Z(n18618) );
  AND U27064 ( .A(n18624), .B(n18625), .Z(n18595) );
  NAND U27065 ( .A(n18626), .B(n18627), .Z(n18625) );
  OR U27066 ( .A(n18628), .B(n18629), .Z(n18626) );
  NANDN U27067 ( .A(n18630), .B(n18628), .Z(n18624) );
  NAND U27068 ( .A(n18631), .B(n18632), .Z(n18599) );
  NANDN U27069 ( .A(n18633), .B(n18634), .Z(n18632) );
  OR U27070 ( .A(n18635), .B(n18636), .Z(n18634) );
  NANDN U27071 ( .A(n18637), .B(n18635), .Z(n18631) );
  IV U27072 ( .A(n18636), .Z(n18637) );
  XNOR U27073 ( .A(n18607), .B(n18638), .Z(n18602) );
  XNOR U27074 ( .A(n18605), .B(n18608), .Z(n18638) );
  NAND U27075 ( .A(n18639), .B(n18640), .Z(n18608) );
  NAND U27076 ( .A(n18641), .B(n18642), .Z(n18640) );
  OR U27077 ( .A(n18643), .B(n18644), .Z(n18641) );
  NANDN U27078 ( .A(n18645), .B(n18643), .Z(n18639) );
  IV U27079 ( .A(n18644), .Z(n18645) );
  NAND U27080 ( .A(n18646), .B(n18647), .Z(n18605) );
  NAND U27081 ( .A(n18648), .B(n18649), .Z(n18647) );
  NANDN U27082 ( .A(n18650), .B(n18651), .Z(n18648) );
  NANDN U27083 ( .A(n18651), .B(n18650), .Z(n18646) );
  AND U27084 ( .A(n18652), .B(n18653), .Z(n18607) );
  NAND U27085 ( .A(n18654), .B(n18655), .Z(n18653) );
  OR U27086 ( .A(n18656), .B(n18657), .Z(n18654) );
  NANDN U27087 ( .A(n18658), .B(n18656), .Z(n18652) );
  XNOR U27088 ( .A(n18633), .B(n18659), .Z(N63739) );
  XOR U27089 ( .A(n18635), .B(n18636), .Z(n18659) );
  XNOR U27090 ( .A(n18649), .B(n18660), .Z(n18636) );
  XOR U27091 ( .A(n18650), .B(n18651), .Z(n18660) );
  XOR U27092 ( .A(n18656), .B(n18661), .Z(n18651) );
  XOR U27093 ( .A(n18655), .B(n18658), .Z(n18661) );
  IV U27094 ( .A(n18657), .Z(n18658) );
  NAND U27095 ( .A(n18662), .B(n18663), .Z(n18657) );
  OR U27096 ( .A(n18664), .B(n18665), .Z(n18663) );
  OR U27097 ( .A(n18666), .B(n18667), .Z(n18662) );
  NAND U27098 ( .A(n18668), .B(n18669), .Z(n18655) );
  OR U27099 ( .A(n18670), .B(n18671), .Z(n18669) );
  OR U27100 ( .A(n18672), .B(n18673), .Z(n18668) );
  NOR U27101 ( .A(n18674), .B(n18675), .Z(n18656) );
  ANDN U27102 ( .B(n18676), .A(n18677), .Z(n18650) );
  XNOR U27103 ( .A(n18643), .B(n18678), .Z(n18649) );
  XNOR U27104 ( .A(n18642), .B(n18644), .Z(n18678) );
  NAND U27105 ( .A(n18679), .B(n18680), .Z(n18644) );
  OR U27106 ( .A(n18681), .B(n18682), .Z(n18680) );
  OR U27107 ( .A(n18683), .B(n18684), .Z(n18679) );
  NAND U27108 ( .A(n18685), .B(n18686), .Z(n18642) );
  OR U27109 ( .A(n18687), .B(n18688), .Z(n18686) );
  OR U27110 ( .A(n18689), .B(n18690), .Z(n18685) );
  ANDN U27111 ( .B(n18691), .A(n18692), .Z(n18643) );
  IV U27112 ( .A(n18693), .Z(n18691) );
  ANDN U27113 ( .B(n18694), .A(n18695), .Z(n18635) );
  XOR U27114 ( .A(n18621), .B(n18696), .Z(n18633) );
  XOR U27115 ( .A(n18622), .B(n18623), .Z(n18696) );
  XOR U27116 ( .A(n18628), .B(n18697), .Z(n18623) );
  XOR U27117 ( .A(n18627), .B(n18630), .Z(n18697) );
  IV U27118 ( .A(n18629), .Z(n18630) );
  NAND U27119 ( .A(n18698), .B(n18699), .Z(n18629) );
  OR U27120 ( .A(n18700), .B(n18701), .Z(n18699) );
  OR U27121 ( .A(n18702), .B(n18703), .Z(n18698) );
  NAND U27122 ( .A(n18704), .B(n18705), .Z(n18627) );
  OR U27123 ( .A(n18706), .B(n18707), .Z(n18705) );
  OR U27124 ( .A(n18708), .B(n18709), .Z(n18704) );
  NOR U27125 ( .A(n18710), .B(n18711), .Z(n18628) );
  ANDN U27126 ( .B(n18712), .A(n18713), .Z(n18622) );
  IV U27127 ( .A(n18714), .Z(n18712) );
  XNOR U27128 ( .A(n18615), .B(n18715), .Z(n18621) );
  XNOR U27129 ( .A(n18614), .B(n18616), .Z(n18715) );
  NAND U27130 ( .A(n18716), .B(n18717), .Z(n18616) );
  OR U27131 ( .A(n18718), .B(n18719), .Z(n18717) );
  OR U27132 ( .A(n18720), .B(n18721), .Z(n18716) );
  NAND U27133 ( .A(n18722), .B(n18723), .Z(n18614) );
  OR U27134 ( .A(n18724), .B(n18725), .Z(n18723) );
  OR U27135 ( .A(n18726), .B(n18727), .Z(n18722) );
  ANDN U27136 ( .B(n18728), .A(n18729), .Z(n18615) );
  IV U27137 ( .A(n18730), .Z(n18728) );
  XNOR U27138 ( .A(n18695), .B(n18694), .Z(N63738) );
  XOR U27139 ( .A(n18714), .B(n18713), .Z(n18694) );
  XNOR U27140 ( .A(n18729), .B(n18730), .Z(n18713) );
  XNOR U27141 ( .A(n18724), .B(n18725), .Z(n18730) );
  XNOR U27142 ( .A(n18726), .B(n18727), .Z(n18725) );
  XNOR U27143 ( .A(y[5821]), .B(x[5821]), .Z(n18727) );
  XNOR U27144 ( .A(y[5822]), .B(x[5822]), .Z(n18726) );
  XNOR U27145 ( .A(y[5820]), .B(x[5820]), .Z(n18724) );
  XNOR U27146 ( .A(n18718), .B(n18719), .Z(n18729) );
  XNOR U27147 ( .A(y[5817]), .B(x[5817]), .Z(n18719) );
  XNOR U27148 ( .A(n18720), .B(n18721), .Z(n18718) );
  XNOR U27149 ( .A(y[5818]), .B(x[5818]), .Z(n18721) );
  XNOR U27150 ( .A(y[5819]), .B(x[5819]), .Z(n18720) );
  XNOR U27151 ( .A(n18711), .B(n18710), .Z(n18714) );
  XNOR U27152 ( .A(n18706), .B(n18707), .Z(n18710) );
  XNOR U27153 ( .A(y[5814]), .B(x[5814]), .Z(n18707) );
  XNOR U27154 ( .A(n18708), .B(n18709), .Z(n18706) );
  XNOR U27155 ( .A(y[5815]), .B(x[5815]), .Z(n18709) );
  XNOR U27156 ( .A(y[5816]), .B(x[5816]), .Z(n18708) );
  XNOR U27157 ( .A(n18700), .B(n18701), .Z(n18711) );
  XNOR U27158 ( .A(y[5811]), .B(x[5811]), .Z(n18701) );
  XNOR U27159 ( .A(n18702), .B(n18703), .Z(n18700) );
  XNOR U27160 ( .A(y[5812]), .B(x[5812]), .Z(n18703) );
  XNOR U27161 ( .A(y[5813]), .B(x[5813]), .Z(n18702) );
  XOR U27162 ( .A(n18676), .B(n18677), .Z(n18695) );
  XNOR U27163 ( .A(n18692), .B(n18693), .Z(n18677) );
  XNOR U27164 ( .A(n18687), .B(n18688), .Z(n18693) );
  XNOR U27165 ( .A(n18689), .B(n18690), .Z(n18688) );
  XNOR U27166 ( .A(y[5809]), .B(x[5809]), .Z(n18690) );
  XNOR U27167 ( .A(y[5810]), .B(x[5810]), .Z(n18689) );
  XNOR U27168 ( .A(y[5808]), .B(x[5808]), .Z(n18687) );
  XNOR U27169 ( .A(n18681), .B(n18682), .Z(n18692) );
  XNOR U27170 ( .A(y[5805]), .B(x[5805]), .Z(n18682) );
  XNOR U27171 ( .A(n18683), .B(n18684), .Z(n18681) );
  XNOR U27172 ( .A(y[5806]), .B(x[5806]), .Z(n18684) );
  XNOR U27173 ( .A(y[5807]), .B(x[5807]), .Z(n18683) );
  XOR U27174 ( .A(n18675), .B(n18674), .Z(n18676) );
  XNOR U27175 ( .A(n18670), .B(n18671), .Z(n18674) );
  XNOR U27176 ( .A(y[5802]), .B(x[5802]), .Z(n18671) );
  XNOR U27177 ( .A(n18672), .B(n18673), .Z(n18670) );
  XNOR U27178 ( .A(y[5803]), .B(x[5803]), .Z(n18673) );
  XNOR U27179 ( .A(y[5804]), .B(x[5804]), .Z(n18672) );
  XNOR U27180 ( .A(n18664), .B(n18665), .Z(n18675) );
  XNOR U27181 ( .A(y[5799]), .B(x[5799]), .Z(n18665) );
  XNOR U27182 ( .A(n18666), .B(n18667), .Z(n18664) );
  XNOR U27183 ( .A(y[5800]), .B(x[5800]), .Z(n18667) );
  XNOR U27184 ( .A(y[5801]), .B(x[5801]), .Z(n18666) );
  NAND U27185 ( .A(n18731), .B(n18732), .Z(N63729) );
  NANDN U27186 ( .A(n18733), .B(n18734), .Z(n18732) );
  OR U27187 ( .A(n18735), .B(n18736), .Z(n18734) );
  NAND U27188 ( .A(n18735), .B(n18736), .Z(n18731) );
  XOR U27189 ( .A(n18735), .B(n18737), .Z(N63728) );
  XNOR U27190 ( .A(n18733), .B(n18736), .Z(n18737) );
  AND U27191 ( .A(n18738), .B(n18739), .Z(n18736) );
  NANDN U27192 ( .A(n18740), .B(n18741), .Z(n18739) );
  NANDN U27193 ( .A(n18742), .B(n18743), .Z(n18741) );
  NANDN U27194 ( .A(n18743), .B(n18742), .Z(n18738) );
  NAND U27195 ( .A(n18744), .B(n18745), .Z(n18733) );
  NANDN U27196 ( .A(n18746), .B(n18747), .Z(n18745) );
  OR U27197 ( .A(n18748), .B(n18749), .Z(n18747) );
  NAND U27198 ( .A(n18749), .B(n18748), .Z(n18744) );
  AND U27199 ( .A(n18750), .B(n18751), .Z(n18735) );
  NANDN U27200 ( .A(n18752), .B(n18753), .Z(n18751) );
  NANDN U27201 ( .A(n18754), .B(n18755), .Z(n18753) );
  NANDN U27202 ( .A(n18755), .B(n18754), .Z(n18750) );
  XOR U27203 ( .A(n18749), .B(n18756), .Z(N63727) );
  XOR U27204 ( .A(n18746), .B(n18748), .Z(n18756) );
  XNOR U27205 ( .A(n18742), .B(n18757), .Z(n18748) );
  XNOR U27206 ( .A(n18740), .B(n18743), .Z(n18757) );
  NAND U27207 ( .A(n18758), .B(n18759), .Z(n18743) );
  NAND U27208 ( .A(n18760), .B(n18761), .Z(n18759) );
  OR U27209 ( .A(n18762), .B(n18763), .Z(n18760) );
  NANDN U27210 ( .A(n18764), .B(n18762), .Z(n18758) );
  IV U27211 ( .A(n18763), .Z(n18764) );
  NAND U27212 ( .A(n18765), .B(n18766), .Z(n18740) );
  NAND U27213 ( .A(n18767), .B(n18768), .Z(n18766) );
  NANDN U27214 ( .A(n18769), .B(n18770), .Z(n18767) );
  NANDN U27215 ( .A(n18770), .B(n18769), .Z(n18765) );
  AND U27216 ( .A(n18771), .B(n18772), .Z(n18742) );
  NAND U27217 ( .A(n18773), .B(n18774), .Z(n18772) );
  OR U27218 ( .A(n18775), .B(n18776), .Z(n18773) );
  NANDN U27219 ( .A(n18777), .B(n18775), .Z(n18771) );
  NAND U27220 ( .A(n18778), .B(n18779), .Z(n18746) );
  NANDN U27221 ( .A(n18780), .B(n18781), .Z(n18779) );
  OR U27222 ( .A(n18782), .B(n18783), .Z(n18781) );
  NANDN U27223 ( .A(n18784), .B(n18782), .Z(n18778) );
  IV U27224 ( .A(n18783), .Z(n18784) );
  XNOR U27225 ( .A(n18754), .B(n18785), .Z(n18749) );
  XNOR U27226 ( .A(n18752), .B(n18755), .Z(n18785) );
  NAND U27227 ( .A(n18786), .B(n18787), .Z(n18755) );
  NAND U27228 ( .A(n18788), .B(n18789), .Z(n18787) );
  OR U27229 ( .A(n18790), .B(n18791), .Z(n18788) );
  NANDN U27230 ( .A(n18792), .B(n18790), .Z(n18786) );
  IV U27231 ( .A(n18791), .Z(n18792) );
  NAND U27232 ( .A(n18793), .B(n18794), .Z(n18752) );
  NAND U27233 ( .A(n18795), .B(n18796), .Z(n18794) );
  NANDN U27234 ( .A(n18797), .B(n18798), .Z(n18795) );
  NANDN U27235 ( .A(n18798), .B(n18797), .Z(n18793) );
  AND U27236 ( .A(n18799), .B(n18800), .Z(n18754) );
  NAND U27237 ( .A(n18801), .B(n18802), .Z(n18800) );
  OR U27238 ( .A(n18803), .B(n18804), .Z(n18801) );
  NANDN U27239 ( .A(n18805), .B(n18803), .Z(n18799) );
  XNOR U27240 ( .A(n18780), .B(n18806), .Z(N63726) );
  XOR U27241 ( .A(n18782), .B(n18783), .Z(n18806) );
  XNOR U27242 ( .A(n18796), .B(n18807), .Z(n18783) );
  XOR U27243 ( .A(n18797), .B(n18798), .Z(n18807) );
  XOR U27244 ( .A(n18803), .B(n18808), .Z(n18798) );
  XOR U27245 ( .A(n18802), .B(n18805), .Z(n18808) );
  IV U27246 ( .A(n18804), .Z(n18805) );
  NAND U27247 ( .A(n18809), .B(n18810), .Z(n18804) );
  OR U27248 ( .A(n18811), .B(n18812), .Z(n18810) );
  OR U27249 ( .A(n18813), .B(n18814), .Z(n18809) );
  NAND U27250 ( .A(n18815), .B(n18816), .Z(n18802) );
  OR U27251 ( .A(n18817), .B(n18818), .Z(n18816) );
  OR U27252 ( .A(n18819), .B(n18820), .Z(n18815) );
  NOR U27253 ( .A(n18821), .B(n18822), .Z(n18803) );
  ANDN U27254 ( .B(n18823), .A(n18824), .Z(n18797) );
  XNOR U27255 ( .A(n18790), .B(n18825), .Z(n18796) );
  XNOR U27256 ( .A(n18789), .B(n18791), .Z(n18825) );
  NAND U27257 ( .A(n18826), .B(n18827), .Z(n18791) );
  OR U27258 ( .A(n18828), .B(n18829), .Z(n18827) );
  OR U27259 ( .A(n18830), .B(n18831), .Z(n18826) );
  NAND U27260 ( .A(n18832), .B(n18833), .Z(n18789) );
  OR U27261 ( .A(n18834), .B(n18835), .Z(n18833) );
  OR U27262 ( .A(n18836), .B(n18837), .Z(n18832) );
  ANDN U27263 ( .B(n18838), .A(n18839), .Z(n18790) );
  IV U27264 ( .A(n18840), .Z(n18838) );
  ANDN U27265 ( .B(n18841), .A(n18842), .Z(n18782) );
  XOR U27266 ( .A(n18768), .B(n18843), .Z(n18780) );
  XOR U27267 ( .A(n18769), .B(n18770), .Z(n18843) );
  XOR U27268 ( .A(n18775), .B(n18844), .Z(n18770) );
  XOR U27269 ( .A(n18774), .B(n18777), .Z(n18844) );
  IV U27270 ( .A(n18776), .Z(n18777) );
  NAND U27271 ( .A(n18845), .B(n18846), .Z(n18776) );
  OR U27272 ( .A(n18847), .B(n18848), .Z(n18846) );
  OR U27273 ( .A(n18849), .B(n18850), .Z(n18845) );
  NAND U27274 ( .A(n18851), .B(n18852), .Z(n18774) );
  OR U27275 ( .A(n18853), .B(n18854), .Z(n18852) );
  OR U27276 ( .A(n18855), .B(n18856), .Z(n18851) );
  NOR U27277 ( .A(n18857), .B(n18858), .Z(n18775) );
  ANDN U27278 ( .B(n18859), .A(n18860), .Z(n18769) );
  IV U27279 ( .A(n18861), .Z(n18859) );
  XNOR U27280 ( .A(n18762), .B(n18862), .Z(n18768) );
  XNOR U27281 ( .A(n18761), .B(n18763), .Z(n18862) );
  NAND U27282 ( .A(n18863), .B(n18864), .Z(n18763) );
  OR U27283 ( .A(n18865), .B(n18866), .Z(n18864) );
  OR U27284 ( .A(n18867), .B(n18868), .Z(n18863) );
  NAND U27285 ( .A(n18869), .B(n18870), .Z(n18761) );
  OR U27286 ( .A(n18871), .B(n18872), .Z(n18870) );
  OR U27287 ( .A(n18873), .B(n18874), .Z(n18869) );
  ANDN U27288 ( .B(n18875), .A(n18876), .Z(n18762) );
  IV U27289 ( .A(n18877), .Z(n18875) );
  XNOR U27290 ( .A(n18842), .B(n18841), .Z(N63725) );
  XOR U27291 ( .A(n18861), .B(n18860), .Z(n18841) );
  XNOR U27292 ( .A(n18876), .B(n18877), .Z(n18860) );
  XNOR U27293 ( .A(n18871), .B(n18872), .Z(n18877) );
  XNOR U27294 ( .A(n18873), .B(n18874), .Z(n18872) );
  XNOR U27295 ( .A(y[5797]), .B(x[5797]), .Z(n18874) );
  XNOR U27296 ( .A(y[5798]), .B(x[5798]), .Z(n18873) );
  XNOR U27297 ( .A(y[5796]), .B(x[5796]), .Z(n18871) );
  XNOR U27298 ( .A(n18865), .B(n18866), .Z(n18876) );
  XNOR U27299 ( .A(y[5793]), .B(x[5793]), .Z(n18866) );
  XNOR U27300 ( .A(n18867), .B(n18868), .Z(n18865) );
  XNOR U27301 ( .A(y[5794]), .B(x[5794]), .Z(n18868) );
  XNOR U27302 ( .A(y[5795]), .B(x[5795]), .Z(n18867) );
  XNOR U27303 ( .A(n18858), .B(n18857), .Z(n18861) );
  XNOR U27304 ( .A(n18853), .B(n18854), .Z(n18857) );
  XNOR U27305 ( .A(y[5790]), .B(x[5790]), .Z(n18854) );
  XNOR U27306 ( .A(n18855), .B(n18856), .Z(n18853) );
  XNOR U27307 ( .A(y[5791]), .B(x[5791]), .Z(n18856) );
  XNOR U27308 ( .A(y[5792]), .B(x[5792]), .Z(n18855) );
  XNOR U27309 ( .A(n18847), .B(n18848), .Z(n18858) );
  XNOR U27310 ( .A(y[5787]), .B(x[5787]), .Z(n18848) );
  XNOR U27311 ( .A(n18849), .B(n18850), .Z(n18847) );
  XNOR U27312 ( .A(y[5788]), .B(x[5788]), .Z(n18850) );
  XNOR U27313 ( .A(y[5789]), .B(x[5789]), .Z(n18849) );
  XOR U27314 ( .A(n18823), .B(n18824), .Z(n18842) );
  XNOR U27315 ( .A(n18839), .B(n18840), .Z(n18824) );
  XNOR U27316 ( .A(n18834), .B(n18835), .Z(n18840) );
  XNOR U27317 ( .A(n18836), .B(n18837), .Z(n18835) );
  XNOR U27318 ( .A(y[5785]), .B(x[5785]), .Z(n18837) );
  XNOR U27319 ( .A(y[5786]), .B(x[5786]), .Z(n18836) );
  XNOR U27320 ( .A(y[5784]), .B(x[5784]), .Z(n18834) );
  XNOR U27321 ( .A(n18828), .B(n18829), .Z(n18839) );
  XNOR U27322 ( .A(y[5781]), .B(x[5781]), .Z(n18829) );
  XNOR U27323 ( .A(n18830), .B(n18831), .Z(n18828) );
  XNOR U27324 ( .A(y[5782]), .B(x[5782]), .Z(n18831) );
  XNOR U27325 ( .A(y[5783]), .B(x[5783]), .Z(n18830) );
  XOR U27326 ( .A(n18822), .B(n18821), .Z(n18823) );
  XNOR U27327 ( .A(n18817), .B(n18818), .Z(n18821) );
  XNOR U27328 ( .A(y[5778]), .B(x[5778]), .Z(n18818) );
  XNOR U27329 ( .A(n18819), .B(n18820), .Z(n18817) );
  XNOR U27330 ( .A(y[5779]), .B(x[5779]), .Z(n18820) );
  XNOR U27331 ( .A(y[5780]), .B(x[5780]), .Z(n18819) );
  XNOR U27332 ( .A(n18811), .B(n18812), .Z(n18822) );
  XNOR U27333 ( .A(y[5775]), .B(x[5775]), .Z(n18812) );
  XNOR U27334 ( .A(n18813), .B(n18814), .Z(n18811) );
  XNOR U27335 ( .A(y[5776]), .B(x[5776]), .Z(n18814) );
  XNOR U27336 ( .A(y[5777]), .B(x[5777]), .Z(n18813) );
  NAND U27337 ( .A(n18878), .B(n18879), .Z(N63716) );
  NANDN U27338 ( .A(n18880), .B(n18881), .Z(n18879) );
  OR U27339 ( .A(n18882), .B(n18883), .Z(n18881) );
  NAND U27340 ( .A(n18882), .B(n18883), .Z(n18878) );
  XOR U27341 ( .A(n18882), .B(n18884), .Z(N63715) );
  XNOR U27342 ( .A(n18880), .B(n18883), .Z(n18884) );
  AND U27343 ( .A(n18885), .B(n18886), .Z(n18883) );
  NANDN U27344 ( .A(n18887), .B(n18888), .Z(n18886) );
  NANDN U27345 ( .A(n18889), .B(n18890), .Z(n18888) );
  NANDN U27346 ( .A(n18890), .B(n18889), .Z(n18885) );
  NAND U27347 ( .A(n18891), .B(n18892), .Z(n18880) );
  NANDN U27348 ( .A(n18893), .B(n18894), .Z(n18892) );
  OR U27349 ( .A(n18895), .B(n18896), .Z(n18894) );
  NAND U27350 ( .A(n18896), .B(n18895), .Z(n18891) );
  AND U27351 ( .A(n18897), .B(n18898), .Z(n18882) );
  NANDN U27352 ( .A(n18899), .B(n18900), .Z(n18898) );
  NANDN U27353 ( .A(n18901), .B(n18902), .Z(n18900) );
  NANDN U27354 ( .A(n18902), .B(n18901), .Z(n18897) );
  XOR U27355 ( .A(n18896), .B(n18903), .Z(N63714) );
  XOR U27356 ( .A(n18893), .B(n18895), .Z(n18903) );
  XNOR U27357 ( .A(n18889), .B(n18904), .Z(n18895) );
  XNOR U27358 ( .A(n18887), .B(n18890), .Z(n18904) );
  NAND U27359 ( .A(n18905), .B(n18906), .Z(n18890) );
  NAND U27360 ( .A(n18907), .B(n18908), .Z(n18906) );
  OR U27361 ( .A(n18909), .B(n18910), .Z(n18907) );
  NANDN U27362 ( .A(n18911), .B(n18909), .Z(n18905) );
  IV U27363 ( .A(n18910), .Z(n18911) );
  NAND U27364 ( .A(n18912), .B(n18913), .Z(n18887) );
  NAND U27365 ( .A(n18914), .B(n18915), .Z(n18913) );
  NANDN U27366 ( .A(n18916), .B(n18917), .Z(n18914) );
  NANDN U27367 ( .A(n18917), .B(n18916), .Z(n18912) );
  AND U27368 ( .A(n18918), .B(n18919), .Z(n18889) );
  NAND U27369 ( .A(n18920), .B(n18921), .Z(n18919) );
  OR U27370 ( .A(n18922), .B(n18923), .Z(n18920) );
  NANDN U27371 ( .A(n18924), .B(n18922), .Z(n18918) );
  NAND U27372 ( .A(n18925), .B(n18926), .Z(n18893) );
  NANDN U27373 ( .A(n18927), .B(n18928), .Z(n18926) );
  OR U27374 ( .A(n18929), .B(n18930), .Z(n18928) );
  NANDN U27375 ( .A(n18931), .B(n18929), .Z(n18925) );
  IV U27376 ( .A(n18930), .Z(n18931) );
  XNOR U27377 ( .A(n18901), .B(n18932), .Z(n18896) );
  XNOR U27378 ( .A(n18899), .B(n18902), .Z(n18932) );
  NAND U27379 ( .A(n18933), .B(n18934), .Z(n18902) );
  NAND U27380 ( .A(n18935), .B(n18936), .Z(n18934) );
  OR U27381 ( .A(n18937), .B(n18938), .Z(n18935) );
  NANDN U27382 ( .A(n18939), .B(n18937), .Z(n18933) );
  IV U27383 ( .A(n18938), .Z(n18939) );
  NAND U27384 ( .A(n18940), .B(n18941), .Z(n18899) );
  NAND U27385 ( .A(n18942), .B(n18943), .Z(n18941) );
  NANDN U27386 ( .A(n18944), .B(n18945), .Z(n18942) );
  NANDN U27387 ( .A(n18945), .B(n18944), .Z(n18940) );
  AND U27388 ( .A(n18946), .B(n18947), .Z(n18901) );
  NAND U27389 ( .A(n18948), .B(n18949), .Z(n18947) );
  OR U27390 ( .A(n18950), .B(n18951), .Z(n18948) );
  NANDN U27391 ( .A(n18952), .B(n18950), .Z(n18946) );
  XNOR U27392 ( .A(n18927), .B(n18953), .Z(N63713) );
  XOR U27393 ( .A(n18929), .B(n18930), .Z(n18953) );
  XNOR U27394 ( .A(n18943), .B(n18954), .Z(n18930) );
  XOR U27395 ( .A(n18944), .B(n18945), .Z(n18954) );
  XOR U27396 ( .A(n18950), .B(n18955), .Z(n18945) );
  XOR U27397 ( .A(n18949), .B(n18952), .Z(n18955) );
  IV U27398 ( .A(n18951), .Z(n18952) );
  NAND U27399 ( .A(n18956), .B(n18957), .Z(n18951) );
  OR U27400 ( .A(n18958), .B(n18959), .Z(n18957) );
  OR U27401 ( .A(n18960), .B(n18961), .Z(n18956) );
  NAND U27402 ( .A(n18962), .B(n18963), .Z(n18949) );
  OR U27403 ( .A(n18964), .B(n18965), .Z(n18963) );
  OR U27404 ( .A(n18966), .B(n18967), .Z(n18962) );
  NOR U27405 ( .A(n18968), .B(n18969), .Z(n18950) );
  ANDN U27406 ( .B(n18970), .A(n18971), .Z(n18944) );
  XNOR U27407 ( .A(n18937), .B(n18972), .Z(n18943) );
  XNOR U27408 ( .A(n18936), .B(n18938), .Z(n18972) );
  NAND U27409 ( .A(n18973), .B(n18974), .Z(n18938) );
  OR U27410 ( .A(n18975), .B(n18976), .Z(n18974) );
  OR U27411 ( .A(n18977), .B(n18978), .Z(n18973) );
  NAND U27412 ( .A(n18979), .B(n18980), .Z(n18936) );
  OR U27413 ( .A(n18981), .B(n18982), .Z(n18980) );
  OR U27414 ( .A(n18983), .B(n18984), .Z(n18979) );
  ANDN U27415 ( .B(n18985), .A(n18986), .Z(n18937) );
  IV U27416 ( .A(n18987), .Z(n18985) );
  ANDN U27417 ( .B(n18988), .A(n18989), .Z(n18929) );
  XOR U27418 ( .A(n18915), .B(n18990), .Z(n18927) );
  XOR U27419 ( .A(n18916), .B(n18917), .Z(n18990) );
  XOR U27420 ( .A(n18922), .B(n18991), .Z(n18917) );
  XOR U27421 ( .A(n18921), .B(n18924), .Z(n18991) );
  IV U27422 ( .A(n18923), .Z(n18924) );
  NAND U27423 ( .A(n18992), .B(n18993), .Z(n18923) );
  OR U27424 ( .A(n18994), .B(n18995), .Z(n18993) );
  OR U27425 ( .A(n18996), .B(n18997), .Z(n18992) );
  NAND U27426 ( .A(n18998), .B(n18999), .Z(n18921) );
  OR U27427 ( .A(n19000), .B(n19001), .Z(n18999) );
  OR U27428 ( .A(n19002), .B(n19003), .Z(n18998) );
  NOR U27429 ( .A(n19004), .B(n19005), .Z(n18922) );
  ANDN U27430 ( .B(n19006), .A(n19007), .Z(n18916) );
  IV U27431 ( .A(n19008), .Z(n19006) );
  XNOR U27432 ( .A(n18909), .B(n19009), .Z(n18915) );
  XNOR U27433 ( .A(n18908), .B(n18910), .Z(n19009) );
  NAND U27434 ( .A(n19010), .B(n19011), .Z(n18910) );
  OR U27435 ( .A(n19012), .B(n19013), .Z(n19011) );
  OR U27436 ( .A(n19014), .B(n19015), .Z(n19010) );
  NAND U27437 ( .A(n19016), .B(n19017), .Z(n18908) );
  OR U27438 ( .A(n19018), .B(n19019), .Z(n19017) );
  OR U27439 ( .A(n19020), .B(n19021), .Z(n19016) );
  ANDN U27440 ( .B(n19022), .A(n19023), .Z(n18909) );
  IV U27441 ( .A(n19024), .Z(n19022) );
  XNOR U27442 ( .A(n18989), .B(n18988), .Z(N63712) );
  XOR U27443 ( .A(n19008), .B(n19007), .Z(n18988) );
  XNOR U27444 ( .A(n19023), .B(n19024), .Z(n19007) );
  XNOR U27445 ( .A(n19018), .B(n19019), .Z(n19024) );
  XNOR U27446 ( .A(n19020), .B(n19021), .Z(n19019) );
  XNOR U27447 ( .A(y[5773]), .B(x[5773]), .Z(n19021) );
  XNOR U27448 ( .A(y[5774]), .B(x[5774]), .Z(n19020) );
  XNOR U27449 ( .A(y[5772]), .B(x[5772]), .Z(n19018) );
  XNOR U27450 ( .A(n19012), .B(n19013), .Z(n19023) );
  XNOR U27451 ( .A(y[5769]), .B(x[5769]), .Z(n19013) );
  XNOR U27452 ( .A(n19014), .B(n19015), .Z(n19012) );
  XNOR U27453 ( .A(y[5770]), .B(x[5770]), .Z(n19015) );
  XNOR U27454 ( .A(y[5771]), .B(x[5771]), .Z(n19014) );
  XNOR U27455 ( .A(n19005), .B(n19004), .Z(n19008) );
  XNOR U27456 ( .A(n19000), .B(n19001), .Z(n19004) );
  XNOR U27457 ( .A(y[5766]), .B(x[5766]), .Z(n19001) );
  XNOR U27458 ( .A(n19002), .B(n19003), .Z(n19000) );
  XNOR U27459 ( .A(y[5767]), .B(x[5767]), .Z(n19003) );
  XNOR U27460 ( .A(y[5768]), .B(x[5768]), .Z(n19002) );
  XNOR U27461 ( .A(n18994), .B(n18995), .Z(n19005) );
  XNOR U27462 ( .A(y[5763]), .B(x[5763]), .Z(n18995) );
  XNOR U27463 ( .A(n18996), .B(n18997), .Z(n18994) );
  XNOR U27464 ( .A(y[5764]), .B(x[5764]), .Z(n18997) );
  XNOR U27465 ( .A(y[5765]), .B(x[5765]), .Z(n18996) );
  XOR U27466 ( .A(n18970), .B(n18971), .Z(n18989) );
  XNOR U27467 ( .A(n18986), .B(n18987), .Z(n18971) );
  XNOR U27468 ( .A(n18981), .B(n18982), .Z(n18987) );
  XNOR U27469 ( .A(n18983), .B(n18984), .Z(n18982) );
  XNOR U27470 ( .A(y[5761]), .B(x[5761]), .Z(n18984) );
  XNOR U27471 ( .A(y[5762]), .B(x[5762]), .Z(n18983) );
  XNOR U27472 ( .A(y[5760]), .B(x[5760]), .Z(n18981) );
  XNOR U27473 ( .A(n18975), .B(n18976), .Z(n18986) );
  XNOR U27474 ( .A(y[5757]), .B(x[5757]), .Z(n18976) );
  XNOR U27475 ( .A(n18977), .B(n18978), .Z(n18975) );
  XNOR U27476 ( .A(y[5758]), .B(x[5758]), .Z(n18978) );
  XNOR U27477 ( .A(y[5759]), .B(x[5759]), .Z(n18977) );
  XOR U27478 ( .A(n18969), .B(n18968), .Z(n18970) );
  XNOR U27479 ( .A(n18964), .B(n18965), .Z(n18968) );
  XNOR U27480 ( .A(y[5754]), .B(x[5754]), .Z(n18965) );
  XNOR U27481 ( .A(n18966), .B(n18967), .Z(n18964) );
  XNOR U27482 ( .A(y[5755]), .B(x[5755]), .Z(n18967) );
  XNOR U27483 ( .A(y[5756]), .B(x[5756]), .Z(n18966) );
  XNOR U27484 ( .A(n18958), .B(n18959), .Z(n18969) );
  XNOR U27485 ( .A(y[5751]), .B(x[5751]), .Z(n18959) );
  XNOR U27486 ( .A(n18960), .B(n18961), .Z(n18958) );
  XNOR U27487 ( .A(y[5752]), .B(x[5752]), .Z(n18961) );
  XNOR U27488 ( .A(y[5753]), .B(x[5753]), .Z(n18960) );
  NAND U27489 ( .A(n19025), .B(n19026), .Z(N63703) );
  NANDN U27490 ( .A(n19027), .B(n19028), .Z(n19026) );
  OR U27491 ( .A(n19029), .B(n19030), .Z(n19028) );
  NAND U27492 ( .A(n19029), .B(n19030), .Z(n19025) );
  XOR U27493 ( .A(n19029), .B(n19031), .Z(N63702) );
  XNOR U27494 ( .A(n19027), .B(n19030), .Z(n19031) );
  AND U27495 ( .A(n19032), .B(n19033), .Z(n19030) );
  NANDN U27496 ( .A(n19034), .B(n19035), .Z(n19033) );
  NANDN U27497 ( .A(n19036), .B(n19037), .Z(n19035) );
  NANDN U27498 ( .A(n19037), .B(n19036), .Z(n19032) );
  NAND U27499 ( .A(n19038), .B(n19039), .Z(n19027) );
  NANDN U27500 ( .A(n19040), .B(n19041), .Z(n19039) );
  OR U27501 ( .A(n19042), .B(n19043), .Z(n19041) );
  NAND U27502 ( .A(n19043), .B(n19042), .Z(n19038) );
  AND U27503 ( .A(n19044), .B(n19045), .Z(n19029) );
  NANDN U27504 ( .A(n19046), .B(n19047), .Z(n19045) );
  NANDN U27505 ( .A(n19048), .B(n19049), .Z(n19047) );
  NANDN U27506 ( .A(n19049), .B(n19048), .Z(n19044) );
  XOR U27507 ( .A(n19043), .B(n19050), .Z(N63701) );
  XOR U27508 ( .A(n19040), .B(n19042), .Z(n19050) );
  XNOR U27509 ( .A(n19036), .B(n19051), .Z(n19042) );
  XNOR U27510 ( .A(n19034), .B(n19037), .Z(n19051) );
  NAND U27511 ( .A(n19052), .B(n19053), .Z(n19037) );
  NAND U27512 ( .A(n19054), .B(n19055), .Z(n19053) );
  OR U27513 ( .A(n19056), .B(n19057), .Z(n19054) );
  NANDN U27514 ( .A(n19058), .B(n19056), .Z(n19052) );
  IV U27515 ( .A(n19057), .Z(n19058) );
  NAND U27516 ( .A(n19059), .B(n19060), .Z(n19034) );
  NAND U27517 ( .A(n19061), .B(n19062), .Z(n19060) );
  NANDN U27518 ( .A(n19063), .B(n19064), .Z(n19061) );
  NANDN U27519 ( .A(n19064), .B(n19063), .Z(n19059) );
  AND U27520 ( .A(n19065), .B(n19066), .Z(n19036) );
  NAND U27521 ( .A(n19067), .B(n19068), .Z(n19066) );
  OR U27522 ( .A(n19069), .B(n19070), .Z(n19067) );
  NANDN U27523 ( .A(n19071), .B(n19069), .Z(n19065) );
  NAND U27524 ( .A(n19072), .B(n19073), .Z(n19040) );
  NANDN U27525 ( .A(n19074), .B(n19075), .Z(n19073) );
  OR U27526 ( .A(n19076), .B(n19077), .Z(n19075) );
  NANDN U27527 ( .A(n19078), .B(n19076), .Z(n19072) );
  IV U27528 ( .A(n19077), .Z(n19078) );
  XNOR U27529 ( .A(n19048), .B(n19079), .Z(n19043) );
  XNOR U27530 ( .A(n19046), .B(n19049), .Z(n19079) );
  NAND U27531 ( .A(n19080), .B(n19081), .Z(n19049) );
  NAND U27532 ( .A(n19082), .B(n19083), .Z(n19081) );
  OR U27533 ( .A(n19084), .B(n19085), .Z(n19082) );
  NANDN U27534 ( .A(n19086), .B(n19084), .Z(n19080) );
  IV U27535 ( .A(n19085), .Z(n19086) );
  NAND U27536 ( .A(n19087), .B(n19088), .Z(n19046) );
  NAND U27537 ( .A(n19089), .B(n19090), .Z(n19088) );
  NANDN U27538 ( .A(n19091), .B(n19092), .Z(n19089) );
  NANDN U27539 ( .A(n19092), .B(n19091), .Z(n19087) );
  AND U27540 ( .A(n19093), .B(n19094), .Z(n19048) );
  NAND U27541 ( .A(n19095), .B(n19096), .Z(n19094) );
  OR U27542 ( .A(n19097), .B(n19098), .Z(n19095) );
  NANDN U27543 ( .A(n19099), .B(n19097), .Z(n19093) );
  XNOR U27544 ( .A(n19074), .B(n19100), .Z(N63700) );
  XOR U27545 ( .A(n19076), .B(n19077), .Z(n19100) );
  XNOR U27546 ( .A(n19090), .B(n19101), .Z(n19077) );
  XOR U27547 ( .A(n19091), .B(n19092), .Z(n19101) );
  XOR U27548 ( .A(n19097), .B(n19102), .Z(n19092) );
  XOR U27549 ( .A(n19096), .B(n19099), .Z(n19102) );
  IV U27550 ( .A(n19098), .Z(n19099) );
  NAND U27551 ( .A(n19103), .B(n19104), .Z(n19098) );
  OR U27552 ( .A(n19105), .B(n19106), .Z(n19104) );
  OR U27553 ( .A(n19107), .B(n19108), .Z(n19103) );
  NAND U27554 ( .A(n19109), .B(n19110), .Z(n19096) );
  OR U27555 ( .A(n19111), .B(n19112), .Z(n19110) );
  OR U27556 ( .A(n19113), .B(n19114), .Z(n19109) );
  NOR U27557 ( .A(n19115), .B(n19116), .Z(n19097) );
  ANDN U27558 ( .B(n19117), .A(n19118), .Z(n19091) );
  XNOR U27559 ( .A(n19084), .B(n19119), .Z(n19090) );
  XNOR U27560 ( .A(n19083), .B(n19085), .Z(n19119) );
  NAND U27561 ( .A(n19120), .B(n19121), .Z(n19085) );
  OR U27562 ( .A(n19122), .B(n19123), .Z(n19121) );
  OR U27563 ( .A(n19124), .B(n19125), .Z(n19120) );
  NAND U27564 ( .A(n19126), .B(n19127), .Z(n19083) );
  OR U27565 ( .A(n19128), .B(n19129), .Z(n19127) );
  OR U27566 ( .A(n19130), .B(n19131), .Z(n19126) );
  ANDN U27567 ( .B(n19132), .A(n19133), .Z(n19084) );
  IV U27568 ( .A(n19134), .Z(n19132) );
  ANDN U27569 ( .B(n19135), .A(n19136), .Z(n19076) );
  XOR U27570 ( .A(n19062), .B(n19137), .Z(n19074) );
  XOR U27571 ( .A(n19063), .B(n19064), .Z(n19137) );
  XOR U27572 ( .A(n19069), .B(n19138), .Z(n19064) );
  XOR U27573 ( .A(n19068), .B(n19071), .Z(n19138) );
  IV U27574 ( .A(n19070), .Z(n19071) );
  NAND U27575 ( .A(n19139), .B(n19140), .Z(n19070) );
  OR U27576 ( .A(n19141), .B(n19142), .Z(n19140) );
  OR U27577 ( .A(n19143), .B(n19144), .Z(n19139) );
  NAND U27578 ( .A(n19145), .B(n19146), .Z(n19068) );
  OR U27579 ( .A(n19147), .B(n19148), .Z(n19146) );
  OR U27580 ( .A(n19149), .B(n19150), .Z(n19145) );
  NOR U27581 ( .A(n19151), .B(n19152), .Z(n19069) );
  ANDN U27582 ( .B(n19153), .A(n19154), .Z(n19063) );
  IV U27583 ( .A(n19155), .Z(n19153) );
  XNOR U27584 ( .A(n19056), .B(n19156), .Z(n19062) );
  XNOR U27585 ( .A(n19055), .B(n19057), .Z(n19156) );
  NAND U27586 ( .A(n19157), .B(n19158), .Z(n19057) );
  OR U27587 ( .A(n19159), .B(n19160), .Z(n19158) );
  OR U27588 ( .A(n19161), .B(n19162), .Z(n19157) );
  NAND U27589 ( .A(n19163), .B(n19164), .Z(n19055) );
  OR U27590 ( .A(n19165), .B(n19166), .Z(n19164) );
  OR U27591 ( .A(n19167), .B(n19168), .Z(n19163) );
  ANDN U27592 ( .B(n19169), .A(n19170), .Z(n19056) );
  IV U27593 ( .A(n19171), .Z(n19169) );
  XNOR U27594 ( .A(n19136), .B(n19135), .Z(N63699) );
  XOR U27595 ( .A(n19155), .B(n19154), .Z(n19135) );
  XNOR U27596 ( .A(n19170), .B(n19171), .Z(n19154) );
  XNOR U27597 ( .A(n19165), .B(n19166), .Z(n19171) );
  XNOR U27598 ( .A(n19167), .B(n19168), .Z(n19166) );
  XNOR U27599 ( .A(y[5749]), .B(x[5749]), .Z(n19168) );
  XNOR U27600 ( .A(y[5750]), .B(x[5750]), .Z(n19167) );
  XNOR U27601 ( .A(y[5748]), .B(x[5748]), .Z(n19165) );
  XNOR U27602 ( .A(n19159), .B(n19160), .Z(n19170) );
  XNOR U27603 ( .A(y[5745]), .B(x[5745]), .Z(n19160) );
  XNOR U27604 ( .A(n19161), .B(n19162), .Z(n19159) );
  XNOR U27605 ( .A(y[5746]), .B(x[5746]), .Z(n19162) );
  XNOR U27606 ( .A(y[5747]), .B(x[5747]), .Z(n19161) );
  XNOR U27607 ( .A(n19152), .B(n19151), .Z(n19155) );
  XNOR U27608 ( .A(n19147), .B(n19148), .Z(n19151) );
  XNOR U27609 ( .A(y[5742]), .B(x[5742]), .Z(n19148) );
  XNOR U27610 ( .A(n19149), .B(n19150), .Z(n19147) );
  XNOR U27611 ( .A(y[5743]), .B(x[5743]), .Z(n19150) );
  XNOR U27612 ( .A(y[5744]), .B(x[5744]), .Z(n19149) );
  XNOR U27613 ( .A(n19141), .B(n19142), .Z(n19152) );
  XNOR U27614 ( .A(y[5739]), .B(x[5739]), .Z(n19142) );
  XNOR U27615 ( .A(n19143), .B(n19144), .Z(n19141) );
  XNOR U27616 ( .A(y[5740]), .B(x[5740]), .Z(n19144) );
  XNOR U27617 ( .A(y[5741]), .B(x[5741]), .Z(n19143) );
  XOR U27618 ( .A(n19117), .B(n19118), .Z(n19136) );
  XNOR U27619 ( .A(n19133), .B(n19134), .Z(n19118) );
  XNOR U27620 ( .A(n19128), .B(n19129), .Z(n19134) );
  XNOR U27621 ( .A(n19130), .B(n19131), .Z(n19129) );
  XNOR U27622 ( .A(y[5737]), .B(x[5737]), .Z(n19131) );
  XNOR U27623 ( .A(y[5738]), .B(x[5738]), .Z(n19130) );
  XNOR U27624 ( .A(y[5736]), .B(x[5736]), .Z(n19128) );
  XNOR U27625 ( .A(n19122), .B(n19123), .Z(n19133) );
  XNOR U27626 ( .A(y[5733]), .B(x[5733]), .Z(n19123) );
  XNOR U27627 ( .A(n19124), .B(n19125), .Z(n19122) );
  XNOR U27628 ( .A(y[5734]), .B(x[5734]), .Z(n19125) );
  XNOR U27629 ( .A(y[5735]), .B(x[5735]), .Z(n19124) );
  XOR U27630 ( .A(n19116), .B(n19115), .Z(n19117) );
  XNOR U27631 ( .A(n19111), .B(n19112), .Z(n19115) );
  XNOR U27632 ( .A(y[5730]), .B(x[5730]), .Z(n19112) );
  XNOR U27633 ( .A(n19113), .B(n19114), .Z(n19111) );
  XNOR U27634 ( .A(y[5731]), .B(x[5731]), .Z(n19114) );
  XNOR U27635 ( .A(y[5732]), .B(x[5732]), .Z(n19113) );
  XNOR U27636 ( .A(n19105), .B(n19106), .Z(n19116) );
  XNOR U27637 ( .A(y[5727]), .B(x[5727]), .Z(n19106) );
  XNOR U27638 ( .A(n19107), .B(n19108), .Z(n19105) );
  XNOR U27639 ( .A(y[5728]), .B(x[5728]), .Z(n19108) );
  XNOR U27640 ( .A(y[5729]), .B(x[5729]), .Z(n19107) );
  NAND U27641 ( .A(n19172), .B(n19173), .Z(N63690) );
  NANDN U27642 ( .A(n19174), .B(n19175), .Z(n19173) );
  OR U27643 ( .A(n19176), .B(n19177), .Z(n19175) );
  NAND U27644 ( .A(n19176), .B(n19177), .Z(n19172) );
  XOR U27645 ( .A(n19176), .B(n19178), .Z(N63689) );
  XNOR U27646 ( .A(n19174), .B(n19177), .Z(n19178) );
  AND U27647 ( .A(n19179), .B(n19180), .Z(n19177) );
  NANDN U27648 ( .A(n19181), .B(n19182), .Z(n19180) );
  NANDN U27649 ( .A(n19183), .B(n19184), .Z(n19182) );
  NANDN U27650 ( .A(n19184), .B(n19183), .Z(n19179) );
  NAND U27651 ( .A(n19185), .B(n19186), .Z(n19174) );
  NANDN U27652 ( .A(n19187), .B(n19188), .Z(n19186) );
  OR U27653 ( .A(n19189), .B(n19190), .Z(n19188) );
  NAND U27654 ( .A(n19190), .B(n19189), .Z(n19185) );
  AND U27655 ( .A(n19191), .B(n19192), .Z(n19176) );
  NANDN U27656 ( .A(n19193), .B(n19194), .Z(n19192) );
  NANDN U27657 ( .A(n19195), .B(n19196), .Z(n19194) );
  NANDN U27658 ( .A(n19196), .B(n19195), .Z(n19191) );
  XOR U27659 ( .A(n19190), .B(n19197), .Z(N63688) );
  XOR U27660 ( .A(n19187), .B(n19189), .Z(n19197) );
  XNOR U27661 ( .A(n19183), .B(n19198), .Z(n19189) );
  XNOR U27662 ( .A(n19181), .B(n19184), .Z(n19198) );
  NAND U27663 ( .A(n19199), .B(n19200), .Z(n19184) );
  NAND U27664 ( .A(n19201), .B(n19202), .Z(n19200) );
  OR U27665 ( .A(n19203), .B(n19204), .Z(n19201) );
  NANDN U27666 ( .A(n19205), .B(n19203), .Z(n19199) );
  IV U27667 ( .A(n19204), .Z(n19205) );
  NAND U27668 ( .A(n19206), .B(n19207), .Z(n19181) );
  NAND U27669 ( .A(n19208), .B(n19209), .Z(n19207) );
  NANDN U27670 ( .A(n19210), .B(n19211), .Z(n19208) );
  NANDN U27671 ( .A(n19211), .B(n19210), .Z(n19206) );
  AND U27672 ( .A(n19212), .B(n19213), .Z(n19183) );
  NAND U27673 ( .A(n19214), .B(n19215), .Z(n19213) );
  OR U27674 ( .A(n19216), .B(n19217), .Z(n19214) );
  NANDN U27675 ( .A(n19218), .B(n19216), .Z(n19212) );
  NAND U27676 ( .A(n19219), .B(n19220), .Z(n19187) );
  NANDN U27677 ( .A(n19221), .B(n19222), .Z(n19220) );
  OR U27678 ( .A(n19223), .B(n19224), .Z(n19222) );
  NANDN U27679 ( .A(n19225), .B(n19223), .Z(n19219) );
  IV U27680 ( .A(n19224), .Z(n19225) );
  XNOR U27681 ( .A(n19195), .B(n19226), .Z(n19190) );
  XNOR U27682 ( .A(n19193), .B(n19196), .Z(n19226) );
  NAND U27683 ( .A(n19227), .B(n19228), .Z(n19196) );
  NAND U27684 ( .A(n19229), .B(n19230), .Z(n19228) );
  OR U27685 ( .A(n19231), .B(n19232), .Z(n19229) );
  NANDN U27686 ( .A(n19233), .B(n19231), .Z(n19227) );
  IV U27687 ( .A(n19232), .Z(n19233) );
  NAND U27688 ( .A(n19234), .B(n19235), .Z(n19193) );
  NAND U27689 ( .A(n19236), .B(n19237), .Z(n19235) );
  NANDN U27690 ( .A(n19238), .B(n19239), .Z(n19236) );
  NANDN U27691 ( .A(n19239), .B(n19238), .Z(n19234) );
  AND U27692 ( .A(n19240), .B(n19241), .Z(n19195) );
  NAND U27693 ( .A(n19242), .B(n19243), .Z(n19241) );
  OR U27694 ( .A(n19244), .B(n19245), .Z(n19242) );
  NANDN U27695 ( .A(n19246), .B(n19244), .Z(n19240) );
  XNOR U27696 ( .A(n19221), .B(n19247), .Z(N63687) );
  XOR U27697 ( .A(n19223), .B(n19224), .Z(n19247) );
  XNOR U27698 ( .A(n19237), .B(n19248), .Z(n19224) );
  XOR U27699 ( .A(n19238), .B(n19239), .Z(n19248) );
  XOR U27700 ( .A(n19244), .B(n19249), .Z(n19239) );
  XOR U27701 ( .A(n19243), .B(n19246), .Z(n19249) );
  IV U27702 ( .A(n19245), .Z(n19246) );
  NAND U27703 ( .A(n19250), .B(n19251), .Z(n19245) );
  OR U27704 ( .A(n19252), .B(n19253), .Z(n19251) );
  OR U27705 ( .A(n19254), .B(n19255), .Z(n19250) );
  NAND U27706 ( .A(n19256), .B(n19257), .Z(n19243) );
  OR U27707 ( .A(n19258), .B(n19259), .Z(n19257) );
  OR U27708 ( .A(n19260), .B(n19261), .Z(n19256) );
  NOR U27709 ( .A(n19262), .B(n19263), .Z(n19244) );
  ANDN U27710 ( .B(n19264), .A(n19265), .Z(n19238) );
  XNOR U27711 ( .A(n19231), .B(n19266), .Z(n19237) );
  XNOR U27712 ( .A(n19230), .B(n19232), .Z(n19266) );
  NAND U27713 ( .A(n19267), .B(n19268), .Z(n19232) );
  OR U27714 ( .A(n19269), .B(n19270), .Z(n19268) );
  OR U27715 ( .A(n19271), .B(n19272), .Z(n19267) );
  NAND U27716 ( .A(n19273), .B(n19274), .Z(n19230) );
  OR U27717 ( .A(n19275), .B(n19276), .Z(n19274) );
  OR U27718 ( .A(n19277), .B(n19278), .Z(n19273) );
  ANDN U27719 ( .B(n19279), .A(n19280), .Z(n19231) );
  IV U27720 ( .A(n19281), .Z(n19279) );
  ANDN U27721 ( .B(n19282), .A(n19283), .Z(n19223) );
  XOR U27722 ( .A(n19209), .B(n19284), .Z(n19221) );
  XOR U27723 ( .A(n19210), .B(n19211), .Z(n19284) );
  XOR U27724 ( .A(n19216), .B(n19285), .Z(n19211) );
  XOR U27725 ( .A(n19215), .B(n19218), .Z(n19285) );
  IV U27726 ( .A(n19217), .Z(n19218) );
  NAND U27727 ( .A(n19286), .B(n19287), .Z(n19217) );
  OR U27728 ( .A(n19288), .B(n19289), .Z(n19287) );
  OR U27729 ( .A(n19290), .B(n19291), .Z(n19286) );
  NAND U27730 ( .A(n19292), .B(n19293), .Z(n19215) );
  OR U27731 ( .A(n19294), .B(n19295), .Z(n19293) );
  OR U27732 ( .A(n19296), .B(n19297), .Z(n19292) );
  NOR U27733 ( .A(n19298), .B(n19299), .Z(n19216) );
  ANDN U27734 ( .B(n19300), .A(n19301), .Z(n19210) );
  IV U27735 ( .A(n19302), .Z(n19300) );
  XNOR U27736 ( .A(n19203), .B(n19303), .Z(n19209) );
  XNOR U27737 ( .A(n19202), .B(n19204), .Z(n19303) );
  NAND U27738 ( .A(n19304), .B(n19305), .Z(n19204) );
  OR U27739 ( .A(n19306), .B(n19307), .Z(n19305) );
  OR U27740 ( .A(n19308), .B(n19309), .Z(n19304) );
  NAND U27741 ( .A(n19310), .B(n19311), .Z(n19202) );
  OR U27742 ( .A(n19312), .B(n19313), .Z(n19311) );
  OR U27743 ( .A(n19314), .B(n19315), .Z(n19310) );
  ANDN U27744 ( .B(n19316), .A(n19317), .Z(n19203) );
  IV U27745 ( .A(n19318), .Z(n19316) );
  XNOR U27746 ( .A(n19283), .B(n19282), .Z(N63686) );
  XOR U27747 ( .A(n19302), .B(n19301), .Z(n19282) );
  XNOR U27748 ( .A(n19317), .B(n19318), .Z(n19301) );
  XNOR U27749 ( .A(n19312), .B(n19313), .Z(n19318) );
  XNOR U27750 ( .A(n19314), .B(n19315), .Z(n19313) );
  XNOR U27751 ( .A(y[5725]), .B(x[5725]), .Z(n19315) );
  XNOR U27752 ( .A(y[5726]), .B(x[5726]), .Z(n19314) );
  XNOR U27753 ( .A(y[5724]), .B(x[5724]), .Z(n19312) );
  XNOR U27754 ( .A(n19306), .B(n19307), .Z(n19317) );
  XNOR U27755 ( .A(y[5721]), .B(x[5721]), .Z(n19307) );
  XNOR U27756 ( .A(n19308), .B(n19309), .Z(n19306) );
  XNOR U27757 ( .A(y[5722]), .B(x[5722]), .Z(n19309) );
  XNOR U27758 ( .A(y[5723]), .B(x[5723]), .Z(n19308) );
  XNOR U27759 ( .A(n19299), .B(n19298), .Z(n19302) );
  XNOR U27760 ( .A(n19294), .B(n19295), .Z(n19298) );
  XNOR U27761 ( .A(y[5718]), .B(x[5718]), .Z(n19295) );
  XNOR U27762 ( .A(n19296), .B(n19297), .Z(n19294) );
  XNOR U27763 ( .A(y[5719]), .B(x[5719]), .Z(n19297) );
  XNOR U27764 ( .A(y[5720]), .B(x[5720]), .Z(n19296) );
  XNOR U27765 ( .A(n19288), .B(n19289), .Z(n19299) );
  XNOR U27766 ( .A(y[5715]), .B(x[5715]), .Z(n19289) );
  XNOR U27767 ( .A(n19290), .B(n19291), .Z(n19288) );
  XNOR U27768 ( .A(y[5716]), .B(x[5716]), .Z(n19291) );
  XNOR U27769 ( .A(y[5717]), .B(x[5717]), .Z(n19290) );
  XOR U27770 ( .A(n19264), .B(n19265), .Z(n19283) );
  XNOR U27771 ( .A(n19280), .B(n19281), .Z(n19265) );
  XNOR U27772 ( .A(n19275), .B(n19276), .Z(n19281) );
  XNOR U27773 ( .A(n19277), .B(n19278), .Z(n19276) );
  XNOR U27774 ( .A(y[5713]), .B(x[5713]), .Z(n19278) );
  XNOR U27775 ( .A(y[5714]), .B(x[5714]), .Z(n19277) );
  XNOR U27776 ( .A(y[5712]), .B(x[5712]), .Z(n19275) );
  XNOR U27777 ( .A(n19269), .B(n19270), .Z(n19280) );
  XNOR U27778 ( .A(y[5709]), .B(x[5709]), .Z(n19270) );
  XNOR U27779 ( .A(n19271), .B(n19272), .Z(n19269) );
  XNOR U27780 ( .A(y[5710]), .B(x[5710]), .Z(n19272) );
  XNOR U27781 ( .A(y[5711]), .B(x[5711]), .Z(n19271) );
  XOR U27782 ( .A(n19263), .B(n19262), .Z(n19264) );
  XNOR U27783 ( .A(n19258), .B(n19259), .Z(n19262) );
  XNOR U27784 ( .A(y[5706]), .B(x[5706]), .Z(n19259) );
  XNOR U27785 ( .A(n19260), .B(n19261), .Z(n19258) );
  XNOR U27786 ( .A(y[5707]), .B(x[5707]), .Z(n19261) );
  XNOR U27787 ( .A(y[5708]), .B(x[5708]), .Z(n19260) );
  XNOR U27788 ( .A(n19252), .B(n19253), .Z(n19263) );
  XNOR U27789 ( .A(y[5703]), .B(x[5703]), .Z(n19253) );
  XNOR U27790 ( .A(n19254), .B(n19255), .Z(n19252) );
  XNOR U27791 ( .A(y[5704]), .B(x[5704]), .Z(n19255) );
  XNOR U27792 ( .A(y[5705]), .B(x[5705]), .Z(n19254) );
  NAND U27793 ( .A(n19319), .B(n19320), .Z(N63677) );
  NANDN U27794 ( .A(n19321), .B(n19322), .Z(n19320) );
  OR U27795 ( .A(n19323), .B(n19324), .Z(n19322) );
  NAND U27796 ( .A(n19323), .B(n19324), .Z(n19319) );
  XOR U27797 ( .A(n19323), .B(n19325), .Z(N63676) );
  XNOR U27798 ( .A(n19321), .B(n19324), .Z(n19325) );
  AND U27799 ( .A(n19326), .B(n19327), .Z(n19324) );
  NANDN U27800 ( .A(n19328), .B(n19329), .Z(n19327) );
  NANDN U27801 ( .A(n19330), .B(n19331), .Z(n19329) );
  NANDN U27802 ( .A(n19331), .B(n19330), .Z(n19326) );
  NAND U27803 ( .A(n19332), .B(n19333), .Z(n19321) );
  NANDN U27804 ( .A(n19334), .B(n19335), .Z(n19333) );
  OR U27805 ( .A(n19336), .B(n19337), .Z(n19335) );
  NAND U27806 ( .A(n19337), .B(n19336), .Z(n19332) );
  AND U27807 ( .A(n19338), .B(n19339), .Z(n19323) );
  NANDN U27808 ( .A(n19340), .B(n19341), .Z(n19339) );
  NANDN U27809 ( .A(n19342), .B(n19343), .Z(n19341) );
  NANDN U27810 ( .A(n19343), .B(n19342), .Z(n19338) );
  XOR U27811 ( .A(n19337), .B(n19344), .Z(N63675) );
  XOR U27812 ( .A(n19334), .B(n19336), .Z(n19344) );
  XNOR U27813 ( .A(n19330), .B(n19345), .Z(n19336) );
  XNOR U27814 ( .A(n19328), .B(n19331), .Z(n19345) );
  NAND U27815 ( .A(n19346), .B(n19347), .Z(n19331) );
  NAND U27816 ( .A(n19348), .B(n19349), .Z(n19347) );
  OR U27817 ( .A(n19350), .B(n19351), .Z(n19348) );
  NANDN U27818 ( .A(n19352), .B(n19350), .Z(n19346) );
  IV U27819 ( .A(n19351), .Z(n19352) );
  NAND U27820 ( .A(n19353), .B(n19354), .Z(n19328) );
  NAND U27821 ( .A(n19355), .B(n19356), .Z(n19354) );
  NANDN U27822 ( .A(n19357), .B(n19358), .Z(n19355) );
  NANDN U27823 ( .A(n19358), .B(n19357), .Z(n19353) );
  AND U27824 ( .A(n19359), .B(n19360), .Z(n19330) );
  NAND U27825 ( .A(n19361), .B(n19362), .Z(n19360) );
  OR U27826 ( .A(n19363), .B(n19364), .Z(n19361) );
  NANDN U27827 ( .A(n19365), .B(n19363), .Z(n19359) );
  NAND U27828 ( .A(n19366), .B(n19367), .Z(n19334) );
  NANDN U27829 ( .A(n19368), .B(n19369), .Z(n19367) );
  OR U27830 ( .A(n19370), .B(n19371), .Z(n19369) );
  NANDN U27831 ( .A(n19372), .B(n19370), .Z(n19366) );
  IV U27832 ( .A(n19371), .Z(n19372) );
  XNOR U27833 ( .A(n19342), .B(n19373), .Z(n19337) );
  XNOR U27834 ( .A(n19340), .B(n19343), .Z(n19373) );
  NAND U27835 ( .A(n19374), .B(n19375), .Z(n19343) );
  NAND U27836 ( .A(n19376), .B(n19377), .Z(n19375) );
  OR U27837 ( .A(n19378), .B(n19379), .Z(n19376) );
  NANDN U27838 ( .A(n19380), .B(n19378), .Z(n19374) );
  IV U27839 ( .A(n19379), .Z(n19380) );
  NAND U27840 ( .A(n19381), .B(n19382), .Z(n19340) );
  NAND U27841 ( .A(n19383), .B(n19384), .Z(n19382) );
  NANDN U27842 ( .A(n19385), .B(n19386), .Z(n19383) );
  NANDN U27843 ( .A(n19386), .B(n19385), .Z(n19381) );
  AND U27844 ( .A(n19387), .B(n19388), .Z(n19342) );
  NAND U27845 ( .A(n19389), .B(n19390), .Z(n19388) );
  OR U27846 ( .A(n19391), .B(n19392), .Z(n19389) );
  NANDN U27847 ( .A(n19393), .B(n19391), .Z(n19387) );
  XNOR U27848 ( .A(n19368), .B(n19394), .Z(N63674) );
  XOR U27849 ( .A(n19370), .B(n19371), .Z(n19394) );
  XNOR U27850 ( .A(n19384), .B(n19395), .Z(n19371) );
  XOR U27851 ( .A(n19385), .B(n19386), .Z(n19395) );
  XOR U27852 ( .A(n19391), .B(n19396), .Z(n19386) );
  XOR U27853 ( .A(n19390), .B(n19393), .Z(n19396) );
  IV U27854 ( .A(n19392), .Z(n19393) );
  NAND U27855 ( .A(n19397), .B(n19398), .Z(n19392) );
  OR U27856 ( .A(n19399), .B(n19400), .Z(n19398) );
  OR U27857 ( .A(n19401), .B(n19402), .Z(n19397) );
  NAND U27858 ( .A(n19403), .B(n19404), .Z(n19390) );
  OR U27859 ( .A(n19405), .B(n19406), .Z(n19404) );
  OR U27860 ( .A(n19407), .B(n19408), .Z(n19403) );
  NOR U27861 ( .A(n19409), .B(n19410), .Z(n19391) );
  ANDN U27862 ( .B(n19411), .A(n19412), .Z(n19385) );
  XNOR U27863 ( .A(n19378), .B(n19413), .Z(n19384) );
  XNOR U27864 ( .A(n19377), .B(n19379), .Z(n19413) );
  NAND U27865 ( .A(n19414), .B(n19415), .Z(n19379) );
  OR U27866 ( .A(n19416), .B(n19417), .Z(n19415) );
  OR U27867 ( .A(n19418), .B(n19419), .Z(n19414) );
  NAND U27868 ( .A(n19420), .B(n19421), .Z(n19377) );
  OR U27869 ( .A(n19422), .B(n19423), .Z(n19421) );
  OR U27870 ( .A(n19424), .B(n19425), .Z(n19420) );
  ANDN U27871 ( .B(n19426), .A(n19427), .Z(n19378) );
  IV U27872 ( .A(n19428), .Z(n19426) );
  ANDN U27873 ( .B(n19429), .A(n19430), .Z(n19370) );
  XOR U27874 ( .A(n19356), .B(n19431), .Z(n19368) );
  XOR U27875 ( .A(n19357), .B(n19358), .Z(n19431) );
  XOR U27876 ( .A(n19363), .B(n19432), .Z(n19358) );
  XOR U27877 ( .A(n19362), .B(n19365), .Z(n19432) );
  IV U27878 ( .A(n19364), .Z(n19365) );
  NAND U27879 ( .A(n19433), .B(n19434), .Z(n19364) );
  OR U27880 ( .A(n19435), .B(n19436), .Z(n19434) );
  OR U27881 ( .A(n19437), .B(n19438), .Z(n19433) );
  NAND U27882 ( .A(n19439), .B(n19440), .Z(n19362) );
  OR U27883 ( .A(n19441), .B(n19442), .Z(n19440) );
  OR U27884 ( .A(n19443), .B(n19444), .Z(n19439) );
  NOR U27885 ( .A(n19445), .B(n19446), .Z(n19363) );
  ANDN U27886 ( .B(n19447), .A(n19448), .Z(n19357) );
  IV U27887 ( .A(n19449), .Z(n19447) );
  XNOR U27888 ( .A(n19350), .B(n19450), .Z(n19356) );
  XNOR U27889 ( .A(n19349), .B(n19351), .Z(n19450) );
  NAND U27890 ( .A(n19451), .B(n19452), .Z(n19351) );
  OR U27891 ( .A(n19453), .B(n19454), .Z(n19452) );
  OR U27892 ( .A(n19455), .B(n19456), .Z(n19451) );
  NAND U27893 ( .A(n19457), .B(n19458), .Z(n19349) );
  OR U27894 ( .A(n19459), .B(n19460), .Z(n19458) );
  OR U27895 ( .A(n19461), .B(n19462), .Z(n19457) );
  ANDN U27896 ( .B(n19463), .A(n19464), .Z(n19350) );
  IV U27897 ( .A(n19465), .Z(n19463) );
  XNOR U27898 ( .A(n19430), .B(n19429), .Z(N63673) );
  XOR U27899 ( .A(n19449), .B(n19448), .Z(n19429) );
  XNOR U27900 ( .A(n19464), .B(n19465), .Z(n19448) );
  XNOR U27901 ( .A(n19459), .B(n19460), .Z(n19465) );
  XNOR U27902 ( .A(n19461), .B(n19462), .Z(n19460) );
  XNOR U27903 ( .A(y[5701]), .B(x[5701]), .Z(n19462) );
  XNOR U27904 ( .A(y[5702]), .B(x[5702]), .Z(n19461) );
  XNOR U27905 ( .A(y[5700]), .B(x[5700]), .Z(n19459) );
  XNOR U27906 ( .A(n19453), .B(n19454), .Z(n19464) );
  XNOR U27907 ( .A(y[5697]), .B(x[5697]), .Z(n19454) );
  XNOR U27908 ( .A(n19455), .B(n19456), .Z(n19453) );
  XNOR U27909 ( .A(y[5698]), .B(x[5698]), .Z(n19456) );
  XNOR U27910 ( .A(y[5699]), .B(x[5699]), .Z(n19455) );
  XNOR U27911 ( .A(n19446), .B(n19445), .Z(n19449) );
  XNOR U27912 ( .A(n19441), .B(n19442), .Z(n19445) );
  XNOR U27913 ( .A(y[5694]), .B(x[5694]), .Z(n19442) );
  XNOR U27914 ( .A(n19443), .B(n19444), .Z(n19441) );
  XNOR U27915 ( .A(y[5695]), .B(x[5695]), .Z(n19444) );
  XNOR U27916 ( .A(y[5696]), .B(x[5696]), .Z(n19443) );
  XNOR U27917 ( .A(n19435), .B(n19436), .Z(n19446) );
  XNOR U27918 ( .A(y[5691]), .B(x[5691]), .Z(n19436) );
  XNOR U27919 ( .A(n19437), .B(n19438), .Z(n19435) );
  XNOR U27920 ( .A(y[5692]), .B(x[5692]), .Z(n19438) );
  XNOR U27921 ( .A(y[5693]), .B(x[5693]), .Z(n19437) );
  XOR U27922 ( .A(n19411), .B(n19412), .Z(n19430) );
  XNOR U27923 ( .A(n19427), .B(n19428), .Z(n19412) );
  XNOR U27924 ( .A(n19422), .B(n19423), .Z(n19428) );
  XNOR U27925 ( .A(n19424), .B(n19425), .Z(n19423) );
  XNOR U27926 ( .A(y[5689]), .B(x[5689]), .Z(n19425) );
  XNOR U27927 ( .A(y[5690]), .B(x[5690]), .Z(n19424) );
  XNOR U27928 ( .A(y[5688]), .B(x[5688]), .Z(n19422) );
  XNOR U27929 ( .A(n19416), .B(n19417), .Z(n19427) );
  XNOR U27930 ( .A(y[5685]), .B(x[5685]), .Z(n19417) );
  XNOR U27931 ( .A(n19418), .B(n19419), .Z(n19416) );
  XNOR U27932 ( .A(y[5686]), .B(x[5686]), .Z(n19419) );
  XNOR U27933 ( .A(y[5687]), .B(x[5687]), .Z(n19418) );
  XOR U27934 ( .A(n19410), .B(n19409), .Z(n19411) );
  XNOR U27935 ( .A(n19405), .B(n19406), .Z(n19409) );
  XNOR U27936 ( .A(y[5682]), .B(x[5682]), .Z(n19406) );
  XNOR U27937 ( .A(n19407), .B(n19408), .Z(n19405) );
  XNOR U27938 ( .A(y[5683]), .B(x[5683]), .Z(n19408) );
  XNOR U27939 ( .A(y[5684]), .B(x[5684]), .Z(n19407) );
  XNOR U27940 ( .A(n19399), .B(n19400), .Z(n19410) );
  XNOR U27941 ( .A(y[5679]), .B(x[5679]), .Z(n19400) );
  XNOR U27942 ( .A(n19401), .B(n19402), .Z(n19399) );
  XNOR U27943 ( .A(y[5680]), .B(x[5680]), .Z(n19402) );
  XNOR U27944 ( .A(y[5681]), .B(x[5681]), .Z(n19401) );
  NAND U27945 ( .A(n19466), .B(n19467), .Z(N63664) );
  NANDN U27946 ( .A(n19468), .B(n19469), .Z(n19467) );
  OR U27947 ( .A(n19470), .B(n19471), .Z(n19469) );
  NAND U27948 ( .A(n19470), .B(n19471), .Z(n19466) );
  XOR U27949 ( .A(n19470), .B(n19472), .Z(N63663) );
  XNOR U27950 ( .A(n19468), .B(n19471), .Z(n19472) );
  AND U27951 ( .A(n19473), .B(n19474), .Z(n19471) );
  NANDN U27952 ( .A(n19475), .B(n19476), .Z(n19474) );
  NANDN U27953 ( .A(n19477), .B(n19478), .Z(n19476) );
  NANDN U27954 ( .A(n19478), .B(n19477), .Z(n19473) );
  NAND U27955 ( .A(n19479), .B(n19480), .Z(n19468) );
  NANDN U27956 ( .A(n19481), .B(n19482), .Z(n19480) );
  OR U27957 ( .A(n19483), .B(n19484), .Z(n19482) );
  NAND U27958 ( .A(n19484), .B(n19483), .Z(n19479) );
  AND U27959 ( .A(n19485), .B(n19486), .Z(n19470) );
  NANDN U27960 ( .A(n19487), .B(n19488), .Z(n19486) );
  NANDN U27961 ( .A(n19489), .B(n19490), .Z(n19488) );
  NANDN U27962 ( .A(n19490), .B(n19489), .Z(n19485) );
  XOR U27963 ( .A(n19484), .B(n19491), .Z(N63662) );
  XOR U27964 ( .A(n19481), .B(n19483), .Z(n19491) );
  XNOR U27965 ( .A(n19477), .B(n19492), .Z(n19483) );
  XNOR U27966 ( .A(n19475), .B(n19478), .Z(n19492) );
  NAND U27967 ( .A(n19493), .B(n19494), .Z(n19478) );
  NAND U27968 ( .A(n19495), .B(n19496), .Z(n19494) );
  OR U27969 ( .A(n19497), .B(n19498), .Z(n19495) );
  NANDN U27970 ( .A(n19499), .B(n19497), .Z(n19493) );
  IV U27971 ( .A(n19498), .Z(n19499) );
  NAND U27972 ( .A(n19500), .B(n19501), .Z(n19475) );
  NAND U27973 ( .A(n19502), .B(n19503), .Z(n19501) );
  NANDN U27974 ( .A(n19504), .B(n19505), .Z(n19502) );
  NANDN U27975 ( .A(n19505), .B(n19504), .Z(n19500) );
  AND U27976 ( .A(n19506), .B(n19507), .Z(n19477) );
  NAND U27977 ( .A(n19508), .B(n19509), .Z(n19507) );
  OR U27978 ( .A(n19510), .B(n19511), .Z(n19508) );
  NANDN U27979 ( .A(n19512), .B(n19510), .Z(n19506) );
  NAND U27980 ( .A(n19513), .B(n19514), .Z(n19481) );
  NANDN U27981 ( .A(n19515), .B(n19516), .Z(n19514) );
  OR U27982 ( .A(n19517), .B(n19518), .Z(n19516) );
  NANDN U27983 ( .A(n19519), .B(n19517), .Z(n19513) );
  IV U27984 ( .A(n19518), .Z(n19519) );
  XNOR U27985 ( .A(n19489), .B(n19520), .Z(n19484) );
  XNOR U27986 ( .A(n19487), .B(n19490), .Z(n19520) );
  NAND U27987 ( .A(n19521), .B(n19522), .Z(n19490) );
  NAND U27988 ( .A(n19523), .B(n19524), .Z(n19522) );
  OR U27989 ( .A(n19525), .B(n19526), .Z(n19523) );
  NANDN U27990 ( .A(n19527), .B(n19525), .Z(n19521) );
  IV U27991 ( .A(n19526), .Z(n19527) );
  NAND U27992 ( .A(n19528), .B(n19529), .Z(n19487) );
  NAND U27993 ( .A(n19530), .B(n19531), .Z(n19529) );
  NANDN U27994 ( .A(n19532), .B(n19533), .Z(n19530) );
  NANDN U27995 ( .A(n19533), .B(n19532), .Z(n19528) );
  AND U27996 ( .A(n19534), .B(n19535), .Z(n19489) );
  NAND U27997 ( .A(n19536), .B(n19537), .Z(n19535) );
  OR U27998 ( .A(n19538), .B(n19539), .Z(n19536) );
  NANDN U27999 ( .A(n19540), .B(n19538), .Z(n19534) );
  XNOR U28000 ( .A(n19515), .B(n19541), .Z(N63661) );
  XOR U28001 ( .A(n19517), .B(n19518), .Z(n19541) );
  XNOR U28002 ( .A(n19531), .B(n19542), .Z(n19518) );
  XOR U28003 ( .A(n19532), .B(n19533), .Z(n19542) );
  XOR U28004 ( .A(n19538), .B(n19543), .Z(n19533) );
  XOR U28005 ( .A(n19537), .B(n19540), .Z(n19543) );
  IV U28006 ( .A(n19539), .Z(n19540) );
  NAND U28007 ( .A(n19544), .B(n19545), .Z(n19539) );
  OR U28008 ( .A(n19546), .B(n19547), .Z(n19545) );
  OR U28009 ( .A(n19548), .B(n19549), .Z(n19544) );
  NAND U28010 ( .A(n19550), .B(n19551), .Z(n19537) );
  OR U28011 ( .A(n19552), .B(n19553), .Z(n19551) );
  OR U28012 ( .A(n19554), .B(n19555), .Z(n19550) );
  NOR U28013 ( .A(n19556), .B(n19557), .Z(n19538) );
  ANDN U28014 ( .B(n19558), .A(n19559), .Z(n19532) );
  XNOR U28015 ( .A(n19525), .B(n19560), .Z(n19531) );
  XNOR U28016 ( .A(n19524), .B(n19526), .Z(n19560) );
  NAND U28017 ( .A(n19561), .B(n19562), .Z(n19526) );
  OR U28018 ( .A(n19563), .B(n19564), .Z(n19562) );
  OR U28019 ( .A(n19565), .B(n19566), .Z(n19561) );
  NAND U28020 ( .A(n19567), .B(n19568), .Z(n19524) );
  OR U28021 ( .A(n19569), .B(n19570), .Z(n19568) );
  OR U28022 ( .A(n19571), .B(n19572), .Z(n19567) );
  ANDN U28023 ( .B(n19573), .A(n19574), .Z(n19525) );
  IV U28024 ( .A(n19575), .Z(n19573) );
  ANDN U28025 ( .B(n19576), .A(n19577), .Z(n19517) );
  XOR U28026 ( .A(n19503), .B(n19578), .Z(n19515) );
  XOR U28027 ( .A(n19504), .B(n19505), .Z(n19578) );
  XOR U28028 ( .A(n19510), .B(n19579), .Z(n19505) );
  XOR U28029 ( .A(n19509), .B(n19512), .Z(n19579) );
  IV U28030 ( .A(n19511), .Z(n19512) );
  NAND U28031 ( .A(n19580), .B(n19581), .Z(n19511) );
  OR U28032 ( .A(n19582), .B(n19583), .Z(n19581) );
  OR U28033 ( .A(n19584), .B(n19585), .Z(n19580) );
  NAND U28034 ( .A(n19586), .B(n19587), .Z(n19509) );
  OR U28035 ( .A(n19588), .B(n19589), .Z(n19587) );
  OR U28036 ( .A(n19590), .B(n19591), .Z(n19586) );
  NOR U28037 ( .A(n19592), .B(n19593), .Z(n19510) );
  ANDN U28038 ( .B(n19594), .A(n19595), .Z(n19504) );
  IV U28039 ( .A(n19596), .Z(n19594) );
  XNOR U28040 ( .A(n19497), .B(n19597), .Z(n19503) );
  XNOR U28041 ( .A(n19496), .B(n19498), .Z(n19597) );
  NAND U28042 ( .A(n19598), .B(n19599), .Z(n19498) );
  OR U28043 ( .A(n19600), .B(n19601), .Z(n19599) );
  OR U28044 ( .A(n19602), .B(n19603), .Z(n19598) );
  NAND U28045 ( .A(n19604), .B(n19605), .Z(n19496) );
  OR U28046 ( .A(n19606), .B(n19607), .Z(n19605) );
  OR U28047 ( .A(n19608), .B(n19609), .Z(n19604) );
  ANDN U28048 ( .B(n19610), .A(n19611), .Z(n19497) );
  IV U28049 ( .A(n19612), .Z(n19610) );
  XNOR U28050 ( .A(n19577), .B(n19576), .Z(N63660) );
  XOR U28051 ( .A(n19596), .B(n19595), .Z(n19576) );
  XNOR U28052 ( .A(n19611), .B(n19612), .Z(n19595) );
  XNOR U28053 ( .A(n19606), .B(n19607), .Z(n19612) );
  XNOR U28054 ( .A(n19608), .B(n19609), .Z(n19607) );
  XNOR U28055 ( .A(y[5677]), .B(x[5677]), .Z(n19609) );
  XNOR U28056 ( .A(y[5678]), .B(x[5678]), .Z(n19608) );
  XNOR U28057 ( .A(y[5676]), .B(x[5676]), .Z(n19606) );
  XNOR U28058 ( .A(n19600), .B(n19601), .Z(n19611) );
  XNOR U28059 ( .A(y[5673]), .B(x[5673]), .Z(n19601) );
  XNOR U28060 ( .A(n19602), .B(n19603), .Z(n19600) );
  XNOR U28061 ( .A(y[5674]), .B(x[5674]), .Z(n19603) );
  XNOR U28062 ( .A(y[5675]), .B(x[5675]), .Z(n19602) );
  XNOR U28063 ( .A(n19593), .B(n19592), .Z(n19596) );
  XNOR U28064 ( .A(n19588), .B(n19589), .Z(n19592) );
  XNOR U28065 ( .A(y[5670]), .B(x[5670]), .Z(n19589) );
  XNOR U28066 ( .A(n19590), .B(n19591), .Z(n19588) );
  XNOR U28067 ( .A(y[5671]), .B(x[5671]), .Z(n19591) );
  XNOR U28068 ( .A(y[5672]), .B(x[5672]), .Z(n19590) );
  XNOR U28069 ( .A(n19582), .B(n19583), .Z(n19593) );
  XNOR U28070 ( .A(y[5667]), .B(x[5667]), .Z(n19583) );
  XNOR U28071 ( .A(n19584), .B(n19585), .Z(n19582) );
  XNOR U28072 ( .A(y[5668]), .B(x[5668]), .Z(n19585) );
  XNOR U28073 ( .A(y[5669]), .B(x[5669]), .Z(n19584) );
  XOR U28074 ( .A(n19558), .B(n19559), .Z(n19577) );
  XNOR U28075 ( .A(n19574), .B(n19575), .Z(n19559) );
  XNOR U28076 ( .A(n19569), .B(n19570), .Z(n19575) );
  XNOR U28077 ( .A(n19571), .B(n19572), .Z(n19570) );
  XNOR U28078 ( .A(y[5665]), .B(x[5665]), .Z(n19572) );
  XNOR U28079 ( .A(y[5666]), .B(x[5666]), .Z(n19571) );
  XNOR U28080 ( .A(y[5664]), .B(x[5664]), .Z(n19569) );
  XNOR U28081 ( .A(n19563), .B(n19564), .Z(n19574) );
  XNOR U28082 ( .A(y[5661]), .B(x[5661]), .Z(n19564) );
  XNOR U28083 ( .A(n19565), .B(n19566), .Z(n19563) );
  XNOR U28084 ( .A(y[5662]), .B(x[5662]), .Z(n19566) );
  XNOR U28085 ( .A(y[5663]), .B(x[5663]), .Z(n19565) );
  XOR U28086 ( .A(n19557), .B(n19556), .Z(n19558) );
  XNOR U28087 ( .A(n19552), .B(n19553), .Z(n19556) );
  XNOR U28088 ( .A(y[5658]), .B(x[5658]), .Z(n19553) );
  XNOR U28089 ( .A(n19554), .B(n19555), .Z(n19552) );
  XNOR U28090 ( .A(y[5659]), .B(x[5659]), .Z(n19555) );
  XNOR U28091 ( .A(y[5660]), .B(x[5660]), .Z(n19554) );
  XNOR U28092 ( .A(n19546), .B(n19547), .Z(n19557) );
  XNOR U28093 ( .A(y[5655]), .B(x[5655]), .Z(n19547) );
  XNOR U28094 ( .A(n19548), .B(n19549), .Z(n19546) );
  XNOR U28095 ( .A(y[5656]), .B(x[5656]), .Z(n19549) );
  XNOR U28096 ( .A(y[5657]), .B(x[5657]), .Z(n19548) );
  NAND U28097 ( .A(n19613), .B(n19614), .Z(N63651) );
  NANDN U28098 ( .A(n19615), .B(n19616), .Z(n19614) );
  OR U28099 ( .A(n19617), .B(n19618), .Z(n19616) );
  NAND U28100 ( .A(n19617), .B(n19618), .Z(n19613) );
  XOR U28101 ( .A(n19617), .B(n19619), .Z(N63650) );
  XNOR U28102 ( .A(n19615), .B(n19618), .Z(n19619) );
  AND U28103 ( .A(n19620), .B(n19621), .Z(n19618) );
  NANDN U28104 ( .A(n19622), .B(n19623), .Z(n19621) );
  NANDN U28105 ( .A(n19624), .B(n19625), .Z(n19623) );
  NANDN U28106 ( .A(n19625), .B(n19624), .Z(n19620) );
  NAND U28107 ( .A(n19626), .B(n19627), .Z(n19615) );
  NANDN U28108 ( .A(n19628), .B(n19629), .Z(n19627) );
  OR U28109 ( .A(n19630), .B(n19631), .Z(n19629) );
  NAND U28110 ( .A(n19631), .B(n19630), .Z(n19626) );
  AND U28111 ( .A(n19632), .B(n19633), .Z(n19617) );
  NANDN U28112 ( .A(n19634), .B(n19635), .Z(n19633) );
  NANDN U28113 ( .A(n19636), .B(n19637), .Z(n19635) );
  NANDN U28114 ( .A(n19637), .B(n19636), .Z(n19632) );
  XOR U28115 ( .A(n19631), .B(n19638), .Z(N63649) );
  XOR U28116 ( .A(n19628), .B(n19630), .Z(n19638) );
  XNOR U28117 ( .A(n19624), .B(n19639), .Z(n19630) );
  XNOR U28118 ( .A(n19622), .B(n19625), .Z(n19639) );
  NAND U28119 ( .A(n19640), .B(n19641), .Z(n19625) );
  NAND U28120 ( .A(n19642), .B(n19643), .Z(n19641) );
  OR U28121 ( .A(n19644), .B(n19645), .Z(n19642) );
  NANDN U28122 ( .A(n19646), .B(n19644), .Z(n19640) );
  IV U28123 ( .A(n19645), .Z(n19646) );
  NAND U28124 ( .A(n19647), .B(n19648), .Z(n19622) );
  NAND U28125 ( .A(n19649), .B(n19650), .Z(n19648) );
  NANDN U28126 ( .A(n19651), .B(n19652), .Z(n19649) );
  NANDN U28127 ( .A(n19652), .B(n19651), .Z(n19647) );
  AND U28128 ( .A(n19653), .B(n19654), .Z(n19624) );
  NAND U28129 ( .A(n19655), .B(n19656), .Z(n19654) );
  OR U28130 ( .A(n19657), .B(n19658), .Z(n19655) );
  NANDN U28131 ( .A(n19659), .B(n19657), .Z(n19653) );
  NAND U28132 ( .A(n19660), .B(n19661), .Z(n19628) );
  NANDN U28133 ( .A(n19662), .B(n19663), .Z(n19661) );
  OR U28134 ( .A(n19664), .B(n19665), .Z(n19663) );
  NANDN U28135 ( .A(n19666), .B(n19664), .Z(n19660) );
  IV U28136 ( .A(n19665), .Z(n19666) );
  XNOR U28137 ( .A(n19636), .B(n19667), .Z(n19631) );
  XNOR U28138 ( .A(n19634), .B(n19637), .Z(n19667) );
  NAND U28139 ( .A(n19668), .B(n19669), .Z(n19637) );
  NAND U28140 ( .A(n19670), .B(n19671), .Z(n19669) );
  OR U28141 ( .A(n19672), .B(n19673), .Z(n19670) );
  NANDN U28142 ( .A(n19674), .B(n19672), .Z(n19668) );
  IV U28143 ( .A(n19673), .Z(n19674) );
  NAND U28144 ( .A(n19675), .B(n19676), .Z(n19634) );
  NAND U28145 ( .A(n19677), .B(n19678), .Z(n19676) );
  NANDN U28146 ( .A(n19679), .B(n19680), .Z(n19677) );
  NANDN U28147 ( .A(n19680), .B(n19679), .Z(n19675) );
  AND U28148 ( .A(n19681), .B(n19682), .Z(n19636) );
  NAND U28149 ( .A(n19683), .B(n19684), .Z(n19682) );
  OR U28150 ( .A(n19685), .B(n19686), .Z(n19683) );
  NANDN U28151 ( .A(n19687), .B(n19685), .Z(n19681) );
  XNOR U28152 ( .A(n19662), .B(n19688), .Z(N63648) );
  XOR U28153 ( .A(n19664), .B(n19665), .Z(n19688) );
  XNOR U28154 ( .A(n19678), .B(n19689), .Z(n19665) );
  XOR U28155 ( .A(n19679), .B(n19680), .Z(n19689) );
  XOR U28156 ( .A(n19685), .B(n19690), .Z(n19680) );
  XOR U28157 ( .A(n19684), .B(n19687), .Z(n19690) );
  IV U28158 ( .A(n19686), .Z(n19687) );
  NAND U28159 ( .A(n19691), .B(n19692), .Z(n19686) );
  OR U28160 ( .A(n19693), .B(n19694), .Z(n19692) );
  OR U28161 ( .A(n19695), .B(n19696), .Z(n19691) );
  NAND U28162 ( .A(n19697), .B(n19698), .Z(n19684) );
  OR U28163 ( .A(n19699), .B(n19700), .Z(n19698) );
  OR U28164 ( .A(n19701), .B(n19702), .Z(n19697) );
  NOR U28165 ( .A(n19703), .B(n19704), .Z(n19685) );
  ANDN U28166 ( .B(n19705), .A(n19706), .Z(n19679) );
  XNOR U28167 ( .A(n19672), .B(n19707), .Z(n19678) );
  XNOR U28168 ( .A(n19671), .B(n19673), .Z(n19707) );
  NAND U28169 ( .A(n19708), .B(n19709), .Z(n19673) );
  OR U28170 ( .A(n19710), .B(n19711), .Z(n19709) );
  OR U28171 ( .A(n19712), .B(n19713), .Z(n19708) );
  NAND U28172 ( .A(n19714), .B(n19715), .Z(n19671) );
  OR U28173 ( .A(n19716), .B(n19717), .Z(n19715) );
  OR U28174 ( .A(n19718), .B(n19719), .Z(n19714) );
  ANDN U28175 ( .B(n19720), .A(n19721), .Z(n19672) );
  IV U28176 ( .A(n19722), .Z(n19720) );
  ANDN U28177 ( .B(n19723), .A(n19724), .Z(n19664) );
  XOR U28178 ( .A(n19650), .B(n19725), .Z(n19662) );
  XOR U28179 ( .A(n19651), .B(n19652), .Z(n19725) );
  XOR U28180 ( .A(n19657), .B(n19726), .Z(n19652) );
  XOR U28181 ( .A(n19656), .B(n19659), .Z(n19726) );
  IV U28182 ( .A(n19658), .Z(n19659) );
  NAND U28183 ( .A(n19727), .B(n19728), .Z(n19658) );
  OR U28184 ( .A(n19729), .B(n19730), .Z(n19728) );
  OR U28185 ( .A(n19731), .B(n19732), .Z(n19727) );
  NAND U28186 ( .A(n19733), .B(n19734), .Z(n19656) );
  OR U28187 ( .A(n19735), .B(n19736), .Z(n19734) );
  OR U28188 ( .A(n19737), .B(n19738), .Z(n19733) );
  NOR U28189 ( .A(n19739), .B(n19740), .Z(n19657) );
  ANDN U28190 ( .B(n19741), .A(n19742), .Z(n19651) );
  IV U28191 ( .A(n19743), .Z(n19741) );
  XNOR U28192 ( .A(n19644), .B(n19744), .Z(n19650) );
  XNOR U28193 ( .A(n19643), .B(n19645), .Z(n19744) );
  NAND U28194 ( .A(n19745), .B(n19746), .Z(n19645) );
  OR U28195 ( .A(n19747), .B(n19748), .Z(n19746) );
  OR U28196 ( .A(n19749), .B(n19750), .Z(n19745) );
  NAND U28197 ( .A(n19751), .B(n19752), .Z(n19643) );
  OR U28198 ( .A(n19753), .B(n19754), .Z(n19752) );
  OR U28199 ( .A(n19755), .B(n19756), .Z(n19751) );
  ANDN U28200 ( .B(n19757), .A(n19758), .Z(n19644) );
  IV U28201 ( .A(n19759), .Z(n19757) );
  XNOR U28202 ( .A(n19724), .B(n19723), .Z(N63647) );
  XOR U28203 ( .A(n19743), .B(n19742), .Z(n19723) );
  XNOR U28204 ( .A(n19758), .B(n19759), .Z(n19742) );
  XNOR U28205 ( .A(n19753), .B(n19754), .Z(n19759) );
  XNOR U28206 ( .A(n19755), .B(n19756), .Z(n19754) );
  XNOR U28207 ( .A(y[5653]), .B(x[5653]), .Z(n19756) );
  XNOR U28208 ( .A(y[5654]), .B(x[5654]), .Z(n19755) );
  XNOR U28209 ( .A(y[5652]), .B(x[5652]), .Z(n19753) );
  XNOR U28210 ( .A(n19747), .B(n19748), .Z(n19758) );
  XNOR U28211 ( .A(y[5649]), .B(x[5649]), .Z(n19748) );
  XNOR U28212 ( .A(n19749), .B(n19750), .Z(n19747) );
  XNOR U28213 ( .A(y[5650]), .B(x[5650]), .Z(n19750) );
  XNOR U28214 ( .A(y[5651]), .B(x[5651]), .Z(n19749) );
  XNOR U28215 ( .A(n19740), .B(n19739), .Z(n19743) );
  XNOR U28216 ( .A(n19735), .B(n19736), .Z(n19739) );
  XNOR U28217 ( .A(y[5646]), .B(x[5646]), .Z(n19736) );
  XNOR U28218 ( .A(n19737), .B(n19738), .Z(n19735) );
  XNOR U28219 ( .A(y[5647]), .B(x[5647]), .Z(n19738) );
  XNOR U28220 ( .A(y[5648]), .B(x[5648]), .Z(n19737) );
  XNOR U28221 ( .A(n19729), .B(n19730), .Z(n19740) );
  XNOR U28222 ( .A(y[5643]), .B(x[5643]), .Z(n19730) );
  XNOR U28223 ( .A(n19731), .B(n19732), .Z(n19729) );
  XNOR U28224 ( .A(y[5644]), .B(x[5644]), .Z(n19732) );
  XNOR U28225 ( .A(y[5645]), .B(x[5645]), .Z(n19731) );
  XOR U28226 ( .A(n19705), .B(n19706), .Z(n19724) );
  XNOR U28227 ( .A(n19721), .B(n19722), .Z(n19706) );
  XNOR U28228 ( .A(n19716), .B(n19717), .Z(n19722) );
  XNOR U28229 ( .A(n19718), .B(n19719), .Z(n19717) );
  XNOR U28230 ( .A(y[5641]), .B(x[5641]), .Z(n19719) );
  XNOR U28231 ( .A(y[5642]), .B(x[5642]), .Z(n19718) );
  XNOR U28232 ( .A(y[5640]), .B(x[5640]), .Z(n19716) );
  XNOR U28233 ( .A(n19710), .B(n19711), .Z(n19721) );
  XNOR U28234 ( .A(y[5637]), .B(x[5637]), .Z(n19711) );
  XNOR U28235 ( .A(n19712), .B(n19713), .Z(n19710) );
  XNOR U28236 ( .A(y[5638]), .B(x[5638]), .Z(n19713) );
  XNOR U28237 ( .A(y[5639]), .B(x[5639]), .Z(n19712) );
  XOR U28238 ( .A(n19704), .B(n19703), .Z(n19705) );
  XNOR U28239 ( .A(n19699), .B(n19700), .Z(n19703) );
  XNOR U28240 ( .A(y[5634]), .B(x[5634]), .Z(n19700) );
  XNOR U28241 ( .A(n19701), .B(n19702), .Z(n19699) );
  XNOR U28242 ( .A(y[5635]), .B(x[5635]), .Z(n19702) );
  XNOR U28243 ( .A(y[5636]), .B(x[5636]), .Z(n19701) );
  XNOR U28244 ( .A(n19693), .B(n19694), .Z(n19704) );
  XNOR U28245 ( .A(y[5631]), .B(x[5631]), .Z(n19694) );
  XNOR U28246 ( .A(n19695), .B(n19696), .Z(n19693) );
  XNOR U28247 ( .A(y[5632]), .B(x[5632]), .Z(n19696) );
  XNOR U28248 ( .A(y[5633]), .B(x[5633]), .Z(n19695) );
  NAND U28249 ( .A(n19760), .B(n19761), .Z(N63638) );
  NANDN U28250 ( .A(n19762), .B(n19763), .Z(n19761) );
  OR U28251 ( .A(n19764), .B(n19765), .Z(n19763) );
  NAND U28252 ( .A(n19764), .B(n19765), .Z(n19760) );
  XOR U28253 ( .A(n19764), .B(n19766), .Z(N63637) );
  XNOR U28254 ( .A(n19762), .B(n19765), .Z(n19766) );
  AND U28255 ( .A(n19767), .B(n19768), .Z(n19765) );
  NANDN U28256 ( .A(n19769), .B(n19770), .Z(n19768) );
  NANDN U28257 ( .A(n19771), .B(n19772), .Z(n19770) );
  NANDN U28258 ( .A(n19772), .B(n19771), .Z(n19767) );
  NAND U28259 ( .A(n19773), .B(n19774), .Z(n19762) );
  NANDN U28260 ( .A(n19775), .B(n19776), .Z(n19774) );
  OR U28261 ( .A(n19777), .B(n19778), .Z(n19776) );
  NAND U28262 ( .A(n19778), .B(n19777), .Z(n19773) );
  AND U28263 ( .A(n19779), .B(n19780), .Z(n19764) );
  NANDN U28264 ( .A(n19781), .B(n19782), .Z(n19780) );
  NANDN U28265 ( .A(n19783), .B(n19784), .Z(n19782) );
  NANDN U28266 ( .A(n19784), .B(n19783), .Z(n19779) );
  XOR U28267 ( .A(n19778), .B(n19785), .Z(N63636) );
  XOR U28268 ( .A(n19775), .B(n19777), .Z(n19785) );
  XNOR U28269 ( .A(n19771), .B(n19786), .Z(n19777) );
  XNOR U28270 ( .A(n19769), .B(n19772), .Z(n19786) );
  NAND U28271 ( .A(n19787), .B(n19788), .Z(n19772) );
  NAND U28272 ( .A(n19789), .B(n19790), .Z(n19788) );
  OR U28273 ( .A(n19791), .B(n19792), .Z(n19789) );
  NANDN U28274 ( .A(n19793), .B(n19791), .Z(n19787) );
  IV U28275 ( .A(n19792), .Z(n19793) );
  NAND U28276 ( .A(n19794), .B(n19795), .Z(n19769) );
  NAND U28277 ( .A(n19796), .B(n19797), .Z(n19795) );
  NANDN U28278 ( .A(n19798), .B(n19799), .Z(n19796) );
  NANDN U28279 ( .A(n19799), .B(n19798), .Z(n19794) );
  AND U28280 ( .A(n19800), .B(n19801), .Z(n19771) );
  NAND U28281 ( .A(n19802), .B(n19803), .Z(n19801) );
  OR U28282 ( .A(n19804), .B(n19805), .Z(n19802) );
  NANDN U28283 ( .A(n19806), .B(n19804), .Z(n19800) );
  NAND U28284 ( .A(n19807), .B(n19808), .Z(n19775) );
  NANDN U28285 ( .A(n19809), .B(n19810), .Z(n19808) );
  OR U28286 ( .A(n19811), .B(n19812), .Z(n19810) );
  NANDN U28287 ( .A(n19813), .B(n19811), .Z(n19807) );
  IV U28288 ( .A(n19812), .Z(n19813) );
  XNOR U28289 ( .A(n19783), .B(n19814), .Z(n19778) );
  XNOR U28290 ( .A(n19781), .B(n19784), .Z(n19814) );
  NAND U28291 ( .A(n19815), .B(n19816), .Z(n19784) );
  NAND U28292 ( .A(n19817), .B(n19818), .Z(n19816) );
  OR U28293 ( .A(n19819), .B(n19820), .Z(n19817) );
  NANDN U28294 ( .A(n19821), .B(n19819), .Z(n19815) );
  IV U28295 ( .A(n19820), .Z(n19821) );
  NAND U28296 ( .A(n19822), .B(n19823), .Z(n19781) );
  NAND U28297 ( .A(n19824), .B(n19825), .Z(n19823) );
  NANDN U28298 ( .A(n19826), .B(n19827), .Z(n19824) );
  NANDN U28299 ( .A(n19827), .B(n19826), .Z(n19822) );
  AND U28300 ( .A(n19828), .B(n19829), .Z(n19783) );
  NAND U28301 ( .A(n19830), .B(n19831), .Z(n19829) );
  OR U28302 ( .A(n19832), .B(n19833), .Z(n19830) );
  NANDN U28303 ( .A(n19834), .B(n19832), .Z(n19828) );
  XNOR U28304 ( .A(n19809), .B(n19835), .Z(N63635) );
  XOR U28305 ( .A(n19811), .B(n19812), .Z(n19835) );
  XNOR U28306 ( .A(n19825), .B(n19836), .Z(n19812) );
  XOR U28307 ( .A(n19826), .B(n19827), .Z(n19836) );
  XOR U28308 ( .A(n19832), .B(n19837), .Z(n19827) );
  XOR U28309 ( .A(n19831), .B(n19834), .Z(n19837) );
  IV U28310 ( .A(n19833), .Z(n19834) );
  NAND U28311 ( .A(n19838), .B(n19839), .Z(n19833) );
  OR U28312 ( .A(n19840), .B(n19841), .Z(n19839) );
  OR U28313 ( .A(n19842), .B(n19843), .Z(n19838) );
  NAND U28314 ( .A(n19844), .B(n19845), .Z(n19831) );
  OR U28315 ( .A(n19846), .B(n19847), .Z(n19845) );
  OR U28316 ( .A(n19848), .B(n19849), .Z(n19844) );
  NOR U28317 ( .A(n19850), .B(n19851), .Z(n19832) );
  ANDN U28318 ( .B(n19852), .A(n19853), .Z(n19826) );
  XNOR U28319 ( .A(n19819), .B(n19854), .Z(n19825) );
  XNOR U28320 ( .A(n19818), .B(n19820), .Z(n19854) );
  NAND U28321 ( .A(n19855), .B(n19856), .Z(n19820) );
  OR U28322 ( .A(n19857), .B(n19858), .Z(n19856) );
  OR U28323 ( .A(n19859), .B(n19860), .Z(n19855) );
  NAND U28324 ( .A(n19861), .B(n19862), .Z(n19818) );
  OR U28325 ( .A(n19863), .B(n19864), .Z(n19862) );
  OR U28326 ( .A(n19865), .B(n19866), .Z(n19861) );
  ANDN U28327 ( .B(n19867), .A(n19868), .Z(n19819) );
  IV U28328 ( .A(n19869), .Z(n19867) );
  ANDN U28329 ( .B(n19870), .A(n19871), .Z(n19811) );
  XOR U28330 ( .A(n19797), .B(n19872), .Z(n19809) );
  XOR U28331 ( .A(n19798), .B(n19799), .Z(n19872) );
  XOR U28332 ( .A(n19804), .B(n19873), .Z(n19799) );
  XOR U28333 ( .A(n19803), .B(n19806), .Z(n19873) );
  IV U28334 ( .A(n19805), .Z(n19806) );
  NAND U28335 ( .A(n19874), .B(n19875), .Z(n19805) );
  OR U28336 ( .A(n19876), .B(n19877), .Z(n19875) );
  OR U28337 ( .A(n19878), .B(n19879), .Z(n19874) );
  NAND U28338 ( .A(n19880), .B(n19881), .Z(n19803) );
  OR U28339 ( .A(n19882), .B(n19883), .Z(n19881) );
  OR U28340 ( .A(n19884), .B(n19885), .Z(n19880) );
  NOR U28341 ( .A(n19886), .B(n19887), .Z(n19804) );
  ANDN U28342 ( .B(n19888), .A(n19889), .Z(n19798) );
  IV U28343 ( .A(n19890), .Z(n19888) );
  XNOR U28344 ( .A(n19791), .B(n19891), .Z(n19797) );
  XNOR U28345 ( .A(n19790), .B(n19792), .Z(n19891) );
  NAND U28346 ( .A(n19892), .B(n19893), .Z(n19792) );
  OR U28347 ( .A(n19894), .B(n19895), .Z(n19893) );
  OR U28348 ( .A(n19896), .B(n19897), .Z(n19892) );
  NAND U28349 ( .A(n19898), .B(n19899), .Z(n19790) );
  OR U28350 ( .A(n19900), .B(n19901), .Z(n19899) );
  OR U28351 ( .A(n19902), .B(n19903), .Z(n19898) );
  ANDN U28352 ( .B(n19904), .A(n19905), .Z(n19791) );
  IV U28353 ( .A(n19906), .Z(n19904) );
  XNOR U28354 ( .A(n19871), .B(n19870), .Z(N63634) );
  XOR U28355 ( .A(n19890), .B(n19889), .Z(n19870) );
  XNOR U28356 ( .A(n19905), .B(n19906), .Z(n19889) );
  XNOR U28357 ( .A(n19900), .B(n19901), .Z(n19906) );
  XNOR U28358 ( .A(n19902), .B(n19903), .Z(n19901) );
  XNOR U28359 ( .A(y[5629]), .B(x[5629]), .Z(n19903) );
  XNOR U28360 ( .A(y[5630]), .B(x[5630]), .Z(n19902) );
  XNOR U28361 ( .A(y[5628]), .B(x[5628]), .Z(n19900) );
  XNOR U28362 ( .A(n19894), .B(n19895), .Z(n19905) );
  XNOR U28363 ( .A(y[5625]), .B(x[5625]), .Z(n19895) );
  XNOR U28364 ( .A(n19896), .B(n19897), .Z(n19894) );
  XNOR U28365 ( .A(y[5626]), .B(x[5626]), .Z(n19897) );
  XNOR U28366 ( .A(y[5627]), .B(x[5627]), .Z(n19896) );
  XNOR U28367 ( .A(n19887), .B(n19886), .Z(n19890) );
  XNOR U28368 ( .A(n19882), .B(n19883), .Z(n19886) );
  XNOR U28369 ( .A(y[5622]), .B(x[5622]), .Z(n19883) );
  XNOR U28370 ( .A(n19884), .B(n19885), .Z(n19882) );
  XNOR U28371 ( .A(y[5623]), .B(x[5623]), .Z(n19885) );
  XNOR U28372 ( .A(y[5624]), .B(x[5624]), .Z(n19884) );
  XNOR U28373 ( .A(n19876), .B(n19877), .Z(n19887) );
  XNOR U28374 ( .A(y[5619]), .B(x[5619]), .Z(n19877) );
  XNOR U28375 ( .A(n19878), .B(n19879), .Z(n19876) );
  XNOR U28376 ( .A(y[5620]), .B(x[5620]), .Z(n19879) );
  XNOR U28377 ( .A(y[5621]), .B(x[5621]), .Z(n19878) );
  XOR U28378 ( .A(n19852), .B(n19853), .Z(n19871) );
  XNOR U28379 ( .A(n19868), .B(n19869), .Z(n19853) );
  XNOR U28380 ( .A(n19863), .B(n19864), .Z(n19869) );
  XNOR U28381 ( .A(n19865), .B(n19866), .Z(n19864) );
  XNOR U28382 ( .A(y[5617]), .B(x[5617]), .Z(n19866) );
  XNOR U28383 ( .A(y[5618]), .B(x[5618]), .Z(n19865) );
  XNOR U28384 ( .A(y[5616]), .B(x[5616]), .Z(n19863) );
  XNOR U28385 ( .A(n19857), .B(n19858), .Z(n19868) );
  XNOR U28386 ( .A(y[5613]), .B(x[5613]), .Z(n19858) );
  XNOR U28387 ( .A(n19859), .B(n19860), .Z(n19857) );
  XNOR U28388 ( .A(y[5614]), .B(x[5614]), .Z(n19860) );
  XNOR U28389 ( .A(y[5615]), .B(x[5615]), .Z(n19859) );
  XOR U28390 ( .A(n19851), .B(n19850), .Z(n19852) );
  XNOR U28391 ( .A(n19846), .B(n19847), .Z(n19850) );
  XNOR U28392 ( .A(y[5610]), .B(x[5610]), .Z(n19847) );
  XNOR U28393 ( .A(n19848), .B(n19849), .Z(n19846) );
  XNOR U28394 ( .A(y[5611]), .B(x[5611]), .Z(n19849) );
  XNOR U28395 ( .A(y[5612]), .B(x[5612]), .Z(n19848) );
  XNOR U28396 ( .A(n19840), .B(n19841), .Z(n19851) );
  XNOR U28397 ( .A(y[5607]), .B(x[5607]), .Z(n19841) );
  XNOR U28398 ( .A(n19842), .B(n19843), .Z(n19840) );
  XNOR U28399 ( .A(y[5608]), .B(x[5608]), .Z(n19843) );
  XNOR U28400 ( .A(y[5609]), .B(x[5609]), .Z(n19842) );
  NAND U28401 ( .A(n19907), .B(n19908), .Z(N63625) );
  NANDN U28402 ( .A(n19909), .B(n19910), .Z(n19908) );
  OR U28403 ( .A(n19911), .B(n19912), .Z(n19910) );
  NAND U28404 ( .A(n19911), .B(n19912), .Z(n19907) );
  XOR U28405 ( .A(n19911), .B(n19913), .Z(N63624) );
  XNOR U28406 ( .A(n19909), .B(n19912), .Z(n19913) );
  AND U28407 ( .A(n19914), .B(n19915), .Z(n19912) );
  NANDN U28408 ( .A(n19916), .B(n19917), .Z(n19915) );
  NANDN U28409 ( .A(n19918), .B(n19919), .Z(n19917) );
  NANDN U28410 ( .A(n19919), .B(n19918), .Z(n19914) );
  NAND U28411 ( .A(n19920), .B(n19921), .Z(n19909) );
  NANDN U28412 ( .A(n19922), .B(n19923), .Z(n19921) );
  OR U28413 ( .A(n19924), .B(n19925), .Z(n19923) );
  NAND U28414 ( .A(n19925), .B(n19924), .Z(n19920) );
  AND U28415 ( .A(n19926), .B(n19927), .Z(n19911) );
  NANDN U28416 ( .A(n19928), .B(n19929), .Z(n19927) );
  NANDN U28417 ( .A(n19930), .B(n19931), .Z(n19929) );
  NANDN U28418 ( .A(n19931), .B(n19930), .Z(n19926) );
  XOR U28419 ( .A(n19925), .B(n19932), .Z(N63623) );
  XOR U28420 ( .A(n19922), .B(n19924), .Z(n19932) );
  XNOR U28421 ( .A(n19918), .B(n19933), .Z(n19924) );
  XNOR U28422 ( .A(n19916), .B(n19919), .Z(n19933) );
  NAND U28423 ( .A(n19934), .B(n19935), .Z(n19919) );
  NAND U28424 ( .A(n19936), .B(n19937), .Z(n19935) );
  OR U28425 ( .A(n19938), .B(n19939), .Z(n19936) );
  NANDN U28426 ( .A(n19940), .B(n19938), .Z(n19934) );
  IV U28427 ( .A(n19939), .Z(n19940) );
  NAND U28428 ( .A(n19941), .B(n19942), .Z(n19916) );
  NAND U28429 ( .A(n19943), .B(n19944), .Z(n19942) );
  NANDN U28430 ( .A(n19945), .B(n19946), .Z(n19943) );
  NANDN U28431 ( .A(n19946), .B(n19945), .Z(n19941) );
  AND U28432 ( .A(n19947), .B(n19948), .Z(n19918) );
  NAND U28433 ( .A(n19949), .B(n19950), .Z(n19948) );
  OR U28434 ( .A(n19951), .B(n19952), .Z(n19949) );
  NANDN U28435 ( .A(n19953), .B(n19951), .Z(n19947) );
  NAND U28436 ( .A(n19954), .B(n19955), .Z(n19922) );
  NANDN U28437 ( .A(n19956), .B(n19957), .Z(n19955) );
  OR U28438 ( .A(n19958), .B(n19959), .Z(n19957) );
  NANDN U28439 ( .A(n19960), .B(n19958), .Z(n19954) );
  IV U28440 ( .A(n19959), .Z(n19960) );
  XNOR U28441 ( .A(n19930), .B(n19961), .Z(n19925) );
  XNOR U28442 ( .A(n19928), .B(n19931), .Z(n19961) );
  NAND U28443 ( .A(n19962), .B(n19963), .Z(n19931) );
  NAND U28444 ( .A(n19964), .B(n19965), .Z(n19963) );
  OR U28445 ( .A(n19966), .B(n19967), .Z(n19964) );
  NANDN U28446 ( .A(n19968), .B(n19966), .Z(n19962) );
  IV U28447 ( .A(n19967), .Z(n19968) );
  NAND U28448 ( .A(n19969), .B(n19970), .Z(n19928) );
  NAND U28449 ( .A(n19971), .B(n19972), .Z(n19970) );
  NANDN U28450 ( .A(n19973), .B(n19974), .Z(n19971) );
  NANDN U28451 ( .A(n19974), .B(n19973), .Z(n19969) );
  AND U28452 ( .A(n19975), .B(n19976), .Z(n19930) );
  NAND U28453 ( .A(n19977), .B(n19978), .Z(n19976) );
  OR U28454 ( .A(n19979), .B(n19980), .Z(n19977) );
  NANDN U28455 ( .A(n19981), .B(n19979), .Z(n19975) );
  XNOR U28456 ( .A(n19956), .B(n19982), .Z(N63622) );
  XOR U28457 ( .A(n19958), .B(n19959), .Z(n19982) );
  XNOR U28458 ( .A(n19972), .B(n19983), .Z(n19959) );
  XOR U28459 ( .A(n19973), .B(n19974), .Z(n19983) );
  XOR U28460 ( .A(n19979), .B(n19984), .Z(n19974) );
  XOR U28461 ( .A(n19978), .B(n19981), .Z(n19984) );
  IV U28462 ( .A(n19980), .Z(n19981) );
  NAND U28463 ( .A(n19985), .B(n19986), .Z(n19980) );
  OR U28464 ( .A(n19987), .B(n19988), .Z(n19986) );
  OR U28465 ( .A(n19989), .B(n19990), .Z(n19985) );
  NAND U28466 ( .A(n19991), .B(n19992), .Z(n19978) );
  OR U28467 ( .A(n19993), .B(n19994), .Z(n19992) );
  OR U28468 ( .A(n19995), .B(n19996), .Z(n19991) );
  NOR U28469 ( .A(n19997), .B(n19998), .Z(n19979) );
  ANDN U28470 ( .B(n19999), .A(n20000), .Z(n19973) );
  XNOR U28471 ( .A(n19966), .B(n20001), .Z(n19972) );
  XNOR U28472 ( .A(n19965), .B(n19967), .Z(n20001) );
  NAND U28473 ( .A(n20002), .B(n20003), .Z(n19967) );
  OR U28474 ( .A(n20004), .B(n20005), .Z(n20003) );
  OR U28475 ( .A(n20006), .B(n20007), .Z(n20002) );
  NAND U28476 ( .A(n20008), .B(n20009), .Z(n19965) );
  OR U28477 ( .A(n20010), .B(n20011), .Z(n20009) );
  OR U28478 ( .A(n20012), .B(n20013), .Z(n20008) );
  ANDN U28479 ( .B(n20014), .A(n20015), .Z(n19966) );
  IV U28480 ( .A(n20016), .Z(n20014) );
  ANDN U28481 ( .B(n20017), .A(n20018), .Z(n19958) );
  XOR U28482 ( .A(n19944), .B(n20019), .Z(n19956) );
  XOR U28483 ( .A(n19945), .B(n19946), .Z(n20019) );
  XOR U28484 ( .A(n19951), .B(n20020), .Z(n19946) );
  XOR U28485 ( .A(n19950), .B(n19953), .Z(n20020) );
  IV U28486 ( .A(n19952), .Z(n19953) );
  NAND U28487 ( .A(n20021), .B(n20022), .Z(n19952) );
  OR U28488 ( .A(n20023), .B(n20024), .Z(n20022) );
  OR U28489 ( .A(n20025), .B(n20026), .Z(n20021) );
  NAND U28490 ( .A(n20027), .B(n20028), .Z(n19950) );
  OR U28491 ( .A(n20029), .B(n20030), .Z(n20028) );
  OR U28492 ( .A(n20031), .B(n20032), .Z(n20027) );
  NOR U28493 ( .A(n20033), .B(n20034), .Z(n19951) );
  ANDN U28494 ( .B(n20035), .A(n20036), .Z(n19945) );
  IV U28495 ( .A(n20037), .Z(n20035) );
  XNOR U28496 ( .A(n19938), .B(n20038), .Z(n19944) );
  XNOR U28497 ( .A(n19937), .B(n19939), .Z(n20038) );
  NAND U28498 ( .A(n20039), .B(n20040), .Z(n19939) );
  OR U28499 ( .A(n20041), .B(n20042), .Z(n20040) );
  OR U28500 ( .A(n20043), .B(n20044), .Z(n20039) );
  NAND U28501 ( .A(n20045), .B(n20046), .Z(n19937) );
  OR U28502 ( .A(n20047), .B(n20048), .Z(n20046) );
  OR U28503 ( .A(n20049), .B(n20050), .Z(n20045) );
  ANDN U28504 ( .B(n20051), .A(n20052), .Z(n19938) );
  IV U28505 ( .A(n20053), .Z(n20051) );
  XNOR U28506 ( .A(n20018), .B(n20017), .Z(N63621) );
  XOR U28507 ( .A(n20037), .B(n20036), .Z(n20017) );
  XNOR U28508 ( .A(n20052), .B(n20053), .Z(n20036) );
  XNOR U28509 ( .A(n20047), .B(n20048), .Z(n20053) );
  XNOR U28510 ( .A(n20049), .B(n20050), .Z(n20048) );
  XNOR U28511 ( .A(y[5605]), .B(x[5605]), .Z(n20050) );
  XNOR U28512 ( .A(y[5606]), .B(x[5606]), .Z(n20049) );
  XNOR U28513 ( .A(y[5604]), .B(x[5604]), .Z(n20047) );
  XNOR U28514 ( .A(n20041), .B(n20042), .Z(n20052) );
  XNOR U28515 ( .A(y[5601]), .B(x[5601]), .Z(n20042) );
  XNOR U28516 ( .A(n20043), .B(n20044), .Z(n20041) );
  XNOR U28517 ( .A(y[5602]), .B(x[5602]), .Z(n20044) );
  XNOR U28518 ( .A(y[5603]), .B(x[5603]), .Z(n20043) );
  XNOR U28519 ( .A(n20034), .B(n20033), .Z(n20037) );
  XNOR U28520 ( .A(n20029), .B(n20030), .Z(n20033) );
  XNOR U28521 ( .A(y[5598]), .B(x[5598]), .Z(n20030) );
  XNOR U28522 ( .A(n20031), .B(n20032), .Z(n20029) );
  XNOR U28523 ( .A(y[5599]), .B(x[5599]), .Z(n20032) );
  XNOR U28524 ( .A(y[5600]), .B(x[5600]), .Z(n20031) );
  XNOR U28525 ( .A(n20023), .B(n20024), .Z(n20034) );
  XNOR U28526 ( .A(y[5595]), .B(x[5595]), .Z(n20024) );
  XNOR U28527 ( .A(n20025), .B(n20026), .Z(n20023) );
  XNOR U28528 ( .A(y[5596]), .B(x[5596]), .Z(n20026) );
  XNOR U28529 ( .A(y[5597]), .B(x[5597]), .Z(n20025) );
  XOR U28530 ( .A(n19999), .B(n20000), .Z(n20018) );
  XNOR U28531 ( .A(n20015), .B(n20016), .Z(n20000) );
  XNOR U28532 ( .A(n20010), .B(n20011), .Z(n20016) );
  XNOR U28533 ( .A(n20012), .B(n20013), .Z(n20011) );
  XNOR U28534 ( .A(y[5593]), .B(x[5593]), .Z(n20013) );
  XNOR U28535 ( .A(y[5594]), .B(x[5594]), .Z(n20012) );
  XNOR U28536 ( .A(y[5592]), .B(x[5592]), .Z(n20010) );
  XNOR U28537 ( .A(n20004), .B(n20005), .Z(n20015) );
  XNOR U28538 ( .A(y[5589]), .B(x[5589]), .Z(n20005) );
  XNOR U28539 ( .A(n20006), .B(n20007), .Z(n20004) );
  XNOR U28540 ( .A(y[5590]), .B(x[5590]), .Z(n20007) );
  XNOR U28541 ( .A(y[5591]), .B(x[5591]), .Z(n20006) );
  XOR U28542 ( .A(n19998), .B(n19997), .Z(n19999) );
  XNOR U28543 ( .A(n19993), .B(n19994), .Z(n19997) );
  XNOR U28544 ( .A(y[5586]), .B(x[5586]), .Z(n19994) );
  XNOR U28545 ( .A(n19995), .B(n19996), .Z(n19993) );
  XNOR U28546 ( .A(y[5587]), .B(x[5587]), .Z(n19996) );
  XNOR U28547 ( .A(y[5588]), .B(x[5588]), .Z(n19995) );
  XNOR U28548 ( .A(n19987), .B(n19988), .Z(n19998) );
  XNOR U28549 ( .A(y[5583]), .B(x[5583]), .Z(n19988) );
  XNOR U28550 ( .A(n19989), .B(n19990), .Z(n19987) );
  XNOR U28551 ( .A(y[5584]), .B(x[5584]), .Z(n19990) );
  XNOR U28552 ( .A(y[5585]), .B(x[5585]), .Z(n19989) );
  NAND U28553 ( .A(n20054), .B(n20055), .Z(N63612) );
  NANDN U28554 ( .A(n20056), .B(n20057), .Z(n20055) );
  OR U28555 ( .A(n20058), .B(n20059), .Z(n20057) );
  NAND U28556 ( .A(n20058), .B(n20059), .Z(n20054) );
  XOR U28557 ( .A(n20058), .B(n20060), .Z(N63611) );
  XNOR U28558 ( .A(n20056), .B(n20059), .Z(n20060) );
  AND U28559 ( .A(n20061), .B(n20062), .Z(n20059) );
  NANDN U28560 ( .A(n20063), .B(n20064), .Z(n20062) );
  NANDN U28561 ( .A(n20065), .B(n20066), .Z(n20064) );
  NANDN U28562 ( .A(n20066), .B(n20065), .Z(n20061) );
  NAND U28563 ( .A(n20067), .B(n20068), .Z(n20056) );
  NANDN U28564 ( .A(n20069), .B(n20070), .Z(n20068) );
  OR U28565 ( .A(n20071), .B(n20072), .Z(n20070) );
  NAND U28566 ( .A(n20072), .B(n20071), .Z(n20067) );
  AND U28567 ( .A(n20073), .B(n20074), .Z(n20058) );
  NANDN U28568 ( .A(n20075), .B(n20076), .Z(n20074) );
  NANDN U28569 ( .A(n20077), .B(n20078), .Z(n20076) );
  NANDN U28570 ( .A(n20078), .B(n20077), .Z(n20073) );
  XOR U28571 ( .A(n20072), .B(n20079), .Z(N63610) );
  XOR U28572 ( .A(n20069), .B(n20071), .Z(n20079) );
  XNOR U28573 ( .A(n20065), .B(n20080), .Z(n20071) );
  XNOR U28574 ( .A(n20063), .B(n20066), .Z(n20080) );
  NAND U28575 ( .A(n20081), .B(n20082), .Z(n20066) );
  NAND U28576 ( .A(n20083), .B(n20084), .Z(n20082) );
  OR U28577 ( .A(n20085), .B(n20086), .Z(n20083) );
  NANDN U28578 ( .A(n20087), .B(n20085), .Z(n20081) );
  IV U28579 ( .A(n20086), .Z(n20087) );
  NAND U28580 ( .A(n20088), .B(n20089), .Z(n20063) );
  NAND U28581 ( .A(n20090), .B(n20091), .Z(n20089) );
  NANDN U28582 ( .A(n20092), .B(n20093), .Z(n20090) );
  NANDN U28583 ( .A(n20093), .B(n20092), .Z(n20088) );
  AND U28584 ( .A(n20094), .B(n20095), .Z(n20065) );
  NAND U28585 ( .A(n20096), .B(n20097), .Z(n20095) );
  OR U28586 ( .A(n20098), .B(n20099), .Z(n20096) );
  NANDN U28587 ( .A(n20100), .B(n20098), .Z(n20094) );
  NAND U28588 ( .A(n20101), .B(n20102), .Z(n20069) );
  NANDN U28589 ( .A(n20103), .B(n20104), .Z(n20102) );
  OR U28590 ( .A(n20105), .B(n20106), .Z(n20104) );
  NANDN U28591 ( .A(n20107), .B(n20105), .Z(n20101) );
  IV U28592 ( .A(n20106), .Z(n20107) );
  XNOR U28593 ( .A(n20077), .B(n20108), .Z(n20072) );
  XNOR U28594 ( .A(n20075), .B(n20078), .Z(n20108) );
  NAND U28595 ( .A(n20109), .B(n20110), .Z(n20078) );
  NAND U28596 ( .A(n20111), .B(n20112), .Z(n20110) );
  OR U28597 ( .A(n20113), .B(n20114), .Z(n20111) );
  NANDN U28598 ( .A(n20115), .B(n20113), .Z(n20109) );
  IV U28599 ( .A(n20114), .Z(n20115) );
  NAND U28600 ( .A(n20116), .B(n20117), .Z(n20075) );
  NAND U28601 ( .A(n20118), .B(n20119), .Z(n20117) );
  NANDN U28602 ( .A(n20120), .B(n20121), .Z(n20118) );
  NANDN U28603 ( .A(n20121), .B(n20120), .Z(n20116) );
  AND U28604 ( .A(n20122), .B(n20123), .Z(n20077) );
  NAND U28605 ( .A(n20124), .B(n20125), .Z(n20123) );
  OR U28606 ( .A(n20126), .B(n20127), .Z(n20124) );
  NANDN U28607 ( .A(n20128), .B(n20126), .Z(n20122) );
  XNOR U28608 ( .A(n20103), .B(n20129), .Z(N63609) );
  XOR U28609 ( .A(n20105), .B(n20106), .Z(n20129) );
  XNOR U28610 ( .A(n20119), .B(n20130), .Z(n20106) );
  XOR U28611 ( .A(n20120), .B(n20121), .Z(n20130) );
  XOR U28612 ( .A(n20126), .B(n20131), .Z(n20121) );
  XOR U28613 ( .A(n20125), .B(n20128), .Z(n20131) );
  IV U28614 ( .A(n20127), .Z(n20128) );
  NAND U28615 ( .A(n20132), .B(n20133), .Z(n20127) );
  OR U28616 ( .A(n20134), .B(n20135), .Z(n20133) );
  OR U28617 ( .A(n20136), .B(n20137), .Z(n20132) );
  NAND U28618 ( .A(n20138), .B(n20139), .Z(n20125) );
  OR U28619 ( .A(n20140), .B(n20141), .Z(n20139) );
  OR U28620 ( .A(n20142), .B(n20143), .Z(n20138) );
  NOR U28621 ( .A(n20144), .B(n20145), .Z(n20126) );
  ANDN U28622 ( .B(n20146), .A(n20147), .Z(n20120) );
  XNOR U28623 ( .A(n20113), .B(n20148), .Z(n20119) );
  XNOR U28624 ( .A(n20112), .B(n20114), .Z(n20148) );
  NAND U28625 ( .A(n20149), .B(n20150), .Z(n20114) );
  OR U28626 ( .A(n20151), .B(n20152), .Z(n20150) );
  OR U28627 ( .A(n20153), .B(n20154), .Z(n20149) );
  NAND U28628 ( .A(n20155), .B(n20156), .Z(n20112) );
  OR U28629 ( .A(n20157), .B(n20158), .Z(n20156) );
  OR U28630 ( .A(n20159), .B(n20160), .Z(n20155) );
  ANDN U28631 ( .B(n20161), .A(n20162), .Z(n20113) );
  IV U28632 ( .A(n20163), .Z(n20161) );
  ANDN U28633 ( .B(n20164), .A(n20165), .Z(n20105) );
  XOR U28634 ( .A(n20091), .B(n20166), .Z(n20103) );
  XOR U28635 ( .A(n20092), .B(n20093), .Z(n20166) );
  XOR U28636 ( .A(n20098), .B(n20167), .Z(n20093) );
  XOR U28637 ( .A(n20097), .B(n20100), .Z(n20167) );
  IV U28638 ( .A(n20099), .Z(n20100) );
  NAND U28639 ( .A(n20168), .B(n20169), .Z(n20099) );
  OR U28640 ( .A(n20170), .B(n20171), .Z(n20169) );
  OR U28641 ( .A(n20172), .B(n20173), .Z(n20168) );
  NAND U28642 ( .A(n20174), .B(n20175), .Z(n20097) );
  OR U28643 ( .A(n20176), .B(n20177), .Z(n20175) );
  OR U28644 ( .A(n20178), .B(n20179), .Z(n20174) );
  NOR U28645 ( .A(n20180), .B(n20181), .Z(n20098) );
  ANDN U28646 ( .B(n20182), .A(n20183), .Z(n20092) );
  IV U28647 ( .A(n20184), .Z(n20182) );
  XNOR U28648 ( .A(n20085), .B(n20185), .Z(n20091) );
  XNOR U28649 ( .A(n20084), .B(n20086), .Z(n20185) );
  NAND U28650 ( .A(n20186), .B(n20187), .Z(n20086) );
  OR U28651 ( .A(n20188), .B(n20189), .Z(n20187) );
  OR U28652 ( .A(n20190), .B(n20191), .Z(n20186) );
  NAND U28653 ( .A(n20192), .B(n20193), .Z(n20084) );
  OR U28654 ( .A(n20194), .B(n20195), .Z(n20193) );
  OR U28655 ( .A(n20196), .B(n20197), .Z(n20192) );
  ANDN U28656 ( .B(n20198), .A(n20199), .Z(n20085) );
  IV U28657 ( .A(n20200), .Z(n20198) );
  XNOR U28658 ( .A(n20165), .B(n20164), .Z(N63608) );
  XOR U28659 ( .A(n20184), .B(n20183), .Z(n20164) );
  XNOR U28660 ( .A(n20199), .B(n20200), .Z(n20183) );
  XNOR U28661 ( .A(n20194), .B(n20195), .Z(n20200) );
  XNOR U28662 ( .A(n20196), .B(n20197), .Z(n20195) );
  XNOR U28663 ( .A(y[5581]), .B(x[5581]), .Z(n20197) );
  XNOR U28664 ( .A(y[5582]), .B(x[5582]), .Z(n20196) );
  XNOR U28665 ( .A(y[5580]), .B(x[5580]), .Z(n20194) );
  XNOR U28666 ( .A(n20188), .B(n20189), .Z(n20199) );
  XNOR U28667 ( .A(y[5577]), .B(x[5577]), .Z(n20189) );
  XNOR U28668 ( .A(n20190), .B(n20191), .Z(n20188) );
  XNOR U28669 ( .A(y[5578]), .B(x[5578]), .Z(n20191) );
  XNOR U28670 ( .A(y[5579]), .B(x[5579]), .Z(n20190) );
  XNOR U28671 ( .A(n20181), .B(n20180), .Z(n20184) );
  XNOR U28672 ( .A(n20176), .B(n20177), .Z(n20180) );
  XNOR U28673 ( .A(y[5574]), .B(x[5574]), .Z(n20177) );
  XNOR U28674 ( .A(n20178), .B(n20179), .Z(n20176) );
  XNOR U28675 ( .A(y[5575]), .B(x[5575]), .Z(n20179) );
  XNOR U28676 ( .A(y[5576]), .B(x[5576]), .Z(n20178) );
  XNOR U28677 ( .A(n20170), .B(n20171), .Z(n20181) );
  XNOR U28678 ( .A(y[5571]), .B(x[5571]), .Z(n20171) );
  XNOR U28679 ( .A(n20172), .B(n20173), .Z(n20170) );
  XNOR U28680 ( .A(y[5572]), .B(x[5572]), .Z(n20173) );
  XNOR U28681 ( .A(y[5573]), .B(x[5573]), .Z(n20172) );
  XOR U28682 ( .A(n20146), .B(n20147), .Z(n20165) );
  XNOR U28683 ( .A(n20162), .B(n20163), .Z(n20147) );
  XNOR U28684 ( .A(n20157), .B(n20158), .Z(n20163) );
  XNOR U28685 ( .A(n20159), .B(n20160), .Z(n20158) );
  XNOR U28686 ( .A(y[5569]), .B(x[5569]), .Z(n20160) );
  XNOR U28687 ( .A(y[5570]), .B(x[5570]), .Z(n20159) );
  XNOR U28688 ( .A(y[5568]), .B(x[5568]), .Z(n20157) );
  XNOR U28689 ( .A(n20151), .B(n20152), .Z(n20162) );
  XNOR U28690 ( .A(y[5565]), .B(x[5565]), .Z(n20152) );
  XNOR U28691 ( .A(n20153), .B(n20154), .Z(n20151) );
  XNOR U28692 ( .A(y[5566]), .B(x[5566]), .Z(n20154) );
  XNOR U28693 ( .A(y[5567]), .B(x[5567]), .Z(n20153) );
  XOR U28694 ( .A(n20145), .B(n20144), .Z(n20146) );
  XNOR U28695 ( .A(n20140), .B(n20141), .Z(n20144) );
  XNOR U28696 ( .A(y[5562]), .B(x[5562]), .Z(n20141) );
  XNOR U28697 ( .A(n20142), .B(n20143), .Z(n20140) );
  XNOR U28698 ( .A(y[5563]), .B(x[5563]), .Z(n20143) );
  XNOR U28699 ( .A(y[5564]), .B(x[5564]), .Z(n20142) );
  XNOR U28700 ( .A(n20134), .B(n20135), .Z(n20145) );
  XNOR U28701 ( .A(y[5559]), .B(x[5559]), .Z(n20135) );
  XNOR U28702 ( .A(n20136), .B(n20137), .Z(n20134) );
  XNOR U28703 ( .A(y[5560]), .B(x[5560]), .Z(n20137) );
  XNOR U28704 ( .A(y[5561]), .B(x[5561]), .Z(n20136) );
  NAND U28705 ( .A(n20201), .B(n20202), .Z(N63599) );
  NANDN U28706 ( .A(n20203), .B(n20204), .Z(n20202) );
  OR U28707 ( .A(n20205), .B(n20206), .Z(n20204) );
  NAND U28708 ( .A(n20205), .B(n20206), .Z(n20201) );
  XOR U28709 ( .A(n20205), .B(n20207), .Z(N63598) );
  XNOR U28710 ( .A(n20203), .B(n20206), .Z(n20207) );
  AND U28711 ( .A(n20208), .B(n20209), .Z(n20206) );
  NANDN U28712 ( .A(n20210), .B(n20211), .Z(n20209) );
  NANDN U28713 ( .A(n20212), .B(n20213), .Z(n20211) );
  NANDN U28714 ( .A(n20213), .B(n20212), .Z(n20208) );
  NAND U28715 ( .A(n20214), .B(n20215), .Z(n20203) );
  NANDN U28716 ( .A(n20216), .B(n20217), .Z(n20215) );
  OR U28717 ( .A(n20218), .B(n20219), .Z(n20217) );
  NAND U28718 ( .A(n20219), .B(n20218), .Z(n20214) );
  AND U28719 ( .A(n20220), .B(n20221), .Z(n20205) );
  NANDN U28720 ( .A(n20222), .B(n20223), .Z(n20221) );
  NANDN U28721 ( .A(n20224), .B(n20225), .Z(n20223) );
  NANDN U28722 ( .A(n20225), .B(n20224), .Z(n20220) );
  XOR U28723 ( .A(n20219), .B(n20226), .Z(N63597) );
  XOR U28724 ( .A(n20216), .B(n20218), .Z(n20226) );
  XNOR U28725 ( .A(n20212), .B(n20227), .Z(n20218) );
  XNOR U28726 ( .A(n20210), .B(n20213), .Z(n20227) );
  NAND U28727 ( .A(n20228), .B(n20229), .Z(n20213) );
  NAND U28728 ( .A(n20230), .B(n20231), .Z(n20229) );
  OR U28729 ( .A(n20232), .B(n20233), .Z(n20230) );
  NANDN U28730 ( .A(n20234), .B(n20232), .Z(n20228) );
  IV U28731 ( .A(n20233), .Z(n20234) );
  NAND U28732 ( .A(n20235), .B(n20236), .Z(n20210) );
  NAND U28733 ( .A(n20237), .B(n20238), .Z(n20236) );
  NANDN U28734 ( .A(n20239), .B(n20240), .Z(n20237) );
  NANDN U28735 ( .A(n20240), .B(n20239), .Z(n20235) );
  AND U28736 ( .A(n20241), .B(n20242), .Z(n20212) );
  NAND U28737 ( .A(n20243), .B(n20244), .Z(n20242) );
  OR U28738 ( .A(n20245), .B(n20246), .Z(n20243) );
  NANDN U28739 ( .A(n20247), .B(n20245), .Z(n20241) );
  NAND U28740 ( .A(n20248), .B(n20249), .Z(n20216) );
  NANDN U28741 ( .A(n20250), .B(n20251), .Z(n20249) );
  OR U28742 ( .A(n20252), .B(n20253), .Z(n20251) );
  NANDN U28743 ( .A(n20254), .B(n20252), .Z(n20248) );
  IV U28744 ( .A(n20253), .Z(n20254) );
  XNOR U28745 ( .A(n20224), .B(n20255), .Z(n20219) );
  XNOR U28746 ( .A(n20222), .B(n20225), .Z(n20255) );
  NAND U28747 ( .A(n20256), .B(n20257), .Z(n20225) );
  NAND U28748 ( .A(n20258), .B(n20259), .Z(n20257) );
  OR U28749 ( .A(n20260), .B(n20261), .Z(n20258) );
  NANDN U28750 ( .A(n20262), .B(n20260), .Z(n20256) );
  IV U28751 ( .A(n20261), .Z(n20262) );
  NAND U28752 ( .A(n20263), .B(n20264), .Z(n20222) );
  NAND U28753 ( .A(n20265), .B(n20266), .Z(n20264) );
  NANDN U28754 ( .A(n20267), .B(n20268), .Z(n20265) );
  NANDN U28755 ( .A(n20268), .B(n20267), .Z(n20263) );
  AND U28756 ( .A(n20269), .B(n20270), .Z(n20224) );
  NAND U28757 ( .A(n20271), .B(n20272), .Z(n20270) );
  OR U28758 ( .A(n20273), .B(n20274), .Z(n20271) );
  NANDN U28759 ( .A(n20275), .B(n20273), .Z(n20269) );
  XNOR U28760 ( .A(n20250), .B(n20276), .Z(N63596) );
  XOR U28761 ( .A(n20252), .B(n20253), .Z(n20276) );
  XNOR U28762 ( .A(n20266), .B(n20277), .Z(n20253) );
  XOR U28763 ( .A(n20267), .B(n20268), .Z(n20277) );
  XOR U28764 ( .A(n20273), .B(n20278), .Z(n20268) );
  XOR U28765 ( .A(n20272), .B(n20275), .Z(n20278) );
  IV U28766 ( .A(n20274), .Z(n20275) );
  NAND U28767 ( .A(n20279), .B(n20280), .Z(n20274) );
  OR U28768 ( .A(n20281), .B(n20282), .Z(n20280) );
  OR U28769 ( .A(n20283), .B(n20284), .Z(n20279) );
  NAND U28770 ( .A(n20285), .B(n20286), .Z(n20272) );
  OR U28771 ( .A(n20287), .B(n20288), .Z(n20286) );
  OR U28772 ( .A(n20289), .B(n20290), .Z(n20285) );
  NOR U28773 ( .A(n20291), .B(n20292), .Z(n20273) );
  ANDN U28774 ( .B(n20293), .A(n20294), .Z(n20267) );
  XNOR U28775 ( .A(n20260), .B(n20295), .Z(n20266) );
  XNOR U28776 ( .A(n20259), .B(n20261), .Z(n20295) );
  NAND U28777 ( .A(n20296), .B(n20297), .Z(n20261) );
  OR U28778 ( .A(n20298), .B(n20299), .Z(n20297) );
  OR U28779 ( .A(n20300), .B(n20301), .Z(n20296) );
  NAND U28780 ( .A(n20302), .B(n20303), .Z(n20259) );
  OR U28781 ( .A(n20304), .B(n20305), .Z(n20303) );
  OR U28782 ( .A(n20306), .B(n20307), .Z(n20302) );
  ANDN U28783 ( .B(n20308), .A(n20309), .Z(n20260) );
  IV U28784 ( .A(n20310), .Z(n20308) );
  ANDN U28785 ( .B(n20311), .A(n20312), .Z(n20252) );
  XOR U28786 ( .A(n20238), .B(n20313), .Z(n20250) );
  XOR U28787 ( .A(n20239), .B(n20240), .Z(n20313) );
  XOR U28788 ( .A(n20245), .B(n20314), .Z(n20240) );
  XOR U28789 ( .A(n20244), .B(n20247), .Z(n20314) );
  IV U28790 ( .A(n20246), .Z(n20247) );
  NAND U28791 ( .A(n20315), .B(n20316), .Z(n20246) );
  OR U28792 ( .A(n20317), .B(n20318), .Z(n20316) );
  OR U28793 ( .A(n20319), .B(n20320), .Z(n20315) );
  NAND U28794 ( .A(n20321), .B(n20322), .Z(n20244) );
  OR U28795 ( .A(n20323), .B(n20324), .Z(n20322) );
  OR U28796 ( .A(n20325), .B(n20326), .Z(n20321) );
  NOR U28797 ( .A(n20327), .B(n20328), .Z(n20245) );
  ANDN U28798 ( .B(n20329), .A(n20330), .Z(n20239) );
  IV U28799 ( .A(n20331), .Z(n20329) );
  XNOR U28800 ( .A(n20232), .B(n20332), .Z(n20238) );
  XNOR U28801 ( .A(n20231), .B(n20233), .Z(n20332) );
  NAND U28802 ( .A(n20333), .B(n20334), .Z(n20233) );
  OR U28803 ( .A(n20335), .B(n20336), .Z(n20334) );
  OR U28804 ( .A(n20337), .B(n20338), .Z(n20333) );
  NAND U28805 ( .A(n20339), .B(n20340), .Z(n20231) );
  OR U28806 ( .A(n20341), .B(n20342), .Z(n20340) );
  OR U28807 ( .A(n20343), .B(n20344), .Z(n20339) );
  ANDN U28808 ( .B(n20345), .A(n20346), .Z(n20232) );
  IV U28809 ( .A(n20347), .Z(n20345) );
  XNOR U28810 ( .A(n20312), .B(n20311), .Z(N63595) );
  XOR U28811 ( .A(n20331), .B(n20330), .Z(n20311) );
  XNOR U28812 ( .A(n20346), .B(n20347), .Z(n20330) );
  XNOR U28813 ( .A(n20341), .B(n20342), .Z(n20347) );
  XNOR U28814 ( .A(n20343), .B(n20344), .Z(n20342) );
  XNOR U28815 ( .A(y[5557]), .B(x[5557]), .Z(n20344) );
  XNOR U28816 ( .A(y[5558]), .B(x[5558]), .Z(n20343) );
  XNOR U28817 ( .A(y[5556]), .B(x[5556]), .Z(n20341) );
  XNOR U28818 ( .A(n20335), .B(n20336), .Z(n20346) );
  XNOR U28819 ( .A(y[5553]), .B(x[5553]), .Z(n20336) );
  XNOR U28820 ( .A(n20337), .B(n20338), .Z(n20335) );
  XNOR U28821 ( .A(y[5554]), .B(x[5554]), .Z(n20338) );
  XNOR U28822 ( .A(y[5555]), .B(x[5555]), .Z(n20337) );
  XNOR U28823 ( .A(n20328), .B(n20327), .Z(n20331) );
  XNOR U28824 ( .A(n20323), .B(n20324), .Z(n20327) );
  XNOR U28825 ( .A(y[5550]), .B(x[5550]), .Z(n20324) );
  XNOR U28826 ( .A(n20325), .B(n20326), .Z(n20323) );
  XNOR U28827 ( .A(y[5551]), .B(x[5551]), .Z(n20326) );
  XNOR U28828 ( .A(y[5552]), .B(x[5552]), .Z(n20325) );
  XNOR U28829 ( .A(n20317), .B(n20318), .Z(n20328) );
  XNOR U28830 ( .A(y[5547]), .B(x[5547]), .Z(n20318) );
  XNOR U28831 ( .A(n20319), .B(n20320), .Z(n20317) );
  XNOR U28832 ( .A(y[5548]), .B(x[5548]), .Z(n20320) );
  XNOR U28833 ( .A(y[5549]), .B(x[5549]), .Z(n20319) );
  XOR U28834 ( .A(n20293), .B(n20294), .Z(n20312) );
  XNOR U28835 ( .A(n20309), .B(n20310), .Z(n20294) );
  XNOR U28836 ( .A(n20304), .B(n20305), .Z(n20310) );
  XNOR U28837 ( .A(n20306), .B(n20307), .Z(n20305) );
  XNOR U28838 ( .A(y[5545]), .B(x[5545]), .Z(n20307) );
  XNOR U28839 ( .A(y[5546]), .B(x[5546]), .Z(n20306) );
  XNOR U28840 ( .A(y[5544]), .B(x[5544]), .Z(n20304) );
  XNOR U28841 ( .A(n20298), .B(n20299), .Z(n20309) );
  XNOR U28842 ( .A(y[5541]), .B(x[5541]), .Z(n20299) );
  XNOR U28843 ( .A(n20300), .B(n20301), .Z(n20298) );
  XNOR U28844 ( .A(y[5542]), .B(x[5542]), .Z(n20301) );
  XNOR U28845 ( .A(y[5543]), .B(x[5543]), .Z(n20300) );
  XOR U28846 ( .A(n20292), .B(n20291), .Z(n20293) );
  XNOR U28847 ( .A(n20287), .B(n20288), .Z(n20291) );
  XNOR U28848 ( .A(y[5538]), .B(x[5538]), .Z(n20288) );
  XNOR U28849 ( .A(n20289), .B(n20290), .Z(n20287) );
  XNOR U28850 ( .A(y[5539]), .B(x[5539]), .Z(n20290) );
  XNOR U28851 ( .A(y[5540]), .B(x[5540]), .Z(n20289) );
  XNOR U28852 ( .A(n20281), .B(n20282), .Z(n20292) );
  XNOR U28853 ( .A(y[5535]), .B(x[5535]), .Z(n20282) );
  XNOR U28854 ( .A(n20283), .B(n20284), .Z(n20281) );
  XNOR U28855 ( .A(y[5536]), .B(x[5536]), .Z(n20284) );
  XNOR U28856 ( .A(y[5537]), .B(x[5537]), .Z(n20283) );
  NAND U28857 ( .A(n20348), .B(n20349), .Z(N63586) );
  NANDN U28858 ( .A(n20350), .B(n20351), .Z(n20349) );
  OR U28859 ( .A(n20352), .B(n20353), .Z(n20351) );
  NAND U28860 ( .A(n20352), .B(n20353), .Z(n20348) );
  XOR U28861 ( .A(n20352), .B(n20354), .Z(N63585) );
  XNOR U28862 ( .A(n20350), .B(n20353), .Z(n20354) );
  AND U28863 ( .A(n20355), .B(n20356), .Z(n20353) );
  NANDN U28864 ( .A(n20357), .B(n20358), .Z(n20356) );
  NANDN U28865 ( .A(n20359), .B(n20360), .Z(n20358) );
  NANDN U28866 ( .A(n20360), .B(n20359), .Z(n20355) );
  NAND U28867 ( .A(n20361), .B(n20362), .Z(n20350) );
  NANDN U28868 ( .A(n20363), .B(n20364), .Z(n20362) );
  OR U28869 ( .A(n20365), .B(n20366), .Z(n20364) );
  NAND U28870 ( .A(n20366), .B(n20365), .Z(n20361) );
  AND U28871 ( .A(n20367), .B(n20368), .Z(n20352) );
  NANDN U28872 ( .A(n20369), .B(n20370), .Z(n20368) );
  NANDN U28873 ( .A(n20371), .B(n20372), .Z(n20370) );
  NANDN U28874 ( .A(n20372), .B(n20371), .Z(n20367) );
  XOR U28875 ( .A(n20366), .B(n20373), .Z(N63584) );
  XOR U28876 ( .A(n20363), .B(n20365), .Z(n20373) );
  XNOR U28877 ( .A(n20359), .B(n20374), .Z(n20365) );
  XNOR U28878 ( .A(n20357), .B(n20360), .Z(n20374) );
  NAND U28879 ( .A(n20375), .B(n20376), .Z(n20360) );
  NAND U28880 ( .A(n20377), .B(n20378), .Z(n20376) );
  OR U28881 ( .A(n20379), .B(n20380), .Z(n20377) );
  NANDN U28882 ( .A(n20381), .B(n20379), .Z(n20375) );
  IV U28883 ( .A(n20380), .Z(n20381) );
  NAND U28884 ( .A(n20382), .B(n20383), .Z(n20357) );
  NAND U28885 ( .A(n20384), .B(n20385), .Z(n20383) );
  NANDN U28886 ( .A(n20386), .B(n20387), .Z(n20384) );
  NANDN U28887 ( .A(n20387), .B(n20386), .Z(n20382) );
  AND U28888 ( .A(n20388), .B(n20389), .Z(n20359) );
  NAND U28889 ( .A(n20390), .B(n20391), .Z(n20389) );
  OR U28890 ( .A(n20392), .B(n20393), .Z(n20390) );
  NANDN U28891 ( .A(n20394), .B(n20392), .Z(n20388) );
  NAND U28892 ( .A(n20395), .B(n20396), .Z(n20363) );
  NANDN U28893 ( .A(n20397), .B(n20398), .Z(n20396) );
  OR U28894 ( .A(n20399), .B(n20400), .Z(n20398) );
  NANDN U28895 ( .A(n20401), .B(n20399), .Z(n20395) );
  IV U28896 ( .A(n20400), .Z(n20401) );
  XNOR U28897 ( .A(n20371), .B(n20402), .Z(n20366) );
  XNOR U28898 ( .A(n20369), .B(n20372), .Z(n20402) );
  NAND U28899 ( .A(n20403), .B(n20404), .Z(n20372) );
  NAND U28900 ( .A(n20405), .B(n20406), .Z(n20404) );
  OR U28901 ( .A(n20407), .B(n20408), .Z(n20405) );
  NANDN U28902 ( .A(n20409), .B(n20407), .Z(n20403) );
  IV U28903 ( .A(n20408), .Z(n20409) );
  NAND U28904 ( .A(n20410), .B(n20411), .Z(n20369) );
  NAND U28905 ( .A(n20412), .B(n20413), .Z(n20411) );
  NANDN U28906 ( .A(n20414), .B(n20415), .Z(n20412) );
  NANDN U28907 ( .A(n20415), .B(n20414), .Z(n20410) );
  AND U28908 ( .A(n20416), .B(n20417), .Z(n20371) );
  NAND U28909 ( .A(n20418), .B(n20419), .Z(n20417) );
  OR U28910 ( .A(n20420), .B(n20421), .Z(n20418) );
  NANDN U28911 ( .A(n20422), .B(n20420), .Z(n20416) );
  XNOR U28912 ( .A(n20397), .B(n20423), .Z(N63583) );
  XOR U28913 ( .A(n20399), .B(n20400), .Z(n20423) );
  XNOR U28914 ( .A(n20413), .B(n20424), .Z(n20400) );
  XOR U28915 ( .A(n20414), .B(n20415), .Z(n20424) );
  XOR U28916 ( .A(n20420), .B(n20425), .Z(n20415) );
  XOR U28917 ( .A(n20419), .B(n20422), .Z(n20425) );
  IV U28918 ( .A(n20421), .Z(n20422) );
  NAND U28919 ( .A(n20426), .B(n20427), .Z(n20421) );
  OR U28920 ( .A(n20428), .B(n20429), .Z(n20427) );
  OR U28921 ( .A(n20430), .B(n20431), .Z(n20426) );
  NAND U28922 ( .A(n20432), .B(n20433), .Z(n20419) );
  OR U28923 ( .A(n20434), .B(n20435), .Z(n20433) );
  OR U28924 ( .A(n20436), .B(n20437), .Z(n20432) );
  NOR U28925 ( .A(n20438), .B(n20439), .Z(n20420) );
  ANDN U28926 ( .B(n20440), .A(n20441), .Z(n20414) );
  XNOR U28927 ( .A(n20407), .B(n20442), .Z(n20413) );
  XNOR U28928 ( .A(n20406), .B(n20408), .Z(n20442) );
  NAND U28929 ( .A(n20443), .B(n20444), .Z(n20408) );
  OR U28930 ( .A(n20445), .B(n20446), .Z(n20444) );
  OR U28931 ( .A(n20447), .B(n20448), .Z(n20443) );
  NAND U28932 ( .A(n20449), .B(n20450), .Z(n20406) );
  OR U28933 ( .A(n20451), .B(n20452), .Z(n20450) );
  OR U28934 ( .A(n20453), .B(n20454), .Z(n20449) );
  ANDN U28935 ( .B(n20455), .A(n20456), .Z(n20407) );
  IV U28936 ( .A(n20457), .Z(n20455) );
  ANDN U28937 ( .B(n20458), .A(n20459), .Z(n20399) );
  XOR U28938 ( .A(n20385), .B(n20460), .Z(n20397) );
  XOR U28939 ( .A(n20386), .B(n20387), .Z(n20460) );
  XOR U28940 ( .A(n20392), .B(n20461), .Z(n20387) );
  XOR U28941 ( .A(n20391), .B(n20394), .Z(n20461) );
  IV U28942 ( .A(n20393), .Z(n20394) );
  NAND U28943 ( .A(n20462), .B(n20463), .Z(n20393) );
  OR U28944 ( .A(n20464), .B(n20465), .Z(n20463) );
  OR U28945 ( .A(n20466), .B(n20467), .Z(n20462) );
  NAND U28946 ( .A(n20468), .B(n20469), .Z(n20391) );
  OR U28947 ( .A(n20470), .B(n20471), .Z(n20469) );
  OR U28948 ( .A(n20472), .B(n20473), .Z(n20468) );
  NOR U28949 ( .A(n20474), .B(n20475), .Z(n20392) );
  ANDN U28950 ( .B(n20476), .A(n20477), .Z(n20386) );
  IV U28951 ( .A(n20478), .Z(n20476) );
  XNOR U28952 ( .A(n20379), .B(n20479), .Z(n20385) );
  XNOR U28953 ( .A(n20378), .B(n20380), .Z(n20479) );
  NAND U28954 ( .A(n20480), .B(n20481), .Z(n20380) );
  OR U28955 ( .A(n20482), .B(n20483), .Z(n20481) );
  OR U28956 ( .A(n20484), .B(n20485), .Z(n20480) );
  NAND U28957 ( .A(n20486), .B(n20487), .Z(n20378) );
  OR U28958 ( .A(n20488), .B(n20489), .Z(n20487) );
  OR U28959 ( .A(n20490), .B(n20491), .Z(n20486) );
  ANDN U28960 ( .B(n20492), .A(n20493), .Z(n20379) );
  IV U28961 ( .A(n20494), .Z(n20492) );
  XNOR U28962 ( .A(n20459), .B(n20458), .Z(N63582) );
  XOR U28963 ( .A(n20478), .B(n20477), .Z(n20458) );
  XNOR U28964 ( .A(n20493), .B(n20494), .Z(n20477) );
  XNOR U28965 ( .A(n20488), .B(n20489), .Z(n20494) );
  XNOR U28966 ( .A(n20490), .B(n20491), .Z(n20489) );
  XNOR U28967 ( .A(y[5533]), .B(x[5533]), .Z(n20491) );
  XNOR U28968 ( .A(y[5534]), .B(x[5534]), .Z(n20490) );
  XNOR U28969 ( .A(y[5532]), .B(x[5532]), .Z(n20488) );
  XNOR U28970 ( .A(n20482), .B(n20483), .Z(n20493) );
  XNOR U28971 ( .A(y[5529]), .B(x[5529]), .Z(n20483) );
  XNOR U28972 ( .A(n20484), .B(n20485), .Z(n20482) );
  XNOR U28973 ( .A(y[5530]), .B(x[5530]), .Z(n20485) );
  XNOR U28974 ( .A(y[5531]), .B(x[5531]), .Z(n20484) );
  XNOR U28975 ( .A(n20475), .B(n20474), .Z(n20478) );
  XNOR U28976 ( .A(n20470), .B(n20471), .Z(n20474) );
  XNOR U28977 ( .A(y[5526]), .B(x[5526]), .Z(n20471) );
  XNOR U28978 ( .A(n20472), .B(n20473), .Z(n20470) );
  XNOR U28979 ( .A(y[5527]), .B(x[5527]), .Z(n20473) );
  XNOR U28980 ( .A(y[5528]), .B(x[5528]), .Z(n20472) );
  XNOR U28981 ( .A(n20464), .B(n20465), .Z(n20475) );
  XNOR U28982 ( .A(y[5523]), .B(x[5523]), .Z(n20465) );
  XNOR U28983 ( .A(n20466), .B(n20467), .Z(n20464) );
  XNOR U28984 ( .A(y[5524]), .B(x[5524]), .Z(n20467) );
  XNOR U28985 ( .A(y[5525]), .B(x[5525]), .Z(n20466) );
  XOR U28986 ( .A(n20440), .B(n20441), .Z(n20459) );
  XNOR U28987 ( .A(n20456), .B(n20457), .Z(n20441) );
  XNOR U28988 ( .A(n20451), .B(n20452), .Z(n20457) );
  XNOR U28989 ( .A(n20453), .B(n20454), .Z(n20452) );
  XNOR U28990 ( .A(y[5521]), .B(x[5521]), .Z(n20454) );
  XNOR U28991 ( .A(y[5522]), .B(x[5522]), .Z(n20453) );
  XNOR U28992 ( .A(y[5520]), .B(x[5520]), .Z(n20451) );
  XNOR U28993 ( .A(n20445), .B(n20446), .Z(n20456) );
  XNOR U28994 ( .A(y[5517]), .B(x[5517]), .Z(n20446) );
  XNOR U28995 ( .A(n20447), .B(n20448), .Z(n20445) );
  XNOR U28996 ( .A(y[5518]), .B(x[5518]), .Z(n20448) );
  XNOR U28997 ( .A(y[5519]), .B(x[5519]), .Z(n20447) );
  XOR U28998 ( .A(n20439), .B(n20438), .Z(n20440) );
  XNOR U28999 ( .A(n20434), .B(n20435), .Z(n20438) );
  XNOR U29000 ( .A(y[5514]), .B(x[5514]), .Z(n20435) );
  XNOR U29001 ( .A(n20436), .B(n20437), .Z(n20434) );
  XNOR U29002 ( .A(y[5515]), .B(x[5515]), .Z(n20437) );
  XNOR U29003 ( .A(y[5516]), .B(x[5516]), .Z(n20436) );
  XNOR U29004 ( .A(n20428), .B(n20429), .Z(n20439) );
  XNOR U29005 ( .A(y[5511]), .B(x[5511]), .Z(n20429) );
  XNOR U29006 ( .A(n20430), .B(n20431), .Z(n20428) );
  XNOR U29007 ( .A(y[5512]), .B(x[5512]), .Z(n20431) );
  XNOR U29008 ( .A(y[5513]), .B(x[5513]), .Z(n20430) );
  NAND U29009 ( .A(n20495), .B(n20496), .Z(N63573) );
  NANDN U29010 ( .A(n20497), .B(n20498), .Z(n20496) );
  OR U29011 ( .A(n20499), .B(n20500), .Z(n20498) );
  NAND U29012 ( .A(n20499), .B(n20500), .Z(n20495) );
  XOR U29013 ( .A(n20499), .B(n20501), .Z(N63572) );
  XNOR U29014 ( .A(n20497), .B(n20500), .Z(n20501) );
  AND U29015 ( .A(n20502), .B(n20503), .Z(n20500) );
  NANDN U29016 ( .A(n20504), .B(n20505), .Z(n20503) );
  NANDN U29017 ( .A(n20506), .B(n20507), .Z(n20505) );
  NANDN U29018 ( .A(n20507), .B(n20506), .Z(n20502) );
  NAND U29019 ( .A(n20508), .B(n20509), .Z(n20497) );
  NANDN U29020 ( .A(n20510), .B(n20511), .Z(n20509) );
  OR U29021 ( .A(n20512), .B(n20513), .Z(n20511) );
  NAND U29022 ( .A(n20513), .B(n20512), .Z(n20508) );
  AND U29023 ( .A(n20514), .B(n20515), .Z(n20499) );
  NANDN U29024 ( .A(n20516), .B(n20517), .Z(n20515) );
  NANDN U29025 ( .A(n20518), .B(n20519), .Z(n20517) );
  NANDN U29026 ( .A(n20519), .B(n20518), .Z(n20514) );
  XOR U29027 ( .A(n20513), .B(n20520), .Z(N63571) );
  XOR U29028 ( .A(n20510), .B(n20512), .Z(n20520) );
  XNOR U29029 ( .A(n20506), .B(n20521), .Z(n20512) );
  XNOR U29030 ( .A(n20504), .B(n20507), .Z(n20521) );
  NAND U29031 ( .A(n20522), .B(n20523), .Z(n20507) );
  NAND U29032 ( .A(n20524), .B(n20525), .Z(n20523) );
  OR U29033 ( .A(n20526), .B(n20527), .Z(n20524) );
  NANDN U29034 ( .A(n20528), .B(n20526), .Z(n20522) );
  IV U29035 ( .A(n20527), .Z(n20528) );
  NAND U29036 ( .A(n20529), .B(n20530), .Z(n20504) );
  NAND U29037 ( .A(n20531), .B(n20532), .Z(n20530) );
  NANDN U29038 ( .A(n20533), .B(n20534), .Z(n20531) );
  NANDN U29039 ( .A(n20534), .B(n20533), .Z(n20529) );
  AND U29040 ( .A(n20535), .B(n20536), .Z(n20506) );
  NAND U29041 ( .A(n20537), .B(n20538), .Z(n20536) );
  OR U29042 ( .A(n20539), .B(n20540), .Z(n20537) );
  NANDN U29043 ( .A(n20541), .B(n20539), .Z(n20535) );
  NAND U29044 ( .A(n20542), .B(n20543), .Z(n20510) );
  NANDN U29045 ( .A(n20544), .B(n20545), .Z(n20543) );
  OR U29046 ( .A(n20546), .B(n20547), .Z(n20545) );
  NANDN U29047 ( .A(n20548), .B(n20546), .Z(n20542) );
  IV U29048 ( .A(n20547), .Z(n20548) );
  XNOR U29049 ( .A(n20518), .B(n20549), .Z(n20513) );
  XNOR U29050 ( .A(n20516), .B(n20519), .Z(n20549) );
  NAND U29051 ( .A(n20550), .B(n20551), .Z(n20519) );
  NAND U29052 ( .A(n20552), .B(n20553), .Z(n20551) );
  OR U29053 ( .A(n20554), .B(n20555), .Z(n20552) );
  NANDN U29054 ( .A(n20556), .B(n20554), .Z(n20550) );
  IV U29055 ( .A(n20555), .Z(n20556) );
  NAND U29056 ( .A(n20557), .B(n20558), .Z(n20516) );
  NAND U29057 ( .A(n20559), .B(n20560), .Z(n20558) );
  NANDN U29058 ( .A(n20561), .B(n20562), .Z(n20559) );
  NANDN U29059 ( .A(n20562), .B(n20561), .Z(n20557) );
  AND U29060 ( .A(n20563), .B(n20564), .Z(n20518) );
  NAND U29061 ( .A(n20565), .B(n20566), .Z(n20564) );
  OR U29062 ( .A(n20567), .B(n20568), .Z(n20565) );
  NANDN U29063 ( .A(n20569), .B(n20567), .Z(n20563) );
  XNOR U29064 ( .A(n20544), .B(n20570), .Z(N63570) );
  XOR U29065 ( .A(n20546), .B(n20547), .Z(n20570) );
  XNOR U29066 ( .A(n20560), .B(n20571), .Z(n20547) );
  XOR U29067 ( .A(n20561), .B(n20562), .Z(n20571) );
  XOR U29068 ( .A(n20567), .B(n20572), .Z(n20562) );
  XOR U29069 ( .A(n20566), .B(n20569), .Z(n20572) );
  IV U29070 ( .A(n20568), .Z(n20569) );
  NAND U29071 ( .A(n20573), .B(n20574), .Z(n20568) );
  OR U29072 ( .A(n20575), .B(n20576), .Z(n20574) );
  OR U29073 ( .A(n20577), .B(n20578), .Z(n20573) );
  NAND U29074 ( .A(n20579), .B(n20580), .Z(n20566) );
  OR U29075 ( .A(n20581), .B(n20582), .Z(n20580) );
  OR U29076 ( .A(n20583), .B(n20584), .Z(n20579) );
  NOR U29077 ( .A(n20585), .B(n20586), .Z(n20567) );
  ANDN U29078 ( .B(n20587), .A(n20588), .Z(n20561) );
  XNOR U29079 ( .A(n20554), .B(n20589), .Z(n20560) );
  XNOR U29080 ( .A(n20553), .B(n20555), .Z(n20589) );
  NAND U29081 ( .A(n20590), .B(n20591), .Z(n20555) );
  OR U29082 ( .A(n20592), .B(n20593), .Z(n20591) );
  OR U29083 ( .A(n20594), .B(n20595), .Z(n20590) );
  NAND U29084 ( .A(n20596), .B(n20597), .Z(n20553) );
  OR U29085 ( .A(n20598), .B(n20599), .Z(n20597) );
  OR U29086 ( .A(n20600), .B(n20601), .Z(n20596) );
  ANDN U29087 ( .B(n20602), .A(n20603), .Z(n20554) );
  IV U29088 ( .A(n20604), .Z(n20602) );
  ANDN U29089 ( .B(n20605), .A(n20606), .Z(n20546) );
  XOR U29090 ( .A(n20532), .B(n20607), .Z(n20544) );
  XOR U29091 ( .A(n20533), .B(n20534), .Z(n20607) );
  XOR U29092 ( .A(n20539), .B(n20608), .Z(n20534) );
  XOR U29093 ( .A(n20538), .B(n20541), .Z(n20608) );
  IV U29094 ( .A(n20540), .Z(n20541) );
  NAND U29095 ( .A(n20609), .B(n20610), .Z(n20540) );
  OR U29096 ( .A(n20611), .B(n20612), .Z(n20610) );
  OR U29097 ( .A(n20613), .B(n20614), .Z(n20609) );
  NAND U29098 ( .A(n20615), .B(n20616), .Z(n20538) );
  OR U29099 ( .A(n20617), .B(n20618), .Z(n20616) );
  OR U29100 ( .A(n20619), .B(n20620), .Z(n20615) );
  NOR U29101 ( .A(n20621), .B(n20622), .Z(n20539) );
  ANDN U29102 ( .B(n20623), .A(n20624), .Z(n20533) );
  IV U29103 ( .A(n20625), .Z(n20623) );
  XNOR U29104 ( .A(n20526), .B(n20626), .Z(n20532) );
  XNOR U29105 ( .A(n20525), .B(n20527), .Z(n20626) );
  NAND U29106 ( .A(n20627), .B(n20628), .Z(n20527) );
  OR U29107 ( .A(n20629), .B(n20630), .Z(n20628) );
  OR U29108 ( .A(n20631), .B(n20632), .Z(n20627) );
  NAND U29109 ( .A(n20633), .B(n20634), .Z(n20525) );
  OR U29110 ( .A(n20635), .B(n20636), .Z(n20634) );
  OR U29111 ( .A(n20637), .B(n20638), .Z(n20633) );
  ANDN U29112 ( .B(n20639), .A(n20640), .Z(n20526) );
  IV U29113 ( .A(n20641), .Z(n20639) );
  XNOR U29114 ( .A(n20606), .B(n20605), .Z(N63569) );
  XOR U29115 ( .A(n20625), .B(n20624), .Z(n20605) );
  XNOR U29116 ( .A(n20640), .B(n20641), .Z(n20624) );
  XNOR U29117 ( .A(n20635), .B(n20636), .Z(n20641) );
  XNOR U29118 ( .A(n20637), .B(n20638), .Z(n20636) );
  XNOR U29119 ( .A(y[5509]), .B(x[5509]), .Z(n20638) );
  XNOR U29120 ( .A(y[5510]), .B(x[5510]), .Z(n20637) );
  XNOR U29121 ( .A(y[5508]), .B(x[5508]), .Z(n20635) );
  XNOR U29122 ( .A(n20629), .B(n20630), .Z(n20640) );
  XNOR U29123 ( .A(y[5505]), .B(x[5505]), .Z(n20630) );
  XNOR U29124 ( .A(n20631), .B(n20632), .Z(n20629) );
  XNOR U29125 ( .A(y[5506]), .B(x[5506]), .Z(n20632) );
  XNOR U29126 ( .A(y[5507]), .B(x[5507]), .Z(n20631) );
  XNOR U29127 ( .A(n20622), .B(n20621), .Z(n20625) );
  XNOR U29128 ( .A(n20617), .B(n20618), .Z(n20621) );
  XNOR U29129 ( .A(y[5502]), .B(x[5502]), .Z(n20618) );
  XNOR U29130 ( .A(n20619), .B(n20620), .Z(n20617) );
  XNOR U29131 ( .A(y[5503]), .B(x[5503]), .Z(n20620) );
  XNOR U29132 ( .A(y[5504]), .B(x[5504]), .Z(n20619) );
  XNOR U29133 ( .A(n20611), .B(n20612), .Z(n20622) );
  XNOR U29134 ( .A(y[5499]), .B(x[5499]), .Z(n20612) );
  XNOR U29135 ( .A(n20613), .B(n20614), .Z(n20611) );
  XNOR U29136 ( .A(y[5500]), .B(x[5500]), .Z(n20614) );
  XNOR U29137 ( .A(y[5501]), .B(x[5501]), .Z(n20613) );
  XOR U29138 ( .A(n20587), .B(n20588), .Z(n20606) );
  XNOR U29139 ( .A(n20603), .B(n20604), .Z(n20588) );
  XNOR U29140 ( .A(n20598), .B(n20599), .Z(n20604) );
  XNOR U29141 ( .A(n20600), .B(n20601), .Z(n20599) );
  XNOR U29142 ( .A(y[5497]), .B(x[5497]), .Z(n20601) );
  XNOR U29143 ( .A(y[5498]), .B(x[5498]), .Z(n20600) );
  XNOR U29144 ( .A(y[5496]), .B(x[5496]), .Z(n20598) );
  XNOR U29145 ( .A(n20592), .B(n20593), .Z(n20603) );
  XNOR U29146 ( .A(y[5493]), .B(x[5493]), .Z(n20593) );
  XNOR U29147 ( .A(n20594), .B(n20595), .Z(n20592) );
  XNOR U29148 ( .A(y[5494]), .B(x[5494]), .Z(n20595) );
  XNOR U29149 ( .A(y[5495]), .B(x[5495]), .Z(n20594) );
  XOR U29150 ( .A(n20586), .B(n20585), .Z(n20587) );
  XNOR U29151 ( .A(n20581), .B(n20582), .Z(n20585) );
  XNOR U29152 ( .A(y[5490]), .B(x[5490]), .Z(n20582) );
  XNOR U29153 ( .A(n20583), .B(n20584), .Z(n20581) );
  XNOR U29154 ( .A(y[5491]), .B(x[5491]), .Z(n20584) );
  XNOR U29155 ( .A(y[5492]), .B(x[5492]), .Z(n20583) );
  XNOR U29156 ( .A(n20575), .B(n20576), .Z(n20586) );
  XNOR U29157 ( .A(y[5487]), .B(x[5487]), .Z(n20576) );
  XNOR U29158 ( .A(n20577), .B(n20578), .Z(n20575) );
  XNOR U29159 ( .A(y[5488]), .B(x[5488]), .Z(n20578) );
  XNOR U29160 ( .A(y[5489]), .B(x[5489]), .Z(n20577) );
  NAND U29161 ( .A(n20642), .B(n20643), .Z(N63560) );
  NANDN U29162 ( .A(n20644), .B(n20645), .Z(n20643) );
  OR U29163 ( .A(n20646), .B(n20647), .Z(n20645) );
  NAND U29164 ( .A(n20646), .B(n20647), .Z(n20642) );
  XOR U29165 ( .A(n20646), .B(n20648), .Z(N63559) );
  XNOR U29166 ( .A(n20644), .B(n20647), .Z(n20648) );
  AND U29167 ( .A(n20649), .B(n20650), .Z(n20647) );
  NANDN U29168 ( .A(n20651), .B(n20652), .Z(n20650) );
  NANDN U29169 ( .A(n20653), .B(n20654), .Z(n20652) );
  NANDN U29170 ( .A(n20654), .B(n20653), .Z(n20649) );
  NAND U29171 ( .A(n20655), .B(n20656), .Z(n20644) );
  NANDN U29172 ( .A(n20657), .B(n20658), .Z(n20656) );
  OR U29173 ( .A(n20659), .B(n20660), .Z(n20658) );
  NAND U29174 ( .A(n20660), .B(n20659), .Z(n20655) );
  AND U29175 ( .A(n20661), .B(n20662), .Z(n20646) );
  NANDN U29176 ( .A(n20663), .B(n20664), .Z(n20662) );
  NANDN U29177 ( .A(n20665), .B(n20666), .Z(n20664) );
  NANDN U29178 ( .A(n20666), .B(n20665), .Z(n20661) );
  XOR U29179 ( .A(n20660), .B(n20667), .Z(N63558) );
  XOR U29180 ( .A(n20657), .B(n20659), .Z(n20667) );
  XNOR U29181 ( .A(n20653), .B(n20668), .Z(n20659) );
  XNOR U29182 ( .A(n20651), .B(n20654), .Z(n20668) );
  NAND U29183 ( .A(n20669), .B(n20670), .Z(n20654) );
  NAND U29184 ( .A(n20671), .B(n20672), .Z(n20670) );
  OR U29185 ( .A(n20673), .B(n20674), .Z(n20671) );
  NANDN U29186 ( .A(n20675), .B(n20673), .Z(n20669) );
  IV U29187 ( .A(n20674), .Z(n20675) );
  NAND U29188 ( .A(n20676), .B(n20677), .Z(n20651) );
  NAND U29189 ( .A(n20678), .B(n20679), .Z(n20677) );
  NANDN U29190 ( .A(n20680), .B(n20681), .Z(n20678) );
  NANDN U29191 ( .A(n20681), .B(n20680), .Z(n20676) );
  AND U29192 ( .A(n20682), .B(n20683), .Z(n20653) );
  NAND U29193 ( .A(n20684), .B(n20685), .Z(n20683) );
  OR U29194 ( .A(n20686), .B(n20687), .Z(n20684) );
  NANDN U29195 ( .A(n20688), .B(n20686), .Z(n20682) );
  NAND U29196 ( .A(n20689), .B(n20690), .Z(n20657) );
  NANDN U29197 ( .A(n20691), .B(n20692), .Z(n20690) );
  OR U29198 ( .A(n20693), .B(n20694), .Z(n20692) );
  NANDN U29199 ( .A(n20695), .B(n20693), .Z(n20689) );
  IV U29200 ( .A(n20694), .Z(n20695) );
  XNOR U29201 ( .A(n20665), .B(n20696), .Z(n20660) );
  XNOR U29202 ( .A(n20663), .B(n20666), .Z(n20696) );
  NAND U29203 ( .A(n20697), .B(n20698), .Z(n20666) );
  NAND U29204 ( .A(n20699), .B(n20700), .Z(n20698) );
  OR U29205 ( .A(n20701), .B(n20702), .Z(n20699) );
  NANDN U29206 ( .A(n20703), .B(n20701), .Z(n20697) );
  IV U29207 ( .A(n20702), .Z(n20703) );
  NAND U29208 ( .A(n20704), .B(n20705), .Z(n20663) );
  NAND U29209 ( .A(n20706), .B(n20707), .Z(n20705) );
  NANDN U29210 ( .A(n20708), .B(n20709), .Z(n20706) );
  NANDN U29211 ( .A(n20709), .B(n20708), .Z(n20704) );
  AND U29212 ( .A(n20710), .B(n20711), .Z(n20665) );
  NAND U29213 ( .A(n20712), .B(n20713), .Z(n20711) );
  OR U29214 ( .A(n20714), .B(n20715), .Z(n20712) );
  NANDN U29215 ( .A(n20716), .B(n20714), .Z(n20710) );
  XNOR U29216 ( .A(n20691), .B(n20717), .Z(N63557) );
  XOR U29217 ( .A(n20693), .B(n20694), .Z(n20717) );
  XNOR U29218 ( .A(n20707), .B(n20718), .Z(n20694) );
  XOR U29219 ( .A(n20708), .B(n20709), .Z(n20718) );
  XOR U29220 ( .A(n20714), .B(n20719), .Z(n20709) );
  XOR U29221 ( .A(n20713), .B(n20716), .Z(n20719) );
  IV U29222 ( .A(n20715), .Z(n20716) );
  NAND U29223 ( .A(n20720), .B(n20721), .Z(n20715) );
  OR U29224 ( .A(n20722), .B(n20723), .Z(n20721) );
  OR U29225 ( .A(n20724), .B(n20725), .Z(n20720) );
  NAND U29226 ( .A(n20726), .B(n20727), .Z(n20713) );
  OR U29227 ( .A(n20728), .B(n20729), .Z(n20727) );
  OR U29228 ( .A(n20730), .B(n20731), .Z(n20726) );
  NOR U29229 ( .A(n20732), .B(n20733), .Z(n20714) );
  ANDN U29230 ( .B(n20734), .A(n20735), .Z(n20708) );
  XNOR U29231 ( .A(n20701), .B(n20736), .Z(n20707) );
  XNOR U29232 ( .A(n20700), .B(n20702), .Z(n20736) );
  NAND U29233 ( .A(n20737), .B(n20738), .Z(n20702) );
  OR U29234 ( .A(n20739), .B(n20740), .Z(n20738) );
  OR U29235 ( .A(n20741), .B(n20742), .Z(n20737) );
  NAND U29236 ( .A(n20743), .B(n20744), .Z(n20700) );
  OR U29237 ( .A(n20745), .B(n20746), .Z(n20744) );
  OR U29238 ( .A(n20747), .B(n20748), .Z(n20743) );
  ANDN U29239 ( .B(n20749), .A(n20750), .Z(n20701) );
  IV U29240 ( .A(n20751), .Z(n20749) );
  ANDN U29241 ( .B(n20752), .A(n20753), .Z(n20693) );
  XOR U29242 ( .A(n20679), .B(n20754), .Z(n20691) );
  XOR U29243 ( .A(n20680), .B(n20681), .Z(n20754) );
  XOR U29244 ( .A(n20686), .B(n20755), .Z(n20681) );
  XOR U29245 ( .A(n20685), .B(n20688), .Z(n20755) );
  IV U29246 ( .A(n20687), .Z(n20688) );
  NAND U29247 ( .A(n20756), .B(n20757), .Z(n20687) );
  OR U29248 ( .A(n20758), .B(n20759), .Z(n20757) );
  OR U29249 ( .A(n20760), .B(n20761), .Z(n20756) );
  NAND U29250 ( .A(n20762), .B(n20763), .Z(n20685) );
  OR U29251 ( .A(n20764), .B(n20765), .Z(n20763) );
  OR U29252 ( .A(n20766), .B(n20767), .Z(n20762) );
  NOR U29253 ( .A(n20768), .B(n20769), .Z(n20686) );
  ANDN U29254 ( .B(n20770), .A(n20771), .Z(n20680) );
  IV U29255 ( .A(n20772), .Z(n20770) );
  XNOR U29256 ( .A(n20673), .B(n20773), .Z(n20679) );
  XNOR U29257 ( .A(n20672), .B(n20674), .Z(n20773) );
  NAND U29258 ( .A(n20774), .B(n20775), .Z(n20674) );
  OR U29259 ( .A(n20776), .B(n20777), .Z(n20775) );
  OR U29260 ( .A(n20778), .B(n20779), .Z(n20774) );
  NAND U29261 ( .A(n20780), .B(n20781), .Z(n20672) );
  OR U29262 ( .A(n20782), .B(n20783), .Z(n20781) );
  OR U29263 ( .A(n20784), .B(n20785), .Z(n20780) );
  ANDN U29264 ( .B(n20786), .A(n20787), .Z(n20673) );
  IV U29265 ( .A(n20788), .Z(n20786) );
  XNOR U29266 ( .A(n20753), .B(n20752), .Z(N63556) );
  XOR U29267 ( .A(n20772), .B(n20771), .Z(n20752) );
  XNOR U29268 ( .A(n20787), .B(n20788), .Z(n20771) );
  XNOR U29269 ( .A(n20782), .B(n20783), .Z(n20788) );
  XNOR U29270 ( .A(n20784), .B(n20785), .Z(n20783) );
  XNOR U29271 ( .A(y[5485]), .B(x[5485]), .Z(n20785) );
  XNOR U29272 ( .A(y[5486]), .B(x[5486]), .Z(n20784) );
  XNOR U29273 ( .A(y[5484]), .B(x[5484]), .Z(n20782) );
  XNOR U29274 ( .A(n20776), .B(n20777), .Z(n20787) );
  XNOR U29275 ( .A(y[5481]), .B(x[5481]), .Z(n20777) );
  XNOR U29276 ( .A(n20778), .B(n20779), .Z(n20776) );
  XNOR U29277 ( .A(y[5482]), .B(x[5482]), .Z(n20779) );
  XNOR U29278 ( .A(y[5483]), .B(x[5483]), .Z(n20778) );
  XNOR U29279 ( .A(n20769), .B(n20768), .Z(n20772) );
  XNOR U29280 ( .A(n20764), .B(n20765), .Z(n20768) );
  XNOR U29281 ( .A(y[5478]), .B(x[5478]), .Z(n20765) );
  XNOR U29282 ( .A(n20766), .B(n20767), .Z(n20764) );
  XNOR U29283 ( .A(y[5479]), .B(x[5479]), .Z(n20767) );
  XNOR U29284 ( .A(y[5480]), .B(x[5480]), .Z(n20766) );
  XNOR U29285 ( .A(n20758), .B(n20759), .Z(n20769) );
  XNOR U29286 ( .A(y[5475]), .B(x[5475]), .Z(n20759) );
  XNOR U29287 ( .A(n20760), .B(n20761), .Z(n20758) );
  XNOR U29288 ( .A(y[5476]), .B(x[5476]), .Z(n20761) );
  XNOR U29289 ( .A(y[5477]), .B(x[5477]), .Z(n20760) );
  XOR U29290 ( .A(n20734), .B(n20735), .Z(n20753) );
  XNOR U29291 ( .A(n20750), .B(n20751), .Z(n20735) );
  XNOR U29292 ( .A(n20745), .B(n20746), .Z(n20751) );
  XNOR U29293 ( .A(n20747), .B(n20748), .Z(n20746) );
  XNOR U29294 ( .A(y[5473]), .B(x[5473]), .Z(n20748) );
  XNOR U29295 ( .A(y[5474]), .B(x[5474]), .Z(n20747) );
  XNOR U29296 ( .A(y[5472]), .B(x[5472]), .Z(n20745) );
  XNOR U29297 ( .A(n20739), .B(n20740), .Z(n20750) );
  XNOR U29298 ( .A(y[5469]), .B(x[5469]), .Z(n20740) );
  XNOR U29299 ( .A(n20741), .B(n20742), .Z(n20739) );
  XNOR U29300 ( .A(y[5470]), .B(x[5470]), .Z(n20742) );
  XNOR U29301 ( .A(y[5471]), .B(x[5471]), .Z(n20741) );
  XOR U29302 ( .A(n20733), .B(n20732), .Z(n20734) );
  XNOR U29303 ( .A(n20728), .B(n20729), .Z(n20732) );
  XNOR U29304 ( .A(y[5466]), .B(x[5466]), .Z(n20729) );
  XNOR U29305 ( .A(n20730), .B(n20731), .Z(n20728) );
  XNOR U29306 ( .A(y[5467]), .B(x[5467]), .Z(n20731) );
  XNOR U29307 ( .A(y[5468]), .B(x[5468]), .Z(n20730) );
  XNOR U29308 ( .A(n20722), .B(n20723), .Z(n20733) );
  XNOR U29309 ( .A(y[5463]), .B(x[5463]), .Z(n20723) );
  XNOR U29310 ( .A(n20724), .B(n20725), .Z(n20722) );
  XNOR U29311 ( .A(y[5464]), .B(x[5464]), .Z(n20725) );
  XNOR U29312 ( .A(y[5465]), .B(x[5465]), .Z(n20724) );
  NAND U29313 ( .A(n20789), .B(n20790), .Z(N63547) );
  NANDN U29314 ( .A(n20791), .B(n20792), .Z(n20790) );
  OR U29315 ( .A(n20793), .B(n20794), .Z(n20792) );
  NAND U29316 ( .A(n20793), .B(n20794), .Z(n20789) );
  XOR U29317 ( .A(n20793), .B(n20795), .Z(N63546) );
  XNOR U29318 ( .A(n20791), .B(n20794), .Z(n20795) );
  AND U29319 ( .A(n20796), .B(n20797), .Z(n20794) );
  NANDN U29320 ( .A(n20798), .B(n20799), .Z(n20797) );
  NANDN U29321 ( .A(n20800), .B(n20801), .Z(n20799) );
  NANDN U29322 ( .A(n20801), .B(n20800), .Z(n20796) );
  NAND U29323 ( .A(n20802), .B(n20803), .Z(n20791) );
  NANDN U29324 ( .A(n20804), .B(n20805), .Z(n20803) );
  OR U29325 ( .A(n20806), .B(n20807), .Z(n20805) );
  NAND U29326 ( .A(n20807), .B(n20806), .Z(n20802) );
  AND U29327 ( .A(n20808), .B(n20809), .Z(n20793) );
  NANDN U29328 ( .A(n20810), .B(n20811), .Z(n20809) );
  NANDN U29329 ( .A(n20812), .B(n20813), .Z(n20811) );
  NANDN U29330 ( .A(n20813), .B(n20812), .Z(n20808) );
  XOR U29331 ( .A(n20807), .B(n20814), .Z(N63545) );
  XOR U29332 ( .A(n20804), .B(n20806), .Z(n20814) );
  XNOR U29333 ( .A(n20800), .B(n20815), .Z(n20806) );
  XNOR U29334 ( .A(n20798), .B(n20801), .Z(n20815) );
  NAND U29335 ( .A(n20816), .B(n20817), .Z(n20801) );
  NAND U29336 ( .A(n20818), .B(n20819), .Z(n20817) );
  OR U29337 ( .A(n20820), .B(n20821), .Z(n20818) );
  NANDN U29338 ( .A(n20822), .B(n20820), .Z(n20816) );
  IV U29339 ( .A(n20821), .Z(n20822) );
  NAND U29340 ( .A(n20823), .B(n20824), .Z(n20798) );
  NAND U29341 ( .A(n20825), .B(n20826), .Z(n20824) );
  NANDN U29342 ( .A(n20827), .B(n20828), .Z(n20825) );
  NANDN U29343 ( .A(n20828), .B(n20827), .Z(n20823) );
  AND U29344 ( .A(n20829), .B(n20830), .Z(n20800) );
  NAND U29345 ( .A(n20831), .B(n20832), .Z(n20830) );
  OR U29346 ( .A(n20833), .B(n20834), .Z(n20831) );
  NANDN U29347 ( .A(n20835), .B(n20833), .Z(n20829) );
  NAND U29348 ( .A(n20836), .B(n20837), .Z(n20804) );
  NANDN U29349 ( .A(n20838), .B(n20839), .Z(n20837) );
  OR U29350 ( .A(n20840), .B(n20841), .Z(n20839) );
  NANDN U29351 ( .A(n20842), .B(n20840), .Z(n20836) );
  IV U29352 ( .A(n20841), .Z(n20842) );
  XNOR U29353 ( .A(n20812), .B(n20843), .Z(n20807) );
  XNOR U29354 ( .A(n20810), .B(n20813), .Z(n20843) );
  NAND U29355 ( .A(n20844), .B(n20845), .Z(n20813) );
  NAND U29356 ( .A(n20846), .B(n20847), .Z(n20845) );
  OR U29357 ( .A(n20848), .B(n20849), .Z(n20846) );
  NANDN U29358 ( .A(n20850), .B(n20848), .Z(n20844) );
  IV U29359 ( .A(n20849), .Z(n20850) );
  NAND U29360 ( .A(n20851), .B(n20852), .Z(n20810) );
  NAND U29361 ( .A(n20853), .B(n20854), .Z(n20852) );
  NANDN U29362 ( .A(n20855), .B(n20856), .Z(n20853) );
  NANDN U29363 ( .A(n20856), .B(n20855), .Z(n20851) );
  AND U29364 ( .A(n20857), .B(n20858), .Z(n20812) );
  NAND U29365 ( .A(n20859), .B(n20860), .Z(n20858) );
  OR U29366 ( .A(n20861), .B(n20862), .Z(n20859) );
  NANDN U29367 ( .A(n20863), .B(n20861), .Z(n20857) );
  XNOR U29368 ( .A(n20838), .B(n20864), .Z(N63544) );
  XOR U29369 ( .A(n20840), .B(n20841), .Z(n20864) );
  XNOR U29370 ( .A(n20854), .B(n20865), .Z(n20841) );
  XOR U29371 ( .A(n20855), .B(n20856), .Z(n20865) );
  XOR U29372 ( .A(n20861), .B(n20866), .Z(n20856) );
  XOR U29373 ( .A(n20860), .B(n20863), .Z(n20866) );
  IV U29374 ( .A(n20862), .Z(n20863) );
  NAND U29375 ( .A(n20867), .B(n20868), .Z(n20862) );
  OR U29376 ( .A(n20869), .B(n20870), .Z(n20868) );
  OR U29377 ( .A(n20871), .B(n20872), .Z(n20867) );
  NAND U29378 ( .A(n20873), .B(n20874), .Z(n20860) );
  OR U29379 ( .A(n20875), .B(n20876), .Z(n20874) );
  OR U29380 ( .A(n20877), .B(n20878), .Z(n20873) );
  NOR U29381 ( .A(n20879), .B(n20880), .Z(n20861) );
  ANDN U29382 ( .B(n20881), .A(n20882), .Z(n20855) );
  XNOR U29383 ( .A(n20848), .B(n20883), .Z(n20854) );
  XNOR U29384 ( .A(n20847), .B(n20849), .Z(n20883) );
  NAND U29385 ( .A(n20884), .B(n20885), .Z(n20849) );
  OR U29386 ( .A(n20886), .B(n20887), .Z(n20885) );
  OR U29387 ( .A(n20888), .B(n20889), .Z(n20884) );
  NAND U29388 ( .A(n20890), .B(n20891), .Z(n20847) );
  OR U29389 ( .A(n20892), .B(n20893), .Z(n20891) );
  OR U29390 ( .A(n20894), .B(n20895), .Z(n20890) );
  ANDN U29391 ( .B(n20896), .A(n20897), .Z(n20848) );
  IV U29392 ( .A(n20898), .Z(n20896) );
  ANDN U29393 ( .B(n20899), .A(n20900), .Z(n20840) );
  XOR U29394 ( .A(n20826), .B(n20901), .Z(n20838) );
  XOR U29395 ( .A(n20827), .B(n20828), .Z(n20901) );
  XOR U29396 ( .A(n20833), .B(n20902), .Z(n20828) );
  XOR U29397 ( .A(n20832), .B(n20835), .Z(n20902) );
  IV U29398 ( .A(n20834), .Z(n20835) );
  NAND U29399 ( .A(n20903), .B(n20904), .Z(n20834) );
  OR U29400 ( .A(n20905), .B(n20906), .Z(n20904) );
  OR U29401 ( .A(n20907), .B(n20908), .Z(n20903) );
  NAND U29402 ( .A(n20909), .B(n20910), .Z(n20832) );
  OR U29403 ( .A(n20911), .B(n20912), .Z(n20910) );
  OR U29404 ( .A(n20913), .B(n20914), .Z(n20909) );
  NOR U29405 ( .A(n20915), .B(n20916), .Z(n20833) );
  ANDN U29406 ( .B(n20917), .A(n20918), .Z(n20827) );
  IV U29407 ( .A(n20919), .Z(n20917) );
  XNOR U29408 ( .A(n20820), .B(n20920), .Z(n20826) );
  XNOR U29409 ( .A(n20819), .B(n20821), .Z(n20920) );
  NAND U29410 ( .A(n20921), .B(n20922), .Z(n20821) );
  OR U29411 ( .A(n20923), .B(n20924), .Z(n20922) );
  OR U29412 ( .A(n20925), .B(n20926), .Z(n20921) );
  NAND U29413 ( .A(n20927), .B(n20928), .Z(n20819) );
  OR U29414 ( .A(n20929), .B(n20930), .Z(n20928) );
  OR U29415 ( .A(n20931), .B(n20932), .Z(n20927) );
  ANDN U29416 ( .B(n20933), .A(n20934), .Z(n20820) );
  IV U29417 ( .A(n20935), .Z(n20933) );
  XNOR U29418 ( .A(n20900), .B(n20899), .Z(N63543) );
  XOR U29419 ( .A(n20919), .B(n20918), .Z(n20899) );
  XNOR U29420 ( .A(n20934), .B(n20935), .Z(n20918) );
  XNOR U29421 ( .A(n20929), .B(n20930), .Z(n20935) );
  XNOR U29422 ( .A(n20931), .B(n20932), .Z(n20930) );
  XNOR U29423 ( .A(y[5461]), .B(x[5461]), .Z(n20932) );
  XNOR U29424 ( .A(y[5462]), .B(x[5462]), .Z(n20931) );
  XNOR U29425 ( .A(y[5460]), .B(x[5460]), .Z(n20929) );
  XNOR U29426 ( .A(n20923), .B(n20924), .Z(n20934) );
  XNOR U29427 ( .A(y[5457]), .B(x[5457]), .Z(n20924) );
  XNOR U29428 ( .A(n20925), .B(n20926), .Z(n20923) );
  XNOR U29429 ( .A(y[5458]), .B(x[5458]), .Z(n20926) );
  XNOR U29430 ( .A(y[5459]), .B(x[5459]), .Z(n20925) );
  XNOR U29431 ( .A(n20916), .B(n20915), .Z(n20919) );
  XNOR U29432 ( .A(n20911), .B(n20912), .Z(n20915) );
  XNOR U29433 ( .A(y[5454]), .B(x[5454]), .Z(n20912) );
  XNOR U29434 ( .A(n20913), .B(n20914), .Z(n20911) );
  XNOR U29435 ( .A(y[5455]), .B(x[5455]), .Z(n20914) );
  XNOR U29436 ( .A(y[5456]), .B(x[5456]), .Z(n20913) );
  XNOR U29437 ( .A(n20905), .B(n20906), .Z(n20916) );
  XNOR U29438 ( .A(y[5451]), .B(x[5451]), .Z(n20906) );
  XNOR U29439 ( .A(n20907), .B(n20908), .Z(n20905) );
  XNOR U29440 ( .A(y[5452]), .B(x[5452]), .Z(n20908) );
  XNOR U29441 ( .A(y[5453]), .B(x[5453]), .Z(n20907) );
  XOR U29442 ( .A(n20881), .B(n20882), .Z(n20900) );
  XNOR U29443 ( .A(n20897), .B(n20898), .Z(n20882) );
  XNOR U29444 ( .A(n20892), .B(n20893), .Z(n20898) );
  XNOR U29445 ( .A(n20894), .B(n20895), .Z(n20893) );
  XNOR U29446 ( .A(y[5449]), .B(x[5449]), .Z(n20895) );
  XNOR U29447 ( .A(y[5450]), .B(x[5450]), .Z(n20894) );
  XNOR U29448 ( .A(y[5448]), .B(x[5448]), .Z(n20892) );
  XNOR U29449 ( .A(n20886), .B(n20887), .Z(n20897) );
  XNOR U29450 ( .A(y[5445]), .B(x[5445]), .Z(n20887) );
  XNOR U29451 ( .A(n20888), .B(n20889), .Z(n20886) );
  XNOR U29452 ( .A(y[5446]), .B(x[5446]), .Z(n20889) );
  XNOR U29453 ( .A(y[5447]), .B(x[5447]), .Z(n20888) );
  XOR U29454 ( .A(n20880), .B(n20879), .Z(n20881) );
  XNOR U29455 ( .A(n20875), .B(n20876), .Z(n20879) );
  XNOR U29456 ( .A(y[5442]), .B(x[5442]), .Z(n20876) );
  XNOR U29457 ( .A(n20877), .B(n20878), .Z(n20875) );
  XNOR U29458 ( .A(y[5443]), .B(x[5443]), .Z(n20878) );
  XNOR U29459 ( .A(y[5444]), .B(x[5444]), .Z(n20877) );
  XNOR U29460 ( .A(n20869), .B(n20870), .Z(n20880) );
  XNOR U29461 ( .A(y[5439]), .B(x[5439]), .Z(n20870) );
  XNOR U29462 ( .A(n20871), .B(n20872), .Z(n20869) );
  XNOR U29463 ( .A(y[5440]), .B(x[5440]), .Z(n20872) );
  XNOR U29464 ( .A(y[5441]), .B(x[5441]), .Z(n20871) );
  NAND U29465 ( .A(n20936), .B(n20937), .Z(N63534) );
  NANDN U29466 ( .A(n20938), .B(n20939), .Z(n20937) );
  OR U29467 ( .A(n20940), .B(n20941), .Z(n20939) );
  NAND U29468 ( .A(n20940), .B(n20941), .Z(n20936) );
  XOR U29469 ( .A(n20940), .B(n20942), .Z(N63533) );
  XNOR U29470 ( .A(n20938), .B(n20941), .Z(n20942) );
  AND U29471 ( .A(n20943), .B(n20944), .Z(n20941) );
  NANDN U29472 ( .A(n20945), .B(n20946), .Z(n20944) );
  NANDN U29473 ( .A(n20947), .B(n20948), .Z(n20946) );
  NANDN U29474 ( .A(n20948), .B(n20947), .Z(n20943) );
  NAND U29475 ( .A(n20949), .B(n20950), .Z(n20938) );
  NANDN U29476 ( .A(n20951), .B(n20952), .Z(n20950) );
  OR U29477 ( .A(n20953), .B(n20954), .Z(n20952) );
  NAND U29478 ( .A(n20954), .B(n20953), .Z(n20949) );
  AND U29479 ( .A(n20955), .B(n20956), .Z(n20940) );
  NANDN U29480 ( .A(n20957), .B(n20958), .Z(n20956) );
  NANDN U29481 ( .A(n20959), .B(n20960), .Z(n20958) );
  NANDN U29482 ( .A(n20960), .B(n20959), .Z(n20955) );
  XOR U29483 ( .A(n20954), .B(n20961), .Z(N63532) );
  XOR U29484 ( .A(n20951), .B(n20953), .Z(n20961) );
  XNOR U29485 ( .A(n20947), .B(n20962), .Z(n20953) );
  XNOR U29486 ( .A(n20945), .B(n20948), .Z(n20962) );
  NAND U29487 ( .A(n20963), .B(n20964), .Z(n20948) );
  NAND U29488 ( .A(n20965), .B(n20966), .Z(n20964) );
  OR U29489 ( .A(n20967), .B(n20968), .Z(n20965) );
  NANDN U29490 ( .A(n20969), .B(n20967), .Z(n20963) );
  IV U29491 ( .A(n20968), .Z(n20969) );
  NAND U29492 ( .A(n20970), .B(n20971), .Z(n20945) );
  NAND U29493 ( .A(n20972), .B(n20973), .Z(n20971) );
  NANDN U29494 ( .A(n20974), .B(n20975), .Z(n20972) );
  NANDN U29495 ( .A(n20975), .B(n20974), .Z(n20970) );
  AND U29496 ( .A(n20976), .B(n20977), .Z(n20947) );
  NAND U29497 ( .A(n20978), .B(n20979), .Z(n20977) );
  OR U29498 ( .A(n20980), .B(n20981), .Z(n20978) );
  NANDN U29499 ( .A(n20982), .B(n20980), .Z(n20976) );
  NAND U29500 ( .A(n20983), .B(n20984), .Z(n20951) );
  NANDN U29501 ( .A(n20985), .B(n20986), .Z(n20984) );
  OR U29502 ( .A(n20987), .B(n20988), .Z(n20986) );
  NANDN U29503 ( .A(n20989), .B(n20987), .Z(n20983) );
  IV U29504 ( .A(n20988), .Z(n20989) );
  XNOR U29505 ( .A(n20959), .B(n20990), .Z(n20954) );
  XNOR U29506 ( .A(n20957), .B(n20960), .Z(n20990) );
  NAND U29507 ( .A(n20991), .B(n20992), .Z(n20960) );
  NAND U29508 ( .A(n20993), .B(n20994), .Z(n20992) );
  OR U29509 ( .A(n20995), .B(n20996), .Z(n20993) );
  NANDN U29510 ( .A(n20997), .B(n20995), .Z(n20991) );
  IV U29511 ( .A(n20996), .Z(n20997) );
  NAND U29512 ( .A(n20998), .B(n20999), .Z(n20957) );
  NAND U29513 ( .A(n21000), .B(n21001), .Z(n20999) );
  NANDN U29514 ( .A(n21002), .B(n21003), .Z(n21000) );
  NANDN U29515 ( .A(n21003), .B(n21002), .Z(n20998) );
  AND U29516 ( .A(n21004), .B(n21005), .Z(n20959) );
  NAND U29517 ( .A(n21006), .B(n21007), .Z(n21005) );
  OR U29518 ( .A(n21008), .B(n21009), .Z(n21006) );
  NANDN U29519 ( .A(n21010), .B(n21008), .Z(n21004) );
  XNOR U29520 ( .A(n20985), .B(n21011), .Z(N63531) );
  XOR U29521 ( .A(n20987), .B(n20988), .Z(n21011) );
  XNOR U29522 ( .A(n21001), .B(n21012), .Z(n20988) );
  XOR U29523 ( .A(n21002), .B(n21003), .Z(n21012) );
  XOR U29524 ( .A(n21008), .B(n21013), .Z(n21003) );
  XOR U29525 ( .A(n21007), .B(n21010), .Z(n21013) );
  IV U29526 ( .A(n21009), .Z(n21010) );
  NAND U29527 ( .A(n21014), .B(n21015), .Z(n21009) );
  OR U29528 ( .A(n21016), .B(n21017), .Z(n21015) );
  OR U29529 ( .A(n21018), .B(n21019), .Z(n21014) );
  NAND U29530 ( .A(n21020), .B(n21021), .Z(n21007) );
  OR U29531 ( .A(n21022), .B(n21023), .Z(n21021) );
  OR U29532 ( .A(n21024), .B(n21025), .Z(n21020) );
  NOR U29533 ( .A(n21026), .B(n21027), .Z(n21008) );
  ANDN U29534 ( .B(n21028), .A(n21029), .Z(n21002) );
  XNOR U29535 ( .A(n20995), .B(n21030), .Z(n21001) );
  XNOR U29536 ( .A(n20994), .B(n20996), .Z(n21030) );
  NAND U29537 ( .A(n21031), .B(n21032), .Z(n20996) );
  OR U29538 ( .A(n21033), .B(n21034), .Z(n21032) );
  OR U29539 ( .A(n21035), .B(n21036), .Z(n21031) );
  NAND U29540 ( .A(n21037), .B(n21038), .Z(n20994) );
  OR U29541 ( .A(n21039), .B(n21040), .Z(n21038) );
  OR U29542 ( .A(n21041), .B(n21042), .Z(n21037) );
  ANDN U29543 ( .B(n21043), .A(n21044), .Z(n20995) );
  IV U29544 ( .A(n21045), .Z(n21043) );
  ANDN U29545 ( .B(n21046), .A(n21047), .Z(n20987) );
  XOR U29546 ( .A(n20973), .B(n21048), .Z(n20985) );
  XOR U29547 ( .A(n20974), .B(n20975), .Z(n21048) );
  XOR U29548 ( .A(n20980), .B(n21049), .Z(n20975) );
  XOR U29549 ( .A(n20979), .B(n20982), .Z(n21049) );
  IV U29550 ( .A(n20981), .Z(n20982) );
  NAND U29551 ( .A(n21050), .B(n21051), .Z(n20981) );
  OR U29552 ( .A(n21052), .B(n21053), .Z(n21051) );
  OR U29553 ( .A(n21054), .B(n21055), .Z(n21050) );
  NAND U29554 ( .A(n21056), .B(n21057), .Z(n20979) );
  OR U29555 ( .A(n21058), .B(n21059), .Z(n21057) );
  OR U29556 ( .A(n21060), .B(n21061), .Z(n21056) );
  NOR U29557 ( .A(n21062), .B(n21063), .Z(n20980) );
  ANDN U29558 ( .B(n21064), .A(n21065), .Z(n20974) );
  IV U29559 ( .A(n21066), .Z(n21064) );
  XNOR U29560 ( .A(n20967), .B(n21067), .Z(n20973) );
  XNOR U29561 ( .A(n20966), .B(n20968), .Z(n21067) );
  NAND U29562 ( .A(n21068), .B(n21069), .Z(n20968) );
  OR U29563 ( .A(n21070), .B(n21071), .Z(n21069) );
  OR U29564 ( .A(n21072), .B(n21073), .Z(n21068) );
  NAND U29565 ( .A(n21074), .B(n21075), .Z(n20966) );
  OR U29566 ( .A(n21076), .B(n21077), .Z(n21075) );
  OR U29567 ( .A(n21078), .B(n21079), .Z(n21074) );
  ANDN U29568 ( .B(n21080), .A(n21081), .Z(n20967) );
  IV U29569 ( .A(n21082), .Z(n21080) );
  XNOR U29570 ( .A(n21047), .B(n21046), .Z(N63530) );
  XOR U29571 ( .A(n21066), .B(n21065), .Z(n21046) );
  XNOR U29572 ( .A(n21081), .B(n21082), .Z(n21065) );
  XNOR U29573 ( .A(n21076), .B(n21077), .Z(n21082) );
  XNOR U29574 ( .A(n21078), .B(n21079), .Z(n21077) );
  XNOR U29575 ( .A(y[5437]), .B(x[5437]), .Z(n21079) );
  XNOR U29576 ( .A(y[5438]), .B(x[5438]), .Z(n21078) );
  XNOR U29577 ( .A(y[5436]), .B(x[5436]), .Z(n21076) );
  XNOR U29578 ( .A(n21070), .B(n21071), .Z(n21081) );
  XNOR U29579 ( .A(y[5433]), .B(x[5433]), .Z(n21071) );
  XNOR U29580 ( .A(n21072), .B(n21073), .Z(n21070) );
  XNOR U29581 ( .A(y[5434]), .B(x[5434]), .Z(n21073) );
  XNOR U29582 ( .A(y[5435]), .B(x[5435]), .Z(n21072) );
  XNOR U29583 ( .A(n21063), .B(n21062), .Z(n21066) );
  XNOR U29584 ( .A(n21058), .B(n21059), .Z(n21062) );
  XNOR U29585 ( .A(y[5430]), .B(x[5430]), .Z(n21059) );
  XNOR U29586 ( .A(n21060), .B(n21061), .Z(n21058) );
  XNOR U29587 ( .A(y[5431]), .B(x[5431]), .Z(n21061) );
  XNOR U29588 ( .A(y[5432]), .B(x[5432]), .Z(n21060) );
  XNOR U29589 ( .A(n21052), .B(n21053), .Z(n21063) );
  XNOR U29590 ( .A(y[5427]), .B(x[5427]), .Z(n21053) );
  XNOR U29591 ( .A(n21054), .B(n21055), .Z(n21052) );
  XNOR U29592 ( .A(y[5428]), .B(x[5428]), .Z(n21055) );
  XNOR U29593 ( .A(y[5429]), .B(x[5429]), .Z(n21054) );
  XOR U29594 ( .A(n21028), .B(n21029), .Z(n21047) );
  XNOR U29595 ( .A(n21044), .B(n21045), .Z(n21029) );
  XNOR U29596 ( .A(n21039), .B(n21040), .Z(n21045) );
  XNOR U29597 ( .A(n21041), .B(n21042), .Z(n21040) );
  XNOR U29598 ( .A(y[5425]), .B(x[5425]), .Z(n21042) );
  XNOR U29599 ( .A(y[5426]), .B(x[5426]), .Z(n21041) );
  XNOR U29600 ( .A(y[5424]), .B(x[5424]), .Z(n21039) );
  XNOR U29601 ( .A(n21033), .B(n21034), .Z(n21044) );
  XNOR U29602 ( .A(y[5421]), .B(x[5421]), .Z(n21034) );
  XNOR U29603 ( .A(n21035), .B(n21036), .Z(n21033) );
  XNOR U29604 ( .A(y[5422]), .B(x[5422]), .Z(n21036) );
  XNOR U29605 ( .A(y[5423]), .B(x[5423]), .Z(n21035) );
  XOR U29606 ( .A(n21027), .B(n21026), .Z(n21028) );
  XNOR U29607 ( .A(n21022), .B(n21023), .Z(n21026) );
  XNOR U29608 ( .A(y[5418]), .B(x[5418]), .Z(n21023) );
  XNOR U29609 ( .A(n21024), .B(n21025), .Z(n21022) );
  XNOR U29610 ( .A(y[5419]), .B(x[5419]), .Z(n21025) );
  XNOR U29611 ( .A(y[5420]), .B(x[5420]), .Z(n21024) );
  XNOR U29612 ( .A(n21016), .B(n21017), .Z(n21027) );
  XNOR U29613 ( .A(y[5415]), .B(x[5415]), .Z(n21017) );
  XNOR U29614 ( .A(n21018), .B(n21019), .Z(n21016) );
  XNOR U29615 ( .A(y[5416]), .B(x[5416]), .Z(n21019) );
  XNOR U29616 ( .A(y[5417]), .B(x[5417]), .Z(n21018) );
  NAND U29617 ( .A(n21083), .B(n21084), .Z(N63521) );
  NANDN U29618 ( .A(n21085), .B(n21086), .Z(n21084) );
  OR U29619 ( .A(n21087), .B(n21088), .Z(n21086) );
  NAND U29620 ( .A(n21087), .B(n21088), .Z(n21083) );
  XOR U29621 ( .A(n21087), .B(n21089), .Z(N63520) );
  XNOR U29622 ( .A(n21085), .B(n21088), .Z(n21089) );
  AND U29623 ( .A(n21090), .B(n21091), .Z(n21088) );
  NANDN U29624 ( .A(n21092), .B(n21093), .Z(n21091) );
  NANDN U29625 ( .A(n21094), .B(n21095), .Z(n21093) );
  NANDN U29626 ( .A(n21095), .B(n21094), .Z(n21090) );
  NAND U29627 ( .A(n21096), .B(n21097), .Z(n21085) );
  NANDN U29628 ( .A(n21098), .B(n21099), .Z(n21097) );
  OR U29629 ( .A(n21100), .B(n21101), .Z(n21099) );
  NAND U29630 ( .A(n21101), .B(n21100), .Z(n21096) );
  AND U29631 ( .A(n21102), .B(n21103), .Z(n21087) );
  NANDN U29632 ( .A(n21104), .B(n21105), .Z(n21103) );
  NANDN U29633 ( .A(n21106), .B(n21107), .Z(n21105) );
  NANDN U29634 ( .A(n21107), .B(n21106), .Z(n21102) );
  XOR U29635 ( .A(n21101), .B(n21108), .Z(N63519) );
  XOR U29636 ( .A(n21098), .B(n21100), .Z(n21108) );
  XNOR U29637 ( .A(n21094), .B(n21109), .Z(n21100) );
  XNOR U29638 ( .A(n21092), .B(n21095), .Z(n21109) );
  NAND U29639 ( .A(n21110), .B(n21111), .Z(n21095) );
  NAND U29640 ( .A(n21112), .B(n21113), .Z(n21111) );
  OR U29641 ( .A(n21114), .B(n21115), .Z(n21112) );
  NANDN U29642 ( .A(n21116), .B(n21114), .Z(n21110) );
  IV U29643 ( .A(n21115), .Z(n21116) );
  NAND U29644 ( .A(n21117), .B(n21118), .Z(n21092) );
  NAND U29645 ( .A(n21119), .B(n21120), .Z(n21118) );
  NANDN U29646 ( .A(n21121), .B(n21122), .Z(n21119) );
  NANDN U29647 ( .A(n21122), .B(n21121), .Z(n21117) );
  AND U29648 ( .A(n21123), .B(n21124), .Z(n21094) );
  NAND U29649 ( .A(n21125), .B(n21126), .Z(n21124) );
  OR U29650 ( .A(n21127), .B(n21128), .Z(n21125) );
  NANDN U29651 ( .A(n21129), .B(n21127), .Z(n21123) );
  NAND U29652 ( .A(n21130), .B(n21131), .Z(n21098) );
  NANDN U29653 ( .A(n21132), .B(n21133), .Z(n21131) );
  OR U29654 ( .A(n21134), .B(n21135), .Z(n21133) );
  NANDN U29655 ( .A(n21136), .B(n21134), .Z(n21130) );
  IV U29656 ( .A(n21135), .Z(n21136) );
  XNOR U29657 ( .A(n21106), .B(n21137), .Z(n21101) );
  XNOR U29658 ( .A(n21104), .B(n21107), .Z(n21137) );
  NAND U29659 ( .A(n21138), .B(n21139), .Z(n21107) );
  NAND U29660 ( .A(n21140), .B(n21141), .Z(n21139) );
  OR U29661 ( .A(n21142), .B(n21143), .Z(n21140) );
  NANDN U29662 ( .A(n21144), .B(n21142), .Z(n21138) );
  IV U29663 ( .A(n21143), .Z(n21144) );
  NAND U29664 ( .A(n21145), .B(n21146), .Z(n21104) );
  NAND U29665 ( .A(n21147), .B(n21148), .Z(n21146) );
  NANDN U29666 ( .A(n21149), .B(n21150), .Z(n21147) );
  NANDN U29667 ( .A(n21150), .B(n21149), .Z(n21145) );
  AND U29668 ( .A(n21151), .B(n21152), .Z(n21106) );
  NAND U29669 ( .A(n21153), .B(n21154), .Z(n21152) );
  OR U29670 ( .A(n21155), .B(n21156), .Z(n21153) );
  NANDN U29671 ( .A(n21157), .B(n21155), .Z(n21151) );
  XNOR U29672 ( .A(n21132), .B(n21158), .Z(N63518) );
  XOR U29673 ( .A(n21134), .B(n21135), .Z(n21158) );
  XNOR U29674 ( .A(n21148), .B(n21159), .Z(n21135) );
  XOR U29675 ( .A(n21149), .B(n21150), .Z(n21159) );
  XOR U29676 ( .A(n21155), .B(n21160), .Z(n21150) );
  XOR U29677 ( .A(n21154), .B(n21157), .Z(n21160) );
  IV U29678 ( .A(n21156), .Z(n21157) );
  NAND U29679 ( .A(n21161), .B(n21162), .Z(n21156) );
  OR U29680 ( .A(n21163), .B(n21164), .Z(n21162) );
  OR U29681 ( .A(n21165), .B(n21166), .Z(n21161) );
  NAND U29682 ( .A(n21167), .B(n21168), .Z(n21154) );
  OR U29683 ( .A(n21169), .B(n21170), .Z(n21168) );
  OR U29684 ( .A(n21171), .B(n21172), .Z(n21167) );
  NOR U29685 ( .A(n21173), .B(n21174), .Z(n21155) );
  ANDN U29686 ( .B(n21175), .A(n21176), .Z(n21149) );
  XNOR U29687 ( .A(n21142), .B(n21177), .Z(n21148) );
  XNOR U29688 ( .A(n21141), .B(n21143), .Z(n21177) );
  NAND U29689 ( .A(n21178), .B(n21179), .Z(n21143) );
  OR U29690 ( .A(n21180), .B(n21181), .Z(n21179) );
  OR U29691 ( .A(n21182), .B(n21183), .Z(n21178) );
  NAND U29692 ( .A(n21184), .B(n21185), .Z(n21141) );
  OR U29693 ( .A(n21186), .B(n21187), .Z(n21185) );
  OR U29694 ( .A(n21188), .B(n21189), .Z(n21184) );
  ANDN U29695 ( .B(n21190), .A(n21191), .Z(n21142) );
  IV U29696 ( .A(n21192), .Z(n21190) );
  ANDN U29697 ( .B(n21193), .A(n21194), .Z(n21134) );
  XOR U29698 ( .A(n21120), .B(n21195), .Z(n21132) );
  XOR U29699 ( .A(n21121), .B(n21122), .Z(n21195) );
  XOR U29700 ( .A(n21127), .B(n21196), .Z(n21122) );
  XOR U29701 ( .A(n21126), .B(n21129), .Z(n21196) );
  IV U29702 ( .A(n21128), .Z(n21129) );
  NAND U29703 ( .A(n21197), .B(n21198), .Z(n21128) );
  OR U29704 ( .A(n21199), .B(n21200), .Z(n21198) );
  OR U29705 ( .A(n21201), .B(n21202), .Z(n21197) );
  NAND U29706 ( .A(n21203), .B(n21204), .Z(n21126) );
  OR U29707 ( .A(n21205), .B(n21206), .Z(n21204) );
  OR U29708 ( .A(n21207), .B(n21208), .Z(n21203) );
  NOR U29709 ( .A(n21209), .B(n21210), .Z(n21127) );
  ANDN U29710 ( .B(n21211), .A(n21212), .Z(n21121) );
  IV U29711 ( .A(n21213), .Z(n21211) );
  XNOR U29712 ( .A(n21114), .B(n21214), .Z(n21120) );
  XNOR U29713 ( .A(n21113), .B(n21115), .Z(n21214) );
  NAND U29714 ( .A(n21215), .B(n21216), .Z(n21115) );
  OR U29715 ( .A(n21217), .B(n21218), .Z(n21216) );
  OR U29716 ( .A(n21219), .B(n21220), .Z(n21215) );
  NAND U29717 ( .A(n21221), .B(n21222), .Z(n21113) );
  OR U29718 ( .A(n21223), .B(n21224), .Z(n21222) );
  OR U29719 ( .A(n21225), .B(n21226), .Z(n21221) );
  ANDN U29720 ( .B(n21227), .A(n21228), .Z(n21114) );
  IV U29721 ( .A(n21229), .Z(n21227) );
  XNOR U29722 ( .A(n21194), .B(n21193), .Z(N63517) );
  XOR U29723 ( .A(n21213), .B(n21212), .Z(n21193) );
  XNOR U29724 ( .A(n21228), .B(n21229), .Z(n21212) );
  XNOR U29725 ( .A(n21223), .B(n21224), .Z(n21229) );
  XNOR U29726 ( .A(n21225), .B(n21226), .Z(n21224) );
  XNOR U29727 ( .A(y[5413]), .B(x[5413]), .Z(n21226) );
  XNOR U29728 ( .A(y[5414]), .B(x[5414]), .Z(n21225) );
  XNOR U29729 ( .A(y[5412]), .B(x[5412]), .Z(n21223) );
  XNOR U29730 ( .A(n21217), .B(n21218), .Z(n21228) );
  XNOR U29731 ( .A(y[5409]), .B(x[5409]), .Z(n21218) );
  XNOR U29732 ( .A(n21219), .B(n21220), .Z(n21217) );
  XNOR U29733 ( .A(y[5410]), .B(x[5410]), .Z(n21220) );
  XNOR U29734 ( .A(y[5411]), .B(x[5411]), .Z(n21219) );
  XNOR U29735 ( .A(n21210), .B(n21209), .Z(n21213) );
  XNOR U29736 ( .A(n21205), .B(n21206), .Z(n21209) );
  XNOR U29737 ( .A(y[5406]), .B(x[5406]), .Z(n21206) );
  XNOR U29738 ( .A(n21207), .B(n21208), .Z(n21205) );
  XNOR U29739 ( .A(y[5407]), .B(x[5407]), .Z(n21208) );
  XNOR U29740 ( .A(y[5408]), .B(x[5408]), .Z(n21207) );
  XNOR U29741 ( .A(n21199), .B(n21200), .Z(n21210) );
  XNOR U29742 ( .A(y[5403]), .B(x[5403]), .Z(n21200) );
  XNOR U29743 ( .A(n21201), .B(n21202), .Z(n21199) );
  XNOR U29744 ( .A(y[5404]), .B(x[5404]), .Z(n21202) );
  XNOR U29745 ( .A(y[5405]), .B(x[5405]), .Z(n21201) );
  XOR U29746 ( .A(n21175), .B(n21176), .Z(n21194) );
  XNOR U29747 ( .A(n21191), .B(n21192), .Z(n21176) );
  XNOR U29748 ( .A(n21186), .B(n21187), .Z(n21192) );
  XNOR U29749 ( .A(n21188), .B(n21189), .Z(n21187) );
  XNOR U29750 ( .A(y[5401]), .B(x[5401]), .Z(n21189) );
  XNOR U29751 ( .A(y[5402]), .B(x[5402]), .Z(n21188) );
  XNOR U29752 ( .A(y[5400]), .B(x[5400]), .Z(n21186) );
  XNOR U29753 ( .A(n21180), .B(n21181), .Z(n21191) );
  XNOR U29754 ( .A(y[5397]), .B(x[5397]), .Z(n21181) );
  XNOR U29755 ( .A(n21182), .B(n21183), .Z(n21180) );
  XNOR U29756 ( .A(y[5398]), .B(x[5398]), .Z(n21183) );
  XNOR U29757 ( .A(y[5399]), .B(x[5399]), .Z(n21182) );
  XOR U29758 ( .A(n21174), .B(n21173), .Z(n21175) );
  XNOR U29759 ( .A(n21169), .B(n21170), .Z(n21173) );
  XNOR U29760 ( .A(y[5394]), .B(x[5394]), .Z(n21170) );
  XNOR U29761 ( .A(n21171), .B(n21172), .Z(n21169) );
  XNOR U29762 ( .A(y[5395]), .B(x[5395]), .Z(n21172) );
  XNOR U29763 ( .A(y[5396]), .B(x[5396]), .Z(n21171) );
  XNOR U29764 ( .A(n21163), .B(n21164), .Z(n21174) );
  XNOR U29765 ( .A(y[5391]), .B(x[5391]), .Z(n21164) );
  XNOR U29766 ( .A(n21165), .B(n21166), .Z(n21163) );
  XNOR U29767 ( .A(y[5392]), .B(x[5392]), .Z(n21166) );
  XNOR U29768 ( .A(y[5393]), .B(x[5393]), .Z(n21165) );
  NAND U29769 ( .A(n21230), .B(n21231), .Z(N63508) );
  NANDN U29770 ( .A(n21232), .B(n21233), .Z(n21231) );
  OR U29771 ( .A(n21234), .B(n21235), .Z(n21233) );
  NAND U29772 ( .A(n21234), .B(n21235), .Z(n21230) );
  XOR U29773 ( .A(n21234), .B(n21236), .Z(N63507) );
  XNOR U29774 ( .A(n21232), .B(n21235), .Z(n21236) );
  AND U29775 ( .A(n21237), .B(n21238), .Z(n21235) );
  NANDN U29776 ( .A(n21239), .B(n21240), .Z(n21238) );
  NANDN U29777 ( .A(n21241), .B(n21242), .Z(n21240) );
  NANDN U29778 ( .A(n21242), .B(n21241), .Z(n21237) );
  NAND U29779 ( .A(n21243), .B(n21244), .Z(n21232) );
  NANDN U29780 ( .A(n21245), .B(n21246), .Z(n21244) );
  OR U29781 ( .A(n21247), .B(n21248), .Z(n21246) );
  NAND U29782 ( .A(n21248), .B(n21247), .Z(n21243) );
  AND U29783 ( .A(n21249), .B(n21250), .Z(n21234) );
  NANDN U29784 ( .A(n21251), .B(n21252), .Z(n21250) );
  NANDN U29785 ( .A(n21253), .B(n21254), .Z(n21252) );
  NANDN U29786 ( .A(n21254), .B(n21253), .Z(n21249) );
  XOR U29787 ( .A(n21248), .B(n21255), .Z(N63506) );
  XOR U29788 ( .A(n21245), .B(n21247), .Z(n21255) );
  XNOR U29789 ( .A(n21241), .B(n21256), .Z(n21247) );
  XNOR U29790 ( .A(n21239), .B(n21242), .Z(n21256) );
  NAND U29791 ( .A(n21257), .B(n21258), .Z(n21242) );
  NAND U29792 ( .A(n21259), .B(n21260), .Z(n21258) );
  OR U29793 ( .A(n21261), .B(n21262), .Z(n21259) );
  NANDN U29794 ( .A(n21263), .B(n21261), .Z(n21257) );
  IV U29795 ( .A(n21262), .Z(n21263) );
  NAND U29796 ( .A(n21264), .B(n21265), .Z(n21239) );
  NAND U29797 ( .A(n21266), .B(n21267), .Z(n21265) );
  NANDN U29798 ( .A(n21268), .B(n21269), .Z(n21266) );
  NANDN U29799 ( .A(n21269), .B(n21268), .Z(n21264) );
  AND U29800 ( .A(n21270), .B(n21271), .Z(n21241) );
  NAND U29801 ( .A(n21272), .B(n21273), .Z(n21271) );
  OR U29802 ( .A(n21274), .B(n21275), .Z(n21272) );
  NANDN U29803 ( .A(n21276), .B(n21274), .Z(n21270) );
  NAND U29804 ( .A(n21277), .B(n21278), .Z(n21245) );
  NANDN U29805 ( .A(n21279), .B(n21280), .Z(n21278) );
  OR U29806 ( .A(n21281), .B(n21282), .Z(n21280) );
  NANDN U29807 ( .A(n21283), .B(n21281), .Z(n21277) );
  IV U29808 ( .A(n21282), .Z(n21283) );
  XNOR U29809 ( .A(n21253), .B(n21284), .Z(n21248) );
  XNOR U29810 ( .A(n21251), .B(n21254), .Z(n21284) );
  NAND U29811 ( .A(n21285), .B(n21286), .Z(n21254) );
  NAND U29812 ( .A(n21287), .B(n21288), .Z(n21286) );
  OR U29813 ( .A(n21289), .B(n21290), .Z(n21287) );
  NANDN U29814 ( .A(n21291), .B(n21289), .Z(n21285) );
  IV U29815 ( .A(n21290), .Z(n21291) );
  NAND U29816 ( .A(n21292), .B(n21293), .Z(n21251) );
  NAND U29817 ( .A(n21294), .B(n21295), .Z(n21293) );
  NANDN U29818 ( .A(n21296), .B(n21297), .Z(n21294) );
  NANDN U29819 ( .A(n21297), .B(n21296), .Z(n21292) );
  AND U29820 ( .A(n21298), .B(n21299), .Z(n21253) );
  NAND U29821 ( .A(n21300), .B(n21301), .Z(n21299) );
  OR U29822 ( .A(n21302), .B(n21303), .Z(n21300) );
  NANDN U29823 ( .A(n21304), .B(n21302), .Z(n21298) );
  XNOR U29824 ( .A(n21279), .B(n21305), .Z(N63505) );
  XOR U29825 ( .A(n21281), .B(n21282), .Z(n21305) );
  XNOR U29826 ( .A(n21295), .B(n21306), .Z(n21282) );
  XOR U29827 ( .A(n21296), .B(n21297), .Z(n21306) );
  XOR U29828 ( .A(n21302), .B(n21307), .Z(n21297) );
  XOR U29829 ( .A(n21301), .B(n21304), .Z(n21307) );
  IV U29830 ( .A(n21303), .Z(n21304) );
  NAND U29831 ( .A(n21308), .B(n21309), .Z(n21303) );
  OR U29832 ( .A(n21310), .B(n21311), .Z(n21309) );
  OR U29833 ( .A(n21312), .B(n21313), .Z(n21308) );
  NAND U29834 ( .A(n21314), .B(n21315), .Z(n21301) );
  OR U29835 ( .A(n21316), .B(n21317), .Z(n21315) );
  OR U29836 ( .A(n21318), .B(n21319), .Z(n21314) );
  NOR U29837 ( .A(n21320), .B(n21321), .Z(n21302) );
  ANDN U29838 ( .B(n21322), .A(n21323), .Z(n21296) );
  XNOR U29839 ( .A(n21289), .B(n21324), .Z(n21295) );
  XNOR U29840 ( .A(n21288), .B(n21290), .Z(n21324) );
  NAND U29841 ( .A(n21325), .B(n21326), .Z(n21290) );
  OR U29842 ( .A(n21327), .B(n21328), .Z(n21326) );
  OR U29843 ( .A(n21329), .B(n21330), .Z(n21325) );
  NAND U29844 ( .A(n21331), .B(n21332), .Z(n21288) );
  OR U29845 ( .A(n21333), .B(n21334), .Z(n21332) );
  OR U29846 ( .A(n21335), .B(n21336), .Z(n21331) );
  ANDN U29847 ( .B(n21337), .A(n21338), .Z(n21289) );
  IV U29848 ( .A(n21339), .Z(n21337) );
  ANDN U29849 ( .B(n21340), .A(n21341), .Z(n21281) );
  XOR U29850 ( .A(n21267), .B(n21342), .Z(n21279) );
  XOR U29851 ( .A(n21268), .B(n21269), .Z(n21342) );
  XOR U29852 ( .A(n21274), .B(n21343), .Z(n21269) );
  XOR U29853 ( .A(n21273), .B(n21276), .Z(n21343) );
  IV U29854 ( .A(n21275), .Z(n21276) );
  NAND U29855 ( .A(n21344), .B(n21345), .Z(n21275) );
  OR U29856 ( .A(n21346), .B(n21347), .Z(n21345) );
  OR U29857 ( .A(n21348), .B(n21349), .Z(n21344) );
  NAND U29858 ( .A(n21350), .B(n21351), .Z(n21273) );
  OR U29859 ( .A(n21352), .B(n21353), .Z(n21351) );
  OR U29860 ( .A(n21354), .B(n21355), .Z(n21350) );
  NOR U29861 ( .A(n21356), .B(n21357), .Z(n21274) );
  ANDN U29862 ( .B(n21358), .A(n21359), .Z(n21268) );
  IV U29863 ( .A(n21360), .Z(n21358) );
  XNOR U29864 ( .A(n21261), .B(n21361), .Z(n21267) );
  XNOR U29865 ( .A(n21260), .B(n21262), .Z(n21361) );
  NAND U29866 ( .A(n21362), .B(n21363), .Z(n21262) );
  OR U29867 ( .A(n21364), .B(n21365), .Z(n21363) );
  OR U29868 ( .A(n21366), .B(n21367), .Z(n21362) );
  NAND U29869 ( .A(n21368), .B(n21369), .Z(n21260) );
  OR U29870 ( .A(n21370), .B(n21371), .Z(n21369) );
  OR U29871 ( .A(n21372), .B(n21373), .Z(n21368) );
  ANDN U29872 ( .B(n21374), .A(n21375), .Z(n21261) );
  IV U29873 ( .A(n21376), .Z(n21374) );
  XNOR U29874 ( .A(n21341), .B(n21340), .Z(N63504) );
  XOR U29875 ( .A(n21360), .B(n21359), .Z(n21340) );
  XNOR U29876 ( .A(n21375), .B(n21376), .Z(n21359) );
  XNOR U29877 ( .A(n21370), .B(n21371), .Z(n21376) );
  XNOR U29878 ( .A(n21372), .B(n21373), .Z(n21371) );
  XNOR U29879 ( .A(y[5389]), .B(x[5389]), .Z(n21373) );
  XNOR U29880 ( .A(y[5390]), .B(x[5390]), .Z(n21372) );
  XNOR U29881 ( .A(y[5388]), .B(x[5388]), .Z(n21370) );
  XNOR U29882 ( .A(n21364), .B(n21365), .Z(n21375) );
  XNOR U29883 ( .A(y[5385]), .B(x[5385]), .Z(n21365) );
  XNOR U29884 ( .A(n21366), .B(n21367), .Z(n21364) );
  XNOR U29885 ( .A(y[5386]), .B(x[5386]), .Z(n21367) );
  XNOR U29886 ( .A(y[5387]), .B(x[5387]), .Z(n21366) );
  XNOR U29887 ( .A(n21357), .B(n21356), .Z(n21360) );
  XNOR U29888 ( .A(n21352), .B(n21353), .Z(n21356) );
  XNOR U29889 ( .A(y[5382]), .B(x[5382]), .Z(n21353) );
  XNOR U29890 ( .A(n21354), .B(n21355), .Z(n21352) );
  XNOR U29891 ( .A(y[5383]), .B(x[5383]), .Z(n21355) );
  XNOR U29892 ( .A(y[5384]), .B(x[5384]), .Z(n21354) );
  XNOR U29893 ( .A(n21346), .B(n21347), .Z(n21357) );
  XNOR U29894 ( .A(y[5379]), .B(x[5379]), .Z(n21347) );
  XNOR U29895 ( .A(n21348), .B(n21349), .Z(n21346) );
  XNOR U29896 ( .A(y[5380]), .B(x[5380]), .Z(n21349) );
  XNOR U29897 ( .A(y[5381]), .B(x[5381]), .Z(n21348) );
  XOR U29898 ( .A(n21322), .B(n21323), .Z(n21341) );
  XNOR U29899 ( .A(n21338), .B(n21339), .Z(n21323) );
  XNOR U29900 ( .A(n21333), .B(n21334), .Z(n21339) );
  XNOR U29901 ( .A(n21335), .B(n21336), .Z(n21334) );
  XNOR U29902 ( .A(y[5377]), .B(x[5377]), .Z(n21336) );
  XNOR U29903 ( .A(y[5378]), .B(x[5378]), .Z(n21335) );
  XNOR U29904 ( .A(y[5376]), .B(x[5376]), .Z(n21333) );
  XNOR U29905 ( .A(n21327), .B(n21328), .Z(n21338) );
  XNOR U29906 ( .A(y[5373]), .B(x[5373]), .Z(n21328) );
  XNOR U29907 ( .A(n21329), .B(n21330), .Z(n21327) );
  XNOR U29908 ( .A(y[5374]), .B(x[5374]), .Z(n21330) );
  XNOR U29909 ( .A(y[5375]), .B(x[5375]), .Z(n21329) );
  XOR U29910 ( .A(n21321), .B(n21320), .Z(n21322) );
  XNOR U29911 ( .A(n21316), .B(n21317), .Z(n21320) );
  XNOR U29912 ( .A(y[5370]), .B(x[5370]), .Z(n21317) );
  XNOR U29913 ( .A(n21318), .B(n21319), .Z(n21316) );
  XNOR U29914 ( .A(y[5371]), .B(x[5371]), .Z(n21319) );
  XNOR U29915 ( .A(y[5372]), .B(x[5372]), .Z(n21318) );
  XNOR U29916 ( .A(n21310), .B(n21311), .Z(n21321) );
  XNOR U29917 ( .A(y[5367]), .B(x[5367]), .Z(n21311) );
  XNOR U29918 ( .A(n21312), .B(n21313), .Z(n21310) );
  XNOR U29919 ( .A(y[5368]), .B(x[5368]), .Z(n21313) );
  XNOR U29920 ( .A(y[5369]), .B(x[5369]), .Z(n21312) );
  NAND U29921 ( .A(n21377), .B(n21378), .Z(N63495) );
  NANDN U29922 ( .A(n21379), .B(n21380), .Z(n21378) );
  OR U29923 ( .A(n21381), .B(n21382), .Z(n21380) );
  NAND U29924 ( .A(n21381), .B(n21382), .Z(n21377) );
  XOR U29925 ( .A(n21381), .B(n21383), .Z(N63494) );
  XNOR U29926 ( .A(n21379), .B(n21382), .Z(n21383) );
  AND U29927 ( .A(n21384), .B(n21385), .Z(n21382) );
  NANDN U29928 ( .A(n21386), .B(n21387), .Z(n21385) );
  NANDN U29929 ( .A(n21388), .B(n21389), .Z(n21387) );
  NANDN U29930 ( .A(n21389), .B(n21388), .Z(n21384) );
  NAND U29931 ( .A(n21390), .B(n21391), .Z(n21379) );
  NANDN U29932 ( .A(n21392), .B(n21393), .Z(n21391) );
  OR U29933 ( .A(n21394), .B(n21395), .Z(n21393) );
  NAND U29934 ( .A(n21395), .B(n21394), .Z(n21390) );
  AND U29935 ( .A(n21396), .B(n21397), .Z(n21381) );
  NANDN U29936 ( .A(n21398), .B(n21399), .Z(n21397) );
  NANDN U29937 ( .A(n21400), .B(n21401), .Z(n21399) );
  NANDN U29938 ( .A(n21401), .B(n21400), .Z(n21396) );
  XOR U29939 ( .A(n21395), .B(n21402), .Z(N63493) );
  XOR U29940 ( .A(n21392), .B(n21394), .Z(n21402) );
  XNOR U29941 ( .A(n21388), .B(n21403), .Z(n21394) );
  XNOR U29942 ( .A(n21386), .B(n21389), .Z(n21403) );
  NAND U29943 ( .A(n21404), .B(n21405), .Z(n21389) );
  NAND U29944 ( .A(n21406), .B(n21407), .Z(n21405) );
  OR U29945 ( .A(n21408), .B(n21409), .Z(n21406) );
  NANDN U29946 ( .A(n21410), .B(n21408), .Z(n21404) );
  IV U29947 ( .A(n21409), .Z(n21410) );
  NAND U29948 ( .A(n21411), .B(n21412), .Z(n21386) );
  NAND U29949 ( .A(n21413), .B(n21414), .Z(n21412) );
  NANDN U29950 ( .A(n21415), .B(n21416), .Z(n21413) );
  NANDN U29951 ( .A(n21416), .B(n21415), .Z(n21411) );
  AND U29952 ( .A(n21417), .B(n21418), .Z(n21388) );
  NAND U29953 ( .A(n21419), .B(n21420), .Z(n21418) );
  OR U29954 ( .A(n21421), .B(n21422), .Z(n21419) );
  NANDN U29955 ( .A(n21423), .B(n21421), .Z(n21417) );
  NAND U29956 ( .A(n21424), .B(n21425), .Z(n21392) );
  NANDN U29957 ( .A(n21426), .B(n21427), .Z(n21425) );
  OR U29958 ( .A(n21428), .B(n21429), .Z(n21427) );
  NANDN U29959 ( .A(n21430), .B(n21428), .Z(n21424) );
  IV U29960 ( .A(n21429), .Z(n21430) );
  XNOR U29961 ( .A(n21400), .B(n21431), .Z(n21395) );
  XNOR U29962 ( .A(n21398), .B(n21401), .Z(n21431) );
  NAND U29963 ( .A(n21432), .B(n21433), .Z(n21401) );
  NAND U29964 ( .A(n21434), .B(n21435), .Z(n21433) );
  OR U29965 ( .A(n21436), .B(n21437), .Z(n21434) );
  NANDN U29966 ( .A(n21438), .B(n21436), .Z(n21432) );
  IV U29967 ( .A(n21437), .Z(n21438) );
  NAND U29968 ( .A(n21439), .B(n21440), .Z(n21398) );
  NAND U29969 ( .A(n21441), .B(n21442), .Z(n21440) );
  NANDN U29970 ( .A(n21443), .B(n21444), .Z(n21441) );
  NANDN U29971 ( .A(n21444), .B(n21443), .Z(n21439) );
  AND U29972 ( .A(n21445), .B(n21446), .Z(n21400) );
  NAND U29973 ( .A(n21447), .B(n21448), .Z(n21446) );
  OR U29974 ( .A(n21449), .B(n21450), .Z(n21447) );
  NANDN U29975 ( .A(n21451), .B(n21449), .Z(n21445) );
  XNOR U29976 ( .A(n21426), .B(n21452), .Z(N63492) );
  XOR U29977 ( .A(n21428), .B(n21429), .Z(n21452) );
  XNOR U29978 ( .A(n21442), .B(n21453), .Z(n21429) );
  XOR U29979 ( .A(n21443), .B(n21444), .Z(n21453) );
  XOR U29980 ( .A(n21449), .B(n21454), .Z(n21444) );
  XOR U29981 ( .A(n21448), .B(n21451), .Z(n21454) );
  IV U29982 ( .A(n21450), .Z(n21451) );
  NAND U29983 ( .A(n21455), .B(n21456), .Z(n21450) );
  OR U29984 ( .A(n21457), .B(n21458), .Z(n21456) );
  OR U29985 ( .A(n21459), .B(n21460), .Z(n21455) );
  NAND U29986 ( .A(n21461), .B(n21462), .Z(n21448) );
  OR U29987 ( .A(n21463), .B(n21464), .Z(n21462) );
  OR U29988 ( .A(n21465), .B(n21466), .Z(n21461) );
  NOR U29989 ( .A(n21467), .B(n21468), .Z(n21449) );
  ANDN U29990 ( .B(n21469), .A(n21470), .Z(n21443) );
  XNOR U29991 ( .A(n21436), .B(n21471), .Z(n21442) );
  XNOR U29992 ( .A(n21435), .B(n21437), .Z(n21471) );
  NAND U29993 ( .A(n21472), .B(n21473), .Z(n21437) );
  OR U29994 ( .A(n21474), .B(n21475), .Z(n21473) );
  OR U29995 ( .A(n21476), .B(n21477), .Z(n21472) );
  NAND U29996 ( .A(n21478), .B(n21479), .Z(n21435) );
  OR U29997 ( .A(n21480), .B(n21481), .Z(n21479) );
  OR U29998 ( .A(n21482), .B(n21483), .Z(n21478) );
  ANDN U29999 ( .B(n21484), .A(n21485), .Z(n21436) );
  IV U30000 ( .A(n21486), .Z(n21484) );
  ANDN U30001 ( .B(n21487), .A(n21488), .Z(n21428) );
  XOR U30002 ( .A(n21414), .B(n21489), .Z(n21426) );
  XOR U30003 ( .A(n21415), .B(n21416), .Z(n21489) );
  XOR U30004 ( .A(n21421), .B(n21490), .Z(n21416) );
  XOR U30005 ( .A(n21420), .B(n21423), .Z(n21490) );
  IV U30006 ( .A(n21422), .Z(n21423) );
  NAND U30007 ( .A(n21491), .B(n21492), .Z(n21422) );
  OR U30008 ( .A(n21493), .B(n21494), .Z(n21492) );
  OR U30009 ( .A(n21495), .B(n21496), .Z(n21491) );
  NAND U30010 ( .A(n21497), .B(n21498), .Z(n21420) );
  OR U30011 ( .A(n21499), .B(n21500), .Z(n21498) );
  OR U30012 ( .A(n21501), .B(n21502), .Z(n21497) );
  NOR U30013 ( .A(n21503), .B(n21504), .Z(n21421) );
  ANDN U30014 ( .B(n21505), .A(n21506), .Z(n21415) );
  IV U30015 ( .A(n21507), .Z(n21505) );
  XNOR U30016 ( .A(n21408), .B(n21508), .Z(n21414) );
  XNOR U30017 ( .A(n21407), .B(n21409), .Z(n21508) );
  NAND U30018 ( .A(n21509), .B(n21510), .Z(n21409) );
  OR U30019 ( .A(n21511), .B(n21512), .Z(n21510) );
  OR U30020 ( .A(n21513), .B(n21514), .Z(n21509) );
  NAND U30021 ( .A(n21515), .B(n21516), .Z(n21407) );
  OR U30022 ( .A(n21517), .B(n21518), .Z(n21516) );
  OR U30023 ( .A(n21519), .B(n21520), .Z(n21515) );
  ANDN U30024 ( .B(n21521), .A(n21522), .Z(n21408) );
  IV U30025 ( .A(n21523), .Z(n21521) );
  XNOR U30026 ( .A(n21488), .B(n21487), .Z(N63491) );
  XOR U30027 ( .A(n21507), .B(n21506), .Z(n21487) );
  XNOR U30028 ( .A(n21522), .B(n21523), .Z(n21506) );
  XNOR U30029 ( .A(n21517), .B(n21518), .Z(n21523) );
  XNOR U30030 ( .A(n21519), .B(n21520), .Z(n21518) );
  XNOR U30031 ( .A(y[5365]), .B(x[5365]), .Z(n21520) );
  XNOR U30032 ( .A(y[5366]), .B(x[5366]), .Z(n21519) );
  XNOR U30033 ( .A(y[5364]), .B(x[5364]), .Z(n21517) );
  XNOR U30034 ( .A(n21511), .B(n21512), .Z(n21522) );
  XNOR U30035 ( .A(y[5361]), .B(x[5361]), .Z(n21512) );
  XNOR U30036 ( .A(n21513), .B(n21514), .Z(n21511) );
  XNOR U30037 ( .A(y[5362]), .B(x[5362]), .Z(n21514) );
  XNOR U30038 ( .A(y[5363]), .B(x[5363]), .Z(n21513) );
  XNOR U30039 ( .A(n21504), .B(n21503), .Z(n21507) );
  XNOR U30040 ( .A(n21499), .B(n21500), .Z(n21503) );
  XNOR U30041 ( .A(y[5358]), .B(x[5358]), .Z(n21500) );
  XNOR U30042 ( .A(n21501), .B(n21502), .Z(n21499) );
  XNOR U30043 ( .A(y[5359]), .B(x[5359]), .Z(n21502) );
  XNOR U30044 ( .A(y[5360]), .B(x[5360]), .Z(n21501) );
  XNOR U30045 ( .A(n21493), .B(n21494), .Z(n21504) );
  XNOR U30046 ( .A(y[5355]), .B(x[5355]), .Z(n21494) );
  XNOR U30047 ( .A(n21495), .B(n21496), .Z(n21493) );
  XNOR U30048 ( .A(y[5356]), .B(x[5356]), .Z(n21496) );
  XNOR U30049 ( .A(y[5357]), .B(x[5357]), .Z(n21495) );
  XOR U30050 ( .A(n21469), .B(n21470), .Z(n21488) );
  XNOR U30051 ( .A(n21485), .B(n21486), .Z(n21470) );
  XNOR U30052 ( .A(n21480), .B(n21481), .Z(n21486) );
  XNOR U30053 ( .A(n21482), .B(n21483), .Z(n21481) );
  XNOR U30054 ( .A(y[5353]), .B(x[5353]), .Z(n21483) );
  XNOR U30055 ( .A(y[5354]), .B(x[5354]), .Z(n21482) );
  XNOR U30056 ( .A(y[5352]), .B(x[5352]), .Z(n21480) );
  XNOR U30057 ( .A(n21474), .B(n21475), .Z(n21485) );
  XNOR U30058 ( .A(y[5349]), .B(x[5349]), .Z(n21475) );
  XNOR U30059 ( .A(n21476), .B(n21477), .Z(n21474) );
  XNOR U30060 ( .A(y[5350]), .B(x[5350]), .Z(n21477) );
  XNOR U30061 ( .A(y[5351]), .B(x[5351]), .Z(n21476) );
  XOR U30062 ( .A(n21468), .B(n21467), .Z(n21469) );
  XNOR U30063 ( .A(n21463), .B(n21464), .Z(n21467) );
  XNOR U30064 ( .A(y[5346]), .B(x[5346]), .Z(n21464) );
  XNOR U30065 ( .A(n21465), .B(n21466), .Z(n21463) );
  XNOR U30066 ( .A(y[5347]), .B(x[5347]), .Z(n21466) );
  XNOR U30067 ( .A(y[5348]), .B(x[5348]), .Z(n21465) );
  XNOR U30068 ( .A(n21457), .B(n21458), .Z(n21468) );
  XNOR U30069 ( .A(y[5343]), .B(x[5343]), .Z(n21458) );
  XNOR U30070 ( .A(n21459), .B(n21460), .Z(n21457) );
  XNOR U30071 ( .A(y[5344]), .B(x[5344]), .Z(n21460) );
  XNOR U30072 ( .A(y[5345]), .B(x[5345]), .Z(n21459) );
  NAND U30073 ( .A(n21524), .B(n21525), .Z(N63482) );
  NANDN U30074 ( .A(n21526), .B(n21527), .Z(n21525) );
  OR U30075 ( .A(n21528), .B(n21529), .Z(n21527) );
  NAND U30076 ( .A(n21528), .B(n21529), .Z(n21524) );
  XOR U30077 ( .A(n21528), .B(n21530), .Z(N63481) );
  XNOR U30078 ( .A(n21526), .B(n21529), .Z(n21530) );
  AND U30079 ( .A(n21531), .B(n21532), .Z(n21529) );
  NANDN U30080 ( .A(n21533), .B(n21534), .Z(n21532) );
  NANDN U30081 ( .A(n21535), .B(n21536), .Z(n21534) );
  NANDN U30082 ( .A(n21536), .B(n21535), .Z(n21531) );
  NAND U30083 ( .A(n21537), .B(n21538), .Z(n21526) );
  NANDN U30084 ( .A(n21539), .B(n21540), .Z(n21538) );
  OR U30085 ( .A(n21541), .B(n21542), .Z(n21540) );
  NAND U30086 ( .A(n21542), .B(n21541), .Z(n21537) );
  AND U30087 ( .A(n21543), .B(n21544), .Z(n21528) );
  NANDN U30088 ( .A(n21545), .B(n21546), .Z(n21544) );
  NANDN U30089 ( .A(n21547), .B(n21548), .Z(n21546) );
  NANDN U30090 ( .A(n21548), .B(n21547), .Z(n21543) );
  XOR U30091 ( .A(n21542), .B(n21549), .Z(N63480) );
  XOR U30092 ( .A(n21539), .B(n21541), .Z(n21549) );
  XNOR U30093 ( .A(n21535), .B(n21550), .Z(n21541) );
  XNOR U30094 ( .A(n21533), .B(n21536), .Z(n21550) );
  NAND U30095 ( .A(n21551), .B(n21552), .Z(n21536) );
  NAND U30096 ( .A(n21553), .B(n21554), .Z(n21552) );
  OR U30097 ( .A(n21555), .B(n21556), .Z(n21553) );
  NANDN U30098 ( .A(n21557), .B(n21555), .Z(n21551) );
  IV U30099 ( .A(n21556), .Z(n21557) );
  NAND U30100 ( .A(n21558), .B(n21559), .Z(n21533) );
  NAND U30101 ( .A(n21560), .B(n21561), .Z(n21559) );
  NANDN U30102 ( .A(n21562), .B(n21563), .Z(n21560) );
  NANDN U30103 ( .A(n21563), .B(n21562), .Z(n21558) );
  AND U30104 ( .A(n21564), .B(n21565), .Z(n21535) );
  NAND U30105 ( .A(n21566), .B(n21567), .Z(n21565) );
  OR U30106 ( .A(n21568), .B(n21569), .Z(n21566) );
  NANDN U30107 ( .A(n21570), .B(n21568), .Z(n21564) );
  NAND U30108 ( .A(n21571), .B(n21572), .Z(n21539) );
  NANDN U30109 ( .A(n21573), .B(n21574), .Z(n21572) );
  OR U30110 ( .A(n21575), .B(n21576), .Z(n21574) );
  NANDN U30111 ( .A(n21577), .B(n21575), .Z(n21571) );
  IV U30112 ( .A(n21576), .Z(n21577) );
  XNOR U30113 ( .A(n21547), .B(n21578), .Z(n21542) );
  XNOR U30114 ( .A(n21545), .B(n21548), .Z(n21578) );
  NAND U30115 ( .A(n21579), .B(n21580), .Z(n21548) );
  NAND U30116 ( .A(n21581), .B(n21582), .Z(n21580) );
  OR U30117 ( .A(n21583), .B(n21584), .Z(n21581) );
  NANDN U30118 ( .A(n21585), .B(n21583), .Z(n21579) );
  IV U30119 ( .A(n21584), .Z(n21585) );
  NAND U30120 ( .A(n21586), .B(n21587), .Z(n21545) );
  NAND U30121 ( .A(n21588), .B(n21589), .Z(n21587) );
  NANDN U30122 ( .A(n21590), .B(n21591), .Z(n21588) );
  NANDN U30123 ( .A(n21591), .B(n21590), .Z(n21586) );
  AND U30124 ( .A(n21592), .B(n21593), .Z(n21547) );
  NAND U30125 ( .A(n21594), .B(n21595), .Z(n21593) );
  OR U30126 ( .A(n21596), .B(n21597), .Z(n21594) );
  NANDN U30127 ( .A(n21598), .B(n21596), .Z(n21592) );
  XNOR U30128 ( .A(n21573), .B(n21599), .Z(N63479) );
  XOR U30129 ( .A(n21575), .B(n21576), .Z(n21599) );
  XNOR U30130 ( .A(n21589), .B(n21600), .Z(n21576) );
  XOR U30131 ( .A(n21590), .B(n21591), .Z(n21600) );
  XOR U30132 ( .A(n21596), .B(n21601), .Z(n21591) );
  XOR U30133 ( .A(n21595), .B(n21598), .Z(n21601) );
  IV U30134 ( .A(n21597), .Z(n21598) );
  NAND U30135 ( .A(n21602), .B(n21603), .Z(n21597) );
  OR U30136 ( .A(n21604), .B(n21605), .Z(n21603) );
  OR U30137 ( .A(n21606), .B(n21607), .Z(n21602) );
  NAND U30138 ( .A(n21608), .B(n21609), .Z(n21595) );
  OR U30139 ( .A(n21610), .B(n21611), .Z(n21609) );
  OR U30140 ( .A(n21612), .B(n21613), .Z(n21608) );
  NOR U30141 ( .A(n21614), .B(n21615), .Z(n21596) );
  ANDN U30142 ( .B(n21616), .A(n21617), .Z(n21590) );
  XNOR U30143 ( .A(n21583), .B(n21618), .Z(n21589) );
  XNOR U30144 ( .A(n21582), .B(n21584), .Z(n21618) );
  NAND U30145 ( .A(n21619), .B(n21620), .Z(n21584) );
  OR U30146 ( .A(n21621), .B(n21622), .Z(n21620) );
  OR U30147 ( .A(n21623), .B(n21624), .Z(n21619) );
  NAND U30148 ( .A(n21625), .B(n21626), .Z(n21582) );
  OR U30149 ( .A(n21627), .B(n21628), .Z(n21626) );
  OR U30150 ( .A(n21629), .B(n21630), .Z(n21625) );
  ANDN U30151 ( .B(n21631), .A(n21632), .Z(n21583) );
  IV U30152 ( .A(n21633), .Z(n21631) );
  ANDN U30153 ( .B(n21634), .A(n21635), .Z(n21575) );
  XOR U30154 ( .A(n21561), .B(n21636), .Z(n21573) );
  XOR U30155 ( .A(n21562), .B(n21563), .Z(n21636) );
  XOR U30156 ( .A(n21568), .B(n21637), .Z(n21563) );
  XOR U30157 ( .A(n21567), .B(n21570), .Z(n21637) );
  IV U30158 ( .A(n21569), .Z(n21570) );
  NAND U30159 ( .A(n21638), .B(n21639), .Z(n21569) );
  OR U30160 ( .A(n21640), .B(n21641), .Z(n21639) );
  OR U30161 ( .A(n21642), .B(n21643), .Z(n21638) );
  NAND U30162 ( .A(n21644), .B(n21645), .Z(n21567) );
  OR U30163 ( .A(n21646), .B(n21647), .Z(n21645) );
  OR U30164 ( .A(n21648), .B(n21649), .Z(n21644) );
  NOR U30165 ( .A(n21650), .B(n21651), .Z(n21568) );
  ANDN U30166 ( .B(n21652), .A(n21653), .Z(n21562) );
  IV U30167 ( .A(n21654), .Z(n21652) );
  XNOR U30168 ( .A(n21555), .B(n21655), .Z(n21561) );
  XNOR U30169 ( .A(n21554), .B(n21556), .Z(n21655) );
  NAND U30170 ( .A(n21656), .B(n21657), .Z(n21556) );
  OR U30171 ( .A(n21658), .B(n21659), .Z(n21657) );
  OR U30172 ( .A(n21660), .B(n21661), .Z(n21656) );
  NAND U30173 ( .A(n21662), .B(n21663), .Z(n21554) );
  OR U30174 ( .A(n21664), .B(n21665), .Z(n21663) );
  OR U30175 ( .A(n21666), .B(n21667), .Z(n21662) );
  ANDN U30176 ( .B(n21668), .A(n21669), .Z(n21555) );
  IV U30177 ( .A(n21670), .Z(n21668) );
  XNOR U30178 ( .A(n21635), .B(n21634), .Z(N63478) );
  XOR U30179 ( .A(n21654), .B(n21653), .Z(n21634) );
  XNOR U30180 ( .A(n21669), .B(n21670), .Z(n21653) );
  XNOR U30181 ( .A(n21664), .B(n21665), .Z(n21670) );
  XNOR U30182 ( .A(n21666), .B(n21667), .Z(n21665) );
  XNOR U30183 ( .A(y[5341]), .B(x[5341]), .Z(n21667) );
  XNOR U30184 ( .A(y[5342]), .B(x[5342]), .Z(n21666) );
  XNOR U30185 ( .A(y[5340]), .B(x[5340]), .Z(n21664) );
  XNOR U30186 ( .A(n21658), .B(n21659), .Z(n21669) );
  XNOR U30187 ( .A(y[5337]), .B(x[5337]), .Z(n21659) );
  XNOR U30188 ( .A(n21660), .B(n21661), .Z(n21658) );
  XNOR U30189 ( .A(y[5338]), .B(x[5338]), .Z(n21661) );
  XNOR U30190 ( .A(y[5339]), .B(x[5339]), .Z(n21660) );
  XNOR U30191 ( .A(n21651), .B(n21650), .Z(n21654) );
  XNOR U30192 ( .A(n21646), .B(n21647), .Z(n21650) );
  XNOR U30193 ( .A(y[5334]), .B(x[5334]), .Z(n21647) );
  XNOR U30194 ( .A(n21648), .B(n21649), .Z(n21646) );
  XNOR U30195 ( .A(y[5335]), .B(x[5335]), .Z(n21649) );
  XNOR U30196 ( .A(y[5336]), .B(x[5336]), .Z(n21648) );
  XNOR U30197 ( .A(n21640), .B(n21641), .Z(n21651) );
  XNOR U30198 ( .A(y[5331]), .B(x[5331]), .Z(n21641) );
  XNOR U30199 ( .A(n21642), .B(n21643), .Z(n21640) );
  XNOR U30200 ( .A(y[5332]), .B(x[5332]), .Z(n21643) );
  XNOR U30201 ( .A(y[5333]), .B(x[5333]), .Z(n21642) );
  XOR U30202 ( .A(n21616), .B(n21617), .Z(n21635) );
  XNOR U30203 ( .A(n21632), .B(n21633), .Z(n21617) );
  XNOR U30204 ( .A(n21627), .B(n21628), .Z(n21633) );
  XNOR U30205 ( .A(n21629), .B(n21630), .Z(n21628) );
  XNOR U30206 ( .A(y[5329]), .B(x[5329]), .Z(n21630) );
  XNOR U30207 ( .A(y[5330]), .B(x[5330]), .Z(n21629) );
  XNOR U30208 ( .A(y[5328]), .B(x[5328]), .Z(n21627) );
  XNOR U30209 ( .A(n21621), .B(n21622), .Z(n21632) );
  XNOR U30210 ( .A(y[5325]), .B(x[5325]), .Z(n21622) );
  XNOR U30211 ( .A(n21623), .B(n21624), .Z(n21621) );
  XNOR U30212 ( .A(y[5326]), .B(x[5326]), .Z(n21624) );
  XNOR U30213 ( .A(y[5327]), .B(x[5327]), .Z(n21623) );
  XOR U30214 ( .A(n21615), .B(n21614), .Z(n21616) );
  XNOR U30215 ( .A(n21610), .B(n21611), .Z(n21614) );
  XNOR U30216 ( .A(y[5322]), .B(x[5322]), .Z(n21611) );
  XNOR U30217 ( .A(n21612), .B(n21613), .Z(n21610) );
  XNOR U30218 ( .A(y[5323]), .B(x[5323]), .Z(n21613) );
  XNOR U30219 ( .A(y[5324]), .B(x[5324]), .Z(n21612) );
  XNOR U30220 ( .A(n21604), .B(n21605), .Z(n21615) );
  XNOR U30221 ( .A(y[5319]), .B(x[5319]), .Z(n21605) );
  XNOR U30222 ( .A(n21606), .B(n21607), .Z(n21604) );
  XNOR U30223 ( .A(y[5320]), .B(x[5320]), .Z(n21607) );
  XNOR U30224 ( .A(y[5321]), .B(x[5321]), .Z(n21606) );
  NAND U30225 ( .A(n21671), .B(n21672), .Z(N63469) );
  NANDN U30226 ( .A(n21673), .B(n21674), .Z(n21672) );
  OR U30227 ( .A(n21675), .B(n21676), .Z(n21674) );
  NAND U30228 ( .A(n21675), .B(n21676), .Z(n21671) );
  XOR U30229 ( .A(n21675), .B(n21677), .Z(N63468) );
  XNOR U30230 ( .A(n21673), .B(n21676), .Z(n21677) );
  AND U30231 ( .A(n21678), .B(n21679), .Z(n21676) );
  NANDN U30232 ( .A(n21680), .B(n21681), .Z(n21679) );
  NANDN U30233 ( .A(n21682), .B(n21683), .Z(n21681) );
  NANDN U30234 ( .A(n21683), .B(n21682), .Z(n21678) );
  NAND U30235 ( .A(n21684), .B(n21685), .Z(n21673) );
  NANDN U30236 ( .A(n21686), .B(n21687), .Z(n21685) );
  OR U30237 ( .A(n21688), .B(n21689), .Z(n21687) );
  NAND U30238 ( .A(n21689), .B(n21688), .Z(n21684) );
  AND U30239 ( .A(n21690), .B(n21691), .Z(n21675) );
  NANDN U30240 ( .A(n21692), .B(n21693), .Z(n21691) );
  NANDN U30241 ( .A(n21694), .B(n21695), .Z(n21693) );
  NANDN U30242 ( .A(n21695), .B(n21694), .Z(n21690) );
  XOR U30243 ( .A(n21689), .B(n21696), .Z(N63467) );
  XOR U30244 ( .A(n21686), .B(n21688), .Z(n21696) );
  XNOR U30245 ( .A(n21682), .B(n21697), .Z(n21688) );
  XNOR U30246 ( .A(n21680), .B(n21683), .Z(n21697) );
  NAND U30247 ( .A(n21698), .B(n21699), .Z(n21683) );
  NAND U30248 ( .A(n21700), .B(n21701), .Z(n21699) );
  OR U30249 ( .A(n21702), .B(n21703), .Z(n21700) );
  NANDN U30250 ( .A(n21704), .B(n21702), .Z(n21698) );
  IV U30251 ( .A(n21703), .Z(n21704) );
  NAND U30252 ( .A(n21705), .B(n21706), .Z(n21680) );
  NAND U30253 ( .A(n21707), .B(n21708), .Z(n21706) );
  NANDN U30254 ( .A(n21709), .B(n21710), .Z(n21707) );
  NANDN U30255 ( .A(n21710), .B(n21709), .Z(n21705) );
  AND U30256 ( .A(n21711), .B(n21712), .Z(n21682) );
  NAND U30257 ( .A(n21713), .B(n21714), .Z(n21712) );
  OR U30258 ( .A(n21715), .B(n21716), .Z(n21713) );
  NANDN U30259 ( .A(n21717), .B(n21715), .Z(n21711) );
  NAND U30260 ( .A(n21718), .B(n21719), .Z(n21686) );
  NANDN U30261 ( .A(n21720), .B(n21721), .Z(n21719) );
  OR U30262 ( .A(n21722), .B(n21723), .Z(n21721) );
  NANDN U30263 ( .A(n21724), .B(n21722), .Z(n21718) );
  IV U30264 ( .A(n21723), .Z(n21724) );
  XNOR U30265 ( .A(n21694), .B(n21725), .Z(n21689) );
  XNOR U30266 ( .A(n21692), .B(n21695), .Z(n21725) );
  NAND U30267 ( .A(n21726), .B(n21727), .Z(n21695) );
  NAND U30268 ( .A(n21728), .B(n21729), .Z(n21727) );
  OR U30269 ( .A(n21730), .B(n21731), .Z(n21728) );
  NANDN U30270 ( .A(n21732), .B(n21730), .Z(n21726) );
  IV U30271 ( .A(n21731), .Z(n21732) );
  NAND U30272 ( .A(n21733), .B(n21734), .Z(n21692) );
  NAND U30273 ( .A(n21735), .B(n21736), .Z(n21734) );
  NANDN U30274 ( .A(n21737), .B(n21738), .Z(n21735) );
  NANDN U30275 ( .A(n21738), .B(n21737), .Z(n21733) );
  AND U30276 ( .A(n21739), .B(n21740), .Z(n21694) );
  NAND U30277 ( .A(n21741), .B(n21742), .Z(n21740) );
  OR U30278 ( .A(n21743), .B(n21744), .Z(n21741) );
  NANDN U30279 ( .A(n21745), .B(n21743), .Z(n21739) );
  XNOR U30280 ( .A(n21720), .B(n21746), .Z(N63466) );
  XOR U30281 ( .A(n21722), .B(n21723), .Z(n21746) );
  XNOR U30282 ( .A(n21736), .B(n21747), .Z(n21723) );
  XOR U30283 ( .A(n21737), .B(n21738), .Z(n21747) );
  XOR U30284 ( .A(n21743), .B(n21748), .Z(n21738) );
  XOR U30285 ( .A(n21742), .B(n21745), .Z(n21748) );
  IV U30286 ( .A(n21744), .Z(n21745) );
  NAND U30287 ( .A(n21749), .B(n21750), .Z(n21744) );
  OR U30288 ( .A(n21751), .B(n21752), .Z(n21750) );
  OR U30289 ( .A(n21753), .B(n21754), .Z(n21749) );
  NAND U30290 ( .A(n21755), .B(n21756), .Z(n21742) );
  OR U30291 ( .A(n21757), .B(n21758), .Z(n21756) );
  OR U30292 ( .A(n21759), .B(n21760), .Z(n21755) );
  NOR U30293 ( .A(n21761), .B(n21762), .Z(n21743) );
  ANDN U30294 ( .B(n21763), .A(n21764), .Z(n21737) );
  XNOR U30295 ( .A(n21730), .B(n21765), .Z(n21736) );
  XNOR U30296 ( .A(n21729), .B(n21731), .Z(n21765) );
  NAND U30297 ( .A(n21766), .B(n21767), .Z(n21731) );
  OR U30298 ( .A(n21768), .B(n21769), .Z(n21767) );
  OR U30299 ( .A(n21770), .B(n21771), .Z(n21766) );
  NAND U30300 ( .A(n21772), .B(n21773), .Z(n21729) );
  OR U30301 ( .A(n21774), .B(n21775), .Z(n21773) );
  OR U30302 ( .A(n21776), .B(n21777), .Z(n21772) );
  ANDN U30303 ( .B(n21778), .A(n21779), .Z(n21730) );
  IV U30304 ( .A(n21780), .Z(n21778) );
  ANDN U30305 ( .B(n21781), .A(n21782), .Z(n21722) );
  XOR U30306 ( .A(n21708), .B(n21783), .Z(n21720) );
  XOR U30307 ( .A(n21709), .B(n21710), .Z(n21783) );
  XOR U30308 ( .A(n21715), .B(n21784), .Z(n21710) );
  XOR U30309 ( .A(n21714), .B(n21717), .Z(n21784) );
  IV U30310 ( .A(n21716), .Z(n21717) );
  NAND U30311 ( .A(n21785), .B(n21786), .Z(n21716) );
  OR U30312 ( .A(n21787), .B(n21788), .Z(n21786) );
  OR U30313 ( .A(n21789), .B(n21790), .Z(n21785) );
  NAND U30314 ( .A(n21791), .B(n21792), .Z(n21714) );
  OR U30315 ( .A(n21793), .B(n21794), .Z(n21792) );
  OR U30316 ( .A(n21795), .B(n21796), .Z(n21791) );
  NOR U30317 ( .A(n21797), .B(n21798), .Z(n21715) );
  ANDN U30318 ( .B(n21799), .A(n21800), .Z(n21709) );
  IV U30319 ( .A(n21801), .Z(n21799) );
  XNOR U30320 ( .A(n21702), .B(n21802), .Z(n21708) );
  XNOR U30321 ( .A(n21701), .B(n21703), .Z(n21802) );
  NAND U30322 ( .A(n21803), .B(n21804), .Z(n21703) );
  OR U30323 ( .A(n21805), .B(n21806), .Z(n21804) );
  OR U30324 ( .A(n21807), .B(n21808), .Z(n21803) );
  NAND U30325 ( .A(n21809), .B(n21810), .Z(n21701) );
  OR U30326 ( .A(n21811), .B(n21812), .Z(n21810) );
  OR U30327 ( .A(n21813), .B(n21814), .Z(n21809) );
  ANDN U30328 ( .B(n21815), .A(n21816), .Z(n21702) );
  IV U30329 ( .A(n21817), .Z(n21815) );
  XNOR U30330 ( .A(n21782), .B(n21781), .Z(N63465) );
  XOR U30331 ( .A(n21801), .B(n21800), .Z(n21781) );
  XNOR U30332 ( .A(n21816), .B(n21817), .Z(n21800) );
  XNOR U30333 ( .A(n21811), .B(n21812), .Z(n21817) );
  XNOR U30334 ( .A(n21813), .B(n21814), .Z(n21812) );
  XNOR U30335 ( .A(y[5317]), .B(x[5317]), .Z(n21814) );
  XNOR U30336 ( .A(y[5318]), .B(x[5318]), .Z(n21813) );
  XNOR U30337 ( .A(y[5316]), .B(x[5316]), .Z(n21811) );
  XNOR U30338 ( .A(n21805), .B(n21806), .Z(n21816) );
  XNOR U30339 ( .A(y[5313]), .B(x[5313]), .Z(n21806) );
  XNOR U30340 ( .A(n21807), .B(n21808), .Z(n21805) );
  XNOR U30341 ( .A(y[5314]), .B(x[5314]), .Z(n21808) );
  XNOR U30342 ( .A(y[5315]), .B(x[5315]), .Z(n21807) );
  XNOR U30343 ( .A(n21798), .B(n21797), .Z(n21801) );
  XNOR U30344 ( .A(n21793), .B(n21794), .Z(n21797) );
  XNOR U30345 ( .A(y[5310]), .B(x[5310]), .Z(n21794) );
  XNOR U30346 ( .A(n21795), .B(n21796), .Z(n21793) );
  XNOR U30347 ( .A(y[5311]), .B(x[5311]), .Z(n21796) );
  XNOR U30348 ( .A(y[5312]), .B(x[5312]), .Z(n21795) );
  XNOR U30349 ( .A(n21787), .B(n21788), .Z(n21798) );
  XNOR U30350 ( .A(y[5307]), .B(x[5307]), .Z(n21788) );
  XNOR U30351 ( .A(n21789), .B(n21790), .Z(n21787) );
  XNOR U30352 ( .A(y[5308]), .B(x[5308]), .Z(n21790) );
  XNOR U30353 ( .A(y[5309]), .B(x[5309]), .Z(n21789) );
  XOR U30354 ( .A(n21763), .B(n21764), .Z(n21782) );
  XNOR U30355 ( .A(n21779), .B(n21780), .Z(n21764) );
  XNOR U30356 ( .A(n21774), .B(n21775), .Z(n21780) );
  XNOR U30357 ( .A(n21776), .B(n21777), .Z(n21775) );
  XNOR U30358 ( .A(y[5305]), .B(x[5305]), .Z(n21777) );
  XNOR U30359 ( .A(y[5306]), .B(x[5306]), .Z(n21776) );
  XNOR U30360 ( .A(y[5304]), .B(x[5304]), .Z(n21774) );
  XNOR U30361 ( .A(n21768), .B(n21769), .Z(n21779) );
  XNOR U30362 ( .A(y[5301]), .B(x[5301]), .Z(n21769) );
  XNOR U30363 ( .A(n21770), .B(n21771), .Z(n21768) );
  XNOR U30364 ( .A(y[5302]), .B(x[5302]), .Z(n21771) );
  XNOR U30365 ( .A(y[5303]), .B(x[5303]), .Z(n21770) );
  XOR U30366 ( .A(n21762), .B(n21761), .Z(n21763) );
  XNOR U30367 ( .A(n21757), .B(n21758), .Z(n21761) );
  XNOR U30368 ( .A(y[5298]), .B(x[5298]), .Z(n21758) );
  XNOR U30369 ( .A(n21759), .B(n21760), .Z(n21757) );
  XNOR U30370 ( .A(y[5299]), .B(x[5299]), .Z(n21760) );
  XNOR U30371 ( .A(y[5300]), .B(x[5300]), .Z(n21759) );
  XNOR U30372 ( .A(n21751), .B(n21752), .Z(n21762) );
  XNOR U30373 ( .A(y[5295]), .B(x[5295]), .Z(n21752) );
  XNOR U30374 ( .A(n21753), .B(n21754), .Z(n21751) );
  XNOR U30375 ( .A(y[5296]), .B(x[5296]), .Z(n21754) );
  XNOR U30376 ( .A(y[5297]), .B(x[5297]), .Z(n21753) );
  NAND U30377 ( .A(n21818), .B(n21819), .Z(N63456) );
  NANDN U30378 ( .A(n21820), .B(n21821), .Z(n21819) );
  OR U30379 ( .A(n21822), .B(n21823), .Z(n21821) );
  NAND U30380 ( .A(n21822), .B(n21823), .Z(n21818) );
  XOR U30381 ( .A(n21822), .B(n21824), .Z(N63455) );
  XNOR U30382 ( .A(n21820), .B(n21823), .Z(n21824) );
  AND U30383 ( .A(n21825), .B(n21826), .Z(n21823) );
  NANDN U30384 ( .A(n21827), .B(n21828), .Z(n21826) );
  NANDN U30385 ( .A(n21829), .B(n21830), .Z(n21828) );
  NANDN U30386 ( .A(n21830), .B(n21829), .Z(n21825) );
  NAND U30387 ( .A(n21831), .B(n21832), .Z(n21820) );
  NANDN U30388 ( .A(n21833), .B(n21834), .Z(n21832) );
  OR U30389 ( .A(n21835), .B(n21836), .Z(n21834) );
  NAND U30390 ( .A(n21836), .B(n21835), .Z(n21831) );
  AND U30391 ( .A(n21837), .B(n21838), .Z(n21822) );
  NANDN U30392 ( .A(n21839), .B(n21840), .Z(n21838) );
  NANDN U30393 ( .A(n21841), .B(n21842), .Z(n21840) );
  NANDN U30394 ( .A(n21842), .B(n21841), .Z(n21837) );
  XOR U30395 ( .A(n21836), .B(n21843), .Z(N63454) );
  XOR U30396 ( .A(n21833), .B(n21835), .Z(n21843) );
  XNOR U30397 ( .A(n21829), .B(n21844), .Z(n21835) );
  XNOR U30398 ( .A(n21827), .B(n21830), .Z(n21844) );
  NAND U30399 ( .A(n21845), .B(n21846), .Z(n21830) );
  NAND U30400 ( .A(n21847), .B(n21848), .Z(n21846) );
  OR U30401 ( .A(n21849), .B(n21850), .Z(n21847) );
  NANDN U30402 ( .A(n21851), .B(n21849), .Z(n21845) );
  IV U30403 ( .A(n21850), .Z(n21851) );
  NAND U30404 ( .A(n21852), .B(n21853), .Z(n21827) );
  NAND U30405 ( .A(n21854), .B(n21855), .Z(n21853) );
  NANDN U30406 ( .A(n21856), .B(n21857), .Z(n21854) );
  NANDN U30407 ( .A(n21857), .B(n21856), .Z(n21852) );
  AND U30408 ( .A(n21858), .B(n21859), .Z(n21829) );
  NAND U30409 ( .A(n21860), .B(n21861), .Z(n21859) );
  OR U30410 ( .A(n21862), .B(n21863), .Z(n21860) );
  NANDN U30411 ( .A(n21864), .B(n21862), .Z(n21858) );
  NAND U30412 ( .A(n21865), .B(n21866), .Z(n21833) );
  NANDN U30413 ( .A(n21867), .B(n21868), .Z(n21866) );
  OR U30414 ( .A(n21869), .B(n21870), .Z(n21868) );
  NANDN U30415 ( .A(n21871), .B(n21869), .Z(n21865) );
  IV U30416 ( .A(n21870), .Z(n21871) );
  XNOR U30417 ( .A(n21841), .B(n21872), .Z(n21836) );
  XNOR U30418 ( .A(n21839), .B(n21842), .Z(n21872) );
  NAND U30419 ( .A(n21873), .B(n21874), .Z(n21842) );
  NAND U30420 ( .A(n21875), .B(n21876), .Z(n21874) );
  OR U30421 ( .A(n21877), .B(n21878), .Z(n21875) );
  NANDN U30422 ( .A(n21879), .B(n21877), .Z(n21873) );
  IV U30423 ( .A(n21878), .Z(n21879) );
  NAND U30424 ( .A(n21880), .B(n21881), .Z(n21839) );
  NAND U30425 ( .A(n21882), .B(n21883), .Z(n21881) );
  NANDN U30426 ( .A(n21884), .B(n21885), .Z(n21882) );
  NANDN U30427 ( .A(n21885), .B(n21884), .Z(n21880) );
  AND U30428 ( .A(n21886), .B(n21887), .Z(n21841) );
  NAND U30429 ( .A(n21888), .B(n21889), .Z(n21887) );
  OR U30430 ( .A(n21890), .B(n21891), .Z(n21888) );
  NANDN U30431 ( .A(n21892), .B(n21890), .Z(n21886) );
  XNOR U30432 ( .A(n21867), .B(n21893), .Z(N63453) );
  XOR U30433 ( .A(n21869), .B(n21870), .Z(n21893) );
  XNOR U30434 ( .A(n21883), .B(n21894), .Z(n21870) );
  XOR U30435 ( .A(n21884), .B(n21885), .Z(n21894) );
  XOR U30436 ( .A(n21890), .B(n21895), .Z(n21885) );
  XOR U30437 ( .A(n21889), .B(n21892), .Z(n21895) );
  IV U30438 ( .A(n21891), .Z(n21892) );
  NAND U30439 ( .A(n21896), .B(n21897), .Z(n21891) );
  OR U30440 ( .A(n21898), .B(n21899), .Z(n21897) );
  OR U30441 ( .A(n21900), .B(n21901), .Z(n21896) );
  NAND U30442 ( .A(n21902), .B(n21903), .Z(n21889) );
  OR U30443 ( .A(n21904), .B(n21905), .Z(n21903) );
  OR U30444 ( .A(n21906), .B(n21907), .Z(n21902) );
  NOR U30445 ( .A(n21908), .B(n21909), .Z(n21890) );
  ANDN U30446 ( .B(n21910), .A(n21911), .Z(n21884) );
  XNOR U30447 ( .A(n21877), .B(n21912), .Z(n21883) );
  XNOR U30448 ( .A(n21876), .B(n21878), .Z(n21912) );
  NAND U30449 ( .A(n21913), .B(n21914), .Z(n21878) );
  OR U30450 ( .A(n21915), .B(n21916), .Z(n21914) );
  OR U30451 ( .A(n21917), .B(n21918), .Z(n21913) );
  NAND U30452 ( .A(n21919), .B(n21920), .Z(n21876) );
  OR U30453 ( .A(n21921), .B(n21922), .Z(n21920) );
  OR U30454 ( .A(n21923), .B(n21924), .Z(n21919) );
  ANDN U30455 ( .B(n21925), .A(n21926), .Z(n21877) );
  IV U30456 ( .A(n21927), .Z(n21925) );
  ANDN U30457 ( .B(n21928), .A(n21929), .Z(n21869) );
  XOR U30458 ( .A(n21855), .B(n21930), .Z(n21867) );
  XOR U30459 ( .A(n21856), .B(n21857), .Z(n21930) );
  XOR U30460 ( .A(n21862), .B(n21931), .Z(n21857) );
  XOR U30461 ( .A(n21861), .B(n21864), .Z(n21931) );
  IV U30462 ( .A(n21863), .Z(n21864) );
  NAND U30463 ( .A(n21932), .B(n21933), .Z(n21863) );
  OR U30464 ( .A(n21934), .B(n21935), .Z(n21933) );
  OR U30465 ( .A(n21936), .B(n21937), .Z(n21932) );
  NAND U30466 ( .A(n21938), .B(n21939), .Z(n21861) );
  OR U30467 ( .A(n21940), .B(n21941), .Z(n21939) );
  OR U30468 ( .A(n21942), .B(n21943), .Z(n21938) );
  NOR U30469 ( .A(n21944), .B(n21945), .Z(n21862) );
  ANDN U30470 ( .B(n21946), .A(n21947), .Z(n21856) );
  IV U30471 ( .A(n21948), .Z(n21946) );
  XNOR U30472 ( .A(n21849), .B(n21949), .Z(n21855) );
  XNOR U30473 ( .A(n21848), .B(n21850), .Z(n21949) );
  NAND U30474 ( .A(n21950), .B(n21951), .Z(n21850) );
  OR U30475 ( .A(n21952), .B(n21953), .Z(n21951) );
  OR U30476 ( .A(n21954), .B(n21955), .Z(n21950) );
  NAND U30477 ( .A(n21956), .B(n21957), .Z(n21848) );
  OR U30478 ( .A(n21958), .B(n21959), .Z(n21957) );
  OR U30479 ( .A(n21960), .B(n21961), .Z(n21956) );
  ANDN U30480 ( .B(n21962), .A(n21963), .Z(n21849) );
  IV U30481 ( .A(n21964), .Z(n21962) );
  XNOR U30482 ( .A(n21929), .B(n21928), .Z(N63452) );
  XOR U30483 ( .A(n21948), .B(n21947), .Z(n21928) );
  XNOR U30484 ( .A(n21963), .B(n21964), .Z(n21947) );
  XNOR U30485 ( .A(n21958), .B(n21959), .Z(n21964) );
  XNOR U30486 ( .A(n21960), .B(n21961), .Z(n21959) );
  XNOR U30487 ( .A(y[5293]), .B(x[5293]), .Z(n21961) );
  XNOR U30488 ( .A(y[5294]), .B(x[5294]), .Z(n21960) );
  XNOR U30489 ( .A(y[5292]), .B(x[5292]), .Z(n21958) );
  XNOR U30490 ( .A(n21952), .B(n21953), .Z(n21963) );
  XNOR U30491 ( .A(y[5289]), .B(x[5289]), .Z(n21953) );
  XNOR U30492 ( .A(n21954), .B(n21955), .Z(n21952) );
  XNOR U30493 ( .A(y[5290]), .B(x[5290]), .Z(n21955) );
  XNOR U30494 ( .A(y[5291]), .B(x[5291]), .Z(n21954) );
  XNOR U30495 ( .A(n21945), .B(n21944), .Z(n21948) );
  XNOR U30496 ( .A(n21940), .B(n21941), .Z(n21944) );
  XNOR U30497 ( .A(y[5286]), .B(x[5286]), .Z(n21941) );
  XNOR U30498 ( .A(n21942), .B(n21943), .Z(n21940) );
  XNOR U30499 ( .A(y[5287]), .B(x[5287]), .Z(n21943) );
  XNOR U30500 ( .A(y[5288]), .B(x[5288]), .Z(n21942) );
  XNOR U30501 ( .A(n21934), .B(n21935), .Z(n21945) );
  XNOR U30502 ( .A(y[5283]), .B(x[5283]), .Z(n21935) );
  XNOR U30503 ( .A(n21936), .B(n21937), .Z(n21934) );
  XNOR U30504 ( .A(y[5284]), .B(x[5284]), .Z(n21937) );
  XNOR U30505 ( .A(y[5285]), .B(x[5285]), .Z(n21936) );
  XOR U30506 ( .A(n21910), .B(n21911), .Z(n21929) );
  XNOR U30507 ( .A(n21926), .B(n21927), .Z(n21911) );
  XNOR U30508 ( .A(n21921), .B(n21922), .Z(n21927) );
  XNOR U30509 ( .A(n21923), .B(n21924), .Z(n21922) );
  XNOR U30510 ( .A(y[5281]), .B(x[5281]), .Z(n21924) );
  XNOR U30511 ( .A(y[5282]), .B(x[5282]), .Z(n21923) );
  XNOR U30512 ( .A(y[5280]), .B(x[5280]), .Z(n21921) );
  XNOR U30513 ( .A(n21915), .B(n21916), .Z(n21926) );
  XNOR U30514 ( .A(y[5277]), .B(x[5277]), .Z(n21916) );
  XNOR U30515 ( .A(n21917), .B(n21918), .Z(n21915) );
  XNOR U30516 ( .A(y[5278]), .B(x[5278]), .Z(n21918) );
  XNOR U30517 ( .A(y[5279]), .B(x[5279]), .Z(n21917) );
  XOR U30518 ( .A(n21909), .B(n21908), .Z(n21910) );
  XNOR U30519 ( .A(n21904), .B(n21905), .Z(n21908) );
  XNOR U30520 ( .A(y[5274]), .B(x[5274]), .Z(n21905) );
  XNOR U30521 ( .A(n21906), .B(n21907), .Z(n21904) );
  XNOR U30522 ( .A(y[5275]), .B(x[5275]), .Z(n21907) );
  XNOR U30523 ( .A(y[5276]), .B(x[5276]), .Z(n21906) );
  XNOR U30524 ( .A(n21898), .B(n21899), .Z(n21909) );
  XNOR U30525 ( .A(y[5271]), .B(x[5271]), .Z(n21899) );
  XNOR U30526 ( .A(n21900), .B(n21901), .Z(n21898) );
  XNOR U30527 ( .A(y[5272]), .B(x[5272]), .Z(n21901) );
  XNOR U30528 ( .A(y[5273]), .B(x[5273]), .Z(n21900) );
  NAND U30529 ( .A(n21965), .B(n21966), .Z(N63443) );
  NANDN U30530 ( .A(n21967), .B(n21968), .Z(n21966) );
  OR U30531 ( .A(n21969), .B(n21970), .Z(n21968) );
  NAND U30532 ( .A(n21969), .B(n21970), .Z(n21965) );
  XOR U30533 ( .A(n21969), .B(n21971), .Z(N63442) );
  XNOR U30534 ( .A(n21967), .B(n21970), .Z(n21971) );
  AND U30535 ( .A(n21972), .B(n21973), .Z(n21970) );
  NANDN U30536 ( .A(n21974), .B(n21975), .Z(n21973) );
  NANDN U30537 ( .A(n21976), .B(n21977), .Z(n21975) );
  NANDN U30538 ( .A(n21977), .B(n21976), .Z(n21972) );
  NAND U30539 ( .A(n21978), .B(n21979), .Z(n21967) );
  NANDN U30540 ( .A(n21980), .B(n21981), .Z(n21979) );
  OR U30541 ( .A(n21982), .B(n21983), .Z(n21981) );
  NAND U30542 ( .A(n21983), .B(n21982), .Z(n21978) );
  AND U30543 ( .A(n21984), .B(n21985), .Z(n21969) );
  NANDN U30544 ( .A(n21986), .B(n21987), .Z(n21985) );
  NANDN U30545 ( .A(n21988), .B(n21989), .Z(n21987) );
  NANDN U30546 ( .A(n21989), .B(n21988), .Z(n21984) );
  XOR U30547 ( .A(n21983), .B(n21990), .Z(N63441) );
  XOR U30548 ( .A(n21980), .B(n21982), .Z(n21990) );
  XNOR U30549 ( .A(n21976), .B(n21991), .Z(n21982) );
  XNOR U30550 ( .A(n21974), .B(n21977), .Z(n21991) );
  NAND U30551 ( .A(n21992), .B(n21993), .Z(n21977) );
  NAND U30552 ( .A(n21994), .B(n21995), .Z(n21993) );
  OR U30553 ( .A(n21996), .B(n21997), .Z(n21994) );
  NANDN U30554 ( .A(n21998), .B(n21996), .Z(n21992) );
  IV U30555 ( .A(n21997), .Z(n21998) );
  NAND U30556 ( .A(n21999), .B(n22000), .Z(n21974) );
  NAND U30557 ( .A(n22001), .B(n22002), .Z(n22000) );
  NANDN U30558 ( .A(n22003), .B(n22004), .Z(n22001) );
  NANDN U30559 ( .A(n22004), .B(n22003), .Z(n21999) );
  AND U30560 ( .A(n22005), .B(n22006), .Z(n21976) );
  NAND U30561 ( .A(n22007), .B(n22008), .Z(n22006) );
  OR U30562 ( .A(n22009), .B(n22010), .Z(n22007) );
  NANDN U30563 ( .A(n22011), .B(n22009), .Z(n22005) );
  NAND U30564 ( .A(n22012), .B(n22013), .Z(n21980) );
  NANDN U30565 ( .A(n22014), .B(n22015), .Z(n22013) );
  OR U30566 ( .A(n22016), .B(n22017), .Z(n22015) );
  NANDN U30567 ( .A(n22018), .B(n22016), .Z(n22012) );
  IV U30568 ( .A(n22017), .Z(n22018) );
  XNOR U30569 ( .A(n21988), .B(n22019), .Z(n21983) );
  XNOR U30570 ( .A(n21986), .B(n21989), .Z(n22019) );
  NAND U30571 ( .A(n22020), .B(n22021), .Z(n21989) );
  NAND U30572 ( .A(n22022), .B(n22023), .Z(n22021) );
  OR U30573 ( .A(n22024), .B(n22025), .Z(n22022) );
  NANDN U30574 ( .A(n22026), .B(n22024), .Z(n22020) );
  IV U30575 ( .A(n22025), .Z(n22026) );
  NAND U30576 ( .A(n22027), .B(n22028), .Z(n21986) );
  NAND U30577 ( .A(n22029), .B(n22030), .Z(n22028) );
  NANDN U30578 ( .A(n22031), .B(n22032), .Z(n22029) );
  NANDN U30579 ( .A(n22032), .B(n22031), .Z(n22027) );
  AND U30580 ( .A(n22033), .B(n22034), .Z(n21988) );
  NAND U30581 ( .A(n22035), .B(n22036), .Z(n22034) );
  OR U30582 ( .A(n22037), .B(n22038), .Z(n22035) );
  NANDN U30583 ( .A(n22039), .B(n22037), .Z(n22033) );
  XNOR U30584 ( .A(n22014), .B(n22040), .Z(N63440) );
  XOR U30585 ( .A(n22016), .B(n22017), .Z(n22040) );
  XNOR U30586 ( .A(n22030), .B(n22041), .Z(n22017) );
  XOR U30587 ( .A(n22031), .B(n22032), .Z(n22041) );
  XOR U30588 ( .A(n22037), .B(n22042), .Z(n22032) );
  XOR U30589 ( .A(n22036), .B(n22039), .Z(n22042) );
  IV U30590 ( .A(n22038), .Z(n22039) );
  NAND U30591 ( .A(n22043), .B(n22044), .Z(n22038) );
  OR U30592 ( .A(n22045), .B(n22046), .Z(n22044) );
  OR U30593 ( .A(n22047), .B(n22048), .Z(n22043) );
  NAND U30594 ( .A(n22049), .B(n22050), .Z(n22036) );
  OR U30595 ( .A(n22051), .B(n22052), .Z(n22050) );
  OR U30596 ( .A(n22053), .B(n22054), .Z(n22049) );
  NOR U30597 ( .A(n22055), .B(n22056), .Z(n22037) );
  ANDN U30598 ( .B(n22057), .A(n22058), .Z(n22031) );
  XNOR U30599 ( .A(n22024), .B(n22059), .Z(n22030) );
  XNOR U30600 ( .A(n22023), .B(n22025), .Z(n22059) );
  NAND U30601 ( .A(n22060), .B(n22061), .Z(n22025) );
  OR U30602 ( .A(n22062), .B(n22063), .Z(n22061) );
  OR U30603 ( .A(n22064), .B(n22065), .Z(n22060) );
  NAND U30604 ( .A(n22066), .B(n22067), .Z(n22023) );
  OR U30605 ( .A(n22068), .B(n22069), .Z(n22067) );
  OR U30606 ( .A(n22070), .B(n22071), .Z(n22066) );
  ANDN U30607 ( .B(n22072), .A(n22073), .Z(n22024) );
  IV U30608 ( .A(n22074), .Z(n22072) );
  ANDN U30609 ( .B(n22075), .A(n22076), .Z(n22016) );
  XOR U30610 ( .A(n22002), .B(n22077), .Z(n22014) );
  XOR U30611 ( .A(n22003), .B(n22004), .Z(n22077) );
  XOR U30612 ( .A(n22009), .B(n22078), .Z(n22004) );
  XOR U30613 ( .A(n22008), .B(n22011), .Z(n22078) );
  IV U30614 ( .A(n22010), .Z(n22011) );
  NAND U30615 ( .A(n22079), .B(n22080), .Z(n22010) );
  OR U30616 ( .A(n22081), .B(n22082), .Z(n22080) );
  OR U30617 ( .A(n22083), .B(n22084), .Z(n22079) );
  NAND U30618 ( .A(n22085), .B(n22086), .Z(n22008) );
  OR U30619 ( .A(n22087), .B(n22088), .Z(n22086) );
  OR U30620 ( .A(n22089), .B(n22090), .Z(n22085) );
  NOR U30621 ( .A(n22091), .B(n22092), .Z(n22009) );
  ANDN U30622 ( .B(n22093), .A(n22094), .Z(n22003) );
  IV U30623 ( .A(n22095), .Z(n22093) );
  XNOR U30624 ( .A(n21996), .B(n22096), .Z(n22002) );
  XNOR U30625 ( .A(n21995), .B(n21997), .Z(n22096) );
  NAND U30626 ( .A(n22097), .B(n22098), .Z(n21997) );
  OR U30627 ( .A(n22099), .B(n22100), .Z(n22098) );
  OR U30628 ( .A(n22101), .B(n22102), .Z(n22097) );
  NAND U30629 ( .A(n22103), .B(n22104), .Z(n21995) );
  OR U30630 ( .A(n22105), .B(n22106), .Z(n22104) );
  OR U30631 ( .A(n22107), .B(n22108), .Z(n22103) );
  ANDN U30632 ( .B(n22109), .A(n22110), .Z(n21996) );
  IV U30633 ( .A(n22111), .Z(n22109) );
  XNOR U30634 ( .A(n22076), .B(n22075), .Z(N63439) );
  XOR U30635 ( .A(n22095), .B(n22094), .Z(n22075) );
  XNOR U30636 ( .A(n22110), .B(n22111), .Z(n22094) );
  XNOR U30637 ( .A(n22105), .B(n22106), .Z(n22111) );
  XNOR U30638 ( .A(n22107), .B(n22108), .Z(n22106) );
  XNOR U30639 ( .A(y[5269]), .B(x[5269]), .Z(n22108) );
  XNOR U30640 ( .A(y[5270]), .B(x[5270]), .Z(n22107) );
  XNOR U30641 ( .A(y[5268]), .B(x[5268]), .Z(n22105) );
  XNOR U30642 ( .A(n22099), .B(n22100), .Z(n22110) );
  XNOR U30643 ( .A(y[5265]), .B(x[5265]), .Z(n22100) );
  XNOR U30644 ( .A(n22101), .B(n22102), .Z(n22099) );
  XNOR U30645 ( .A(y[5266]), .B(x[5266]), .Z(n22102) );
  XNOR U30646 ( .A(y[5267]), .B(x[5267]), .Z(n22101) );
  XNOR U30647 ( .A(n22092), .B(n22091), .Z(n22095) );
  XNOR U30648 ( .A(n22087), .B(n22088), .Z(n22091) );
  XNOR U30649 ( .A(y[5262]), .B(x[5262]), .Z(n22088) );
  XNOR U30650 ( .A(n22089), .B(n22090), .Z(n22087) );
  XNOR U30651 ( .A(y[5263]), .B(x[5263]), .Z(n22090) );
  XNOR U30652 ( .A(y[5264]), .B(x[5264]), .Z(n22089) );
  XNOR U30653 ( .A(n22081), .B(n22082), .Z(n22092) );
  XNOR U30654 ( .A(y[5259]), .B(x[5259]), .Z(n22082) );
  XNOR U30655 ( .A(n22083), .B(n22084), .Z(n22081) );
  XNOR U30656 ( .A(y[5260]), .B(x[5260]), .Z(n22084) );
  XNOR U30657 ( .A(y[5261]), .B(x[5261]), .Z(n22083) );
  XOR U30658 ( .A(n22057), .B(n22058), .Z(n22076) );
  XNOR U30659 ( .A(n22073), .B(n22074), .Z(n22058) );
  XNOR U30660 ( .A(n22068), .B(n22069), .Z(n22074) );
  XNOR U30661 ( .A(n22070), .B(n22071), .Z(n22069) );
  XNOR U30662 ( .A(y[5257]), .B(x[5257]), .Z(n22071) );
  XNOR U30663 ( .A(y[5258]), .B(x[5258]), .Z(n22070) );
  XNOR U30664 ( .A(y[5256]), .B(x[5256]), .Z(n22068) );
  XNOR U30665 ( .A(n22062), .B(n22063), .Z(n22073) );
  XNOR U30666 ( .A(y[5253]), .B(x[5253]), .Z(n22063) );
  XNOR U30667 ( .A(n22064), .B(n22065), .Z(n22062) );
  XNOR U30668 ( .A(y[5254]), .B(x[5254]), .Z(n22065) );
  XNOR U30669 ( .A(y[5255]), .B(x[5255]), .Z(n22064) );
  XOR U30670 ( .A(n22056), .B(n22055), .Z(n22057) );
  XNOR U30671 ( .A(n22051), .B(n22052), .Z(n22055) );
  XNOR U30672 ( .A(y[5250]), .B(x[5250]), .Z(n22052) );
  XNOR U30673 ( .A(n22053), .B(n22054), .Z(n22051) );
  XNOR U30674 ( .A(y[5251]), .B(x[5251]), .Z(n22054) );
  XNOR U30675 ( .A(y[5252]), .B(x[5252]), .Z(n22053) );
  XNOR U30676 ( .A(n22045), .B(n22046), .Z(n22056) );
  XNOR U30677 ( .A(y[5247]), .B(x[5247]), .Z(n22046) );
  XNOR U30678 ( .A(n22047), .B(n22048), .Z(n22045) );
  XNOR U30679 ( .A(y[5248]), .B(x[5248]), .Z(n22048) );
  XNOR U30680 ( .A(y[5249]), .B(x[5249]), .Z(n22047) );
  NAND U30681 ( .A(n22112), .B(n22113), .Z(N63430) );
  NANDN U30682 ( .A(n22114), .B(n22115), .Z(n22113) );
  OR U30683 ( .A(n22116), .B(n22117), .Z(n22115) );
  NAND U30684 ( .A(n22116), .B(n22117), .Z(n22112) );
  XOR U30685 ( .A(n22116), .B(n22118), .Z(N63429) );
  XNOR U30686 ( .A(n22114), .B(n22117), .Z(n22118) );
  AND U30687 ( .A(n22119), .B(n22120), .Z(n22117) );
  NANDN U30688 ( .A(n22121), .B(n22122), .Z(n22120) );
  NANDN U30689 ( .A(n22123), .B(n22124), .Z(n22122) );
  NANDN U30690 ( .A(n22124), .B(n22123), .Z(n22119) );
  NAND U30691 ( .A(n22125), .B(n22126), .Z(n22114) );
  NANDN U30692 ( .A(n22127), .B(n22128), .Z(n22126) );
  OR U30693 ( .A(n22129), .B(n22130), .Z(n22128) );
  NAND U30694 ( .A(n22130), .B(n22129), .Z(n22125) );
  AND U30695 ( .A(n22131), .B(n22132), .Z(n22116) );
  NANDN U30696 ( .A(n22133), .B(n22134), .Z(n22132) );
  NANDN U30697 ( .A(n22135), .B(n22136), .Z(n22134) );
  NANDN U30698 ( .A(n22136), .B(n22135), .Z(n22131) );
  XOR U30699 ( .A(n22130), .B(n22137), .Z(N63428) );
  XOR U30700 ( .A(n22127), .B(n22129), .Z(n22137) );
  XNOR U30701 ( .A(n22123), .B(n22138), .Z(n22129) );
  XNOR U30702 ( .A(n22121), .B(n22124), .Z(n22138) );
  NAND U30703 ( .A(n22139), .B(n22140), .Z(n22124) );
  NAND U30704 ( .A(n22141), .B(n22142), .Z(n22140) );
  OR U30705 ( .A(n22143), .B(n22144), .Z(n22141) );
  NANDN U30706 ( .A(n22145), .B(n22143), .Z(n22139) );
  IV U30707 ( .A(n22144), .Z(n22145) );
  NAND U30708 ( .A(n22146), .B(n22147), .Z(n22121) );
  NAND U30709 ( .A(n22148), .B(n22149), .Z(n22147) );
  NANDN U30710 ( .A(n22150), .B(n22151), .Z(n22148) );
  NANDN U30711 ( .A(n22151), .B(n22150), .Z(n22146) );
  AND U30712 ( .A(n22152), .B(n22153), .Z(n22123) );
  NAND U30713 ( .A(n22154), .B(n22155), .Z(n22153) );
  OR U30714 ( .A(n22156), .B(n22157), .Z(n22154) );
  NANDN U30715 ( .A(n22158), .B(n22156), .Z(n22152) );
  NAND U30716 ( .A(n22159), .B(n22160), .Z(n22127) );
  NANDN U30717 ( .A(n22161), .B(n22162), .Z(n22160) );
  OR U30718 ( .A(n22163), .B(n22164), .Z(n22162) );
  NANDN U30719 ( .A(n22165), .B(n22163), .Z(n22159) );
  IV U30720 ( .A(n22164), .Z(n22165) );
  XNOR U30721 ( .A(n22135), .B(n22166), .Z(n22130) );
  XNOR U30722 ( .A(n22133), .B(n22136), .Z(n22166) );
  NAND U30723 ( .A(n22167), .B(n22168), .Z(n22136) );
  NAND U30724 ( .A(n22169), .B(n22170), .Z(n22168) );
  OR U30725 ( .A(n22171), .B(n22172), .Z(n22169) );
  NANDN U30726 ( .A(n22173), .B(n22171), .Z(n22167) );
  IV U30727 ( .A(n22172), .Z(n22173) );
  NAND U30728 ( .A(n22174), .B(n22175), .Z(n22133) );
  NAND U30729 ( .A(n22176), .B(n22177), .Z(n22175) );
  NANDN U30730 ( .A(n22178), .B(n22179), .Z(n22176) );
  NANDN U30731 ( .A(n22179), .B(n22178), .Z(n22174) );
  AND U30732 ( .A(n22180), .B(n22181), .Z(n22135) );
  NAND U30733 ( .A(n22182), .B(n22183), .Z(n22181) );
  OR U30734 ( .A(n22184), .B(n22185), .Z(n22182) );
  NANDN U30735 ( .A(n22186), .B(n22184), .Z(n22180) );
  XNOR U30736 ( .A(n22161), .B(n22187), .Z(N63427) );
  XOR U30737 ( .A(n22163), .B(n22164), .Z(n22187) );
  XNOR U30738 ( .A(n22177), .B(n22188), .Z(n22164) );
  XOR U30739 ( .A(n22178), .B(n22179), .Z(n22188) );
  XOR U30740 ( .A(n22184), .B(n22189), .Z(n22179) );
  XOR U30741 ( .A(n22183), .B(n22186), .Z(n22189) );
  IV U30742 ( .A(n22185), .Z(n22186) );
  NAND U30743 ( .A(n22190), .B(n22191), .Z(n22185) );
  OR U30744 ( .A(n22192), .B(n22193), .Z(n22191) );
  OR U30745 ( .A(n22194), .B(n22195), .Z(n22190) );
  NAND U30746 ( .A(n22196), .B(n22197), .Z(n22183) );
  OR U30747 ( .A(n22198), .B(n22199), .Z(n22197) );
  OR U30748 ( .A(n22200), .B(n22201), .Z(n22196) );
  NOR U30749 ( .A(n22202), .B(n22203), .Z(n22184) );
  ANDN U30750 ( .B(n22204), .A(n22205), .Z(n22178) );
  XNOR U30751 ( .A(n22171), .B(n22206), .Z(n22177) );
  XNOR U30752 ( .A(n22170), .B(n22172), .Z(n22206) );
  NAND U30753 ( .A(n22207), .B(n22208), .Z(n22172) );
  OR U30754 ( .A(n22209), .B(n22210), .Z(n22208) );
  OR U30755 ( .A(n22211), .B(n22212), .Z(n22207) );
  NAND U30756 ( .A(n22213), .B(n22214), .Z(n22170) );
  OR U30757 ( .A(n22215), .B(n22216), .Z(n22214) );
  OR U30758 ( .A(n22217), .B(n22218), .Z(n22213) );
  ANDN U30759 ( .B(n22219), .A(n22220), .Z(n22171) );
  IV U30760 ( .A(n22221), .Z(n22219) );
  ANDN U30761 ( .B(n22222), .A(n22223), .Z(n22163) );
  XOR U30762 ( .A(n22149), .B(n22224), .Z(n22161) );
  XOR U30763 ( .A(n22150), .B(n22151), .Z(n22224) );
  XOR U30764 ( .A(n22156), .B(n22225), .Z(n22151) );
  XOR U30765 ( .A(n22155), .B(n22158), .Z(n22225) );
  IV U30766 ( .A(n22157), .Z(n22158) );
  NAND U30767 ( .A(n22226), .B(n22227), .Z(n22157) );
  OR U30768 ( .A(n22228), .B(n22229), .Z(n22227) );
  OR U30769 ( .A(n22230), .B(n22231), .Z(n22226) );
  NAND U30770 ( .A(n22232), .B(n22233), .Z(n22155) );
  OR U30771 ( .A(n22234), .B(n22235), .Z(n22233) );
  OR U30772 ( .A(n22236), .B(n22237), .Z(n22232) );
  NOR U30773 ( .A(n22238), .B(n22239), .Z(n22156) );
  ANDN U30774 ( .B(n22240), .A(n22241), .Z(n22150) );
  IV U30775 ( .A(n22242), .Z(n22240) );
  XNOR U30776 ( .A(n22143), .B(n22243), .Z(n22149) );
  XNOR U30777 ( .A(n22142), .B(n22144), .Z(n22243) );
  NAND U30778 ( .A(n22244), .B(n22245), .Z(n22144) );
  OR U30779 ( .A(n22246), .B(n22247), .Z(n22245) );
  OR U30780 ( .A(n22248), .B(n22249), .Z(n22244) );
  NAND U30781 ( .A(n22250), .B(n22251), .Z(n22142) );
  OR U30782 ( .A(n22252), .B(n22253), .Z(n22251) );
  OR U30783 ( .A(n22254), .B(n22255), .Z(n22250) );
  ANDN U30784 ( .B(n22256), .A(n22257), .Z(n22143) );
  IV U30785 ( .A(n22258), .Z(n22256) );
  XNOR U30786 ( .A(n22223), .B(n22222), .Z(N63426) );
  XOR U30787 ( .A(n22242), .B(n22241), .Z(n22222) );
  XNOR U30788 ( .A(n22257), .B(n22258), .Z(n22241) );
  XNOR U30789 ( .A(n22252), .B(n22253), .Z(n22258) );
  XNOR U30790 ( .A(n22254), .B(n22255), .Z(n22253) );
  XNOR U30791 ( .A(y[5245]), .B(x[5245]), .Z(n22255) );
  XNOR U30792 ( .A(y[5246]), .B(x[5246]), .Z(n22254) );
  XNOR U30793 ( .A(y[5244]), .B(x[5244]), .Z(n22252) );
  XNOR U30794 ( .A(n22246), .B(n22247), .Z(n22257) );
  XNOR U30795 ( .A(y[5241]), .B(x[5241]), .Z(n22247) );
  XNOR U30796 ( .A(n22248), .B(n22249), .Z(n22246) );
  XNOR U30797 ( .A(y[5242]), .B(x[5242]), .Z(n22249) );
  XNOR U30798 ( .A(y[5243]), .B(x[5243]), .Z(n22248) );
  XNOR U30799 ( .A(n22239), .B(n22238), .Z(n22242) );
  XNOR U30800 ( .A(n22234), .B(n22235), .Z(n22238) );
  XNOR U30801 ( .A(y[5238]), .B(x[5238]), .Z(n22235) );
  XNOR U30802 ( .A(n22236), .B(n22237), .Z(n22234) );
  XNOR U30803 ( .A(y[5239]), .B(x[5239]), .Z(n22237) );
  XNOR U30804 ( .A(y[5240]), .B(x[5240]), .Z(n22236) );
  XNOR U30805 ( .A(n22228), .B(n22229), .Z(n22239) );
  XNOR U30806 ( .A(y[5235]), .B(x[5235]), .Z(n22229) );
  XNOR U30807 ( .A(n22230), .B(n22231), .Z(n22228) );
  XNOR U30808 ( .A(y[5236]), .B(x[5236]), .Z(n22231) );
  XNOR U30809 ( .A(y[5237]), .B(x[5237]), .Z(n22230) );
  XOR U30810 ( .A(n22204), .B(n22205), .Z(n22223) );
  XNOR U30811 ( .A(n22220), .B(n22221), .Z(n22205) );
  XNOR U30812 ( .A(n22215), .B(n22216), .Z(n22221) );
  XNOR U30813 ( .A(n22217), .B(n22218), .Z(n22216) );
  XNOR U30814 ( .A(y[5233]), .B(x[5233]), .Z(n22218) );
  XNOR U30815 ( .A(y[5234]), .B(x[5234]), .Z(n22217) );
  XNOR U30816 ( .A(y[5232]), .B(x[5232]), .Z(n22215) );
  XNOR U30817 ( .A(n22209), .B(n22210), .Z(n22220) );
  XNOR U30818 ( .A(y[5229]), .B(x[5229]), .Z(n22210) );
  XNOR U30819 ( .A(n22211), .B(n22212), .Z(n22209) );
  XNOR U30820 ( .A(y[5230]), .B(x[5230]), .Z(n22212) );
  XNOR U30821 ( .A(y[5231]), .B(x[5231]), .Z(n22211) );
  XOR U30822 ( .A(n22203), .B(n22202), .Z(n22204) );
  XNOR U30823 ( .A(n22198), .B(n22199), .Z(n22202) );
  XNOR U30824 ( .A(y[5226]), .B(x[5226]), .Z(n22199) );
  XNOR U30825 ( .A(n22200), .B(n22201), .Z(n22198) );
  XNOR U30826 ( .A(y[5227]), .B(x[5227]), .Z(n22201) );
  XNOR U30827 ( .A(y[5228]), .B(x[5228]), .Z(n22200) );
  XNOR U30828 ( .A(n22192), .B(n22193), .Z(n22203) );
  XNOR U30829 ( .A(y[5223]), .B(x[5223]), .Z(n22193) );
  XNOR U30830 ( .A(n22194), .B(n22195), .Z(n22192) );
  XNOR U30831 ( .A(y[5224]), .B(x[5224]), .Z(n22195) );
  XNOR U30832 ( .A(y[5225]), .B(x[5225]), .Z(n22194) );
  NAND U30833 ( .A(n22259), .B(n22260), .Z(N63417) );
  NANDN U30834 ( .A(n22261), .B(n22262), .Z(n22260) );
  OR U30835 ( .A(n22263), .B(n22264), .Z(n22262) );
  NAND U30836 ( .A(n22263), .B(n22264), .Z(n22259) );
  XOR U30837 ( .A(n22263), .B(n22265), .Z(N63416) );
  XNOR U30838 ( .A(n22261), .B(n22264), .Z(n22265) );
  AND U30839 ( .A(n22266), .B(n22267), .Z(n22264) );
  NANDN U30840 ( .A(n22268), .B(n22269), .Z(n22267) );
  NANDN U30841 ( .A(n22270), .B(n22271), .Z(n22269) );
  NANDN U30842 ( .A(n22271), .B(n22270), .Z(n22266) );
  NAND U30843 ( .A(n22272), .B(n22273), .Z(n22261) );
  NANDN U30844 ( .A(n22274), .B(n22275), .Z(n22273) );
  OR U30845 ( .A(n22276), .B(n22277), .Z(n22275) );
  NAND U30846 ( .A(n22277), .B(n22276), .Z(n22272) );
  AND U30847 ( .A(n22278), .B(n22279), .Z(n22263) );
  NANDN U30848 ( .A(n22280), .B(n22281), .Z(n22279) );
  NANDN U30849 ( .A(n22282), .B(n22283), .Z(n22281) );
  NANDN U30850 ( .A(n22283), .B(n22282), .Z(n22278) );
  XOR U30851 ( .A(n22277), .B(n22284), .Z(N63415) );
  XOR U30852 ( .A(n22274), .B(n22276), .Z(n22284) );
  XNOR U30853 ( .A(n22270), .B(n22285), .Z(n22276) );
  XNOR U30854 ( .A(n22268), .B(n22271), .Z(n22285) );
  NAND U30855 ( .A(n22286), .B(n22287), .Z(n22271) );
  NAND U30856 ( .A(n22288), .B(n22289), .Z(n22287) );
  OR U30857 ( .A(n22290), .B(n22291), .Z(n22288) );
  NANDN U30858 ( .A(n22292), .B(n22290), .Z(n22286) );
  IV U30859 ( .A(n22291), .Z(n22292) );
  NAND U30860 ( .A(n22293), .B(n22294), .Z(n22268) );
  NAND U30861 ( .A(n22295), .B(n22296), .Z(n22294) );
  NANDN U30862 ( .A(n22297), .B(n22298), .Z(n22295) );
  NANDN U30863 ( .A(n22298), .B(n22297), .Z(n22293) );
  AND U30864 ( .A(n22299), .B(n22300), .Z(n22270) );
  NAND U30865 ( .A(n22301), .B(n22302), .Z(n22300) );
  OR U30866 ( .A(n22303), .B(n22304), .Z(n22301) );
  NANDN U30867 ( .A(n22305), .B(n22303), .Z(n22299) );
  NAND U30868 ( .A(n22306), .B(n22307), .Z(n22274) );
  NANDN U30869 ( .A(n22308), .B(n22309), .Z(n22307) );
  OR U30870 ( .A(n22310), .B(n22311), .Z(n22309) );
  NANDN U30871 ( .A(n22312), .B(n22310), .Z(n22306) );
  IV U30872 ( .A(n22311), .Z(n22312) );
  XNOR U30873 ( .A(n22282), .B(n22313), .Z(n22277) );
  XNOR U30874 ( .A(n22280), .B(n22283), .Z(n22313) );
  NAND U30875 ( .A(n22314), .B(n22315), .Z(n22283) );
  NAND U30876 ( .A(n22316), .B(n22317), .Z(n22315) );
  OR U30877 ( .A(n22318), .B(n22319), .Z(n22316) );
  NANDN U30878 ( .A(n22320), .B(n22318), .Z(n22314) );
  IV U30879 ( .A(n22319), .Z(n22320) );
  NAND U30880 ( .A(n22321), .B(n22322), .Z(n22280) );
  NAND U30881 ( .A(n22323), .B(n22324), .Z(n22322) );
  NANDN U30882 ( .A(n22325), .B(n22326), .Z(n22323) );
  NANDN U30883 ( .A(n22326), .B(n22325), .Z(n22321) );
  AND U30884 ( .A(n22327), .B(n22328), .Z(n22282) );
  NAND U30885 ( .A(n22329), .B(n22330), .Z(n22328) );
  OR U30886 ( .A(n22331), .B(n22332), .Z(n22329) );
  NANDN U30887 ( .A(n22333), .B(n22331), .Z(n22327) );
  XNOR U30888 ( .A(n22308), .B(n22334), .Z(N63414) );
  XOR U30889 ( .A(n22310), .B(n22311), .Z(n22334) );
  XNOR U30890 ( .A(n22324), .B(n22335), .Z(n22311) );
  XOR U30891 ( .A(n22325), .B(n22326), .Z(n22335) );
  XOR U30892 ( .A(n22331), .B(n22336), .Z(n22326) );
  XOR U30893 ( .A(n22330), .B(n22333), .Z(n22336) );
  IV U30894 ( .A(n22332), .Z(n22333) );
  NAND U30895 ( .A(n22337), .B(n22338), .Z(n22332) );
  OR U30896 ( .A(n22339), .B(n22340), .Z(n22338) );
  OR U30897 ( .A(n22341), .B(n22342), .Z(n22337) );
  NAND U30898 ( .A(n22343), .B(n22344), .Z(n22330) );
  OR U30899 ( .A(n22345), .B(n22346), .Z(n22344) );
  OR U30900 ( .A(n22347), .B(n22348), .Z(n22343) );
  NOR U30901 ( .A(n22349), .B(n22350), .Z(n22331) );
  ANDN U30902 ( .B(n22351), .A(n22352), .Z(n22325) );
  XNOR U30903 ( .A(n22318), .B(n22353), .Z(n22324) );
  XNOR U30904 ( .A(n22317), .B(n22319), .Z(n22353) );
  NAND U30905 ( .A(n22354), .B(n22355), .Z(n22319) );
  OR U30906 ( .A(n22356), .B(n22357), .Z(n22355) );
  OR U30907 ( .A(n22358), .B(n22359), .Z(n22354) );
  NAND U30908 ( .A(n22360), .B(n22361), .Z(n22317) );
  OR U30909 ( .A(n22362), .B(n22363), .Z(n22361) );
  OR U30910 ( .A(n22364), .B(n22365), .Z(n22360) );
  ANDN U30911 ( .B(n22366), .A(n22367), .Z(n22318) );
  IV U30912 ( .A(n22368), .Z(n22366) );
  ANDN U30913 ( .B(n22369), .A(n22370), .Z(n22310) );
  XOR U30914 ( .A(n22296), .B(n22371), .Z(n22308) );
  XOR U30915 ( .A(n22297), .B(n22298), .Z(n22371) );
  XOR U30916 ( .A(n22303), .B(n22372), .Z(n22298) );
  XOR U30917 ( .A(n22302), .B(n22305), .Z(n22372) );
  IV U30918 ( .A(n22304), .Z(n22305) );
  NAND U30919 ( .A(n22373), .B(n22374), .Z(n22304) );
  OR U30920 ( .A(n22375), .B(n22376), .Z(n22374) );
  OR U30921 ( .A(n22377), .B(n22378), .Z(n22373) );
  NAND U30922 ( .A(n22379), .B(n22380), .Z(n22302) );
  OR U30923 ( .A(n22381), .B(n22382), .Z(n22380) );
  OR U30924 ( .A(n22383), .B(n22384), .Z(n22379) );
  NOR U30925 ( .A(n22385), .B(n22386), .Z(n22303) );
  ANDN U30926 ( .B(n22387), .A(n22388), .Z(n22297) );
  IV U30927 ( .A(n22389), .Z(n22387) );
  XNOR U30928 ( .A(n22290), .B(n22390), .Z(n22296) );
  XNOR U30929 ( .A(n22289), .B(n22291), .Z(n22390) );
  NAND U30930 ( .A(n22391), .B(n22392), .Z(n22291) );
  OR U30931 ( .A(n22393), .B(n22394), .Z(n22392) );
  OR U30932 ( .A(n22395), .B(n22396), .Z(n22391) );
  NAND U30933 ( .A(n22397), .B(n22398), .Z(n22289) );
  OR U30934 ( .A(n22399), .B(n22400), .Z(n22398) );
  OR U30935 ( .A(n22401), .B(n22402), .Z(n22397) );
  ANDN U30936 ( .B(n22403), .A(n22404), .Z(n22290) );
  IV U30937 ( .A(n22405), .Z(n22403) );
  XNOR U30938 ( .A(n22370), .B(n22369), .Z(N63413) );
  XOR U30939 ( .A(n22389), .B(n22388), .Z(n22369) );
  XNOR U30940 ( .A(n22404), .B(n22405), .Z(n22388) );
  XNOR U30941 ( .A(n22399), .B(n22400), .Z(n22405) );
  XNOR U30942 ( .A(n22401), .B(n22402), .Z(n22400) );
  XNOR U30943 ( .A(y[5221]), .B(x[5221]), .Z(n22402) );
  XNOR U30944 ( .A(y[5222]), .B(x[5222]), .Z(n22401) );
  XNOR U30945 ( .A(y[5220]), .B(x[5220]), .Z(n22399) );
  XNOR U30946 ( .A(n22393), .B(n22394), .Z(n22404) );
  XNOR U30947 ( .A(y[5217]), .B(x[5217]), .Z(n22394) );
  XNOR U30948 ( .A(n22395), .B(n22396), .Z(n22393) );
  XNOR U30949 ( .A(y[5218]), .B(x[5218]), .Z(n22396) );
  XNOR U30950 ( .A(y[5219]), .B(x[5219]), .Z(n22395) );
  XNOR U30951 ( .A(n22386), .B(n22385), .Z(n22389) );
  XNOR U30952 ( .A(n22381), .B(n22382), .Z(n22385) );
  XNOR U30953 ( .A(y[5214]), .B(x[5214]), .Z(n22382) );
  XNOR U30954 ( .A(n22383), .B(n22384), .Z(n22381) );
  XNOR U30955 ( .A(y[5215]), .B(x[5215]), .Z(n22384) );
  XNOR U30956 ( .A(y[5216]), .B(x[5216]), .Z(n22383) );
  XNOR U30957 ( .A(n22375), .B(n22376), .Z(n22386) );
  XNOR U30958 ( .A(y[5211]), .B(x[5211]), .Z(n22376) );
  XNOR U30959 ( .A(n22377), .B(n22378), .Z(n22375) );
  XNOR U30960 ( .A(y[5212]), .B(x[5212]), .Z(n22378) );
  XNOR U30961 ( .A(y[5213]), .B(x[5213]), .Z(n22377) );
  XOR U30962 ( .A(n22351), .B(n22352), .Z(n22370) );
  XNOR U30963 ( .A(n22367), .B(n22368), .Z(n22352) );
  XNOR U30964 ( .A(n22362), .B(n22363), .Z(n22368) );
  XNOR U30965 ( .A(n22364), .B(n22365), .Z(n22363) );
  XNOR U30966 ( .A(y[5209]), .B(x[5209]), .Z(n22365) );
  XNOR U30967 ( .A(y[5210]), .B(x[5210]), .Z(n22364) );
  XNOR U30968 ( .A(y[5208]), .B(x[5208]), .Z(n22362) );
  XNOR U30969 ( .A(n22356), .B(n22357), .Z(n22367) );
  XNOR U30970 ( .A(y[5205]), .B(x[5205]), .Z(n22357) );
  XNOR U30971 ( .A(n22358), .B(n22359), .Z(n22356) );
  XNOR U30972 ( .A(y[5206]), .B(x[5206]), .Z(n22359) );
  XNOR U30973 ( .A(y[5207]), .B(x[5207]), .Z(n22358) );
  XOR U30974 ( .A(n22350), .B(n22349), .Z(n22351) );
  XNOR U30975 ( .A(n22345), .B(n22346), .Z(n22349) );
  XNOR U30976 ( .A(y[5202]), .B(x[5202]), .Z(n22346) );
  XNOR U30977 ( .A(n22347), .B(n22348), .Z(n22345) );
  XNOR U30978 ( .A(y[5203]), .B(x[5203]), .Z(n22348) );
  XNOR U30979 ( .A(y[5204]), .B(x[5204]), .Z(n22347) );
  XNOR U30980 ( .A(n22339), .B(n22340), .Z(n22350) );
  XNOR U30981 ( .A(y[5199]), .B(x[5199]), .Z(n22340) );
  XNOR U30982 ( .A(n22341), .B(n22342), .Z(n22339) );
  XNOR U30983 ( .A(y[5200]), .B(x[5200]), .Z(n22342) );
  XNOR U30984 ( .A(y[5201]), .B(x[5201]), .Z(n22341) );
  NAND U30985 ( .A(n22406), .B(n22407), .Z(N63404) );
  NANDN U30986 ( .A(n22408), .B(n22409), .Z(n22407) );
  OR U30987 ( .A(n22410), .B(n22411), .Z(n22409) );
  NAND U30988 ( .A(n22410), .B(n22411), .Z(n22406) );
  XOR U30989 ( .A(n22410), .B(n22412), .Z(N63403) );
  XNOR U30990 ( .A(n22408), .B(n22411), .Z(n22412) );
  AND U30991 ( .A(n22413), .B(n22414), .Z(n22411) );
  NANDN U30992 ( .A(n22415), .B(n22416), .Z(n22414) );
  NANDN U30993 ( .A(n22417), .B(n22418), .Z(n22416) );
  NANDN U30994 ( .A(n22418), .B(n22417), .Z(n22413) );
  NAND U30995 ( .A(n22419), .B(n22420), .Z(n22408) );
  NANDN U30996 ( .A(n22421), .B(n22422), .Z(n22420) );
  OR U30997 ( .A(n22423), .B(n22424), .Z(n22422) );
  NAND U30998 ( .A(n22424), .B(n22423), .Z(n22419) );
  AND U30999 ( .A(n22425), .B(n22426), .Z(n22410) );
  NANDN U31000 ( .A(n22427), .B(n22428), .Z(n22426) );
  NANDN U31001 ( .A(n22429), .B(n22430), .Z(n22428) );
  NANDN U31002 ( .A(n22430), .B(n22429), .Z(n22425) );
  XOR U31003 ( .A(n22424), .B(n22431), .Z(N63402) );
  XOR U31004 ( .A(n22421), .B(n22423), .Z(n22431) );
  XNOR U31005 ( .A(n22417), .B(n22432), .Z(n22423) );
  XNOR U31006 ( .A(n22415), .B(n22418), .Z(n22432) );
  NAND U31007 ( .A(n22433), .B(n22434), .Z(n22418) );
  NAND U31008 ( .A(n22435), .B(n22436), .Z(n22434) );
  OR U31009 ( .A(n22437), .B(n22438), .Z(n22435) );
  NANDN U31010 ( .A(n22439), .B(n22437), .Z(n22433) );
  IV U31011 ( .A(n22438), .Z(n22439) );
  NAND U31012 ( .A(n22440), .B(n22441), .Z(n22415) );
  NAND U31013 ( .A(n22442), .B(n22443), .Z(n22441) );
  NANDN U31014 ( .A(n22444), .B(n22445), .Z(n22442) );
  NANDN U31015 ( .A(n22445), .B(n22444), .Z(n22440) );
  AND U31016 ( .A(n22446), .B(n22447), .Z(n22417) );
  NAND U31017 ( .A(n22448), .B(n22449), .Z(n22447) );
  OR U31018 ( .A(n22450), .B(n22451), .Z(n22448) );
  NANDN U31019 ( .A(n22452), .B(n22450), .Z(n22446) );
  NAND U31020 ( .A(n22453), .B(n22454), .Z(n22421) );
  NANDN U31021 ( .A(n22455), .B(n22456), .Z(n22454) );
  OR U31022 ( .A(n22457), .B(n22458), .Z(n22456) );
  NANDN U31023 ( .A(n22459), .B(n22457), .Z(n22453) );
  IV U31024 ( .A(n22458), .Z(n22459) );
  XNOR U31025 ( .A(n22429), .B(n22460), .Z(n22424) );
  XNOR U31026 ( .A(n22427), .B(n22430), .Z(n22460) );
  NAND U31027 ( .A(n22461), .B(n22462), .Z(n22430) );
  NAND U31028 ( .A(n22463), .B(n22464), .Z(n22462) );
  OR U31029 ( .A(n22465), .B(n22466), .Z(n22463) );
  NANDN U31030 ( .A(n22467), .B(n22465), .Z(n22461) );
  IV U31031 ( .A(n22466), .Z(n22467) );
  NAND U31032 ( .A(n22468), .B(n22469), .Z(n22427) );
  NAND U31033 ( .A(n22470), .B(n22471), .Z(n22469) );
  NANDN U31034 ( .A(n22472), .B(n22473), .Z(n22470) );
  NANDN U31035 ( .A(n22473), .B(n22472), .Z(n22468) );
  AND U31036 ( .A(n22474), .B(n22475), .Z(n22429) );
  NAND U31037 ( .A(n22476), .B(n22477), .Z(n22475) );
  OR U31038 ( .A(n22478), .B(n22479), .Z(n22476) );
  NANDN U31039 ( .A(n22480), .B(n22478), .Z(n22474) );
  XNOR U31040 ( .A(n22455), .B(n22481), .Z(N63401) );
  XOR U31041 ( .A(n22457), .B(n22458), .Z(n22481) );
  XNOR U31042 ( .A(n22471), .B(n22482), .Z(n22458) );
  XOR U31043 ( .A(n22472), .B(n22473), .Z(n22482) );
  XOR U31044 ( .A(n22478), .B(n22483), .Z(n22473) );
  XOR U31045 ( .A(n22477), .B(n22480), .Z(n22483) );
  IV U31046 ( .A(n22479), .Z(n22480) );
  NAND U31047 ( .A(n22484), .B(n22485), .Z(n22479) );
  OR U31048 ( .A(n22486), .B(n22487), .Z(n22485) );
  OR U31049 ( .A(n22488), .B(n22489), .Z(n22484) );
  NAND U31050 ( .A(n22490), .B(n22491), .Z(n22477) );
  OR U31051 ( .A(n22492), .B(n22493), .Z(n22491) );
  OR U31052 ( .A(n22494), .B(n22495), .Z(n22490) );
  NOR U31053 ( .A(n22496), .B(n22497), .Z(n22478) );
  ANDN U31054 ( .B(n22498), .A(n22499), .Z(n22472) );
  XNOR U31055 ( .A(n22465), .B(n22500), .Z(n22471) );
  XNOR U31056 ( .A(n22464), .B(n22466), .Z(n22500) );
  NAND U31057 ( .A(n22501), .B(n22502), .Z(n22466) );
  OR U31058 ( .A(n22503), .B(n22504), .Z(n22502) );
  OR U31059 ( .A(n22505), .B(n22506), .Z(n22501) );
  NAND U31060 ( .A(n22507), .B(n22508), .Z(n22464) );
  OR U31061 ( .A(n22509), .B(n22510), .Z(n22508) );
  OR U31062 ( .A(n22511), .B(n22512), .Z(n22507) );
  ANDN U31063 ( .B(n22513), .A(n22514), .Z(n22465) );
  IV U31064 ( .A(n22515), .Z(n22513) );
  ANDN U31065 ( .B(n22516), .A(n22517), .Z(n22457) );
  XOR U31066 ( .A(n22443), .B(n22518), .Z(n22455) );
  XOR U31067 ( .A(n22444), .B(n22445), .Z(n22518) );
  XOR U31068 ( .A(n22450), .B(n22519), .Z(n22445) );
  XOR U31069 ( .A(n22449), .B(n22452), .Z(n22519) );
  IV U31070 ( .A(n22451), .Z(n22452) );
  NAND U31071 ( .A(n22520), .B(n22521), .Z(n22451) );
  OR U31072 ( .A(n22522), .B(n22523), .Z(n22521) );
  OR U31073 ( .A(n22524), .B(n22525), .Z(n22520) );
  NAND U31074 ( .A(n22526), .B(n22527), .Z(n22449) );
  OR U31075 ( .A(n22528), .B(n22529), .Z(n22527) );
  OR U31076 ( .A(n22530), .B(n22531), .Z(n22526) );
  NOR U31077 ( .A(n22532), .B(n22533), .Z(n22450) );
  ANDN U31078 ( .B(n22534), .A(n22535), .Z(n22444) );
  IV U31079 ( .A(n22536), .Z(n22534) );
  XNOR U31080 ( .A(n22437), .B(n22537), .Z(n22443) );
  XNOR U31081 ( .A(n22436), .B(n22438), .Z(n22537) );
  NAND U31082 ( .A(n22538), .B(n22539), .Z(n22438) );
  OR U31083 ( .A(n22540), .B(n22541), .Z(n22539) );
  OR U31084 ( .A(n22542), .B(n22543), .Z(n22538) );
  NAND U31085 ( .A(n22544), .B(n22545), .Z(n22436) );
  OR U31086 ( .A(n22546), .B(n22547), .Z(n22545) );
  OR U31087 ( .A(n22548), .B(n22549), .Z(n22544) );
  ANDN U31088 ( .B(n22550), .A(n22551), .Z(n22437) );
  IV U31089 ( .A(n22552), .Z(n22550) );
  XNOR U31090 ( .A(n22517), .B(n22516), .Z(N63400) );
  XOR U31091 ( .A(n22536), .B(n22535), .Z(n22516) );
  XNOR U31092 ( .A(n22551), .B(n22552), .Z(n22535) );
  XNOR U31093 ( .A(n22546), .B(n22547), .Z(n22552) );
  XNOR U31094 ( .A(n22548), .B(n22549), .Z(n22547) );
  XNOR U31095 ( .A(y[5197]), .B(x[5197]), .Z(n22549) );
  XNOR U31096 ( .A(y[5198]), .B(x[5198]), .Z(n22548) );
  XNOR U31097 ( .A(y[5196]), .B(x[5196]), .Z(n22546) );
  XNOR U31098 ( .A(n22540), .B(n22541), .Z(n22551) );
  XNOR U31099 ( .A(y[5193]), .B(x[5193]), .Z(n22541) );
  XNOR U31100 ( .A(n22542), .B(n22543), .Z(n22540) );
  XNOR U31101 ( .A(y[5194]), .B(x[5194]), .Z(n22543) );
  XNOR U31102 ( .A(y[5195]), .B(x[5195]), .Z(n22542) );
  XNOR U31103 ( .A(n22533), .B(n22532), .Z(n22536) );
  XNOR U31104 ( .A(n22528), .B(n22529), .Z(n22532) );
  XNOR U31105 ( .A(y[5190]), .B(x[5190]), .Z(n22529) );
  XNOR U31106 ( .A(n22530), .B(n22531), .Z(n22528) );
  XNOR U31107 ( .A(y[5191]), .B(x[5191]), .Z(n22531) );
  XNOR U31108 ( .A(y[5192]), .B(x[5192]), .Z(n22530) );
  XNOR U31109 ( .A(n22522), .B(n22523), .Z(n22533) );
  XNOR U31110 ( .A(y[5187]), .B(x[5187]), .Z(n22523) );
  XNOR U31111 ( .A(n22524), .B(n22525), .Z(n22522) );
  XNOR U31112 ( .A(y[5188]), .B(x[5188]), .Z(n22525) );
  XNOR U31113 ( .A(y[5189]), .B(x[5189]), .Z(n22524) );
  XOR U31114 ( .A(n22498), .B(n22499), .Z(n22517) );
  XNOR U31115 ( .A(n22514), .B(n22515), .Z(n22499) );
  XNOR U31116 ( .A(n22509), .B(n22510), .Z(n22515) );
  XNOR U31117 ( .A(n22511), .B(n22512), .Z(n22510) );
  XNOR U31118 ( .A(y[5185]), .B(x[5185]), .Z(n22512) );
  XNOR U31119 ( .A(y[5186]), .B(x[5186]), .Z(n22511) );
  XNOR U31120 ( .A(y[5184]), .B(x[5184]), .Z(n22509) );
  XNOR U31121 ( .A(n22503), .B(n22504), .Z(n22514) );
  XNOR U31122 ( .A(y[5181]), .B(x[5181]), .Z(n22504) );
  XNOR U31123 ( .A(n22505), .B(n22506), .Z(n22503) );
  XNOR U31124 ( .A(y[5182]), .B(x[5182]), .Z(n22506) );
  XNOR U31125 ( .A(y[5183]), .B(x[5183]), .Z(n22505) );
  XOR U31126 ( .A(n22497), .B(n22496), .Z(n22498) );
  XNOR U31127 ( .A(n22492), .B(n22493), .Z(n22496) );
  XNOR U31128 ( .A(y[5178]), .B(x[5178]), .Z(n22493) );
  XNOR U31129 ( .A(n22494), .B(n22495), .Z(n22492) );
  XNOR U31130 ( .A(y[5179]), .B(x[5179]), .Z(n22495) );
  XNOR U31131 ( .A(y[5180]), .B(x[5180]), .Z(n22494) );
  XNOR U31132 ( .A(n22486), .B(n22487), .Z(n22497) );
  XNOR U31133 ( .A(y[5175]), .B(x[5175]), .Z(n22487) );
  XNOR U31134 ( .A(n22488), .B(n22489), .Z(n22486) );
  XNOR U31135 ( .A(y[5176]), .B(x[5176]), .Z(n22489) );
  XNOR U31136 ( .A(y[5177]), .B(x[5177]), .Z(n22488) );
  NAND U31137 ( .A(n22553), .B(n22554), .Z(N63391) );
  NANDN U31138 ( .A(n22555), .B(n22556), .Z(n22554) );
  OR U31139 ( .A(n22557), .B(n22558), .Z(n22556) );
  NAND U31140 ( .A(n22557), .B(n22558), .Z(n22553) );
  XOR U31141 ( .A(n22557), .B(n22559), .Z(N63390) );
  XNOR U31142 ( .A(n22555), .B(n22558), .Z(n22559) );
  AND U31143 ( .A(n22560), .B(n22561), .Z(n22558) );
  NANDN U31144 ( .A(n22562), .B(n22563), .Z(n22561) );
  NANDN U31145 ( .A(n22564), .B(n22565), .Z(n22563) );
  NANDN U31146 ( .A(n22565), .B(n22564), .Z(n22560) );
  NAND U31147 ( .A(n22566), .B(n22567), .Z(n22555) );
  NANDN U31148 ( .A(n22568), .B(n22569), .Z(n22567) );
  OR U31149 ( .A(n22570), .B(n22571), .Z(n22569) );
  NAND U31150 ( .A(n22571), .B(n22570), .Z(n22566) );
  AND U31151 ( .A(n22572), .B(n22573), .Z(n22557) );
  NANDN U31152 ( .A(n22574), .B(n22575), .Z(n22573) );
  NANDN U31153 ( .A(n22576), .B(n22577), .Z(n22575) );
  NANDN U31154 ( .A(n22577), .B(n22576), .Z(n22572) );
  XOR U31155 ( .A(n22571), .B(n22578), .Z(N63389) );
  XOR U31156 ( .A(n22568), .B(n22570), .Z(n22578) );
  XNOR U31157 ( .A(n22564), .B(n22579), .Z(n22570) );
  XNOR U31158 ( .A(n22562), .B(n22565), .Z(n22579) );
  NAND U31159 ( .A(n22580), .B(n22581), .Z(n22565) );
  NAND U31160 ( .A(n22582), .B(n22583), .Z(n22581) );
  OR U31161 ( .A(n22584), .B(n22585), .Z(n22582) );
  NANDN U31162 ( .A(n22586), .B(n22584), .Z(n22580) );
  IV U31163 ( .A(n22585), .Z(n22586) );
  NAND U31164 ( .A(n22587), .B(n22588), .Z(n22562) );
  NAND U31165 ( .A(n22589), .B(n22590), .Z(n22588) );
  NANDN U31166 ( .A(n22591), .B(n22592), .Z(n22589) );
  NANDN U31167 ( .A(n22592), .B(n22591), .Z(n22587) );
  AND U31168 ( .A(n22593), .B(n22594), .Z(n22564) );
  NAND U31169 ( .A(n22595), .B(n22596), .Z(n22594) );
  OR U31170 ( .A(n22597), .B(n22598), .Z(n22595) );
  NANDN U31171 ( .A(n22599), .B(n22597), .Z(n22593) );
  NAND U31172 ( .A(n22600), .B(n22601), .Z(n22568) );
  NANDN U31173 ( .A(n22602), .B(n22603), .Z(n22601) );
  OR U31174 ( .A(n22604), .B(n22605), .Z(n22603) );
  NANDN U31175 ( .A(n22606), .B(n22604), .Z(n22600) );
  IV U31176 ( .A(n22605), .Z(n22606) );
  XNOR U31177 ( .A(n22576), .B(n22607), .Z(n22571) );
  XNOR U31178 ( .A(n22574), .B(n22577), .Z(n22607) );
  NAND U31179 ( .A(n22608), .B(n22609), .Z(n22577) );
  NAND U31180 ( .A(n22610), .B(n22611), .Z(n22609) );
  OR U31181 ( .A(n22612), .B(n22613), .Z(n22610) );
  NANDN U31182 ( .A(n22614), .B(n22612), .Z(n22608) );
  IV U31183 ( .A(n22613), .Z(n22614) );
  NAND U31184 ( .A(n22615), .B(n22616), .Z(n22574) );
  NAND U31185 ( .A(n22617), .B(n22618), .Z(n22616) );
  NANDN U31186 ( .A(n22619), .B(n22620), .Z(n22617) );
  NANDN U31187 ( .A(n22620), .B(n22619), .Z(n22615) );
  AND U31188 ( .A(n22621), .B(n22622), .Z(n22576) );
  NAND U31189 ( .A(n22623), .B(n22624), .Z(n22622) );
  OR U31190 ( .A(n22625), .B(n22626), .Z(n22623) );
  NANDN U31191 ( .A(n22627), .B(n22625), .Z(n22621) );
  XNOR U31192 ( .A(n22602), .B(n22628), .Z(N63388) );
  XOR U31193 ( .A(n22604), .B(n22605), .Z(n22628) );
  XNOR U31194 ( .A(n22618), .B(n22629), .Z(n22605) );
  XOR U31195 ( .A(n22619), .B(n22620), .Z(n22629) );
  XOR U31196 ( .A(n22625), .B(n22630), .Z(n22620) );
  XOR U31197 ( .A(n22624), .B(n22627), .Z(n22630) );
  IV U31198 ( .A(n22626), .Z(n22627) );
  NAND U31199 ( .A(n22631), .B(n22632), .Z(n22626) );
  OR U31200 ( .A(n22633), .B(n22634), .Z(n22632) );
  OR U31201 ( .A(n22635), .B(n22636), .Z(n22631) );
  NAND U31202 ( .A(n22637), .B(n22638), .Z(n22624) );
  OR U31203 ( .A(n22639), .B(n22640), .Z(n22638) );
  OR U31204 ( .A(n22641), .B(n22642), .Z(n22637) );
  NOR U31205 ( .A(n22643), .B(n22644), .Z(n22625) );
  ANDN U31206 ( .B(n22645), .A(n22646), .Z(n22619) );
  XNOR U31207 ( .A(n22612), .B(n22647), .Z(n22618) );
  XNOR U31208 ( .A(n22611), .B(n22613), .Z(n22647) );
  NAND U31209 ( .A(n22648), .B(n22649), .Z(n22613) );
  OR U31210 ( .A(n22650), .B(n22651), .Z(n22649) );
  OR U31211 ( .A(n22652), .B(n22653), .Z(n22648) );
  NAND U31212 ( .A(n22654), .B(n22655), .Z(n22611) );
  OR U31213 ( .A(n22656), .B(n22657), .Z(n22655) );
  OR U31214 ( .A(n22658), .B(n22659), .Z(n22654) );
  ANDN U31215 ( .B(n22660), .A(n22661), .Z(n22612) );
  IV U31216 ( .A(n22662), .Z(n22660) );
  ANDN U31217 ( .B(n22663), .A(n22664), .Z(n22604) );
  XOR U31218 ( .A(n22590), .B(n22665), .Z(n22602) );
  XOR U31219 ( .A(n22591), .B(n22592), .Z(n22665) );
  XOR U31220 ( .A(n22597), .B(n22666), .Z(n22592) );
  XOR U31221 ( .A(n22596), .B(n22599), .Z(n22666) );
  IV U31222 ( .A(n22598), .Z(n22599) );
  NAND U31223 ( .A(n22667), .B(n22668), .Z(n22598) );
  OR U31224 ( .A(n22669), .B(n22670), .Z(n22668) );
  OR U31225 ( .A(n22671), .B(n22672), .Z(n22667) );
  NAND U31226 ( .A(n22673), .B(n22674), .Z(n22596) );
  OR U31227 ( .A(n22675), .B(n22676), .Z(n22674) );
  OR U31228 ( .A(n22677), .B(n22678), .Z(n22673) );
  NOR U31229 ( .A(n22679), .B(n22680), .Z(n22597) );
  ANDN U31230 ( .B(n22681), .A(n22682), .Z(n22591) );
  IV U31231 ( .A(n22683), .Z(n22681) );
  XNOR U31232 ( .A(n22584), .B(n22684), .Z(n22590) );
  XNOR U31233 ( .A(n22583), .B(n22585), .Z(n22684) );
  NAND U31234 ( .A(n22685), .B(n22686), .Z(n22585) );
  OR U31235 ( .A(n22687), .B(n22688), .Z(n22686) );
  OR U31236 ( .A(n22689), .B(n22690), .Z(n22685) );
  NAND U31237 ( .A(n22691), .B(n22692), .Z(n22583) );
  OR U31238 ( .A(n22693), .B(n22694), .Z(n22692) );
  OR U31239 ( .A(n22695), .B(n22696), .Z(n22691) );
  ANDN U31240 ( .B(n22697), .A(n22698), .Z(n22584) );
  IV U31241 ( .A(n22699), .Z(n22697) );
  XNOR U31242 ( .A(n22664), .B(n22663), .Z(N63387) );
  XOR U31243 ( .A(n22683), .B(n22682), .Z(n22663) );
  XNOR U31244 ( .A(n22698), .B(n22699), .Z(n22682) );
  XNOR U31245 ( .A(n22693), .B(n22694), .Z(n22699) );
  XNOR U31246 ( .A(n22695), .B(n22696), .Z(n22694) );
  XNOR U31247 ( .A(y[5173]), .B(x[5173]), .Z(n22696) );
  XNOR U31248 ( .A(y[5174]), .B(x[5174]), .Z(n22695) );
  XNOR U31249 ( .A(y[5172]), .B(x[5172]), .Z(n22693) );
  XNOR U31250 ( .A(n22687), .B(n22688), .Z(n22698) );
  XNOR U31251 ( .A(y[5169]), .B(x[5169]), .Z(n22688) );
  XNOR U31252 ( .A(n22689), .B(n22690), .Z(n22687) );
  XNOR U31253 ( .A(y[5170]), .B(x[5170]), .Z(n22690) );
  XNOR U31254 ( .A(y[5171]), .B(x[5171]), .Z(n22689) );
  XNOR U31255 ( .A(n22680), .B(n22679), .Z(n22683) );
  XNOR U31256 ( .A(n22675), .B(n22676), .Z(n22679) );
  XNOR U31257 ( .A(y[5166]), .B(x[5166]), .Z(n22676) );
  XNOR U31258 ( .A(n22677), .B(n22678), .Z(n22675) );
  XNOR U31259 ( .A(y[5167]), .B(x[5167]), .Z(n22678) );
  XNOR U31260 ( .A(y[5168]), .B(x[5168]), .Z(n22677) );
  XNOR U31261 ( .A(n22669), .B(n22670), .Z(n22680) );
  XNOR U31262 ( .A(y[5163]), .B(x[5163]), .Z(n22670) );
  XNOR U31263 ( .A(n22671), .B(n22672), .Z(n22669) );
  XNOR U31264 ( .A(y[5164]), .B(x[5164]), .Z(n22672) );
  XNOR U31265 ( .A(y[5165]), .B(x[5165]), .Z(n22671) );
  XOR U31266 ( .A(n22645), .B(n22646), .Z(n22664) );
  XNOR U31267 ( .A(n22661), .B(n22662), .Z(n22646) );
  XNOR U31268 ( .A(n22656), .B(n22657), .Z(n22662) );
  XNOR U31269 ( .A(n22658), .B(n22659), .Z(n22657) );
  XNOR U31270 ( .A(y[5161]), .B(x[5161]), .Z(n22659) );
  XNOR U31271 ( .A(y[5162]), .B(x[5162]), .Z(n22658) );
  XNOR U31272 ( .A(y[5160]), .B(x[5160]), .Z(n22656) );
  XNOR U31273 ( .A(n22650), .B(n22651), .Z(n22661) );
  XNOR U31274 ( .A(y[5157]), .B(x[5157]), .Z(n22651) );
  XNOR U31275 ( .A(n22652), .B(n22653), .Z(n22650) );
  XNOR U31276 ( .A(y[5158]), .B(x[5158]), .Z(n22653) );
  XNOR U31277 ( .A(y[5159]), .B(x[5159]), .Z(n22652) );
  XOR U31278 ( .A(n22644), .B(n22643), .Z(n22645) );
  XNOR U31279 ( .A(n22639), .B(n22640), .Z(n22643) );
  XNOR U31280 ( .A(y[5154]), .B(x[5154]), .Z(n22640) );
  XNOR U31281 ( .A(n22641), .B(n22642), .Z(n22639) );
  XNOR U31282 ( .A(y[5155]), .B(x[5155]), .Z(n22642) );
  XNOR U31283 ( .A(y[5156]), .B(x[5156]), .Z(n22641) );
  XNOR U31284 ( .A(n22633), .B(n22634), .Z(n22644) );
  XNOR U31285 ( .A(y[5151]), .B(x[5151]), .Z(n22634) );
  XNOR U31286 ( .A(n22635), .B(n22636), .Z(n22633) );
  XNOR U31287 ( .A(y[5152]), .B(x[5152]), .Z(n22636) );
  XNOR U31288 ( .A(y[5153]), .B(x[5153]), .Z(n22635) );
  NAND U31289 ( .A(n22700), .B(n22701), .Z(N63378) );
  NANDN U31290 ( .A(n22702), .B(n22703), .Z(n22701) );
  OR U31291 ( .A(n22704), .B(n22705), .Z(n22703) );
  NAND U31292 ( .A(n22704), .B(n22705), .Z(n22700) );
  XOR U31293 ( .A(n22704), .B(n22706), .Z(N63377) );
  XNOR U31294 ( .A(n22702), .B(n22705), .Z(n22706) );
  AND U31295 ( .A(n22707), .B(n22708), .Z(n22705) );
  NANDN U31296 ( .A(n22709), .B(n22710), .Z(n22708) );
  NANDN U31297 ( .A(n22711), .B(n22712), .Z(n22710) );
  NANDN U31298 ( .A(n22712), .B(n22711), .Z(n22707) );
  NAND U31299 ( .A(n22713), .B(n22714), .Z(n22702) );
  NANDN U31300 ( .A(n22715), .B(n22716), .Z(n22714) );
  OR U31301 ( .A(n22717), .B(n22718), .Z(n22716) );
  NAND U31302 ( .A(n22718), .B(n22717), .Z(n22713) );
  AND U31303 ( .A(n22719), .B(n22720), .Z(n22704) );
  NANDN U31304 ( .A(n22721), .B(n22722), .Z(n22720) );
  NANDN U31305 ( .A(n22723), .B(n22724), .Z(n22722) );
  NANDN U31306 ( .A(n22724), .B(n22723), .Z(n22719) );
  XOR U31307 ( .A(n22718), .B(n22725), .Z(N63376) );
  XOR U31308 ( .A(n22715), .B(n22717), .Z(n22725) );
  XNOR U31309 ( .A(n22711), .B(n22726), .Z(n22717) );
  XNOR U31310 ( .A(n22709), .B(n22712), .Z(n22726) );
  NAND U31311 ( .A(n22727), .B(n22728), .Z(n22712) );
  NAND U31312 ( .A(n22729), .B(n22730), .Z(n22728) );
  OR U31313 ( .A(n22731), .B(n22732), .Z(n22729) );
  NANDN U31314 ( .A(n22733), .B(n22731), .Z(n22727) );
  IV U31315 ( .A(n22732), .Z(n22733) );
  NAND U31316 ( .A(n22734), .B(n22735), .Z(n22709) );
  NAND U31317 ( .A(n22736), .B(n22737), .Z(n22735) );
  NANDN U31318 ( .A(n22738), .B(n22739), .Z(n22736) );
  NANDN U31319 ( .A(n22739), .B(n22738), .Z(n22734) );
  AND U31320 ( .A(n22740), .B(n22741), .Z(n22711) );
  NAND U31321 ( .A(n22742), .B(n22743), .Z(n22741) );
  OR U31322 ( .A(n22744), .B(n22745), .Z(n22742) );
  NANDN U31323 ( .A(n22746), .B(n22744), .Z(n22740) );
  NAND U31324 ( .A(n22747), .B(n22748), .Z(n22715) );
  NANDN U31325 ( .A(n22749), .B(n22750), .Z(n22748) );
  OR U31326 ( .A(n22751), .B(n22752), .Z(n22750) );
  NANDN U31327 ( .A(n22753), .B(n22751), .Z(n22747) );
  IV U31328 ( .A(n22752), .Z(n22753) );
  XNOR U31329 ( .A(n22723), .B(n22754), .Z(n22718) );
  XNOR U31330 ( .A(n22721), .B(n22724), .Z(n22754) );
  NAND U31331 ( .A(n22755), .B(n22756), .Z(n22724) );
  NAND U31332 ( .A(n22757), .B(n22758), .Z(n22756) );
  OR U31333 ( .A(n22759), .B(n22760), .Z(n22757) );
  NANDN U31334 ( .A(n22761), .B(n22759), .Z(n22755) );
  IV U31335 ( .A(n22760), .Z(n22761) );
  NAND U31336 ( .A(n22762), .B(n22763), .Z(n22721) );
  NAND U31337 ( .A(n22764), .B(n22765), .Z(n22763) );
  NANDN U31338 ( .A(n22766), .B(n22767), .Z(n22764) );
  NANDN U31339 ( .A(n22767), .B(n22766), .Z(n22762) );
  AND U31340 ( .A(n22768), .B(n22769), .Z(n22723) );
  NAND U31341 ( .A(n22770), .B(n22771), .Z(n22769) );
  OR U31342 ( .A(n22772), .B(n22773), .Z(n22770) );
  NANDN U31343 ( .A(n22774), .B(n22772), .Z(n22768) );
  XNOR U31344 ( .A(n22749), .B(n22775), .Z(N63375) );
  XOR U31345 ( .A(n22751), .B(n22752), .Z(n22775) );
  XNOR U31346 ( .A(n22765), .B(n22776), .Z(n22752) );
  XOR U31347 ( .A(n22766), .B(n22767), .Z(n22776) );
  XOR U31348 ( .A(n22772), .B(n22777), .Z(n22767) );
  XOR U31349 ( .A(n22771), .B(n22774), .Z(n22777) );
  IV U31350 ( .A(n22773), .Z(n22774) );
  NAND U31351 ( .A(n22778), .B(n22779), .Z(n22773) );
  OR U31352 ( .A(n22780), .B(n22781), .Z(n22779) );
  OR U31353 ( .A(n22782), .B(n22783), .Z(n22778) );
  NAND U31354 ( .A(n22784), .B(n22785), .Z(n22771) );
  OR U31355 ( .A(n22786), .B(n22787), .Z(n22785) );
  OR U31356 ( .A(n22788), .B(n22789), .Z(n22784) );
  NOR U31357 ( .A(n22790), .B(n22791), .Z(n22772) );
  ANDN U31358 ( .B(n22792), .A(n22793), .Z(n22766) );
  XNOR U31359 ( .A(n22759), .B(n22794), .Z(n22765) );
  XNOR U31360 ( .A(n22758), .B(n22760), .Z(n22794) );
  NAND U31361 ( .A(n22795), .B(n22796), .Z(n22760) );
  OR U31362 ( .A(n22797), .B(n22798), .Z(n22796) );
  OR U31363 ( .A(n22799), .B(n22800), .Z(n22795) );
  NAND U31364 ( .A(n22801), .B(n22802), .Z(n22758) );
  OR U31365 ( .A(n22803), .B(n22804), .Z(n22802) );
  OR U31366 ( .A(n22805), .B(n22806), .Z(n22801) );
  ANDN U31367 ( .B(n22807), .A(n22808), .Z(n22759) );
  IV U31368 ( .A(n22809), .Z(n22807) );
  ANDN U31369 ( .B(n22810), .A(n22811), .Z(n22751) );
  XOR U31370 ( .A(n22737), .B(n22812), .Z(n22749) );
  XOR U31371 ( .A(n22738), .B(n22739), .Z(n22812) );
  XOR U31372 ( .A(n22744), .B(n22813), .Z(n22739) );
  XOR U31373 ( .A(n22743), .B(n22746), .Z(n22813) );
  IV U31374 ( .A(n22745), .Z(n22746) );
  NAND U31375 ( .A(n22814), .B(n22815), .Z(n22745) );
  OR U31376 ( .A(n22816), .B(n22817), .Z(n22815) );
  OR U31377 ( .A(n22818), .B(n22819), .Z(n22814) );
  NAND U31378 ( .A(n22820), .B(n22821), .Z(n22743) );
  OR U31379 ( .A(n22822), .B(n22823), .Z(n22821) );
  OR U31380 ( .A(n22824), .B(n22825), .Z(n22820) );
  NOR U31381 ( .A(n22826), .B(n22827), .Z(n22744) );
  ANDN U31382 ( .B(n22828), .A(n22829), .Z(n22738) );
  IV U31383 ( .A(n22830), .Z(n22828) );
  XNOR U31384 ( .A(n22731), .B(n22831), .Z(n22737) );
  XNOR U31385 ( .A(n22730), .B(n22732), .Z(n22831) );
  NAND U31386 ( .A(n22832), .B(n22833), .Z(n22732) );
  OR U31387 ( .A(n22834), .B(n22835), .Z(n22833) );
  OR U31388 ( .A(n22836), .B(n22837), .Z(n22832) );
  NAND U31389 ( .A(n22838), .B(n22839), .Z(n22730) );
  OR U31390 ( .A(n22840), .B(n22841), .Z(n22839) );
  OR U31391 ( .A(n22842), .B(n22843), .Z(n22838) );
  ANDN U31392 ( .B(n22844), .A(n22845), .Z(n22731) );
  IV U31393 ( .A(n22846), .Z(n22844) );
  XNOR U31394 ( .A(n22811), .B(n22810), .Z(N63374) );
  XOR U31395 ( .A(n22830), .B(n22829), .Z(n22810) );
  XNOR U31396 ( .A(n22845), .B(n22846), .Z(n22829) );
  XNOR U31397 ( .A(n22840), .B(n22841), .Z(n22846) );
  XNOR U31398 ( .A(n22842), .B(n22843), .Z(n22841) );
  XNOR U31399 ( .A(y[5149]), .B(x[5149]), .Z(n22843) );
  XNOR U31400 ( .A(y[5150]), .B(x[5150]), .Z(n22842) );
  XNOR U31401 ( .A(y[5148]), .B(x[5148]), .Z(n22840) );
  XNOR U31402 ( .A(n22834), .B(n22835), .Z(n22845) );
  XNOR U31403 ( .A(y[5145]), .B(x[5145]), .Z(n22835) );
  XNOR U31404 ( .A(n22836), .B(n22837), .Z(n22834) );
  XNOR U31405 ( .A(y[5146]), .B(x[5146]), .Z(n22837) );
  XNOR U31406 ( .A(y[5147]), .B(x[5147]), .Z(n22836) );
  XNOR U31407 ( .A(n22827), .B(n22826), .Z(n22830) );
  XNOR U31408 ( .A(n22822), .B(n22823), .Z(n22826) );
  XNOR U31409 ( .A(y[5142]), .B(x[5142]), .Z(n22823) );
  XNOR U31410 ( .A(n22824), .B(n22825), .Z(n22822) );
  XNOR U31411 ( .A(y[5143]), .B(x[5143]), .Z(n22825) );
  XNOR U31412 ( .A(y[5144]), .B(x[5144]), .Z(n22824) );
  XNOR U31413 ( .A(n22816), .B(n22817), .Z(n22827) );
  XNOR U31414 ( .A(y[5139]), .B(x[5139]), .Z(n22817) );
  XNOR U31415 ( .A(n22818), .B(n22819), .Z(n22816) );
  XNOR U31416 ( .A(y[5140]), .B(x[5140]), .Z(n22819) );
  XNOR U31417 ( .A(y[5141]), .B(x[5141]), .Z(n22818) );
  XOR U31418 ( .A(n22792), .B(n22793), .Z(n22811) );
  XNOR U31419 ( .A(n22808), .B(n22809), .Z(n22793) );
  XNOR U31420 ( .A(n22803), .B(n22804), .Z(n22809) );
  XNOR U31421 ( .A(n22805), .B(n22806), .Z(n22804) );
  XNOR U31422 ( .A(y[5137]), .B(x[5137]), .Z(n22806) );
  XNOR U31423 ( .A(y[5138]), .B(x[5138]), .Z(n22805) );
  XNOR U31424 ( .A(y[5136]), .B(x[5136]), .Z(n22803) );
  XNOR U31425 ( .A(n22797), .B(n22798), .Z(n22808) );
  XNOR U31426 ( .A(y[5133]), .B(x[5133]), .Z(n22798) );
  XNOR U31427 ( .A(n22799), .B(n22800), .Z(n22797) );
  XNOR U31428 ( .A(y[5134]), .B(x[5134]), .Z(n22800) );
  XNOR U31429 ( .A(y[5135]), .B(x[5135]), .Z(n22799) );
  XOR U31430 ( .A(n22791), .B(n22790), .Z(n22792) );
  XNOR U31431 ( .A(n22786), .B(n22787), .Z(n22790) );
  XNOR U31432 ( .A(y[5130]), .B(x[5130]), .Z(n22787) );
  XNOR U31433 ( .A(n22788), .B(n22789), .Z(n22786) );
  XNOR U31434 ( .A(y[5131]), .B(x[5131]), .Z(n22789) );
  XNOR U31435 ( .A(y[5132]), .B(x[5132]), .Z(n22788) );
  XNOR U31436 ( .A(n22780), .B(n22781), .Z(n22791) );
  XNOR U31437 ( .A(y[5127]), .B(x[5127]), .Z(n22781) );
  XNOR U31438 ( .A(n22782), .B(n22783), .Z(n22780) );
  XNOR U31439 ( .A(y[5128]), .B(x[5128]), .Z(n22783) );
  XNOR U31440 ( .A(y[5129]), .B(x[5129]), .Z(n22782) );
  NAND U31441 ( .A(n22847), .B(n22848), .Z(N63365) );
  NANDN U31442 ( .A(n22849), .B(n22850), .Z(n22848) );
  OR U31443 ( .A(n22851), .B(n22852), .Z(n22850) );
  NAND U31444 ( .A(n22851), .B(n22852), .Z(n22847) );
  XOR U31445 ( .A(n22851), .B(n22853), .Z(N63364) );
  XNOR U31446 ( .A(n22849), .B(n22852), .Z(n22853) );
  AND U31447 ( .A(n22854), .B(n22855), .Z(n22852) );
  NANDN U31448 ( .A(n22856), .B(n22857), .Z(n22855) );
  NANDN U31449 ( .A(n22858), .B(n22859), .Z(n22857) );
  NANDN U31450 ( .A(n22859), .B(n22858), .Z(n22854) );
  NAND U31451 ( .A(n22860), .B(n22861), .Z(n22849) );
  NANDN U31452 ( .A(n22862), .B(n22863), .Z(n22861) );
  OR U31453 ( .A(n22864), .B(n22865), .Z(n22863) );
  NAND U31454 ( .A(n22865), .B(n22864), .Z(n22860) );
  AND U31455 ( .A(n22866), .B(n22867), .Z(n22851) );
  NANDN U31456 ( .A(n22868), .B(n22869), .Z(n22867) );
  NANDN U31457 ( .A(n22870), .B(n22871), .Z(n22869) );
  NANDN U31458 ( .A(n22871), .B(n22870), .Z(n22866) );
  XOR U31459 ( .A(n22865), .B(n22872), .Z(N63363) );
  XOR U31460 ( .A(n22862), .B(n22864), .Z(n22872) );
  XNOR U31461 ( .A(n22858), .B(n22873), .Z(n22864) );
  XNOR U31462 ( .A(n22856), .B(n22859), .Z(n22873) );
  NAND U31463 ( .A(n22874), .B(n22875), .Z(n22859) );
  NAND U31464 ( .A(n22876), .B(n22877), .Z(n22875) );
  OR U31465 ( .A(n22878), .B(n22879), .Z(n22876) );
  NANDN U31466 ( .A(n22880), .B(n22878), .Z(n22874) );
  IV U31467 ( .A(n22879), .Z(n22880) );
  NAND U31468 ( .A(n22881), .B(n22882), .Z(n22856) );
  NAND U31469 ( .A(n22883), .B(n22884), .Z(n22882) );
  NANDN U31470 ( .A(n22885), .B(n22886), .Z(n22883) );
  NANDN U31471 ( .A(n22886), .B(n22885), .Z(n22881) );
  AND U31472 ( .A(n22887), .B(n22888), .Z(n22858) );
  NAND U31473 ( .A(n22889), .B(n22890), .Z(n22888) );
  OR U31474 ( .A(n22891), .B(n22892), .Z(n22889) );
  NANDN U31475 ( .A(n22893), .B(n22891), .Z(n22887) );
  NAND U31476 ( .A(n22894), .B(n22895), .Z(n22862) );
  NANDN U31477 ( .A(n22896), .B(n22897), .Z(n22895) );
  OR U31478 ( .A(n22898), .B(n22899), .Z(n22897) );
  NANDN U31479 ( .A(n22900), .B(n22898), .Z(n22894) );
  IV U31480 ( .A(n22899), .Z(n22900) );
  XNOR U31481 ( .A(n22870), .B(n22901), .Z(n22865) );
  XNOR U31482 ( .A(n22868), .B(n22871), .Z(n22901) );
  NAND U31483 ( .A(n22902), .B(n22903), .Z(n22871) );
  NAND U31484 ( .A(n22904), .B(n22905), .Z(n22903) );
  OR U31485 ( .A(n22906), .B(n22907), .Z(n22904) );
  NANDN U31486 ( .A(n22908), .B(n22906), .Z(n22902) );
  IV U31487 ( .A(n22907), .Z(n22908) );
  NAND U31488 ( .A(n22909), .B(n22910), .Z(n22868) );
  NAND U31489 ( .A(n22911), .B(n22912), .Z(n22910) );
  NANDN U31490 ( .A(n22913), .B(n22914), .Z(n22911) );
  NANDN U31491 ( .A(n22914), .B(n22913), .Z(n22909) );
  AND U31492 ( .A(n22915), .B(n22916), .Z(n22870) );
  NAND U31493 ( .A(n22917), .B(n22918), .Z(n22916) );
  OR U31494 ( .A(n22919), .B(n22920), .Z(n22917) );
  NANDN U31495 ( .A(n22921), .B(n22919), .Z(n22915) );
  XNOR U31496 ( .A(n22896), .B(n22922), .Z(N63362) );
  XOR U31497 ( .A(n22898), .B(n22899), .Z(n22922) );
  XNOR U31498 ( .A(n22912), .B(n22923), .Z(n22899) );
  XOR U31499 ( .A(n22913), .B(n22914), .Z(n22923) );
  XOR U31500 ( .A(n22919), .B(n22924), .Z(n22914) );
  XOR U31501 ( .A(n22918), .B(n22921), .Z(n22924) );
  IV U31502 ( .A(n22920), .Z(n22921) );
  NAND U31503 ( .A(n22925), .B(n22926), .Z(n22920) );
  OR U31504 ( .A(n22927), .B(n22928), .Z(n22926) );
  OR U31505 ( .A(n22929), .B(n22930), .Z(n22925) );
  NAND U31506 ( .A(n22931), .B(n22932), .Z(n22918) );
  OR U31507 ( .A(n22933), .B(n22934), .Z(n22932) );
  OR U31508 ( .A(n22935), .B(n22936), .Z(n22931) );
  NOR U31509 ( .A(n22937), .B(n22938), .Z(n22919) );
  ANDN U31510 ( .B(n22939), .A(n22940), .Z(n22913) );
  XNOR U31511 ( .A(n22906), .B(n22941), .Z(n22912) );
  XNOR U31512 ( .A(n22905), .B(n22907), .Z(n22941) );
  NAND U31513 ( .A(n22942), .B(n22943), .Z(n22907) );
  OR U31514 ( .A(n22944), .B(n22945), .Z(n22943) );
  OR U31515 ( .A(n22946), .B(n22947), .Z(n22942) );
  NAND U31516 ( .A(n22948), .B(n22949), .Z(n22905) );
  OR U31517 ( .A(n22950), .B(n22951), .Z(n22949) );
  OR U31518 ( .A(n22952), .B(n22953), .Z(n22948) );
  ANDN U31519 ( .B(n22954), .A(n22955), .Z(n22906) );
  IV U31520 ( .A(n22956), .Z(n22954) );
  ANDN U31521 ( .B(n22957), .A(n22958), .Z(n22898) );
  XOR U31522 ( .A(n22884), .B(n22959), .Z(n22896) );
  XOR U31523 ( .A(n22885), .B(n22886), .Z(n22959) );
  XOR U31524 ( .A(n22891), .B(n22960), .Z(n22886) );
  XOR U31525 ( .A(n22890), .B(n22893), .Z(n22960) );
  IV U31526 ( .A(n22892), .Z(n22893) );
  NAND U31527 ( .A(n22961), .B(n22962), .Z(n22892) );
  OR U31528 ( .A(n22963), .B(n22964), .Z(n22962) );
  OR U31529 ( .A(n22965), .B(n22966), .Z(n22961) );
  NAND U31530 ( .A(n22967), .B(n22968), .Z(n22890) );
  OR U31531 ( .A(n22969), .B(n22970), .Z(n22968) );
  OR U31532 ( .A(n22971), .B(n22972), .Z(n22967) );
  NOR U31533 ( .A(n22973), .B(n22974), .Z(n22891) );
  ANDN U31534 ( .B(n22975), .A(n22976), .Z(n22885) );
  IV U31535 ( .A(n22977), .Z(n22975) );
  XNOR U31536 ( .A(n22878), .B(n22978), .Z(n22884) );
  XNOR U31537 ( .A(n22877), .B(n22879), .Z(n22978) );
  NAND U31538 ( .A(n22979), .B(n22980), .Z(n22879) );
  OR U31539 ( .A(n22981), .B(n22982), .Z(n22980) );
  OR U31540 ( .A(n22983), .B(n22984), .Z(n22979) );
  NAND U31541 ( .A(n22985), .B(n22986), .Z(n22877) );
  OR U31542 ( .A(n22987), .B(n22988), .Z(n22986) );
  OR U31543 ( .A(n22989), .B(n22990), .Z(n22985) );
  ANDN U31544 ( .B(n22991), .A(n22992), .Z(n22878) );
  IV U31545 ( .A(n22993), .Z(n22991) );
  XNOR U31546 ( .A(n22958), .B(n22957), .Z(N63361) );
  XOR U31547 ( .A(n22977), .B(n22976), .Z(n22957) );
  XNOR U31548 ( .A(n22992), .B(n22993), .Z(n22976) );
  XNOR U31549 ( .A(n22987), .B(n22988), .Z(n22993) );
  XNOR U31550 ( .A(n22989), .B(n22990), .Z(n22988) );
  XNOR U31551 ( .A(y[5125]), .B(x[5125]), .Z(n22990) );
  XNOR U31552 ( .A(y[5126]), .B(x[5126]), .Z(n22989) );
  XNOR U31553 ( .A(y[5124]), .B(x[5124]), .Z(n22987) );
  XNOR U31554 ( .A(n22981), .B(n22982), .Z(n22992) );
  XNOR U31555 ( .A(y[5121]), .B(x[5121]), .Z(n22982) );
  XNOR U31556 ( .A(n22983), .B(n22984), .Z(n22981) );
  XNOR U31557 ( .A(y[5122]), .B(x[5122]), .Z(n22984) );
  XNOR U31558 ( .A(y[5123]), .B(x[5123]), .Z(n22983) );
  XNOR U31559 ( .A(n22974), .B(n22973), .Z(n22977) );
  XNOR U31560 ( .A(n22969), .B(n22970), .Z(n22973) );
  XNOR U31561 ( .A(y[5118]), .B(x[5118]), .Z(n22970) );
  XNOR U31562 ( .A(n22971), .B(n22972), .Z(n22969) );
  XNOR U31563 ( .A(y[5119]), .B(x[5119]), .Z(n22972) );
  XNOR U31564 ( .A(y[5120]), .B(x[5120]), .Z(n22971) );
  XNOR U31565 ( .A(n22963), .B(n22964), .Z(n22974) );
  XNOR U31566 ( .A(y[5115]), .B(x[5115]), .Z(n22964) );
  XNOR U31567 ( .A(n22965), .B(n22966), .Z(n22963) );
  XNOR U31568 ( .A(y[5116]), .B(x[5116]), .Z(n22966) );
  XNOR U31569 ( .A(y[5117]), .B(x[5117]), .Z(n22965) );
  XOR U31570 ( .A(n22939), .B(n22940), .Z(n22958) );
  XNOR U31571 ( .A(n22955), .B(n22956), .Z(n22940) );
  XNOR U31572 ( .A(n22950), .B(n22951), .Z(n22956) );
  XNOR U31573 ( .A(n22952), .B(n22953), .Z(n22951) );
  XNOR U31574 ( .A(y[5113]), .B(x[5113]), .Z(n22953) );
  XNOR U31575 ( .A(y[5114]), .B(x[5114]), .Z(n22952) );
  XNOR U31576 ( .A(y[5112]), .B(x[5112]), .Z(n22950) );
  XNOR U31577 ( .A(n22944), .B(n22945), .Z(n22955) );
  XNOR U31578 ( .A(y[5109]), .B(x[5109]), .Z(n22945) );
  XNOR U31579 ( .A(n22946), .B(n22947), .Z(n22944) );
  XNOR U31580 ( .A(y[5110]), .B(x[5110]), .Z(n22947) );
  XNOR U31581 ( .A(y[5111]), .B(x[5111]), .Z(n22946) );
  XOR U31582 ( .A(n22938), .B(n22937), .Z(n22939) );
  XNOR U31583 ( .A(n22933), .B(n22934), .Z(n22937) );
  XNOR U31584 ( .A(y[5106]), .B(x[5106]), .Z(n22934) );
  XNOR U31585 ( .A(n22935), .B(n22936), .Z(n22933) );
  XNOR U31586 ( .A(y[5107]), .B(x[5107]), .Z(n22936) );
  XNOR U31587 ( .A(y[5108]), .B(x[5108]), .Z(n22935) );
  XNOR U31588 ( .A(n22927), .B(n22928), .Z(n22938) );
  XNOR U31589 ( .A(y[5103]), .B(x[5103]), .Z(n22928) );
  XNOR U31590 ( .A(n22929), .B(n22930), .Z(n22927) );
  XNOR U31591 ( .A(y[5104]), .B(x[5104]), .Z(n22930) );
  XNOR U31592 ( .A(y[5105]), .B(x[5105]), .Z(n22929) );
  NAND U31593 ( .A(n22994), .B(n22995), .Z(N63352) );
  NANDN U31594 ( .A(n22996), .B(n22997), .Z(n22995) );
  OR U31595 ( .A(n22998), .B(n22999), .Z(n22997) );
  NAND U31596 ( .A(n22998), .B(n22999), .Z(n22994) );
  XOR U31597 ( .A(n22998), .B(n23000), .Z(N63351) );
  XNOR U31598 ( .A(n22996), .B(n22999), .Z(n23000) );
  AND U31599 ( .A(n23001), .B(n23002), .Z(n22999) );
  NANDN U31600 ( .A(n23003), .B(n23004), .Z(n23002) );
  NANDN U31601 ( .A(n23005), .B(n23006), .Z(n23004) );
  NANDN U31602 ( .A(n23006), .B(n23005), .Z(n23001) );
  NAND U31603 ( .A(n23007), .B(n23008), .Z(n22996) );
  NANDN U31604 ( .A(n23009), .B(n23010), .Z(n23008) );
  OR U31605 ( .A(n23011), .B(n23012), .Z(n23010) );
  NAND U31606 ( .A(n23012), .B(n23011), .Z(n23007) );
  AND U31607 ( .A(n23013), .B(n23014), .Z(n22998) );
  NANDN U31608 ( .A(n23015), .B(n23016), .Z(n23014) );
  NANDN U31609 ( .A(n23017), .B(n23018), .Z(n23016) );
  NANDN U31610 ( .A(n23018), .B(n23017), .Z(n23013) );
  XOR U31611 ( .A(n23012), .B(n23019), .Z(N63350) );
  XOR U31612 ( .A(n23009), .B(n23011), .Z(n23019) );
  XNOR U31613 ( .A(n23005), .B(n23020), .Z(n23011) );
  XNOR U31614 ( .A(n23003), .B(n23006), .Z(n23020) );
  NAND U31615 ( .A(n23021), .B(n23022), .Z(n23006) );
  NAND U31616 ( .A(n23023), .B(n23024), .Z(n23022) );
  OR U31617 ( .A(n23025), .B(n23026), .Z(n23023) );
  NANDN U31618 ( .A(n23027), .B(n23025), .Z(n23021) );
  IV U31619 ( .A(n23026), .Z(n23027) );
  NAND U31620 ( .A(n23028), .B(n23029), .Z(n23003) );
  NAND U31621 ( .A(n23030), .B(n23031), .Z(n23029) );
  NANDN U31622 ( .A(n23032), .B(n23033), .Z(n23030) );
  NANDN U31623 ( .A(n23033), .B(n23032), .Z(n23028) );
  AND U31624 ( .A(n23034), .B(n23035), .Z(n23005) );
  NAND U31625 ( .A(n23036), .B(n23037), .Z(n23035) );
  OR U31626 ( .A(n23038), .B(n23039), .Z(n23036) );
  NANDN U31627 ( .A(n23040), .B(n23038), .Z(n23034) );
  NAND U31628 ( .A(n23041), .B(n23042), .Z(n23009) );
  NANDN U31629 ( .A(n23043), .B(n23044), .Z(n23042) );
  OR U31630 ( .A(n23045), .B(n23046), .Z(n23044) );
  NANDN U31631 ( .A(n23047), .B(n23045), .Z(n23041) );
  IV U31632 ( .A(n23046), .Z(n23047) );
  XNOR U31633 ( .A(n23017), .B(n23048), .Z(n23012) );
  XNOR U31634 ( .A(n23015), .B(n23018), .Z(n23048) );
  NAND U31635 ( .A(n23049), .B(n23050), .Z(n23018) );
  NAND U31636 ( .A(n23051), .B(n23052), .Z(n23050) );
  OR U31637 ( .A(n23053), .B(n23054), .Z(n23051) );
  NANDN U31638 ( .A(n23055), .B(n23053), .Z(n23049) );
  IV U31639 ( .A(n23054), .Z(n23055) );
  NAND U31640 ( .A(n23056), .B(n23057), .Z(n23015) );
  NAND U31641 ( .A(n23058), .B(n23059), .Z(n23057) );
  NANDN U31642 ( .A(n23060), .B(n23061), .Z(n23058) );
  NANDN U31643 ( .A(n23061), .B(n23060), .Z(n23056) );
  AND U31644 ( .A(n23062), .B(n23063), .Z(n23017) );
  NAND U31645 ( .A(n23064), .B(n23065), .Z(n23063) );
  OR U31646 ( .A(n23066), .B(n23067), .Z(n23064) );
  NANDN U31647 ( .A(n23068), .B(n23066), .Z(n23062) );
  XNOR U31648 ( .A(n23043), .B(n23069), .Z(N63349) );
  XOR U31649 ( .A(n23045), .B(n23046), .Z(n23069) );
  XNOR U31650 ( .A(n23059), .B(n23070), .Z(n23046) );
  XOR U31651 ( .A(n23060), .B(n23061), .Z(n23070) );
  XOR U31652 ( .A(n23066), .B(n23071), .Z(n23061) );
  XOR U31653 ( .A(n23065), .B(n23068), .Z(n23071) );
  IV U31654 ( .A(n23067), .Z(n23068) );
  NAND U31655 ( .A(n23072), .B(n23073), .Z(n23067) );
  OR U31656 ( .A(n23074), .B(n23075), .Z(n23073) );
  OR U31657 ( .A(n23076), .B(n23077), .Z(n23072) );
  NAND U31658 ( .A(n23078), .B(n23079), .Z(n23065) );
  OR U31659 ( .A(n23080), .B(n23081), .Z(n23079) );
  OR U31660 ( .A(n23082), .B(n23083), .Z(n23078) );
  NOR U31661 ( .A(n23084), .B(n23085), .Z(n23066) );
  ANDN U31662 ( .B(n23086), .A(n23087), .Z(n23060) );
  XNOR U31663 ( .A(n23053), .B(n23088), .Z(n23059) );
  XNOR U31664 ( .A(n23052), .B(n23054), .Z(n23088) );
  NAND U31665 ( .A(n23089), .B(n23090), .Z(n23054) );
  OR U31666 ( .A(n23091), .B(n23092), .Z(n23090) );
  OR U31667 ( .A(n23093), .B(n23094), .Z(n23089) );
  NAND U31668 ( .A(n23095), .B(n23096), .Z(n23052) );
  OR U31669 ( .A(n23097), .B(n23098), .Z(n23096) );
  OR U31670 ( .A(n23099), .B(n23100), .Z(n23095) );
  ANDN U31671 ( .B(n23101), .A(n23102), .Z(n23053) );
  IV U31672 ( .A(n23103), .Z(n23101) );
  ANDN U31673 ( .B(n23104), .A(n23105), .Z(n23045) );
  XOR U31674 ( .A(n23031), .B(n23106), .Z(n23043) );
  XOR U31675 ( .A(n23032), .B(n23033), .Z(n23106) );
  XOR U31676 ( .A(n23038), .B(n23107), .Z(n23033) );
  XOR U31677 ( .A(n23037), .B(n23040), .Z(n23107) );
  IV U31678 ( .A(n23039), .Z(n23040) );
  NAND U31679 ( .A(n23108), .B(n23109), .Z(n23039) );
  OR U31680 ( .A(n23110), .B(n23111), .Z(n23109) );
  OR U31681 ( .A(n23112), .B(n23113), .Z(n23108) );
  NAND U31682 ( .A(n23114), .B(n23115), .Z(n23037) );
  OR U31683 ( .A(n23116), .B(n23117), .Z(n23115) );
  OR U31684 ( .A(n23118), .B(n23119), .Z(n23114) );
  NOR U31685 ( .A(n23120), .B(n23121), .Z(n23038) );
  ANDN U31686 ( .B(n23122), .A(n23123), .Z(n23032) );
  IV U31687 ( .A(n23124), .Z(n23122) );
  XNOR U31688 ( .A(n23025), .B(n23125), .Z(n23031) );
  XNOR U31689 ( .A(n23024), .B(n23026), .Z(n23125) );
  NAND U31690 ( .A(n23126), .B(n23127), .Z(n23026) );
  OR U31691 ( .A(n23128), .B(n23129), .Z(n23127) );
  OR U31692 ( .A(n23130), .B(n23131), .Z(n23126) );
  NAND U31693 ( .A(n23132), .B(n23133), .Z(n23024) );
  OR U31694 ( .A(n23134), .B(n23135), .Z(n23133) );
  OR U31695 ( .A(n23136), .B(n23137), .Z(n23132) );
  ANDN U31696 ( .B(n23138), .A(n23139), .Z(n23025) );
  IV U31697 ( .A(n23140), .Z(n23138) );
  XNOR U31698 ( .A(n23105), .B(n23104), .Z(N63348) );
  XOR U31699 ( .A(n23124), .B(n23123), .Z(n23104) );
  XNOR U31700 ( .A(n23139), .B(n23140), .Z(n23123) );
  XNOR U31701 ( .A(n23134), .B(n23135), .Z(n23140) );
  XNOR U31702 ( .A(n23136), .B(n23137), .Z(n23135) );
  XNOR U31703 ( .A(y[5101]), .B(x[5101]), .Z(n23137) );
  XNOR U31704 ( .A(y[5102]), .B(x[5102]), .Z(n23136) );
  XNOR U31705 ( .A(y[5100]), .B(x[5100]), .Z(n23134) );
  XNOR U31706 ( .A(n23128), .B(n23129), .Z(n23139) );
  XNOR U31707 ( .A(y[5097]), .B(x[5097]), .Z(n23129) );
  XNOR U31708 ( .A(n23130), .B(n23131), .Z(n23128) );
  XNOR U31709 ( .A(y[5098]), .B(x[5098]), .Z(n23131) );
  XNOR U31710 ( .A(y[5099]), .B(x[5099]), .Z(n23130) );
  XNOR U31711 ( .A(n23121), .B(n23120), .Z(n23124) );
  XNOR U31712 ( .A(n23116), .B(n23117), .Z(n23120) );
  XNOR U31713 ( .A(y[5094]), .B(x[5094]), .Z(n23117) );
  XNOR U31714 ( .A(n23118), .B(n23119), .Z(n23116) );
  XNOR U31715 ( .A(y[5095]), .B(x[5095]), .Z(n23119) );
  XNOR U31716 ( .A(y[5096]), .B(x[5096]), .Z(n23118) );
  XNOR U31717 ( .A(n23110), .B(n23111), .Z(n23121) );
  XNOR U31718 ( .A(y[5091]), .B(x[5091]), .Z(n23111) );
  XNOR U31719 ( .A(n23112), .B(n23113), .Z(n23110) );
  XNOR U31720 ( .A(y[5092]), .B(x[5092]), .Z(n23113) );
  XNOR U31721 ( .A(y[5093]), .B(x[5093]), .Z(n23112) );
  XOR U31722 ( .A(n23086), .B(n23087), .Z(n23105) );
  XNOR U31723 ( .A(n23102), .B(n23103), .Z(n23087) );
  XNOR U31724 ( .A(n23097), .B(n23098), .Z(n23103) );
  XNOR U31725 ( .A(n23099), .B(n23100), .Z(n23098) );
  XNOR U31726 ( .A(y[5089]), .B(x[5089]), .Z(n23100) );
  XNOR U31727 ( .A(y[5090]), .B(x[5090]), .Z(n23099) );
  XNOR U31728 ( .A(y[5088]), .B(x[5088]), .Z(n23097) );
  XNOR U31729 ( .A(n23091), .B(n23092), .Z(n23102) );
  XNOR U31730 ( .A(y[5085]), .B(x[5085]), .Z(n23092) );
  XNOR U31731 ( .A(n23093), .B(n23094), .Z(n23091) );
  XNOR U31732 ( .A(y[5086]), .B(x[5086]), .Z(n23094) );
  XNOR U31733 ( .A(y[5087]), .B(x[5087]), .Z(n23093) );
  XOR U31734 ( .A(n23085), .B(n23084), .Z(n23086) );
  XNOR U31735 ( .A(n23080), .B(n23081), .Z(n23084) );
  XNOR U31736 ( .A(y[5082]), .B(x[5082]), .Z(n23081) );
  XNOR U31737 ( .A(n23082), .B(n23083), .Z(n23080) );
  XNOR U31738 ( .A(y[5083]), .B(x[5083]), .Z(n23083) );
  XNOR U31739 ( .A(y[5084]), .B(x[5084]), .Z(n23082) );
  XNOR U31740 ( .A(n23074), .B(n23075), .Z(n23085) );
  XNOR U31741 ( .A(y[5079]), .B(x[5079]), .Z(n23075) );
  XNOR U31742 ( .A(n23076), .B(n23077), .Z(n23074) );
  XNOR U31743 ( .A(y[5080]), .B(x[5080]), .Z(n23077) );
  XNOR U31744 ( .A(y[5081]), .B(x[5081]), .Z(n23076) );
  NAND U31745 ( .A(n23141), .B(n23142), .Z(N63339) );
  NANDN U31746 ( .A(n23143), .B(n23144), .Z(n23142) );
  OR U31747 ( .A(n23145), .B(n23146), .Z(n23144) );
  NAND U31748 ( .A(n23145), .B(n23146), .Z(n23141) );
  XOR U31749 ( .A(n23145), .B(n23147), .Z(N63338) );
  XNOR U31750 ( .A(n23143), .B(n23146), .Z(n23147) );
  AND U31751 ( .A(n23148), .B(n23149), .Z(n23146) );
  NANDN U31752 ( .A(n23150), .B(n23151), .Z(n23149) );
  NANDN U31753 ( .A(n23152), .B(n23153), .Z(n23151) );
  NANDN U31754 ( .A(n23153), .B(n23152), .Z(n23148) );
  NAND U31755 ( .A(n23154), .B(n23155), .Z(n23143) );
  NANDN U31756 ( .A(n23156), .B(n23157), .Z(n23155) );
  OR U31757 ( .A(n23158), .B(n23159), .Z(n23157) );
  NAND U31758 ( .A(n23159), .B(n23158), .Z(n23154) );
  AND U31759 ( .A(n23160), .B(n23161), .Z(n23145) );
  NANDN U31760 ( .A(n23162), .B(n23163), .Z(n23161) );
  NANDN U31761 ( .A(n23164), .B(n23165), .Z(n23163) );
  NANDN U31762 ( .A(n23165), .B(n23164), .Z(n23160) );
  XOR U31763 ( .A(n23159), .B(n23166), .Z(N63337) );
  XOR U31764 ( .A(n23156), .B(n23158), .Z(n23166) );
  XNOR U31765 ( .A(n23152), .B(n23167), .Z(n23158) );
  XNOR U31766 ( .A(n23150), .B(n23153), .Z(n23167) );
  NAND U31767 ( .A(n23168), .B(n23169), .Z(n23153) );
  NAND U31768 ( .A(n23170), .B(n23171), .Z(n23169) );
  OR U31769 ( .A(n23172), .B(n23173), .Z(n23170) );
  NANDN U31770 ( .A(n23174), .B(n23172), .Z(n23168) );
  IV U31771 ( .A(n23173), .Z(n23174) );
  NAND U31772 ( .A(n23175), .B(n23176), .Z(n23150) );
  NAND U31773 ( .A(n23177), .B(n23178), .Z(n23176) );
  NANDN U31774 ( .A(n23179), .B(n23180), .Z(n23177) );
  NANDN U31775 ( .A(n23180), .B(n23179), .Z(n23175) );
  AND U31776 ( .A(n23181), .B(n23182), .Z(n23152) );
  NAND U31777 ( .A(n23183), .B(n23184), .Z(n23182) );
  OR U31778 ( .A(n23185), .B(n23186), .Z(n23183) );
  NANDN U31779 ( .A(n23187), .B(n23185), .Z(n23181) );
  NAND U31780 ( .A(n23188), .B(n23189), .Z(n23156) );
  NANDN U31781 ( .A(n23190), .B(n23191), .Z(n23189) );
  OR U31782 ( .A(n23192), .B(n23193), .Z(n23191) );
  NANDN U31783 ( .A(n23194), .B(n23192), .Z(n23188) );
  IV U31784 ( .A(n23193), .Z(n23194) );
  XNOR U31785 ( .A(n23164), .B(n23195), .Z(n23159) );
  XNOR U31786 ( .A(n23162), .B(n23165), .Z(n23195) );
  NAND U31787 ( .A(n23196), .B(n23197), .Z(n23165) );
  NAND U31788 ( .A(n23198), .B(n23199), .Z(n23197) );
  OR U31789 ( .A(n23200), .B(n23201), .Z(n23198) );
  NANDN U31790 ( .A(n23202), .B(n23200), .Z(n23196) );
  IV U31791 ( .A(n23201), .Z(n23202) );
  NAND U31792 ( .A(n23203), .B(n23204), .Z(n23162) );
  NAND U31793 ( .A(n23205), .B(n23206), .Z(n23204) );
  NANDN U31794 ( .A(n23207), .B(n23208), .Z(n23205) );
  NANDN U31795 ( .A(n23208), .B(n23207), .Z(n23203) );
  AND U31796 ( .A(n23209), .B(n23210), .Z(n23164) );
  NAND U31797 ( .A(n23211), .B(n23212), .Z(n23210) );
  OR U31798 ( .A(n23213), .B(n23214), .Z(n23211) );
  NANDN U31799 ( .A(n23215), .B(n23213), .Z(n23209) );
  XNOR U31800 ( .A(n23190), .B(n23216), .Z(N63336) );
  XOR U31801 ( .A(n23192), .B(n23193), .Z(n23216) );
  XNOR U31802 ( .A(n23206), .B(n23217), .Z(n23193) );
  XOR U31803 ( .A(n23207), .B(n23208), .Z(n23217) );
  XOR U31804 ( .A(n23213), .B(n23218), .Z(n23208) );
  XOR U31805 ( .A(n23212), .B(n23215), .Z(n23218) );
  IV U31806 ( .A(n23214), .Z(n23215) );
  NAND U31807 ( .A(n23219), .B(n23220), .Z(n23214) );
  OR U31808 ( .A(n23221), .B(n23222), .Z(n23220) );
  OR U31809 ( .A(n23223), .B(n23224), .Z(n23219) );
  NAND U31810 ( .A(n23225), .B(n23226), .Z(n23212) );
  OR U31811 ( .A(n23227), .B(n23228), .Z(n23226) );
  OR U31812 ( .A(n23229), .B(n23230), .Z(n23225) );
  NOR U31813 ( .A(n23231), .B(n23232), .Z(n23213) );
  ANDN U31814 ( .B(n23233), .A(n23234), .Z(n23207) );
  XNOR U31815 ( .A(n23200), .B(n23235), .Z(n23206) );
  XNOR U31816 ( .A(n23199), .B(n23201), .Z(n23235) );
  NAND U31817 ( .A(n23236), .B(n23237), .Z(n23201) );
  OR U31818 ( .A(n23238), .B(n23239), .Z(n23237) );
  OR U31819 ( .A(n23240), .B(n23241), .Z(n23236) );
  NAND U31820 ( .A(n23242), .B(n23243), .Z(n23199) );
  OR U31821 ( .A(n23244), .B(n23245), .Z(n23243) );
  OR U31822 ( .A(n23246), .B(n23247), .Z(n23242) );
  ANDN U31823 ( .B(n23248), .A(n23249), .Z(n23200) );
  IV U31824 ( .A(n23250), .Z(n23248) );
  ANDN U31825 ( .B(n23251), .A(n23252), .Z(n23192) );
  XOR U31826 ( .A(n23178), .B(n23253), .Z(n23190) );
  XOR U31827 ( .A(n23179), .B(n23180), .Z(n23253) );
  XOR U31828 ( .A(n23185), .B(n23254), .Z(n23180) );
  XOR U31829 ( .A(n23184), .B(n23187), .Z(n23254) );
  IV U31830 ( .A(n23186), .Z(n23187) );
  NAND U31831 ( .A(n23255), .B(n23256), .Z(n23186) );
  OR U31832 ( .A(n23257), .B(n23258), .Z(n23256) );
  OR U31833 ( .A(n23259), .B(n23260), .Z(n23255) );
  NAND U31834 ( .A(n23261), .B(n23262), .Z(n23184) );
  OR U31835 ( .A(n23263), .B(n23264), .Z(n23262) );
  OR U31836 ( .A(n23265), .B(n23266), .Z(n23261) );
  NOR U31837 ( .A(n23267), .B(n23268), .Z(n23185) );
  ANDN U31838 ( .B(n23269), .A(n23270), .Z(n23179) );
  IV U31839 ( .A(n23271), .Z(n23269) );
  XNOR U31840 ( .A(n23172), .B(n23272), .Z(n23178) );
  XNOR U31841 ( .A(n23171), .B(n23173), .Z(n23272) );
  NAND U31842 ( .A(n23273), .B(n23274), .Z(n23173) );
  OR U31843 ( .A(n23275), .B(n23276), .Z(n23274) );
  OR U31844 ( .A(n23277), .B(n23278), .Z(n23273) );
  NAND U31845 ( .A(n23279), .B(n23280), .Z(n23171) );
  OR U31846 ( .A(n23281), .B(n23282), .Z(n23280) );
  OR U31847 ( .A(n23283), .B(n23284), .Z(n23279) );
  ANDN U31848 ( .B(n23285), .A(n23286), .Z(n23172) );
  IV U31849 ( .A(n23287), .Z(n23285) );
  XNOR U31850 ( .A(n23252), .B(n23251), .Z(N63335) );
  XOR U31851 ( .A(n23271), .B(n23270), .Z(n23251) );
  XNOR U31852 ( .A(n23286), .B(n23287), .Z(n23270) );
  XNOR U31853 ( .A(n23281), .B(n23282), .Z(n23287) );
  XNOR U31854 ( .A(n23283), .B(n23284), .Z(n23282) );
  XNOR U31855 ( .A(y[5077]), .B(x[5077]), .Z(n23284) );
  XNOR U31856 ( .A(y[5078]), .B(x[5078]), .Z(n23283) );
  XNOR U31857 ( .A(y[5076]), .B(x[5076]), .Z(n23281) );
  XNOR U31858 ( .A(n23275), .B(n23276), .Z(n23286) );
  XNOR U31859 ( .A(y[5073]), .B(x[5073]), .Z(n23276) );
  XNOR U31860 ( .A(n23277), .B(n23278), .Z(n23275) );
  XNOR U31861 ( .A(y[5074]), .B(x[5074]), .Z(n23278) );
  XNOR U31862 ( .A(y[5075]), .B(x[5075]), .Z(n23277) );
  XNOR U31863 ( .A(n23268), .B(n23267), .Z(n23271) );
  XNOR U31864 ( .A(n23263), .B(n23264), .Z(n23267) );
  XNOR U31865 ( .A(y[5070]), .B(x[5070]), .Z(n23264) );
  XNOR U31866 ( .A(n23265), .B(n23266), .Z(n23263) );
  XNOR U31867 ( .A(y[5071]), .B(x[5071]), .Z(n23266) );
  XNOR U31868 ( .A(y[5072]), .B(x[5072]), .Z(n23265) );
  XNOR U31869 ( .A(n23257), .B(n23258), .Z(n23268) );
  XNOR U31870 ( .A(y[5067]), .B(x[5067]), .Z(n23258) );
  XNOR U31871 ( .A(n23259), .B(n23260), .Z(n23257) );
  XNOR U31872 ( .A(y[5068]), .B(x[5068]), .Z(n23260) );
  XNOR U31873 ( .A(y[5069]), .B(x[5069]), .Z(n23259) );
  XOR U31874 ( .A(n23233), .B(n23234), .Z(n23252) );
  XNOR U31875 ( .A(n23249), .B(n23250), .Z(n23234) );
  XNOR U31876 ( .A(n23244), .B(n23245), .Z(n23250) );
  XNOR U31877 ( .A(n23246), .B(n23247), .Z(n23245) );
  XNOR U31878 ( .A(y[5065]), .B(x[5065]), .Z(n23247) );
  XNOR U31879 ( .A(y[5066]), .B(x[5066]), .Z(n23246) );
  XNOR U31880 ( .A(y[5064]), .B(x[5064]), .Z(n23244) );
  XNOR U31881 ( .A(n23238), .B(n23239), .Z(n23249) );
  XNOR U31882 ( .A(y[5061]), .B(x[5061]), .Z(n23239) );
  XNOR U31883 ( .A(n23240), .B(n23241), .Z(n23238) );
  XNOR U31884 ( .A(y[5062]), .B(x[5062]), .Z(n23241) );
  XNOR U31885 ( .A(y[5063]), .B(x[5063]), .Z(n23240) );
  XOR U31886 ( .A(n23232), .B(n23231), .Z(n23233) );
  XNOR U31887 ( .A(n23227), .B(n23228), .Z(n23231) );
  XNOR U31888 ( .A(y[5058]), .B(x[5058]), .Z(n23228) );
  XNOR U31889 ( .A(n23229), .B(n23230), .Z(n23227) );
  XNOR U31890 ( .A(y[5059]), .B(x[5059]), .Z(n23230) );
  XNOR U31891 ( .A(y[5060]), .B(x[5060]), .Z(n23229) );
  XNOR U31892 ( .A(n23221), .B(n23222), .Z(n23232) );
  XNOR U31893 ( .A(y[5055]), .B(x[5055]), .Z(n23222) );
  XNOR U31894 ( .A(n23223), .B(n23224), .Z(n23221) );
  XNOR U31895 ( .A(y[5056]), .B(x[5056]), .Z(n23224) );
  XNOR U31896 ( .A(y[5057]), .B(x[5057]), .Z(n23223) );
  NAND U31897 ( .A(n23288), .B(n23289), .Z(N63326) );
  NANDN U31898 ( .A(n23290), .B(n23291), .Z(n23289) );
  OR U31899 ( .A(n23292), .B(n23293), .Z(n23291) );
  NAND U31900 ( .A(n23292), .B(n23293), .Z(n23288) );
  XOR U31901 ( .A(n23292), .B(n23294), .Z(N63325) );
  XNOR U31902 ( .A(n23290), .B(n23293), .Z(n23294) );
  AND U31903 ( .A(n23295), .B(n23296), .Z(n23293) );
  NANDN U31904 ( .A(n23297), .B(n23298), .Z(n23296) );
  NANDN U31905 ( .A(n23299), .B(n23300), .Z(n23298) );
  NANDN U31906 ( .A(n23300), .B(n23299), .Z(n23295) );
  NAND U31907 ( .A(n23301), .B(n23302), .Z(n23290) );
  NANDN U31908 ( .A(n23303), .B(n23304), .Z(n23302) );
  OR U31909 ( .A(n23305), .B(n23306), .Z(n23304) );
  NAND U31910 ( .A(n23306), .B(n23305), .Z(n23301) );
  AND U31911 ( .A(n23307), .B(n23308), .Z(n23292) );
  NANDN U31912 ( .A(n23309), .B(n23310), .Z(n23308) );
  NANDN U31913 ( .A(n23311), .B(n23312), .Z(n23310) );
  NANDN U31914 ( .A(n23312), .B(n23311), .Z(n23307) );
  XOR U31915 ( .A(n23306), .B(n23313), .Z(N63324) );
  XOR U31916 ( .A(n23303), .B(n23305), .Z(n23313) );
  XNOR U31917 ( .A(n23299), .B(n23314), .Z(n23305) );
  XNOR U31918 ( .A(n23297), .B(n23300), .Z(n23314) );
  NAND U31919 ( .A(n23315), .B(n23316), .Z(n23300) );
  NAND U31920 ( .A(n23317), .B(n23318), .Z(n23316) );
  OR U31921 ( .A(n23319), .B(n23320), .Z(n23317) );
  NANDN U31922 ( .A(n23321), .B(n23319), .Z(n23315) );
  IV U31923 ( .A(n23320), .Z(n23321) );
  NAND U31924 ( .A(n23322), .B(n23323), .Z(n23297) );
  NAND U31925 ( .A(n23324), .B(n23325), .Z(n23323) );
  NANDN U31926 ( .A(n23326), .B(n23327), .Z(n23324) );
  NANDN U31927 ( .A(n23327), .B(n23326), .Z(n23322) );
  AND U31928 ( .A(n23328), .B(n23329), .Z(n23299) );
  NAND U31929 ( .A(n23330), .B(n23331), .Z(n23329) );
  OR U31930 ( .A(n23332), .B(n23333), .Z(n23330) );
  NANDN U31931 ( .A(n23334), .B(n23332), .Z(n23328) );
  NAND U31932 ( .A(n23335), .B(n23336), .Z(n23303) );
  NANDN U31933 ( .A(n23337), .B(n23338), .Z(n23336) );
  OR U31934 ( .A(n23339), .B(n23340), .Z(n23338) );
  NANDN U31935 ( .A(n23341), .B(n23339), .Z(n23335) );
  IV U31936 ( .A(n23340), .Z(n23341) );
  XNOR U31937 ( .A(n23311), .B(n23342), .Z(n23306) );
  XNOR U31938 ( .A(n23309), .B(n23312), .Z(n23342) );
  NAND U31939 ( .A(n23343), .B(n23344), .Z(n23312) );
  NAND U31940 ( .A(n23345), .B(n23346), .Z(n23344) );
  OR U31941 ( .A(n23347), .B(n23348), .Z(n23345) );
  NANDN U31942 ( .A(n23349), .B(n23347), .Z(n23343) );
  IV U31943 ( .A(n23348), .Z(n23349) );
  NAND U31944 ( .A(n23350), .B(n23351), .Z(n23309) );
  NAND U31945 ( .A(n23352), .B(n23353), .Z(n23351) );
  NANDN U31946 ( .A(n23354), .B(n23355), .Z(n23352) );
  NANDN U31947 ( .A(n23355), .B(n23354), .Z(n23350) );
  AND U31948 ( .A(n23356), .B(n23357), .Z(n23311) );
  NAND U31949 ( .A(n23358), .B(n23359), .Z(n23357) );
  OR U31950 ( .A(n23360), .B(n23361), .Z(n23358) );
  NANDN U31951 ( .A(n23362), .B(n23360), .Z(n23356) );
  XNOR U31952 ( .A(n23337), .B(n23363), .Z(N63323) );
  XOR U31953 ( .A(n23339), .B(n23340), .Z(n23363) );
  XNOR U31954 ( .A(n23353), .B(n23364), .Z(n23340) );
  XOR U31955 ( .A(n23354), .B(n23355), .Z(n23364) );
  XOR U31956 ( .A(n23360), .B(n23365), .Z(n23355) );
  XOR U31957 ( .A(n23359), .B(n23362), .Z(n23365) );
  IV U31958 ( .A(n23361), .Z(n23362) );
  NAND U31959 ( .A(n23366), .B(n23367), .Z(n23361) );
  OR U31960 ( .A(n23368), .B(n23369), .Z(n23367) );
  OR U31961 ( .A(n23370), .B(n23371), .Z(n23366) );
  NAND U31962 ( .A(n23372), .B(n23373), .Z(n23359) );
  OR U31963 ( .A(n23374), .B(n23375), .Z(n23373) );
  OR U31964 ( .A(n23376), .B(n23377), .Z(n23372) );
  NOR U31965 ( .A(n23378), .B(n23379), .Z(n23360) );
  ANDN U31966 ( .B(n23380), .A(n23381), .Z(n23354) );
  XNOR U31967 ( .A(n23347), .B(n23382), .Z(n23353) );
  XNOR U31968 ( .A(n23346), .B(n23348), .Z(n23382) );
  NAND U31969 ( .A(n23383), .B(n23384), .Z(n23348) );
  OR U31970 ( .A(n23385), .B(n23386), .Z(n23384) );
  OR U31971 ( .A(n23387), .B(n23388), .Z(n23383) );
  NAND U31972 ( .A(n23389), .B(n23390), .Z(n23346) );
  OR U31973 ( .A(n23391), .B(n23392), .Z(n23390) );
  OR U31974 ( .A(n23393), .B(n23394), .Z(n23389) );
  ANDN U31975 ( .B(n23395), .A(n23396), .Z(n23347) );
  IV U31976 ( .A(n23397), .Z(n23395) );
  ANDN U31977 ( .B(n23398), .A(n23399), .Z(n23339) );
  XOR U31978 ( .A(n23325), .B(n23400), .Z(n23337) );
  XOR U31979 ( .A(n23326), .B(n23327), .Z(n23400) );
  XOR U31980 ( .A(n23332), .B(n23401), .Z(n23327) );
  XOR U31981 ( .A(n23331), .B(n23334), .Z(n23401) );
  IV U31982 ( .A(n23333), .Z(n23334) );
  NAND U31983 ( .A(n23402), .B(n23403), .Z(n23333) );
  OR U31984 ( .A(n23404), .B(n23405), .Z(n23403) );
  OR U31985 ( .A(n23406), .B(n23407), .Z(n23402) );
  NAND U31986 ( .A(n23408), .B(n23409), .Z(n23331) );
  OR U31987 ( .A(n23410), .B(n23411), .Z(n23409) );
  OR U31988 ( .A(n23412), .B(n23413), .Z(n23408) );
  NOR U31989 ( .A(n23414), .B(n23415), .Z(n23332) );
  ANDN U31990 ( .B(n23416), .A(n23417), .Z(n23326) );
  IV U31991 ( .A(n23418), .Z(n23416) );
  XNOR U31992 ( .A(n23319), .B(n23419), .Z(n23325) );
  XNOR U31993 ( .A(n23318), .B(n23320), .Z(n23419) );
  NAND U31994 ( .A(n23420), .B(n23421), .Z(n23320) );
  OR U31995 ( .A(n23422), .B(n23423), .Z(n23421) );
  OR U31996 ( .A(n23424), .B(n23425), .Z(n23420) );
  NAND U31997 ( .A(n23426), .B(n23427), .Z(n23318) );
  OR U31998 ( .A(n23428), .B(n23429), .Z(n23427) );
  OR U31999 ( .A(n23430), .B(n23431), .Z(n23426) );
  ANDN U32000 ( .B(n23432), .A(n23433), .Z(n23319) );
  IV U32001 ( .A(n23434), .Z(n23432) );
  XNOR U32002 ( .A(n23399), .B(n23398), .Z(N63322) );
  XOR U32003 ( .A(n23418), .B(n23417), .Z(n23398) );
  XNOR U32004 ( .A(n23433), .B(n23434), .Z(n23417) );
  XNOR U32005 ( .A(n23428), .B(n23429), .Z(n23434) );
  XNOR U32006 ( .A(n23430), .B(n23431), .Z(n23429) );
  XNOR U32007 ( .A(y[5053]), .B(x[5053]), .Z(n23431) );
  XNOR U32008 ( .A(y[5054]), .B(x[5054]), .Z(n23430) );
  XNOR U32009 ( .A(y[5052]), .B(x[5052]), .Z(n23428) );
  XNOR U32010 ( .A(n23422), .B(n23423), .Z(n23433) );
  XNOR U32011 ( .A(y[5049]), .B(x[5049]), .Z(n23423) );
  XNOR U32012 ( .A(n23424), .B(n23425), .Z(n23422) );
  XNOR U32013 ( .A(y[5050]), .B(x[5050]), .Z(n23425) );
  XNOR U32014 ( .A(y[5051]), .B(x[5051]), .Z(n23424) );
  XNOR U32015 ( .A(n23415), .B(n23414), .Z(n23418) );
  XNOR U32016 ( .A(n23410), .B(n23411), .Z(n23414) );
  XNOR U32017 ( .A(y[5046]), .B(x[5046]), .Z(n23411) );
  XNOR U32018 ( .A(n23412), .B(n23413), .Z(n23410) );
  XNOR U32019 ( .A(y[5047]), .B(x[5047]), .Z(n23413) );
  XNOR U32020 ( .A(y[5048]), .B(x[5048]), .Z(n23412) );
  XNOR U32021 ( .A(n23404), .B(n23405), .Z(n23415) );
  XNOR U32022 ( .A(y[5043]), .B(x[5043]), .Z(n23405) );
  XNOR U32023 ( .A(n23406), .B(n23407), .Z(n23404) );
  XNOR U32024 ( .A(y[5044]), .B(x[5044]), .Z(n23407) );
  XNOR U32025 ( .A(y[5045]), .B(x[5045]), .Z(n23406) );
  XOR U32026 ( .A(n23380), .B(n23381), .Z(n23399) );
  XNOR U32027 ( .A(n23396), .B(n23397), .Z(n23381) );
  XNOR U32028 ( .A(n23391), .B(n23392), .Z(n23397) );
  XNOR U32029 ( .A(n23393), .B(n23394), .Z(n23392) );
  XNOR U32030 ( .A(y[5041]), .B(x[5041]), .Z(n23394) );
  XNOR U32031 ( .A(y[5042]), .B(x[5042]), .Z(n23393) );
  XNOR U32032 ( .A(y[5040]), .B(x[5040]), .Z(n23391) );
  XNOR U32033 ( .A(n23385), .B(n23386), .Z(n23396) );
  XNOR U32034 ( .A(y[5037]), .B(x[5037]), .Z(n23386) );
  XNOR U32035 ( .A(n23387), .B(n23388), .Z(n23385) );
  XNOR U32036 ( .A(y[5038]), .B(x[5038]), .Z(n23388) );
  XNOR U32037 ( .A(y[5039]), .B(x[5039]), .Z(n23387) );
  XOR U32038 ( .A(n23379), .B(n23378), .Z(n23380) );
  XNOR U32039 ( .A(n23374), .B(n23375), .Z(n23378) );
  XNOR U32040 ( .A(y[5034]), .B(x[5034]), .Z(n23375) );
  XNOR U32041 ( .A(n23376), .B(n23377), .Z(n23374) );
  XNOR U32042 ( .A(y[5035]), .B(x[5035]), .Z(n23377) );
  XNOR U32043 ( .A(y[5036]), .B(x[5036]), .Z(n23376) );
  XNOR U32044 ( .A(n23368), .B(n23369), .Z(n23379) );
  XNOR U32045 ( .A(y[5031]), .B(x[5031]), .Z(n23369) );
  XNOR U32046 ( .A(n23370), .B(n23371), .Z(n23368) );
  XNOR U32047 ( .A(y[5032]), .B(x[5032]), .Z(n23371) );
  XNOR U32048 ( .A(y[5033]), .B(x[5033]), .Z(n23370) );
  NAND U32049 ( .A(n23435), .B(n23436), .Z(N63313) );
  NANDN U32050 ( .A(n23437), .B(n23438), .Z(n23436) );
  OR U32051 ( .A(n23439), .B(n23440), .Z(n23438) );
  NAND U32052 ( .A(n23439), .B(n23440), .Z(n23435) );
  XOR U32053 ( .A(n23439), .B(n23441), .Z(N63312) );
  XNOR U32054 ( .A(n23437), .B(n23440), .Z(n23441) );
  AND U32055 ( .A(n23442), .B(n23443), .Z(n23440) );
  NANDN U32056 ( .A(n23444), .B(n23445), .Z(n23443) );
  NANDN U32057 ( .A(n23446), .B(n23447), .Z(n23445) );
  NANDN U32058 ( .A(n23447), .B(n23446), .Z(n23442) );
  NAND U32059 ( .A(n23448), .B(n23449), .Z(n23437) );
  NANDN U32060 ( .A(n23450), .B(n23451), .Z(n23449) );
  OR U32061 ( .A(n23452), .B(n23453), .Z(n23451) );
  NAND U32062 ( .A(n23453), .B(n23452), .Z(n23448) );
  AND U32063 ( .A(n23454), .B(n23455), .Z(n23439) );
  NANDN U32064 ( .A(n23456), .B(n23457), .Z(n23455) );
  NANDN U32065 ( .A(n23458), .B(n23459), .Z(n23457) );
  NANDN U32066 ( .A(n23459), .B(n23458), .Z(n23454) );
  XOR U32067 ( .A(n23453), .B(n23460), .Z(N63311) );
  XOR U32068 ( .A(n23450), .B(n23452), .Z(n23460) );
  XNOR U32069 ( .A(n23446), .B(n23461), .Z(n23452) );
  XNOR U32070 ( .A(n23444), .B(n23447), .Z(n23461) );
  NAND U32071 ( .A(n23462), .B(n23463), .Z(n23447) );
  NAND U32072 ( .A(n23464), .B(n23465), .Z(n23463) );
  OR U32073 ( .A(n23466), .B(n23467), .Z(n23464) );
  NANDN U32074 ( .A(n23468), .B(n23466), .Z(n23462) );
  IV U32075 ( .A(n23467), .Z(n23468) );
  NAND U32076 ( .A(n23469), .B(n23470), .Z(n23444) );
  NAND U32077 ( .A(n23471), .B(n23472), .Z(n23470) );
  NANDN U32078 ( .A(n23473), .B(n23474), .Z(n23471) );
  NANDN U32079 ( .A(n23474), .B(n23473), .Z(n23469) );
  AND U32080 ( .A(n23475), .B(n23476), .Z(n23446) );
  NAND U32081 ( .A(n23477), .B(n23478), .Z(n23476) );
  OR U32082 ( .A(n23479), .B(n23480), .Z(n23477) );
  NANDN U32083 ( .A(n23481), .B(n23479), .Z(n23475) );
  NAND U32084 ( .A(n23482), .B(n23483), .Z(n23450) );
  NANDN U32085 ( .A(n23484), .B(n23485), .Z(n23483) );
  OR U32086 ( .A(n23486), .B(n23487), .Z(n23485) );
  NANDN U32087 ( .A(n23488), .B(n23486), .Z(n23482) );
  IV U32088 ( .A(n23487), .Z(n23488) );
  XNOR U32089 ( .A(n23458), .B(n23489), .Z(n23453) );
  XNOR U32090 ( .A(n23456), .B(n23459), .Z(n23489) );
  NAND U32091 ( .A(n23490), .B(n23491), .Z(n23459) );
  NAND U32092 ( .A(n23492), .B(n23493), .Z(n23491) );
  OR U32093 ( .A(n23494), .B(n23495), .Z(n23492) );
  NANDN U32094 ( .A(n23496), .B(n23494), .Z(n23490) );
  IV U32095 ( .A(n23495), .Z(n23496) );
  NAND U32096 ( .A(n23497), .B(n23498), .Z(n23456) );
  NAND U32097 ( .A(n23499), .B(n23500), .Z(n23498) );
  NANDN U32098 ( .A(n23501), .B(n23502), .Z(n23499) );
  NANDN U32099 ( .A(n23502), .B(n23501), .Z(n23497) );
  AND U32100 ( .A(n23503), .B(n23504), .Z(n23458) );
  NAND U32101 ( .A(n23505), .B(n23506), .Z(n23504) );
  OR U32102 ( .A(n23507), .B(n23508), .Z(n23505) );
  NANDN U32103 ( .A(n23509), .B(n23507), .Z(n23503) );
  XNOR U32104 ( .A(n23484), .B(n23510), .Z(N63310) );
  XOR U32105 ( .A(n23486), .B(n23487), .Z(n23510) );
  XNOR U32106 ( .A(n23500), .B(n23511), .Z(n23487) );
  XOR U32107 ( .A(n23501), .B(n23502), .Z(n23511) );
  XOR U32108 ( .A(n23507), .B(n23512), .Z(n23502) );
  XOR U32109 ( .A(n23506), .B(n23509), .Z(n23512) );
  IV U32110 ( .A(n23508), .Z(n23509) );
  NAND U32111 ( .A(n23513), .B(n23514), .Z(n23508) );
  OR U32112 ( .A(n23515), .B(n23516), .Z(n23514) );
  OR U32113 ( .A(n23517), .B(n23518), .Z(n23513) );
  NAND U32114 ( .A(n23519), .B(n23520), .Z(n23506) );
  OR U32115 ( .A(n23521), .B(n23522), .Z(n23520) );
  OR U32116 ( .A(n23523), .B(n23524), .Z(n23519) );
  NOR U32117 ( .A(n23525), .B(n23526), .Z(n23507) );
  ANDN U32118 ( .B(n23527), .A(n23528), .Z(n23501) );
  XNOR U32119 ( .A(n23494), .B(n23529), .Z(n23500) );
  XNOR U32120 ( .A(n23493), .B(n23495), .Z(n23529) );
  NAND U32121 ( .A(n23530), .B(n23531), .Z(n23495) );
  OR U32122 ( .A(n23532), .B(n23533), .Z(n23531) );
  OR U32123 ( .A(n23534), .B(n23535), .Z(n23530) );
  NAND U32124 ( .A(n23536), .B(n23537), .Z(n23493) );
  OR U32125 ( .A(n23538), .B(n23539), .Z(n23537) );
  OR U32126 ( .A(n23540), .B(n23541), .Z(n23536) );
  ANDN U32127 ( .B(n23542), .A(n23543), .Z(n23494) );
  IV U32128 ( .A(n23544), .Z(n23542) );
  ANDN U32129 ( .B(n23545), .A(n23546), .Z(n23486) );
  XOR U32130 ( .A(n23472), .B(n23547), .Z(n23484) );
  XOR U32131 ( .A(n23473), .B(n23474), .Z(n23547) );
  XOR U32132 ( .A(n23479), .B(n23548), .Z(n23474) );
  XOR U32133 ( .A(n23478), .B(n23481), .Z(n23548) );
  IV U32134 ( .A(n23480), .Z(n23481) );
  NAND U32135 ( .A(n23549), .B(n23550), .Z(n23480) );
  OR U32136 ( .A(n23551), .B(n23552), .Z(n23550) );
  OR U32137 ( .A(n23553), .B(n23554), .Z(n23549) );
  NAND U32138 ( .A(n23555), .B(n23556), .Z(n23478) );
  OR U32139 ( .A(n23557), .B(n23558), .Z(n23556) );
  OR U32140 ( .A(n23559), .B(n23560), .Z(n23555) );
  NOR U32141 ( .A(n23561), .B(n23562), .Z(n23479) );
  ANDN U32142 ( .B(n23563), .A(n23564), .Z(n23473) );
  IV U32143 ( .A(n23565), .Z(n23563) );
  XNOR U32144 ( .A(n23466), .B(n23566), .Z(n23472) );
  XNOR U32145 ( .A(n23465), .B(n23467), .Z(n23566) );
  NAND U32146 ( .A(n23567), .B(n23568), .Z(n23467) );
  OR U32147 ( .A(n23569), .B(n23570), .Z(n23568) );
  OR U32148 ( .A(n23571), .B(n23572), .Z(n23567) );
  NAND U32149 ( .A(n23573), .B(n23574), .Z(n23465) );
  OR U32150 ( .A(n23575), .B(n23576), .Z(n23574) );
  OR U32151 ( .A(n23577), .B(n23578), .Z(n23573) );
  ANDN U32152 ( .B(n23579), .A(n23580), .Z(n23466) );
  IV U32153 ( .A(n23581), .Z(n23579) );
  XNOR U32154 ( .A(n23546), .B(n23545), .Z(N63309) );
  XOR U32155 ( .A(n23565), .B(n23564), .Z(n23545) );
  XNOR U32156 ( .A(n23580), .B(n23581), .Z(n23564) );
  XNOR U32157 ( .A(n23575), .B(n23576), .Z(n23581) );
  XNOR U32158 ( .A(n23577), .B(n23578), .Z(n23576) );
  XNOR U32159 ( .A(y[5029]), .B(x[5029]), .Z(n23578) );
  XNOR U32160 ( .A(y[5030]), .B(x[5030]), .Z(n23577) );
  XNOR U32161 ( .A(y[5028]), .B(x[5028]), .Z(n23575) );
  XNOR U32162 ( .A(n23569), .B(n23570), .Z(n23580) );
  XNOR U32163 ( .A(y[5025]), .B(x[5025]), .Z(n23570) );
  XNOR U32164 ( .A(n23571), .B(n23572), .Z(n23569) );
  XNOR U32165 ( .A(y[5026]), .B(x[5026]), .Z(n23572) );
  XNOR U32166 ( .A(y[5027]), .B(x[5027]), .Z(n23571) );
  XNOR U32167 ( .A(n23562), .B(n23561), .Z(n23565) );
  XNOR U32168 ( .A(n23557), .B(n23558), .Z(n23561) );
  XNOR U32169 ( .A(y[5022]), .B(x[5022]), .Z(n23558) );
  XNOR U32170 ( .A(n23559), .B(n23560), .Z(n23557) );
  XNOR U32171 ( .A(y[5023]), .B(x[5023]), .Z(n23560) );
  XNOR U32172 ( .A(y[5024]), .B(x[5024]), .Z(n23559) );
  XNOR U32173 ( .A(n23551), .B(n23552), .Z(n23562) );
  XNOR U32174 ( .A(y[5019]), .B(x[5019]), .Z(n23552) );
  XNOR U32175 ( .A(n23553), .B(n23554), .Z(n23551) );
  XNOR U32176 ( .A(y[5020]), .B(x[5020]), .Z(n23554) );
  XNOR U32177 ( .A(y[5021]), .B(x[5021]), .Z(n23553) );
  XOR U32178 ( .A(n23527), .B(n23528), .Z(n23546) );
  XNOR U32179 ( .A(n23543), .B(n23544), .Z(n23528) );
  XNOR U32180 ( .A(n23538), .B(n23539), .Z(n23544) );
  XNOR U32181 ( .A(n23540), .B(n23541), .Z(n23539) );
  XNOR U32182 ( .A(y[5017]), .B(x[5017]), .Z(n23541) );
  XNOR U32183 ( .A(y[5018]), .B(x[5018]), .Z(n23540) );
  XNOR U32184 ( .A(y[5016]), .B(x[5016]), .Z(n23538) );
  XNOR U32185 ( .A(n23532), .B(n23533), .Z(n23543) );
  XNOR U32186 ( .A(y[5013]), .B(x[5013]), .Z(n23533) );
  XNOR U32187 ( .A(n23534), .B(n23535), .Z(n23532) );
  XNOR U32188 ( .A(y[5014]), .B(x[5014]), .Z(n23535) );
  XNOR U32189 ( .A(y[5015]), .B(x[5015]), .Z(n23534) );
  XOR U32190 ( .A(n23526), .B(n23525), .Z(n23527) );
  XNOR U32191 ( .A(n23521), .B(n23522), .Z(n23525) );
  XNOR U32192 ( .A(y[5010]), .B(x[5010]), .Z(n23522) );
  XNOR U32193 ( .A(n23523), .B(n23524), .Z(n23521) );
  XNOR U32194 ( .A(y[5011]), .B(x[5011]), .Z(n23524) );
  XNOR U32195 ( .A(y[5012]), .B(x[5012]), .Z(n23523) );
  XNOR U32196 ( .A(n23515), .B(n23516), .Z(n23526) );
  XNOR U32197 ( .A(y[5007]), .B(x[5007]), .Z(n23516) );
  XNOR U32198 ( .A(n23517), .B(n23518), .Z(n23515) );
  XNOR U32199 ( .A(y[5008]), .B(x[5008]), .Z(n23518) );
  XNOR U32200 ( .A(y[5009]), .B(x[5009]), .Z(n23517) );
  NAND U32201 ( .A(n23582), .B(n23583), .Z(N63300) );
  NANDN U32202 ( .A(n23584), .B(n23585), .Z(n23583) );
  OR U32203 ( .A(n23586), .B(n23587), .Z(n23585) );
  NAND U32204 ( .A(n23586), .B(n23587), .Z(n23582) );
  XOR U32205 ( .A(n23586), .B(n23588), .Z(N63299) );
  XNOR U32206 ( .A(n23584), .B(n23587), .Z(n23588) );
  AND U32207 ( .A(n23589), .B(n23590), .Z(n23587) );
  NANDN U32208 ( .A(n23591), .B(n23592), .Z(n23590) );
  NANDN U32209 ( .A(n23593), .B(n23594), .Z(n23592) );
  NANDN U32210 ( .A(n23594), .B(n23593), .Z(n23589) );
  NAND U32211 ( .A(n23595), .B(n23596), .Z(n23584) );
  NANDN U32212 ( .A(n23597), .B(n23598), .Z(n23596) );
  OR U32213 ( .A(n23599), .B(n23600), .Z(n23598) );
  NAND U32214 ( .A(n23600), .B(n23599), .Z(n23595) );
  AND U32215 ( .A(n23601), .B(n23602), .Z(n23586) );
  NANDN U32216 ( .A(n23603), .B(n23604), .Z(n23602) );
  NANDN U32217 ( .A(n23605), .B(n23606), .Z(n23604) );
  NANDN U32218 ( .A(n23606), .B(n23605), .Z(n23601) );
  XOR U32219 ( .A(n23600), .B(n23607), .Z(N63298) );
  XOR U32220 ( .A(n23597), .B(n23599), .Z(n23607) );
  XNOR U32221 ( .A(n23593), .B(n23608), .Z(n23599) );
  XNOR U32222 ( .A(n23591), .B(n23594), .Z(n23608) );
  NAND U32223 ( .A(n23609), .B(n23610), .Z(n23594) );
  NAND U32224 ( .A(n23611), .B(n23612), .Z(n23610) );
  OR U32225 ( .A(n23613), .B(n23614), .Z(n23611) );
  NANDN U32226 ( .A(n23615), .B(n23613), .Z(n23609) );
  IV U32227 ( .A(n23614), .Z(n23615) );
  NAND U32228 ( .A(n23616), .B(n23617), .Z(n23591) );
  NAND U32229 ( .A(n23618), .B(n23619), .Z(n23617) );
  NANDN U32230 ( .A(n23620), .B(n23621), .Z(n23618) );
  NANDN U32231 ( .A(n23621), .B(n23620), .Z(n23616) );
  AND U32232 ( .A(n23622), .B(n23623), .Z(n23593) );
  NAND U32233 ( .A(n23624), .B(n23625), .Z(n23623) );
  OR U32234 ( .A(n23626), .B(n23627), .Z(n23624) );
  NANDN U32235 ( .A(n23628), .B(n23626), .Z(n23622) );
  NAND U32236 ( .A(n23629), .B(n23630), .Z(n23597) );
  NANDN U32237 ( .A(n23631), .B(n23632), .Z(n23630) );
  OR U32238 ( .A(n23633), .B(n23634), .Z(n23632) );
  NANDN U32239 ( .A(n23635), .B(n23633), .Z(n23629) );
  IV U32240 ( .A(n23634), .Z(n23635) );
  XNOR U32241 ( .A(n23605), .B(n23636), .Z(n23600) );
  XNOR U32242 ( .A(n23603), .B(n23606), .Z(n23636) );
  NAND U32243 ( .A(n23637), .B(n23638), .Z(n23606) );
  NAND U32244 ( .A(n23639), .B(n23640), .Z(n23638) );
  OR U32245 ( .A(n23641), .B(n23642), .Z(n23639) );
  NANDN U32246 ( .A(n23643), .B(n23641), .Z(n23637) );
  IV U32247 ( .A(n23642), .Z(n23643) );
  NAND U32248 ( .A(n23644), .B(n23645), .Z(n23603) );
  NAND U32249 ( .A(n23646), .B(n23647), .Z(n23645) );
  NANDN U32250 ( .A(n23648), .B(n23649), .Z(n23646) );
  NANDN U32251 ( .A(n23649), .B(n23648), .Z(n23644) );
  AND U32252 ( .A(n23650), .B(n23651), .Z(n23605) );
  NAND U32253 ( .A(n23652), .B(n23653), .Z(n23651) );
  OR U32254 ( .A(n23654), .B(n23655), .Z(n23652) );
  NANDN U32255 ( .A(n23656), .B(n23654), .Z(n23650) );
  XNOR U32256 ( .A(n23631), .B(n23657), .Z(N63297) );
  XOR U32257 ( .A(n23633), .B(n23634), .Z(n23657) );
  XNOR U32258 ( .A(n23647), .B(n23658), .Z(n23634) );
  XOR U32259 ( .A(n23648), .B(n23649), .Z(n23658) );
  XOR U32260 ( .A(n23654), .B(n23659), .Z(n23649) );
  XOR U32261 ( .A(n23653), .B(n23656), .Z(n23659) );
  IV U32262 ( .A(n23655), .Z(n23656) );
  NAND U32263 ( .A(n23660), .B(n23661), .Z(n23655) );
  OR U32264 ( .A(n23662), .B(n23663), .Z(n23661) );
  OR U32265 ( .A(n23664), .B(n23665), .Z(n23660) );
  NAND U32266 ( .A(n23666), .B(n23667), .Z(n23653) );
  OR U32267 ( .A(n23668), .B(n23669), .Z(n23667) );
  OR U32268 ( .A(n23670), .B(n23671), .Z(n23666) );
  NOR U32269 ( .A(n23672), .B(n23673), .Z(n23654) );
  ANDN U32270 ( .B(n23674), .A(n23675), .Z(n23648) );
  XNOR U32271 ( .A(n23641), .B(n23676), .Z(n23647) );
  XNOR U32272 ( .A(n23640), .B(n23642), .Z(n23676) );
  NAND U32273 ( .A(n23677), .B(n23678), .Z(n23642) );
  OR U32274 ( .A(n23679), .B(n23680), .Z(n23678) );
  OR U32275 ( .A(n23681), .B(n23682), .Z(n23677) );
  NAND U32276 ( .A(n23683), .B(n23684), .Z(n23640) );
  OR U32277 ( .A(n23685), .B(n23686), .Z(n23684) );
  OR U32278 ( .A(n23687), .B(n23688), .Z(n23683) );
  ANDN U32279 ( .B(n23689), .A(n23690), .Z(n23641) );
  IV U32280 ( .A(n23691), .Z(n23689) );
  ANDN U32281 ( .B(n23692), .A(n23693), .Z(n23633) );
  XOR U32282 ( .A(n23619), .B(n23694), .Z(n23631) );
  XOR U32283 ( .A(n23620), .B(n23621), .Z(n23694) );
  XOR U32284 ( .A(n23626), .B(n23695), .Z(n23621) );
  XOR U32285 ( .A(n23625), .B(n23628), .Z(n23695) );
  IV U32286 ( .A(n23627), .Z(n23628) );
  NAND U32287 ( .A(n23696), .B(n23697), .Z(n23627) );
  OR U32288 ( .A(n23698), .B(n23699), .Z(n23697) );
  OR U32289 ( .A(n23700), .B(n23701), .Z(n23696) );
  NAND U32290 ( .A(n23702), .B(n23703), .Z(n23625) );
  OR U32291 ( .A(n23704), .B(n23705), .Z(n23703) );
  OR U32292 ( .A(n23706), .B(n23707), .Z(n23702) );
  NOR U32293 ( .A(n23708), .B(n23709), .Z(n23626) );
  ANDN U32294 ( .B(n23710), .A(n23711), .Z(n23620) );
  IV U32295 ( .A(n23712), .Z(n23710) );
  XNOR U32296 ( .A(n23613), .B(n23713), .Z(n23619) );
  XNOR U32297 ( .A(n23612), .B(n23614), .Z(n23713) );
  NAND U32298 ( .A(n23714), .B(n23715), .Z(n23614) );
  OR U32299 ( .A(n23716), .B(n23717), .Z(n23715) );
  OR U32300 ( .A(n23718), .B(n23719), .Z(n23714) );
  NAND U32301 ( .A(n23720), .B(n23721), .Z(n23612) );
  OR U32302 ( .A(n23722), .B(n23723), .Z(n23721) );
  OR U32303 ( .A(n23724), .B(n23725), .Z(n23720) );
  ANDN U32304 ( .B(n23726), .A(n23727), .Z(n23613) );
  IV U32305 ( .A(n23728), .Z(n23726) );
  XNOR U32306 ( .A(n23693), .B(n23692), .Z(N63296) );
  XOR U32307 ( .A(n23712), .B(n23711), .Z(n23692) );
  XNOR U32308 ( .A(n23727), .B(n23728), .Z(n23711) );
  XNOR U32309 ( .A(n23722), .B(n23723), .Z(n23728) );
  XNOR U32310 ( .A(n23724), .B(n23725), .Z(n23723) );
  XNOR U32311 ( .A(y[5005]), .B(x[5005]), .Z(n23725) );
  XNOR U32312 ( .A(y[5006]), .B(x[5006]), .Z(n23724) );
  XNOR U32313 ( .A(y[5004]), .B(x[5004]), .Z(n23722) );
  XNOR U32314 ( .A(n23716), .B(n23717), .Z(n23727) );
  XNOR U32315 ( .A(y[5001]), .B(x[5001]), .Z(n23717) );
  XNOR U32316 ( .A(n23718), .B(n23719), .Z(n23716) );
  XNOR U32317 ( .A(y[5002]), .B(x[5002]), .Z(n23719) );
  XNOR U32318 ( .A(y[5003]), .B(x[5003]), .Z(n23718) );
  XNOR U32319 ( .A(n23709), .B(n23708), .Z(n23712) );
  XNOR U32320 ( .A(n23704), .B(n23705), .Z(n23708) );
  XNOR U32321 ( .A(y[4998]), .B(x[4998]), .Z(n23705) );
  XNOR U32322 ( .A(n23706), .B(n23707), .Z(n23704) );
  XNOR U32323 ( .A(y[4999]), .B(x[4999]), .Z(n23707) );
  XNOR U32324 ( .A(y[5000]), .B(x[5000]), .Z(n23706) );
  XNOR U32325 ( .A(n23698), .B(n23699), .Z(n23709) );
  XNOR U32326 ( .A(y[4995]), .B(x[4995]), .Z(n23699) );
  XNOR U32327 ( .A(n23700), .B(n23701), .Z(n23698) );
  XNOR U32328 ( .A(y[4996]), .B(x[4996]), .Z(n23701) );
  XNOR U32329 ( .A(y[4997]), .B(x[4997]), .Z(n23700) );
  XOR U32330 ( .A(n23674), .B(n23675), .Z(n23693) );
  XNOR U32331 ( .A(n23690), .B(n23691), .Z(n23675) );
  XNOR U32332 ( .A(n23685), .B(n23686), .Z(n23691) );
  XNOR U32333 ( .A(n23687), .B(n23688), .Z(n23686) );
  XNOR U32334 ( .A(y[4993]), .B(x[4993]), .Z(n23688) );
  XNOR U32335 ( .A(y[4994]), .B(x[4994]), .Z(n23687) );
  XNOR U32336 ( .A(y[4992]), .B(x[4992]), .Z(n23685) );
  XNOR U32337 ( .A(n23679), .B(n23680), .Z(n23690) );
  XNOR U32338 ( .A(y[4989]), .B(x[4989]), .Z(n23680) );
  XNOR U32339 ( .A(n23681), .B(n23682), .Z(n23679) );
  XNOR U32340 ( .A(y[4990]), .B(x[4990]), .Z(n23682) );
  XNOR U32341 ( .A(y[4991]), .B(x[4991]), .Z(n23681) );
  XOR U32342 ( .A(n23673), .B(n23672), .Z(n23674) );
  XNOR U32343 ( .A(n23668), .B(n23669), .Z(n23672) );
  XNOR U32344 ( .A(y[4986]), .B(x[4986]), .Z(n23669) );
  XNOR U32345 ( .A(n23670), .B(n23671), .Z(n23668) );
  XNOR U32346 ( .A(y[4987]), .B(x[4987]), .Z(n23671) );
  XNOR U32347 ( .A(y[4988]), .B(x[4988]), .Z(n23670) );
  XNOR U32348 ( .A(n23662), .B(n23663), .Z(n23673) );
  XNOR U32349 ( .A(y[4983]), .B(x[4983]), .Z(n23663) );
  XNOR U32350 ( .A(n23664), .B(n23665), .Z(n23662) );
  XNOR U32351 ( .A(y[4984]), .B(x[4984]), .Z(n23665) );
  XNOR U32352 ( .A(y[4985]), .B(x[4985]), .Z(n23664) );
  NAND U32353 ( .A(n23729), .B(n23730), .Z(N63287) );
  NANDN U32354 ( .A(n23731), .B(n23732), .Z(n23730) );
  OR U32355 ( .A(n23733), .B(n23734), .Z(n23732) );
  NAND U32356 ( .A(n23733), .B(n23734), .Z(n23729) );
  XOR U32357 ( .A(n23733), .B(n23735), .Z(N63286) );
  XNOR U32358 ( .A(n23731), .B(n23734), .Z(n23735) );
  AND U32359 ( .A(n23736), .B(n23737), .Z(n23734) );
  NANDN U32360 ( .A(n23738), .B(n23739), .Z(n23737) );
  NANDN U32361 ( .A(n23740), .B(n23741), .Z(n23739) );
  NANDN U32362 ( .A(n23741), .B(n23740), .Z(n23736) );
  NAND U32363 ( .A(n23742), .B(n23743), .Z(n23731) );
  NANDN U32364 ( .A(n23744), .B(n23745), .Z(n23743) );
  OR U32365 ( .A(n23746), .B(n23747), .Z(n23745) );
  NAND U32366 ( .A(n23747), .B(n23746), .Z(n23742) );
  AND U32367 ( .A(n23748), .B(n23749), .Z(n23733) );
  NANDN U32368 ( .A(n23750), .B(n23751), .Z(n23749) );
  NANDN U32369 ( .A(n23752), .B(n23753), .Z(n23751) );
  NANDN U32370 ( .A(n23753), .B(n23752), .Z(n23748) );
  XOR U32371 ( .A(n23747), .B(n23754), .Z(N63285) );
  XOR U32372 ( .A(n23744), .B(n23746), .Z(n23754) );
  XNOR U32373 ( .A(n23740), .B(n23755), .Z(n23746) );
  XNOR U32374 ( .A(n23738), .B(n23741), .Z(n23755) );
  NAND U32375 ( .A(n23756), .B(n23757), .Z(n23741) );
  NAND U32376 ( .A(n23758), .B(n23759), .Z(n23757) );
  OR U32377 ( .A(n23760), .B(n23761), .Z(n23758) );
  NANDN U32378 ( .A(n23762), .B(n23760), .Z(n23756) );
  IV U32379 ( .A(n23761), .Z(n23762) );
  NAND U32380 ( .A(n23763), .B(n23764), .Z(n23738) );
  NAND U32381 ( .A(n23765), .B(n23766), .Z(n23764) );
  NANDN U32382 ( .A(n23767), .B(n23768), .Z(n23765) );
  NANDN U32383 ( .A(n23768), .B(n23767), .Z(n23763) );
  AND U32384 ( .A(n23769), .B(n23770), .Z(n23740) );
  NAND U32385 ( .A(n23771), .B(n23772), .Z(n23770) );
  OR U32386 ( .A(n23773), .B(n23774), .Z(n23771) );
  NANDN U32387 ( .A(n23775), .B(n23773), .Z(n23769) );
  NAND U32388 ( .A(n23776), .B(n23777), .Z(n23744) );
  NANDN U32389 ( .A(n23778), .B(n23779), .Z(n23777) );
  OR U32390 ( .A(n23780), .B(n23781), .Z(n23779) );
  NANDN U32391 ( .A(n23782), .B(n23780), .Z(n23776) );
  IV U32392 ( .A(n23781), .Z(n23782) );
  XNOR U32393 ( .A(n23752), .B(n23783), .Z(n23747) );
  XNOR U32394 ( .A(n23750), .B(n23753), .Z(n23783) );
  NAND U32395 ( .A(n23784), .B(n23785), .Z(n23753) );
  NAND U32396 ( .A(n23786), .B(n23787), .Z(n23785) );
  OR U32397 ( .A(n23788), .B(n23789), .Z(n23786) );
  NANDN U32398 ( .A(n23790), .B(n23788), .Z(n23784) );
  IV U32399 ( .A(n23789), .Z(n23790) );
  NAND U32400 ( .A(n23791), .B(n23792), .Z(n23750) );
  NAND U32401 ( .A(n23793), .B(n23794), .Z(n23792) );
  NANDN U32402 ( .A(n23795), .B(n23796), .Z(n23793) );
  NANDN U32403 ( .A(n23796), .B(n23795), .Z(n23791) );
  AND U32404 ( .A(n23797), .B(n23798), .Z(n23752) );
  NAND U32405 ( .A(n23799), .B(n23800), .Z(n23798) );
  OR U32406 ( .A(n23801), .B(n23802), .Z(n23799) );
  NANDN U32407 ( .A(n23803), .B(n23801), .Z(n23797) );
  XNOR U32408 ( .A(n23778), .B(n23804), .Z(N63284) );
  XOR U32409 ( .A(n23780), .B(n23781), .Z(n23804) );
  XNOR U32410 ( .A(n23794), .B(n23805), .Z(n23781) );
  XOR U32411 ( .A(n23795), .B(n23796), .Z(n23805) );
  XOR U32412 ( .A(n23801), .B(n23806), .Z(n23796) );
  XOR U32413 ( .A(n23800), .B(n23803), .Z(n23806) );
  IV U32414 ( .A(n23802), .Z(n23803) );
  NAND U32415 ( .A(n23807), .B(n23808), .Z(n23802) );
  OR U32416 ( .A(n23809), .B(n23810), .Z(n23808) );
  OR U32417 ( .A(n23811), .B(n23812), .Z(n23807) );
  NAND U32418 ( .A(n23813), .B(n23814), .Z(n23800) );
  OR U32419 ( .A(n23815), .B(n23816), .Z(n23814) );
  OR U32420 ( .A(n23817), .B(n23818), .Z(n23813) );
  NOR U32421 ( .A(n23819), .B(n23820), .Z(n23801) );
  ANDN U32422 ( .B(n23821), .A(n23822), .Z(n23795) );
  XNOR U32423 ( .A(n23788), .B(n23823), .Z(n23794) );
  XNOR U32424 ( .A(n23787), .B(n23789), .Z(n23823) );
  NAND U32425 ( .A(n23824), .B(n23825), .Z(n23789) );
  OR U32426 ( .A(n23826), .B(n23827), .Z(n23825) );
  OR U32427 ( .A(n23828), .B(n23829), .Z(n23824) );
  NAND U32428 ( .A(n23830), .B(n23831), .Z(n23787) );
  OR U32429 ( .A(n23832), .B(n23833), .Z(n23831) );
  OR U32430 ( .A(n23834), .B(n23835), .Z(n23830) );
  ANDN U32431 ( .B(n23836), .A(n23837), .Z(n23788) );
  IV U32432 ( .A(n23838), .Z(n23836) );
  ANDN U32433 ( .B(n23839), .A(n23840), .Z(n23780) );
  XOR U32434 ( .A(n23766), .B(n23841), .Z(n23778) );
  XOR U32435 ( .A(n23767), .B(n23768), .Z(n23841) );
  XOR U32436 ( .A(n23773), .B(n23842), .Z(n23768) );
  XOR U32437 ( .A(n23772), .B(n23775), .Z(n23842) );
  IV U32438 ( .A(n23774), .Z(n23775) );
  NAND U32439 ( .A(n23843), .B(n23844), .Z(n23774) );
  OR U32440 ( .A(n23845), .B(n23846), .Z(n23844) );
  OR U32441 ( .A(n23847), .B(n23848), .Z(n23843) );
  NAND U32442 ( .A(n23849), .B(n23850), .Z(n23772) );
  OR U32443 ( .A(n23851), .B(n23852), .Z(n23850) );
  OR U32444 ( .A(n23853), .B(n23854), .Z(n23849) );
  NOR U32445 ( .A(n23855), .B(n23856), .Z(n23773) );
  ANDN U32446 ( .B(n23857), .A(n23858), .Z(n23767) );
  IV U32447 ( .A(n23859), .Z(n23857) );
  XNOR U32448 ( .A(n23760), .B(n23860), .Z(n23766) );
  XNOR U32449 ( .A(n23759), .B(n23761), .Z(n23860) );
  NAND U32450 ( .A(n23861), .B(n23862), .Z(n23761) );
  OR U32451 ( .A(n23863), .B(n23864), .Z(n23862) );
  OR U32452 ( .A(n23865), .B(n23866), .Z(n23861) );
  NAND U32453 ( .A(n23867), .B(n23868), .Z(n23759) );
  OR U32454 ( .A(n23869), .B(n23870), .Z(n23868) );
  OR U32455 ( .A(n23871), .B(n23872), .Z(n23867) );
  ANDN U32456 ( .B(n23873), .A(n23874), .Z(n23760) );
  IV U32457 ( .A(n23875), .Z(n23873) );
  XNOR U32458 ( .A(n23840), .B(n23839), .Z(N63283) );
  XOR U32459 ( .A(n23859), .B(n23858), .Z(n23839) );
  XNOR U32460 ( .A(n23874), .B(n23875), .Z(n23858) );
  XNOR U32461 ( .A(n23869), .B(n23870), .Z(n23875) );
  XNOR U32462 ( .A(n23871), .B(n23872), .Z(n23870) );
  XNOR U32463 ( .A(y[4981]), .B(x[4981]), .Z(n23872) );
  XNOR U32464 ( .A(y[4982]), .B(x[4982]), .Z(n23871) );
  XNOR U32465 ( .A(y[4980]), .B(x[4980]), .Z(n23869) );
  XNOR U32466 ( .A(n23863), .B(n23864), .Z(n23874) );
  XNOR U32467 ( .A(y[4977]), .B(x[4977]), .Z(n23864) );
  XNOR U32468 ( .A(n23865), .B(n23866), .Z(n23863) );
  XNOR U32469 ( .A(y[4978]), .B(x[4978]), .Z(n23866) );
  XNOR U32470 ( .A(y[4979]), .B(x[4979]), .Z(n23865) );
  XNOR U32471 ( .A(n23856), .B(n23855), .Z(n23859) );
  XNOR U32472 ( .A(n23851), .B(n23852), .Z(n23855) );
  XNOR U32473 ( .A(y[4974]), .B(x[4974]), .Z(n23852) );
  XNOR U32474 ( .A(n23853), .B(n23854), .Z(n23851) );
  XNOR U32475 ( .A(y[4975]), .B(x[4975]), .Z(n23854) );
  XNOR U32476 ( .A(y[4976]), .B(x[4976]), .Z(n23853) );
  XNOR U32477 ( .A(n23845), .B(n23846), .Z(n23856) );
  XNOR U32478 ( .A(y[4971]), .B(x[4971]), .Z(n23846) );
  XNOR U32479 ( .A(n23847), .B(n23848), .Z(n23845) );
  XNOR U32480 ( .A(y[4972]), .B(x[4972]), .Z(n23848) );
  XNOR U32481 ( .A(y[4973]), .B(x[4973]), .Z(n23847) );
  XOR U32482 ( .A(n23821), .B(n23822), .Z(n23840) );
  XNOR U32483 ( .A(n23837), .B(n23838), .Z(n23822) );
  XNOR U32484 ( .A(n23832), .B(n23833), .Z(n23838) );
  XNOR U32485 ( .A(n23834), .B(n23835), .Z(n23833) );
  XNOR U32486 ( .A(y[4969]), .B(x[4969]), .Z(n23835) );
  XNOR U32487 ( .A(y[4970]), .B(x[4970]), .Z(n23834) );
  XNOR U32488 ( .A(y[4968]), .B(x[4968]), .Z(n23832) );
  XNOR U32489 ( .A(n23826), .B(n23827), .Z(n23837) );
  XNOR U32490 ( .A(y[4965]), .B(x[4965]), .Z(n23827) );
  XNOR U32491 ( .A(n23828), .B(n23829), .Z(n23826) );
  XNOR U32492 ( .A(y[4966]), .B(x[4966]), .Z(n23829) );
  XNOR U32493 ( .A(y[4967]), .B(x[4967]), .Z(n23828) );
  XOR U32494 ( .A(n23820), .B(n23819), .Z(n23821) );
  XNOR U32495 ( .A(n23815), .B(n23816), .Z(n23819) );
  XNOR U32496 ( .A(y[4962]), .B(x[4962]), .Z(n23816) );
  XNOR U32497 ( .A(n23817), .B(n23818), .Z(n23815) );
  XNOR U32498 ( .A(y[4963]), .B(x[4963]), .Z(n23818) );
  XNOR U32499 ( .A(y[4964]), .B(x[4964]), .Z(n23817) );
  XNOR U32500 ( .A(n23809), .B(n23810), .Z(n23820) );
  XNOR U32501 ( .A(y[4959]), .B(x[4959]), .Z(n23810) );
  XNOR U32502 ( .A(n23811), .B(n23812), .Z(n23809) );
  XNOR U32503 ( .A(y[4960]), .B(x[4960]), .Z(n23812) );
  XNOR U32504 ( .A(y[4961]), .B(x[4961]), .Z(n23811) );
  NAND U32505 ( .A(n23876), .B(n23877), .Z(N63274) );
  NANDN U32506 ( .A(n23878), .B(n23879), .Z(n23877) );
  OR U32507 ( .A(n23880), .B(n23881), .Z(n23879) );
  NAND U32508 ( .A(n23880), .B(n23881), .Z(n23876) );
  XOR U32509 ( .A(n23880), .B(n23882), .Z(N63273) );
  XNOR U32510 ( .A(n23878), .B(n23881), .Z(n23882) );
  AND U32511 ( .A(n23883), .B(n23884), .Z(n23881) );
  NANDN U32512 ( .A(n23885), .B(n23886), .Z(n23884) );
  NANDN U32513 ( .A(n23887), .B(n23888), .Z(n23886) );
  NANDN U32514 ( .A(n23888), .B(n23887), .Z(n23883) );
  NAND U32515 ( .A(n23889), .B(n23890), .Z(n23878) );
  NANDN U32516 ( .A(n23891), .B(n23892), .Z(n23890) );
  OR U32517 ( .A(n23893), .B(n23894), .Z(n23892) );
  NAND U32518 ( .A(n23894), .B(n23893), .Z(n23889) );
  AND U32519 ( .A(n23895), .B(n23896), .Z(n23880) );
  NANDN U32520 ( .A(n23897), .B(n23898), .Z(n23896) );
  NANDN U32521 ( .A(n23899), .B(n23900), .Z(n23898) );
  NANDN U32522 ( .A(n23900), .B(n23899), .Z(n23895) );
  XOR U32523 ( .A(n23894), .B(n23901), .Z(N63272) );
  XOR U32524 ( .A(n23891), .B(n23893), .Z(n23901) );
  XNOR U32525 ( .A(n23887), .B(n23902), .Z(n23893) );
  XNOR U32526 ( .A(n23885), .B(n23888), .Z(n23902) );
  NAND U32527 ( .A(n23903), .B(n23904), .Z(n23888) );
  NAND U32528 ( .A(n23905), .B(n23906), .Z(n23904) );
  OR U32529 ( .A(n23907), .B(n23908), .Z(n23905) );
  NANDN U32530 ( .A(n23909), .B(n23907), .Z(n23903) );
  IV U32531 ( .A(n23908), .Z(n23909) );
  NAND U32532 ( .A(n23910), .B(n23911), .Z(n23885) );
  NAND U32533 ( .A(n23912), .B(n23913), .Z(n23911) );
  NANDN U32534 ( .A(n23914), .B(n23915), .Z(n23912) );
  NANDN U32535 ( .A(n23915), .B(n23914), .Z(n23910) );
  AND U32536 ( .A(n23916), .B(n23917), .Z(n23887) );
  NAND U32537 ( .A(n23918), .B(n23919), .Z(n23917) );
  OR U32538 ( .A(n23920), .B(n23921), .Z(n23918) );
  NANDN U32539 ( .A(n23922), .B(n23920), .Z(n23916) );
  NAND U32540 ( .A(n23923), .B(n23924), .Z(n23891) );
  NANDN U32541 ( .A(n23925), .B(n23926), .Z(n23924) );
  OR U32542 ( .A(n23927), .B(n23928), .Z(n23926) );
  NANDN U32543 ( .A(n23929), .B(n23927), .Z(n23923) );
  IV U32544 ( .A(n23928), .Z(n23929) );
  XNOR U32545 ( .A(n23899), .B(n23930), .Z(n23894) );
  XNOR U32546 ( .A(n23897), .B(n23900), .Z(n23930) );
  NAND U32547 ( .A(n23931), .B(n23932), .Z(n23900) );
  NAND U32548 ( .A(n23933), .B(n23934), .Z(n23932) );
  OR U32549 ( .A(n23935), .B(n23936), .Z(n23933) );
  NANDN U32550 ( .A(n23937), .B(n23935), .Z(n23931) );
  IV U32551 ( .A(n23936), .Z(n23937) );
  NAND U32552 ( .A(n23938), .B(n23939), .Z(n23897) );
  NAND U32553 ( .A(n23940), .B(n23941), .Z(n23939) );
  NANDN U32554 ( .A(n23942), .B(n23943), .Z(n23940) );
  NANDN U32555 ( .A(n23943), .B(n23942), .Z(n23938) );
  AND U32556 ( .A(n23944), .B(n23945), .Z(n23899) );
  NAND U32557 ( .A(n23946), .B(n23947), .Z(n23945) );
  OR U32558 ( .A(n23948), .B(n23949), .Z(n23946) );
  NANDN U32559 ( .A(n23950), .B(n23948), .Z(n23944) );
  XNOR U32560 ( .A(n23925), .B(n23951), .Z(N63271) );
  XOR U32561 ( .A(n23927), .B(n23928), .Z(n23951) );
  XNOR U32562 ( .A(n23941), .B(n23952), .Z(n23928) );
  XOR U32563 ( .A(n23942), .B(n23943), .Z(n23952) );
  XOR U32564 ( .A(n23948), .B(n23953), .Z(n23943) );
  XOR U32565 ( .A(n23947), .B(n23950), .Z(n23953) );
  IV U32566 ( .A(n23949), .Z(n23950) );
  NAND U32567 ( .A(n23954), .B(n23955), .Z(n23949) );
  OR U32568 ( .A(n23956), .B(n23957), .Z(n23955) );
  OR U32569 ( .A(n23958), .B(n23959), .Z(n23954) );
  NAND U32570 ( .A(n23960), .B(n23961), .Z(n23947) );
  OR U32571 ( .A(n23962), .B(n23963), .Z(n23961) );
  OR U32572 ( .A(n23964), .B(n23965), .Z(n23960) );
  NOR U32573 ( .A(n23966), .B(n23967), .Z(n23948) );
  ANDN U32574 ( .B(n23968), .A(n23969), .Z(n23942) );
  XNOR U32575 ( .A(n23935), .B(n23970), .Z(n23941) );
  XNOR U32576 ( .A(n23934), .B(n23936), .Z(n23970) );
  NAND U32577 ( .A(n23971), .B(n23972), .Z(n23936) );
  OR U32578 ( .A(n23973), .B(n23974), .Z(n23972) );
  OR U32579 ( .A(n23975), .B(n23976), .Z(n23971) );
  NAND U32580 ( .A(n23977), .B(n23978), .Z(n23934) );
  OR U32581 ( .A(n23979), .B(n23980), .Z(n23978) );
  OR U32582 ( .A(n23981), .B(n23982), .Z(n23977) );
  ANDN U32583 ( .B(n23983), .A(n23984), .Z(n23935) );
  IV U32584 ( .A(n23985), .Z(n23983) );
  ANDN U32585 ( .B(n23986), .A(n23987), .Z(n23927) );
  XOR U32586 ( .A(n23913), .B(n23988), .Z(n23925) );
  XOR U32587 ( .A(n23914), .B(n23915), .Z(n23988) );
  XOR U32588 ( .A(n23920), .B(n23989), .Z(n23915) );
  XOR U32589 ( .A(n23919), .B(n23922), .Z(n23989) );
  IV U32590 ( .A(n23921), .Z(n23922) );
  NAND U32591 ( .A(n23990), .B(n23991), .Z(n23921) );
  OR U32592 ( .A(n23992), .B(n23993), .Z(n23991) );
  OR U32593 ( .A(n23994), .B(n23995), .Z(n23990) );
  NAND U32594 ( .A(n23996), .B(n23997), .Z(n23919) );
  OR U32595 ( .A(n23998), .B(n23999), .Z(n23997) );
  OR U32596 ( .A(n24000), .B(n24001), .Z(n23996) );
  NOR U32597 ( .A(n24002), .B(n24003), .Z(n23920) );
  ANDN U32598 ( .B(n24004), .A(n24005), .Z(n23914) );
  IV U32599 ( .A(n24006), .Z(n24004) );
  XNOR U32600 ( .A(n23907), .B(n24007), .Z(n23913) );
  XNOR U32601 ( .A(n23906), .B(n23908), .Z(n24007) );
  NAND U32602 ( .A(n24008), .B(n24009), .Z(n23908) );
  OR U32603 ( .A(n24010), .B(n24011), .Z(n24009) );
  OR U32604 ( .A(n24012), .B(n24013), .Z(n24008) );
  NAND U32605 ( .A(n24014), .B(n24015), .Z(n23906) );
  OR U32606 ( .A(n24016), .B(n24017), .Z(n24015) );
  OR U32607 ( .A(n24018), .B(n24019), .Z(n24014) );
  ANDN U32608 ( .B(n24020), .A(n24021), .Z(n23907) );
  IV U32609 ( .A(n24022), .Z(n24020) );
  XNOR U32610 ( .A(n23987), .B(n23986), .Z(N63270) );
  XOR U32611 ( .A(n24006), .B(n24005), .Z(n23986) );
  XNOR U32612 ( .A(n24021), .B(n24022), .Z(n24005) );
  XNOR U32613 ( .A(n24016), .B(n24017), .Z(n24022) );
  XNOR U32614 ( .A(n24018), .B(n24019), .Z(n24017) );
  XNOR U32615 ( .A(y[4957]), .B(x[4957]), .Z(n24019) );
  XNOR U32616 ( .A(y[4958]), .B(x[4958]), .Z(n24018) );
  XNOR U32617 ( .A(y[4956]), .B(x[4956]), .Z(n24016) );
  XNOR U32618 ( .A(n24010), .B(n24011), .Z(n24021) );
  XNOR U32619 ( .A(y[4953]), .B(x[4953]), .Z(n24011) );
  XNOR U32620 ( .A(n24012), .B(n24013), .Z(n24010) );
  XNOR U32621 ( .A(y[4954]), .B(x[4954]), .Z(n24013) );
  XNOR U32622 ( .A(y[4955]), .B(x[4955]), .Z(n24012) );
  XNOR U32623 ( .A(n24003), .B(n24002), .Z(n24006) );
  XNOR U32624 ( .A(n23998), .B(n23999), .Z(n24002) );
  XNOR U32625 ( .A(y[4950]), .B(x[4950]), .Z(n23999) );
  XNOR U32626 ( .A(n24000), .B(n24001), .Z(n23998) );
  XNOR U32627 ( .A(y[4951]), .B(x[4951]), .Z(n24001) );
  XNOR U32628 ( .A(y[4952]), .B(x[4952]), .Z(n24000) );
  XNOR U32629 ( .A(n23992), .B(n23993), .Z(n24003) );
  XNOR U32630 ( .A(y[4947]), .B(x[4947]), .Z(n23993) );
  XNOR U32631 ( .A(n23994), .B(n23995), .Z(n23992) );
  XNOR U32632 ( .A(y[4948]), .B(x[4948]), .Z(n23995) );
  XNOR U32633 ( .A(y[4949]), .B(x[4949]), .Z(n23994) );
  XOR U32634 ( .A(n23968), .B(n23969), .Z(n23987) );
  XNOR U32635 ( .A(n23984), .B(n23985), .Z(n23969) );
  XNOR U32636 ( .A(n23979), .B(n23980), .Z(n23985) );
  XNOR U32637 ( .A(n23981), .B(n23982), .Z(n23980) );
  XNOR U32638 ( .A(y[4945]), .B(x[4945]), .Z(n23982) );
  XNOR U32639 ( .A(y[4946]), .B(x[4946]), .Z(n23981) );
  XNOR U32640 ( .A(y[4944]), .B(x[4944]), .Z(n23979) );
  XNOR U32641 ( .A(n23973), .B(n23974), .Z(n23984) );
  XNOR U32642 ( .A(y[4941]), .B(x[4941]), .Z(n23974) );
  XNOR U32643 ( .A(n23975), .B(n23976), .Z(n23973) );
  XNOR U32644 ( .A(y[4942]), .B(x[4942]), .Z(n23976) );
  XNOR U32645 ( .A(y[4943]), .B(x[4943]), .Z(n23975) );
  XOR U32646 ( .A(n23967), .B(n23966), .Z(n23968) );
  XNOR U32647 ( .A(n23962), .B(n23963), .Z(n23966) );
  XNOR U32648 ( .A(y[4938]), .B(x[4938]), .Z(n23963) );
  XNOR U32649 ( .A(n23964), .B(n23965), .Z(n23962) );
  XNOR U32650 ( .A(y[4939]), .B(x[4939]), .Z(n23965) );
  XNOR U32651 ( .A(y[4940]), .B(x[4940]), .Z(n23964) );
  XNOR U32652 ( .A(n23956), .B(n23957), .Z(n23967) );
  XNOR U32653 ( .A(y[4935]), .B(x[4935]), .Z(n23957) );
  XNOR U32654 ( .A(n23958), .B(n23959), .Z(n23956) );
  XNOR U32655 ( .A(y[4936]), .B(x[4936]), .Z(n23959) );
  XNOR U32656 ( .A(y[4937]), .B(x[4937]), .Z(n23958) );
  NAND U32657 ( .A(n24023), .B(n24024), .Z(N63261) );
  NANDN U32658 ( .A(n24025), .B(n24026), .Z(n24024) );
  OR U32659 ( .A(n24027), .B(n24028), .Z(n24026) );
  NAND U32660 ( .A(n24027), .B(n24028), .Z(n24023) );
  XOR U32661 ( .A(n24027), .B(n24029), .Z(N63260) );
  XNOR U32662 ( .A(n24025), .B(n24028), .Z(n24029) );
  AND U32663 ( .A(n24030), .B(n24031), .Z(n24028) );
  NANDN U32664 ( .A(n24032), .B(n24033), .Z(n24031) );
  NANDN U32665 ( .A(n24034), .B(n24035), .Z(n24033) );
  NANDN U32666 ( .A(n24035), .B(n24034), .Z(n24030) );
  NAND U32667 ( .A(n24036), .B(n24037), .Z(n24025) );
  NANDN U32668 ( .A(n24038), .B(n24039), .Z(n24037) );
  OR U32669 ( .A(n24040), .B(n24041), .Z(n24039) );
  NAND U32670 ( .A(n24041), .B(n24040), .Z(n24036) );
  AND U32671 ( .A(n24042), .B(n24043), .Z(n24027) );
  NANDN U32672 ( .A(n24044), .B(n24045), .Z(n24043) );
  NANDN U32673 ( .A(n24046), .B(n24047), .Z(n24045) );
  NANDN U32674 ( .A(n24047), .B(n24046), .Z(n24042) );
  XOR U32675 ( .A(n24041), .B(n24048), .Z(N63259) );
  XOR U32676 ( .A(n24038), .B(n24040), .Z(n24048) );
  XNOR U32677 ( .A(n24034), .B(n24049), .Z(n24040) );
  XNOR U32678 ( .A(n24032), .B(n24035), .Z(n24049) );
  NAND U32679 ( .A(n24050), .B(n24051), .Z(n24035) );
  NAND U32680 ( .A(n24052), .B(n24053), .Z(n24051) );
  OR U32681 ( .A(n24054), .B(n24055), .Z(n24052) );
  NANDN U32682 ( .A(n24056), .B(n24054), .Z(n24050) );
  IV U32683 ( .A(n24055), .Z(n24056) );
  NAND U32684 ( .A(n24057), .B(n24058), .Z(n24032) );
  NAND U32685 ( .A(n24059), .B(n24060), .Z(n24058) );
  NANDN U32686 ( .A(n24061), .B(n24062), .Z(n24059) );
  NANDN U32687 ( .A(n24062), .B(n24061), .Z(n24057) );
  AND U32688 ( .A(n24063), .B(n24064), .Z(n24034) );
  NAND U32689 ( .A(n24065), .B(n24066), .Z(n24064) );
  OR U32690 ( .A(n24067), .B(n24068), .Z(n24065) );
  NANDN U32691 ( .A(n24069), .B(n24067), .Z(n24063) );
  NAND U32692 ( .A(n24070), .B(n24071), .Z(n24038) );
  NANDN U32693 ( .A(n24072), .B(n24073), .Z(n24071) );
  OR U32694 ( .A(n24074), .B(n24075), .Z(n24073) );
  NANDN U32695 ( .A(n24076), .B(n24074), .Z(n24070) );
  IV U32696 ( .A(n24075), .Z(n24076) );
  XNOR U32697 ( .A(n24046), .B(n24077), .Z(n24041) );
  XNOR U32698 ( .A(n24044), .B(n24047), .Z(n24077) );
  NAND U32699 ( .A(n24078), .B(n24079), .Z(n24047) );
  NAND U32700 ( .A(n24080), .B(n24081), .Z(n24079) );
  OR U32701 ( .A(n24082), .B(n24083), .Z(n24080) );
  NANDN U32702 ( .A(n24084), .B(n24082), .Z(n24078) );
  IV U32703 ( .A(n24083), .Z(n24084) );
  NAND U32704 ( .A(n24085), .B(n24086), .Z(n24044) );
  NAND U32705 ( .A(n24087), .B(n24088), .Z(n24086) );
  NANDN U32706 ( .A(n24089), .B(n24090), .Z(n24087) );
  NANDN U32707 ( .A(n24090), .B(n24089), .Z(n24085) );
  AND U32708 ( .A(n24091), .B(n24092), .Z(n24046) );
  NAND U32709 ( .A(n24093), .B(n24094), .Z(n24092) );
  OR U32710 ( .A(n24095), .B(n24096), .Z(n24093) );
  NANDN U32711 ( .A(n24097), .B(n24095), .Z(n24091) );
  XNOR U32712 ( .A(n24072), .B(n24098), .Z(N63258) );
  XOR U32713 ( .A(n24074), .B(n24075), .Z(n24098) );
  XNOR U32714 ( .A(n24088), .B(n24099), .Z(n24075) );
  XOR U32715 ( .A(n24089), .B(n24090), .Z(n24099) );
  XOR U32716 ( .A(n24095), .B(n24100), .Z(n24090) );
  XOR U32717 ( .A(n24094), .B(n24097), .Z(n24100) );
  IV U32718 ( .A(n24096), .Z(n24097) );
  NAND U32719 ( .A(n24101), .B(n24102), .Z(n24096) );
  OR U32720 ( .A(n24103), .B(n24104), .Z(n24102) );
  OR U32721 ( .A(n24105), .B(n24106), .Z(n24101) );
  NAND U32722 ( .A(n24107), .B(n24108), .Z(n24094) );
  OR U32723 ( .A(n24109), .B(n24110), .Z(n24108) );
  OR U32724 ( .A(n24111), .B(n24112), .Z(n24107) );
  NOR U32725 ( .A(n24113), .B(n24114), .Z(n24095) );
  ANDN U32726 ( .B(n24115), .A(n24116), .Z(n24089) );
  XNOR U32727 ( .A(n24082), .B(n24117), .Z(n24088) );
  XNOR U32728 ( .A(n24081), .B(n24083), .Z(n24117) );
  NAND U32729 ( .A(n24118), .B(n24119), .Z(n24083) );
  OR U32730 ( .A(n24120), .B(n24121), .Z(n24119) );
  OR U32731 ( .A(n24122), .B(n24123), .Z(n24118) );
  NAND U32732 ( .A(n24124), .B(n24125), .Z(n24081) );
  OR U32733 ( .A(n24126), .B(n24127), .Z(n24125) );
  OR U32734 ( .A(n24128), .B(n24129), .Z(n24124) );
  ANDN U32735 ( .B(n24130), .A(n24131), .Z(n24082) );
  IV U32736 ( .A(n24132), .Z(n24130) );
  ANDN U32737 ( .B(n24133), .A(n24134), .Z(n24074) );
  XOR U32738 ( .A(n24060), .B(n24135), .Z(n24072) );
  XOR U32739 ( .A(n24061), .B(n24062), .Z(n24135) );
  XOR U32740 ( .A(n24067), .B(n24136), .Z(n24062) );
  XOR U32741 ( .A(n24066), .B(n24069), .Z(n24136) );
  IV U32742 ( .A(n24068), .Z(n24069) );
  NAND U32743 ( .A(n24137), .B(n24138), .Z(n24068) );
  OR U32744 ( .A(n24139), .B(n24140), .Z(n24138) );
  OR U32745 ( .A(n24141), .B(n24142), .Z(n24137) );
  NAND U32746 ( .A(n24143), .B(n24144), .Z(n24066) );
  OR U32747 ( .A(n24145), .B(n24146), .Z(n24144) );
  OR U32748 ( .A(n24147), .B(n24148), .Z(n24143) );
  NOR U32749 ( .A(n24149), .B(n24150), .Z(n24067) );
  ANDN U32750 ( .B(n24151), .A(n24152), .Z(n24061) );
  IV U32751 ( .A(n24153), .Z(n24151) );
  XNOR U32752 ( .A(n24054), .B(n24154), .Z(n24060) );
  XNOR U32753 ( .A(n24053), .B(n24055), .Z(n24154) );
  NAND U32754 ( .A(n24155), .B(n24156), .Z(n24055) );
  OR U32755 ( .A(n24157), .B(n24158), .Z(n24156) );
  OR U32756 ( .A(n24159), .B(n24160), .Z(n24155) );
  NAND U32757 ( .A(n24161), .B(n24162), .Z(n24053) );
  OR U32758 ( .A(n24163), .B(n24164), .Z(n24162) );
  OR U32759 ( .A(n24165), .B(n24166), .Z(n24161) );
  ANDN U32760 ( .B(n24167), .A(n24168), .Z(n24054) );
  IV U32761 ( .A(n24169), .Z(n24167) );
  XNOR U32762 ( .A(n24134), .B(n24133), .Z(N63257) );
  XOR U32763 ( .A(n24153), .B(n24152), .Z(n24133) );
  XNOR U32764 ( .A(n24168), .B(n24169), .Z(n24152) );
  XNOR U32765 ( .A(n24163), .B(n24164), .Z(n24169) );
  XNOR U32766 ( .A(n24165), .B(n24166), .Z(n24164) );
  XNOR U32767 ( .A(y[4933]), .B(x[4933]), .Z(n24166) );
  XNOR U32768 ( .A(y[4934]), .B(x[4934]), .Z(n24165) );
  XNOR U32769 ( .A(y[4932]), .B(x[4932]), .Z(n24163) );
  XNOR U32770 ( .A(n24157), .B(n24158), .Z(n24168) );
  XNOR U32771 ( .A(y[4929]), .B(x[4929]), .Z(n24158) );
  XNOR U32772 ( .A(n24159), .B(n24160), .Z(n24157) );
  XNOR U32773 ( .A(y[4930]), .B(x[4930]), .Z(n24160) );
  XNOR U32774 ( .A(y[4931]), .B(x[4931]), .Z(n24159) );
  XNOR U32775 ( .A(n24150), .B(n24149), .Z(n24153) );
  XNOR U32776 ( .A(n24145), .B(n24146), .Z(n24149) );
  XNOR U32777 ( .A(y[4926]), .B(x[4926]), .Z(n24146) );
  XNOR U32778 ( .A(n24147), .B(n24148), .Z(n24145) );
  XNOR U32779 ( .A(y[4927]), .B(x[4927]), .Z(n24148) );
  XNOR U32780 ( .A(y[4928]), .B(x[4928]), .Z(n24147) );
  XNOR U32781 ( .A(n24139), .B(n24140), .Z(n24150) );
  XNOR U32782 ( .A(y[4923]), .B(x[4923]), .Z(n24140) );
  XNOR U32783 ( .A(n24141), .B(n24142), .Z(n24139) );
  XNOR U32784 ( .A(y[4924]), .B(x[4924]), .Z(n24142) );
  XNOR U32785 ( .A(y[4925]), .B(x[4925]), .Z(n24141) );
  XOR U32786 ( .A(n24115), .B(n24116), .Z(n24134) );
  XNOR U32787 ( .A(n24131), .B(n24132), .Z(n24116) );
  XNOR U32788 ( .A(n24126), .B(n24127), .Z(n24132) );
  XNOR U32789 ( .A(n24128), .B(n24129), .Z(n24127) );
  XNOR U32790 ( .A(y[4921]), .B(x[4921]), .Z(n24129) );
  XNOR U32791 ( .A(y[4922]), .B(x[4922]), .Z(n24128) );
  XNOR U32792 ( .A(y[4920]), .B(x[4920]), .Z(n24126) );
  XNOR U32793 ( .A(n24120), .B(n24121), .Z(n24131) );
  XNOR U32794 ( .A(y[4917]), .B(x[4917]), .Z(n24121) );
  XNOR U32795 ( .A(n24122), .B(n24123), .Z(n24120) );
  XNOR U32796 ( .A(y[4918]), .B(x[4918]), .Z(n24123) );
  XNOR U32797 ( .A(y[4919]), .B(x[4919]), .Z(n24122) );
  XOR U32798 ( .A(n24114), .B(n24113), .Z(n24115) );
  XNOR U32799 ( .A(n24109), .B(n24110), .Z(n24113) );
  XNOR U32800 ( .A(y[4914]), .B(x[4914]), .Z(n24110) );
  XNOR U32801 ( .A(n24111), .B(n24112), .Z(n24109) );
  XNOR U32802 ( .A(y[4915]), .B(x[4915]), .Z(n24112) );
  XNOR U32803 ( .A(y[4916]), .B(x[4916]), .Z(n24111) );
  XNOR U32804 ( .A(n24103), .B(n24104), .Z(n24114) );
  XNOR U32805 ( .A(y[4911]), .B(x[4911]), .Z(n24104) );
  XNOR U32806 ( .A(n24105), .B(n24106), .Z(n24103) );
  XNOR U32807 ( .A(y[4912]), .B(x[4912]), .Z(n24106) );
  XNOR U32808 ( .A(y[4913]), .B(x[4913]), .Z(n24105) );
  NAND U32809 ( .A(n24170), .B(n24171), .Z(N63248) );
  NANDN U32810 ( .A(n24172), .B(n24173), .Z(n24171) );
  OR U32811 ( .A(n24174), .B(n24175), .Z(n24173) );
  NAND U32812 ( .A(n24174), .B(n24175), .Z(n24170) );
  XOR U32813 ( .A(n24174), .B(n24176), .Z(N63247) );
  XNOR U32814 ( .A(n24172), .B(n24175), .Z(n24176) );
  AND U32815 ( .A(n24177), .B(n24178), .Z(n24175) );
  NANDN U32816 ( .A(n24179), .B(n24180), .Z(n24178) );
  NANDN U32817 ( .A(n24181), .B(n24182), .Z(n24180) );
  NANDN U32818 ( .A(n24182), .B(n24181), .Z(n24177) );
  NAND U32819 ( .A(n24183), .B(n24184), .Z(n24172) );
  NANDN U32820 ( .A(n24185), .B(n24186), .Z(n24184) );
  OR U32821 ( .A(n24187), .B(n24188), .Z(n24186) );
  NAND U32822 ( .A(n24188), .B(n24187), .Z(n24183) );
  AND U32823 ( .A(n24189), .B(n24190), .Z(n24174) );
  NANDN U32824 ( .A(n24191), .B(n24192), .Z(n24190) );
  NANDN U32825 ( .A(n24193), .B(n24194), .Z(n24192) );
  NANDN U32826 ( .A(n24194), .B(n24193), .Z(n24189) );
  XOR U32827 ( .A(n24188), .B(n24195), .Z(N63246) );
  XOR U32828 ( .A(n24185), .B(n24187), .Z(n24195) );
  XNOR U32829 ( .A(n24181), .B(n24196), .Z(n24187) );
  XNOR U32830 ( .A(n24179), .B(n24182), .Z(n24196) );
  NAND U32831 ( .A(n24197), .B(n24198), .Z(n24182) );
  NAND U32832 ( .A(n24199), .B(n24200), .Z(n24198) );
  OR U32833 ( .A(n24201), .B(n24202), .Z(n24199) );
  NANDN U32834 ( .A(n24203), .B(n24201), .Z(n24197) );
  IV U32835 ( .A(n24202), .Z(n24203) );
  NAND U32836 ( .A(n24204), .B(n24205), .Z(n24179) );
  NAND U32837 ( .A(n24206), .B(n24207), .Z(n24205) );
  NANDN U32838 ( .A(n24208), .B(n24209), .Z(n24206) );
  NANDN U32839 ( .A(n24209), .B(n24208), .Z(n24204) );
  AND U32840 ( .A(n24210), .B(n24211), .Z(n24181) );
  NAND U32841 ( .A(n24212), .B(n24213), .Z(n24211) );
  OR U32842 ( .A(n24214), .B(n24215), .Z(n24212) );
  NANDN U32843 ( .A(n24216), .B(n24214), .Z(n24210) );
  NAND U32844 ( .A(n24217), .B(n24218), .Z(n24185) );
  NANDN U32845 ( .A(n24219), .B(n24220), .Z(n24218) );
  OR U32846 ( .A(n24221), .B(n24222), .Z(n24220) );
  NANDN U32847 ( .A(n24223), .B(n24221), .Z(n24217) );
  IV U32848 ( .A(n24222), .Z(n24223) );
  XNOR U32849 ( .A(n24193), .B(n24224), .Z(n24188) );
  XNOR U32850 ( .A(n24191), .B(n24194), .Z(n24224) );
  NAND U32851 ( .A(n24225), .B(n24226), .Z(n24194) );
  NAND U32852 ( .A(n24227), .B(n24228), .Z(n24226) );
  OR U32853 ( .A(n24229), .B(n24230), .Z(n24227) );
  NANDN U32854 ( .A(n24231), .B(n24229), .Z(n24225) );
  IV U32855 ( .A(n24230), .Z(n24231) );
  NAND U32856 ( .A(n24232), .B(n24233), .Z(n24191) );
  NAND U32857 ( .A(n24234), .B(n24235), .Z(n24233) );
  NANDN U32858 ( .A(n24236), .B(n24237), .Z(n24234) );
  NANDN U32859 ( .A(n24237), .B(n24236), .Z(n24232) );
  AND U32860 ( .A(n24238), .B(n24239), .Z(n24193) );
  NAND U32861 ( .A(n24240), .B(n24241), .Z(n24239) );
  OR U32862 ( .A(n24242), .B(n24243), .Z(n24240) );
  NANDN U32863 ( .A(n24244), .B(n24242), .Z(n24238) );
  XNOR U32864 ( .A(n24219), .B(n24245), .Z(N63245) );
  XOR U32865 ( .A(n24221), .B(n24222), .Z(n24245) );
  XNOR U32866 ( .A(n24235), .B(n24246), .Z(n24222) );
  XOR U32867 ( .A(n24236), .B(n24237), .Z(n24246) );
  XOR U32868 ( .A(n24242), .B(n24247), .Z(n24237) );
  XOR U32869 ( .A(n24241), .B(n24244), .Z(n24247) );
  IV U32870 ( .A(n24243), .Z(n24244) );
  NAND U32871 ( .A(n24248), .B(n24249), .Z(n24243) );
  OR U32872 ( .A(n24250), .B(n24251), .Z(n24249) );
  OR U32873 ( .A(n24252), .B(n24253), .Z(n24248) );
  NAND U32874 ( .A(n24254), .B(n24255), .Z(n24241) );
  OR U32875 ( .A(n24256), .B(n24257), .Z(n24255) );
  OR U32876 ( .A(n24258), .B(n24259), .Z(n24254) );
  NOR U32877 ( .A(n24260), .B(n24261), .Z(n24242) );
  ANDN U32878 ( .B(n24262), .A(n24263), .Z(n24236) );
  XNOR U32879 ( .A(n24229), .B(n24264), .Z(n24235) );
  XNOR U32880 ( .A(n24228), .B(n24230), .Z(n24264) );
  NAND U32881 ( .A(n24265), .B(n24266), .Z(n24230) );
  OR U32882 ( .A(n24267), .B(n24268), .Z(n24266) );
  OR U32883 ( .A(n24269), .B(n24270), .Z(n24265) );
  NAND U32884 ( .A(n24271), .B(n24272), .Z(n24228) );
  OR U32885 ( .A(n24273), .B(n24274), .Z(n24272) );
  OR U32886 ( .A(n24275), .B(n24276), .Z(n24271) );
  ANDN U32887 ( .B(n24277), .A(n24278), .Z(n24229) );
  IV U32888 ( .A(n24279), .Z(n24277) );
  ANDN U32889 ( .B(n24280), .A(n24281), .Z(n24221) );
  XOR U32890 ( .A(n24207), .B(n24282), .Z(n24219) );
  XOR U32891 ( .A(n24208), .B(n24209), .Z(n24282) );
  XOR U32892 ( .A(n24214), .B(n24283), .Z(n24209) );
  XOR U32893 ( .A(n24213), .B(n24216), .Z(n24283) );
  IV U32894 ( .A(n24215), .Z(n24216) );
  NAND U32895 ( .A(n24284), .B(n24285), .Z(n24215) );
  OR U32896 ( .A(n24286), .B(n24287), .Z(n24285) );
  OR U32897 ( .A(n24288), .B(n24289), .Z(n24284) );
  NAND U32898 ( .A(n24290), .B(n24291), .Z(n24213) );
  OR U32899 ( .A(n24292), .B(n24293), .Z(n24291) );
  OR U32900 ( .A(n24294), .B(n24295), .Z(n24290) );
  NOR U32901 ( .A(n24296), .B(n24297), .Z(n24214) );
  ANDN U32902 ( .B(n24298), .A(n24299), .Z(n24208) );
  IV U32903 ( .A(n24300), .Z(n24298) );
  XNOR U32904 ( .A(n24201), .B(n24301), .Z(n24207) );
  XNOR U32905 ( .A(n24200), .B(n24202), .Z(n24301) );
  NAND U32906 ( .A(n24302), .B(n24303), .Z(n24202) );
  OR U32907 ( .A(n24304), .B(n24305), .Z(n24303) );
  OR U32908 ( .A(n24306), .B(n24307), .Z(n24302) );
  NAND U32909 ( .A(n24308), .B(n24309), .Z(n24200) );
  OR U32910 ( .A(n24310), .B(n24311), .Z(n24309) );
  OR U32911 ( .A(n24312), .B(n24313), .Z(n24308) );
  ANDN U32912 ( .B(n24314), .A(n24315), .Z(n24201) );
  IV U32913 ( .A(n24316), .Z(n24314) );
  XNOR U32914 ( .A(n24281), .B(n24280), .Z(N63244) );
  XOR U32915 ( .A(n24300), .B(n24299), .Z(n24280) );
  XNOR U32916 ( .A(n24315), .B(n24316), .Z(n24299) );
  XNOR U32917 ( .A(n24310), .B(n24311), .Z(n24316) );
  XNOR U32918 ( .A(n24312), .B(n24313), .Z(n24311) );
  XNOR U32919 ( .A(y[4909]), .B(x[4909]), .Z(n24313) );
  XNOR U32920 ( .A(y[4910]), .B(x[4910]), .Z(n24312) );
  XNOR U32921 ( .A(y[4908]), .B(x[4908]), .Z(n24310) );
  XNOR U32922 ( .A(n24304), .B(n24305), .Z(n24315) );
  XNOR U32923 ( .A(y[4905]), .B(x[4905]), .Z(n24305) );
  XNOR U32924 ( .A(n24306), .B(n24307), .Z(n24304) );
  XNOR U32925 ( .A(y[4906]), .B(x[4906]), .Z(n24307) );
  XNOR U32926 ( .A(y[4907]), .B(x[4907]), .Z(n24306) );
  XNOR U32927 ( .A(n24297), .B(n24296), .Z(n24300) );
  XNOR U32928 ( .A(n24292), .B(n24293), .Z(n24296) );
  XNOR U32929 ( .A(y[4902]), .B(x[4902]), .Z(n24293) );
  XNOR U32930 ( .A(n24294), .B(n24295), .Z(n24292) );
  XNOR U32931 ( .A(y[4903]), .B(x[4903]), .Z(n24295) );
  XNOR U32932 ( .A(y[4904]), .B(x[4904]), .Z(n24294) );
  XNOR U32933 ( .A(n24286), .B(n24287), .Z(n24297) );
  XNOR U32934 ( .A(y[4899]), .B(x[4899]), .Z(n24287) );
  XNOR U32935 ( .A(n24288), .B(n24289), .Z(n24286) );
  XNOR U32936 ( .A(y[4900]), .B(x[4900]), .Z(n24289) );
  XNOR U32937 ( .A(y[4901]), .B(x[4901]), .Z(n24288) );
  XOR U32938 ( .A(n24262), .B(n24263), .Z(n24281) );
  XNOR U32939 ( .A(n24278), .B(n24279), .Z(n24263) );
  XNOR U32940 ( .A(n24273), .B(n24274), .Z(n24279) );
  XNOR U32941 ( .A(n24275), .B(n24276), .Z(n24274) );
  XNOR U32942 ( .A(y[4897]), .B(x[4897]), .Z(n24276) );
  XNOR U32943 ( .A(y[4898]), .B(x[4898]), .Z(n24275) );
  XNOR U32944 ( .A(y[4896]), .B(x[4896]), .Z(n24273) );
  XNOR U32945 ( .A(n24267), .B(n24268), .Z(n24278) );
  XNOR U32946 ( .A(y[4893]), .B(x[4893]), .Z(n24268) );
  XNOR U32947 ( .A(n24269), .B(n24270), .Z(n24267) );
  XNOR U32948 ( .A(y[4894]), .B(x[4894]), .Z(n24270) );
  XNOR U32949 ( .A(y[4895]), .B(x[4895]), .Z(n24269) );
  XOR U32950 ( .A(n24261), .B(n24260), .Z(n24262) );
  XNOR U32951 ( .A(n24256), .B(n24257), .Z(n24260) );
  XNOR U32952 ( .A(y[4890]), .B(x[4890]), .Z(n24257) );
  XNOR U32953 ( .A(n24258), .B(n24259), .Z(n24256) );
  XNOR U32954 ( .A(y[4891]), .B(x[4891]), .Z(n24259) );
  XNOR U32955 ( .A(y[4892]), .B(x[4892]), .Z(n24258) );
  XNOR U32956 ( .A(n24250), .B(n24251), .Z(n24261) );
  XNOR U32957 ( .A(y[4887]), .B(x[4887]), .Z(n24251) );
  XNOR U32958 ( .A(n24252), .B(n24253), .Z(n24250) );
  XNOR U32959 ( .A(y[4888]), .B(x[4888]), .Z(n24253) );
  XNOR U32960 ( .A(y[4889]), .B(x[4889]), .Z(n24252) );
  NAND U32961 ( .A(n24317), .B(n24318), .Z(N63235) );
  NANDN U32962 ( .A(n24319), .B(n24320), .Z(n24318) );
  OR U32963 ( .A(n24321), .B(n24322), .Z(n24320) );
  NAND U32964 ( .A(n24321), .B(n24322), .Z(n24317) );
  XOR U32965 ( .A(n24321), .B(n24323), .Z(N63234) );
  XNOR U32966 ( .A(n24319), .B(n24322), .Z(n24323) );
  AND U32967 ( .A(n24324), .B(n24325), .Z(n24322) );
  NANDN U32968 ( .A(n24326), .B(n24327), .Z(n24325) );
  NANDN U32969 ( .A(n24328), .B(n24329), .Z(n24327) );
  NANDN U32970 ( .A(n24329), .B(n24328), .Z(n24324) );
  NAND U32971 ( .A(n24330), .B(n24331), .Z(n24319) );
  NANDN U32972 ( .A(n24332), .B(n24333), .Z(n24331) );
  OR U32973 ( .A(n24334), .B(n24335), .Z(n24333) );
  NAND U32974 ( .A(n24335), .B(n24334), .Z(n24330) );
  AND U32975 ( .A(n24336), .B(n24337), .Z(n24321) );
  NANDN U32976 ( .A(n24338), .B(n24339), .Z(n24337) );
  NANDN U32977 ( .A(n24340), .B(n24341), .Z(n24339) );
  NANDN U32978 ( .A(n24341), .B(n24340), .Z(n24336) );
  XOR U32979 ( .A(n24335), .B(n24342), .Z(N63233) );
  XOR U32980 ( .A(n24332), .B(n24334), .Z(n24342) );
  XNOR U32981 ( .A(n24328), .B(n24343), .Z(n24334) );
  XNOR U32982 ( .A(n24326), .B(n24329), .Z(n24343) );
  NAND U32983 ( .A(n24344), .B(n24345), .Z(n24329) );
  NAND U32984 ( .A(n24346), .B(n24347), .Z(n24345) );
  OR U32985 ( .A(n24348), .B(n24349), .Z(n24346) );
  NANDN U32986 ( .A(n24350), .B(n24348), .Z(n24344) );
  IV U32987 ( .A(n24349), .Z(n24350) );
  NAND U32988 ( .A(n24351), .B(n24352), .Z(n24326) );
  NAND U32989 ( .A(n24353), .B(n24354), .Z(n24352) );
  NANDN U32990 ( .A(n24355), .B(n24356), .Z(n24353) );
  NANDN U32991 ( .A(n24356), .B(n24355), .Z(n24351) );
  AND U32992 ( .A(n24357), .B(n24358), .Z(n24328) );
  NAND U32993 ( .A(n24359), .B(n24360), .Z(n24358) );
  OR U32994 ( .A(n24361), .B(n24362), .Z(n24359) );
  NANDN U32995 ( .A(n24363), .B(n24361), .Z(n24357) );
  NAND U32996 ( .A(n24364), .B(n24365), .Z(n24332) );
  NANDN U32997 ( .A(n24366), .B(n24367), .Z(n24365) );
  OR U32998 ( .A(n24368), .B(n24369), .Z(n24367) );
  NANDN U32999 ( .A(n24370), .B(n24368), .Z(n24364) );
  IV U33000 ( .A(n24369), .Z(n24370) );
  XNOR U33001 ( .A(n24340), .B(n24371), .Z(n24335) );
  XNOR U33002 ( .A(n24338), .B(n24341), .Z(n24371) );
  NAND U33003 ( .A(n24372), .B(n24373), .Z(n24341) );
  NAND U33004 ( .A(n24374), .B(n24375), .Z(n24373) );
  OR U33005 ( .A(n24376), .B(n24377), .Z(n24374) );
  NANDN U33006 ( .A(n24378), .B(n24376), .Z(n24372) );
  IV U33007 ( .A(n24377), .Z(n24378) );
  NAND U33008 ( .A(n24379), .B(n24380), .Z(n24338) );
  NAND U33009 ( .A(n24381), .B(n24382), .Z(n24380) );
  NANDN U33010 ( .A(n24383), .B(n24384), .Z(n24381) );
  NANDN U33011 ( .A(n24384), .B(n24383), .Z(n24379) );
  AND U33012 ( .A(n24385), .B(n24386), .Z(n24340) );
  NAND U33013 ( .A(n24387), .B(n24388), .Z(n24386) );
  OR U33014 ( .A(n24389), .B(n24390), .Z(n24387) );
  NANDN U33015 ( .A(n24391), .B(n24389), .Z(n24385) );
  XNOR U33016 ( .A(n24366), .B(n24392), .Z(N63232) );
  XOR U33017 ( .A(n24368), .B(n24369), .Z(n24392) );
  XNOR U33018 ( .A(n24382), .B(n24393), .Z(n24369) );
  XOR U33019 ( .A(n24383), .B(n24384), .Z(n24393) );
  XOR U33020 ( .A(n24389), .B(n24394), .Z(n24384) );
  XOR U33021 ( .A(n24388), .B(n24391), .Z(n24394) );
  IV U33022 ( .A(n24390), .Z(n24391) );
  NAND U33023 ( .A(n24395), .B(n24396), .Z(n24390) );
  OR U33024 ( .A(n24397), .B(n24398), .Z(n24396) );
  OR U33025 ( .A(n24399), .B(n24400), .Z(n24395) );
  NAND U33026 ( .A(n24401), .B(n24402), .Z(n24388) );
  OR U33027 ( .A(n24403), .B(n24404), .Z(n24402) );
  OR U33028 ( .A(n24405), .B(n24406), .Z(n24401) );
  NOR U33029 ( .A(n24407), .B(n24408), .Z(n24389) );
  ANDN U33030 ( .B(n24409), .A(n24410), .Z(n24383) );
  XNOR U33031 ( .A(n24376), .B(n24411), .Z(n24382) );
  XNOR U33032 ( .A(n24375), .B(n24377), .Z(n24411) );
  NAND U33033 ( .A(n24412), .B(n24413), .Z(n24377) );
  OR U33034 ( .A(n24414), .B(n24415), .Z(n24413) );
  OR U33035 ( .A(n24416), .B(n24417), .Z(n24412) );
  NAND U33036 ( .A(n24418), .B(n24419), .Z(n24375) );
  OR U33037 ( .A(n24420), .B(n24421), .Z(n24419) );
  OR U33038 ( .A(n24422), .B(n24423), .Z(n24418) );
  ANDN U33039 ( .B(n24424), .A(n24425), .Z(n24376) );
  IV U33040 ( .A(n24426), .Z(n24424) );
  ANDN U33041 ( .B(n24427), .A(n24428), .Z(n24368) );
  XOR U33042 ( .A(n24354), .B(n24429), .Z(n24366) );
  XOR U33043 ( .A(n24355), .B(n24356), .Z(n24429) );
  XOR U33044 ( .A(n24361), .B(n24430), .Z(n24356) );
  XOR U33045 ( .A(n24360), .B(n24363), .Z(n24430) );
  IV U33046 ( .A(n24362), .Z(n24363) );
  NAND U33047 ( .A(n24431), .B(n24432), .Z(n24362) );
  OR U33048 ( .A(n24433), .B(n24434), .Z(n24432) );
  OR U33049 ( .A(n24435), .B(n24436), .Z(n24431) );
  NAND U33050 ( .A(n24437), .B(n24438), .Z(n24360) );
  OR U33051 ( .A(n24439), .B(n24440), .Z(n24438) );
  OR U33052 ( .A(n24441), .B(n24442), .Z(n24437) );
  NOR U33053 ( .A(n24443), .B(n24444), .Z(n24361) );
  ANDN U33054 ( .B(n24445), .A(n24446), .Z(n24355) );
  IV U33055 ( .A(n24447), .Z(n24445) );
  XNOR U33056 ( .A(n24348), .B(n24448), .Z(n24354) );
  XNOR U33057 ( .A(n24347), .B(n24349), .Z(n24448) );
  NAND U33058 ( .A(n24449), .B(n24450), .Z(n24349) );
  OR U33059 ( .A(n24451), .B(n24452), .Z(n24450) );
  OR U33060 ( .A(n24453), .B(n24454), .Z(n24449) );
  NAND U33061 ( .A(n24455), .B(n24456), .Z(n24347) );
  OR U33062 ( .A(n24457), .B(n24458), .Z(n24456) );
  OR U33063 ( .A(n24459), .B(n24460), .Z(n24455) );
  ANDN U33064 ( .B(n24461), .A(n24462), .Z(n24348) );
  IV U33065 ( .A(n24463), .Z(n24461) );
  XNOR U33066 ( .A(n24428), .B(n24427), .Z(N63231) );
  XOR U33067 ( .A(n24447), .B(n24446), .Z(n24427) );
  XNOR U33068 ( .A(n24462), .B(n24463), .Z(n24446) );
  XNOR U33069 ( .A(n24457), .B(n24458), .Z(n24463) );
  XNOR U33070 ( .A(n24459), .B(n24460), .Z(n24458) );
  XNOR U33071 ( .A(y[4885]), .B(x[4885]), .Z(n24460) );
  XNOR U33072 ( .A(y[4886]), .B(x[4886]), .Z(n24459) );
  XNOR U33073 ( .A(y[4884]), .B(x[4884]), .Z(n24457) );
  XNOR U33074 ( .A(n24451), .B(n24452), .Z(n24462) );
  XNOR U33075 ( .A(y[4881]), .B(x[4881]), .Z(n24452) );
  XNOR U33076 ( .A(n24453), .B(n24454), .Z(n24451) );
  XNOR U33077 ( .A(y[4882]), .B(x[4882]), .Z(n24454) );
  XNOR U33078 ( .A(y[4883]), .B(x[4883]), .Z(n24453) );
  XNOR U33079 ( .A(n24444), .B(n24443), .Z(n24447) );
  XNOR U33080 ( .A(n24439), .B(n24440), .Z(n24443) );
  XNOR U33081 ( .A(y[4878]), .B(x[4878]), .Z(n24440) );
  XNOR U33082 ( .A(n24441), .B(n24442), .Z(n24439) );
  XNOR U33083 ( .A(y[4879]), .B(x[4879]), .Z(n24442) );
  XNOR U33084 ( .A(y[4880]), .B(x[4880]), .Z(n24441) );
  XNOR U33085 ( .A(n24433), .B(n24434), .Z(n24444) );
  XNOR U33086 ( .A(y[4875]), .B(x[4875]), .Z(n24434) );
  XNOR U33087 ( .A(n24435), .B(n24436), .Z(n24433) );
  XNOR U33088 ( .A(y[4876]), .B(x[4876]), .Z(n24436) );
  XNOR U33089 ( .A(y[4877]), .B(x[4877]), .Z(n24435) );
  XOR U33090 ( .A(n24409), .B(n24410), .Z(n24428) );
  XNOR U33091 ( .A(n24425), .B(n24426), .Z(n24410) );
  XNOR U33092 ( .A(n24420), .B(n24421), .Z(n24426) );
  XNOR U33093 ( .A(n24422), .B(n24423), .Z(n24421) );
  XNOR U33094 ( .A(y[4873]), .B(x[4873]), .Z(n24423) );
  XNOR U33095 ( .A(y[4874]), .B(x[4874]), .Z(n24422) );
  XNOR U33096 ( .A(y[4872]), .B(x[4872]), .Z(n24420) );
  XNOR U33097 ( .A(n24414), .B(n24415), .Z(n24425) );
  XNOR U33098 ( .A(y[4869]), .B(x[4869]), .Z(n24415) );
  XNOR U33099 ( .A(n24416), .B(n24417), .Z(n24414) );
  XNOR U33100 ( .A(y[4870]), .B(x[4870]), .Z(n24417) );
  XNOR U33101 ( .A(y[4871]), .B(x[4871]), .Z(n24416) );
  XOR U33102 ( .A(n24408), .B(n24407), .Z(n24409) );
  XNOR U33103 ( .A(n24403), .B(n24404), .Z(n24407) );
  XNOR U33104 ( .A(y[4866]), .B(x[4866]), .Z(n24404) );
  XNOR U33105 ( .A(n24405), .B(n24406), .Z(n24403) );
  XNOR U33106 ( .A(y[4867]), .B(x[4867]), .Z(n24406) );
  XNOR U33107 ( .A(y[4868]), .B(x[4868]), .Z(n24405) );
  XNOR U33108 ( .A(n24397), .B(n24398), .Z(n24408) );
  XNOR U33109 ( .A(y[4863]), .B(x[4863]), .Z(n24398) );
  XNOR U33110 ( .A(n24399), .B(n24400), .Z(n24397) );
  XNOR U33111 ( .A(y[4864]), .B(x[4864]), .Z(n24400) );
  XNOR U33112 ( .A(y[4865]), .B(x[4865]), .Z(n24399) );
  NAND U33113 ( .A(n24464), .B(n24465), .Z(N63222) );
  NANDN U33114 ( .A(n24466), .B(n24467), .Z(n24465) );
  OR U33115 ( .A(n24468), .B(n24469), .Z(n24467) );
  NAND U33116 ( .A(n24468), .B(n24469), .Z(n24464) );
  XOR U33117 ( .A(n24468), .B(n24470), .Z(N63221) );
  XNOR U33118 ( .A(n24466), .B(n24469), .Z(n24470) );
  AND U33119 ( .A(n24471), .B(n24472), .Z(n24469) );
  NANDN U33120 ( .A(n24473), .B(n24474), .Z(n24472) );
  NANDN U33121 ( .A(n24475), .B(n24476), .Z(n24474) );
  NANDN U33122 ( .A(n24476), .B(n24475), .Z(n24471) );
  NAND U33123 ( .A(n24477), .B(n24478), .Z(n24466) );
  NANDN U33124 ( .A(n24479), .B(n24480), .Z(n24478) );
  OR U33125 ( .A(n24481), .B(n24482), .Z(n24480) );
  NAND U33126 ( .A(n24482), .B(n24481), .Z(n24477) );
  AND U33127 ( .A(n24483), .B(n24484), .Z(n24468) );
  NANDN U33128 ( .A(n24485), .B(n24486), .Z(n24484) );
  NANDN U33129 ( .A(n24487), .B(n24488), .Z(n24486) );
  NANDN U33130 ( .A(n24488), .B(n24487), .Z(n24483) );
  XOR U33131 ( .A(n24482), .B(n24489), .Z(N63220) );
  XOR U33132 ( .A(n24479), .B(n24481), .Z(n24489) );
  XNOR U33133 ( .A(n24475), .B(n24490), .Z(n24481) );
  XNOR U33134 ( .A(n24473), .B(n24476), .Z(n24490) );
  NAND U33135 ( .A(n24491), .B(n24492), .Z(n24476) );
  NAND U33136 ( .A(n24493), .B(n24494), .Z(n24492) );
  OR U33137 ( .A(n24495), .B(n24496), .Z(n24493) );
  NANDN U33138 ( .A(n24497), .B(n24495), .Z(n24491) );
  IV U33139 ( .A(n24496), .Z(n24497) );
  NAND U33140 ( .A(n24498), .B(n24499), .Z(n24473) );
  NAND U33141 ( .A(n24500), .B(n24501), .Z(n24499) );
  NANDN U33142 ( .A(n24502), .B(n24503), .Z(n24500) );
  NANDN U33143 ( .A(n24503), .B(n24502), .Z(n24498) );
  AND U33144 ( .A(n24504), .B(n24505), .Z(n24475) );
  NAND U33145 ( .A(n24506), .B(n24507), .Z(n24505) );
  OR U33146 ( .A(n24508), .B(n24509), .Z(n24506) );
  NANDN U33147 ( .A(n24510), .B(n24508), .Z(n24504) );
  NAND U33148 ( .A(n24511), .B(n24512), .Z(n24479) );
  NANDN U33149 ( .A(n24513), .B(n24514), .Z(n24512) );
  OR U33150 ( .A(n24515), .B(n24516), .Z(n24514) );
  NANDN U33151 ( .A(n24517), .B(n24515), .Z(n24511) );
  IV U33152 ( .A(n24516), .Z(n24517) );
  XNOR U33153 ( .A(n24487), .B(n24518), .Z(n24482) );
  XNOR U33154 ( .A(n24485), .B(n24488), .Z(n24518) );
  NAND U33155 ( .A(n24519), .B(n24520), .Z(n24488) );
  NAND U33156 ( .A(n24521), .B(n24522), .Z(n24520) );
  OR U33157 ( .A(n24523), .B(n24524), .Z(n24521) );
  NANDN U33158 ( .A(n24525), .B(n24523), .Z(n24519) );
  IV U33159 ( .A(n24524), .Z(n24525) );
  NAND U33160 ( .A(n24526), .B(n24527), .Z(n24485) );
  NAND U33161 ( .A(n24528), .B(n24529), .Z(n24527) );
  NANDN U33162 ( .A(n24530), .B(n24531), .Z(n24528) );
  NANDN U33163 ( .A(n24531), .B(n24530), .Z(n24526) );
  AND U33164 ( .A(n24532), .B(n24533), .Z(n24487) );
  NAND U33165 ( .A(n24534), .B(n24535), .Z(n24533) );
  OR U33166 ( .A(n24536), .B(n24537), .Z(n24534) );
  NANDN U33167 ( .A(n24538), .B(n24536), .Z(n24532) );
  XNOR U33168 ( .A(n24513), .B(n24539), .Z(N63219) );
  XOR U33169 ( .A(n24515), .B(n24516), .Z(n24539) );
  XNOR U33170 ( .A(n24529), .B(n24540), .Z(n24516) );
  XOR U33171 ( .A(n24530), .B(n24531), .Z(n24540) );
  XOR U33172 ( .A(n24536), .B(n24541), .Z(n24531) );
  XOR U33173 ( .A(n24535), .B(n24538), .Z(n24541) );
  IV U33174 ( .A(n24537), .Z(n24538) );
  NAND U33175 ( .A(n24542), .B(n24543), .Z(n24537) );
  OR U33176 ( .A(n24544), .B(n24545), .Z(n24543) );
  OR U33177 ( .A(n24546), .B(n24547), .Z(n24542) );
  NAND U33178 ( .A(n24548), .B(n24549), .Z(n24535) );
  OR U33179 ( .A(n24550), .B(n24551), .Z(n24549) );
  OR U33180 ( .A(n24552), .B(n24553), .Z(n24548) );
  NOR U33181 ( .A(n24554), .B(n24555), .Z(n24536) );
  ANDN U33182 ( .B(n24556), .A(n24557), .Z(n24530) );
  XNOR U33183 ( .A(n24523), .B(n24558), .Z(n24529) );
  XNOR U33184 ( .A(n24522), .B(n24524), .Z(n24558) );
  NAND U33185 ( .A(n24559), .B(n24560), .Z(n24524) );
  OR U33186 ( .A(n24561), .B(n24562), .Z(n24560) );
  OR U33187 ( .A(n24563), .B(n24564), .Z(n24559) );
  NAND U33188 ( .A(n24565), .B(n24566), .Z(n24522) );
  OR U33189 ( .A(n24567), .B(n24568), .Z(n24566) );
  OR U33190 ( .A(n24569), .B(n24570), .Z(n24565) );
  ANDN U33191 ( .B(n24571), .A(n24572), .Z(n24523) );
  IV U33192 ( .A(n24573), .Z(n24571) );
  ANDN U33193 ( .B(n24574), .A(n24575), .Z(n24515) );
  XOR U33194 ( .A(n24501), .B(n24576), .Z(n24513) );
  XOR U33195 ( .A(n24502), .B(n24503), .Z(n24576) );
  XOR U33196 ( .A(n24508), .B(n24577), .Z(n24503) );
  XOR U33197 ( .A(n24507), .B(n24510), .Z(n24577) );
  IV U33198 ( .A(n24509), .Z(n24510) );
  NAND U33199 ( .A(n24578), .B(n24579), .Z(n24509) );
  OR U33200 ( .A(n24580), .B(n24581), .Z(n24579) );
  OR U33201 ( .A(n24582), .B(n24583), .Z(n24578) );
  NAND U33202 ( .A(n24584), .B(n24585), .Z(n24507) );
  OR U33203 ( .A(n24586), .B(n24587), .Z(n24585) );
  OR U33204 ( .A(n24588), .B(n24589), .Z(n24584) );
  NOR U33205 ( .A(n24590), .B(n24591), .Z(n24508) );
  ANDN U33206 ( .B(n24592), .A(n24593), .Z(n24502) );
  IV U33207 ( .A(n24594), .Z(n24592) );
  XNOR U33208 ( .A(n24495), .B(n24595), .Z(n24501) );
  XNOR U33209 ( .A(n24494), .B(n24496), .Z(n24595) );
  NAND U33210 ( .A(n24596), .B(n24597), .Z(n24496) );
  OR U33211 ( .A(n24598), .B(n24599), .Z(n24597) );
  OR U33212 ( .A(n24600), .B(n24601), .Z(n24596) );
  NAND U33213 ( .A(n24602), .B(n24603), .Z(n24494) );
  OR U33214 ( .A(n24604), .B(n24605), .Z(n24603) );
  OR U33215 ( .A(n24606), .B(n24607), .Z(n24602) );
  ANDN U33216 ( .B(n24608), .A(n24609), .Z(n24495) );
  IV U33217 ( .A(n24610), .Z(n24608) );
  XNOR U33218 ( .A(n24575), .B(n24574), .Z(N63218) );
  XOR U33219 ( .A(n24594), .B(n24593), .Z(n24574) );
  XNOR U33220 ( .A(n24609), .B(n24610), .Z(n24593) );
  XNOR U33221 ( .A(n24604), .B(n24605), .Z(n24610) );
  XNOR U33222 ( .A(n24606), .B(n24607), .Z(n24605) );
  XNOR U33223 ( .A(y[4861]), .B(x[4861]), .Z(n24607) );
  XNOR U33224 ( .A(y[4862]), .B(x[4862]), .Z(n24606) );
  XNOR U33225 ( .A(y[4860]), .B(x[4860]), .Z(n24604) );
  XNOR U33226 ( .A(n24598), .B(n24599), .Z(n24609) );
  XNOR U33227 ( .A(y[4857]), .B(x[4857]), .Z(n24599) );
  XNOR U33228 ( .A(n24600), .B(n24601), .Z(n24598) );
  XNOR U33229 ( .A(y[4858]), .B(x[4858]), .Z(n24601) );
  XNOR U33230 ( .A(y[4859]), .B(x[4859]), .Z(n24600) );
  XNOR U33231 ( .A(n24591), .B(n24590), .Z(n24594) );
  XNOR U33232 ( .A(n24586), .B(n24587), .Z(n24590) );
  XNOR U33233 ( .A(y[4854]), .B(x[4854]), .Z(n24587) );
  XNOR U33234 ( .A(n24588), .B(n24589), .Z(n24586) );
  XNOR U33235 ( .A(y[4855]), .B(x[4855]), .Z(n24589) );
  XNOR U33236 ( .A(y[4856]), .B(x[4856]), .Z(n24588) );
  XNOR U33237 ( .A(n24580), .B(n24581), .Z(n24591) );
  XNOR U33238 ( .A(y[4851]), .B(x[4851]), .Z(n24581) );
  XNOR U33239 ( .A(n24582), .B(n24583), .Z(n24580) );
  XNOR U33240 ( .A(y[4852]), .B(x[4852]), .Z(n24583) );
  XNOR U33241 ( .A(y[4853]), .B(x[4853]), .Z(n24582) );
  XOR U33242 ( .A(n24556), .B(n24557), .Z(n24575) );
  XNOR U33243 ( .A(n24572), .B(n24573), .Z(n24557) );
  XNOR U33244 ( .A(n24567), .B(n24568), .Z(n24573) );
  XNOR U33245 ( .A(n24569), .B(n24570), .Z(n24568) );
  XNOR U33246 ( .A(y[4849]), .B(x[4849]), .Z(n24570) );
  XNOR U33247 ( .A(y[4850]), .B(x[4850]), .Z(n24569) );
  XNOR U33248 ( .A(y[4848]), .B(x[4848]), .Z(n24567) );
  XNOR U33249 ( .A(n24561), .B(n24562), .Z(n24572) );
  XNOR U33250 ( .A(y[4845]), .B(x[4845]), .Z(n24562) );
  XNOR U33251 ( .A(n24563), .B(n24564), .Z(n24561) );
  XNOR U33252 ( .A(y[4846]), .B(x[4846]), .Z(n24564) );
  XNOR U33253 ( .A(y[4847]), .B(x[4847]), .Z(n24563) );
  XOR U33254 ( .A(n24555), .B(n24554), .Z(n24556) );
  XNOR U33255 ( .A(n24550), .B(n24551), .Z(n24554) );
  XNOR U33256 ( .A(y[4842]), .B(x[4842]), .Z(n24551) );
  XNOR U33257 ( .A(n24552), .B(n24553), .Z(n24550) );
  XNOR U33258 ( .A(y[4843]), .B(x[4843]), .Z(n24553) );
  XNOR U33259 ( .A(y[4844]), .B(x[4844]), .Z(n24552) );
  XNOR U33260 ( .A(n24544), .B(n24545), .Z(n24555) );
  XNOR U33261 ( .A(y[4839]), .B(x[4839]), .Z(n24545) );
  XNOR U33262 ( .A(n24546), .B(n24547), .Z(n24544) );
  XNOR U33263 ( .A(y[4840]), .B(x[4840]), .Z(n24547) );
  XNOR U33264 ( .A(y[4841]), .B(x[4841]), .Z(n24546) );
  NAND U33265 ( .A(n24611), .B(n24612), .Z(N63209) );
  NANDN U33266 ( .A(n24613), .B(n24614), .Z(n24612) );
  OR U33267 ( .A(n24615), .B(n24616), .Z(n24614) );
  NAND U33268 ( .A(n24615), .B(n24616), .Z(n24611) );
  XOR U33269 ( .A(n24615), .B(n24617), .Z(N63208) );
  XNOR U33270 ( .A(n24613), .B(n24616), .Z(n24617) );
  AND U33271 ( .A(n24618), .B(n24619), .Z(n24616) );
  NANDN U33272 ( .A(n24620), .B(n24621), .Z(n24619) );
  NANDN U33273 ( .A(n24622), .B(n24623), .Z(n24621) );
  NANDN U33274 ( .A(n24623), .B(n24622), .Z(n24618) );
  NAND U33275 ( .A(n24624), .B(n24625), .Z(n24613) );
  NANDN U33276 ( .A(n24626), .B(n24627), .Z(n24625) );
  OR U33277 ( .A(n24628), .B(n24629), .Z(n24627) );
  NAND U33278 ( .A(n24629), .B(n24628), .Z(n24624) );
  AND U33279 ( .A(n24630), .B(n24631), .Z(n24615) );
  NANDN U33280 ( .A(n24632), .B(n24633), .Z(n24631) );
  NANDN U33281 ( .A(n24634), .B(n24635), .Z(n24633) );
  NANDN U33282 ( .A(n24635), .B(n24634), .Z(n24630) );
  XOR U33283 ( .A(n24629), .B(n24636), .Z(N63207) );
  XOR U33284 ( .A(n24626), .B(n24628), .Z(n24636) );
  XNOR U33285 ( .A(n24622), .B(n24637), .Z(n24628) );
  XNOR U33286 ( .A(n24620), .B(n24623), .Z(n24637) );
  NAND U33287 ( .A(n24638), .B(n24639), .Z(n24623) );
  NAND U33288 ( .A(n24640), .B(n24641), .Z(n24639) );
  OR U33289 ( .A(n24642), .B(n24643), .Z(n24640) );
  NANDN U33290 ( .A(n24644), .B(n24642), .Z(n24638) );
  IV U33291 ( .A(n24643), .Z(n24644) );
  NAND U33292 ( .A(n24645), .B(n24646), .Z(n24620) );
  NAND U33293 ( .A(n24647), .B(n24648), .Z(n24646) );
  NANDN U33294 ( .A(n24649), .B(n24650), .Z(n24647) );
  NANDN U33295 ( .A(n24650), .B(n24649), .Z(n24645) );
  AND U33296 ( .A(n24651), .B(n24652), .Z(n24622) );
  NAND U33297 ( .A(n24653), .B(n24654), .Z(n24652) );
  OR U33298 ( .A(n24655), .B(n24656), .Z(n24653) );
  NANDN U33299 ( .A(n24657), .B(n24655), .Z(n24651) );
  NAND U33300 ( .A(n24658), .B(n24659), .Z(n24626) );
  NANDN U33301 ( .A(n24660), .B(n24661), .Z(n24659) );
  OR U33302 ( .A(n24662), .B(n24663), .Z(n24661) );
  NANDN U33303 ( .A(n24664), .B(n24662), .Z(n24658) );
  IV U33304 ( .A(n24663), .Z(n24664) );
  XNOR U33305 ( .A(n24634), .B(n24665), .Z(n24629) );
  XNOR U33306 ( .A(n24632), .B(n24635), .Z(n24665) );
  NAND U33307 ( .A(n24666), .B(n24667), .Z(n24635) );
  NAND U33308 ( .A(n24668), .B(n24669), .Z(n24667) );
  OR U33309 ( .A(n24670), .B(n24671), .Z(n24668) );
  NANDN U33310 ( .A(n24672), .B(n24670), .Z(n24666) );
  IV U33311 ( .A(n24671), .Z(n24672) );
  NAND U33312 ( .A(n24673), .B(n24674), .Z(n24632) );
  NAND U33313 ( .A(n24675), .B(n24676), .Z(n24674) );
  NANDN U33314 ( .A(n24677), .B(n24678), .Z(n24675) );
  NANDN U33315 ( .A(n24678), .B(n24677), .Z(n24673) );
  AND U33316 ( .A(n24679), .B(n24680), .Z(n24634) );
  NAND U33317 ( .A(n24681), .B(n24682), .Z(n24680) );
  OR U33318 ( .A(n24683), .B(n24684), .Z(n24681) );
  NANDN U33319 ( .A(n24685), .B(n24683), .Z(n24679) );
  XNOR U33320 ( .A(n24660), .B(n24686), .Z(N63206) );
  XOR U33321 ( .A(n24662), .B(n24663), .Z(n24686) );
  XNOR U33322 ( .A(n24676), .B(n24687), .Z(n24663) );
  XOR U33323 ( .A(n24677), .B(n24678), .Z(n24687) );
  XOR U33324 ( .A(n24683), .B(n24688), .Z(n24678) );
  XOR U33325 ( .A(n24682), .B(n24685), .Z(n24688) );
  IV U33326 ( .A(n24684), .Z(n24685) );
  NAND U33327 ( .A(n24689), .B(n24690), .Z(n24684) );
  OR U33328 ( .A(n24691), .B(n24692), .Z(n24690) );
  OR U33329 ( .A(n24693), .B(n24694), .Z(n24689) );
  NAND U33330 ( .A(n24695), .B(n24696), .Z(n24682) );
  OR U33331 ( .A(n24697), .B(n24698), .Z(n24696) );
  OR U33332 ( .A(n24699), .B(n24700), .Z(n24695) );
  NOR U33333 ( .A(n24701), .B(n24702), .Z(n24683) );
  ANDN U33334 ( .B(n24703), .A(n24704), .Z(n24677) );
  XNOR U33335 ( .A(n24670), .B(n24705), .Z(n24676) );
  XNOR U33336 ( .A(n24669), .B(n24671), .Z(n24705) );
  NAND U33337 ( .A(n24706), .B(n24707), .Z(n24671) );
  OR U33338 ( .A(n24708), .B(n24709), .Z(n24707) );
  OR U33339 ( .A(n24710), .B(n24711), .Z(n24706) );
  NAND U33340 ( .A(n24712), .B(n24713), .Z(n24669) );
  OR U33341 ( .A(n24714), .B(n24715), .Z(n24713) );
  OR U33342 ( .A(n24716), .B(n24717), .Z(n24712) );
  ANDN U33343 ( .B(n24718), .A(n24719), .Z(n24670) );
  IV U33344 ( .A(n24720), .Z(n24718) );
  ANDN U33345 ( .B(n24721), .A(n24722), .Z(n24662) );
  XOR U33346 ( .A(n24648), .B(n24723), .Z(n24660) );
  XOR U33347 ( .A(n24649), .B(n24650), .Z(n24723) );
  XOR U33348 ( .A(n24655), .B(n24724), .Z(n24650) );
  XOR U33349 ( .A(n24654), .B(n24657), .Z(n24724) );
  IV U33350 ( .A(n24656), .Z(n24657) );
  NAND U33351 ( .A(n24725), .B(n24726), .Z(n24656) );
  OR U33352 ( .A(n24727), .B(n24728), .Z(n24726) );
  OR U33353 ( .A(n24729), .B(n24730), .Z(n24725) );
  NAND U33354 ( .A(n24731), .B(n24732), .Z(n24654) );
  OR U33355 ( .A(n24733), .B(n24734), .Z(n24732) );
  OR U33356 ( .A(n24735), .B(n24736), .Z(n24731) );
  NOR U33357 ( .A(n24737), .B(n24738), .Z(n24655) );
  ANDN U33358 ( .B(n24739), .A(n24740), .Z(n24649) );
  IV U33359 ( .A(n24741), .Z(n24739) );
  XNOR U33360 ( .A(n24642), .B(n24742), .Z(n24648) );
  XNOR U33361 ( .A(n24641), .B(n24643), .Z(n24742) );
  NAND U33362 ( .A(n24743), .B(n24744), .Z(n24643) );
  OR U33363 ( .A(n24745), .B(n24746), .Z(n24744) );
  OR U33364 ( .A(n24747), .B(n24748), .Z(n24743) );
  NAND U33365 ( .A(n24749), .B(n24750), .Z(n24641) );
  OR U33366 ( .A(n24751), .B(n24752), .Z(n24750) );
  OR U33367 ( .A(n24753), .B(n24754), .Z(n24749) );
  ANDN U33368 ( .B(n24755), .A(n24756), .Z(n24642) );
  IV U33369 ( .A(n24757), .Z(n24755) );
  XNOR U33370 ( .A(n24722), .B(n24721), .Z(N63205) );
  XOR U33371 ( .A(n24741), .B(n24740), .Z(n24721) );
  XNOR U33372 ( .A(n24756), .B(n24757), .Z(n24740) );
  XNOR U33373 ( .A(n24751), .B(n24752), .Z(n24757) );
  XNOR U33374 ( .A(n24753), .B(n24754), .Z(n24752) );
  XNOR U33375 ( .A(y[4837]), .B(x[4837]), .Z(n24754) );
  XNOR U33376 ( .A(y[4838]), .B(x[4838]), .Z(n24753) );
  XNOR U33377 ( .A(y[4836]), .B(x[4836]), .Z(n24751) );
  XNOR U33378 ( .A(n24745), .B(n24746), .Z(n24756) );
  XNOR U33379 ( .A(y[4833]), .B(x[4833]), .Z(n24746) );
  XNOR U33380 ( .A(n24747), .B(n24748), .Z(n24745) );
  XNOR U33381 ( .A(y[4834]), .B(x[4834]), .Z(n24748) );
  XNOR U33382 ( .A(y[4835]), .B(x[4835]), .Z(n24747) );
  XNOR U33383 ( .A(n24738), .B(n24737), .Z(n24741) );
  XNOR U33384 ( .A(n24733), .B(n24734), .Z(n24737) );
  XNOR U33385 ( .A(y[4830]), .B(x[4830]), .Z(n24734) );
  XNOR U33386 ( .A(n24735), .B(n24736), .Z(n24733) );
  XNOR U33387 ( .A(y[4831]), .B(x[4831]), .Z(n24736) );
  XNOR U33388 ( .A(y[4832]), .B(x[4832]), .Z(n24735) );
  XNOR U33389 ( .A(n24727), .B(n24728), .Z(n24738) );
  XNOR U33390 ( .A(y[4827]), .B(x[4827]), .Z(n24728) );
  XNOR U33391 ( .A(n24729), .B(n24730), .Z(n24727) );
  XNOR U33392 ( .A(y[4828]), .B(x[4828]), .Z(n24730) );
  XNOR U33393 ( .A(y[4829]), .B(x[4829]), .Z(n24729) );
  XOR U33394 ( .A(n24703), .B(n24704), .Z(n24722) );
  XNOR U33395 ( .A(n24719), .B(n24720), .Z(n24704) );
  XNOR U33396 ( .A(n24714), .B(n24715), .Z(n24720) );
  XNOR U33397 ( .A(n24716), .B(n24717), .Z(n24715) );
  XNOR U33398 ( .A(y[4825]), .B(x[4825]), .Z(n24717) );
  XNOR U33399 ( .A(y[4826]), .B(x[4826]), .Z(n24716) );
  XNOR U33400 ( .A(y[4824]), .B(x[4824]), .Z(n24714) );
  XNOR U33401 ( .A(n24708), .B(n24709), .Z(n24719) );
  XNOR U33402 ( .A(y[4821]), .B(x[4821]), .Z(n24709) );
  XNOR U33403 ( .A(n24710), .B(n24711), .Z(n24708) );
  XNOR U33404 ( .A(y[4822]), .B(x[4822]), .Z(n24711) );
  XNOR U33405 ( .A(y[4823]), .B(x[4823]), .Z(n24710) );
  XOR U33406 ( .A(n24702), .B(n24701), .Z(n24703) );
  XNOR U33407 ( .A(n24697), .B(n24698), .Z(n24701) );
  XNOR U33408 ( .A(y[4818]), .B(x[4818]), .Z(n24698) );
  XNOR U33409 ( .A(n24699), .B(n24700), .Z(n24697) );
  XNOR U33410 ( .A(y[4819]), .B(x[4819]), .Z(n24700) );
  XNOR U33411 ( .A(y[4820]), .B(x[4820]), .Z(n24699) );
  XNOR U33412 ( .A(n24691), .B(n24692), .Z(n24702) );
  XNOR U33413 ( .A(y[4815]), .B(x[4815]), .Z(n24692) );
  XNOR U33414 ( .A(n24693), .B(n24694), .Z(n24691) );
  XNOR U33415 ( .A(y[4816]), .B(x[4816]), .Z(n24694) );
  XNOR U33416 ( .A(y[4817]), .B(x[4817]), .Z(n24693) );
  NAND U33417 ( .A(n24758), .B(n24759), .Z(N63196) );
  NANDN U33418 ( .A(n24760), .B(n24761), .Z(n24759) );
  OR U33419 ( .A(n24762), .B(n24763), .Z(n24761) );
  NAND U33420 ( .A(n24762), .B(n24763), .Z(n24758) );
  XOR U33421 ( .A(n24762), .B(n24764), .Z(N63195) );
  XNOR U33422 ( .A(n24760), .B(n24763), .Z(n24764) );
  AND U33423 ( .A(n24765), .B(n24766), .Z(n24763) );
  NANDN U33424 ( .A(n24767), .B(n24768), .Z(n24766) );
  NANDN U33425 ( .A(n24769), .B(n24770), .Z(n24768) );
  NANDN U33426 ( .A(n24770), .B(n24769), .Z(n24765) );
  NAND U33427 ( .A(n24771), .B(n24772), .Z(n24760) );
  NANDN U33428 ( .A(n24773), .B(n24774), .Z(n24772) );
  OR U33429 ( .A(n24775), .B(n24776), .Z(n24774) );
  NAND U33430 ( .A(n24776), .B(n24775), .Z(n24771) );
  AND U33431 ( .A(n24777), .B(n24778), .Z(n24762) );
  NANDN U33432 ( .A(n24779), .B(n24780), .Z(n24778) );
  NANDN U33433 ( .A(n24781), .B(n24782), .Z(n24780) );
  NANDN U33434 ( .A(n24782), .B(n24781), .Z(n24777) );
  XOR U33435 ( .A(n24776), .B(n24783), .Z(N63194) );
  XOR U33436 ( .A(n24773), .B(n24775), .Z(n24783) );
  XNOR U33437 ( .A(n24769), .B(n24784), .Z(n24775) );
  XNOR U33438 ( .A(n24767), .B(n24770), .Z(n24784) );
  NAND U33439 ( .A(n24785), .B(n24786), .Z(n24770) );
  NAND U33440 ( .A(n24787), .B(n24788), .Z(n24786) );
  OR U33441 ( .A(n24789), .B(n24790), .Z(n24787) );
  NANDN U33442 ( .A(n24791), .B(n24789), .Z(n24785) );
  IV U33443 ( .A(n24790), .Z(n24791) );
  NAND U33444 ( .A(n24792), .B(n24793), .Z(n24767) );
  NAND U33445 ( .A(n24794), .B(n24795), .Z(n24793) );
  NANDN U33446 ( .A(n24796), .B(n24797), .Z(n24794) );
  NANDN U33447 ( .A(n24797), .B(n24796), .Z(n24792) );
  AND U33448 ( .A(n24798), .B(n24799), .Z(n24769) );
  NAND U33449 ( .A(n24800), .B(n24801), .Z(n24799) );
  OR U33450 ( .A(n24802), .B(n24803), .Z(n24800) );
  NANDN U33451 ( .A(n24804), .B(n24802), .Z(n24798) );
  NAND U33452 ( .A(n24805), .B(n24806), .Z(n24773) );
  NANDN U33453 ( .A(n24807), .B(n24808), .Z(n24806) );
  OR U33454 ( .A(n24809), .B(n24810), .Z(n24808) );
  NANDN U33455 ( .A(n24811), .B(n24809), .Z(n24805) );
  IV U33456 ( .A(n24810), .Z(n24811) );
  XNOR U33457 ( .A(n24781), .B(n24812), .Z(n24776) );
  XNOR U33458 ( .A(n24779), .B(n24782), .Z(n24812) );
  NAND U33459 ( .A(n24813), .B(n24814), .Z(n24782) );
  NAND U33460 ( .A(n24815), .B(n24816), .Z(n24814) );
  OR U33461 ( .A(n24817), .B(n24818), .Z(n24815) );
  NANDN U33462 ( .A(n24819), .B(n24817), .Z(n24813) );
  IV U33463 ( .A(n24818), .Z(n24819) );
  NAND U33464 ( .A(n24820), .B(n24821), .Z(n24779) );
  NAND U33465 ( .A(n24822), .B(n24823), .Z(n24821) );
  NANDN U33466 ( .A(n24824), .B(n24825), .Z(n24822) );
  NANDN U33467 ( .A(n24825), .B(n24824), .Z(n24820) );
  AND U33468 ( .A(n24826), .B(n24827), .Z(n24781) );
  NAND U33469 ( .A(n24828), .B(n24829), .Z(n24827) );
  OR U33470 ( .A(n24830), .B(n24831), .Z(n24828) );
  NANDN U33471 ( .A(n24832), .B(n24830), .Z(n24826) );
  XNOR U33472 ( .A(n24807), .B(n24833), .Z(N63193) );
  XOR U33473 ( .A(n24809), .B(n24810), .Z(n24833) );
  XNOR U33474 ( .A(n24823), .B(n24834), .Z(n24810) );
  XOR U33475 ( .A(n24824), .B(n24825), .Z(n24834) );
  XOR U33476 ( .A(n24830), .B(n24835), .Z(n24825) );
  XOR U33477 ( .A(n24829), .B(n24832), .Z(n24835) );
  IV U33478 ( .A(n24831), .Z(n24832) );
  NAND U33479 ( .A(n24836), .B(n24837), .Z(n24831) );
  OR U33480 ( .A(n24838), .B(n24839), .Z(n24837) );
  OR U33481 ( .A(n24840), .B(n24841), .Z(n24836) );
  NAND U33482 ( .A(n24842), .B(n24843), .Z(n24829) );
  OR U33483 ( .A(n24844), .B(n24845), .Z(n24843) );
  OR U33484 ( .A(n24846), .B(n24847), .Z(n24842) );
  NOR U33485 ( .A(n24848), .B(n24849), .Z(n24830) );
  ANDN U33486 ( .B(n24850), .A(n24851), .Z(n24824) );
  XNOR U33487 ( .A(n24817), .B(n24852), .Z(n24823) );
  XNOR U33488 ( .A(n24816), .B(n24818), .Z(n24852) );
  NAND U33489 ( .A(n24853), .B(n24854), .Z(n24818) );
  OR U33490 ( .A(n24855), .B(n24856), .Z(n24854) );
  OR U33491 ( .A(n24857), .B(n24858), .Z(n24853) );
  NAND U33492 ( .A(n24859), .B(n24860), .Z(n24816) );
  OR U33493 ( .A(n24861), .B(n24862), .Z(n24860) );
  OR U33494 ( .A(n24863), .B(n24864), .Z(n24859) );
  ANDN U33495 ( .B(n24865), .A(n24866), .Z(n24817) );
  IV U33496 ( .A(n24867), .Z(n24865) );
  ANDN U33497 ( .B(n24868), .A(n24869), .Z(n24809) );
  XOR U33498 ( .A(n24795), .B(n24870), .Z(n24807) );
  XOR U33499 ( .A(n24796), .B(n24797), .Z(n24870) );
  XOR U33500 ( .A(n24802), .B(n24871), .Z(n24797) );
  XOR U33501 ( .A(n24801), .B(n24804), .Z(n24871) );
  IV U33502 ( .A(n24803), .Z(n24804) );
  NAND U33503 ( .A(n24872), .B(n24873), .Z(n24803) );
  OR U33504 ( .A(n24874), .B(n24875), .Z(n24873) );
  OR U33505 ( .A(n24876), .B(n24877), .Z(n24872) );
  NAND U33506 ( .A(n24878), .B(n24879), .Z(n24801) );
  OR U33507 ( .A(n24880), .B(n24881), .Z(n24879) );
  OR U33508 ( .A(n24882), .B(n24883), .Z(n24878) );
  NOR U33509 ( .A(n24884), .B(n24885), .Z(n24802) );
  ANDN U33510 ( .B(n24886), .A(n24887), .Z(n24796) );
  IV U33511 ( .A(n24888), .Z(n24886) );
  XNOR U33512 ( .A(n24789), .B(n24889), .Z(n24795) );
  XNOR U33513 ( .A(n24788), .B(n24790), .Z(n24889) );
  NAND U33514 ( .A(n24890), .B(n24891), .Z(n24790) );
  OR U33515 ( .A(n24892), .B(n24893), .Z(n24891) );
  OR U33516 ( .A(n24894), .B(n24895), .Z(n24890) );
  NAND U33517 ( .A(n24896), .B(n24897), .Z(n24788) );
  OR U33518 ( .A(n24898), .B(n24899), .Z(n24897) );
  OR U33519 ( .A(n24900), .B(n24901), .Z(n24896) );
  ANDN U33520 ( .B(n24902), .A(n24903), .Z(n24789) );
  IV U33521 ( .A(n24904), .Z(n24902) );
  XNOR U33522 ( .A(n24869), .B(n24868), .Z(N63192) );
  XOR U33523 ( .A(n24888), .B(n24887), .Z(n24868) );
  XNOR U33524 ( .A(n24903), .B(n24904), .Z(n24887) );
  XNOR U33525 ( .A(n24898), .B(n24899), .Z(n24904) );
  XNOR U33526 ( .A(n24900), .B(n24901), .Z(n24899) );
  XNOR U33527 ( .A(y[4813]), .B(x[4813]), .Z(n24901) );
  XNOR U33528 ( .A(y[4814]), .B(x[4814]), .Z(n24900) );
  XNOR U33529 ( .A(y[4812]), .B(x[4812]), .Z(n24898) );
  XNOR U33530 ( .A(n24892), .B(n24893), .Z(n24903) );
  XNOR U33531 ( .A(y[4809]), .B(x[4809]), .Z(n24893) );
  XNOR U33532 ( .A(n24894), .B(n24895), .Z(n24892) );
  XNOR U33533 ( .A(y[4810]), .B(x[4810]), .Z(n24895) );
  XNOR U33534 ( .A(y[4811]), .B(x[4811]), .Z(n24894) );
  XNOR U33535 ( .A(n24885), .B(n24884), .Z(n24888) );
  XNOR U33536 ( .A(n24880), .B(n24881), .Z(n24884) );
  XNOR U33537 ( .A(y[4806]), .B(x[4806]), .Z(n24881) );
  XNOR U33538 ( .A(n24882), .B(n24883), .Z(n24880) );
  XNOR U33539 ( .A(y[4807]), .B(x[4807]), .Z(n24883) );
  XNOR U33540 ( .A(y[4808]), .B(x[4808]), .Z(n24882) );
  XNOR U33541 ( .A(n24874), .B(n24875), .Z(n24885) );
  XNOR U33542 ( .A(y[4803]), .B(x[4803]), .Z(n24875) );
  XNOR U33543 ( .A(n24876), .B(n24877), .Z(n24874) );
  XNOR U33544 ( .A(y[4804]), .B(x[4804]), .Z(n24877) );
  XNOR U33545 ( .A(y[4805]), .B(x[4805]), .Z(n24876) );
  XOR U33546 ( .A(n24850), .B(n24851), .Z(n24869) );
  XNOR U33547 ( .A(n24866), .B(n24867), .Z(n24851) );
  XNOR U33548 ( .A(n24861), .B(n24862), .Z(n24867) );
  XNOR U33549 ( .A(n24863), .B(n24864), .Z(n24862) );
  XNOR U33550 ( .A(y[4801]), .B(x[4801]), .Z(n24864) );
  XNOR U33551 ( .A(y[4802]), .B(x[4802]), .Z(n24863) );
  XNOR U33552 ( .A(y[4800]), .B(x[4800]), .Z(n24861) );
  XNOR U33553 ( .A(n24855), .B(n24856), .Z(n24866) );
  XNOR U33554 ( .A(y[4797]), .B(x[4797]), .Z(n24856) );
  XNOR U33555 ( .A(n24857), .B(n24858), .Z(n24855) );
  XNOR U33556 ( .A(y[4798]), .B(x[4798]), .Z(n24858) );
  XNOR U33557 ( .A(y[4799]), .B(x[4799]), .Z(n24857) );
  XOR U33558 ( .A(n24849), .B(n24848), .Z(n24850) );
  XNOR U33559 ( .A(n24844), .B(n24845), .Z(n24848) );
  XNOR U33560 ( .A(y[4794]), .B(x[4794]), .Z(n24845) );
  XNOR U33561 ( .A(n24846), .B(n24847), .Z(n24844) );
  XNOR U33562 ( .A(y[4795]), .B(x[4795]), .Z(n24847) );
  XNOR U33563 ( .A(y[4796]), .B(x[4796]), .Z(n24846) );
  XNOR U33564 ( .A(n24838), .B(n24839), .Z(n24849) );
  XNOR U33565 ( .A(y[4791]), .B(x[4791]), .Z(n24839) );
  XNOR U33566 ( .A(n24840), .B(n24841), .Z(n24838) );
  XNOR U33567 ( .A(y[4792]), .B(x[4792]), .Z(n24841) );
  XNOR U33568 ( .A(y[4793]), .B(x[4793]), .Z(n24840) );
  NAND U33569 ( .A(n24905), .B(n24906), .Z(N63183) );
  NANDN U33570 ( .A(n24907), .B(n24908), .Z(n24906) );
  OR U33571 ( .A(n24909), .B(n24910), .Z(n24908) );
  NAND U33572 ( .A(n24909), .B(n24910), .Z(n24905) );
  XOR U33573 ( .A(n24909), .B(n24911), .Z(N63182) );
  XNOR U33574 ( .A(n24907), .B(n24910), .Z(n24911) );
  AND U33575 ( .A(n24912), .B(n24913), .Z(n24910) );
  NANDN U33576 ( .A(n24914), .B(n24915), .Z(n24913) );
  NANDN U33577 ( .A(n24916), .B(n24917), .Z(n24915) );
  NANDN U33578 ( .A(n24917), .B(n24916), .Z(n24912) );
  NAND U33579 ( .A(n24918), .B(n24919), .Z(n24907) );
  NANDN U33580 ( .A(n24920), .B(n24921), .Z(n24919) );
  OR U33581 ( .A(n24922), .B(n24923), .Z(n24921) );
  NAND U33582 ( .A(n24923), .B(n24922), .Z(n24918) );
  AND U33583 ( .A(n24924), .B(n24925), .Z(n24909) );
  NANDN U33584 ( .A(n24926), .B(n24927), .Z(n24925) );
  NANDN U33585 ( .A(n24928), .B(n24929), .Z(n24927) );
  NANDN U33586 ( .A(n24929), .B(n24928), .Z(n24924) );
  XOR U33587 ( .A(n24923), .B(n24930), .Z(N63181) );
  XOR U33588 ( .A(n24920), .B(n24922), .Z(n24930) );
  XNOR U33589 ( .A(n24916), .B(n24931), .Z(n24922) );
  XNOR U33590 ( .A(n24914), .B(n24917), .Z(n24931) );
  NAND U33591 ( .A(n24932), .B(n24933), .Z(n24917) );
  NAND U33592 ( .A(n24934), .B(n24935), .Z(n24933) );
  OR U33593 ( .A(n24936), .B(n24937), .Z(n24934) );
  NANDN U33594 ( .A(n24938), .B(n24936), .Z(n24932) );
  IV U33595 ( .A(n24937), .Z(n24938) );
  NAND U33596 ( .A(n24939), .B(n24940), .Z(n24914) );
  NAND U33597 ( .A(n24941), .B(n24942), .Z(n24940) );
  NANDN U33598 ( .A(n24943), .B(n24944), .Z(n24941) );
  NANDN U33599 ( .A(n24944), .B(n24943), .Z(n24939) );
  AND U33600 ( .A(n24945), .B(n24946), .Z(n24916) );
  NAND U33601 ( .A(n24947), .B(n24948), .Z(n24946) );
  OR U33602 ( .A(n24949), .B(n24950), .Z(n24947) );
  NANDN U33603 ( .A(n24951), .B(n24949), .Z(n24945) );
  NAND U33604 ( .A(n24952), .B(n24953), .Z(n24920) );
  NANDN U33605 ( .A(n24954), .B(n24955), .Z(n24953) );
  OR U33606 ( .A(n24956), .B(n24957), .Z(n24955) );
  NANDN U33607 ( .A(n24958), .B(n24956), .Z(n24952) );
  IV U33608 ( .A(n24957), .Z(n24958) );
  XNOR U33609 ( .A(n24928), .B(n24959), .Z(n24923) );
  XNOR U33610 ( .A(n24926), .B(n24929), .Z(n24959) );
  NAND U33611 ( .A(n24960), .B(n24961), .Z(n24929) );
  NAND U33612 ( .A(n24962), .B(n24963), .Z(n24961) );
  OR U33613 ( .A(n24964), .B(n24965), .Z(n24962) );
  NANDN U33614 ( .A(n24966), .B(n24964), .Z(n24960) );
  IV U33615 ( .A(n24965), .Z(n24966) );
  NAND U33616 ( .A(n24967), .B(n24968), .Z(n24926) );
  NAND U33617 ( .A(n24969), .B(n24970), .Z(n24968) );
  NANDN U33618 ( .A(n24971), .B(n24972), .Z(n24969) );
  NANDN U33619 ( .A(n24972), .B(n24971), .Z(n24967) );
  AND U33620 ( .A(n24973), .B(n24974), .Z(n24928) );
  NAND U33621 ( .A(n24975), .B(n24976), .Z(n24974) );
  OR U33622 ( .A(n24977), .B(n24978), .Z(n24975) );
  NANDN U33623 ( .A(n24979), .B(n24977), .Z(n24973) );
  XNOR U33624 ( .A(n24954), .B(n24980), .Z(N63180) );
  XOR U33625 ( .A(n24956), .B(n24957), .Z(n24980) );
  XNOR U33626 ( .A(n24970), .B(n24981), .Z(n24957) );
  XOR U33627 ( .A(n24971), .B(n24972), .Z(n24981) );
  XOR U33628 ( .A(n24977), .B(n24982), .Z(n24972) );
  XOR U33629 ( .A(n24976), .B(n24979), .Z(n24982) );
  IV U33630 ( .A(n24978), .Z(n24979) );
  NAND U33631 ( .A(n24983), .B(n24984), .Z(n24978) );
  OR U33632 ( .A(n24985), .B(n24986), .Z(n24984) );
  OR U33633 ( .A(n24987), .B(n24988), .Z(n24983) );
  NAND U33634 ( .A(n24989), .B(n24990), .Z(n24976) );
  OR U33635 ( .A(n24991), .B(n24992), .Z(n24990) );
  OR U33636 ( .A(n24993), .B(n24994), .Z(n24989) );
  NOR U33637 ( .A(n24995), .B(n24996), .Z(n24977) );
  ANDN U33638 ( .B(n24997), .A(n24998), .Z(n24971) );
  XNOR U33639 ( .A(n24964), .B(n24999), .Z(n24970) );
  XNOR U33640 ( .A(n24963), .B(n24965), .Z(n24999) );
  NAND U33641 ( .A(n25000), .B(n25001), .Z(n24965) );
  OR U33642 ( .A(n25002), .B(n25003), .Z(n25001) );
  OR U33643 ( .A(n25004), .B(n25005), .Z(n25000) );
  NAND U33644 ( .A(n25006), .B(n25007), .Z(n24963) );
  OR U33645 ( .A(n25008), .B(n25009), .Z(n25007) );
  OR U33646 ( .A(n25010), .B(n25011), .Z(n25006) );
  ANDN U33647 ( .B(n25012), .A(n25013), .Z(n24964) );
  IV U33648 ( .A(n25014), .Z(n25012) );
  ANDN U33649 ( .B(n25015), .A(n25016), .Z(n24956) );
  XOR U33650 ( .A(n24942), .B(n25017), .Z(n24954) );
  XOR U33651 ( .A(n24943), .B(n24944), .Z(n25017) );
  XOR U33652 ( .A(n24949), .B(n25018), .Z(n24944) );
  XOR U33653 ( .A(n24948), .B(n24951), .Z(n25018) );
  IV U33654 ( .A(n24950), .Z(n24951) );
  NAND U33655 ( .A(n25019), .B(n25020), .Z(n24950) );
  OR U33656 ( .A(n25021), .B(n25022), .Z(n25020) );
  OR U33657 ( .A(n25023), .B(n25024), .Z(n25019) );
  NAND U33658 ( .A(n25025), .B(n25026), .Z(n24948) );
  OR U33659 ( .A(n25027), .B(n25028), .Z(n25026) );
  OR U33660 ( .A(n25029), .B(n25030), .Z(n25025) );
  NOR U33661 ( .A(n25031), .B(n25032), .Z(n24949) );
  ANDN U33662 ( .B(n25033), .A(n25034), .Z(n24943) );
  IV U33663 ( .A(n25035), .Z(n25033) );
  XNOR U33664 ( .A(n24936), .B(n25036), .Z(n24942) );
  XNOR U33665 ( .A(n24935), .B(n24937), .Z(n25036) );
  NAND U33666 ( .A(n25037), .B(n25038), .Z(n24937) );
  OR U33667 ( .A(n25039), .B(n25040), .Z(n25038) );
  OR U33668 ( .A(n25041), .B(n25042), .Z(n25037) );
  NAND U33669 ( .A(n25043), .B(n25044), .Z(n24935) );
  OR U33670 ( .A(n25045), .B(n25046), .Z(n25044) );
  OR U33671 ( .A(n25047), .B(n25048), .Z(n25043) );
  ANDN U33672 ( .B(n25049), .A(n25050), .Z(n24936) );
  IV U33673 ( .A(n25051), .Z(n25049) );
  XNOR U33674 ( .A(n25016), .B(n25015), .Z(N63179) );
  XOR U33675 ( .A(n25035), .B(n25034), .Z(n25015) );
  XNOR U33676 ( .A(n25050), .B(n25051), .Z(n25034) );
  XNOR U33677 ( .A(n25045), .B(n25046), .Z(n25051) );
  XNOR U33678 ( .A(n25047), .B(n25048), .Z(n25046) );
  XNOR U33679 ( .A(y[4789]), .B(x[4789]), .Z(n25048) );
  XNOR U33680 ( .A(y[4790]), .B(x[4790]), .Z(n25047) );
  XNOR U33681 ( .A(y[4788]), .B(x[4788]), .Z(n25045) );
  XNOR U33682 ( .A(n25039), .B(n25040), .Z(n25050) );
  XNOR U33683 ( .A(y[4785]), .B(x[4785]), .Z(n25040) );
  XNOR U33684 ( .A(n25041), .B(n25042), .Z(n25039) );
  XNOR U33685 ( .A(y[4786]), .B(x[4786]), .Z(n25042) );
  XNOR U33686 ( .A(y[4787]), .B(x[4787]), .Z(n25041) );
  XNOR U33687 ( .A(n25032), .B(n25031), .Z(n25035) );
  XNOR U33688 ( .A(n25027), .B(n25028), .Z(n25031) );
  XNOR U33689 ( .A(y[4782]), .B(x[4782]), .Z(n25028) );
  XNOR U33690 ( .A(n25029), .B(n25030), .Z(n25027) );
  XNOR U33691 ( .A(y[4783]), .B(x[4783]), .Z(n25030) );
  XNOR U33692 ( .A(y[4784]), .B(x[4784]), .Z(n25029) );
  XNOR U33693 ( .A(n25021), .B(n25022), .Z(n25032) );
  XNOR U33694 ( .A(y[4779]), .B(x[4779]), .Z(n25022) );
  XNOR U33695 ( .A(n25023), .B(n25024), .Z(n25021) );
  XNOR U33696 ( .A(y[4780]), .B(x[4780]), .Z(n25024) );
  XNOR U33697 ( .A(y[4781]), .B(x[4781]), .Z(n25023) );
  XOR U33698 ( .A(n24997), .B(n24998), .Z(n25016) );
  XNOR U33699 ( .A(n25013), .B(n25014), .Z(n24998) );
  XNOR U33700 ( .A(n25008), .B(n25009), .Z(n25014) );
  XNOR U33701 ( .A(n25010), .B(n25011), .Z(n25009) );
  XNOR U33702 ( .A(y[4777]), .B(x[4777]), .Z(n25011) );
  XNOR U33703 ( .A(y[4778]), .B(x[4778]), .Z(n25010) );
  XNOR U33704 ( .A(y[4776]), .B(x[4776]), .Z(n25008) );
  XNOR U33705 ( .A(n25002), .B(n25003), .Z(n25013) );
  XNOR U33706 ( .A(y[4773]), .B(x[4773]), .Z(n25003) );
  XNOR U33707 ( .A(n25004), .B(n25005), .Z(n25002) );
  XNOR U33708 ( .A(y[4774]), .B(x[4774]), .Z(n25005) );
  XNOR U33709 ( .A(y[4775]), .B(x[4775]), .Z(n25004) );
  XOR U33710 ( .A(n24996), .B(n24995), .Z(n24997) );
  XNOR U33711 ( .A(n24991), .B(n24992), .Z(n24995) );
  XNOR U33712 ( .A(y[4770]), .B(x[4770]), .Z(n24992) );
  XNOR U33713 ( .A(n24993), .B(n24994), .Z(n24991) );
  XNOR U33714 ( .A(y[4771]), .B(x[4771]), .Z(n24994) );
  XNOR U33715 ( .A(y[4772]), .B(x[4772]), .Z(n24993) );
  XNOR U33716 ( .A(n24985), .B(n24986), .Z(n24996) );
  XNOR U33717 ( .A(y[4767]), .B(x[4767]), .Z(n24986) );
  XNOR U33718 ( .A(n24987), .B(n24988), .Z(n24985) );
  XNOR U33719 ( .A(y[4768]), .B(x[4768]), .Z(n24988) );
  XNOR U33720 ( .A(y[4769]), .B(x[4769]), .Z(n24987) );
  NAND U33721 ( .A(n25052), .B(n25053), .Z(N63170) );
  NANDN U33722 ( .A(n25054), .B(n25055), .Z(n25053) );
  OR U33723 ( .A(n25056), .B(n25057), .Z(n25055) );
  NAND U33724 ( .A(n25056), .B(n25057), .Z(n25052) );
  XOR U33725 ( .A(n25056), .B(n25058), .Z(N63169) );
  XNOR U33726 ( .A(n25054), .B(n25057), .Z(n25058) );
  AND U33727 ( .A(n25059), .B(n25060), .Z(n25057) );
  NANDN U33728 ( .A(n25061), .B(n25062), .Z(n25060) );
  NANDN U33729 ( .A(n25063), .B(n25064), .Z(n25062) );
  NANDN U33730 ( .A(n25064), .B(n25063), .Z(n25059) );
  NAND U33731 ( .A(n25065), .B(n25066), .Z(n25054) );
  NANDN U33732 ( .A(n25067), .B(n25068), .Z(n25066) );
  OR U33733 ( .A(n25069), .B(n25070), .Z(n25068) );
  NAND U33734 ( .A(n25070), .B(n25069), .Z(n25065) );
  AND U33735 ( .A(n25071), .B(n25072), .Z(n25056) );
  NANDN U33736 ( .A(n25073), .B(n25074), .Z(n25072) );
  NANDN U33737 ( .A(n25075), .B(n25076), .Z(n25074) );
  NANDN U33738 ( .A(n25076), .B(n25075), .Z(n25071) );
  XOR U33739 ( .A(n25070), .B(n25077), .Z(N63168) );
  XOR U33740 ( .A(n25067), .B(n25069), .Z(n25077) );
  XNOR U33741 ( .A(n25063), .B(n25078), .Z(n25069) );
  XNOR U33742 ( .A(n25061), .B(n25064), .Z(n25078) );
  NAND U33743 ( .A(n25079), .B(n25080), .Z(n25064) );
  NAND U33744 ( .A(n25081), .B(n25082), .Z(n25080) );
  OR U33745 ( .A(n25083), .B(n25084), .Z(n25081) );
  NANDN U33746 ( .A(n25085), .B(n25083), .Z(n25079) );
  IV U33747 ( .A(n25084), .Z(n25085) );
  NAND U33748 ( .A(n25086), .B(n25087), .Z(n25061) );
  NAND U33749 ( .A(n25088), .B(n25089), .Z(n25087) );
  NANDN U33750 ( .A(n25090), .B(n25091), .Z(n25088) );
  NANDN U33751 ( .A(n25091), .B(n25090), .Z(n25086) );
  AND U33752 ( .A(n25092), .B(n25093), .Z(n25063) );
  NAND U33753 ( .A(n25094), .B(n25095), .Z(n25093) );
  OR U33754 ( .A(n25096), .B(n25097), .Z(n25094) );
  NANDN U33755 ( .A(n25098), .B(n25096), .Z(n25092) );
  NAND U33756 ( .A(n25099), .B(n25100), .Z(n25067) );
  NANDN U33757 ( .A(n25101), .B(n25102), .Z(n25100) );
  OR U33758 ( .A(n25103), .B(n25104), .Z(n25102) );
  NANDN U33759 ( .A(n25105), .B(n25103), .Z(n25099) );
  IV U33760 ( .A(n25104), .Z(n25105) );
  XNOR U33761 ( .A(n25075), .B(n25106), .Z(n25070) );
  XNOR U33762 ( .A(n25073), .B(n25076), .Z(n25106) );
  NAND U33763 ( .A(n25107), .B(n25108), .Z(n25076) );
  NAND U33764 ( .A(n25109), .B(n25110), .Z(n25108) );
  OR U33765 ( .A(n25111), .B(n25112), .Z(n25109) );
  NANDN U33766 ( .A(n25113), .B(n25111), .Z(n25107) );
  IV U33767 ( .A(n25112), .Z(n25113) );
  NAND U33768 ( .A(n25114), .B(n25115), .Z(n25073) );
  NAND U33769 ( .A(n25116), .B(n25117), .Z(n25115) );
  NANDN U33770 ( .A(n25118), .B(n25119), .Z(n25116) );
  NANDN U33771 ( .A(n25119), .B(n25118), .Z(n25114) );
  AND U33772 ( .A(n25120), .B(n25121), .Z(n25075) );
  NAND U33773 ( .A(n25122), .B(n25123), .Z(n25121) );
  OR U33774 ( .A(n25124), .B(n25125), .Z(n25122) );
  NANDN U33775 ( .A(n25126), .B(n25124), .Z(n25120) );
  XNOR U33776 ( .A(n25101), .B(n25127), .Z(N63167) );
  XOR U33777 ( .A(n25103), .B(n25104), .Z(n25127) );
  XNOR U33778 ( .A(n25117), .B(n25128), .Z(n25104) );
  XOR U33779 ( .A(n25118), .B(n25119), .Z(n25128) );
  XOR U33780 ( .A(n25124), .B(n25129), .Z(n25119) );
  XOR U33781 ( .A(n25123), .B(n25126), .Z(n25129) );
  IV U33782 ( .A(n25125), .Z(n25126) );
  NAND U33783 ( .A(n25130), .B(n25131), .Z(n25125) );
  OR U33784 ( .A(n25132), .B(n25133), .Z(n25131) );
  OR U33785 ( .A(n25134), .B(n25135), .Z(n25130) );
  NAND U33786 ( .A(n25136), .B(n25137), .Z(n25123) );
  OR U33787 ( .A(n25138), .B(n25139), .Z(n25137) );
  OR U33788 ( .A(n25140), .B(n25141), .Z(n25136) );
  NOR U33789 ( .A(n25142), .B(n25143), .Z(n25124) );
  ANDN U33790 ( .B(n25144), .A(n25145), .Z(n25118) );
  XNOR U33791 ( .A(n25111), .B(n25146), .Z(n25117) );
  XNOR U33792 ( .A(n25110), .B(n25112), .Z(n25146) );
  NAND U33793 ( .A(n25147), .B(n25148), .Z(n25112) );
  OR U33794 ( .A(n25149), .B(n25150), .Z(n25148) );
  OR U33795 ( .A(n25151), .B(n25152), .Z(n25147) );
  NAND U33796 ( .A(n25153), .B(n25154), .Z(n25110) );
  OR U33797 ( .A(n25155), .B(n25156), .Z(n25154) );
  OR U33798 ( .A(n25157), .B(n25158), .Z(n25153) );
  ANDN U33799 ( .B(n25159), .A(n25160), .Z(n25111) );
  IV U33800 ( .A(n25161), .Z(n25159) );
  ANDN U33801 ( .B(n25162), .A(n25163), .Z(n25103) );
  XOR U33802 ( .A(n25089), .B(n25164), .Z(n25101) );
  XOR U33803 ( .A(n25090), .B(n25091), .Z(n25164) );
  XOR U33804 ( .A(n25096), .B(n25165), .Z(n25091) );
  XOR U33805 ( .A(n25095), .B(n25098), .Z(n25165) );
  IV U33806 ( .A(n25097), .Z(n25098) );
  NAND U33807 ( .A(n25166), .B(n25167), .Z(n25097) );
  OR U33808 ( .A(n25168), .B(n25169), .Z(n25167) );
  OR U33809 ( .A(n25170), .B(n25171), .Z(n25166) );
  NAND U33810 ( .A(n25172), .B(n25173), .Z(n25095) );
  OR U33811 ( .A(n25174), .B(n25175), .Z(n25173) );
  OR U33812 ( .A(n25176), .B(n25177), .Z(n25172) );
  NOR U33813 ( .A(n25178), .B(n25179), .Z(n25096) );
  ANDN U33814 ( .B(n25180), .A(n25181), .Z(n25090) );
  IV U33815 ( .A(n25182), .Z(n25180) );
  XNOR U33816 ( .A(n25083), .B(n25183), .Z(n25089) );
  XNOR U33817 ( .A(n25082), .B(n25084), .Z(n25183) );
  NAND U33818 ( .A(n25184), .B(n25185), .Z(n25084) );
  OR U33819 ( .A(n25186), .B(n25187), .Z(n25185) );
  OR U33820 ( .A(n25188), .B(n25189), .Z(n25184) );
  NAND U33821 ( .A(n25190), .B(n25191), .Z(n25082) );
  OR U33822 ( .A(n25192), .B(n25193), .Z(n25191) );
  OR U33823 ( .A(n25194), .B(n25195), .Z(n25190) );
  ANDN U33824 ( .B(n25196), .A(n25197), .Z(n25083) );
  IV U33825 ( .A(n25198), .Z(n25196) );
  XNOR U33826 ( .A(n25163), .B(n25162), .Z(N63166) );
  XOR U33827 ( .A(n25182), .B(n25181), .Z(n25162) );
  XNOR U33828 ( .A(n25197), .B(n25198), .Z(n25181) );
  XNOR U33829 ( .A(n25192), .B(n25193), .Z(n25198) );
  XNOR U33830 ( .A(n25194), .B(n25195), .Z(n25193) );
  XNOR U33831 ( .A(y[4765]), .B(x[4765]), .Z(n25195) );
  XNOR U33832 ( .A(y[4766]), .B(x[4766]), .Z(n25194) );
  XNOR U33833 ( .A(y[4764]), .B(x[4764]), .Z(n25192) );
  XNOR U33834 ( .A(n25186), .B(n25187), .Z(n25197) );
  XNOR U33835 ( .A(y[4761]), .B(x[4761]), .Z(n25187) );
  XNOR U33836 ( .A(n25188), .B(n25189), .Z(n25186) );
  XNOR U33837 ( .A(y[4762]), .B(x[4762]), .Z(n25189) );
  XNOR U33838 ( .A(y[4763]), .B(x[4763]), .Z(n25188) );
  XNOR U33839 ( .A(n25179), .B(n25178), .Z(n25182) );
  XNOR U33840 ( .A(n25174), .B(n25175), .Z(n25178) );
  XNOR U33841 ( .A(y[4758]), .B(x[4758]), .Z(n25175) );
  XNOR U33842 ( .A(n25176), .B(n25177), .Z(n25174) );
  XNOR U33843 ( .A(y[4759]), .B(x[4759]), .Z(n25177) );
  XNOR U33844 ( .A(y[4760]), .B(x[4760]), .Z(n25176) );
  XNOR U33845 ( .A(n25168), .B(n25169), .Z(n25179) );
  XNOR U33846 ( .A(y[4755]), .B(x[4755]), .Z(n25169) );
  XNOR U33847 ( .A(n25170), .B(n25171), .Z(n25168) );
  XNOR U33848 ( .A(y[4756]), .B(x[4756]), .Z(n25171) );
  XNOR U33849 ( .A(y[4757]), .B(x[4757]), .Z(n25170) );
  XOR U33850 ( .A(n25144), .B(n25145), .Z(n25163) );
  XNOR U33851 ( .A(n25160), .B(n25161), .Z(n25145) );
  XNOR U33852 ( .A(n25155), .B(n25156), .Z(n25161) );
  XNOR U33853 ( .A(n25157), .B(n25158), .Z(n25156) );
  XNOR U33854 ( .A(y[4753]), .B(x[4753]), .Z(n25158) );
  XNOR U33855 ( .A(y[4754]), .B(x[4754]), .Z(n25157) );
  XNOR U33856 ( .A(y[4752]), .B(x[4752]), .Z(n25155) );
  XNOR U33857 ( .A(n25149), .B(n25150), .Z(n25160) );
  XNOR U33858 ( .A(y[4749]), .B(x[4749]), .Z(n25150) );
  XNOR U33859 ( .A(n25151), .B(n25152), .Z(n25149) );
  XNOR U33860 ( .A(y[4750]), .B(x[4750]), .Z(n25152) );
  XNOR U33861 ( .A(y[4751]), .B(x[4751]), .Z(n25151) );
  XOR U33862 ( .A(n25143), .B(n25142), .Z(n25144) );
  XNOR U33863 ( .A(n25138), .B(n25139), .Z(n25142) );
  XNOR U33864 ( .A(y[4746]), .B(x[4746]), .Z(n25139) );
  XNOR U33865 ( .A(n25140), .B(n25141), .Z(n25138) );
  XNOR U33866 ( .A(y[4747]), .B(x[4747]), .Z(n25141) );
  XNOR U33867 ( .A(y[4748]), .B(x[4748]), .Z(n25140) );
  XNOR U33868 ( .A(n25132), .B(n25133), .Z(n25143) );
  XNOR U33869 ( .A(y[4743]), .B(x[4743]), .Z(n25133) );
  XNOR U33870 ( .A(n25134), .B(n25135), .Z(n25132) );
  XNOR U33871 ( .A(y[4744]), .B(x[4744]), .Z(n25135) );
  XNOR U33872 ( .A(y[4745]), .B(x[4745]), .Z(n25134) );
  NAND U33873 ( .A(n25199), .B(n25200), .Z(N63157) );
  NANDN U33874 ( .A(n25201), .B(n25202), .Z(n25200) );
  OR U33875 ( .A(n25203), .B(n25204), .Z(n25202) );
  NAND U33876 ( .A(n25203), .B(n25204), .Z(n25199) );
  XOR U33877 ( .A(n25203), .B(n25205), .Z(N63156) );
  XNOR U33878 ( .A(n25201), .B(n25204), .Z(n25205) );
  AND U33879 ( .A(n25206), .B(n25207), .Z(n25204) );
  NANDN U33880 ( .A(n25208), .B(n25209), .Z(n25207) );
  NANDN U33881 ( .A(n25210), .B(n25211), .Z(n25209) );
  NANDN U33882 ( .A(n25211), .B(n25210), .Z(n25206) );
  NAND U33883 ( .A(n25212), .B(n25213), .Z(n25201) );
  NANDN U33884 ( .A(n25214), .B(n25215), .Z(n25213) );
  OR U33885 ( .A(n25216), .B(n25217), .Z(n25215) );
  NAND U33886 ( .A(n25217), .B(n25216), .Z(n25212) );
  AND U33887 ( .A(n25218), .B(n25219), .Z(n25203) );
  NANDN U33888 ( .A(n25220), .B(n25221), .Z(n25219) );
  NANDN U33889 ( .A(n25222), .B(n25223), .Z(n25221) );
  NANDN U33890 ( .A(n25223), .B(n25222), .Z(n25218) );
  XOR U33891 ( .A(n25217), .B(n25224), .Z(N63155) );
  XOR U33892 ( .A(n25214), .B(n25216), .Z(n25224) );
  XNOR U33893 ( .A(n25210), .B(n25225), .Z(n25216) );
  XNOR U33894 ( .A(n25208), .B(n25211), .Z(n25225) );
  NAND U33895 ( .A(n25226), .B(n25227), .Z(n25211) );
  NAND U33896 ( .A(n25228), .B(n25229), .Z(n25227) );
  OR U33897 ( .A(n25230), .B(n25231), .Z(n25228) );
  NANDN U33898 ( .A(n25232), .B(n25230), .Z(n25226) );
  IV U33899 ( .A(n25231), .Z(n25232) );
  NAND U33900 ( .A(n25233), .B(n25234), .Z(n25208) );
  NAND U33901 ( .A(n25235), .B(n25236), .Z(n25234) );
  NANDN U33902 ( .A(n25237), .B(n25238), .Z(n25235) );
  NANDN U33903 ( .A(n25238), .B(n25237), .Z(n25233) );
  AND U33904 ( .A(n25239), .B(n25240), .Z(n25210) );
  NAND U33905 ( .A(n25241), .B(n25242), .Z(n25240) );
  OR U33906 ( .A(n25243), .B(n25244), .Z(n25241) );
  NANDN U33907 ( .A(n25245), .B(n25243), .Z(n25239) );
  NAND U33908 ( .A(n25246), .B(n25247), .Z(n25214) );
  NANDN U33909 ( .A(n25248), .B(n25249), .Z(n25247) );
  OR U33910 ( .A(n25250), .B(n25251), .Z(n25249) );
  NANDN U33911 ( .A(n25252), .B(n25250), .Z(n25246) );
  IV U33912 ( .A(n25251), .Z(n25252) );
  XNOR U33913 ( .A(n25222), .B(n25253), .Z(n25217) );
  XNOR U33914 ( .A(n25220), .B(n25223), .Z(n25253) );
  NAND U33915 ( .A(n25254), .B(n25255), .Z(n25223) );
  NAND U33916 ( .A(n25256), .B(n25257), .Z(n25255) );
  OR U33917 ( .A(n25258), .B(n25259), .Z(n25256) );
  NANDN U33918 ( .A(n25260), .B(n25258), .Z(n25254) );
  IV U33919 ( .A(n25259), .Z(n25260) );
  NAND U33920 ( .A(n25261), .B(n25262), .Z(n25220) );
  NAND U33921 ( .A(n25263), .B(n25264), .Z(n25262) );
  NANDN U33922 ( .A(n25265), .B(n25266), .Z(n25263) );
  NANDN U33923 ( .A(n25266), .B(n25265), .Z(n25261) );
  AND U33924 ( .A(n25267), .B(n25268), .Z(n25222) );
  NAND U33925 ( .A(n25269), .B(n25270), .Z(n25268) );
  OR U33926 ( .A(n25271), .B(n25272), .Z(n25269) );
  NANDN U33927 ( .A(n25273), .B(n25271), .Z(n25267) );
  XNOR U33928 ( .A(n25248), .B(n25274), .Z(N63154) );
  XOR U33929 ( .A(n25250), .B(n25251), .Z(n25274) );
  XNOR U33930 ( .A(n25264), .B(n25275), .Z(n25251) );
  XOR U33931 ( .A(n25265), .B(n25266), .Z(n25275) );
  XOR U33932 ( .A(n25271), .B(n25276), .Z(n25266) );
  XOR U33933 ( .A(n25270), .B(n25273), .Z(n25276) );
  IV U33934 ( .A(n25272), .Z(n25273) );
  NAND U33935 ( .A(n25277), .B(n25278), .Z(n25272) );
  OR U33936 ( .A(n25279), .B(n25280), .Z(n25278) );
  OR U33937 ( .A(n25281), .B(n25282), .Z(n25277) );
  NAND U33938 ( .A(n25283), .B(n25284), .Z(n25270) );
  OR U33939 ( .A(n25285), .B(n25286), .Z(n25284) );
  OR U33940 ( .A(n25287), .B(n25288), .Z(n25283) );
  NOR U33941 ( .A(n25289), .B(n25290), .Z(n25271) );
  ANDN U33942 ( .B(n25291), .A(n25292), .Z(n25265) );
  XNOR U33943 ( .A(n25258), .B(n25293), .Z(n25264) );
  XNOR U33944 ( .A(n25257), .B(n25259), .Z(n25293) );
  NAND U33945 ( .A(n25294), .B(n25295), .Z(n25259) );
  OR U33946 ( .A(n25296), .B(n25297), .Z(n25295) );
  OR U33947 ( .A(n25298), .B(n25299), .Z(n25294) );
  NAND U33948 ( .A(n25300), .B(n25301), .Z(n25257) );
  OR U33949 ( .A(n25302), .B(n25303), .Z(n25301) );
  OR U33950 ( .A(n25304), .B(n25305), .Z(n25300) );
  ANDN U33951 ( .B(n25306), .A(n25307), .Z(n25258) );
  IV U33952 ( .A(n25308), .Z(n25306) );
  ANDN U33953 ( .B(n25309), .A(n25310), .Z(n25250) );
  XOR U33954 ( .A(n25236), .B(n25311), .Z(n25248) );
  XOR U33955 ( .A(n25237), .B(n25238), .Z(n25311) );
  XOR U33956 ( .A(n25243), .B(n25312), .Z(n25238) );
  XOR U33957 ( .A(n25242), .B(n25245), .Z(n25312) );
  IV U33958 ( .A(n25244), .Z(n25245) );
  NAND U33959 ( .A(n25313), .B(n25314), .Z(n25244) );
  OR U33960 ( .A(n25315), .B(n25316), .Z(n25314) );
  OR U33961 ( .A(n25317), .B(n25318), .Z(n25313) );
  NAND U33962 ( .A(n25319), .B(n25320), .Z(n25242) );
  OR U33963 ( .A(n25321), .B(n25322), .Z(n25320) );
  OR U33964 ( .A(n25323), .B(n25324), .Z(n25319) );
  NOR U33965 ( .A(n25325), .B(n25326), .Z(n25243) );
  ANDN U33966 ( .B(n25327), .A(n25328), .Z(n25237) );
  IV U33967 ( .A(n25329), .Z(n25327) );
  XNOR U33968 ( .A(n25230), .B(n25330), .Z(n25236) );
  XNOR U33969 ( .A(n25229), .B(n25231), .Z(n25330) );
  NAND U33970 ( .A(n25331), .B(n25332), .Z(n25231) );
  OR U33971 ( .A(n25333), .B(n25334), .Z(n25332) );
  OR U33972 ( .A(n25335), .B(n25336), .Z(n25331) );
  NAND U33973 ( .A(n25337), .B(n25338), .Z(n25229) );
  OR U33974 ( .A(n25339), .B(n25340), .Z(n25338) );
  OR U33975 ( .A(n25341), .B(n25342), .Z(n25337) );
  ANDN U33976 ( .B(n25343), .A(n25344), .Z(n25230) );
  IV U33977 ( .A(n25345), .Z(n25343) );
  XNOR U33978 ( .A(n25310), .B(n25309), .Z(N63153) );
  XOR U33979 ( .A(n25329), .B(n25328), .Z(n25309) );
  XNOR U33980 ( .A(n25344), .B(n25345), .Z(n25328) );
  XNOR U33981 ( .A(n25339), .B(n25340), .Z(n25345) );
  XNOR U33982 ( .A(n25341), .B(n25342), .Z(n25340) );
  XNOR U33983 ( .A(y[4741]), .B(x[4741]), .Z(n25342) );
  XNOR U33984 ( .A(y[4742]), .B(x[4742]), .Z(n25341) );
  XNOR U33985 ( .A(y[4740]), .B(x[4740]), .Z(n25339) );
  XNOR U33986 ( .A(n25333), .B(n25334), .Z(n25344) );
  XNOR U33987 ( .A(y[4737]), .B(x[4737]), .Z(n25334) );
  XNOR U33988 ( .A(n25335), .B(n25336), .Z(n25333) );
  XNOR U33989 ( .A(y[4738]), .B(x[4738]), .Z(n25336) );
  XNOR U33990 ( .A(y[4739]), .B(x[4739]), .Z(n25335) );
  XNOR U33991 ( .A(n25326), .B(n25325), .Z(n25329) );
  XNOR U33992 ( .A(n25321), .B(n25322), .Z(n25325) );
  XNOR U33993 ( .A(y[4734]), .B(x[4734]), .Z(n25322) );
  XNOR U33994 ( .A(n25323), .B(n25324), .Z(n25321) );
  XNOR U33995 ( .A(y[4735]), .B(x[4735]), .Z(n25324) );
  XNOR U33996 ( .A(y[4736]), .B(x[4736]), .Z(n25323) );
  XNOR U33997 ( .A(n25315), .B(n25316), .Z(n25326) );
  XNOR U33998 ( .A(y[4731]), .B(x[4731]), .Z(n25316) );
  XNOR U33999 ( .A(n25317), .B(n25318), .Z(n25315) );
  XNOR U34000 ( .A(y[4732]), .B(x[4732]), .Z(n25318) );
  XNOR U34001 ( .A(y[4733]), .B(x[4733]), .Z(n25317) );
  XOR U34002 ( .A(n25291), .B(n25292), .Z(n25310) );
  XNOR U34003 ( .A(n25307), .B(n25308), .Z(n25292) );
  XNOR U34004 ( .A(n25302), .B(n25303), .Z(n25308) );
  XNOR U34005 ( .A(n25304), .B(n25305), .Z(n25303) );
  XNOR U34006 ( .A(y[4729]), .B(x[4729]), .Z(n25305) );
  XNOR U34007 ( .A(y[4730]), .B(x[4730]), .Z(n25304) );
  XNOR U34008 ( .A(y[4728]), .B(x[4728]), .Z(n25302) );
  XNOR U34009 ( .A(n25296), .B(n25297), .Z(n25307) );
  XNOR U34010 ( .A(y[4725]), .B(x[4725]), .Z(n25297) );
  XNOR U34011 ( .A(n25298), .B(n25299), .Z(n25296) );
  XNOR U34012 ( .A(y[4726]), .B(x[4726]), .Z(n25299) );
  XNOR U34013 ( .A(y[4727]), .B(x[4727]), .Z(n25298) );
  XOR U34014 ( .A(n25290), .B(n25289), .Z(n25291) );
  XNOR U34015 ( .A(n25285), .B(n25286), .Z(n25289) );
  XNOR U34016 ( .A(y[4722]), .B(x[4722]), .Z(n25286) );
  XNOR U34017 ( .A(n25287), .B(n25288), .Z(n25285) );
  XNOR U34018 ( .A(y[4723]), .B(x[4723]), .Z(n25288) );
  XNOR U34019 ( .A(y[4724]), .B(x[4724]), .Z(n25287) );
  XNOR U34020 ( .A(n25279), .B(n25280), .Z(n25290) );
  XNOR U34021 ( .A(y[4719]), .B(x[4719]), .Z(n25280) );
  XNOR U34022 ( .A(n25281), .B(n25282), .Z(n25279) );
  XNOR U34023 ( .A(y[4720]), .B(x[4720]), .Z(n25282) );
  XNOR U34024 ( .A(y[4721]), .B(x[4721]), .Z(n25281) );
  NAND U34025 ( .A(n25346), .B(n25347), .Z(N63144) );
  NANDN U34026 ( .A(n25348), .B(n25349), .Z(n25347) );
  OR U34027 ( .A(n25350), .B(n25351), .Z(n25349) );
  NAND U34028 ( .A(n25350), .B(n25351), .Z(n25346) );
  XOR U34029 ( .A(n25350), .B(n25352), .Z(N63143) );
  XNOR U34030 ( .A(n25348), .B(n25351), .Z(n25352) );
  AND U34031 ( .A(n25353), .B(n25354), .Z(n25351) );
  NANDN U34032 ( .A(n25355), .B(n25356), .Z(n25354) );
  NANDN U34033 ( .A(n25357), .B(n25358), .Z(n25356) );
  NANDN U34034 ( .A(n25358), .B(n25357), .Z(n25353) );
  NAND U34035 ( .A(n25359), .B(n25360), .Z(n25348) );
  NANDN U34036 ( .A(n25361), .B(n25362), .Z(n25360) );
  OR U34037 ( .A(n25363), .B(n25364), .Z(n25362) );
  NAND U34038 ( .A(n25364), .B(n25363), .Z(n25359) );
  AND U34039 ( .A(n25365), .B(n25366), .Z(n25350) );
  NANDN U34040 ( .A(n25367), .B(n25368), .Z(n25366) );
  NANDN U34041 ( .A(n25369), .B(n25370), .Z(n25368) );
  NANDN U34042 ( .A(n25370), .B(n25369), .Z(n25365) );
  XOR U34043 ( .A(n25364), .B(n25371), .Z(N63142) );
  XOR U34044 ( .A(n25361), .B(n25363), .Z(n25371) );
  XNOR U34045 ( .A(n25357), .B(n25372), .Z(n25363) );
  XNOR U34046 ( .A(n25355), .B(n25358), .Z(n25372) );
  NAND U34047 ( .A(n25373), .B(n25374), .Z(n25358) );
  NAND U34048 ( .A(n25375), .B(n25376), .Z(n25374) );
  OR U34049 ( .A(n25377), .B(n25378), .Z(n25375) );
  NANDN U34050 ( .A(n25379), .B(n25377), .Z(n25373) );
  IV U34051 ( .A(n25378), .Z(n25379) );
  NAND U34052 ( .A(n25380), .B(n25381), .Z(n25355) );
  NAND U34053 ( .A(n25382), .B(n25383), .Z(n25381) );
  NANDN U34054 ( .A(n25384), .B(n25385), .Z(n25382) );
  NANDN U34055 ( .A(n25385), .B(n25384), .Z(n25380) );
  AND U34056 ( .A(n25386), .B(n25387), .Z(n25357) );
  NAND U34057 ( .A(n25388), .B(n25389), .Z(n25387) );
  OR U34058 ( .A(n25390), .B(n25391), .Z(n25388) );
  NANDN U34059 ( .A(n25392), .B(n25390), .Z(n25386) );
  NAND U34060 ( .A(n25393), .B(n25394), .Z(n25361) );
  NANDN U34061 ( .A(n25395), .B(n25396), .Z(n25394) );
  OR U34062 ( .A(n25397), .B(n25398), .Z(n25396) );
  NANDN U34063 ( .A(n25399), .B(n25397), .Z(n25393) );
  IV U34064 ( .A(n25398), .Z(n25399) );
  XNOR U34065 ( .A(n25369), .B(n25400), .Z(n25364) );
  XNOR U34066 ( .A(n25367), .B(n25370), .Z(n25400) );
  NAND U34067 ( .A(n25401), .B(n25402), .Z(n25370) );
  NAND U34068 ( .A(n25403), .B(n25404), .Z(n25402) );
  OR U34069 ( .A(n25405), .B(n25406), .Z(n25403) );
  NANDN U34070 ( .A(n25407), .B(n25405), .Z(n25401) );
  IV U34071 ( .A(n25406), .Z(n25407) );
  NAND U34072 ( .A(n25408), .B(n25409), .Z(n25367) );
  NAND U34073 ( .A(n25410), .B(n25411), .Z(n25409) );
  NANDN U34074 ( .A(n25412), .B(n25413), .Z(n25410) );
  NANDN U34075 ( .A(n25413), .B(n25412), .Z(n25408) );
  AND U34076 ( .A(n25414), .B(n25415), .Z(n25369) );
  NAND U34077 ( .A(n25416), .B(n25417), .Z(n25415) );
  OR U34078 ( .A(n25418), .B(n25419), .Z(n25416) );
  NANDN U34079 ( .A(n25420), .B(n25418), .Z(n25414) );
  XNOR U34080 ( .A(n25395), .B(n25421), .Z(N63141) );
  XOR U34081 ( .A(n25397), .B(n25398), .Z(n25421) );
  XNOR U34082 ( .A(n25411), .B(n25422), .Z(n25398) );
  XOR U34083 ( .A(n25412), .B(n25413), .Z(n25422) );
  XOR U34084 ( .A(n25418), .B(n25423), .Z(n25413) );
  XOR U34085 ( .A(n25417), .B(n25420), .Z(n25423) );
  IV U34086 ( .A(n25419), .Z(n25420) );
  NAND U34087 ( .A(n25424), .B(n25425), .Z(n25419) );
  OR U34088 ( .A(n25426), .B(n25427), .Z(n25425) );
  OR U34089 ( .A(n25428), .B(n25429), .Z(n25424) );
  NAND U34090 ( .A(n25430), .B(n25431), .Z(n25417) );
  OR U34091 ( .A(n25432), .B(n25433), .Z(n25431) );
  OR U34092 ( .A(n25434), .B(n25435), .Z(n25430) );
  NOR U34093 ( .A(n25436), .B(n25437), .Z(n25418) );
  ANDN U34094 ( .B(n25438), .A(n25439), .Z(n25412) );
  XNOR U34095 ( .A(n25405), .B(n25440), .Z(n25411) );
  XNOR U34096 ( .A(n25404), .B(n25406), .Z(n25440) );
  NAND U34097 ( .A(n25441), .B(n25442), .Z(n25406) );
  OR U34098 ( .A(n25443), .B(n25444), .Z(n25442) );
  OR U34099 ( .A(n25445), .B(n25446), .Z(n25441) );
  NAND U34100 ( .A(n25447), .B(n25448), .Z(n25404) );
  OR U34101 ( .A(n25449), .B(n25450), .Z(n25448) );
  OR U34102 ( .A(n25451), .B(n25452), .Z(n25447) );
  ANDN U34103 ( .B(n25453), .A(n25454), .Z(n25405) );
  IV U34104 ( .A(n25455), .Z(n25453) );
  ANDN U34105 ( .B(n25456), .A(n25457), .Z(n25397) );
  XOR U34106 ( .A(n25383), .B(n25458), .Z(n25395) );
  XOR U34107 ( .A(n25384), .B(n25385), .Z(n25458) );
  XOR U34108 ( .A(n25390), .B(n25459), .Z(n25385) );
  XOR U34109 ( .A(n25389), .B(n25392), .Z(n25459) );
  IV U34110 ( .A(n25391), .Z(n25392) );
  NAND U34111 ( .A(n25460), .B(n25461), .Z(n25391) );
  OR U34112 ( .A(n25462), .B(n25463), .Z(n25461) );
  OR U34113 ( .A(n25464), .B(n25465), .Z(n25460) );
  NAND U34114 ( .A(n25466), .B(n25467), .Z(n25389) );
  OR U34115 ( .A(n25468), .B(n25469), .Z(n25467) );
  OR U34116 ( .A(n25470), .B(n25471), .Z(n25466) );
  NOR U34117 ( .A(n25472), .B(n25473), .Z(n25390) );
  ANDN U34118 ( .B(n25474), .A(n25475), .Z(n25384) );
  IV U34119 ( .A(n25476), .Z(n25474) );
  XNOR U34120 ( .A(n25377), .B(n25477), .Z(n25383) );
  XNOR U34121 ( .A(n25376), .B(n25378), .Z(n25477) );
  NAND U34122 ( .A(n25478), .B(n25479), .Z(n25378) );
  OR U34123 ( .A(n25480), .B(n25481), .Z(n25479) );
  OR U34124 ( .A(n25482), .B(n25483), .Z(n25478) );
  NAND U34125 ( .A(n25484), .B(n25485), .Z(n25376) );
  OR U34126 ( .A(n25486), .B(n25487), .Z(n25485) );
  OR U34127 ( .A(n25488), .B(n25489), .Z(n25484) );
  ANDN U34128 ( .B(n25490), .A(n25491), .Z(n25377) );
  IV U34129 ( .A(n25492), .Z(n25490) );
  XNOR U34130 ( .A(n25457), .B(n25456), .Z(N63140) );
  XOR U34131 ( .A(n25476), .B(n25475), .Z(n25456) );
  XNOR U34132 ( .A(n25491), .B(n25492), .Z(n25475) );
  XNOR U34133 ( .A(n25486), .B(n25487), .Z(n25492) );
  XNOR U34134 ( .A(n25488), .B(n25489), .Z(n25487) );
  XNOR U34135 ( .A(y[4717]), .B(x[4717]), .Z(n25489) );
  XNOR U34136 ( .A(y[4718]), .B(x[4718]), .Z(n25488) );
  XNOR U34137 ( .A(y[4716]), .B(x[4716]), .Z(n25486) );
  XNOR U34138 ( .A(n25480), .B(n25481), .Z(n25491) );
  XNOR U34139 ( .A(y[4713]), .B(x[4713]), .Z(n25481) );
  XNOR U34140 ( .A(n25482), .B(n25483), .Z(n25480) );
  XNOR U34141 ( .A(y[4714]), .B(x[4714]), .Z(n25483) );
  XNOR U34142 ( .A(y[4715]), .B(x[4715]), .Z(n25482) );
  XNOR U34143 ( .A(n25473), .B(n25472), .Z(n25476) );
  XNOR U34144 ( .A(n25468), .B(n25469), .Z(n25472) );
  XNOR U34145 ( .A(y[4710]), .B(x[4710]), .Z(n25469) );
  XNOR U34146 ( .A(n25470), .B(n25471), .Z(n25468) );
  XNOR U34147 ( .A(y[4711]), .B(x[4711]), .Z(n25471) );
  XNOR U34148 ( .A(y[4712]), .B(x[4712]), .Z(n25470) );
  XNOR U34149 ( .A(n25462), .B(n25463), .Z(n25473) );
  XNOR U34150 ( .A(y[4707]), .B(x[4707]), .Z(n25463) );
  XNOR U34151 ( .A(n25464), .B(n25465), .Z(n25462) );
  XNOR U34152 ( .A(y[4708]), .B(x[4708]), .Z(n25465) );
  XNOR U34153 ( .A(y[4709]), .B(x[4709]), .Z(n25464) );
  XOR U34154 ( .A(n25438), .B(n25439), .Z(n25457) );
  XNOR U34155 ( .A(n25454), .B(n25455), .Z(n25439) );
  XNOR U34156 ( .A(n25449), .B(n25450), .Z(n25455) );
  XNOR U34157 ( .A(n25451), .B(n25452), .Z(n25450) );
  XNOR U34158 ( .A(y[4705]), .B(x[4705]), .Z(n25452) );
  XNOR U34159 ( .A(y[4706]), .B(x[4706]), .Z(n25451) );
  XNOR U34160 ( .A(y[4704]), .B(x[4704]), .Z(n25449) );
  XNOR U34161 ( .A(n25443), .B(n25444), .Z(n25454) );
  XNOR U34162 ( .A(y[4701]), .B(x[4701]), .Z(n25444) );
  XNOR U34163 ( .A(n25445), .B(n25446), .Z(n25443) );
  XNOR U34164 ( .A(y[4702]), .B(x[4702]), .Z(n25446) );
  XNOR U34165 ( .A(y[4703]), .B(x[4703]), .Z(n25445) );
  XOR U34166 ( .A(n25437), .B(n25436), .Z(n25438) );
  XNOR U34167 ( .A(n25432), .B(n25433), .Z(n25436) );
  XNOR U34168 ( .A(y[4698]), .B(x[4698]), .Z(n25433) );
  XNOR U34169 ( .A(n25434), .B(n25435), .Z(n25432) );
  XNOR U34170 ( .A(y[4699]), .B(x[4699]), .Z(n25435) );
  XNOR U34171 ( .A(y[4700]), .B(x[4700]), .Z(n25434) );
  XNOR U34172 ( .A(n25426), .B(n25427), .Z(n25437) );
  XNOR U34173 ( .A(y[4695]), .B(x[4695]), .Z(n25427) );
  XNOR U34174 ( .A(n25428), .B(n25429), .Z(n25426) );
  XNOR U34175 ( .A(y[4696]), .B(x[4696]), .Z(n25429) );
  XNOR U34176 ( .A(y[4697]), .B(x[4697]), .Z(n25428) );
  NAND U34177 ( .A(n25493), .B(n25494), .Z(N63131) );
  NANDN U34178 ( .A(n25495), .B(n25496), .Z(n25494) );
  OR U34179 ( .A(n25497), .B(n25498), .Z(n25496) );
  NAND U34180 ( .A(n25497), .B(n25498), .Z(n25493) );
  XOR U34181 ( .A(n25497), .B(n25499), .Z(N63130) );
  XNOR U34182 ( .A(n25495), .B(n25498), .Z(n25499) );
  AND U34183 ( .A(n25500), .B(n25501), .Z(n25498) );
  NANDN U34184 ( .A(n25502), .B(n25503), .Z(n25501) );
  NANDN U34185 ( .A(n25504), .B(n25505), .Z(n25503) );
  NANDN U34186 ( .A(n25505), .B(n25504), .Z(n25500) );
  NAND U34187 ( .A(n25506), .B(n25507), .Z(n25495) );
  NANDN U34188 ( .A(n25508), .B(n25509), .Z(n25507) );
  OR U34189 ( .A(n25510), .B(n25511), .Z(n25509) );
  NAND U34190 ( .A(n25511), .B(n25510), .Z(n25506) );
  AND U34191 ( .A(n25512), .B(n25513), .Z(n25497) );
  NANDN U34192 ( .A(n25514), .B(n25515), .Z(n25513) );
  NANDN U34193 ( .A(n25516), .B(n25517), .Z(n25515) );
  NANDN U34194 ( .A(n25517), .B(n25516), .Z(n25512) );
  XOR U34195 ( .A(n25511), .B(n25518), .Z(N63129) );
  XOR U34196 ( .A(n25508), .B(n25510), .Z(n25518) );
  XNOR U34197 ( .A(n25504), .B(n25519), .Z(n25510) );
  XNOR U34198 ( .A(n25502), .B(n25505), .Z(n25519) );
  NAND U34199 ( .A(n25520), .B(n25521), .Z(n25505) );
  NAND U34200 ( .A(n25522), .B(n25523), .Z(n25521) );
  OR U34201 ( .A(n25524), .B(n25525), .Z(n25522) );
  NANDN U34202 ( .A(n25526), .B(n25524), .Z(n25520) );
  IV U34203 ( .A(n25525), .Z(n25526) );
  NAND U34204 ( .A(n25527), .B(n25528), .Z(n25502) );
  NAND U34205 ( .A(n25529), .B(n25530), .Z(n25528) );
  NANDN U34206 ( .A(n25531), .B(n25532), .Z(n25529) );
  NANDN U34207 ( .A(n25532), .B(n25531), .Z(n25527) );
  AND U34208 ( .A(n25533), .B(n25534), .Z(n25504) );
  NAND U34209 ( .A(n25535), .B(n25536), .Z(n25534) );
  OR U34210 ( .A(n25537), .B(n25538), .Z(n25535) );
  NANDN U34211 ( .A(n25539), .B(n25537), .Z(n25533) );
  NAND U34212 ( .A(n25540), .B(n25541), .Z(n25508) );
  NANDN U34213 ( .A(n25542), .B(n25543), .Z(n25541) );
  OR U34214 ( .A(n25544), .B(n25545), .Z(n25543) );
  NANDN U34215 ( .A(n25546), .B(n25544), .Z(n25540) );
  IV U34216 ( .A(n25545), .Z(n25546) );
  XNOR U34217 ( .A(n25516), .B(n25547), .Z(n25511) );
  XNOR U34218 ( .A(n25514), .B(n25517), .Z(n25547) );
  NAND U34219 ( .A(n25548), .B(n25549), .Z(n25517) );
  NAND U34220 ( .A(n25550), .B(n25551), .Z(n25549) );
  OR U34221 ( .A(n25552), .B(n25553), .Z(n25550) );
  NANDN U34222 ( .A(n25554), .B(n25552), .Z(n25548) );
  IV U34223 ( .A(n25553), .Z(n25554) );
  NAND U34224 ( .A(n25555), .B(n25556), .Z(n25514) );
  NAND U34225 ( .A(n25557), .B(n25558), .Z(n25556) );
  NANDN U34226 ( .A(n25559), .B(n25560), .Z(n25557) );
  NANDN U34227 ( .A(n25560), .B(n25559), .Z(n25555) );
  AND U34228 ( .A(n25561), .B(n25562), .Z(n25516) );
  NAND U34229 ( .A(n25563), .B(n25564), .Z(n25562) );
  OR U34230 ( .A(n25565), .B(n25566), .Z(n25563) );
  NANDN U34231 ( .A(n25567), .B(n25565), .Z(n25561) );
  XNOR U34232 ( .A(n25542), .B(n25568), .Z(N63128) );
  XOR U34233 ( .A(n25544), .B(n25545), .Z(n25568) );
  XNOR U34234 ( .A(n25558), .B(n25569), .Z(n25545) );
  XOR U34235 ( .A(n25559), .B(n25560), .Z(n25569) );
  XOR U34236 ( .A(n25565), .B(n25570), .Z(n25560) );
  XOR U34237 ( .A(n25564), .B(n25567), .Z(n25570) );
  IV U34238 ( .A(n25566), .Z(n25567) );
  NAND U34239 ( .A(n25571), .B(n25572), .Z(n25566) );
  OR U34240 ( .A(n25573), .B(n25574), .Z(n25572) );
  OR U34241 ( .A(n25575), .B(n25576), .Z(n25571) );
  NAND U34242 ( .A(n25577), .B(n25578), .Z(n25564) );
  OR U34243 ( .A(n25579), .B(n25580), .Z(n25578) );
  OR U34244 ( .A(n25581), .B(n25582), .Z(n25577) );
  NOR U34245 ( .A(n25583), .B(n25584), .Z(n25565) );
  ANDN U34246 ( .B(n25585), .A(n25586), .Z(n25559) );
  XNOR U34247 ( .A(n25552), .B(n25587), .Z(n25558) );
  XNOR U34248 ( .A(n25551), .B(n25553), .Z(n25587) );
  NAND U34249 ( .A(n25588), .B(n25589), .Z(n25553) );
  OR U34250 ( .A(n25590), .B(n25591), .Z(n25589) );
  OR U34251 ( .A(n25592), .B(n25593), .Z(n25588) );
  NAND U34252 ( .A(n25594), .B(n25595), .Z(n25551) );
  OR U34253 ( .A(n25596), .B(n25597), .Z(n25595) );
  OR U34254 ( .A(n25598), .B(n25599), .Z(n25594) );
  ANDN U34255 ( .B(n25600), .A(n25601), .Z(n25552) );
  IV U34256 ( .A(n25602), .Z(n25600) );
  ANDN U34257 ( .B(n25603), .A(n25604), .Z(n25544) );
  XOR U34258 ( .A(n25530), .B(n25605), .Z(n25542) );
  XOR U34259 ( .A(n25531), .B(n25532), .Z(n25605) );
  XOR U34260 ( .A(n25537), .B(n25606), .Z(n25532) );
  XOR U34261 ( .A(n25536), .B(n25539), .Z(n25606) );
  IV U34262 ( .A(n25538), .Z(n25539) );
  NAND U34263 ( .A(n25607), .B(n25608), .Z(n25538) );
  OR U34264 ( .A(n25609), .B(n25610), .Z(n25608) );
  OR U34265 ( .A(n25611), .B(n25612), .Z(n25607) );
  NAND U34266 ( .A(n25613), .B(n25614), .Z(n25536) );
  OR U34267 ( .A(n25615), .B(n25616), .Z(n25614) );
  OR U34268 ( .A(n25617), .B(n25618), .Z(n25613) );
  NOR U34269 ( .A(n25619), .B(n25620), .Z(n25537) );
  ANDN U34270 ( .B(n25621), .A(n25622), .Z(n25531) );
  IV U34271 ( .A(n25623), .Z(n25621) );
  XNOR U34272 ( .A(n25524), .B(n25624), .Z(n25530) );
  XNOR U34273 ( .A(n25523), .B(n25525), .Z(n25624) );
  NAND U34274 ( .A(n25625), .B(n25626), .Z(n25525) );
  OR U34275 ( .A(n25627), .B(n25628), .Z(n25626) );
  OR U34276 ( .A(n25629), .B(n25630), .Z(n25625) );
  NAND U34277 ( .A(n25631), .B(n25632), .Z(n25523) );
  OR U34278 ( .A(n25633), .B(n25634), .Z(n25632) );
  OR U34279 ( .A(n25635), .B(n25636), .Z(n25631) );
  ANDN U34280 ( .B(n25637), .A(n25638), .Z(n25524) );
  IV U34281 ( .A(n25639), .Z(n25637) );
  XNOR U34282 ( .A(n25604), .B(n25603), .Z(N63127) );
  XOR U34283 ( .A(n25623), .B(n25622), .Z(n25603) );
  XNOR U34284 ( .A(n25638), .B(n25639), .Z(n25622) );
  XNOR U34285 ( .A(n25633), .B(n25634), .Z(n25639) );
  XNOR U34286 ( .A(n25635), .B(n25636), .Z(n25634) );
  XNOR U34287 ( .A(y[4693]), .B(x[4693]), .Z(n25636) );
  XNOR U34288 ( .A(y[4694]), .B(x[4694]), .Z(n25635) );
  XNOR U34289 ( .A(y[4692]), .B(x[4692]), .Z(n25633) );
  XNOR U34290 ( .A(n25627), .B(n25628), .Z(n25638) );
  XNOR U34291 ( .A(y[4689]), .B(x[4689]), .Z(n25628) );
  XNOR U34292 ( .A(n25629), .B(n25630), .Z(n25627) );
  XNOR U34293 ( .A(y[4690]), .B(x[4690]), .Z(n25630) );
  XNOR U34294 ( .A(y[4691]), .B(x[4691]), .Z(n25629) );
  XNOR U34295 ( .A(n25620), .B(n25619), .Z(n25623) );
  XNOR U34296 ( .A(n25615), .B(n25616), .Z(n25619) );
  XNOR U34297 ( .A(y[4686]), .B(x[4686]), .Z(n25616) );
  XNOR U34298 ( .A(n25617), .B(n25618), .Z(n25615) );
  XNOR U34299 ( .A(y[4687]), .B(x[4687]), .Z(n25618) );
  XNOR U34300 ( .A(y[4688]), .B(x[4688]), .Z(n25617) );
  XNOR U34301 ( .A(n25609), .B(n25610), .Z(n25620) );
  XNOR U34302 ( .A(y[4683]), .B(x[4683]), .Z(n25610) );
  XNOR U34303 ( .A(n25611), .B(n25612), .Z(n25609) );
  XNOR U34304 ( .A(y[4684]), .B(x[4684]), .Z(n25612) );
  XNOR U34305 ( .A(y[4685]), .B(x[4685]), .Z(n25611) );
  XOR U34306 ( .A(n25585), .B(n25586), .Z(n25604) );
  XNOR U34307 ( .A(n25601), .B(n25602), .Z(n25586) );
  XNOR U34308 ( .A(n25596), .B(n25597), .Z(n25602) );
  XNOR U34309 ( .A(n25598), .B(n25599), .Z(n25597) );
  XNOR U34310 ( .A(y[4681]), .B(x[4681]), .Z(n25599) );
  XNOR U34311 ( .A(y[4682]), .B(x[4682]), .Z(n25598) );
  XNOR U34312 ( .A(y[4680]), .B(x[4680]), .Z(n25596) );
  XNOR U34313 ( .A(n25590), .B(n25591), .Z(n25601) );
  XNOR U34314 ( .A(y[4677]), .B(x[4677]), .Z(n25591) );
  XNOR U34315 ( .A(n25592), .B(n25593), .Z(n25590) );
  XNOR U34316 ( .A(y[4678]), .B(x[4678]), .Z(n25593) );
  XNOR U34317 ( .A(y[4679]), .B(x[4679]), .Z(n25592) );
  XOR U34318 ( .A(n25584), .B(n25583), .Z(n25585) );
  XNOR U34319 ( .A(n25579), .B(n25580), .Z(n25583) );
  XNOR U34320 ( .A(y[4674]), .B(x[4674]), .Z(n25580) );
  XNOR U34321 ( .A(n25581), .B(n25582), .Z(n25579) );
  XNOR U34322 ( .A(y[4675]), .B(x[4675]), .Z(n25582) );
  XNOR U34323 ( .A(y[4676]), .B(x[4676]), .Z(n25581) );
  XNOR U34324 ( .A(n25573), .B(n25574), .Z(n25584) );
  XNOR U34325 ( .A(y[4671]), .B(x[4671]), .Z(n25574) );
  XNOR U34326 ( .A(n25575), .B(n25576), .Z(n25573) );
  XNOR U34327 ( .A(y[4672]), .B(x[4672]), .Z(n25576) );
  XNOR U34328 ( .A(y[4673]), .B(x[4673]), .Z(n25575) );
  NAND U34329 ( .A(n25640), .B(n25641), .Z(N63118) );
  NANDN U34330 ( .A(n25642), .B(n25643), .Z(n25641) );
  OR U34331 ( .A(n25644), .B(n25645), .Z(n25643) );
  NAND U34332 ( .A(n25644), .B(n25645), .Z(n25640) );
  XOR U34333 ( .A(n25644), .B(n25646), .Z(N63117) );
  XNOR U34334 ( .A(n25642), .B(n25645), .Z(n25646) );
  AND U34335 ( .A(n25647), .B(n25648), .Z(n25645) );
  NANDN U34336 ( .A(n25649), .B(n25650), .Z(n25648) );
  NANDN U34337 ( .A(n25651), .B(n25652), .Z(n25650) );
  NANDN U34338 ( .A(n25652), .B(n25651), .Z(n25647) );
  NAND U34339 ( .A(n25653), .B(n25654), .Z(n25642) );
  NANDN U34340 ( .A(n25655), .B(n25656), .Z(n25654) );
  OR U34341 ( .A(n25657), .B(n25658), .Z(n25656) );
  NAND U34342 ( .A(n25658), .B(n25657), .Z(n25653) );
  AND U34343 ( .A(n25659), .B(n25660), .Z(n25644) );
  NANDN U34344 ( .A(n25661), .B(n25662), .Z(n25660) );
  NANDN U34345 ( .A(n25663), .B(n25664), .Z(n25662) );
  NANDN U34346 ( .A(n25664), .B(n25663), .Z(n25659) );
  XOR U34347 ( .A(n25658), .B(n25665), .Z(N63116) );
  XOR U34348 ( .A(n25655), .B(n25657), .Z(n25665) );
  XNOR U34349 ( .A(n25651), .B(n25666), .Z(n25657) );
  XNOR U34350 ( .A(n25649), .B(n25652), .Z(n25666) );
  NAND U34351 ( .A(n25667), .B(n25668), .Z(n25652) );
  NAND U34352 ( .A(n25669), .B(n25670), .Z(n25668) );
  OR U34353 ( .A(n25671), .B(n25672), .Z(n25669) );
  NANDN U34354 ( .A(n25673), .B(n25671), .Z(n25667) );
  IV U34355 ( .A(n25672), .Z(n25673) );
  NAND U34356 ( .A(n25674), .B(n25675), .Z(n25649) );
  NAND U34357 ( .A(n25676), .B(n25677), .Z(n25675) );
  NANDN U34358 ( .A(n25678), .B(n25679), .Z(n25676) );
  NANDN U34359 ( .A(n25679), .B(n25678), .Z(n25674) );
  AND U34360 ( .A(n25680), .B(n25681), .Z(n25651) );
  NAND U34361 ( .A(n25682), .B(n25683), .Z(n25681) );
  OR U34362 ( .A(n25684), .B(n25685), .Z(n25682) );
  NANDN U34363 ( .A(n25686), .B(n25684), .Z(n25680) );
  NAND U34364 ( .A(n25687), .B(n25688), .Z(n25655) );
  NANDN U34365 ( .A(n25689), .B(n25690), .Z(n25688) );
  OR U34366 ( .A(n25691), .B(n25692), .Z(n25690) );
  NANDN U34367 ( .A(n25693), .B(n25691), .Z(n25687) );
  IV U34368 ( .A(n25692), .Z(n25693) );
  XNOR U34369 ( .A(n25663), .B(n25694), .Z(n25658) );
  XNOR U34370 ( .A(n25661), .B(n25664), .Z(n25694) );
  NAND U34371 ( .A(n25695), .B(n25696), .Z(n25664) );
  NAND U34372 ( .A(n25697), .B(n25698), .Z(n25696) );
  OR U34373 ( .A(n25699), .B(n25700), .Z(n25697) );
  NANDN U34374 ( .A(n25701), .B(n25699), .Z(n25695) );
  IV U34375 ( .A(n25700), .Z(n25701) );
  NAND U34376 ( .A(n25702), .B(n25703), .Z(n25661) );
  NAND U34377 ( .A(n25704), .B(n25705), .Z(n25703) );
  NANDN U34378 ( .A(n25706), .B(n25707), .Z(n25704) );
  NANDN U34379 ( .A(n25707), .B(n25706), .Z(n25702) );
  AND U34380 ( .A(n25708), .B(n25709), .Z(n25663) );
  NAND U34381 ( .A(n25710), .B(n25711), .Z(n25709) );
  OR U34382 ( .A(n25712), .B(n25713), .Z(n25710) );
  NANDN U34383 ( .A(n25714), .B(n25712), .Z(n25708) );
  XNOR U34384 ( .A(n25689), .B(n25715), .Z(N63115) );
  XOR U34385 ( .A(n25691), .B(n25692), .Z(n25715) );
  XNOR U34386 ( .A(n25705), .B(n25716), .Z(n25692) );
  XOR U34387 ( .A(n25706), .B(n25707), .Z(n25716) );
  XOR U34388 ( .A(n25712), .B(n25717), .Z(n25707) );
  XOR U34389 ( .A(n25711), .B(n25714), .Z(n25717) );
  IV U34390 ( .A(n25713), .Z(n25714) );
  NAND U34391 ( .A(n25718), .B(n25719), .Z(n25713) );
  OR U34392 ( .A(n25720), .B(n25721), .Z(n25719) );
  OR U34393 ( .A(n25722), .B(n25723), .Z(n25718) );
  NAND U34394 ( .A(n25724), .B(n25725), .Z(n25711) );
  OR U34395 ( .A(n25726), .B(n25727), .Z(n25725) );
  OR U34396 ( .A(n25728), .B(n25729), .Z(n25724) );
  NOR U34397 ( .A(n25730), .B(n25731), .Z(n25712) );
  ANDN U34398 ( .B(n25732), .A(n25733), .Z(n25706) );
  XNOR U34399 ( .A(n25699), .B(n25734), .Z(n25705) );
  XNOR U34400 ( .A(n25698), .B(n25700), .Z(n25734) );
  NAND U34401 ( .A(n25735), .B(n25736), .Z(n25700) );
  OR U34402 ( .A(n25737), .B(n25738), .Z(n25736) );
  OR U34403 ( .A(n25739), .B(n25740), .Z(n25735) );
  NAND U34404 ( .A(n25741), .B(n25742), .Z(n25698) );
  OR U34405 ( .A(n25743), .B(n25744), .Z(n25742) );
  OR U34406 ( .A(n25745), .B(n25746), .Z(n25741) );
  ANDN U34407 ( .B(n25747), .A(n25748), .Z(n25699) );
  IV U34408 ( .A(n25749), .Z(n25747) );
  ANDN U34409 ( .B(n25750), .A(n25751), .Z(n25691) );
  XOR U34410 ( .A(n25677), .B(n25752), .Z(n25689) );
  XOR U34411 ( .A(n25678), .B(n25679), .Z(n25752) );
  XOR U34412 ( .A(n25684), .B(n25753), .Z(n25679) );
  XOR U34413 ( .A(n25683), .B(n25686), .Z(n25753) );
  IV U34414 ( .A(n25685), .Z(n25686) );
  NAND U34415 ( .A(n25754), .B(n25755), .Z(n25685) );
  OR U34416 ( .A(n25756), .B(n25757), .Z(n25755) );
  OR U34417 ( .A(n25758), .B(n25759), .Z(n25754) );
  NAND U34418 ( .A(n25760), .B(n25761), .Z(n25683) );
  OR U34419 ( .A(n25762), .B(n25763), .Z(n25761) );
  OR U34420 ( .A(n25764), .B(n25765), .Z(n25760) );
  NOR U34421 ( .A(n25766), .B(n25767), .Z(n25684) );
  ANDN U34422 ( .B(n25768), .A(n25769), .Z(n25678) );
  IV U34423 ( .A(n25770), .Z(n25768) );
  XNOR U34424 ( .A(n25671), .B(n25771), .Z(n25677) );
  XNOR U34425 ( .A(n25670), .B(n25672), .Z(n25771) );
  NAND U34426 ( .A(n25772), .B(n25773), .Z(n25672) );
  OR U34427 ( .A(n25774), .B(n25775), .Z(n25773) );
  OR U34428 ( .A(n25776), .B(n25777), .Z(n25772) );
  NAND U34429 ( .A(n25778), .B(n25779), .Z(n25670) );
  OR U34430 ( .A(n25780), .B(n25781), .Z(n25779) );
  OR U34431 ( .A(n25782), .B(n25783), .Z(n25778) );
  ANDN U34432 ( .B(n25784), .A(n25785), .Z(n25671) );
  IV U34433 ( .A(n25786), .Z(n25784) );
  XNOR U34434 ( .A(n25751), .B(n25750), .Z(N63114) );
  XOR U34435 ( .A(n25770), .B(n25769), .Z(n25750) );
  XNOR U34436 ( .A(n25785), .B(n25786), .Z(n25769) );
  XNOR U34437 ( .A(n25780), .B(n25781), .Z(n25786) );
  XNOR U34438 ( .A(n25782), .B(n25783), .Z(n25781) );
  XNOR U34439 ( .A(y[4669]), .B(x[4669]), .Z(n25783) );
  XNOR U34440 ( .A(y[4670]), .B(x[4670]), .Z(n25782) );
  XNOR U34441 ( .A(y[4668]), .B(x[4668]), .Z(n25780) );
  XNOR U34442 ( .A(n25774), .B(n25775), .Z(n25785) );
  XNOR U34443 ( .A(y[4665]), .B(x[4665]), .Z(n25775) );
  XNOR U34444 ( .A(n25776), .B(n25777), .Z(n25774) );
  XNOR U34445 ( .A(y[4666]), .B(x[4666]), .Z(n25777) );
  XNOR U34446 ( .A(y[4667]), .B(x[4667]), .Z(n25776) );
  XNOR U34447 ( .A(n25767), .B(n25766), .Z(n25770) );
  XNOR U34448 ( .A(n25762), .B(n25763), .Z(n25766) );
  XNOR U34449 ( .A(y[4662]), .B(x[4662]), .Z(n25763) );
  XNOR U34450 ( .A(n25764), .B(n25765), .Z(n25762) );
  XNOR U34451 ( .A(y[4663]), .B(x[4663]), .Z(n25765) );
  XNOR U34452 ( .A(y[4664]), .B(x[4664]), .Z(n25764) );
  XNOR U34453 ( .A(n25756), .B(n25757), .Z(n25767) );
  XNOR U34454 ( .A(y[4659]), .B(x[4659]), .Z(n25757) );
  XNOR U34455 ( .A(n25758), .B(n25759), .Z(n25756) );
  XNOR U34456 ( .A(y[4660]), .B(x[4660]), .Z(n25759) );
  XNOR U34457 ( .A(y[4661]), .B(x[4661]), .Z(n25758) );
  XOR U34458 ( .A(n25732), .B(n25733), .Z(n25751) );
  XNOR U34459 ( .A(n25748), .B(n25749), .Z(n25733) );
  XNOR U34460 ( .A(n25743), .B(n25744), .Z(n25749) );
  XNOR U34461 ( .A(n25745), .B(n25746), .Z(n25744) );
  XNOR U34462 ( .A(y[4657]), .B(x[4657]), .Z(n25746) );
  XNOR U34463 ( .A(y[4658]), .B(x[4658]), .Z(n25745) );
  XNOR U34464 ( .A(y[4656]), .B(x[4656]), .Z(n25743) );
  XNOR U34465 ( .A(n25737), .B(n25738), .Z(n25748) );
  XNOR U34466 ( .A(y[4653]), .B(x[4653]), .Z(n25738) );
  XNOR U34467 ( .A(n25739), .B(n25740), .Z(n25737) );
  XNOR U34468 ( .A(y[4654]), .B(x[4654]), .Z(n25740) );
  XNOR U34469 ( .A(y[4655]), .B(x[4655]), .Z(n25739) );
  XOR U34470 ( .A(n25731), .B(n25730), .Z(n25732) );
  XNOR U34471 ( .A(n25726), .B(n25727), .Z(n25730) );
  XNOR U34472 ( .A(y[4650]), .B(x[4650]), .Z(n25727) );
  XNOR U34473 ( .A(n25728), .B(n25729), .Z(n25726) );
  XNOR U34474 ( .A(y[4651]), .B(x[4651]), .Z(n25729) );
  XNOR U34475 ( .A(y[4652]), .B(x[4652]), .Z(n25728) );
  XNOR U34476 ( .A(n25720), .B(n25721), .Z(n25731) );
  XNOR U34477 ( .A(y[4647]), .B(x[4647]), .Z(n25721) );
  XNOR U34478 ( .A(n25722), .B(n25723), .Z(n25720) );
  XNOR U34479 ( .A(y[4648]), .B(x[4648]), .Z(n25723) );
  XNOR U34480 ( .A(y[4649]), .B(x[4649]), .Z(n25722) );
  NAND U34481 ( .A(n25787), .B(n25788), .Z(N63105) );
  NANDN U34482 ( .A(n25789), .B(n25790), .Z(n25788) );
  OR U34483 ( .A(n25791), .B(n25792), .Z(n25790) );
  NAND U34484 ( .A(n25791), .B(n25792), .Z(n25787) );
  XOR U34485 ( .A(n25791), .B(n25793), .Z(N63104) );
  XNOR U34486 ( .A(n25789), .B(n25792), .Z(n25793) );
  AND U34487 ( .A(n25794), .B(n25795), .Z(n25792) );
  NANDN U34488 ( .A(n25796), .B(n25797), .Z(n25795) );
  NANDN U34489 ( .A(n25798), .B(n25799), .Z(n25797) );
  NANDN U34490 ( .A(n25799), .B(n25798), .Z(n25794) );
  NAND U34491 ( .A(n25800), .B(n25801), .Z(n25789) );
  NANDN U34492 ( .A(n25802), .B(n25803), .Z(n25801) );
  OR U34493 ( .A(n25804), .B(n25805), .Z(n25803) );
  NAND U34494 ( .A(n25805), .B(n25804), .Z(n25800) );
  AND U34495 ( .A(n25806), .B(n25807), .Z(n25791) );
  NANDN U34496 ( .A(n25808), .B(n25809), .Z(n25807) );
  NANDN U34497 ( .A(n25810), .B(n25811), .Z(n25809) );
  NANDN U34498 ( .A(n25811), .B(n25810), .Z(n25806) );
  XOR U34499 ( .A(n25805), .B(n25812), .Z(N63103) );
  XOR U34500 ( .A(n25802), .B(n25804), .Z(n25812) );
  XNOR U34501 ( .A(n25798), .B(n25813), .Z(n25804) );
  XNOR U34502 ( .A(n25796), .B(n25799), .Z(n25813) );
  NAND U34503 ( .A(n25814), .B(n25815), .Z(n25799) );
  NAND U34504 ( .A(n25816), .B(n25817), .Z(n25815) );
  OR U34505 ( .A(n25818), .B(n25819), .Z(n25816) );
  NANDN U34506 ( .A(n25820), .B(n25818), .Z(n25814) );
  IV U34507 ( .A(n25819), .Z(n25820) );
  NAND U34508 ( .A(n25821), .B(n25822), .Z(n25796) );
  NAND U34509 ( .A(n25823), .B(n25824), .Z(n25822) );
  NANDN U34510 ( .A(n25825), .B(n25826), .Z(n25823) );
  NANDN U34511 ( .A(n25826), .B(n25825), .Z(n25821) );
  AND U34512 ( .A(n25827), .B(n25828), .Z(n25798) );
  NAND U34513 ( .A(n25829), .B(n25830), .Z(n25828) );
  OR U34514 ( .A(n25831), .B(n25832), .Z(n25829) );
  NANDN U34515 ( .A(n25833), .B(n25831), .Z(n25827) );
  NAND U34516 ( .A(n25834), .B(n25835), .Z(n25802) );
  NANDN U34517 ( .A(n25836), .B(n25837), .Z(n25835) );
  OR U34518 ( .A(n25838), .B(n25839), .Z(n25837) );
  NANDN U34519 ( .A(n25840), .B(n25838), .Z(n25834) );
  IV U34520 ( .A(n25839), .Z(n25840) );
  XNOR U34521 ( .A(n25810), .B(n25841), .Z(n25805) );
  XNOR U34522 ( .A(n25808), .B(n25811), .Z(n25841) );
  NAND U34523 ( .A(n25842), .B(n25843), .Z(n25811) );
  NAND U34524 ( .A(n25844), .B(n25845), .Z(n25843) );
  OR U34525 ( .A(n25846), .B(n25847), .Z(n25844) );
  NANDN U34526 ( .A(n25848), .B(n25846), .Z(n25842) );
  IV U34527 ( .A(n25847), .Z(n25848) );
  NAND U34528 ( .A(n25849), .B(n25850), .Z(n25808) );
  NAND U34529 ( .A(n25851), .B(n25852), .Z(n25850) );
  NANDN U34530 ( .A(n25853), .B(n25854), .Z(n25851) );
  NANDN U34531 ( .A(n25854), .B(n25853), .Z(n25849) );
  AND U34532 ( .A(n25855), .B(n25856), .Z(n25810) );
  NAND U34533 ( .A(n25857), .B(n25858), .Z(n25856) );
  OR U34534 ( .A(n25859), .B(n25860), .Z(n25857) );
  NANDN U34535 ( .A(n25861), .B(n25859), .Z(n25855) );
  XNOR U34536 ( .A(n25836), .B(n25862), .Z(N63102) );
  XOR U34537 ( .A(n25838), .B(n25839), .Z(n25862) );
  XNOR U34538 ( .A(n25852), .B(n25863), .Z(n25839) );
  XOR U34539 ( .A(n25853), .B(n25854), .Z(n25863) );
  XOR U34540 ( .A(n25859), .B(n25864), .Z(n25854) );
  XOR U34541 ( .A(n25858), .B(n25861), .Z(n25864) );
  IV U34542 ( .A(n25860), .Z(n25861) );
  NAND U34543 ( .A(n25865), .B(n25866), .Z(n25860) );
  OR U34544 ( .A(n25867), .B(n25868), .Z(n25866) );
  OR U34545 ( .A(n25869), .B(n25870), .Z(n25865) );
  NAND U34546 ( .A(n25871), .B(n25872), .Z(n25858) );
  OR U34547 ( .A(n25873), .B(n25874), .Z(n25872) );
  OR U34548 ( .A(n25875), .B(n25876), .Z(n25871) );
  NOR U34549 ( .A(n25877), .B(n25878), .Z(n25859) );
  ANDN U34550 ( .B(n25879), .A(n25880), .Z(n25853) );
  XNOR U34551 ( .A(n25846), .B(n25881), .Z(n25852) );
  XNOR U34552 ( .A(n25845), .B(n25847), .Z(n25881) );
  NAND U34553 ( .A(n25882), .B(n25883), .Z(n25847) );
  OR U34554 ( .A(n25884), .B(n25885), .Z(n25883) );
  OR U34555 ( .A(n25886), .B(n25887), .Z(n25882) );
  NAND U34556 ( .A(n25888), .B(n25889), .Z(n25845) );
  OR U34557 ( .A(n25890), .B(n25891), .Z(n25889) );
  OR U34558 ( .A(n25892), .B(n25893), .Z(n25888) );
  ANDN U34559 ( .B(n25894), .A(n25895), .Z(n25846) );
  IV U34560 ( .A(n25896), .Z(n25894) );
  ANDN U34561 ( .B(n25897), .A(n25898), .Z(n25838) );
  XOR U34562 ( .A(n25824), .B(n25899), .Z(n25836) );
  XOR U34563 ( .A(n25825), .B(n25826), .Z(n25899) );
  XOR U34564 ( .A(n25831), .B(n25900), .Z(n25826) );
  XOR U34565 ( .A(n25830), .B(n25833), .Z(n25900) );
  IV U34566 ( .A(n25832), .Z(n25833) );
  NAND U34567 ( .A(n25901), .B(n25902), .Z(n25832) );
  OR U34568 ( .A(n25903), .B(n25904), .Z(n25902) );
  OR U34569 ( .A(n25905), .B(n25906), .Z(n25901) );
  NAND U34570 ( .A(n25907), .B(n25908), .Z(n25830) );
  OR U34571 ( .A(n25909), .B(n25910), .Z(n25908) );
  OR U34572 ( .A(n25911), .B(n25912), .Z(n25907) );
  NOR U34573 ( .A(n25913), .B(n25914), .Z(n25831) );
  ANDN U34574 ( .B(n25915), .A(n25916), .Z(n25825) );
  IV U34575 ( .A(n25917), .Z(n25915) );
  XNOR U34576 ( .A(n25818), .B(n25918), .Z(n25824) );
  XNOR U34577 ( .A(n25817), .B(n25819), .Z(n25918) );
  NAND U34578 ( .A(n25919), .B(n25920), .Z(n25819) );
  OR U34579 ( .A(n25921), .B(n25922), .Z(n25920) );
  OR U34580 ( .A(n25923), .B(n25924), .Z(n25919) );
  NAND U34581 ( .A(n25925), .B(n25926), .Z(n25817) );
  OR U34582 ( .A(n25927), .B(n25928), .Z(n25926) );
  OR U34583 ( .A(n25929), .B(n25930), .Z(n25925) );
  ANDN U34584 ( .B(n25931), .A(n25932), .Z(n25818) );
  IV U34585 ( .A(n25933), .Z(n25931) );
  XNOR U34586 ( .A(n25898), .B(n25897), .Z(N63101) );
  XOR U34587 ( .A(n25917), .B(n25916), .Z(n25897) );
  XNOR U34588 ( .A(n25932), .B(n25933), .Z(n25916) );
  XNOR U34589 ( .A(n25927), .B(n25928), .Z(n25933) );
  XNOR U34590 ( .A(n25929), .B(n25930), .Z(n25928) );
  XNOR U34591 ( .A(y[4645]), .B(x[4645]), .Z(n25930) );
  XNOR U34592 ( .A(y[4646]), .B(x[4646]), .Z(n25929) );
  XNOR U34593 ( .A(y[4644]), .B(x[4644]), .Z(n25927) );
  XNOR U34594 ( .A(n25921), .B(n25922), .Z(n25932) );
  XNOR U34595 ( .A(y[4641]), .B(x[4641]), .Z(n25922) );
  XNOR U34596 ( .A(n25923), .B(n25924), .Z(n25921) );
  XNOR U34597 ( .A(y[4642]), .B(x[4642]), .Z(n25924) );
  XNOR U34598 ( .A(y[4643]), .B(x[4643]), .Z(n25923) );
  XNOR U34599 ( .A(n25914), .B(n25913), .Z(n25917) );
  XNOR U34600 ( .A(n25909), .B(n25910), .Z(n25913) );
  XNOR U34601 ( .A(y[4638]), .B(x[4638]), .Z(n25910) );
  XNOR U34602 ( .A(n25911), .B(n25912), .Z(n25909) );
  XNOR U34603 ( .A(y[4639]), .B(x[4639]), .Z(n25912) );
  XNOR U34604 ( .A(y[4640]), .B(x[4640]), .Z(n25911) );
  XNOR U34605 ( .A(n25903), .B(n25904), .Z(n25914) );
  XNOR U34606 ( .A(y[4635]), .B(x[4635]), .Z(n25904) );
  XNOR U34607 ( .A(n25905), .B(n25906), .Z(n25903) );
  XNOR U34608 ( .A(y[4636]), .B(x[4636]), .Z(n25906) );
  XNOR U34609 ( .A(y[4637]), .B(x[4637]), .Z(n25905) );
  XOR U34610 ( .A(n25879), .B(n25880), .Z(n25898) );
  XNOR U34611 ( .A(n25895), .B(n25896), .Z(n25880) );
  XNOR U34612 ( .A(n25890), .B(n25891), .Z(n25896) );
  XNOR U34613 ( .A(n25892), .B(n25893), .Z(n25891) );
  XNOR U34614 ( .A(y[4633]), .B(x[4633]), .Z(n25893) );
  XNOR U34615 ( .A(y[4634]), .B(x[4634]), .Z(n25892) );
  XNOR U34616 ( .A(y[4632]), .B(x[4632]), .Z(n25890) );
  XNOR U34617 ( .A(n25884), .B(n25885), .Z(n25895) );
  XNOR U34618 ( .A(y[4629]), .B(x[4629]), .Z(n25885) );
  XNOR U34619 ( .A(n25886), .B(n25887), .Z(n25884) );
  XNOR U34620 ( .A(y[4630]), .B(x[4630]), .Z(n25887) );
  XNOR U34621 ( .A(y[4631]), .B(x[4631]), .Z(n25886) );
  XOR U34622 ( .A(n25878), .B(n25877), .Z(n25879) );
  XNOR U34623 ( .A(n25873), .B(n25874), .Z(n25877) );
  XNOR U34624 ( .A(y[4626]), .B(x[4626]), .Z(n25874) );
  XNOR U34625 ( .A(n25875), .B(n25876), .Z(n25873) );
  XNOR U34626 ( .A(y[4627]), .B(x[4627]), .Z(n25876) );
  XNOR U34627 ( .A(y[4628]), .B(x[4628]), .Z(n25875) );
  XNOR U34628 ( .A(n25867), .B(n25868), .Z(n25878) );
  XNOR U34629 ( .A(y[4623]), .B(x[4623]), .Z(n25868) );
  XNOR U34630 ( .A(n25869), .B(n25870), .Z(n25867) );
  XNOR U34631 ( .A(y[4624]), .B(x[4624]), .Z(n25870) );
  XNOR U34632 ( .A(y[4625]), .B(x[4625]), .Z(n25869) );
  NAND U34633 ( .A(n25934), .B(n25935), .Z(N63092) );
  NANDN U34634 ( .A(n25936), .B(n25937), .Z(n25935) );
  OR U34635 ( .A(n25938), .B(n25939), .Z(n25937) );
  NAND U34636 ( .A(n25938), .B(n25939), .Z(n25934) );
  XOR U34637 ( .A(n25938), .B(n25940), .Z(N63091) );
  XNOR U34638 ( .A(n25936), .B(n25939), .Z(n25940) );
  AND U34639 ( .A(n25941), .B(n25942), .Z(n25939) );
  NANDN U34640 ( .A(n25943), .B(n25944), .Z(n25942) );
  NANDN U34641 ( .A(n25945), .B(n25946), .Z(n25944) );
  NANDN U34642 ( .A(n25946), .B(n25945), .Z(n25941) );
  NAND U34643 ( .A(n25947), .B(n25948), .Z(n25936) );
  NANDN U34644 ( .A(n25949), .B(n25950), .Z(n25948) );
  OR U34645 ( .A(n25951), .B(n25952), .Z(n25950) );
  NAND U34646 ( .A(n25952), .B(n25951), .Z(n25947) );
  AND U34647 ( .A(n25953), .B(n25954), .Z(n25938) );
  NANDN U34648 ( .A(n25955), .B(n25956), .Z(n25954) );
  NANDN U34649 ( .A(n25957), .B(n25958), .Z(n25956) );
  NANDN U34650 ( .A(n25958), .B(n25957), .Z(n25953) );
  XOR U34651 ( .A(n25952), .B(n25959), .Z(N63090) );
  XOR U34652 ( .A(n25949), .B(n25951), .Z(n25959) );
  XNOR U34653 ( .A(n25945), .B(n25960), .Z(n25951) );
  XNOR U34654 ( .A(n25943), .B(n25946), .Z(n25960) );
  NAND U34655 ( .A(n25961), .B(n25962), .Z(n25946) );
  NAND U34656 ( .A(n25963), .B(n25964), .Z(n25962) );
  OR U34657 ( .A(n25965), .B(n25966), .Z(n25963) );
  NANDN U34658 ( .A(n25967), .B(n25965), .Z(n25961) );
  IV U34659 ( .A(n25966), .Z(n25967) );
  NAND U34660 ( .A(n25968), .B(n25969), .Z(n25943) );
  NAND U34661 ( .A(n25970), .B(n25971), .Z(n25969) );
  NANDN U34662 ( .A(n25972), .B(n25973), .Z(n25970) );
  NANDN U34663 ( .A(n25973), .B(n25972), .Z(n25968) );
  AND U34664 ( .A(n25974), .B(n25975), .Z(n25945) );
  NAND U34665 ( .A(n25976), .B(n25977), .Z(n25975) );
  OR U34666 ( .A(n25978), .B(n25979), .Z(n25976) );
  NANDN U34667 ( .A(n25980), .B(n25978), .Z(n25974) );
  NAND U34668 ( .A(n25981), .B(n25982), .Z(n25949) );
  NANDN U34669 ( .A(n25983), .B(n25984), .Z(n25982) );
  OR U34670 ( .A(n25985), .B(n25986), .Z(n25984) );
  NANDN U34671 ( .A(n25987), .B(n25985), .Z(n25981) );
  IV U34672 ( .A(n25986), .Z(n25987) );
  XNOR U34673 ( .A(n25957), .B(n25988), .Z(n25952) );
  XNOR U34674 ( .A(n25955), .B(n25958), .Z(n25988) );
  NAND U34675 ( .A(n25989), .B(n25990), .Z(n25958) );
  NAND U34676 ( .A(n25991), .B(n25992), .Z(n25990) );
  OR U34677 ( .A(n25993), .B(n25994), .Z(n25991) );
  NANDN U34678 ( .A(n25995), .B(n25993), .Z(n25989) );
  IV U34679 ( .A(n25994), .Z(n25995) );
  NAND U34680 ( .A(n25996), .B(n25997), .Z(n25955) );
  NAND U34681 ( .A(n25998), .B(n25999), .Z(n25997) );
  NANDN U34682 ( .A(n26000), .B(n26001), .Z(n25998) );
  NANDN U34683 ( .A(n26001), .B(n26000), .Z(n25996) );
  AND U34684 ( .A(n26002), .B(n26003), .Z(n25957) );
  NAND U34685 ( .A(n26004), .B(n26005), .Z(n26003) );
  OR U34686 ( .A(n26006), .B(n26007), .Z(n26004) );
  NANDN U34687 ( .A(n26008), .B(n26006), .Z(n26002) );
  XNOR U34688 ( .A(n25983), .B(n26009), .Z(N63089) );
  XOR U34689 ( .A(n25985), .B(n25986), .Z(n26009) );
  XNOR U34690 ( .A(n25999), .B(n26010), .Z(n25986) );
  XOR U34691 ( .A(n26000), .B(n26001), .Z(n26010) );
  XOR U34692 ( .A(n26006), .B(n26011), .Z(n26001) );
  XOR U34693 ( .A(n26005), .B(n26008), .Z(n26011) );
  IV U34694 ( .A(n26007), .Z(n26008) );
  NAND U34695 ( .A(n26012), .B(n26013), .Z(n26007) );
  OR U34696 ( .A(n26014), .B(n26015), .Z(n26013) );
  OR U34697 ( .A(n26016), .B(n26017), .Z(n26012) );
  NAND U34698 ( .A(n26018), .B(n26019), .Z(n26005) );
  OR U34699 ( .A(n26020), .B(n26021), .Z(n26019) );
  OR U34700 ( .A(n26022), .B(n26023), .Z(n26018) );
  NOR U34701 ( .A(n26024), .B(n26025), .Z(n26006) );
  ANDN U34702 ( .B(n26026), .A(n26027), .Z(n26000) );
  XNOR U34703 ( .A(n25993), .B(n26028), .Z(n25999) );
  XNOR U34704 ( .A(n25992), .B(n25994), .Z(n26028) );
  NAND U34705 ( .A(n26029), .B(n26030), .Z(n25994) );
  OR U34706 ( .A(n26031), .B(n26032), .Z(n26030) );
  OR U34707 ( .A(n26033), .B(n26034), .Z(n26029) );
  NAND U34708 ( .A(n26035), .B(n26036), .Z(n25992) );
  OR U34709 ( .A(n26037), .B(n26038), .Z(n26036) );
  OR U34710 ( .A(n26039), .B(n26040), .Z(n26035) );
  ANDN U34711 ( .B(n26041), .A(n26042), .Z(n25993) );
  IV U34712 ( .A(n26043), .Z(n26041) );
  ANDN U34713 ( .B(n26044), .A(n26045), .Z(n25985) );
  XOR U34714 ( .A(n25971), .B(n26046), .Z(n25983) );
  XOR U34715 ( .A(n25972), .B(n25973), .Z(n26046) );
  XOR U34716 ( .A(n25978), .B(n26047), .Z(n25973) );
  XOR U34717 ( .A(n25977), .B(n25980), .Z(n26047) );
  IV U34718 ( .A(n25979), .Z(n25980) );
  NAND U34719 ( .A(n26048), .B(n26049), .Z(n25979) );
  OR U34720 ( .A(n26050), .B(n26051), .Z(n26049) );
  OR U34721 ( .A(n26052), .B(n26053), .Z(n26048) );
  NAND U34722 ( .A(n26054), .B(n26055), .Z(n25977) );
  OR U34723 ( .A(n26056), .B(n26057), .Z(n26055) );
  OR U34724 ( .A(n26058), .B(n26059), .Z(n26054) );
  NOR U34725 ( .A(n26060), .B(n26061), .Z(n25978) );
  ANDN U34726 ( .B(n26062), .A(n26063), .Z(n25972) );
  IV U34727 ( .A(n26064), .Z(n26062) );
  XNOR U34728 ( .A(n25965), .B(n26065), .Z(n25971) );
  XNOR U34729 ( .A(n25964), .B(n25966), .Z(n26065) );
  NAND U34730 ( .A(n26066), .B(n26067), .Z(n25966) );
  OR U34731 ( .A(n26068), .B(n26069), .Z(n26067) );
  OR U34732 ( .A(n26070), .B(n26071), .Z(n26066) );
  NAND U34733 ( .A(n26072), .B(n26073), .Z(n25964) );
  OR U34734 ( .A(n26074), .B(n26075), .Z(n26073) );
  OR U34735 ( .A(n26076), .B(n26077), .Z(n26072) );
  ANDN U34736 ( .B(n26078), .A(n26079), .Z(n25965) );
  IV U34737 ( .A(n26080), .Z(n26078) );
  XNOR U34738 ( .A(n26045), .B(n26044), .Z(N63088) );
  XOR U34739 ( .A(n26064), .B(n26063), .Z(n26044) );
  XNOR U34740 ( .A(n26079), .B(n26080), .Z(n26063) );
  XNOR U34741 ( .A(n26074), .B(n26075), .Z(n26080) );
  XNOR U34742 ( .A(n26076), .B(n26077), .Z(n26075) );
  XNOR U34743 ( .A(y[4621]), .B(x[4621]), .Z(n26077) );
  XNOR U34744 ( .A(y[4622]), .B(x[4622]), .Z(n26076) );
  XNOR U34745 ( .A(y[4620]), .B(x[4620]), .Z(n26074) );
  XNOR U34746 ( .A(n26068), .B(n26069), .Z(n26079) );
  XNOR U34747 ( .A(y[4617]), .B(x[4617]), .Z(n26069) );
  XNOR U34748 ( .A(n26070), .B(n26071), .Z(n26068) );
  XNOR U34749 ( .A(y[4618]), .B(x[4618]), .Z(n26071) );
  XNOR U34750 ( .A(y[4619]), .B(x[4619]), .Z(n26070) );
  XNOR U34751 ( .A(n26061), .B(n26060), .Z(n26064) );
  XNOR U34752 ( .A(n26056), .B(n26057), .Z(n26060) );
  XNOR U34753 ( .A(y[4614]), .B(x[4614]), .Z(n26057) );
  XNOR U34754 ( .A(n26058), .B(n26059), .Z(n26056) );
  XNOR U34755 ( .A(y[4615]), .B(x[4615]), .Z(n26059) );
  XNOR U34756 ( .A(y[4616]), .B(x[4616]), .Z(n26058) );
  XNOR U34757 ( .A(n26050), .B(n26051), .Z(n26061) );
  XNOR U34758 ( .A(y[4611]), .B(x[4611]), .Z(n26051) );
  XNOR U34759 ( .A(n26052), .B(n26053), .Z(n26050) );
  XNOR U34760 ( .A(y[4612]), .B(x[4612]), .Z(n26053) );
  XNOR U34761 ( .A(y[4613]), .B(x[4613]), .Z(n26052) );
  XOR U34762 ( .A(n26026), .B(n26027), .Z(n26045) );
  XNOR U34763 ( .A(n26042), .B(n26043), .Z(n26027) );
  XNOR U34764 ( .A(n26037), .B(n26038), .Z(n26043) );
  XNOR U34765 ( .A(n26039), .B(n26040), .Z(n26038) );
  XNOR U34766 ( .A(y[4609]), .B(x[4609]), .Z(n26040) );
  XNOR U34767 ( .A(y[4610]), .B(x[4610]), .Z(n26039) );
  XNOR U34768 ( .A(y[4608]), .B(x[4608]), .Z(n26037) );
  XNOR U34769 ( .A(n26031), .B(n26032), .Z(n26042) );
  XNOR U34770 ( .A(y[4605]), .B(x[4605]), .Z(n26032) );
  XNOR U34771 ( .A(n26033), .B(n26034), .Z(n26031) );
  XNOR U34772 ( .A(y[4606]), .B(x[4606]), .Z(n26034) );
  XNOR U34773 ( .A(y[4607]), .B(x[4607]), .Z(n26033) );
  XOR U34774 ( .A(n26025), .B(n26024), .Z(n26026) );
  XNOR U34775 ( .A(n26020), .B(n26021), .Z(n26024) );
  XNOR U34776 ( .A(y[4602]), .B(x[4602]), .Z(n26021) );
  XNOR U34777 ( .A(n26022), .B(n26023), .Z(n26020) );
  XNOR U34778 ( .A(y[4603]), .B(x[4603]), .Z(n26023) );
  XNOR U34779 ( .A(y[4604]), .B(x[4604]), .Z(n26022) );
  XNOR U34780 ( .A(n26014), .B(n26015), .Z(n26025) );
  XNOR U34781 ( .A(y[4599]), .B(x[4599]), .Z(n26015) );
  XNOR U34782 ( .A(n26016), .B(n26017), .Z(n26014) );
  XNOR U34783 ( .A(y[4600]), .B(x[4600]), .Z(n26017) );
  XNOR U34784 ( .A(y[4601]), .B(x[4601]), .Z(n26016) );
  NAND U34785 ( .A(n26081), .B(n26082), .Z(N63079) );
  NANDN U34786 ( .A(n26083), .B(n26084), .Z(n26082) );
  OR U34787 ( .A(n26085), .B(n26086), .Z(n26084) );
  NAND U34788 ( .A(n26085), .B(n26086), .Z(n26081) );
  XOR U34789 ( .A(n26085), .B(n26087), .Z(N63078) );
  XNOR U34790 ( .A(n26083), .B(n26086), .Z(n26087) );
  AND U34791 ( .A(n26088), .B(n26089), .Z(n26086) );
  NANDN U34792 ( .A(n26090), .B(n26091), .Z(n26089) );
  NANDN U34793 ( .A(n26092), .B(n26093), .Z(n26091) );
  NANDN U34794 ( .A(n26093), .B(n26092), .Z(n26088) );
  NAND U34795 ( .A(n26094), .B(n26095), .Z(n26083) );
  NANDN U34796 ( .A(n26096), .B(n26097), .Z(n26095) );
  OR U34797 ( .A(n26098), .B(n26099), .Z(n26097) );
  NAND U34798 ( .A(n26099), .B(n26098), .Z(n26094) );
  AND U34799 ( .A(n26100), .B(n26101), .Z(n26085) );
  NANDN U34800 ( .A(n26102), .B(n26103), .Z(n26101) );
  NANDN U34801 ( .A(n26104), .B(n26105), .Z(n26103) );
  NANDN U34802 ( .A(n26105), .B(n26104), .Z(n26100) );
  XOR U34803 ( .A(n26099), .B(n26106), .Z(N63077) );
  XOR U34804 ( .A(n26096), .B(n26098), .Z(n26106) );
  XNOR U34805 ( .A(n26092), .B(n26107), .Z(n26098) );
  XNOR U34806 ( .A(n26090), .B(n26093), .Z(n26107) );
  NAND U34807 ( .A(n26108), .B(n26109), .Z(n26093) );
  NAND U34808 ( .A(n26110), .B(n26111), .Z(n26109) );
  OR U34809 ( .A(n26112), .B(n26113), .Z(n26110) );
  NANDN U34810 ( .A(n26114), .B(n26112), .Z(n26108) );
  IV U34811 ( .A(n26113), .Z(n26114) );
  NAND U34812 ( .A(n26115), .B(n26116), .Z(n26090) );
  NAND U34813 ( .A(n26117), .B(n26118), .Z(n26116) );
  NANDN U34814 ( .A(n26119), .B(n26120), .Z(n26117) );
  NANDN U34815 ( .A(n26120), .B(n26119), .Z(n26115) );
  AND U34816 ( .A(n26121), .B(n26122), .Z(n26092) );
  NAND U34817 ( .A(n26123), .B(n26124), .Z(n26122) );
  OR U34818 ( .A(n26125), .B(n26126), .Z(n26123) );
  NANDN U34819 ( .A(n26127), .B(n26125), .Z(n26121) );
  NAND U34820 ( .A(n26128), .B(n26129), .Z(n26096) );
  NANDN U34821 ( .A(n26130), .B(n26131), .Z(n26129) );
  OR U34822 ( .A(n26132), .B(n26133), .Z(n26131) );
  NANDN U34823 ( .A(n26134), .B(n26132), .Z(n26128) );
  IV U34824 ( .A(n26133), .Z(n26134) );
  XNOR U34825 ( .A(n26104), .B(n26135), .Z(n26099) );
  XNOR U34826 ( .A(n26102), .B(n26105), .Z(n26135) );
  NAND U34827 ( .A(n26136), .B(n26137), .Z(n26105) );
  NAND U34828 ( .A(n26138), .B(n26139), .Z(n26137) );
  OR U34829 ( .A(n26140), .B(n26141), .Z(n26138) );
  NANDN U34830 ( .A(n26142), .B(n26140), .Z(n26136) );
  IV U34831 ( .A(n26141), .Z(n26142) );
  NAND U34832 ( .A(n26143), .B(n26144), .Z(n26102) );
  NAND U34833 ( .A(n26145), .B(n26146), .Z(n26144) );
  NANDN U34834 ( .A(n26147), .B(n26148), .Z(n26145) );
  NANDN U34835 ( .A(n26148), .B(n26147), .Z(n26143) );
  AND U34836 ( .A(n26149), .B(n26150), .Z(n26104) );
  NAND U34837 ( .A(n26151), .B(n26152), .Z(n26150) );
  OR U34838 ( .A(n26153), .B(n26154), .Z(n26151) );
  NANDN U34839 ( .A(n26155), .B(n26153), .Z(n26149) );
  XNOR U34840 ( .A(n26130), .B(n26156), .Z(N63076) );
  XOR U34841 ( .A(n26132), .B(n26133), .Z(n26156) );
  XNOR U34842 ( .A(n26146), .B(n26157), .Z(n26133) );
  XOR U34843 ( .A(n26147), .B(n26148), .Z(n26157) );
  XOR U34844 ( .A(n26153), .B(n26158), .Z(n26148) );
  XOR U34845 ( .A(n26152), .B(n26155), .Z(n26158) );
  IV U34846 ( .A(n26154), .Z(n26155) );
  NAND U34847 ( .A(n26159), .B(n26160), .Z(n26154) );
  OR U34848 ( .A(n26161), .B(n26162), .Z(n26160) );
  OR U34849 ( .A(n26163), .B(n26164), .Z(n26159) );
  NAND U34850 ( .A(n26165), .B(n26166), .Z(n26152) );
  OR U34851 ( .A(n26167), .B(n26168), .Z(n26166) );
  OR U34852 ( .A(n26169), .B(n26170), .Z(n26165) );
  NOR U34853 ( .A(n26171), .B(n26172), .Z(n26153) );
  ANDN U34854 ( .B(n26173), .A(n26174), .Z(n26147) );
  XNOR U34855 ( .A(n26140), .B(n26175), .Z(n26146) );
  XNOR U34856 ( .A(n26139), .B(n26141), .Z(n26175) );
  NAND U34857 ( .A(n26176), .B(n26177), .Z(n26141) );
  OR U34858 ( .A(n26178), .B(n26179), .Z(n26177) );
  OR U34859 ( .A(n26180), .B(n26181), .Z(n26176) );
  NAND U34860 ( .A(n26182), .B(n26183), .Z(n26139) );
  OR U34861 ( .A(n26184), .B(n26185), .Z(n26183) );
  OR U34862 ( .A(n26186), .B(n26187), .Z(n26182) );
  ANDN U34863 ( .B(n26188), .A(n26189), .Z(n26140) );
  IV U34864 ( .A(n26190), .Z(n26188) );
  ANDN U34865 ( .B(n26191), .A(n26192), .Z(n26132) );
  XOR U34866 ( .A(n26118), .B(n26193), .Z(n26130) );
  XOR U34867 ( .A(n26119), .B(n26120), .Z(n26193) );
  XOR U34868 ( .A(n26125), .B(n26194), .Z(n26120) );
  XOR U34869 ( .A(n26124), .B(n26127), .Z(n26194) );
  IV U34870 ( .A(n26126), .Z(n26127) );
  NAND U34871 ( .A(n26195), .B(n26196), .Z(n26126) );
  OR U34872 ( .A(n26197), .B(n26198), .Z(n26196) );
  OR U34873 ( .A(n26199), .B(n26200), .Z(n26195) );
  NAND U34874 ( .A(n26201), .B(n26202), .Z(n26124) );
  OR U34875 ( .A(n26203), .B(n26204), .Z(n26202) );
  OR U34876 ( .A(n26205), .B(n26206), .Z(n26201) );
  NOR U34877 ( .A(n26207), .B(n26208), .Z(n26125) );
  ANDN U34878 ( .B(n26209), .A(n26210), .Z(n26119) );
  IV U34879 ( .A(n26211), .Z(n26209) );
  XNOR U34880 ( .A(n26112), .B(n26212), .Z(n26118) );
  XNOR U34881 ( .A(n26111), .B(n26113), .Z(n26212) );
  NAND U34882 ( .A(n26213), .B(n26214), .Z(n26113) );
  OR U34883 ( .A(n26215), .B(n26216), .Z(n26214) );
  OR U34884 ( .A(n26217), .B(n26218), .Z(n26213) );
  NAND U34885 ( .A(n26219), .B(n26220), .Z(n26111) );
  OR U34886 ( .A(n26221), .B(n26222), .Z(n26220) );
  OR U34887 ( .A(n26223), .B(n26224), .Z(n26219) );
  ANDN U34888 ( .B(n26225), .A(n26226), .Z(n26112) );
  IV U34889 ( .A(n26227), .Z(n26225) );
  XNOR U34890 ( .A(n26192), .B(n26191), .Z(N63075) );
  XOR U34891 ( .A(n26211), .B(n26210), .Z(n26191) );
  XNOR U34892 ( .A(n26226), .B(n26227), .Z(n26210) );
  XNOR U34893 ( .A(n26221), .B(n26222), .Z(n26227) );
  XNOR U34894 ( .A(n26223), .B(n26224), .Z(n26222) );
  XNOR U34895 ( .A(y[4597]), .B(x[4597]), .Z(n26224) );
  XNOR U34896 ( .A(y[4598]), .B(x[4598]), .Z(n26223) );
  XNOR U34897 ( .A(y[4596]), .B(x[4596]), .Z(n26221) );
  XNOR U34898 ( .A(n26215), .B(n26216), .Z(n26226) );
  XNOR U34899 ( .A(y[4593]), .B(x[4593]), .Z(n26216) );
  XNOR U34900 ( .A(n26217), .B(n26218), .Z(n26215) );
  XNOR U34901 ( .A(y[4594]), .B(x[4594]), .Z(n26218) );
  XNOR U34902 ( .A(y[4595]), .B(x[4595]), .Z(n26217) );
  XNOR U34903 ( .A(n26208), .B(n26207), .Z(n26211) );
  XNOR U34904 ( .A(n26203), .B(n26204), .Z(n26207) );
  XNOR U34905 ( .A(y[4590]), .B(x[4590]), .Z(n26204) );
  XNOR U34906 ( .A(n26205), .B(n26206), .Z(n26203) );
  XNOR U34907 ( .A(y[4591]), .B(x[4591]), .Z(n26206) );
  XNOR U34908 ( .A(y[4592]), .B(x[4592]), .Z(n26205) );
  XNOR U34909 ( .A(n26197), .B(n26198), .Z(n26208) );
  XNOR U34910 ( .A(y[4587]), .B(x[4587]), .Z(n26198) );
  XNOR U34911 ( .A(n26199), .B(n26200), .Z(n26197) );
  XNOR U34912 ( .A(y[4588]), .B(x[4588]), .Z(n26200) );
  XNOR U34913 ( .A(y[4589]), .B(x[4589]), .Z(n26199) );
  XOR U34914 ( .A(n26173), .B(n26174), .Z(n26192) );
  XNOR U34915 ( .A(n26189), .B(n26190), .Z(n26174) );
  XNOR U34916 ( .A(n26184), .B(n26185), .Z(n26190) );
  XNOR U34917 ( .A(n26186), .B(n26187), .Z(n26185) );
  XNOR U34918 ( .A(y[4585]), .B(x[4585]), .Z(n26187) );
  XNOR U34919 ( .A(y[4586]), .B(x[4586]), .Z(n26186) );
  XNOR U34920 ( .A(y[4584]), .B(x[4584]), .Z(n26184) );
  XNOR U34921 ( .A(n26178), .B(n26179), .Z(n26189) );
  XNOR U34922 ( .A(y[4581]), .B(x[4581]), .Z(n26179) );
  XNOR U34923 ( .A(n26180), .B(n26181), .Z(n26178) );
  XNOR U34924 ( .A(y[4582]), .B(x[4582]), .Z(n26181) );
  XNOR U34925 ( .A(y[4583]), .B(x[4583]), .Z(n26180) );
  XOR U34926 ( .A(n26172), .B(n26171), .Z(n26173) );
  XNOR U34927 ( .A(n26167), .B(n26168), .Z(n26171) );
  XNOR U34928 ( .A(y[4578]), .B(x[4578]), .Z(n26168) );
  XNOR U34929 ( .A(n26169), .B(n26170), .Z(n26167) );
  XNOR U34930 ( .A(y[4579]), .B(x[4579]), .Z(n26170) );
  XNOR U34931 ( .A(y[4580]), .B(x[4580]), .Z(n26169) );
  XNOR U34932 ( .A(n26161), .B(n26162), .Z(n26172) );
  XNOR U34933 ( .A(y[4575]), .B(x[4575]), .Z(n26162) );
  XNOR U34934 ( .A(n26163), .B(n26164), .Z(n26161) );
  XNOR U34935 ( .A(y[4576]), .B(x[4576]), .Z(n26164) );
  XNOR U34936 ( .A(y[4577]), .B(x[4577]), .Z(n26163) );
  NAND U34937 ( .A(n26228), .B(n26229), .Z(N63066) );
  NANDN U34938 ( .A(n26230), .B(n26231), .Z(n26229) );
  OR U34939 ( .A(n26232), .B(n26233), .Z(n26231) );
  NAND U34940 ( .A(n26232), .B(n26233), .Z(n26228) );
  XOR U34941 ( .A(n26232), .B(n26234), .Z(N63065) );
  XNOR U34942 ( .A(n26230), .B(n26233), .Z(n26234) );
  AND U34943 ( .A(n26235), .B(n26236), .Z(n26233) );
  NANDN U34944 ( .A(n26237), .B(n26238), .Z(n26236) );
  NANDN U34945 ( .A(n26239), .B(n26240), .Z(n26238) );
  NANDN U34946 ( .A(n26240), .B(n26239), .Z(n26235) );
  NAND U34947 ( .A(n26241), .B(n26242), .Z(n26230) );
  NANDN U34948 ( .A(n26243), .B(n26244), .Z(n26242) );
  OR U34949 ( .A(n26245), .B(n26246), .Z(n26244) );
  NAND U34950 ( .A(n26246), .B(n26245), .Z(n26241) );
  AND U34951 ( .A(n26247), .B(n26248), .Z(n26232) );
  NANDN U34952 ( .A(n26249), .B(n26250), .Z(n26248) );
  NANDN U34953 ( .A(n26251), .B(n26252), .Z(n26250) );
  NANDN U34954 ( .A(n26252), .B(n26251), .Z(n26247) );
  XOR U34955 ( .A(n26246), .B(n26253), .Z(N63064) );
  XOR U34956 ( .A(n26243), .B(n26245), .Z(n26253) );
  XNOR U34957 ( .A(n26239), .B(n26254), .Z(n26245) );
  XNOR U34958 ( .A(n26237), .B(n26240), .Z(n26254) );
  NAND U34959 ( .A(n26255), .B(n26256), .Z(n26240) );
  NAND U34960 ( .A(n26257), .B(n26258), .Z(n26256) );
  OR U34961 ( .A(n26259), .B(n26260), .Z(n26257) );
  NANDN U34962 ( .A(n26261), .B(n26259), .Z(n26255) );
  IV U34963 ( .A(n26260), .Z(n26261) );
  NAND U34964 ( .A(n26262), .B(n26263), .Z(n26237) );
  NAND U34965 ( .A(n26264), .B(n26265), .Z(n26263) );
  NANDN U34966 ( .A(n26266), .B(n26267), .Z(n26264) );
  NANDN U34967 ( .A(n26267), .B(n26266), .Z(n26262) );
  AND U34968 ( .A(n26268), .B(n26269), .Z(n26239) );
  NAND U34969 ( .A(n26270), .B(n26271), .Z(n26269) );
  OR U34970 ( .A(n26272), .B(n26273), .Z(n26270) );
  NANDN U34971 ( .A(n26274), .B(n26272), .Z(n26268) );
  NAND U34972 ( .A(n26275), .B(n26276), .Z(n26243) );
  NANDN U34973 ( .A(n26277), .B(n26278), .Z(n26276) );
  OR U34974 ( .A(n26279), .B(n26280), .Z(n26278) );
  NANDN U34975 ( .A(n26281), .B(n26279), .Z(n26275) );
  IV U34976 ( .A(n26280), .Z(n26281) );
  XNOR U34977 ( .A(n26251), .B(n26282), .Z(n26246) );
  XNOR U34978 ( .A(n26249), .B(n26252), .Z(n26282) );
  NAND U34979 ( .A(n26283), .B(n26284), .Z(n26252) );
  NAND U34980 ( .A(n26285), .B(n26286), .Z(n26284) );
  OR U34981 ( .A(n26287), .B(n26288), .Z(n26285) );
  NANDN U34982 ( .A(n26289), .B(n26287), .Z(n26283) );
  IV U34983 ( .A(n26288), .Z(n26289) );
  NAND U34984 ( .A(n26290), .B(n26291), .Z(n26249) );
  NAND U34985 ( .A(n26292), .B(n26293), .Z(n26291) );
  NANDN U34986 ( .A(n26294), .B(n26295), .Z(n26292) );
  NANDN U34987 ( .A(n26295), .B(n26294), .Z(n26290) );
  AND U34988 ( .A(n26296), .B(n26297), .Z(n26251) );
  NAND U34989 ( .A(n26298), .B(n26299), .Z(n26297) );
  OR U34990 ( .A(n26300), .B(n26301), .Z(n26298) );
  NANDN U34991 ( .A(n26302), .B(n26300), .Z(n26296) );
  XNOR U34992 ( .A(n26277), .B(n26303), .Z(N63063) );
  XOR U34993 ( .A(n26279), .B(n26280), .Z(n26303) );
  XNOR U34994 ( .A(n26293), .B(n26304), .Z(n26280) );
  XOR U34995 ( .A(n26294), .B(n26295), .Z(n26304) );
  XOR U34996 ( .A(n26300), .B(n26305), .Z(n26295) );
  XOR U34997 ( .A(n26299), .B(n26302), .Z(n26305) );
  IV U34998 ( .A(n26301), .Z(n26302) );
  NAND U34999 ( .A(n26306), .B(n26307), .Z(n26301) );
  OR U35000 ( .A(n26308), .B(n26309), .Z(n26307) );
  OR U35001 ( .A(n26310), .B(n26311), .Z(n26306) );
  NAND U35002 ( .A(n26312), .B(n26313), .Z(n26299) );
  OR U35003 ( .A(n26314), .B(n26315), .Z(n26313) );
  OR U35004 ( .A(n26316), .B(n26317), .Z(n26312) );
  NOR U35005 ( .A(n26318), .B(n26319), .Z(n26300) );
  ANDN U35006 ( .B(n26320), .A(n26321), .Z(n26294) );
  XNOR U35007 ( .A(n26287), .B(n26322), .Z(n26293) );
  XNOR U35008 ( .A(n26286), .B(n26288), .Z(n26322) );
  NAND U35009 ( .A(n26323), .B(n26324), .Z(n26288) );
  OR U35010 ( .A(n26325), .B(n26326), .Z(n26324) );
  OR U35011 ( .A(n26327), .B(n26328), .Z(n26323) );
  NAND U35012 ( .A(n26329), .B(n26330), .Z(n26286) );
  OR U35013 ( .A(n26331), .B(n26332), .Z(n26330) );
  OR U35014 ( .A(n26333), .B(n26334), .Z(n26329) );
  ANDN U35015 ( .B(n26335), .A(n26336), .Z(n26287) );
  IV U35016 ( .A(n26337), .Z(n26335) );
  ANDN U35017 ( .B(n26338), .A(n26339), .Z(n26279) );
  XOR U35018 ( .A(n26265), .B(n26340), .Z(n26277) );
  XOR U35019 ( .A(n26266), .B(n26267), .Z(n26340) );
  XOR U35020 ( .A(n26272), .B(n26341), .Z(n26267) );
  XOR U35021 ( .A(n26271), .B(n26274), .Z(n26341) );
  IV U35022 ( .A(n26273), .Z(n26274) );
  NAND U35023 ( .A(n26342), .B(n26343), .Z(n26273) );
  OR U35024 ( .A(n26344), .B(n26345), .Z(n26343) );
  OR U35025 ( .A(n26346), .B(n26347), .Z(n26342) );
  NAND U35026 ( .A(n26348), .B(n26349), .Z(n26271) );
  OR U35027 ( .A(n26350), .B(n26351), .Z(n26349) );
  OR U35028 ( .A(n26352), .B(n26353), .Z(n26348) );
  NOR U35029 ( .A(n26354), .B(n26355), .Z(n26272) );
  ANDN U35030 ( .B(n26356), .A(n26357), .Z(n26266) );
  IV U35031 ( .A(n26358), .Z(n26356) );
  XNOR U35032 ( .A(n26259), .B(n26359), .Z(n26265) );
  XNOR U35033 ( .A(n26258), .B(n26260), .Z(n26359) );
  NAND U35034 ( .A(n26360), .B(n26361), .Z(n26260) );
  OR U35035 ( .A(n26362), .B(n26363), .Z(n26361) );
  OR U35036 ( .A(n26364), .B(n26365), .Z(n26360) );
  NAND U35037 ( .A(n26366), .B(n26367), .Z(n26258) );
  OR U35038 ( .A(n26368), .B(n26369), .Z(n26367) );
  OR U35039 ( .A(n26370), .B(n26371), .Z(n26366) );
  ANDN U35040 ( .B(n26372), .A(n26373), .Z(n26259) );
  IV U35041 ( .A(n26374), .Z(n26372) );
  XNOR U35042 ( .A(n26339), .B(n26338), .Z(N63062) );
  XOR U35043 ( .A(n26358), .B(n26357), .Z(n26338) );
  XNOR U35044 ( .A(n26373), .B(n26374), .Z(n26357) );
  XNOR U35045 ( .A(n26368), .B(n26369), .Z(n26374) );
  XNOR U35046 ( .A(n26370), .B(n26371), .Z(n26369) );
  XNOR U35047 ( .A(y[4573]), .B(x[4573]), .Z(n26371) );
  XNOR U35048 ( .A(y[4574]), .B(x[4574]), .Z(n26370) );
  XNOR U35049 ( .A(y[4572]), .B(x[4572]), .Z(n26368) );
  XNOR U35050 ( .A(n26362), .B(n26363), .Z(n26373) );
  XNOR U35051 ( .A(y[4569]), .B(x[4569]), .Z(n26363) );
  XNOR U35052 ( .A(n26364), .B(n26365), .Z(n26362) );
  XNOR U35053 ( .A(y[4570]), .B(x[4570]), .Z(n26365) );
  XNOR U35054 ( .A(y[4571]), .B(x[4571]), .Z(n26364) );
  XNOR U35055 ( .A(n26355), .B(n26354), .Z(n26358) );
  XNOR U35056 ( .A(n26350), .B(n26351), .Z(n26354) );
  XNOR U35057 ( .A(y[4566]), .B(x[4566]), .Z(n26351) );
  XNOR U35058 ( .A(n26352), .B(n26353), .Z(n26350) );
  XNOR U35059 ( .A(y[4567]), .B(x[4567]), .Z(n26353) );
  XNOR U35060 ( .A(y[4568]), .B(x[4568]), .Z(n26352) );
  XNOR U35061 ( .A(n26344), .B(n26345), .Z(n26355) );
  XNOR U35062 ( .A(y[4563]), .B(x[4563]), .Z(n26345) );
  XNOR U35063 ( .A(n26346), .B(n26347), .Z(n26344) );
  XNOR U35064 ( .A(y[4564]), .B(x[4564]), .Z(n26347) );
  XNOR U35065 ( .A(y[4565]), .B(x[4565]), .Z(n26346) );
  XOR U35066 ( .A(n26320), .B(n26321), .Z(n26339) );
  XNOR U35067 ( .A(n26336), .B(n26337), .Z(n26321) );
  XNOR U35068 ( .A(n26331), .B(n26332), .Z(n26337) );
  XNOR U35069 ( .A(n26333), .B(n26334), .Z(n26332) );
  XNOR U35070 ( .A(y[4561]), .B(x[4561]), .Z(n26334) );
  XNOR U35071 ( .A(y[4562]), .B(x[4562]), .Z(n26333) );
  XNOR U35072 ( .A(y[4560]), .B(x[4560]), .Z(n26331) );
  XNOR U35073 ( .A(n26325), .B(n26326), .Z(n26336) );
  XNOR U35074 ( .A(y[4557]), .B(x[4557]), .Z(n26326) );
  XNOR U35075 ( .A(n26327), .B(n26328), .Z(n26325) );
  XNOR U35076 ( .A(y[4558]), .B(x[4558]), .Z(n26328) );
  XNOR U35077 ( .A(y[4559]), .B(x[4559]), .Z(n26327) );
  XOR U35078 ( .A(n26319), .B(n26318), .Z(n26320) );
  XNOR U35079 ( .A(n26314), .B(n26315), .Z(n26318) );
  XNOR U35080 ( .A(y[4554]), .B(x[4554]), .Z(n26315) );
  XNOR U35081 ( .A(n26316), .B(n26317), .Z(n26314) );
  XNOR U35082 ( .A(y[4555]), .B(x[4555]), .Z(n26317) );
  XNOR U35083 ( .A(y[4556]), .B(x[4556]), .Z(n26316) );
  XNOR U35084 ( .A(n26308), .B(n26309), .Z(n26319) );
  XNOR U35085 ( .A(y[4551]), .B(x[4551]), .Z(n26309) );
  XNOR U35086 ( .A(n26310), .B(n26311), .Z(n26308) );
  XNOR U35087 ( .A(y[4552]), .B(x[4552]), .Z(n26311) );
  XNOR U35088 ( .A(y[4553]), .B(x[4553]), .Z(n26310) );
  NAND U35089 ( .A(n26375), .B(n26376), .Z(N63053) );
  NANDN U35090 ( .A(n26377), .B(n26378), .Z(n26376) );
  OR U35091 ( .A(n26379), .B(n26380), .Z(n26378) );
  NAND U35092 ( .A(n26379), .B(n26380), .Z(n26375) );
  XOR U35093 ( .A(n26379), .B(n26381), .Z(N63052) );
  XNOR U35094 ( .A(n26377), .B(n26380), .Z(n26381) );
  AND U35095 ( .A(n26382), .B(n26383), .Z(n26380) );
  NANDN U35096 ( .A(n26384), .B(n26385), .Z(n26383) );
  NANDN U35097 ( .A(n26386), .B(n26387), .Z(n26385) );
  NANDN U35098 ( .A(n26387), .B(n26386), .Z(n26382) );
  NAND U35099 ( .A(n26388), .B(n26389), .Z(n26377) );
  NANDN U35100 ( .A(n26390), .B(n26391), .Z(n26389) );
  OR U35101 ( .A(n26392), .B(n26393), .Z(n26391) );
  NAND U35102 ( .A(n26393), .B(n26392), .Z(n26388) );
  AND U35103 ( .A(n26394), .B(n26395), .Z(n26379) );
  NANDN U35104 ( .A(n26396), .B(n26397), .Z(n26395) );
  NANDN U35105 ( .A(n26398), .B(n26399), .Z(n26397) );
  NANDN U35106 ( .A(n26399), .B(n26398), .Z(n26394) );
  XOR U35107 ( .A(n26393), .B(n26400), .Z(N63051) );
  XOR U35108 ( .A(n26390), .B(n26392), .Z(n26400) );
  XNOR U35109 ( .A(n26386), .B(n26401), .Z(n26392) );
  XNOR U35110 ( .A(n26384), .B(n26387), .Z(n26401) );
  NAND U35111 ( .A(n26402), .B(n26403), .Z(n26387) );
  NAND U35112 ( .A(n26404), .B(n26405), .Z(n26403) );
  OR U35113 ( .A(n26406), .B(n26407), .Z(n26404) );
  NANDN U35114 ( .A(n26408), .B(n26406), .Z(n26402) );
  IV U35115 ( .A(n26407), .Z(n26408) );
  NAND U35116 ( .A(n26409), .B(n26410), .Z(n26384) );
  NAND U35117 ( .A(n26411), .B(n26412), .Z(n26410) );
  NANDN U35118 ( .A(n26413), .B(n26414), .Z(n26411) );
  NANDN U35119 ( .A(n26414), .B(n26413), .Z(n26409) );
  AND U35120 ( .A(n26415), .B(n26416), .Z(n26386) );
  NAND U35121 ( .A(n26417), .B(n26418), .Z(n26416) );
  OR U35122 ( .A(n26419), .B(n26420), .Z(n26417) );
  NANDN U35123 ( .A(n26421), .B(n26419), .Z(n26415) );
  NAND U35124 ( .A(n26422), .B(n26423), .Z(n26390) );
  NANDN U35125 ( .A(n26424), .B(n26425), .Z(n26423) );
  OR U35126 ( .A(n26426), .B(n26427), .Z(n26425) );
  NANDN U35127 ( .A(n26428), .B(n26426), .Z(n26422) );
  IV U35128 ( .A(n26427), .Z(n26428) );
  XNOR U35129 ( .A(n26398), .B(n26429), .Z(n26393) );
  XNOR U35130 ( .A(n26396), .B(n26399), .Z(n26429) );
  NAND U35131 ( .A(n26430), .B(n26431), .Z(n26399) );
  NAND U35132 ( .A(n26432), .B(n26433), .Z(n26431) );
  OR U35133 ( .A(n26434), .B(n26435), .Z(n26432) );
  NANDN U35134 ( .A(n26436), .B(n26434), .Z(n26430) );
  IV U35135 ( .A(n26435), .Z(n26436) );
  NAND U35136 ( .A(n26437), .B(n26438), .Z(n26396) );
  NAND U35137 ( .A(n26439), .B(n26440), .Z(n26438) );
  NANDN U35138 ( .A(n26441), .B(n26442), .Z(n26439) );
  NANDN U35139 ( .A(n26442), .B(n26441), .Z(n26437) );
  AND U35140 ( .A(n26443), .B(n26444), .Z(n26398) );
  NAND U35141 ( .A(n26445), .B(n26446), .Z(n26444) );
  OR U35142 ( .A(n26447), .B(n26448), .Z(n26445) );
  NANDN U35143 ( .A(n26449), .B(n26447), .Z(n26443) );
  XNOR U35144 ( .A(n26424), .B(n26450), .Z(N63050) );
  XOR U35145 ( .A(n26426), .B(n26427), .Z(n26450) );
  XNOR U35146 ( .A(n26440), .B(n26451), .Z(n26427) );
  XOR U35147 ( .A(n26441), .B(n26442), .Z(n26451) );
  XOR U35148 ( .A(n26447), .B(n26452), .Z(n26442) );
  XOR U35149 ( .A(n26446), .B(n26449), .Z(n26452) );
  IV U35150 ( .A(n26448), .Z(n26449) );
  NAND U35151 ( .A(n26453), .B(n26454), .Z(n26448) );
  OR U35152 ( .A(n26455), .B(n26456), .Z(n26454) );
  OR U35153 ( .A(n26457), .B(n26458), .Z(n26453) );
  NAND U35154 ( .A(n26459), .B(n26460), .Z(n26446) );
  OR U35155 ( .A(n26461), .B(n26462), .Z(n26460) );
  OR U35156 ( .A(n26463), .B(n26464), .Z(n26459) );
  NOR U35157 ( .A(n26465), .B(n26466), .Z(n26447) );
  ANDN U35158 ( .B(n26467), .A(n26468), .Z(n26441) );
  XNOR U35159 ( .A(n26434), .B(n26469), .Z(n26440) );
  XNOR U35160 ( .A(n26433), .B(n26435), .Z(n26469) );
  NAND U35161 ( .A(n26470), .B(n26471), .Z(n26435) );
  OR U35162 ( .A(n26472), .B(n26473), .Z(n26471) );
  OR U35163 ( .A(n26474), .B(n26475), .Z(n26470) );
  NAND U35164 ( .A(n26476), .B(n26477), .Z(n26433) );
  OR U35165 ( .A(n26478), .B(n26479), .Z(n26477) );
  OR U35166 ( .A(n26480), .B(n26481), .Z(n26476) );
  ANDN U35167 ( .B(n26482), .A(n26483), .Z(n26434) );
  IV U35168 ( .A(n26484), .Z(n26482) );
  ANDN U35169 ( .B(n26485), .A(n26486), .Z(n26426) );
  XOR U35170 ( .A(n26412), .B(n26487), .Z(n26424) );
  XOR U35171 ( .A(n26413), .B(n26414), .Z(n26487) );
  XOR U35172 ( .A(n26419), .B(n26488), .Z(n26414) );
  XOR U35173 ( .A(n26418), .B(n26421), .Z(n26488) );
  IV U35174 ( .A(n26420), .Z(n26421) );
  NAND U35175 ( .A(n26489), .B(n26490), .Z(n26420) );
  OR U35176 ( .A(n26491), .B(n26492), .Z(n26490) );
  OR U35177 ( .A(n26493), .B(n26494), .Z(n26489) );
  NAND U35178 ( .A(n26495), .B(n26496), .Z(n26418) );
  OR U35179 ( .A(n26497), .B(n26498), .Z(n26496) );
  OR U35180 ( .A(n26499), .B(n26500), .Z(n26495) );
  NOR U35181 ( .A(n26501), .B(n26502), .Z(n26419) );
  ANDN U35182 ( .B(n26503), .A(n26504), .Z(n26413) );
  IV U35183 ( .A(n26505), .Z(n26503) );
  XNOR U35184 ( .A(n26406), .B(n26506), .Z(n26412) );
  XNOR U35185 ( .A(n26405), .B(n26407), .Z(n26506) );
  NAND U35186 ( .A(n26507), .B(n26508), .Z(n26407) );
  OR U35187 ( .A(n26509), .B(n26510), .Z(n26508) );
  OR U35188 ( .A(n26511), .B(n26512), .Z(n26507) );
  NAND U35189 ( .A(n26513), .B(n26514), .Z(n26405) );
  OR U35190 ( .A(n26515), .B(n26516), .Z(n26514) );
  OR U35191 ( .A(n26517), .B(n26518), .Z(n26513) );
  ANDN U35192 ( .B(n26519), .A(n26520), .Z(n26406) );
  IV U35193 ( .A(n26521), .Z(n26519) );
  XNOR U35194 ( .A(n26486), .B(n26485), .Z(N63049) );
  XOR U35195 ( .A(n26505), .B(n26504), .Z(n26485) );
  XNOR U35196 ( .A(n26520), .B(n26521), .Z(n26504) );
  XNOR U35197 ( .A(n26515), .B(n26516), .Z(n26521) );
  XNOR U35198 ( .A(n26517), .B(n26518), .Z(n26516) );
  XNOR U35199 ( .A(y[4549]), .B(x[4549]), .Z(n26518) );
  XNOR U35200 ( .A(y[4550]), .B(x[4550]), .Z(n26517) );
  XNOR U35201 ( .A(y[4548]), .B(x[4548]), .Z(n26515) );
  XNOR U35202 ( .A(n26509), .B(n26510), .Z(n26520) );
  XNOR U35203 ( .A(y[4545]), .B(x[4545]), .Z(n26510) );
  XNOR U35204 ( .A(n26511), .B(n26512), .Z(n26509) );
  XNOR U35205 ( .A(y[4546]), .B(x[4546]), .Z(n26512) );
  XNOR U35206 ( .A(y[4547]), .B(x[4547]), .Z(n26511) );
  XNOR U35207 ( .A(n26502), .B(n26501), .Z(n26505) );
  XNOR U35208 ( .A(n26497), .B(n26498), .Z(n26501) );
  XNOR U35209 ( .A(y[4542]), .B(x[4542]), .Z(n26498) );
  XNOR U35210 ( .A(n26499), .B(n26500), .Z(n26497) );
  XNOR U35211 ( .A(y[4543]), .B(x[4543]), .Z(n26500) );
  XNOR U35212 ( .A(y[4544]), .B(x[4544]), .Z(n26499) );
  XNOR U35213 ( .A(n26491), .B(n26492), .Z(n26502) );
  XNOR U35214 ( .A(y[4539]), .B(x[4539]), .Z(n26492) );
  XNOR U35215 ( .A(n26493), .B(n26494), .Z(n26491) );
  XNOR U35216 ( .A(y[4540]), .B(x[4540]), .Z(n26494) );
  XNOR U35217 ( .A(y[4541]), .B(x[4541]), .Z(n26493) );
  XOR U35218 ( .A(n26467), .B(n26468), .Z(n26486) );
  XNOR U35219 ( .A(n26483), .B(n26484), .Z(n26468) );
  XNOR U35220 ( .A(n26478), .B(n26479), .Z(n26484) );
  XNOR U35221 ( .A(n26480), .B(n26481), .Z(n26479) );
  XNOR U35222 ( .A(y[4537]), .B(x[4537]), .Z(n26481) );
  XNOR U35223 ( .A(y[4538]), .B(x[4538]), .Z(n26480) );
  XNOR U35224 ( .A(y[4536]), .B(x[4536]), .Z(n26478) );
  XNOR U35225 ( .A(n26472), .B(n26473), .Z(n26483) );
  XNOR U35226 ( .A(y[4533]), .B(x[4533]), .Z(n26473) );
  XNOR U35227 ( .A(n26474), .B(n26475), .Z(n26472) );
  XNOR U35228 ( .A(y[4534]), .B(x[4534]), .Z(n26475) );
  XNOR U35229 ( .A(y[4535]), .B(x[4535]), .Z(n26474) );
  XOR U35230 ( .A(n26466), .B(n26465), .Z(n26467) );
  XNOR U35231 ( .A(n26461), .B(n26462), .Z(n26465) );
  XNOR U35232 ( .A(y[4530]), .B(x[4530]), .Z(n26462) );
  XNOR U35233 ( .A(n26463), .B(n26464), .Z(n26461) );
  XNOR U35234 ( .A(y[4531]), .B(x[4531]), .Z(n26464) );
  XNOR U35235 ( .A(y[4532]), .B(x[4532]), .Z(n26463) );
  XNOR U35236 ( .A(n26455), .B(n26456), .Z(n26466) );
  XNOR U35237 ( .A(y[4527]), .B(x[4527]), .Z(n26456) );
  XNOR U35238 ( .A(n26457), .B(n26458), .Z(n26455) );
  XNOR U35239 ( .A(y[4528]), .B(x[4528]), .Z(n26458) );
  XNOR U35240 ( .A(y[4529]), .B(x[4529]), .Z(n26457) );
  NAND U35241 ( .A(n26522), .B(n26523), .Z(N63040) );
  NANDN U35242 ( .A(n26524), .B(n26525), .Z(n26523) );
  OR U35243 ( .A(n26526), .B(n26527), .Z(n26525) );
  NAND U35244 ( .A(n26526), .B(n26527), .Z(n26522) );
  XOR U35245 ( .A(n26526), .B(n26528), .Z(N63039) );
  XNOR U35246 ( .A(n26524), .B(n26527), .Z(n26528) );
  AND U35247 ( .A(n26529), .B(n26530), .Z(n26527) );
  NANDN U35248 ( .A(n26531), .B(n26532), .Z(n26530) );
  NANDN U35249 ( .A(n26533), .B(n26534), .Z(n26532) );
  NANDN U35250 ( .A(n26534), .B(n26533), .Z(n26529) );
  NAND U35251 ( .A(n26535), .B(n26536), .Z(n26524) );
  NANDN U35252 ( .A(n26537), .B(n26538), .Z(n26536) );
  OR U35253 ( .A(n26539), .B(n26540), .Z(n26538) );
  NAND U35254 ( .A(n26540), .B(n26539), .Z(n26535) );
  AND U35255 ( .A(n26541), .B(n26542), .Z(n26526) );
  NANDN U35256 ( .A(n26543), .B(n26544), .Z(n26542) );
  NANDN U35257 ( .A(n26545), .B(n26546), .Z(n26544) );
  NANDN U35258 ( .A(n26546), .B(n26545), .Z(n26541) );
  XOR U35259 ( .A(n26540), .B(n26547), .Z(N63038) );
  XOR U35260 ( .A(n26537), .B(n26539), .Z(n26547) );
  XNOR U35261 ( .A(n26533), .B(n26548), .Z(n26539) );
  XNOR U35262 ( .A(n26531), .B(n26534), .Z(n26548) );
  NAND U35263 ( .A(n26549), .B(n26550), .Z(n26534) );
  NAND U35264 ( .A(n26551), .B(n26552), .Z(n26550) );
  OR U35265 ( .A(n26553), .B(n26554), .Z(n26551) );
  NANDN U35266 ( .A(n26555), .B(n26553), .Z(n26549) );
  IV U35267 ( .A(n26554), .Z(n26555) );
  NAND U35268 ( .A(n26556), .B(n26557), .Z(n26531) );
  NAND U35269 ( .A(n26558), .B(n26559), .Z(n26557) );
  NANDN U35270 ( .A(n26560), .B(n26561), .Z(n26558) );
  NANDN U35271 ( .A(n26561), .B(n26560), .Z(n26556) );
  AND U35272 ( .A(n26562), .B(n26563), .Z(n26533) );
  NAND U35273 ( .A(n26564), .B(n26565), .Z(n26563) );
  OR U35274 ( .A(n26566), .B(n26567), .Z(n26564) );
  NANDN U35275 ( .A(n26568), .B(n26566), .Z(n26562) );
  NAND U35276 ( .A(n26569), .B(n26570), .Z(n26537) );
  NANDN U35277 ( .A(n26571), .B(n26572), .Z(n26570) );
  OR U35278 ( .A(n26573), .B(n26574), .Z(n26572) );
  NANDN U35279 ( .A(n26575), .B(n26573), .Z(n26569) );
  IV U35280 ( .A(n26574), .Z(n26575) );
  XNOR U35281 ( .A(n26545), .B(n26576), .Z(n26540) );
  XNOR U35282 ( .A(n26543), .B(n26546), .Z(n26576) );
  NAND U35283 ( .A(n26577), .B(n26578), .Z(n26546) );
  NAND U35284 ( .A(n26579), .B(n26580), .Z(n26578) );
  OR U35285 ( .A(n26581), .B(n26582), .Z(n26579) );
  NANDN U35286 ( .A(n26583), .B(n26581), .Z(n26577) );
  IV U35287 ( .A(n26582), .Z(n26583) );
  NAND U35288 ( .A(n26584), .B(n26585), .Z(n26543) );
  NAND U35289 ( .A(n26586), .B(n26587), .Z(n26585) );
  NANDN U35290 ( .A(n26588), .B(n26589), .Z(n26586) );
  NANDN U35291 ( .A(n26589), .B(n26588), .Z(n26584) );
  AND U35292 ( .A(n26590), .B(n26591), .Z(n26545) );
  NAND U35293 ( .A(n26592), .B(n26593), .Z(n26591) );
  OR U35294 ( .A(n26594), .B(n26595), .Z(n26592) );
  NANDN U35295 ( .A(n26596), .B(n26594), .Z(n26590) );
  XNOR U35296 ( .A(n26571), .B(n26597), .Z(N63037) );
  XOR U35297 ( .A(n26573), .B(n26574), .Z(n26597) );
  XNOR U35298 ( .A(n26587), .B(n26598), .Z(n26574) );
  XOR U35299 ( .A(n26588), .B(n26589), .Z(n26598) );
  XOR U35300 ( .A(n26594), .B(n26599), .Z(n26589) );
  XOR U35301 ( .A(n26593), .B(n26596), .Z(n26599) );
  IV U35302 ( .A(n26595), .Z(n26596) );
  NAND U35303 ( .A(n26600), .B(n26601), .Z(n26595) );
  OR U35304 ( .A(n26602), .B(n26603), .Z(n26601) );
  OR U35305 ( .A(n26604), .B(n26605), .Z(n26600) );
  NAND U35306 ( .A(n26606), .B(n26607), .Z(n26593) );
  OR U35307 ( .A(n26608), .B(n26609), .Z(n26607) );
  OR U35308 ( .A(n26610), .B(n26611), .Z(n26606) );
  NOR U35309 ( .A(n26612), .B(n26613), .Z(n26594) );
  ANDN U35310 ( .B(n26614), .A(n26615), .Z(n26588) );
  XNOR U35311 ( .A(n26581), .B(n26616), .Z(n26587) );
  XNOR U35312 ( .A(n26580), .B(n26582), .Z(n26616) );
  NAND U35313 ( .A(n26617), .B(n26618), .Z(n26582) );
  OR U35314 ( .A(n26619), .B(n26620), .Z(n26618) );
  OR U35315 ( .A(n26621), .B(n26622), .Z(n26617) );
  NAND U35316 ( .A(n26623), .B(n26624), .Z(n26580) );
  OR U35317 ( .A(n26625), .B(n26626), .Z(n26624) );
  OR U35318 ( .A(n26627), .B(n26628), .Z(n26623) );
  ANDN U35319 ( .B(n26629), .A(n26630), .Z(n26581) );
  IV U35320 ( .A(n26631), .Z(n26629) );
  ANDN U35321 ( .B(n26632), .A(n26633), .Z(n26573) );
  XOR U35322 ( .A(n26559), .B(n26634), .Z(n26571) );
  XOR U35323 ( .A(n26560), .B(n26561), .Z(n26634) );
  XOR U35324 ( .A(n26566), .B(n26635), .Z(n26561) );
  XOR U35325 ( .A(n26565), .B(n26568), .Z(n26635) );
  IV U35326 ( .A(n26567), .Z(n26568) );
  NAND U35327 ( .A(n26636), .B(n26637), .Z(n26567) );
  OR U35328 ( .A(n26638), .B(n26639), .Z(n26637) );
  OR U35329 ( .A(n26640), .B(n26641), .Z(n26636) );
  NAND U35330 ( .A(n26642), .B(n26643), .Z(n26565) );
  OR U35331 ( .A(n26644), .B(n26645), .Z(n26643) );
  OR U35332 ( .A(n26646), .B(n26647), .Z(n26642) );
  NOR U35333 ( .A(n26648), .B(n26649), .Z(n26566) );
  ANDN U35334 ( .B(n26650), .A(n26651), .Z(n26560) );
  IV U35335 ( .A(n26652), .Z(n26650) );
  XNOR U35336 ( .A(n26553), .B(n26653), .Z(n26559) );
  XNOR U35337 ( .A(n26552), .B(n26554), .Z(n26653) );
  NAND U35338 ( .A(n26654), .B(n26655), .Z(n26554) );
  OR U35339 ( .A(n26656), .B(n26657), .Z(n26655) );
  OR U35340 ( .A(n26658), .B(n26659), .Z(n26654) );
  NAND U35341 ( .A(n26660), .B(n26661), .Z(n26552) );
  OR U35342 ( .A(n26662), .B(n26663), .Z(n26661) );
  OR U35343 ( .A(n26664), .B(n26665), .Z(n26660) );
  ANDN U35344 ( .B(n26666), .A(n26667), .Z(n26553) );
  IV U35345 ( .A(n26668), .Z(n26666) );
  XNOR U35346 ( .A(n26633), .B(n26632), .Z(N63036) );
  XOR U35347 ( .A(n26652), .B(n26651), .Z(n26632) );
  XNOR U35348 ( .A(n26667), .B(n26668), .Z(n26651) );
  XNOR U35349 ( .A(n26662), .B(n26663), .Z(n26668) );
  XNOR U35350 ( .A(n26664), .B(n26665), .Z(n26663) );
  XNOR U35351 ( .A(y[4525]), .B(x[4525]), .Z(n26665) );
  XNOR U35352 ( .A(y[4526]), .B(x[4526]), .Z(n26664) );
  XNOR U35353 ( .A(y[4524]), .B(x[4524]), .Z(n26662) );
  XNOR U35354 ( .A(n26656), .B(n26657), .Z(n26667) );
  XNOR U35355 ( .A(y[4521]), .B(x[4521]), .Z(n26657) );
  XNOR U35356 ( .A(n26658), .B(n26659), .Z(n26656) );
  XNOR U35357 ( .A(y[4522]), .B(x[4522]), .Z(n26659) );
  XNOR U35358 ( .A(y[4523]), .B(x[4523]), .Z(n26658) );
  XNOR U35359 ( .A(n26649), .B(n26648), .Z(n26652) );
  XNOR U35360 ( .A(n26644), .B(n26645), .Z(n26648) );
  XNOR U35361 ( .A(y[4518]), .B(x[4518]), .Z(n26645) );
  XNOR U35362 ( .A(n26646), .B(n26647), .Z(n26644) );
  XNOR U35363 ( .A(y[4519]), .B(x[4519]), .Z(n26647) );
  XNOR U35364 ( .A(y[4520]), .B(x[4520]), .Z(n26646) );
  XNOR U35365 ( .A(n26638), .B(n26639), .Z(n26649) );
  XNOR U35366 ( .A(y[4515]), .B(x[4515]), .Z(n26639) );
  XNOR U35367 ( .A(n26640), .B(n26641), .Z(n26638) );
  XNOR U35368 ( .A(y[4516]), .B(x[4516]), .Z(n26641) );
  XNOR U35369 ( .A(y[4517]), .B(x[4517]), .Z(n26640) );
  XOR U35370 ( .A(n26614), .B(n26615), .Z(n26633) );
  XNOR U35371 ( .A(n26630), .B(n26631), .Z(n26615) );
  XNOR U35372 ( .A(n26625), .B(n26626), .Z(n26631) );
  XNOR U35373 ( .A(n26627), .B(n26628), .Z(n26626) );
  XNOR U35374 ( .A(y[4513]), .B(x[4513]), .Z(n26628) );
  XNOR U35375 ( .A(y[4514]), .B(x[4514]), .Z(n26627) );
  XNOR U35376 ( .A(y[4512]), .B(x[4512]), .Z(n26625) );
  XNOR U35377 ( .A(n26619), .B(n26620), .Z(n26630) );
  XNOR U35378 ( .A(y[4509]), .B(x[4509]), .Z(n26620) );
  XNOR U35379 ( .A(n26621), .B(n26622), .Z(n26619) );
  XNOR U35380 ( .A(y[4510]), .B(x[4510]), .Z(n26622) );
  XNOR U35381 ( .A(y[4511]), .B(x[4511]), .Z(n26621) );
  XOR U35382 ( .A(n26613), .B(n26612), .Z(n26614) );
  XNOR U35383 ( .A(n26608), .B(n26609), .Z(n26612) );
  XNOR U35384 ( .A(y[4506]), .B(x[4506]), .Z(n26609) );
  XNOR U35385 ( .A(n26610), .B(n26611), .Z(n26608) );
  XNOR U35386 ( .A(y[4507]), .B(x[4507]), .Z(n26611) );
  XNOR U35387 ( .A(y[4508]), .B(x[4508]), .Z(n26610) );
  XNOR U35388 ( .A(n26602), .B(n26603), .Z(n26613) );
  XNOR U35389 ( .A(y[4503]), .B(x[4503]), .Z(n26603) );
  XNOR U35390 ( .A(n26604), .B(n26605), .Z(n26602) );
  XNOR U35391 ( .A(y[4504]), .B(x[4504]), .Z(n26605) );
  XNOR U35392 ( .A(y[4505]), .B(x[4505]), .Z(n26604) );
  NAND U35393 ( .A(n26669), .B(n26670), .Z(N63027) );
  NANDN U35394 ( .A(n26671), .B(n26672), .Z(n26670) );
  OR U35395 ( .A(n26673), .B(n26674), .Z(n26672) );
  NAND U35396 ( .A(n26673), .B(n26674), .Z(n26669) );
  XOR U35397 ( .A(n26673), .B(n26675), .Z(N63026) );
  XNOR U35398 ( .A(n26671), .B(n26674), .Z(n26675) );
  AND U35399 ( .A(n26676), .B(n26677), .Z(n26674) );
  NANDN U35400 ( .A(n26678), .B(n26679), .Z(n26677) );
  NANDN U35401 ( .A(n26680), .B(n26681), .Z(n26679) );
  NANDN U35402 ( .A(n26681), .B(n26680), .Z(n26676) );
  NAND U35403 ( .A(n26682), .B(n26683), .Z(n26671) );
  NANDN U35404 ( .A(n26684), .B(n26685), .Z(n26683) );
  OR U35405 ( .A(n26686), .B(n26687), .Z(n26685) );
  NAND U35406 ( .A(n26687), .B(n26686), .Z(n26682) );
  AND U35407 ( .A(n26688), .B(n26689), .Z(n26673) );
  NANDN U35408 ( .A(n26690), .B(n26691), .Z(n26689) );
  NANDN U35409 ( .A(n26692), .B(n26693), .Z(n26691) );
  NANDN U35410 ( .A(n26693), .B(n26692), .Z(n26688) );
  XOR U35411 ( .A(n26687), .B(n26694), .Z(N63025) );
  XOR U35412 ( .A(n26684), .B(n26686), .Z(n26694) );
  XNOR U35413 ( .A(n26680), .B(n26695), .Z(n26686) );
  XNOR U35414 ( .A(n26678), .B(n26681), .Z(n26695) );
  NAND U35415 ( .A(n26696), .B(n26697), .Z(n26681) );
  NAND U35416 ( .A(n26698), .B(n26699), .Z(n26697) );
  OR U35417 ( .A(n26700), .B(n26701), .Z(n26698) );
  NANDN U35418 ( .A(n26702), .B(n26700), .Z(n26696) );
  IV U35419 ( .A(n26701), .Z(n26702) );
  NAND U35420 ( .A(n26703), .B(n26704), .Z(n26678) );
  NAND U35421 ( .A(n26705), .B(n26706), .Z(n26704) );
  NANDN U35422 ( .A(n26707), .B(n26708), .Z(n26705) );
  NANDN U35423 ( .A(n26708), .B(n26707), .Z(n26703) );
  AND U35424 ( .A(n26709), .B(n26710), .Z(n26680) );
  NAND U35425 ( .A(n26711), .B(n26712), .Z(n26710) );
  OR U35426 ( .A(n26713), .B(n26714), .Z(n26711) );
  NANDN U35427 ( .A(n26715), .B(n26713), .Z(n26709) );
  NAND U35428 ( .A(n26716), .B(n26717), .Z(n26684) );
  NANDN U35429 ( .A(n26718), .B(n26719), .Z(n26717) );
  OR U35430 ( .A(n26720), .B(n26721), .Z(n26719) );
  NANDN U35431 ( .A(n26722), .B(n26720), .Z(n26716) );
  IV U35432 ( .A(n26721), .Z(n26722) );
  XNOR U35433 ( .A(n26692), .B(n26723), .Z(n26687) );
  XNOR U35434 ( .A(n26690), .B(n26693), .Z(n26723) );
  NAND U35435 ( .A(n26724), .B(n26725), .Z(n26693) );
  NAND U35436 ( .A(n26726), .B(n26727), .Z(n26725) );
  OR U35437 ( .A(n26728), .B(n26729), .Z(n26726) );
  NANDN U35438 ( .A(n26730), .B(n26728), .Z(n26724) );
  IV U35439 ( .A(n26729), .Z(n26730) );
  NAND U35440 ( .A(n26731), .B(n26732), .Z(n26690) );
  NAND U35441 ( .A(n26733), .B(n26734), .Z(n26732) );
  NANDN U35442 ( .A(n26735), .B(n26736), .Z(n26733) );
  NANDN U35443 ( .A(n26736), .B(n26735), .Z(n26731) );
  AND U35444 ( .A(n26737), .B(n26738), .Z(n26692) );
  NAND U35445 ( .A(n26739), .B(n26740), .Z(n26738) );
  OR U35446 ( .A(n26741), .B(n26742), .Z(n26739) );
  NANDN U35447 ( .A(n26743), .B(n26741), .Z(n26737) );
  XNOR U35448 ( .A(n26718), .B(n26744), .Z(N63024) );
  XOR U35449 ( .A(n26720), .B(n26721), .Z(n26744) );
  XNOR U35450 ( .A(n26734), .B(n26745), .Z(n26721) );
  XOR U35451 ( .A(n26735), .B(n26736), .Z(n26745) );
  XOR U35452 ( .A(n26741), .B(n26746), .Z(n26736) );
  XOR U35453 ( .A(n26740), .B(n26743), .Z(n26746) );
  IV U35454 ( .A(n26742), .Z(n26743) );
  NAND U35455 ( .A(n26747), .B(n26748), .Z(n26742) );
  OR U35456 ( .A(n26749), .B(n26750), .Z(n26748) );
  OR U35457 ( .A(n26751), .B(n26752), .Z(n26747) );
  NAND U35458 ( .A(n26753), .B(n26754), .Z(n26740) );
  OR U35459 ( .A(n26755), .B(n26756), .Z(n26754) );
  OR U35460 ( .A(n26757), .B(n26758), .Z(n26753) );
  NOR U35461 ( .A(n26759), .B(n26760), .Z(n26741) );
  ANDN U35462 ( .B(n26761), .A(n26762), .Z(n26735) );
  XNOR U35463 ( .A(n26728), .B(n26763), .Z(n26734) );
  XNOR U35464 ( .A(n26727), .B(n26729), .Z(n26763) );
  NAND U35465 ( .A(n26764), .B(n26765), .Z(n26729) );
  OR U35466 ( .A(n26766), .B(n26767), .Z(n26765) );
  OR U35467 ( .A(n26768), .B(n26769), .Z(n26764) );
  NAND U35468 ( .A(n26770), .B(n26771), .Z(n26727) );
  OR U35469 ( .A(n26772), .B(n26773), .Z(n26771) );
  OR U35470 ( .A(n26774), .B(n26775), .Z(n26770) );
  ANDN U35471 ( .B(n26776), .A(n26777), .Z(n26728) );
  IV U35472 ( .A(n26778), .Z(n26776) );
  ANDN U35473 ( .B(n26779), .A(n26780), .Z(n26720) );
  XOR U35474 ( .A(n26706), .B(n26781), .Z(n26718) );
  XOR U35475 ( .A(n26707), .B(n26708), .Z(n26781) );
  XOR U35476 ( .A(n26713), .B(n26782), .Z(n26708) );
  XOR U35477 ( .A(n26712), .B(n26715), .Z(n26782) );
  IV U35478 ( .A(n26714), .Z(n26715) );
  NAND U35479 ( .A(n26783), .B(n26784), .Z(n26714) );
  OR U35480 ( .A(n26785), .B(n26786), .Z(n26784) );
  OR U35481 ( .A(n26787), .B(n26788), .Z(n26783) );
  NAND U35482 ( .A(n26789), .B(n26790), .Z(n26712) );
  OR U35483 ( .A(n26791), .B(n26792), .Z(n26790) );
  OR U35484 ( .A(n26793), .B(n26794), .Z(n26789) );
  NOR U35485 ( .A(n26795), .B(n26796), .Z(n26713) );
  ANDN U35486 ( .B(n26797), .A(n26798), .Z(n26707) );
  IV U35487 ( .A(n26799), .Z(n26797) );
  XNOR U35488 ( .A(n26700), .B(n26800), .Z(n26706) );
  XNOR U35489 ( .A(n26699), .B(n26701), .Z(n26800) );
  NAND U35490 ( .A(n26801), .B(n26802), .Z(n26701) );
  OR U35491 ( .A(n26803), .B(n26804), .Z(n26802) );
  OR U35492 ( .A(n26805), .B(n26806), .Z(n26801) );
  NAND U35493 ( .A(n26807), .B(n26808), .Z(n26699) );
  OR U35494 ( .A(n26809), .B(n26810), .Z(n26808) );
  OR U35495 ( .A(n26811), .B(n26812), .Z(n26807) );
  ANDN U35496 ( .B(n26813), .A(n26814), .Z(n26700) );
  IV U35497 ( .A(n26815), .Z(n26813) );
  XNOR U35498 ( .A(n26780), .B(n26779), .Z(N63023) );
  XOR U35499 ( .A(n26799), .B(n26798), .Z(n26779) );
  XNOR U35500 ( .A(n26814), .B(n26815), .Z(n26798) );
  XNOR U35501 ( .A(n26809), .B(n26810), .Z(n26815) );
  XNOR U35502 ( .A(n26811), .B(n26812), .Z(n26810) );
  XNOR U35503 ( .A(y[4501]), .B(x[4501]), .Z(n26812) );
  XNOR U35504 ( .A(y[4502]), .B(x[4502]), .Z(n26811) );
  XNOR U35505 ( .A(y[4500]), .B(x[4500]), .Z(n26809) );
  XNOR U35506 ( .A(n26803), .B(n26804), .Z(n26814) );
  XNOR U35507 ( .A(y[4497]), .B(x[4497]), .Z(n26804) );
  XNOR U35508 ( .A(n26805), .B(n26806), .Z(n26803) );
  XNOR U35509 ( .A(y[4498]), .B(x[4498]), .Z(n26806) );
  XNOR U35510 ( .A(y[4499]), .B(x[4499]), .Z(n26805) );
  XNOR U35511 ( .A(n26796), .B(n26795), .Z(n26799) );
  XNOR U35512 ( .A(n26791), .B(n26792), .Z(n26795) );
  XNOR U35513 ( .A(y[4494]), .B(x[4494]), .Z(n26792) );
  XNOR U35514 ( .A(n26793), .B(n26794), .Z(n26791) );
  XNOR U35515 ( .A(y[4495]), .B(x[4495]), .Z(n26794) );
  XNOR U35516 ( .A(y[4496]), .B(x[4496]), .Z(n26793) );
  XNOR U35517 ( .A(n26785), .B(n26786), .Z(n26796) );
  XNOR U35518 ( .A(y[4491]), .B(x[4491]), .Z(n26786) );
  XNOR U35519 ( .A(n26787), .B(n26788), .Z(n26785) );
  XNOR U35520 ( .A(y[4492]), .B(x[4492]), .Z(n26788) );
  XNOR U35521 ( .A(y[4493]), .B(x[4493]), .Z(n26787) );
  XOR U35522 ( .A(n26761), .B(n26762), .Z(n26780) );
  XNOR U35523 ( .A(n26777), .B(n26778), .Z(n26762) );
  XNOR U35524 ( .A(n26772), .B(n26773), .Z(n26778) );
  XNOR U35525 ( .A(n26774), .B(n26775), .Z(n26773) );
  XNOR U35526 ( .A(y[4489]), .B(x[4489]), .Z(n26775) );
  XNOR U35527 ( .A(y[4490]), .B(x[4490]), .Z(n26774) );
  XNOR U35528 ( .A(y[4488]), .B(x[4488]), .Z(n26772) );
  XNOR U35529 ( .A(n26766), .B(n26767), .Z(n26777) );
  XNOR U35530 ( .A(y[4485]), .B(x[4485]), .Z(n26767) );
  XNOR U35531 ( .A(n26768), .B(n26769), .Z(n26766) );
  XNOR U35532 ( .A(y[4486]), .B(x[4486]), .Z(n26769) );
  XNOR U35533 ( .A(y[4487]), .B(x[4487]), .Z(n26768) );
  XOR U35534 ( .A(n26760), .B(n26759), .Z(n26761) );
  XNOR U35535 ( .A(n26755), .B(n26756), .Z(n26759) );
  XNOR U35536 ( .A(y[4482]), .B(x[4482]), .Z(n26756) );
  XNOR U35537 ( .A(n26757), .B(n26758), .Z(n26755) );
  XNOR U35538 ( .A(y[4483]), .B(x[4483]), .Z(n26758) );
  XNOR U35539 ( .A(y[4484]), .B(x[4484]), .Z(n26757) );
  XNOR U35540 ( .A(n26749), .B(n26750), .Z(n26760) );
  XNOR U35541 ( .A(y[4479]), .B(x[4479]), .Z(n26750) );
  XNOR U35542 ( .A(n26751), .B(n26752), .Z(n26749) );
  XNOR U35543 ( .A(y[4480]), .B(x[4480]), .Z(n26752) );
  XNOR U35544 ( .A(y[4481]), .B(x[4481]), .Z(n26751) );
  NAND U35545 ( .A(n26816), .B(n26817), .Z(N63014) );
  NANDN U35546 ( .A(n26818), .B(n26819), .Z(n26817) );
  OR U35547 ( .A(n26820), .B(n26821), .Z(n26819) );
  NAND U35548 ( .A(n26820), .B(n26821), .Z(n26816) );
  XOR U35549 ( .A(n26820), .B(n26822), .Z(N63013) );
  XNOR U35550 ( .A(n26818), .B(n26821), .Z(n26822) );
  AND U35551 ( .A(n26823), .B(n26824), .Z(n26821) );
  NANDN U35552 ( .A(n26825), .B(n26826), .Z(n26824) );
  NANDN U35553 ( .A(n26827), .B(n26828), .Z(n26826) );
  NANDN U35554 ( .A(n26828), .B(n26827), .Z(n26823) );
  NAND U35555 ( .A(n26829), .B(n26830), .Z(n26818) );
  NANDN U35556 ( .A(n26831), .B(n26832), .Z(n26830) );
  OR U35557 ( .A(n26833), .B(n26834), .Z(n26832) );
  NAND U35558 ( .A(n26834), .B(n26833), .Z(n26829) );
  AND U35559 ( .A(n26835), .B(n26836), .Z(n26820) );
  NANDN U35560 ( .A(n26837), .B(n26838), .Z(n26836) );
  NANDN U35561 ( .A(n26839), .B(n26840), .Z(n26838) );
  NANDN U35562 ( .A(n26840), .B(n26839), .Z(n26835) );
  XOR U35563 ( .A(n26834), .B(n26841), .Z(N63012) );
  XOR U35564 ( .A(n26831), .B(n26833), .Z(n26841) );
  XNOR U35565 ( .A(n26827), .B(n26842), .Z(n26833) );
  XNOR U35566 ( .A(n26825), .B(n26828), .Z(n26842) );
  NAND U35567 ( .A(n26843), .B(n26844), .Z(n26828) );
  NAND U35568 ( .A(n26845), .B(n26846), .Z(n26844) );
  OR U35569 ( .A(n26847), .B(n26848), .Z(n26845) );
  NANDN U35570 ( .A(n26849), .B(n26847), .Z(n26843) );
  IV U35571 ( .A(n26848), .Z(n26849) );
  NAND U35572 ( .A(n26850), .B(n26851), .Z(n26825) );
  NAND U35573 ( .A(n26852), .B(n26853), .Z(n26851) );
  NANDN U35574 ( .A(n26854), .B(n26855), .Z(n26852) );
  NANDN U35575 ( .A(n26855), .B(n26854), .Z(n26850) );
  AND U35576 ( .A(n26856), .B(n26857), .Z(n26827) );
  NAND U35577 ( .A(n26858), .B(n26859), .Z(n26857) );
  OR U35578 ( .A(n26860), .B(n26861), .Z(n26858) );
  NANDN U35579 ( .A(n26862), .B(n26860), .Z(n26856) );
  NAND U35580 ( .A(n26863), .B(n26864), .Z(n26831) );
  NANDN U35581 ( .A(n26865), .B(n26866), .Z(n26864) );
  OR U35582 ( .A(n26867), .B(n26868), .Z(n26866) );
  NANDN U35583 ( .A(n26869), .B(n26867), .Z(n26863) );
  IV U35584 ( .A(n26868), .Z(n26869) );
  XNOR U35585 ( .A(n26839), .B(n26870), .Z(n26834) );
  XNOR U35586 ( .A(n26837), .B(n26840), .Z(n26870) );
  NAND U35587 ( .A(n26871), .B(n26872), .Z(n26840) );
  NAND U35588 ( .A(n26873), .B(n26874), .Z(n26872) );
  OR U35589 ( .A(n26875), .B(n26876), .Z(n26873) );
  NANDN U35590 ( .A(n26877), .B(n26875), .Z(n26871) );
  IV U35591 ( .A(n26876), .Z(n26877) );
  NAND U35592 ( .A(n26878), .B(n26879), .Z(n26837) );
  NAND U35593 ( .A(n26880), .B(n26881), .Z(n26879) );
  NANDN U35594 ( .A(n26882), .B(n26883), .Z(n26880) );
  NANDN U35595 ( .A(n26883), .B(n26882), .Z(n26878) );
  AND U35596 ( .A(n26884), .B(n26885), .Z(n26839) );
  NAND U35597 ( .A(n26886), .B(n26887), .Z(n26885) );
  OR U35598 ( .A(n26888), .B(n26889), .Z(n26886) );
  NANDN U35599 ( .A(n26890), .B(n26888), .Z(n26884) );
  XNOR U35600 ( .A(n26865), .B(n26891), .Z(N63011) );
  XOR U35601 ( .A(n26867), .B(n26868), .Z(n26891) );
  XNOR U35602 ( .A(n26881), .B(n26892), .Z(n26868) );
  XOR U35603 ( .A(n26882), .B(n26883), .Z(n26892) );
  XOR U35604 ( .A(n26888), .B(n26893), .Z(n26883) );
  XOR U35605 ( .A(n26887), .B(n26890), .Z(n26893) );
  IV U35606 ( .A(n26889), .Z(n26890) );
  NAND U35607 ( .A(n26894), .B(n26895), .Z(n26889) );
  OR U35608 ( .A(n26896), .B(n26897), .Z(n26895) );
  OR U35609 ( .A(n26898), .B(n26899), .Z(n26894) );
  NAND U35610 ( .A(n26900), .B(n26901), .Z(n26887) );
  OR U35611 ( .A(n26902), .B(n26903), .Z(n26901) );
  OR U35612 ( .A(n26904), .B(n26905), .Z(n26900) );
  NOR U35613 ( .A(n26906), .B(n26907), .Z(n26888) );
  ANDN U35614 ( .B(n26908), .A(n26909), .Z(n26882) );
  XNOR U35615 ( .A(n26875), .B(n26910), .Z(n26881) );
  XNOR U35616 ( .A(n26874), .B(n26876), .Z(n26910) );
  NAND U35617 ( .A(n26911), .B(n26912), .Z(n26876) );
  OR U35618 ( .A(n26913), .B(n26914), .Z(n26912) );
  OR U35619 ( .A(n26915), .B(n26916), .Z(n26911) );
  NAND U35620 ( .A(n26917), .B(n26918), .Z(n26874) );
  OR U35621 ( .A(n26919), .B(n26920), .Z(n26918) );
  OR U35622 ( .A(n26921), .B(n26922), .Z(n26917) );
  ANDN U35623 ( .B(n26923), .A(n26924), .Z(n26875) );
  IV U35624 ( .A(n26925), .Z(n26923) );
  ANDN U35625 ( .B(n26926), .A(n26927), .Z(n26867) );
  XOR U35626 ( .A(n26853), .B(n26928), .Z(n26865) );
  XOR U35627 ( .A(n26854), .B(n26855), .Z(n26928) );
  XOR U35628 ( .A(n26860), .B(n26929), .Z(n26855) );
  XOR U35629 ( .A(n26859), .B(n26862), .Z(n26929) );
  IV U35630 ( .A(n26861), .Z(n26862) );
  NAND U35631 ( .A(n26930), .B(n26931), .Z(n26861) );
  OR U35632 ( .A(n26932), .B(n26933), .Z(n26931) );
  OR U35633 ( .A(n26934), .B(n26935), .Z(n26930) );
  NAND U35634 ( .A(n26936), .B(n26937), .Z(n26859) );
  OR U35635 ( .A(n26938), .B(n26939), .Z(n26937) );
  OR U35636 ( .A(n26940), .B(n26941), .Z(n26936) );
  NOR U35637 ( .A(n26942), .B(n26943), .Z(n26860) );
  ANDN U35638 ( .B(n26944), .A(n26945), .Z(n26854) );
  IV U35639 ( .A(n26946), .Z(n26944) );
  XNOR U35640 ( .A(n26847), .B(n26947), .Z(n26853) );
  XNOR U35641 ( .A(n26846), .B(n26848), .Z(n26947) );
  NAND U35642 ( .A(n26948), .B(n26949), .Z(n26848) );
  OR U35643 ( .A(n26950), .B(n26951), .Z(n26949) );
  OR U35644 ( .A(n26952), .B(n26953), .Z(n26948) );
  NAND U35645 ( .A(n26954), .B(n26955), .Z(n26846) );
  OR U35646 ( .A(n26956), .B(n26957), .Z(n26955) );
  OR U35647 ( .A(n26958), .B(n26959), .Z(n26954) );
  ANDN U35648 ( .B(n26960), .A(n26961), .Z(n26847) );
  IV U35649 ( .A(n26962), .Z(n26960) );
  XNOR U35650 ( .A(n26927), .B(n26926), .Z(N63010) );
  XOR U35651 ( .A(n26946), .B(n26945), .Z(n26926) );
  XNOR U35652 ( .A(n26961), .B(n26962), .Z(n26945) );
  XNOR U35653 ( .A(n26956), .B(n26957), .Z(n26962) );
  XNOR U35654 ( .A(n26958), .B(n26959), .Z(n26957) );
  XNOR U35655 ( .A(y[4477]), .B(x[4477]), .Z(n26959) );
  XNOR U35656 ( .A(y[4478]), .B(x[4478]), .Z(n26958) );
  XNOR U35657 ( .A(y[4476]), .B(x[4476]), .Z(n26956) );
  XNOR U35658 ( .A(n26950), .B(n26951), .Z(n26961) );
  XNOR U35659 ( .A(y[4473]), .B(x[4473]), .Z(n26951) );
  XNOR U35660 ( .A(n26952), .B(n26953), .Z(n26950) );
  XNOR U35661 ( .A(y[4474]), .B(x[4474]), .Z(n26953) );
  XNOR U35662 ( .A(y[4475]), .B(x[4475]), .Z(n26952) );
  XNOR U35663 ( .A(n26943), .B(n26942), .Z(n26946) );
  XNOR U35664 ( .A(n26938), .B(n26939), .Z(n26942) );
  XNOR U35665 ( .A(y[4470]), .B(x[4470]), .Z(n26939) );
  XNOR U35666 ( .A(n26940), .B(n26941), .Z(n26938) );
  XNOR U35667 ( .A(y[4471]), .B(x[4471]), .Z(n26941) );
  XNOR U35668 ( .A(y[4472]), .B(x[4472]), .Z(n26940) );
  XNOR U35669 ( .A(n26932), .B(n26933), .Z(n26943) );
  XNOR U35670 ( .A(y[4467]), .B(x[4467]), .Z(n26933) );
  XNOR U35671 ( .A(n26934), .B(n26935), .Z(n26932) );
  XNOR U35672 ( .A(y[4468]), .B(x[4468]), .Z(n26935) );
  XNOR U35673 ( .A(y[4469]), .B(x[4469]), .Z(n26934) );
  XOR U35674 ( .A(n26908), .B(n26909), .Z(n26927) );
  XNOR U35675 ( .A(n26924), .B(n26925), .Z(n26909) );
  XNOR U35676 ( .A(n26919), .B(n26920), .Z(n26925) );
  XNOR U35677 ( .A(n26921), .B(n26922), .Z(n26920) );
  XNOR U35678 ( .A(y[4465]), .B(x[4465]), .Z(n26922) );
  XNOR U35679 ( .A(y[4466]), .B(x[4466]), .Z(n26921) );
  XNOR U35680 ( .A(y[4464]), .B(x[4464]), .Z(n26919) );
  XNOR U35681 ( .A(n26913), .B(n26914), .Z(n26924) );
  XNOR U35682 ( .A(y[4461]), .B(x[4461]), .Z(n26914) );
  XNOR U35683 ( .A(n26915), .B(n26916), .Z(n26913) );
  XNOR U35684 ( .A(y[4462]), .B(x[4462]), .Z(n26916) );
  XNOR U35685 ( .A(y[4463]), .B(x[4463]), .Z(n26915) );
  XOR U35686 ( .A(n26907), .B(n26906), .Z(n26908) );
  XNOR U35687 ( .A(n26902), .B(n26903), .Z(n26906) );
  XNOR U35688 ( .A(y[4458]), .B(x[4458]), .Z(n26903) );
  XNOR U35689 ( .A(n26904), .B(n26905), .Z(n26902) );
  XNOR U35690 ( .A(y[4459]), .B(x[4459]), .Z(n26905) );
  XNOR U35691 ( .A(y[4460]), .B(x[4460]), .Z(n26904) );
  XNOR U35692 ( .A(n26896), .B(n26897), .Z(n26907) );
  XNOR U35693 ( .A(y[4455]), .B(x[4455]), .Z(n26897) );
  XNOR U35694 ( .A(n26898), .B(n26899), .Z(n26896) );
  XNOR U35695 ( .A(y[4456]), .B(x[4456]), .Z(n26899) );
  XNOR U35696 ( .A(y[4457]), .B(x[4457]), .Z(n26898) );
  NAND U35697 ( .A(n26963), .B(n26964), .Z(N63001) );
  NANDN U35698 ( .A(n26965), .B(n26966), .Z(n26964) );
  OR U35699 ( .A(n26967), .B(n26968), .Z(n26966) );
  NAND U35700 ( .A(n26967), .B(n26968), .Z(n26963) );
  XOR U35701 ( .A(n26967), .B(n26969), .Z(N63000) );
  XNOR U35702 ( .A(n26965), .B(n26968), .Z(n26969) );
  AND U35703 ( .A(n26970), .B(n26971), .Z(n26968) );
  NANDN U35704 ( .A(n26972), .B(n26973), .Z(n26971) );
  NANDN U35705 ( .A(n26974), .B(n26975), .Z(n26973) );
  NANDN U35706 ( .A(n26975), .B(n26974), .Z(n26970) );
  NAND U35707 ( .A(n26976), .B(n26977), .Z(n26965) );
  NANDN U35708 ( .A(n26978), .B(n26979), .Z(n26977) );
  OR U35709 ( .A(n26980), .B(n26981), .Z(n26979) );
  NAND U35710 ( .A(n26981), .B(n26980), .Z(n26976) );
  AND U35711 ( .A(n26982), .B(n26983), .Z(n26967) );
  NANDN U35712 ( .A(n26984), .B(n26985), .Z(n26983) );
  NANDN U35713 ( .A(n26986), .B(n26987), .Z(n26985) );
  NANDN U35714 ( .A(n26987), .B(n26986), .Z(n26982) );
  XOR U35715 ( .A(n26981), .B(n26988), .Z(N62999) );
  XOR U35716 ( .A(n26978), .B(n26980), .Z(n26988) );
  XNOR U35717 ( .A(n26974), .B(n26989), .Z(n26980) );
  XNOR U35718 ( .A(n26972), .B(n26975), .Z(n26989) );
  NAND U35719 ( .A(n26990), .B(n26991), .Z(n26975) );
  NAND U35720 ( .A(n26992), .B(n26993), .Z(n26991) );
  OR U35721 ( .A(n26994), .B(n26995), .Z(n26992) );
  NANDN U35722 ( .A(n26996), .B(n26994), .Z(n26990) );
  IV U35723 ( .A(n26995), .Z(n26996) );
  NAND U35724 ( .A(n26997), .B(n26998), .Z(n26972) );
  NAND U35725 ( .A(n26999), .B(n27000), .Z(n26998) );
  NANDN U35726 ( .A(n27001), .B(n27002), .Z(n26999) );
  NANDN U35727 ( .A(n27002), .B(n27001), .Z(n26997) );
  AND U35728 ( .A(n27003), .B(n27004), .Z(n26974) );
  NAND U35729 ( .A(n27005), .B(n27006), .Z(n27004) );
  OR U35730 ( .A(n27007), .B(n27008), .Z(n27005) );
  NANDN U35731 ( .A(n27009), .B(n27007), .Z(n27003) );
  NAND U35732 ( .A(n27010), .B(n27011), .Z(n26978) );
  NANDN U35733 ( .A(n27012), .B(n27013), .Z(n27011) );
  OR U35734 ( .A(n27014), .B(n27015), .Z(n27013) );
  NANDN U35735 ( .A(n27016), .B(n27014), .Z(n27010) );
  IV U35736 ( .A(n27015), .Z(n27016) );
  XNOR U35737 ( .A(n26986), .B(n27017), .Z(n26981) );
  XNOR U35738 ( .A(n26984), .B(n26987), .Z(n27017) );
  NAND U35739 ( .A(n27018), .B(n27019), .Z(n26987) );
  NAND U35740 ( .A(n27020), .B(n27021), .Z(n27019) );
  OR U35741 ( .A(n27022), .B(n27023), .Z(n27020) );
  NANDN U35742 ( .A(n27024), .B(n27022), .Z(n27018) );
  IV U35743 ( .A(n27023), .Z(n27024) );
  NAND U35744 ( .A(n27025), .B(n27026), .Z(n26984) );
  NAND U35745 ( .A(n27027), .B(n27028), .Z(n27026) );
  NANDN U35746 ( .A(n27029), .B(n27030), .Z(n27027) );
  NANDN U35747 ( .A(n27030), .B(n27029), .Z(n27025) );
  AND U35748 ( .A(n27031), .B(n27032), .Z(n26986) );
  NAND U35749 ( .A(n27033), .B(n27034), .Z(n27032) );
  OR U35750 ( .A(n27035), .B(n27036), .Z(n27033) );
  NANDN U35751 ( .A(n27037), .B(n27035), .Z(n27031) );
  XNOR U35752 ( .A(n27012), .B(n27038), .Z(N62998) );
  XOR U35753 ( .A(n27014), .B(n27015), .Z(n27038) );
  XNOR U35754 ( .A(n27028), .B(n27039), .Z(n27015) );
  XOR U35755 ( .A(n27029), .B(n27030), .Z(n27039) );
  XOR U35756 ( .A(n27035), .B(n27040), .Z(n27030) );
  XOR U35757 ( .A(n27034), .B(n27037), .Z(n27040) );
  IV U35758 ( .A(n27036), .Z(n27037) );
  NAND U35759 ( .A(n27041), .B(n27042), .Z(n27036) );
  OR U35760 ( .A(n27043), .B(n27044), .Z(n27042) );
  OR U35761 ( .A(n27045), .B(n27046), .Z(n27041) );
  NAND U35762 ( .A(n27047), .B(n27048), .Z(n27034) );
  OR U35763 ( .A(n27049), .B(n27050), .Z(n27048) );
  OR U35764 ( .A(n27051), .B(n27052), .Z(n27047) );
  NOR U35765 ( .A(n27053), .B(n27054), .Z(n27035) );
  ANDN U35766 ( .B(n27055), .A(n27056), .Z(n27029) );
  XNOR U35767 ( .A(n27022), .B(n27057), .Z(n27028) );
  XNOR U35768 ( .A(n27021), .B(n27023), .Z(n27057) );
  NAND U35769 ( .A(n27058), .B(n27059), .Z(n27023) );
  OR U35770 ( .A(n27060), .B(n27061), .Z(n27059) );
  OR U35771 ( .A(n27062), .B(n27063), .Z(n27058) );
  NAND U35772 ( .A(n27064), .B(n27065), .Z(n27021) );
  OR U35773 ( .A(n27066), .B(n27067), .Z(n27065) );
  OR U35774 ( .A(n27068), .B(n27069), .Z(n27064) );
  ANDN U35775 ( .B(n27070), .A(n27071), .Z(n27022) );
  IV U35776 ( .A(n27072), .Z(n27070) );
  ANDN U35777 ( .B(n27073), .A(n27074), .Z(n27014) );
  XOR U35778 ( .A(n27000), .B(n27075), .Z(n27012) );
  XOR U35779 ( .A(n27001), .B(n27002), .Z(n27075) );
  XOR U35780 ( .A(n27007), .B(n27076), .Z(n27002) );
  XOR U35781 ( .A(n27006), .B(n27009), .Z(n27076) );
  IV U35782 ( .A(n27008), .Z(n27009) );
  NAND U35783 ( .A(n27077), .B(n27078), .Z(n27008) );
  OR U35784 ( .A(n27079), .B(n27080), .Z(n27078) );
  OR U35785 ( .A(n27081), .B(n27082), .Z(n27077) );
  NAND U35786 ( .A(n27083), .B(n27084), .Z(n27006) );
  OR U35787 ( .A(n27085), .B(n27086), .Z(n27084) );
  OR U35788 ( .A(n27087), .B(n27088), .Z(n27083) );
  NOR U35789 ( .A(n27089), .B(n27090), .Z(n27007) );
  ANDN U35790 ( .B(n27091), .A(n27092), .Z(n27001) );
  IV U35791 ( .A(n27093), .Z(n27091) );
  XNOR U35792 ( .A(n26994), .B(n27094), .Z(n27000) );
  XNOR U35793 ( .A(n26993), .B(n26995), .Z(n27094) );
  NAND U35794 ( .A(n27095), .B(n27096), .Z(n26995) );
  OR U35795 ( .A(n27097), .B(n27098), .Z(n27096) );
  OR U35796 ( .A(n27099), .B(n27100), .Z(n27095) );
  NAND U35797 ( .A(n27101), .B(n27102), .Z(n26993) );
  OR U35798 ( .A(n27103), .B(n27104), .Z(n27102) );
  OR U35799 ( .A(n27105), .B(n27106), .Z(n27101) );
  ANDN U35800 ( .B(n27107), .A(n27108), .Z(n26994) );
  IV U35801 ( .A(n27109), .Z(n27107) );
  XNOR U35802 ( .A(n27074), .B(n27073), .Z(N62997) );
  XOR U35803 ( .A(n27093), .B(n27092), .Z(n27073) );
  XNOR U35804 ( .A(n27108), .B(n27109), .Z(n27092) );
  XNOR U35805 ( .A(n27103), .B(n27104), .Z(n27109) );
  XNOR U35806 ( .A(n27105), .B(n27106), .Z(n27104) );
  XNOR U35807 ( .A(y[4453]), .B(x[4453]), .Z(n27106) );
  XNOR U35808 ( .A(y[4454]), .B(x[4454]), .Z(n27105) );
  XNOR U35809 ( .A(y[4452]), .B(x[4452]), .Z(n27103) );
  XNOR U35810 ( .A(n27097), .B(n27098), .Z(n27108) );
  XNOR U35811 ( .A(y[4449]), .B(x[4449]), .Z(n27098) );
  XNOR U35812 ( .A(n27099), .B(n27100), .Z(n27097) );
  XNOR U35813 ( .A(y[4450]), .B(x[4450]), .Z(n27100) );
  XNOR U35814 ( .A(y[4451]), .B(x[4451]), .Z(n27099) );
  XNOR U35815 ( .A(n27090), .B(n27089), .Z(n27093) );
  XNOR U35816 ( .A(n27085), .B(n27086), .Z(n27089) );
  XNOR U35817 ( .A(y[4446]), .B(x[4446]), .Z(n27086) );
  XNOR U35818 ( .A(n27087), .B(n27088), .Z(n27085) );
  XNOR U35819 ( .A(y[4447]), .B(x[4447]), .Z(n27088) );
  XNOR U35820 ( .A(y[4448]), .B(x[4448]), .Z(n27087) );
  XNOR U35821 ( .A(n27079), .B(n27080), .Z(n27090) );
  XNOR U35822 ( .A(y[4443]), .B(x[4443]), .Z(n27080) );
  XNOR U35823 ( .A(n27081), .B(n27082), .Z(n27079) );
  XNOR U35824 ( .A(y[4444]), .B(x[4444]), .Z(n27082) );
  XNOR U35825 ( .A(y[4445]), .B(x[4445]), .Z(n27081) );
  XOR U35826 ( .A(n27055), .B(n27056), .Z(n27074) );
  XNOR U35827 ( .A(n27071), .B(n27072), .Z(n27056) );
  XNOR U35828 ( .A(n27066), .B(n27067), .Z(n27072) );
  XNOR U35829 ( .A(n27068), .B(n27069), .Z(n27067) );
  XNOR U35830 ( .A(y[4441]), .B(x[4441]), .Z(n27069) );
  XNOR U35831 ( .A(y[4442]), .B(x[4442]), .Z(n27068) );
  XNOR U35832 ( .A(y[4440]), .B(x[4440]), .Z(n27066) );
  XNOR U35833 ( .A(n27060), .B(n27061), .Z(n27071) );
  XNOR U35834 ( .A(y[4437]), .B(x[4437]), .Z(n27061) );
  XNOR U35835 ( .A(n27062), .B(n27063), .Z(n27060) );
  XNOR U35836 ( .A(y[4438]), .B(x[4438]), .Z(n27063) );
  XNOR U35837 ( .A(y[4439]), .B(x[4439]), .Z(n27062) );
  XOR U35838 ( .A(n27054), .B(n27053), .Z(n27055) );
  XNOR U35839 ( .A(n27049), .B(n27050), .Z(n27053) );
  XNOR U35840 ( .A(y[4434]), .B(x[4434]), .Z(n27050) );
  XNOR U35841 ( .A(n27051), .B(n27052), .Z(n27049) );
  XNOR U35842 ( .A(y[4435]), .B(x[4435]), .Z(n27052) );
  XNOR U35843 ( .A(y[4436]), .B(x[4436]), .Z(n27051) );
  XNOR U35844 ( .A(n27043), .B(n27044), .Z(n27054) );
  XNOR U35845 ( .A(y[4431]), .B(x[4431]), .Z(n27044) );
  XNOR U35846 ( .A(n27045), .B(n27046), .Z(n27043) );
  XNOR U35847 ( .A(y[4432]), .B(x[4432]), .Z(n27046) );
  XNOR U35848 ( .A(y[4433]), .B(x[4433]), .Z(n27045) );
  NAND U35849 ( .A(n27110), .B(n27111), .Z(N62988) );
  NANDN U35850 ( .A(n27112), .B(n27113), .Z(n27111) );
  OR U35851 ( .A(n27114), .B(n27115), .Z(n27113) );
  NAND U35852 ( .A(n27114), .B(n27115), .Z(n27110) );
  XOR U35853 ( .A(n27114), .B(n27116), .Z(N62987) );
  XNOR U35854 ( .A(n27112), .B(n27115), .Z(n27116) );
  AND U35855 ( .A(n27117), .B(n27118), .Z(n27115) );
  NANDN U35856 ( .A(n27119), .B(n27120), .Z(n27118) );
  NANDN U35857 ( .A(n27121), .B(n27122), .Z(n27120) );
  NANDN U35858 ( .A(n27122), .B(n27121), .Z(n27117) );
  NAND U35859 ( .A(n27123), .B(n27124), .Z(n27112) );
  NANDN U35860 ( .A(n27125), .B(n27126), .Z(n27124) );
  OR U35861 ( .A(n27127), .B(n27128), .Z(n27126) );
  NAND U35862 ( .A(n27128), .B(n27127), .Z(n27123) );
  AND U35863 ( .A(n27129), .B(n27130), .Z(n27114) );
  NANDN U35864 ( .A(n27131), .B(n27132), .Z(n27130) );
  NANDN U35865 ( .A(n27133), .B(n27134), .Z(n27132) );
  NANDN U35866 ( .A(n27134), .B(n27133), .Z(n27129) );
  XOR U35867 ( .A(n27128), .B(n27135), .Z(N62986) );
  XOR U35868 ( .A(n27125), .B(n27127), .Z(n27135) );
  XNOR U35869 ( .A(n27121), .B(n27136), .Z(n27127) );
  XNOR U35870 ( .A(n27119), .B(n27122), .Z(n27136) );
  NAND U35871 ( .A(n27137), .B(n27138), .Z(n27122) );
  NAND U35872 ( .A(n27139), .B(n27140), .Z(n27138) );
  OR U35873 ( .A(n27141), .B(n27142), .Z(n27139) );
  NANDN U35874 ( .A(n27143), .B(n27141), .Z(n27137) );
  IV U35875 ( .A(n27142), .Z(n27143) );
  NAND U35876 ( .A(n27144), .B(n27145), .Z(n27119) );
  NAND U35877 ( .A(n27146), .B(n27147), .Z(n27145) );
  NANDN U35878 ( .A(n27148), .B(n27149), .Z(n27146) );
  NANDN U35879 ( .A(n27149), .B(n27148), .Z(n27144) );
  AND U35880 ( .A(n27150), .B(n27151), .Z(n27121) );
  NAND U35881 ( .A(n27152), .B(n27153), .Z(n27151) );
  OR U35882 ( .A(n27154), .B(n27155), .Z(n27152) );
  NANDN U35883 ( .A(n27156), .B(n27154), .Z(n27150) );
  NAND U35884 ( .A(n27157), .B(n27158), .Z(n27125) );
  NANDN U35885 ( .A(n27159), .B(n27160), .Z(n27158) );
  OR U35886 ( .A(n27161), .B(n27162), .Z(n27160) );
  NANDN U35887 ( .A(n27163), .B(n27161), .Z(n27157) );
  IV U35888 ( .A(n27162), .Z(n27163) );
  XNOR U35889 ( .A(n27133), .B(n27164), .Z(n27128) );
  XNOR U35890 ( .A(n27131), .B(n27134), .Z(n27164) );
  NAND U35891 ( .A(n27165), .B(n27166), .Z(n27134) );
  NAND U35892 ( .A(n27167), .B(n27168), .Z(n27166) );
  OR U35893 ( .A(n27169), .B(n27170), .Z(n27167) );
  NANDN U35894 ( .A(n27171), .B(n27169), .Z(n27165) );
  IV U35895 ( .A(n27170), .Z(n27171) );
  NAND U35896 ( .A(n27172), .B(n27173), .Z(n27131) );
  NAND U35897 ( .A(n27174), .B(n27175), .Z(n27173) );
  NANDN U35898 ( .A(n27176), .B(n27177), .Z(n27174) );
  NANDN U35899 ( .A(n27177), .B(n27176), .Z(n27172) );
  AND U35900 ( .A(n27178), .B(n27179), .Z(n27133) );
  NAND U35901 ( .A(n27180), .B(n27181), .Z(n27179) );
  OR U35902 ( .A(n27182), .B(n27183), .Z(n27180) );
  NANDN U35903 ( .A(n27184), .B(n27182), .Z(n27178) );
  XNOR U35904 ( .A(n27159), .B(n27185), .Z(N62985) );
  XOR U35905 ( .A(n27161), .B(n27162), .Z(n27185) );
  XNOR U35906 ( .A(n27175), .B(n27186), .Z(n27162) );
  XOR U35907 ( .A(n27176), .B(n27177), .Z(n27186) );
  XOR U35908 ( .A(n27182), .B(n27187), .Z(n27177) );
  XOR U35909 ( .A(n27181), .B(n27184), .Z(n27187) );
  IV U35910 ( .A(n27183), .Z(n27184) );
  NAND U35911 ( .A(n27188), .B(n27189), .Z(n27183) );
  OR U35912 ( .A(n27190), .B(n27191), .Z(n27189) );
  OR U35913 ( .A(n27192), .B(n27193), .Z(n27188) );
  NAND U35914 ( .A(n27194), .B(n27195), .Z(n27181) );
  OR U35915 ( .A(n27196), .B(n27197), .Z(n27195) );
  OR U35916 ( .A(n27198), .B(n27199), .Z(n27194) );
  NOR U35917 ( .A(n27200), .B(n27201), .Z(n27182) );
  ANDN U35918 ( .B(n27202), .A(n27203), .Z(n27176) );
  XNOR U35919 ( .A(n27169), .B(n27204), .Z(n27175) );
  XNOR U35920 ( .A(n27168), .B(n27170), .Z(n27204) );
  NAND U35921 ( .A(n27205), .B(n27206), .Z(n27170) );
  OR U35922 ( .A(n27207), .B(n27208), .Z(n27206) );
  OR U35923 ( .A(n27209), .B(n27210), .Z(n27205) );
  NAND U35924 ( .A(n27211), .B(n27212), .Z(n27168) );
  OR U35925 ( .A(n27213), .B(n27214), .Z(n27212) );
  OR U35926 ( .A(n27215), .B(n27216), .Z(n27211) );
  ANDN U35927 ( .B(n27217), .A(n27218), .Z(n27169) );
  IV U35928 ( .A(n27219), .Z(n27217) );
  ANDN U35929 ( .B(n27220), .A(n27221), .Z(n27161) );
  XOR U35930 ( .A(n27147), .B(n27222), .Z(n27159) );
  XOR U35931 ( .A(n27148), .B(n27149), .Z(n27222) );
  XOR U35932 ( .A(n27154), .B(n27223), .Z(n27149) );
  XOR U35933 ( .A(n27153), .B(n27156), .Z(n27223) );
  IV U35934 ( .A(n27155), .Z(n27156) );
  NAND U35935 ( .A(n27224), .B(n27225), .Z(n27155) );
  OR U35936 ( .A(n27226), .B(n27227), .Z(n27225) );
  OR U35937 ( .A(n27228), .B(n27229), .Z(n27224) );
  NAND U35938 ( .A(n27230), .B(n27231), .Z(n27153) );
  OR U35939 ( .A(n27232), .B(n27233), .Z(n27231) );
  OR U35940 ( .A(n27234), .B(n27235), .Z(n27230) );
  NOR U35941 ( .A(n27236), .B(n27237), .Z(n27154) );
  ANDN U35942 ( .B(n27238), .A(n27239), .Z(n27148) );
  IV U35943 ( .A(n27240), .Z(n27238) );
  XNOR U35944 ( .A(n27141), .B(n27241), .Z(n27147) );
  XNOR U35945 ( .A(n27140), .B(n27142), .Z(n27241) );
  NAND U35946 ( .A(n27242), .B(n27243), .Z(n27142) );
  OR U35947 ( .A(n27244), .B(n27245), .Z(n27243) );
  OR U35948 ( .A(n27246), .B(n27247), .Z(n27242) );
  NAND U35949 ( .A(n27248), .B(n27249), .Z(n27140) );
  OR U35950 ( .A(n27250), .B(n27251), .Z(n27249) );
  OR U35951 ( .A(n27252), .B(n27253), .Z(n27248) );
  ANDN U35952 ( .B(n27254), .A(n27255), .Z(n27141) );
  IV U35953 ( .A(n27256), .Z(n27254) );
  XNOR U35954 ( .A(n27221), .B(n27220), .Z(N62984) );
  XOR U35955 ( .A(n27240), .B(n27239), .Z(n27220) );
  XNOR U35956 ( .A(n27255), .B(n27256), .Z(n27239) );
  XNOR U35957 ( .A(n27250), .B(n27251), .Z(n27256) );
  XNOR U35958 ( .A(n27252), .B(n27253), .Z(n27251) );
  XNOR U35959 ( .A(y[4429]), .B(x[4429]), .Z(n27253) );
  XNOR U35960 ( .A(y[4430]), .B(x[4430]), .Z(n27252) );
  XNOR U35961 ( .A(y[4428]), .B(x[4428]), .Z(n27250) );
  XNOR U35962 ( .A(n27244), .B(n27245), .Z(n27255) );
  XNOR U35963 ( .A(y[4425]), .B(x[4425]), .Z(n27245) );
  XNOR U35964 ( .A(n27246), .B(n27247), .Z(n27244) );
  XNOR U35965 ( .A(y[4426]), .B(x[4426]), .Z(n27247) );
  XNOR U35966 ( .A(y[4427]), .B(x[4427]), .Z(n27246) );
  XNOR U35967 ( .A(n27237), .B(n27236), .Z(n27240) );
  XNOR U35968 ( .A(n27232), .B(n27233), .Z(n27236) );
  XNOR U35969 ( .A(y[4422]), .B(x[4422]), .Z(n27233) );
  XNOR U35970 ( .A(n27234), .B(n27235), .Z(n27232) );
  XNOR U35971 ( .A(y[4423]), .B(x[4423]), .Z(n27235) );
  XNOR U35972 ( .A(y[4424]), .B(x[4424]), .Z(n27234) );
  XNOR U35973 ( .A(n27226), .B(n27227), .Z(n27237) );
  XNOR U35974 ( .A(y[4419]), .B(x[4419]), .Z(n27227) );
  XNOR U35975 ( .A(n27228), .B(n27229), .Z(n27226) );
  XNOR U35976 ( .A(y[4420]), .B(x[4420]), .Z(n27229) );
  XNOR U35977 ( .A(y[4421]), .B(x[4421]), .Z(n27228) );
  XOR U35978 ( .A(n27202), .B(n27203), .Z(n27221) );
  XNOR U35979 ( .A(n27218), .B(n27219), .Z(n27203) );
  XNOR U35980 ( .A(n27213), .B(n27214), .Z(n27219) );
  XNOR U35981 ( .A(n27215), .B(n27216), .Z(n27214) );
  XNOR U35982 ( .A(y[4417]), .B(x[4417]), .Z(n27216) );
  XNOR U35983 ( .A(y[4418]), .B(x[4418]), .Z(n27215) );
  XNOR U35984 ( .A(y[4416]), .B(x[4416]), .Z(n27213) );
  XNOR U35985 ( .A(n27207), .B(n27208), .Z(n27218) );
  XNOR U35986 ( .A(y[4413]), .B(x[4413]), .Z(n27208) );
  XNOR U35987 ( .A(n27209), .B(n27210), .Z(n27207) );
  XNOR U35988 ( .A(y[4414]), .B(x[4414]), .Z(n27210) );
  XNOR U35989 ( .A(y[4415]), .B(x[4415]), .Z(n27209) );
  XOR U35990 ( .A(n27201), .B(n27200), .Z(n27202) );
  XNOR U35991 ( .A(n27196), .B(n27197), .Z(n27200) );
  XNOR U35992 ( .A(y[4410]), .B(x[4410]), .Z(n27197) );
  XNOR U35993 ( .A(n27198), .B(n27199), .Z(n27196) );
  XNOR U35994 ( .A(y[4411]), .B(x[4411]), .Z(n27199) );
  XNOR U35995 ( .A(y[4412]), .B(x[4412]), .Z(n27198) );
  XNOR U35996 ( .A(n27190), .B(n27191), .Z(n27201) );
  XNOR U35997 ( .A(y[4407]), .B(x[4407]), .Z(n27191) );
  XNOR U35998 ( .A(n27192), .B(n27193), .Z(n27190) );
  XNOR U35999 ( .A(y[4408]), .B(x[4408]), .Z(n27193) );
  XNOR U36000 ( .A(y[4409]), .B(x[4409]), .Z(n27192) );
  NAND U36001 ( .A(n27257), .B(n27258), .Z(N62975) );
  NANDN U36002 ( .A(n27259), .B(n27260), .Z(n27258) );
  OR U36003 ( .A(n27261), .B(n27262), .Z(n27260) );
  NAND U36004 ( .A(n27261), .B(n27262), .Z(n27257) );
  XOR U36005 ( .A(n27261), .B(n27263), .Z(N62974) );
  XNOR U36006 ( .A(n27259), .B(n27262), .Z(n27263) );
  AND U36007 ( .A(n27264), .B(n27265), .Z(n27262) );
  NANDN U36008 ( .A(n27266), .B(n27267), .Z(n27265) );
  NANDN U36009 ( .A(n27268), .B(n27269), .Z(n27267) );
  NANDN U36010 ( .A(n27269), .B(n27268), .Z(n27264) );
  NAND U36011 ( .A(n27270), .B(n27271), .Z(n27259) );
  NANDN U36012 ( .A(n27272), .B(n27273), .Z(n27271) );
  OR U36013 ( .A(n27274), .B(n27275), .Z(n27273) );
  NAND U36014 ( .A(n27275), .B(n27274), .Z(n27270) );
  AND U36015 ( .A(n27276), .B(n27277), .Z(n27261) );
  NANDN U36016 ( .A(n27278), .B(n27279), .Z(n27277) );
  NANDN U36017 ( .A(n27280), .B(n27281), .Z(n27279) );
  NANDN U36018 ( .A(n27281), .B(n27280), .Z(n27276) );
  XOR U36019 ( .A(n27275), .B(n27282), .Z(N62973) );
  XOR U36020 ( .A(n27272), .B(n27274), .Z(n27282) );
  XNOR U36021 ( .A(n27268), .B(n27283), .Z(n27274) );
  XNOR U36022 ( .A(n27266), .B(n27269), .Z(n27283) );
  NAND U36023 ( .A(n27284), .B(n27285), .Z(n27269) );
  NAND U36024 ( .A(n27286), .B(n27287), .Z(n27285) );
  OR U36025 ( .A(n27288), .B(n27289), .Z(n27286) );
  NANDN U36026 ( .A(n27290), .B(n27288), .Z(n27284) );
  IV U36027 ( .A(n27289), .Z(n27290) );
  NAND U36028 ( .A(n27291), .B(n27292), .Z(n27266) );
  NAND U36029 ( .A(n27293), .B(n27294), .Z(n27292) );
  NANDN U36030 ( .A(n27295), .B(n27296), .Z(n27293) );
  NANDN U36031 ( .A(n27296), .B(n27295), .Z(n27291) );
  AND U36032 ( .A(n27297), .B(n27298), .Z(n27268) );
  NAND U36033 ( .A(n27299), .B(n27300), .Z(n27298) );
  OR U36034 ( .A(n27301), .B(n27302), .Z(n27299) );
  NANDN U36035 ( .A(n27303), .B(n27301), .Z(n27297) );
  NAND U36036 ( .A(n27304), .B(n27305), .Z(n27272) );
  NANDN U36037 ( .A(n27306), .B(n27307), .Z(n27305) );
  OR U36038 ( .A(n27308), .B(n27309), .Z(n27307) );
  NANDN U36039 ( .A(n27310), .B(n27308), .Z(n27304) );
  IV U36040 ( .A(n27309), .Z(n27310) );
  XNOR U36041 ( .A(n27280), .B(n27311), .Z(n27275) );
  XNOR U36042 ( .A(n27278), .B(n27281), .Z(n27311) );
  NAND U36043 ( .A(n27312), .B(n27313), .Z(n27281) );
  NAND U36044 ( .A(n27314), .B(n27315), .Z(n27313) );
  OR U36045 ( .A(n27316), .B(n27317), .Z(n27314) );
  NANDN U36046 ( .A(n27318), .B(n27316), .Z(n27312) );
  IV U36047 ( .A(n27317), .Z(n27318) );
  NAND U36048 ( .A(n27319), .B(n27320), .Z(n27278) );
  NAND U36049 ( .A(n27321), .B(n27322), .Z(n27320) );
  NANDN U36050 ( .A(n27323), .B(n27324), .Z(n27321) );
  NANDN U36051 ( .A(n27324), .B(n27323), .Z(n27319) );
  AND U36052 ( .A(n27325), .B(n27326), .Z(n27280) );
  NAND U36053 ( .A(n27327), .B(n27328), .Z(n27326) );
  OR U36054 ( .A(n27329), .B(n27330), .Z(n27327) );
  NANDN U36055 ( .A(n27331), .B(n27329), .Z(n27325) );
  XNOR U36056 ( .A(n27306), .B(n27332), .Z(N62972) );
  XOR U36057 ( .A(n27308), .B(n27309), .Z(n27332) );
  XNOR U36058 ( .A(n27322), .B(n27333), .Z(n27309) );
  XOR U36059 ( .A(n27323), .B(n27324), .Z(n27333) );
  XOR U36060 ( .A(n27329), .B(n27334), .Z(n27324) );
  XOR U36061 ( .A(n27328), .B(n27331), .Z(n27334) );
  IV U36062 ( .A(n27330), .Z(n27331) );
  NAND U36063 ( .A(n27335), .B(n27336), .Z(n27330) );
  OR U36064 ( .A(n27337), .B(n27338), .Z(n27336) );
  OR U36065 ( .A(n27339), .B(n27340), .Z(n27335) );
  NAND U36066 ( .A(n27341), .B(n27342), .Z(n27328) );
  OR U36067 ( .A(n27343), .B(n27344), .Z(n27342) );
  OR U36068 ( .A(n27345), .B(n27346), .Z(n27341) );
  NOR U36069 ( .A(n27347), .B(n27348), .Z(n27329) );
  ANDN U36070 ( .B(n27349), .A(n27350), .Z(n27323) );
  XNOR U36071 ( .A(n27316), .B(n27351), .Z(n27322) );
  XNOR U36072 ( .A(n27315), .B(n27317), .Z(n27351) );
  NAND U36073 ( .A(n27352), .B(n27353), .Z(n27317) );
  OR U36074 ( .A(n27354), .B(n27355), .Z(n27353) );
  OR U36075 ( .A(n27356), .B(n27357), .Z(n27352) );
  NAND U36076 ( .A(n27358), .B(n27359), .Z(n27315) );
  OR U36077 ( .A(n27360), .B(n27361), .Z(n27359) );
  OR U36078 ( .A(n27362), .B(n27363), .Z(n27358) );
  ANDN U36079 ( .B(n27364), .A(n27365), .Z(n27316) );
  IV U36080 ( .A(n27366), .Z(n27364) );
  ANDN U36081 ( .B(n27367), .A(n27368), .Z(n27308) );
  XOR U36082 ( .A(n27294), .B(n27369), .Z(n27306) );
  XOR U36083 ( .A(n27295), .B(n27296), .Z(n27369) );
  XOR U36084 ( .A(n27301), .B(n27370), .Z(n27296) );
  XOR U36085 ( .A(n27300), .B(n27303), .Z(n27370) );
  IV U36086 ( .A(n27302), .Z(n27303) );
  NAND U36087 ( .A(n27371), .B(n27372), .Z(n27302) );
  OR U36088 ( .A(n27373), .B(n27374), .Z(n27372) );
  OR U36089 ( .A(n27375), .B(n27376), .Z(n27371) );
  NAND U36090 ( .A(n27377), .B(n27378), .Z(n27300) );
  OR U36091 ( .A(n27379), .B(n27380), .Z(n27378) );
  OR U36092 ( .A(n27381), .B(n27382), .Z(n27377) );
  NOR U36093 ( .A(n27383), .B(n27384), .Z(n27301) );
  ANDN U36094 ( .B(n27385), .A(n27386), .Z(n27295) );
  IV U36095 ( .A(n27387), .Z(n27385) );
  XNOR U36096 ( .A(n27288), .B(n27388), .Z(n27294) );
  XNOR U36097 ( .A(n27287), .B(n27289), .Z(n27388) );
  NAND U36098 ( .A(n27389), .B(n27390), .Z(n27289) );
  OR U36099 ( .A(n27391), .B(n27392), .Z(n27390) );
  OR U36100 ( .A(n27393), .B(n27394), .Z(n27389) );
  NAND U36101 ( .A(n27395), .B(n27396), .Z(n27287) );
  OR U36102 ( .A(n27397), .B(n27398), .Z(n27396) );
  OR U36103 ( .A(n27399), .B(n27400), .Z(n27395) );
  ANDN U36104 ( .B(n27401), .A(n27402), .Z(n27288) );
  IV U36105 ( .A(n27403), .Z(n27401) );
  XNOR U36106 ( .A(n27368), .B(n27367), .Z(N62971) );
  XOR U36107 ( .A(n27387), .B(n27386), .Z(n27367) );
  XNOR U36108 ( .A(n27402), .B(n27403), .Z(n27386) );
  XNOR U36109 ( .A(n27397), .B(n27398), .Z(n27403) );
  XNOR U36110 ( .A(n27399), .B(n27400), .Z(n27398) );
  XNOR U36111 ( .A(y[4405]), .B(x[4405]), .Z(n27400) );
  XNOR U36112 ( .A(y[4406]), .B(x[4406]), .Z(n27399) );
  XNOR U36113 ( .A(y[4404]), .B(x[4404]), .Z(n27397) );
  XNOR U36114 ( .A(n27391), .B(n27392), .Z(n27402) );
  XNOR U36115 ( .A(y[4401]), .B(x[4401]), .Z(n27392) );
  XNOR U36116 ( .A(n27393), .B(n27394), .Z(n27391) );
  XNOR U36117 ( .A(y[4402]), .B(x[4402]), .Z(n27394) );
  XNOR U36118 ( .A(y[4403]), .B(x[4403]), .Z(n27393) );
  XNOR U36119 ( .A(n27384), .B(n27383), .Z(n27387) );
  XNOR U36120 ( .A(n27379), .B(n27380), .Z(n27383) );
  XNOR U36121 ( .A(y[4398]), .B(x[4398]), .Z(n27380) );
  XNOR U36122 ( .A(n27381), .B(n27382), .Z(n27379) );
  XNOR U36123 ( .A(y[4399]), .B(x[4399]), .Z(n27382) );
  XNOR U36124 ( .A(y[4400]), .B(x[4400]), .Z(n27381) );
  XNOR U36125 ( .A(n27373), .B(n27374), .Z(n27384) );
  XNOR U36126 ( .A(y[4395]), .B(x[4395]), .Z(n27374) );
  XNOR U36127 ( .A(n27375), .B(n27376), .Z(n27373) );
  XNOR U36128 ( .A(y[4396]), .B(x[4396]), .Z(n27376) );
  XNOR U36129 ( .A(y[4397]), .B(x[4397]), .Z(n27375) );
  XOR U36130 ( .A(n27349), .B(n27350), .Z(n27368) );
  XNOR U36131 ( .A(n27365), .B(n27366), .Z(n27350) );
  XNOR U36132 ( .A(n27360), .B(n27361), .Z(n27366) );
  XNOR U36133 ( .A(n27362), .B(n27363), .Z(n27361) );
  XNOR U36134 ( .A(y[4393]), .B(x[4393]), .Z(n27363) );
  XNOR U36135 ( .A(y[4394]), .B(x[4394]), .Z(n27362) );
  XNOR U36136 ( .A(y[4392]), .B(x[4392]), .Z(n27360) );
  XNOR U36137 ( .A(n27354), .B(n27355), .Z(n27365) );
  XNOR U36138 ( .A(y[4389]), .B(x[4389]), .Z(n27355) );
  XNOR U36139 ( .A(n27356), .B(n27357), .Z(n27354) );
  XNOR U36140 ( .A(y[4390]), .B(x[4390]), .Z(n27357) );
  XNOR U36141 ( .A(y[4391]), .B(x[4391]), .Z(n27356) );
  XOR U36142 ( .A(n27348), .B(n27347), .Z(n27349) );
  XNOR U36143 ( .A(n27343), .B(n27344), .Z(n27347) );
  XNOR U36144 ( .A(y[4386]), .B(x[4386]), .Z(n27344) );
  XNOR U36145 ( .A(n27345), .B(n27346), .Z(n27343) );
  XNOR U36146 ( .A(y[4387]), .B(x[4387]), .Z(n27346) );
  XNOR U36147 ( .A(y[4388]), .B(x[4388]), .Z(n27345) );
  XNOR U36148 ( .A(n27337), .B(n27338), .Z(n27348) );
  XNOR U36149 ( .A(y[4383]), .B(x[4383]), .Z(n27338) );
  XNOR U36150 ( .A(n27339), .B(n27340), .Z(n27337) );
  XNOR U36151 ( .A(y[4384]), .B(x[4384]), .Z(n27340) );
  XNOR U36152 ( .A(y[4385]), .B(x[4385]), .Z(n27339) );
  NAND U36153 ( .A(n27404), .B(n27405), .Z(N62962) );
  NANDN U36154 ( .A(n27406), .B(n27407), .Z(n27405) );
  OR U36155 ( .A(n27408), .B(n27409), .Z(n27407) );
  NAND U36156 ( .A(n27408), .B(n27409), .Z(n27404) );
  XOR U36157 ( .A(n27408), .B(n27410), .Z(N62961) );
  XNOR U36158 ( .A(n27406), .B(n27409), .Z(n27410) );
  AND U36159 ( .A(n27411), .B(n27412), .Z(n27409) );
  NANDN U36160 ( .A(n27413), .B(n27414), .Z(n27412) );
  NANDN U36161 ( .A(n27415), .B(n27416), .Z(n27414) );
  NANDN U36162 ( .A(n27416), .B(n27415), .Z(n27411) );
  NAND U36163 ( .A(n27417), .B(n27418), .Z(n27406) );
  NANDN U36164 ( .A(n27419), .B(n27420), .Z(n27418) );
  OR U36165 ( .A(n27421), .B(n27422), .Z(n27420) );
  NAND U36166 ( .A(n27422), .B(n27421), .Z(n27417) );
  AND U36167 ( .A(n27423), .B(n27424), .Z(n27408) );
  NANDN U36168 ( .A(n27425), .B(n27426), .Z(n27424) );
  NANDN U36169 ( .A(n27427), .B(n27428), .Z(n27426) );
  NANDN U36170 ( .A(n27428), .B(n27427), .Z(n27423) );
  XOR U36171 ( .A(n27422), .B(n27429), .Z(N62960) );
  XOR U36172 ( .A(n27419), .B(n27421), .Z(n27429) );
  XNOR U36173 ( .A(n27415), .B(n27430), .Z(n27421) );
  XNOR U36174 ( .A(n27413), .B(n27416), .Z(n27430) );
  NAND U36175 ( .A(n27431), .B(n27432), .Z(n27416) );
  NAND U36176 ( .A(n27433), .B(n27434), .Z(n27432) );
  OR U36177 ( .A(n27435), .B(n27436), .Z(n27433) );
  NANDN U36178 ( .A(n27437), .B(n27435), .Z(n27431) );
  IV U36179 ( .A(n27436), .Z(n27437) );
  NAND U36180 ( .A(n27438), .B(n27439), .Z(n27413) );
  NAND U36181 ( .A(n27440), .B(n27441), .Z(n27439) );
  NANDN U36182 ( .A(n27442), .B(n27443), .Z(n27440) );
  NANDN U36183 ( .A(n27443), .B(n27442), .Z(n27438) );
  AND U36184 ( .A(n27444), .B(n27445), .Z(n27415) );
  NAND U36185 ( .A(n27446), .B(n27447), .Z(n27445) );
  OR U36186 ( .A(n27448), .B(n27449), .Z(n27446) );
  NANDN U36187 ( .A(n27450), .B(n27448), .Z(n27444) );
  NAND U36188 ( .A(n27451), .B(n27452), .Z(n27419) );
  NANDN U36189 ( .A(n27453), .B(n27454), .Z(n27452) );
  OR U36190 ( .A(n27455), .B(n27456), .Z(n27454) );
  NANDN U36191 ( .A(n27457), .B(n27455), .Z(n27451) );
  IV U36192 ( .A(n27456), .Z(n27457) );
  XNOR U36193 ( .A(n27427), .B(n27458), .Z(n27422) );
  XNOR U36194 ( .A(n27425), .B(n27428), .Z(n27458) );
  NAND U36195 ( .A(n27459), .B(n27460), .Z(n27428) );
  NAND U36196 ( .A(n27461), .B(n27462), .Z(n27460) );
  OR U36197 ( .A(n27463), .B(n27464), .Z(n27461) );
  NANDN U36198 ( .A(n27465), .B(n27463), .Z(n27459) );
  IV U36199 ( .A(n27464), .Z(n27465) );
  NAND U36200 ( .A(n27466), .B(n27467), .Z(n27425) );
  NAND U36201 ( .A(n27468), .B(n27469), .Z(n27467) );
  NANDN U36202 ( .A(n27470), .B(n27471), .Z(n27468) );
  NANDN U36203 ( .A(n27471), .B(n27470), .Z(n27466) );
  AND U36204 ( .A(n27472), .B(n27473), .Z(n27427) );
  NAND U36205 ( .A(n27474), .B(n27475), .Z(n27473) );
  OR U36206 ( .A(n27476), .B(n27477), .Z(n27474) );
  NANDN U36207 ( .A(n27478), .B(n27476), .Z(n27472) );
  XNOR U36208 ( .A(n27453), .B(n27479), .Z(N62959) );
  XOR U36209 ( .A(n27455), .B(n27456), .Z(n27479) );
  XNOR U36210 ( .A(n27469), .B(n27480), .Z(n27456) );
  XOR U36211 ( .A(n27470), .B(n27471), .Z(n27480) );
  XOR U36212 ( .A(n27476), .B(n27481), .Z(n27471) );
  XOR U36213 ( .A(n27475), .B(n27478), .Z(n27481) );
  IV U36214 ( .A(n27477), .Z(n27478) );
  NAND U36215 ( .A(n27482), .B(n27483), .Z(n27477) );
  OR U36216 ( .A(n27484), .B(n27485), .Z(n27483) );
  OR U36217 ( .A(n27486), .B(n27487), .Z(n27482) );
  NAND U36218 ( .A(n27488), .B(n27489), .Z(n27475) );
  OR U36219 ( .A(n27490), .B(n27491), .Z(n27489) );
  OR U36220 ( .A(n27492), .B(n27493), .Z(n27488) );
  NOR U36221 ( .A(n27494), .B(n27495), .Z(n27476) );
  ANDN U36222 ( .B(n27496), .A(n27497), .Z(n27470) );
  XNOR U36223 ( .A(n27463), .B(n27498), .Z(n27469) );
  XNOR U36224 ( .A(n27462), .B(n27464), .Z(n27498) );
  NAND U36225 ( .A(n27499), .B(n27500), .Z(n27464) );
  OR U36226 ( .A(n27501), .B(n27502), .Z(n27500) );
  OR U36227 ( .A(n27503), .B(n27504), .Z(n27499) );
  NAND U36228 ( .A(n27505), .B(n27506), .Z(n27462) );
  OR U36229 ( .A(n27507), .B(n27508), .Z(n27506) );
  OR U36230 ( .A(n27509), .B(n27510), .Z(n27505) );
  ANDN U36231 ( .B(n27511), .A(n27512), .Z(n27463) );
  IV U36232 ( .A(n27513), .Z(n27511) );
  ANDN U36233 ( .B(n27514), .A(n27515), .Z(n27455) );
  XOR U36234 ( .A(n27441), .B(n27516), .Z(n27453) );
  XOR U36235 ( .A(n27442), .B(n27443), .Z(n27516) );
  XOR U36236 ( .A(n27448), .B(n27517), .Z(n27443) );
  XOR U36237 ( .A(n27447), .B(n27450), .Z(n27517) );
  IV U36238 ( .A(n27449), .Z(n27450) );
  NAND U36239 ( .A(n27518), .B(n27519), .Z(n27449) );
  OR U36240 ( .A(n27520), .B(n27521), .Z(n27519) );
  OR U36241 ( .A(n27522), .B(n27523), .Z(n27518) );
  NAND U36242 ( .A(n27524), .B(n27525), .Z(n27447) );
  OR U36243 ( .A(n27526), .B(n27527), .Z(n27525) );
  OR U36244 ( .A(n27528), .B(n27529), .Z(n27524) );
  NOR U36245 ( .A(n27530), .B(n27531), .Z(n27448) );
  ANDN U36246 ( .B(n27532), .A(n27533), .Z(n27442) );
  IV U36247 ( .A(n27534), .Z(n27532) );
  XNOR U36248 ( .A(n27435), .B(n27535), .Z(n27441) );
  XNOR U36249 ( .A(n27434), .B(n27436), .Z(n27535) );
  NAND U36250 ( .A(n27536), .B(n27537), .Z(n27436) );
  OR U36251 ( .A(n27538), .B(n27539), .Z(n27537) );
  OR U36252 ( .A(n27540), .B(n27541), .Z(n27536) );
  NAND U36253 ( .A(n27542), .B(n27543), .Z(n27434) );
  OR U36254 ( .A(n27544), .B(n27545), .Z(n27543) );
  OR U36255 ( .A(n27546), .B(n27547), .Z(n27542) );
  ANDN U36256 ( .B(n27548), .A(n27549), .Z(n27435) );
  IV U36257 ( .A(n27550), .Z(n27548) );
  XNOR U36258 ( .A(n27515), .B(n27514), .Z(N62958) );
  XOR U36259 ( .A(n27534), .B(n27533), .Z(n27514) );
  XNOR U36260 ( .A(n27549), .B(n27550), .Z(n27533) );
  XNOR U36261 ( .A(n27544), .B(n27545), .Z(n27550) );
  XNOR U36262 ( .A(n27546), .B(n27547), .Z(n27545) );
  XNOR U36263 ( .A(y[4381]), .B(x[4381]), .Z(n27547) );
  XNOR U36264 ( .A(y[4382]), .B(x[4382]), .Z(n27546) );
  XNOR U36265 ( .A(y[4380]), .B(x[4380]), .Z(n27544) );
  XNOR U36266 ( .A(n27538), .B(n27539), .Z(n27549) );
  XNOR U36267 ( .A(y[4377]), .B(x[4377]), .Z(n27539) );
  XNOR U36268 ( .A(n27540), .B(n27541), .Z(n27538) );
  XNOR U36269 ( .A(y[4378]), .B(x[4378]), .Z(n27541) );
  XNOR U36270 ( .A(y[4379]), .B(x[4379]), .Z(n27540) );
  XNOR U36271 ( .A(n27531), .B(n27530), .Z(n27534) );
  XNOR U36272 ( .A(n27526), .B(n27527), .Z(n27530) );
  XNOR U36273 ( .A(y[4374]), .B(x[4374]), .Z(n27527) );
  XNOR U36274 ( .A(n27528), .B(n27529), .Z(n27526) );
  XNOR U36275 ( .A(y[4375]), .B(x[4375]), .Z(n27529) );
  XNOR U36276 ( .A(y[4376]), .B(x[4376]), .Z(n27528) );
  XNOR U36277 ( .A(n27520), .B(n27521), .Z(n27531) );
  XNOR U36278 ( .A(y[4371]), .B(x[4371]), .Z(n27521) );
  XNOR U36279 ( .A(n27522), .B(n27523), .Z(n27520) );
  XNOR U36280 ( .A(y[4372]), .B(x[4372]), .Z(n27523) );
  XNOR U36281 ( .A(y[4373]), .B(x[4373]), .Z(n27522) );
  XOR U36282 ( .A(n27496), .B(n27497), .Z(n27515) );
  XNOR U36283 ( .A(n27512), .B(n27513), .Z(n27497) );
  XNOR U36284 ( .A(n27507), .B(n27508), .Z(n27513) );
  XNOR U36285 ( .A(n27509), .B(n27510), .Z(n27508) );
  XNOR U36286 ( .A(y[4369]), .B(x[4369]), .Z(n27510) );
  XNOR U36287 ( .A(y[4370]), .B(x[4370]), .Z(n27509) );
  XNOR U36288 ( .A(y[4368]), .B(x[4368]), .Z(n27507) );
  XNOR U36289 ( .A(n27501), .B(n27502), .Z(n27512) );
  XNOR U36290 ( .A(y[4365]), .B(x[4365]), .Z(n27502) );
  XNOR U36291 ( .A(n27503), .B(n27504), .Z(n27501) );
  XNOR U36292 ( .A(y[4366]), .B(x[4366]), .Z(n27504) );
  XNOR U36293 ( .A(y[4367]), .B(x[4367]), .Z(n27503) );
  XOR U36294 ( .A(n27495), .B(n27494), .Z(n27496) );
  XNOR U36295 ( .A(n27490), .B(n27491), .Z(n27494) );
  XNOR U36296 ( .A(y[4362]), .B(x[4362]), .Z(n27491) );
  XNOR U36297 ( .A(n27492), .B(n27493), .Z(n27490) );
  XNOR U36298 ( .A(y[4363]), .B(x[4363]), .Z(n27493) );
  XNOR U36299 ( .A(y[4364]), .B(x[4364]), .Z(n27492) );
  XNOR U36300 ( .A(n27484), .B(n27485), .Z(n27495) );
  XNOR U36301 ( .A(y[4359]), .B(x[4359]), .Z(n27485) );
  XNOR U36302 ( .A(n27486), .B(n27487), .Z(n27484) );
  XNOR U36303 ( .A(y[4360]), .B(x[4360]), .Z(n27487) );
  XNOR U36304 ( .A(y[4361]), .B(x[4361]), .Z(n27486) );
  NAND U36305 ( .A(n27551), .B(n27552), .Z(N62949) );
  NANDN U36306 ( .A(n27553), .B(n27554), .Z(n27552) );
  OR U36307 ( .A(n27555), .B(n27556), .Z(n27554) );
  NAND U36308 ( .A(n27555), .B(n27556), .Z(n27551) );
  XOR U36309 ( .A(n27555), .B(n27557), .Z(N62948) );
  XNOR U36310 ( .A(n27553), .B(n27556), .Z(n27557) );
  AND U36311 ( .A(n27558), .B(n27559), .Z(n27556) );
  NANDN U36312 ( .A(n27560), .B(n27561), .Z(n27559) );
  NANDN U36313 ( .A(n27562), .B(n27563), .Z(n27561) );
  NANDN U36314 ( .A(n27563), .B(n27562), .Z(n27558) );
  NAND U36315 ( .A(n27564), .B(n27565), .Z(n27553) );
  NANDN U36316 ( .A(n27566), .B(n27567), .Z(n27565) );
  OR U36317 ( .A(n27568), .B(n27569), .Z(n27567) );
  NAND U36318 ( .A(n27569), .B(n27568), .Z(n27564) );
  AND U36319 ( .A(n27570), .B(n27571), .Z(n27555) );
  NANDN U36320 ( .A(n27572), .B(n27573), .Z(n27571) );
  NANDN U36321 ( .A(n27574), .B(n27575), .Z(n27573) );
  NANDN U36322 ( .A(n27575), .B(n27574), .Z(n27570) );
  XOR U36323 ( .A(n27569), .B(n27576), .Z(N62947) );
  XOR U36324 ( .A(n27566), .B(n27568), .Z(n27576) );
  XNOR U36325 ( .A(n27562), .B(n27577), .Z(n27568) );
  XNOR U36326 ( .A(n27560), .B(n27563), .Z(n27577) );
  NAND U36327 ( .A(n27578), .B(n27579), .Z(n27563) );
  NAND U36328 ( .A(n27580), .B(n27581), .Z(n27579) );
  OR U36329 ( .A(n27582), .B(n27583), .Z(n27580) );
  NANDN U36330 ( .A(n27584), .B(n27582), .Z(n27578) );
  IV U36331 ( .A(n27583), .Z(n27584) );
  NAND U36332 ( .A(n27585), .B(n27586), .Z(n27560) );
  NAND U36333 ( .A(n27587), .B(n27588), .Z(n27586) );
  NANDN U36334 ( .A(n27589), .B(n27590), .Z(n27587) );
  NANDN U36335 ( .A(n27590), .B(n27589), .Z(n27585) );
  AND U36336 ( .A(n27591), .B(n27592), .Z(n27562) );
  NAND U36337 ( .A(n27593), .B(n27594), .Z(n27592) );
  OR U36338 ( .A(n27595), .B(n27596), .Z(n27593) );
  NANDN U36339 ( .A(n27597), .B(n27595), .Z(n27591) );
  NAND U36340 ( .A(n27598), .B(n27599), .Z(n27566) );
  NANDN U36341 ( .A(n27600), .B(n27601), .Z(n27599) );
  OR U36342 ( .A(n27602), .B(n27603), .Z(n27601) );
  NANDN U36343 ( .A(n27604), .B(n27602), .Z(n27598) );
  IV U36344 ( .A(n27603), .Z(n27604) );
  XNOR U36345 ( .A(n27574), .B(n27605), .Z(n27569) );
  XNOR U36346 ( .A(n27572), .B(n27575), .Z(n27605) );
  NAND U36347 ( .A(n27606), .B(n27607), .Z(n27575) );
  NAND U36348 ( .A(n27608), .B(n27609), .Z(n27607) );
  OR U36349 ( .A(n27610), .B(n27611), .Z(n27608) );
  NANDN U36350 ( .A(n27612), .B(n27610), .Z(n27606) );
  IV U36351 ( .A(n27611), .Z(n27612) );
  NAND U36352 ( .A(n27613), .B(n27614), .Z(n27572) );
  NAND U36353 ( .A(n27615), .B(n27616), .Z(n27614) );
  NANDN U36354 ( .A(n27617), .B(n27618), .Z(n27615) );
  NANDN U36355 ( .A(n27618), .B(n27617), .Z(n27613) );
  AND U36356 ( .A(n27619), .B(n27620), .Z(n27574) );
  NAND U36357 ( .A(n27621), .B(n27622), .Z(n27620) );
  OR U36358 ( .A(n27623), .B(n27624), .Z(n27621) );
  NANDN U36359 ( .A(n27625), .B(n27623), .Z(n27619) );
  XNOR U36360 ( .A(n27600), .B(n27626), .Z(N62946) );
  XOR U36361 ( .A(n27602), .B(n27603), .Z(n27626) );
  XNOR U36362 ( .A(n27616), .B(n27627), .Z(n27603) );
  XOR U36363 ( .A(n27617), .B(n27618), .Z(n27627) );
  XOR U36364 ( .A(n27623), .B(n27628), .Z(n27618) );
  XOR U36365 ( .A(n27622), .B(n27625), .Z(n27628) );
  IV U36366 ( .A(n27624), .Z(n27625) );
  NAND U36367 ( .A(n27629), .B(n27630), .Z(n27624) );
  OR U36368 ( .A(n27631), .B(n27632), .Z(n27630) );
  OR U36369 ( .A(n27633), .B(n27634), .Z(n27629) );
  NAND U36370 ( .A(n27635), .B(n27636), .Z(n27622) );
  OR U36371 ( .A(n27637), .B(n27638), .Z(n27636) );
  OR U36372 ( .A(n27639), .B(n27640), .Z(n27635) );
  NOR U36373 ( .A(n27641), .B(n27642), .Z(n27623) );
  ANDN U36374 ( .B(n27643), .A(n27644), .Z(n27617) );
  XNOR U36375 ( .A(n27610), .B(n27645), .Z(n27616) );
  XNOR U36376 ( .A(n27609), .B(n27611), .Z(n27645) );
  NAND U36377 ( .A(n27646), .B(n27647), .Z(n27611) );
  OR U36378 ( .A(n27648), .B(n27649), .Z(n27647) );
  OR U36379 ( .A(n27650), .B(n27651), .Z(n27646) );
  NAND U36380 ( .A(n27652), .B(n27653), .Z(n27609) );
  OR U36381 ( .A(n27654), .B(n27655), .Z(n27653) );
  OR U36382 ( .A(n27656), .B(n27657), .Z(n27652) );
  ANDN U36383 ( .B(n27658), .A(n27659), .Z(n27610) );
  IV U36384 ( .A(n27660), .Z(n27658) );
  ANDN U36385 ( .B(n27661), .A(n27662), .Z(n27602) );
  XOR U36386 ( .A(n27588), .B(n27663), .Z(n27600) );
  XOR U36387 ( .A(n27589), .B(n27590), .Z(n27663) );
  XOR U36388 ( .A(n27595), .B(n27664), .Z(n27590) );
  XOR U36389 ( .A(n27594), .B(n27597), .Z(n27664) );
  IV U36390 ( .A(n27596), .Z(n27597) );
  NAND U36391 ( .A(n27665), .B(n27666), .Z(n27596) );
  OR U36392 ( .A(n27667), .B(n27668), .Z(n27666) );
  OR U36393 ( .A(n27669), .B(n27670), .Z(n27665) );
  NAND U36394 ( .A(n27671), .B(n27672), .Z(n27594) );
  OR U36395 ( .A(n27673), .B(n27674), .Z(n27672) );
  OR U36396 ( .A(n27675), .B(n27676), .Z(n27671) );
  NOR U36397 ( .A(n27677), .B(n27678), .Z(n27595) );
  ANDN U36398 ( .B(n27679), .A(n27680), .Z(n27589) );
  IV U36399 ( .A(n27681), .Z(n27679) );
  XNOR U36400 ( .A(n27582), .B(n27682), .Z(n27588) );
  XNOR U36401 ( .A(n27581), .B(n27583), .Z(n27682) );
  NAND U36402 ( .A(n27683), .B(n27684), .Z(n27583) );
  OR U36403 ( .A(n27685), .B(n27686), .Z(n27684) );
  OR U36404 ( .A(n27687), .B(n27688), .Z(n27683) );
  NAND U36405 ( .A(n27689), .B(n27690), .Z(n27581) );
  OR U36406 ( .A(n27691), .B(n27692), .Z(n27690) );
  OR U36407 ( .A(n27693), .B(n27694), .Z(n27689) );
  ANDN U36408 ( .B(n27695), .A(n27696), .Z(n27582) );
  IV U36409 ( .A(n27697), .Z(n27695) );
  XNOR U36410 ( .A(n27662), .B(n27661), .Z(N62945) );
  XOR U36411 ( .A(n27681), .B(n27680), .Z(n27661) );
  XNOR U36412 ( .A(n27696), .B(n27697), .Z(n27680) );
  XNOR U36413 ( .A(n27691), .B(n27692), .Z(n27697) );
  XNOR U36414 ( .A(n27693), .B(n27694), .Z(n27692) );
  XNOR U36415 ( .A(y[4357]), .B(x[4357]), .Z(n27694) );
  XNOR U36416 ( .A(y[4358]), .B(x[4358]), .Z(n27693) );
  XNOR U36417 ( .A(y[4356]), .B(x[4356]), .Z(n27691) );
  XNOR U36418 ( .A(n27685), .B(n27686), .Z(n27696) );
  XNOR U36419 ( .A(y[4353]), .B(x[4353]), .Z(n27686) );
  XNOR U36420 ( .A(n27687), .B(n27688), .Z(n27685) );
  XNOR U36421 ( .A(y[4354]), .B(x[4354]), .Z(n27688) );
  XNOR U36422 ( .A(y[4355]), .B(x[4355]), .Z(n27687) );
  XNOR U36423 ( .A(n27678), .B(n27677), .Z(n27681) );
  XNOR U36424 ( .A(n27673), .B(n27674), .Z(n27677) );
  XNOR U36425 ( .A(y[4350]), .B(x[4350]), .Z(n27674) );
  XNOR U36426 ( .A(n27675), .B(n27676), .Z(n27673) );
  XNOR U36427 ( .A(y[4351]), .B(x[4351]), .Z(n27676) );
  XNOR U36428 ( .A(y[4352]), .B(x[4352]), .Z(n27675) );
  XNOR U36429 ( .A(n27667), .B(n27668), .Z(n27678) );
  XNOR U36430 ( .A(y[4347]), .B(x[4347]), .Z(n27668) );
  XNOR U36431 ( .A(n27669), .B(n27670), .Z(n27667) );
  XNOR U36432 ( .A(y[4348]), .B(x[4348]), .Z(n27670) );
  XNOR U36433 ( .A(y[4349]), .B(x[4349]), .Z(n27669) );
  XOR U36434 ( .A(n27643), .B(n27644), .Z(n27662) );
  XNOR U36435 ( .A(n27659), .B(n27660), .Z(n27644) );
  XNOR U36436 ( .A(n27654), .B(n27655), .Z(n27660) );
  XNOR U36437 ( .A(n27656), .B(n27657), .Z(n27655) );
  XNOR U36438 ( .A(y[4345]), .B(x[4345]), .Z(n27657) );
  XNOR U36439 ( .A(y[4346]), .B(x[4346]), .Z(n27656) );
  XNOR U36440 ( .A(y[4344]), .B(x[4344]), .Z(n27654) );
  XNOR U36441 ( .A(n27648), .B(n27649), .Z(n27659) );
  XNOR U36442 ( .A(y[4341]), .B(x[4341]), .Z(n27649) );
  XNOR U36443 ( .A(n27650), .B(n27651), .Z(n27648) );
  XNOR U36444 ( .A(y[4342]), .B(x[4342]), .Z(n27651) );
  XNOR U36445 ( .A(y[4343]), .B(x[4343]), .Z(n27650) );
  XOR U36446 ( .A(n27642), .B(n27641), .Z(n27643) );
  XNOR U36447 ( .A(n27637), .B(n27638), .Z(n27641) );
  XNOR U36448 ( .A(y[4338]), .B(x[4338]), .Z(n27638) );
  XNOR U36449 ( .A(n27639), .B(n27640), .Z(n27637) );
  XNOR U36450 ( .A(y[4339]), .B(x[4339]), .Z(n27640) );
  XNOR U36451 ( .A(y[4340]), .B(x[4340]), .Z(n27639) );
  XNOR U36452 ( .A(n27631), .B(n27632), .Z(n27642) );
  XNOR U36453 ( .A(y[4335]), .B(x[4335]), .Z(n27632) );
  XNOR U36454 ( .A(n27633), .B(n27634), .Z(n27631) );
  XNOR U36455 ( .A(y[4336]), .B(x[4336]), .Z(n27634) );
  XNOR U36456 ( .A(y[4337]), .B(x[4337]), .Z(n27633) );
  NAND U36457 ( .A(n27698), .B(n27699), .Z(N62936) );
  NANDN U36458 ( .A(n27700), .B(n27701), .Z(n27699) );
  OR U36459 ( .A(n27702), .B(n27703), .Z(n27701) );
  NAND U36460 ( .A(n27702), .B(n27703), .Z(n27698) );
  XOR U36461 ( .A(n27702), .B(n27704), .Z(N62935) );
  XNOR U36462 ( .A(n27700), .B(n27703), .Z(n27704) );
  AND U36463 ( .A(n27705), .B(n27706), .Z(n27703) );
  NANDN U36464 ( .A(n27707), .B(n27708), .Z(n27706) );
  NANDN U36465 ( .A(n27709), .B(n27710), .Z(n27708) );
  NANDN U36466 ( .A(n27710), .B(n27709), .Z(n27705) );
  NAND U36467 ( .A(n27711), .B(n27712), .Z(n27700) );
  NANDN U36468 ( .A(n27713), .B(n27714), .Z(n27712) );
  OR U36469 ( .A(n27715), .B(n27716), .Z(n27714) );
  NAND U36470 ( .A(n27716), .B(n27715), .Z(n27711) );
  AND U36471 ( .A(n27717), .B(n27718), .Z(n27702) );
  NANDN U36472 ( .A(n27719), .B(n27720), .Z(n27718) );
  NANDN U36473 ( .A(n27721), .B(n27722), .Z(n27720) );
  NANDN U36474 ( .A(n27722), .B(n27721), .Z(n27717) );
  XOR U36475 ( .A(n27716), .B(n27723), .Z(N62934) );
  XOR U36476 ( .A(n27713), .B(n27715), .Z(n27723) );
  XNOR U36477 ( .A(n27709), .B(n27724), .Z(n27715) );
  XNOR U36478 ( .A(n27707), .B(n27710), .Z(n27724) );
  NAND U36479 ( .A(n27725), .B(n27726), .Z(n27710) );
  NAND U36480 ( .A(n27727), .B(n27728), .Z(n27726) );
  OR U36481 ( .A(n27729), .B(n27730), .Z(n27727) );
  NANDN U36482 ( .A(n27731), .B(n27729), .Z(n27725) );
  IV U36483 ( .A(n27730), .Z(n27731) );
  NAND U36484 ( .A(n27732), .B(n27733), .Z(n27707) );
  NAND U36485 ( .A(n27734), .B(n27735), .Z(n27733) );
  NANDN U36486 ( .A(n27736), .B(n27737), .Z(n27734) );
  NANDN U36487 ( .A(n27737), .B(n27736), .Z(n27732) );
  AND U36488 ( .A(n27738), .B(n27739), .Z(n27709) );
  NAND U36489 ( .A(n27740), .B(n27741), .Z(n27739) );
  OR U36490 ( .A(n27742), .B(n27743), .Z(n27740) );
  NANDN U36491 ( .A(n27744), .B(n27742), .Z(n27738) );
  NAND U36492 ( .A(n27745), .B(n27746), .Z(n27713) );
  NANDN U36493 ( .A(n27747), .B(n27748), .Z(n27746) );
  OR U36494 ( .A(n27749), .B(n27750), .Z(n27748) );
  NANDN U36495 ( .A(n27751), .B(n27749), .Z(n27745) );
  IV U36496 ( .A(n27750), .Z(n27751) );
  XNOR U36497 ( .A(n27721), .B(n27752), .Z(n27716) );
  XNOR U36498 ( .A(n27719), .B(n27722), .Z(n27752) );
  NAND U36499 ( .A(n27753), .B(n27754), .Z(n27722) );
  NAND U36500 ( .A(n27755), .B(n27756), .Z(n27754) );
  OR U36501 ( .A(n27757), .B(n27758), .Z(n27755) );
  NANDN U36502 ( .A(n27759), .B(n27757), .Z(n27753) );
  IV U36503 ( .A(n27758), .Z(n27759) );
  NAND U36504 ( .A(n27760), .B(n27761), .Z(n27719) );
  NAND U36505 ( .A(n27762), .B(n27763), .Z(n27761) );
  NANDN U36506 ( .A(n27764), .B(n27765), .Z(n27762) );
  NANDN U36507 ( .A(n27765), .B(n27764), .Z(n27760) );
  AND U36508 ( .A(n27766), .B(n27767), .Z(n27721) );
  NAND U36509 ( .A(n27768), .B(n27769), .Z(n27767) );
  OR U36510 ( .A(n27770), .B(n27771), .Z(n27768) );
  NANDN U36511 ( .A(n27772), .B(n27770), .Z(n27766) );
  XNOR U36512 ( .A(n27747), .B(n27773), .Z(N62933) );
  XOR U36513 ( .A(n27749), .B(n27750), .Z(n27773) );
  XNOR U36514 ( .A(n27763), .B(n27774), .Z(n27750) );
  XOR U36515 ( .A(n27764), .B(n27765), .Z(n27774) );
  XOR U36516 ( .A(n27770), .B(n27775), .Z(n27765) );
  XOR U36517 ( .A(n27769), .B(n27772), .Z(n27775) );
  IV U36518 ( .A(n27771), .Z(n27772) );
  NAND U36519 ( .A(n27776), .B(n27777), .Z(n27771) );
  OR U36520 ( .A(n27778), .B(n27779), .Z(n27777) );
  OR U36521 ( .A(n27780), .B(n27781), .Z(n27776) );
  NAND U36522 ( .A(n27782), .B(n27783), .Z(n27769) );
  OR U36523 ( .A(n27784), .B(n27785), .Z(n27783) );
  OR U36524 ( .A(n27786), .B(n27787), .Z(n27782) );
  NOR U36525 ( .A(n27788), .B(n27789), .Z(n27770) );
  ANDN U36526 ( .B(n27790), .A(n27791), .Z(n27764) );
  XNOR U36527 ( .A(n27757), .B(n27792), .Z(n27763) );
  XNOR U36528 ( .A(n27756), .B(n27758), .Z(n27792) );
  NAND U36529 ( .A(n27793), .B(n27794), .Z(n27758) );
  OR U36530 ( .A(n27795), .B(n27796), .Z(n27794) );
  OR U36531 ( .A(n27797), .B(n27798), .Z(n27793) );
  NAND U36532 ( .A(n27799), .B(n27800), .Z(n27756) );
  OR U36533 ( .A(n27801), .B(n27802), .Z(n27800) );
  OR U36534 ( .A(n27803), .B(n27804), .Z(n27799) );
  ANDN U36535 ( .B(n27805), .A(n27806), .Z(n27757) );
  IV U36536 ( .A(n27807), .Z(n27805) );
  ANDN U36537 ( .B(n27808), .A(n27809), .Z(n27749) );
  XOR U36538 ( .A(n27735), .B(n27810), .Z(n27747) );
  XOR U36539 ( .A(n27736), .B(n27737), .Z(n27810) );
  XOR U36540 ( .A(n27742), .B(n27811), .Z(n27737) );
  XOR U36541 ( .A(n27741), .B(n27744), .Z(n27811) );
  IV U36542 ( .A(n27743), .Z(n27744) );
  NAND U36543 ( .A(n27812), .B(n27813), .Z(n27743) );
  OR U36544 ( .A(n27814), .B(n27815), .Z(n27813) );
  OR U36545 ( .A(n27816), .B(n27817), .Z(n27812) );
  NAND U36546 ( .A(n27818), .B(n27819), .Z(n27741) );
  OR U36547 ( .A(n27820), .B(n27821), .Z(n27819) );
  OR U36548 ( .A(n27822), .B(n27823), .Z(n27818) );
  NOR U36549 ( .A(n27824), .B(n27825), .Z(n27742) );
  ANDN U36550 ( .B(n27826), .A(n27827), .Z(n27736) );
  IV U36551 ( .A(n27828), .Z(n27826) );
  XNOR U36552 ( .A(n27729), .B(n27829), .Z(n27735) );
  XNOR U36553 ( .A(n27728), .B(n27730), .Z(n27829) );
  NAND U36554 ( .A(n27830), .B(n27831), .Z(n27730) );
  OR U36555 ( .A(n27832), .B(n27833), .Z(n27831) );
  OR U36556 ( .A(n27834), .B(n27835), .Z(n27830) );
  NAND U36557 ( .A(n27836), .B(n27837), .Z(n27728) );
  OR U36558 ( .A(n27838), .B(n27839), .Z(n27837) );
  OR U36559 ( .A(n27840), .B(n27841), .Z(n27836) );
  ANDN U36560 ( .B(n27842), .A(n27843), .Z(n27729) );
  IV U36561 ( .A(n27844), .Z(n27842) );
  XNOR U36562 ( .A(n27809), .B(n27808), .Z(N62932) );
  XOR U36563 ( .A(n27828), .B(n27827), .Z(n27808) );
  XNOR U36564 ( .A(n27843), .B(n27844), .Z(n27827) );
  XNOR U36565 ( .A(n27838), .B(n27839), .Z(n27844) );
  XNOR U36566 ( .A(n27840), .B(n27841), .Z(n27839) );
  XNOR U36567 ( .A(y[4333]), .B(x[4333]), .Z(n27841) );
  XNOR U36568 ( .A(y[4334]), .B(x[4334]), .Z(n27840) );
  XNOR U36569 ( .A(y[4332]), .B(x[4332]), .Z(n27838) );
  XNOR U36570 ( .A(n27832), .B(n27833), .Z(n27843) );
  XNOR U36571 ( .A(y[4329]), .B(x[4329]), .Z(n27833) );
  XNOR U36572 ( .A(n27834), .B(n27835), .Z(n27832) );
  XNOR U36573 ( .A(y[4330]), .B(x[4330]), .Z(n27835) );
  XNOR U36574 ( .A(y[4331]), .B(x[4331]), .Z(n27834) );
  XNOR U36575 ( .A(n27825), .B(n27824), .Z(n27828) );
  XNOR U36576 ( .A(n27820), .B(n27821), .Z(n27824) );
  XNOR U36577 ( .A(y[4326]), .B(x[4326]), .Z(n27821) );
  XNOR U36578 ( .A(n27822), .B(n27823), .Z(n27820) );
  XNOR U36579 ( .A(y[4327]), .B(x[4327]), .Z(n27823) );
  XNOR U36580 ( .A(y[4328]), .B(x[4328]), .Z(n27822) );
  XNOR U36581 ( .A(n27814), .B(n27815), .Z(n27825) );
  XNOR U36582 ( .A(y[4323]), .B(x[4323]), .Z(n27815) );
  XNOR U36583 ( .A(n27816), .B(n27817), .Z(n27814) );
  XNOR U36584 ( .A(y[4324]), .B(x[4324]), .Z(n27817) );
  XNOR U36585 ( .A(y[4325]), .B(x[4325]), .Z(n27816) );
  XOR U36586 ( .A(n27790), .B(n27791), .Z(n27809) );
  XNOR U36587 ( .A(n27806), .B(n27807), .Z(n27791) );
  XNOR U36588 ( .A(n27801), .B(n27802), .Z(n27807) );
  XNOR U36589 ( .A(n27803), .B(n27804), .Z(n27802) );
  XNOR U36590 ( .A(y[4321]), .B(x[4321]), .Z(n27804) );
  XNOR U36591 ( .A(y[4322]), .B(x[4322]), .Z(n27803) );
  XNOR U36592 ( .A(y[4320]), .B(x[4320]), .Z(n27801) );
  XNOR U36593 ( .A(n27795), .B(n27796), .Z(n27806) );
  XNOR U36594 ( .A(y[4317]), .B(x[4317]), .Z(n27796) );
  XNOR U36595 ( .A(n27797), .B(n27798), .Z(n27795) );
  XNOR U36596 ( .A(y[4318]), .B(x[4318]), .Z(n27798) );
  XNOR U36597 ( .A(y[4319]), .B(x[4319]), .Z(n27797) );
  XOR U36598 ( .A(n27789), .B(n27788), .Z(n27790) );
  XNOR U36599 ( .A(n27784), .B(n27785), .Z(n27788) );
  XNOR U36600 ( .A(y[4314]), .B(x[4314]), .Z(n27785) );
  XNOR U36601 ( .A(n27786), .B(n27787), .Z(n27784) );
  XNOR U36602 ( .A(y[4315]), .B(x[4315]), .Z(n27787) );
  XNOR U36603 ( .A(y[4316]), .B(x[4316]), .Z(n27786) );
  XNOR U36604 ( .A(n27778), .B(n27779), .Z(n27789) );
  XNOR U36605 ( .A(y[4311]), .B(x[4311]), .Z(n27779) );
  XNOR U36606 ( .A(n27780), .B(n27781), .Z(n27778) );
  XNOR U36607 ( .A(y[4312]), .B(x[4312]), .Z(n27781) );
  XNOR U36608 ( .A(y[4313]), .B(x[4313]), .Z(n27780) );
  NAND U36609 ( .A(n27845), .B(n27846), .Z(N62923) );
  NANDN U36610 ( .A(n27847), .B(n27848), .Z(n27846) );
  OR U36611 ( .A(n27849), .B(n27850), .Z(n27848) );
  NAND U36612 ( .A(n27849), .B(n27850), .Z(n27845) );
  XOR U36613 ( .A(n27849), .B(n27851), .Z(N62922) );
  XNOR U36614 ( .A(n27847), .B(n27850), .Z(n27851) );
  AND U36615 ( .A(n27852), .B(n27853), .Z(n27850) );
  NANDN U36616 ( .A(n27854), .B(n27855), .Z(n27853) );
  NANDN U36617 ( .A(n27856), .B(n27857), .Z(n27855) );
  NANDN U36618 ( .A(n27857), .B(n27856), .Z(n27852) );
  NAND U36619 ( .A(n27858), .B(n27859), .Z(n27847) );
  NANDN U36620 ( .A(n27860), .B(n27861), .Z(n27859) );
  OR U36621 ( .A(n27862), .B(n27863), .Z(n27861) );
  NAND U36622 ( .A(n27863), .B(n27862), .Z(n27858) );
  AND U36623 ( .A(n27864), .B(n27865), .Z(n27849) );
  NANDN U36624 ( .A(n27866), .B(n27867), .Z(n27865) );
  NANDN U36625 ( .A(n27868), .B(n27869), .Z(n27867) );
  NANDN U36626 ( .A(n27869), .B(n27868), .Z(n27864) );
  XOR U36627 ( .A(n27863), .B(n27870), .Z(N62921) );
  XOR U36628 ( .A(n27860), .B(n27862), .Z(n27870) );
  XNOR U36629 ( .A(n27856), .B(n27871), .Z(n27862) );
  XNOR U36630 ( .A(n27854), .B(n27857), .Z(n27871) );
  NAND U36631 ( .A(n27872), .B(n27873), .Z(n27857) );
  NAND U36632 ( .A(n27874), .B(n27875), .Z(n27873) );
  OR U36633 ( .A(n27876), .B(n27877), .Z(n27874) );
  NANDN U36634 ( .A(n27878), .B(n27876), .Z(n27872) );
  IV U36635 ( .A(n27877), .Z(n27878) );
  NAND U36636 ( .A(n27879), .B(n27880), .Z(n27854) );
  NAND U36637 ( .A(n27881), .B(n27882), .Z(n27880) );
  NANDN U36638 ( .A(n27883), .B(n27884), .Z(n27881) );
  NANDN U36639 ( .A(n27884), .B(n27883), .Z(n27879) );
  AND U36640 ( .A(n27885), .B(n27886), .Z(n27856) );
  NAND U36641 ( .A(n27887), .B(n27888), .Z(n27886) );
  OR U36642 ( .A(n27889), .B(n27890), .Z(n27887) );
  NANDN U36643 ( .A(n27891), .B(n27889), .Z(n27885) );
  NAND U36644 ( .A(n27892), .B(n27893), .Z(n27860) );
  NANDN U36645 ( .A(n27894), .B(n27895), .Z(n27893) );
  OR U36646 ( .A(n27896), .B(n27897), .Z(n27895) );
  NANDN U36647 ( .A(n27898), .B(n27896), .Z(n27892) );
  IV U36648 ( .A(n27897), .Z(n27898) );
  XNOR U36649 ( .A(n27868), .B(n27899), .Z(n27863) );
  XNOR U36650 ( .A(n27866), .B(n27869), .Z(n27899) );
  NAND U36651 ( .A(n27900), .B(n27901), .Z(n27869) );
  NAND U36652 ( .A(n27902), .B(n27903), .Z(n27901) );
  OR U36653 ( .A(n27904), .B(n27905), .Z(n27902) );
  NANDN U36654 ( .A(n27906), .B(n27904), .Z(n27900) );
  IV U36655 ( .A(n27905), .Z(n27906) );
  NAND U36656 ( .A(n27907), .B(n27908), .Z(n27866) );
  NAND U36657 ( .A(n27909), .B(n27910), .Z(n27908) );
  NANDN U36658 ( .A(n27911), .B(n27912), .Z(n27909) );
  NANDN U36659 ( .A(n27912), .B(n27911), .Z(n27907) );
  AND U36660 ( .A(n27913), .B(n27914), .Z(n27868) );
  NAND U36661 ( .A(n27915), .B(n27916), .Z(n27914) );
  OR U36662 ( .A(n27917), .B(n27918), .Z(n27915) );
  NANDN U36663 ( .A(n27919), .B(n27917), .Z(n27913) );
  XNOR U36664 ( .A(n27894), .B(n27920), .Z(N62920) );
  XOR U36665 ( .A(n27896), .B(n27897), .Z(n27920) );
  XNOR U36666 ( .A(n27910), .B(n27921), .Z(n27897) );
  XOR U36667 ( .A(n27911), .B(n27912), .Z(n27921) );
  XOR U36668 ( .A(n27917), .B(n27922), .Z(n27912) );
  XOR U36669 ( .A(n27916), .B(n27919), .Z(n27922) );
  IV U36670 ( .A(n27918), .Z(n27919) );
  NAND U36671 ( .A(n27923), .B(n27924), .Z(n27918) );
  OR U36672 ( .A(n27925), .B(n27926), .Z(n27924) );
  OR U36673 ( .A(n27927), .B(n27928), .Z(n27923) );
  NAND U36674 ( .A(n27929), .B(n27930), .Z(n27916) );
  OR U36675 ( .A(n27931), .B(n27932), .Z(n27930) );
  OR U36676 ( .A(n27933), .B(n27934), .Z(n27929) );
  NOR U36677 ( .A(n27935), .B(n27936), .Z(n27917) );
  ANDN U36678 ( .B(n27937), .A(n27938), .Z(n27911) );
  XNOR U36679 ( .A(n27904), .B(n27939), .Z(n27910) );
  XNOR U36680 ( .A(n27903), .B(n27905), .Z(n27939) );
  NAND U36681 ( .A(n27940), .B(n27941), .Z(n27905) );
  OR U36682 ( .A(n27942), .B(n27943), .Z(n27941) );
  OR U36683 ( .A(n27944), .B(n27945), .Z(n27940) );
  NAND U36684 ( .A(n27946), .B(n27947), .Z(n27903) );
  OR U36685 ( .A(n27948), .B(n27949), .Z(n27947) );
  OR U36686 ( .A(n27950), .B(n27951), .Z(n27946) );
  ANDN U36687 ( .B(n27952), .A(n27953), .Z(n27904) );
  IV U36688 ( .A(n27954), .Z(n27952) );
  ANDN U36689 ( .B(n27955), .A(n27956), .Z(n27896) );
  XOR U36690 ( .A(n27882), .B(n27957), .Z(n27894) );
  XOR U36691 ( .A(n27883), .B(n27884), .Z(n27957) );
  XOR U36692 ( .A(n27889), .B(n27958), .Z(n27884) );
  XOR U36693 ( .A(n27888), .B(n27891), .Z(n27958) );
  IV U36694 ( .A(n27890), .Z(n27891) );
  NAND U36695 ( .A(n27959), .B(n27960), .Z(n27890) );
  OR U36696 ( .A(n27961), .B(n27962), .Z(n27960) );
  OR U36697 ( .A(n27963), .B(n27964), .Z(n27959) );
  NAND U36698 ( .A(n27965), .B(n27966), .Z(n27888) );
  OR U36699 ( .A(n27967), .B(n27968), .Z(n27966) );
  OR U36700 ( .A(n27969), .B(n27970), .Z(n27965) );
  NOR U36701 ( .A(n27971), .B(n27972), .Z(n27889) );
  ANDN U36702 ( .B(n27973), .A(n27974), .Z(n27883) );
  IV U36703 ( .A(n27975), .Z(n27973) );
  XNOR U36704 ( .A(n27876), .B(n27976), .Z(n27882) );
  XNOR U36705 ( .A(n27875), .B(n27877), .Z(n27976) );
  NAND U36706 ( .A(n27977), .B(n27978), .Z(n27877) );
  OR U36707 ( .A(n27979), .B(n27980), .Z(n27978) );
  OR U36708 ( .A(n27981), .B(n27982), .Z(n27977) );
  NAND U36709 ( .A(n27983), .B(n27984), .Z(n27875) );
  OR U36710 ( .A(n27985), .B(n27986), .Z(n27984) );
  OR U36711 ( .A(n27987), .B(n27988), .Z(n27983) );
  ANDN U36712 ( .B(n27989), .A(n27990), .Z(n27876) );
  IV U36713 ( .A(n27991), .Z(n27989) );
  XNOR U36714 ( .A(n27956), .B(n27955), .Z(N62919) );
  XOR U36715 ( .A(n27975), .B(n27974), .Z(n27955) );
  XNOR U36716 ( .A(n27990), .B(n27991), .Z(n27974) );
  XNOR U36717 ( .A(n27985), .B(n27986), .Z(n27991) );
  XNOR U36718 ( .A(n27987), .B(n27988), .Z(n27986) );
  XNOR U36719 ( .A(y[4309]), .B(x[4309]), .Z(n27988) );
  XNOR U36720 ( .A(y[4310]), .B(x[4310]), .Z(n27987) );
  XNOR U36721 ( .A(y[4308]), .B(x[4308]), .Z(n27985) );
  XNOR U36722 ( .A(n27979), .B(n27980), .Z(n27990) );
  XNOR U36723 ( .A(y[4305]), .B(x[4305]), .Z(n27980) );
  XNOR U36724 ( .A(n27981), .B(n27982), .Z(n27979) );
  XNOR U36725 ( .A(y[4306]), .B(x[4306]), .Z(n27982) );
  XNOR U36726 ( .A(y[4307]), .B(x[4307]), .Z(n27981) );
  XNOR U36727 ( .A(n27972), .B(n27971), .Z(n27975) );
  XNOR U36728 ( .A(n27967), .B(n27968), .Z(n27971) );
  XNOR U36729 ( .A(y[4302]), .B(x[4302]), .Z(n27968) );
  XNOR U36730 ( .A(n27969), .B(n27970), .Z(n27967) );
  XNOR U36731 ( .A(y[4303]), .B(x[4303]), .Z(n27970) );
  XNOR U36732 ( .A(y[4304]), .B(x[4304]), .Z(n27969) );
  XNOR U36733 ( .A(n27961), .B(n27962), .Z(n27972) );
  XNOR U36734 ( .A(y[4299]), .B(x[4299]), .Z(n27962) );
  XNOR U36735 ( .A(n27963), .B(n27964), .Z(n27961) );
  XNOR U36736 ( .A(y[4300]), .B(x[4300]), .Z(n27964) );
  XNOR U36737 ( .A(y[4301]), .B(x[4301]), .Z(n27963) );
  XOR U36738 ( .A(n27937), .B(n27938), .Z(n27956) );
  XNOR U36739 ( .A(n27953), .B(n27954), .Z(n27938) );
  XNOR U36740 ( .A(n27948), .B(n27949), .Z(n27954) );
  XNOR U36741 ( .A(n27950), .B(n27951), .Z(n27949) );
  XNOR U36742 ( .A(y[4297]), .B(x[4297]), .Z(n27951) );
  XNOR U36743 ( .A(y[4298]), .B(x[4298]), .Z(n27950) );
  XNOR U36744 ( .A(y[4296]), .B(x[4296]), .Z(n27948) );
  XNOR U36745 ( .A(n27942), .B(n27943), .Z(n27953) );
  XNOR U36746 ( .A(y[4293]), .B(x[4293]), .Z(n27943) );
  XNOR U36747 ( .A(n27944), .B(n27945), .Z(n27942) );
  XNOR U36748 ( .A(y[4294]), .B(x[4294]), .Z(n27945) );
  XNOR U36749 ( .A(y[4295]), .B(x[4295]), .Z(n27944) );
  XOR U36750 ( .A(n27936), .B(n27935), .Z(n27937) );
  XNOR U36751 ( .A(n27931), .B(n27932), .Z(n27935) );
  XNOR U36752 ( .A(y[4290]), .B(x[4290]), .Z(n27932) );
  XNOR U36753 ( .A(n27933), .B(n27934), .Z(n27931) );
  XNOR U36754 ( .A(y[4291]), .B(x[4291]), .Z(n27934) );
  XNOR U36755 ( .A(y[4292]), .B(x[4292]), .Z(n27933) );
  XNOR U36756 ( .A(n27925), .B(n27926), .Z(n27936) );
  XNOR U36757 ( .A(y[4287]), .B(x[4287]), .Z(n27926) );
  XNOR U36758 ( .A(n27927), .B(n27928), .Z(n27925) );
  XNOR U36759 ( .A(y[4288]), .B(x[4288]), .Z(n27928) );
  XNOR U36760 ( .A(y[4289]), .B(x[4289]), .Z(n27927) );
  NAND U36761 ( .A(n27992), .B(n27993), .Z(N62910) );
  NANDN U36762 ( .A(n27994), .B(n27995), .Z(n27993) );
  OR U36763 ( .A(n27996), .B(n27997), .Z(n27995) );
  NAND U36764 ( .A(n27996), .B(n27997), .Z(n27992) );
  XOR U36765 ( .A(n27996), .B(n27998), .Z(N62909) );
  XNOR U36766 ( .A(n27994), .B(n27997), .Z(n27998) );
  AND U36767 ( .A(n27999), .B(n28000), .Z(n27997) );
  NANDN U36768 ( .A(n28001), .B(n28002), .Z(n28000) );
  NANDN U36769 ( .A(n28003), .B(n28004), .Z(n28002) );
  NANDN U36770 ( .A(n28004), .B(n28003), .Z(n27999) );
  NAND U36771 ( .A(n28005), .B(n28006), .Z(n27994) );
  NANDN U36772 ( .A(n28007), .B(n28008), .Z(n28006) );
  OR U36773 ( .A(n28009), .B(n28010), .Z(n28008) );
  NAND U36774 ( .A(n28010), .B(n28009), .Z(n28005) );
  AND U36775 ( .A(n28011), .B(n28012), .Z(n27996) );
  NANDN U36776 ( .A(n28013), .B(n28014), .Z(n28012) );
  NANDN U36777 ( .A(n28015), .B(n28016), .Z(n28014) );
  NANDN U36778 ( .A(n28016), .B(n28015), .Z(n28011) );
  XOR U36779 ( .A(n28010), .B(n28017), .Z(N62908) );
  XOR U36780 ( .A(n28007), .B(n28009), .Z(n28017) );
  XNOR U36781 ( .A(n28003), .B(n28018), .Z(n28009) );
  XNOR U36782 ( .A(n28001), .B(n28004), .Z(n28018) );
  NAND U36783 ( .A(n28019), .B(n28020), .Z(n28004) );
  NAND U36784 ( .A(n28021), .B(n28022), .Z(n28020) );
  OR U36785 ( .A(n28023), .B(n28024), .Z(n28021) );
  NANDN U36786 ( .A(n28025), .B(n28023), .Z(n28019) );
  IV U36787 ( .A(n28024), .Z(n28025) );
  NAND U36788 ( .A(n28026), .B(n28027), .Z(n28001) );
  NAND U36789 ( .A(n28028), .B(n28029), .Z(n28027) );
  NANDN U36790 ( .A(n28030), .B(n28031), .Z(n28028) );
  NANDN U36791 ( .A(n28031), .B(n28030), .Z(n28026) );
  AND U36792 ( .A(n28032), .B(n28033), .Z(n28003) );
  NAND U36793 ( .A(n28034), .B(n28035), .Z(n28033) );
  OR U36794 ( .A(n28036), .B(n28037), .Z(n28034) );
  NANDN U36795 ( .A(n28038), .B(n28036), .Z(n28032) );
  NAND U36796 ( .A(n28039), .B(n28040), .Z(n28007) );
  NANDN U36797 ( .A(n28041), .B(n28042), .Z(n28040) );
  OR U36798 ( .A(n28043), .B(n28044), .Z(n28042) );
  NANDN U36799 ( .A(n28045), .B(n28043), .Z(n28039) );
  IV U36800 ( .A(n28044), .Z(n28045) );
  XNOR U36801 ( .A(n28015), .B(n28046), .Z(n28010) );
  XNOR U36802 ( .A(n28013), .B(n28016), .Z(n28046) );
  NAND U36803 ( .A(n28047), .B(n28048), .Z(n28016) );
  NAND U36804 ( .A(n28049), .B(n28050), .Z(n28048) );
  OR U36805 ( .A(n28051), .B(n28052), .Z(n28049) );
  NANDN U36806 ( .A(n28053), .B(n28051), .Z(n28047) );
  IV U36807 ( .A(n28052), .Z(n28053) );
  NAND U36808 ( .A(n28054), .B(n28055), .Z(n28013) );
  NAND U36809 ( .A(n28056), .B(n28057), .Z(n28055) );
  NANDN U36810 ( .A(n28058), .B(n28059), .Z(n28056) );
  NANDN U36811 ( .A(n28059), .B(n28058), .Z(n28054) );
  AND U36812 ( .A(n28060), .B(n28061), .Z(n28015) );
  NAND U36813 ( .A(n28062), .B(n28063), .Z(n28061) );
  OR U36814 ( .A(n28064), .B(n28065), .Z(n28062) );
  NANDN U36815 ( .A(n28066), .B(n28064), .Z(n28060) );
  XNOR U36816 ( .A(n28041), .B(n28067), .Z(N62907) );
  XOR U36817 ( .A(n28043), .B(n28044), .Z(n28067) );
  XNOR U36818 ( .A(n28057), .B(n28068), .Z(n28044) );
  XOR U36819 ( .A(n28058), .B(n28059), .Z(n28068) );
  XOR U36820 ( .A(n28064), .B(n28069), .Z(n28059) );
  XOR U36821 ( .A(n28063), .B(n28066), .Z(n28069) );
  IV U36822 ( .A(n28065), .Z(n28066) );
  NAND U36823 ( .A(n28070), .B(n28071), .Z(n28065) );
  OR U36824 ( .A(n28072), .B(n28073), .Z(n28071) );
  OR U36825 ( .A(n28074), .B(n28075), .Z(n28070) );
  NAND U36826 ( .A(n28076), .B(n28077), .Z(n28063) );
  OR U36827 ( .A(n28078), .B(n28079), .Z(n28077) );
  OR U36828 ( .A(n28080), .B(n28081), .Z(n28076) );
  NOR U36829 ( .A(n28082), .B(n28083), .Z(n28064) );
  ANDN U36830 ( .B(n28084), .A(n28085), .Z(n28058) );
  XNOR U36831 ( .A(n28051), .B(n28086), .Z(n28057) );
  XNOR U36832 ( .A(n28050), .B(n28052), .Z(n28086) );
  NAND U36833 ( .A(n28087), .B(n28088), .Z(n28052) );
  OR U36834 ( .A(n28089), .B(n28090), .Z(n28088) );
  OR U36835 ( .A(n28091), .B(n28092), .Z(n28087) );
  NAND U36836 ( .A(n28093), .B(n28094), .Z(n28050) );
  OR U36837 ( .A(n28095), .B(n28096), .Z(n28094) );
  OR U36838 ( .A(n28097), .B(n28098), .Z(n28093) );
  ANDN U36839 ( .B(n28099), .A(n28100), .Z(n28051) );
  IV U36840 ( .A(n28101), .Z(n28099) );
  ANDN U36841 ( .B(n28102), .A(n28103), .Z(n28043) );
  XOR U36842 ( .A(n28029), .B(n28104), .Z(n28041) );
  XOR U36843 ( .A(n28030), .B(n28031), .Z(n28104) );
  XOR U36844 ( .A(n28036), .B(n28105), .Z(n28031) );
  XOR U36845 ( .A(n28035), .B(n28038), .Z(n28105) );
  IV U36846 ( .A(n28037), .Z(n28038) );
  NAND U36847 ( .A(n28106), .B(n28107), .Z(n28037) );
  OR U36848 ( .A(n28108), .B(n28109), .Z(n28107) );
  OR U36849 ( .A(n28110), .B(n28111), .Z(n28106) );
  NAND U36850 ( .A(n28112), .B(n28113), .Z(n28035) );
  OR U36851 ( .A(n28114), .B(n28115), .Z(n28113) );
  OR U36852 ( .A(n28116), .B(n28117), .Z(n28112) );
  NOR U36853 ( .A(n28118), .B(n28119), .Z(n28036) );
  ANDN U36854 ( .B(n28120), .A(n28121), .Z(n28030) );
  IV U36855 ( .A(n28122), .Z(n28120) );
  XNOR U36856 ( .A(n28023), .B(n28123), .Z(n28029) );
  XNOR U36857 ( .A(n28022), .B(n28024), .Z(n28123) );
  NAND U36858 ( .A(n28124), .B(n28125), .Z(n28024) );
  OR U36859 ( .A(n28126), .B(n28127), .Z(n28125) );
  OR U36860 ( .A(n28128), .B(n28129), .Z(n28124) );
  NAND U36861 ( .A(n28130), .B(n28131), .Z(n28022) );
  OR U36862 ( .A(n28132), .B(n28133), .Z(n28131) );
  OR U36863 ( .A(n28134), .B(n28135), .Z(n28130) );
  ANDN U36864 ( .B(n28136), .A(n28137), .Z(n28023) );
  IV U36865 ( .A(n28138), .Z(n28136) );
  XNOR U36866 ( .A(n28103), .B(n28102), .Z(N62906) );
  XOR U36867 ( .A(n28122), .B(n28121), .Z(n28102) );
  XNOR U36868 ( .A(n28137), .B(n28138), .Z(n28121) );
  XNOR U36869 ( .A(n28132), .B(n28133), .Z(n28138) );
  XNOR U36870 ( .A(n28134), .B(n28135), .Z(n28133) );
  XNOR U36871 ( .A(y[4285]), .B(x[4285]), .Z(n28135) );
  XNOR U36872 ( .A(y[4286]), .B(x[4286]), .Z(n28134) );
  XNOR U36873 ( .A(y[4284]), .B(x[4284]), .Z(n28132) );
  XNOR U36874 ( .A(n28126), .B(n28127), .Z(n28137) );
  XNOR U36875 ( .A(y[4281]), .B(x[4281]), .Z(n28127) );
  XNOR U36876 ( .A(n28128), .B(n28129), .Z(n28126) );
  XNOR U36877 ( .A(y[4282]), .B(x[4282]), .Z(n28129) );
  XNOR U36878 ( .A(y[4283]), .B(x[4283]), .Z(n28128) );
  XNOR U36879 ( .A(n28119), .B(n28118), .Z(n28122) );
  XNOR U36880 ( .A(n28114), .B(n28115), .Z(n28118) );
  XNOR U36881 ( .A(y[4278]), .B(x[4278]), .Z(n28115) );
  XNOR U36882 ( .A(n28116), .B(n28117), .Z(n28114) );
  XNOR U36883 ( .A(y[4279]), .B(x[4279]), .Z(n28117) );
  XNOR U36884 ( .A(y[4280]), .B(x[4280]), .Z(n28116) );
  XNOR U36885 ( .A(n28108), .B(n28109), .Z(n28119) );
  XNOR U36886 ( .A(y[4275]), .B(x[4275]), .Z(n28109) );
  XNOR U36887 ( .A(n28110), .B(n28111), .Z(n28108) );
  XNOR U36888 ( .A(y[4276]), .B(x[4276]), .Z(n28111) );
  XNOR U36889 ( .A(y[4277]), .B(x[4277]), .Z(n28110) );
  XOR U36890 ( .A(n28084), .B(n28085), .Z(n28103) );
  XNOR U36891 ( .A(n28100), .B(n28101), .Z(n28085) );
  XNOR U36892 ( .A(n28095), .B(n28096), .Z(n28101) );
  XNOR U36893 ( .A(n28097), .B(n28098), .Z(n28096) );
  XNOR U36894 ( .A(y[4273]), .B(x[4273]), .Z(n28098) );
  XNOR U36895 ( .A(y[4274]), .B(x[4274]), .Z(n28097) );
  XNOR U36896 ( .A(y[4272]), .B(x[4272]), .Z(n28095) );
  XNOR U36897 ( .A(n28089), .B(n28090), .Z(n28100) );
  XNOR U36898 ( .A(y[4269]), .B(x[4269]), .Z(n28090) );
  XNOR U36899 ( .A(n28091), .B(n28092), .Z(n28089) );
  XNOR U36900 ( .A(y[4270]), .B(x[4270]), .Z(n28092) );
  XNOR U36901 ( .A(y[4271]), .B(x[4271]), .Z(n28091) );
  XOR U36902 ( .A(n28083), .B(n28082), .Z(n28084) );
  XNOR U36903 ( .A(n28078), .B(n28079), .Z(n28082) );
  XNOR U36904 ( .A(y[4266]), .B(x[4266]), .Z(n28079) );
  XNOR U36905 ( .A(n28080), .B(n28081), .Z(n28078) );
  XNOR U36906 ( .A(y[4267]), .B(x[4267]), .Z(n28081) );
  XNOR U36907 ( .A(y[4268]), .B(x[4268]), .Z(n28080) );
  XNOR U36908 ( .A(n28072), .B(n28073), .Z(n28083) );
  XNOR U36909 ( .A(y[4263]), .B(x[4263]), .Z(n28073) );
  XNOR U36910 ( .A(n28074), .B(n28075), .Z(n28072) );
  XNOR U36911 ( .A(y[4264]), .B(x[4264]), .Z(n28075) );
  XNOR U36912 ( .A(y[4265]), .B(x[4265]), .Z(n28074) );
  NAND U36913 ( .A(n28139), .B(n28140), .Z(N62897) );
  NANDN U36914 ( .A(n28141), .B(n28142), .Z(n28140) );
  OR U36915 ( .A(n28143), .B(n28144), .Z(n28142) );
  NAND U36916 ( .A(n28143), .B(n28144), .Z(n28139) );
  XOR U36917 ( .A(n28143), .B(n28145), .Z(N62896) );
  XNOR U36918 ( .A(n28141), .B(n28144), .Z(n28145) );
  AND U36919 ( .A(n28146), .B(n28147), .Z(n28144) );
  NANDN U36920 ( .A(n28148), .B(n28149), .Z(n28147) );
  NANDN U36921 ( .A(n28150), .B(n28151), .Z(n28149) );
  NANDN U36922 ( .A(n28151), .B(n28150), .Z(n28146) );
  NAND U36923 ( .A(n28152), .B(n28153), .Z(n28141) );
  NANDN U36924 ( .A(n28154), .B(n28155), .Z(n28153) );
  OR U36925 ( .A(n28156), .B(n28157), .Z(n28155) );
  NAND U36926 ( .A(n28157), .B(n28156), .Z(n28152) );
  AND U36927 ( .A(n28158), .B(n28159), .Z(n28143) );
  NANDN U36928 ( .A(n28160), .B(n28161), .Z(n28159) );
  NANDN U36929 ( .A(n28162), .B(n28163), .Z(n28161) );
  NANDN U36930 ( .A(n28163), .B(n28162), .Z(n28158) );
  XOR U36931 ( .A(n28157), .B(n28164), .Z(N62895) );
  XOR U36932 ( .A(n28154), .B(n28156), .Z(n28164) );
  XNOR U36933 ( .A(n28150), .B(n28165), .Z(n28156) );
  XNOR U36934 ( .A(n28148), .B(n28151), .Z(n28165) );
  NAND U36935 ( .A(n28166), .B(n28167), .Z(n28151) );
  NAND U36936 ( .A(n28168), .B(n28169), .Z(n28167) );
  OR U36937 ( .A(n28170), .B(n28171), .Z(n28168) );
  NANDN U36938 ( .A(n28172), .B(n28170), .Z(n28166) );
  IV U36939 ( .A(n28171), .Z(n28172) );
  NAND U36940 ( .A(n28173), .B(n28174), .Z(n28148) );
  NAND U36941 ( .A(n28175), .B(n28176), .Z(n28174) );
  NANDN U36942 ( .A(n28177), .B(n28178), .Z(n28175) );
  NANDN U36943 ( .A(n28178), .B(n28177), .Z(n28173) );
  AND U36944 ( .A(n28179), .B(n28180), .Z(n28150) );
  NAND U36945 ( .A(n28181), .B(n28182), .Z(n28180) );
  OR U36946 ( .A(n28183), .B(n28184), .Z(n28181) );
  NANDN U36947 ( .A(n28185), .B(n28183), .Z(n28179) );
  NAND U36948 ( .A(n28186), .B(n28187), .Z(n28154) );
  NANDN U36949 ( .A(n28188), .B(n28189), .Z(n28187) );
  OR U36950 ( .A(n28190), .B(n28191), .Z(n28189) );
  NANDN U36951 ( .A(n28192), .B(n28190), .Z(n28186) );
  IV U36952 ( .A(n28191), .Z(n28192) );
  XNOR U36953 ( .A(n28162), .B(n28193), .Z(n28157) );
  XNOR U36954 ( .A(n28160), .B(n28163), .Z(n28193) );
  NAND U36955 ( .A(n28194), .B(n28195), .Z(n28163) );
  NAND U36956 ( .A(n28196), .B(n28197), .Z(n28195) );
  OR U36957 ( .A(n28198), .B(n28199), .Z(n28196) );
  NANDN U36958 ( .A(n28200), .B(n28198), .Z(n28194) );
  IV U36959 ( .A(n28199), .Z(n28200) );
  NAND U36960 ( .A(n28201), .B(n28202), .Z(n28160) );
  NAND U36961 ( .A(n28203), .B(n28204), .Z(n28202) );
  NANDN U36962 ( .A(n28205), .B(n28206), .Z(n28203) );
  NANDN U36963 ( .A(n28206), .B(n28205), .Z(n28201) );
  AND U36964 ( .A(n28207), .B(n28208), .Z(n28162) );
  NAND U36965 ( .A(n28209), .B(n28210), .Z(n28208) );
  OR U36966 ( .A(n28211), .B(n28212), .Z(n28209) );
  NANDN U36967 ( .A(n28213), .B(n28211), .Z(n28207) );
  XNOR U36968 ( .A(n28188), .B(n28214), .Z(N62894) );
  XOR U36969 ( .A(n28190), .B(n28191), .Z(n28214) );
  XNOR U36970 ( .A(n28204), .B(n28215), .Z(n28191) );
  XOR U36971 ( .A(n28205), .B(n28206), .Z(n28215) );
  XOR U36972 ( .A(n28211), .B(n28216), .Z(n28206) );
  XOR U36973 ( .A(n28210), .B(n28213), .Z(n28216) );
  IV U36974 ( .A(n28212), .Z(n28213) );
  NAND U36975 ( .A(n28217), .B(n28218), .Z(n28212) );
  OR U36976 ( .A(n28219), .B(n28220), .Z(n28218) );
  OR U36977 ( .A(n28221), .B(n28222), .Z(n28217) );
  NAND U36978 ( .A(n28223), .B(n28224), .Z(n28210) );
  OR U36979 ( .A(n28225), .B(n28226), .Z(n28224) );
  OR U36980 ( .A(n28227), .B(n28228), .Z(n28223) );
  NOR U36981 ( .A(n28229), .B(n28230), .Z(n28211) );
  ANDN U36982 ( .B(n28231), .A(n28232), .Z(n28205) );
  XNOR U36983 ( .A(n28198), .B(n28233), .Z(n28204) );
  XNOR U36984 ( .A(n28197), .B(n28199), .Z(n28233) );
  NAND U36985 ( .A(n28234), .B(n28235), .Z(n28199) );
  OR U36986 ( .A(n28236), .B(n28237), .Z(n28235) );
  OR U36987 ( .A(n28238), .B(n28239), .Z(n28234) );
  NAND U36988 ( .A(n28240), .B(n28241), .Z(n28197) );
  OR U36989 ( .A(n28242), .B(n28243), .Z(n28241) );
  OR U36990 ( .A(n28244), .B(n28245), .Z(n28240) );
  ANDN U36991 ( .B(n28246), .A(n28247), .Z(n28198) );
  IV U36992 ( .A(n28248), .Z(n28246) );
  ANDN U36993 ( .B(n28249), .A(n28250), .Z(n28190) );
  XOR U36994 ( .A(n28176), .B(n28251), .Z(n28188) );
  XOR U36995 ( .A(n28177), .B(n28178), .Z(n28251) );
  XOR U36996 ( .A(n28183), .B(n28252), .Z(n28178) );
  XOR U36997 ( .A(n28182), .B(n28185), .Z(n28252) );
  IV U36998 ( .A(n28184), .Z(n28185) );
  NAND U36999 ( .A(n28253), .B(n28254), .Z(n28184) );
  OR U37000 ( .A(n28255), .B(n28256), .Z(n28254) );
  OR U37001 ( .A(n28257), .B(n28258), .Z(n28253) );
  NAND U37002 ( .A(n28259), .B(n28260), .Z(n28182) );
  OR U37003 ( .A(n28261), .B(n28262), .Z(n28260) );
  OR U37004 ( .A(n28263), .B(n28264), .Z(n28259) );
  NOR U37005 ( .A(n28265), .B(n28266), .Z(n28183) );
  ANDN U37006 ( .B(n28267), .A(n28268), .Z(n28177) );
  IV U37007 ( .A(n28269), .Z(n28267) );
  XNOR U37008 ( .A(n28170), .B(n28270), .Z(n28176) );
  XNOR U37009 ( .A(n28169), .B(n28171), .Z(n28270) );
  NAND U37010 ( .A(n28271), .B(n28272), .Z(n28171) );
  OR U37011 ( .A(n28273), .B(n28274), .Z(n28272) );
  OR U37012 ( .A(n28275), .B(n28276), .Z(n28271) );
  NAND U37013 ( .A(n28277), .B(n28278), .Z(n28169) );
  OR U37014 ( .A(n28279), .B(n28280), .Z(n28278) );
  OR U37015 ( .A(n28281), .B(n28282), .Z(n28277) );
  ANDN U37016 ( .B(n28283), .A(n28284), .Z(n28170) );
  IV U37017 ( .A(n28285), .Z(n28283) );
  XNOR U37018 ( .A(n28250), .B(n28249), .Z(N62893) );
  XOR U37019 ( .A(n28269), .B(n28268), .Z(n28249) );
  XNOR U37020 ( .A(n28284), .B(n28285), .Z(n28268) );
  XNOR U37021 ( .A(n28279), .B(n28280), .Z(n28285) );
  XNOR U37022 ( .A(n28281), .B(n28282), .Z(n28280) );
  XNOR U37023 ( .A(y[4261]), .B(x[4261]), .Z(n28282) );
  XNOR U37024 ( .A(y[4262]), .B(x[4262]), .Z(n28281) );
  XNOR U37025 ( .A(y[4260]), .B(x[4260]), .Z(n28279) );
  XNOR U37026 ( .A(n28273), .B(n28274), .Z(n28284) );
  XNOR U37027 ( .A(y[4257]), .B(x[4257]), .Z(n28274) );
  XNOR U37028 ( .A(n28275), .B(n28276), .Z(n28273) );
  XNOR U37029 ( .A(y[4258]), .B(x[4258]), .Z(n28276) );
  XNOR U37030 ( .A(y[4259]), .B(x[4259]), .Z(n28275) );
  XNOR U37031 ( .A(n28266), .B(n28265), .Z(n28269) );
  XNOR U37032 ( .A(n28261), .B(n28262), .Z(n28265) );
  XNOR U37033 ( .A(y[4254]), .B(x[4254]), .Z(n28262) );
  XNOR U37034 ( .A(n28263), .B(n28264), .Z(n28261) );
  XNOR U37035 ( .A(y[4255]), .B(x[4255]), .Z(n28264) );
  XNOR U37036 ( .A(y[4256]), .B(x[4256]), .Z(n28263) );
  XNOR U37037 ( .A(n28255), .B(n28256), .Z(n28266) );
  XNOR U37038 ( .A(y[4251]), .B(x[4251]), .Z(n28256) );
  XNOR U37039 ( .A(n28257), .B(n28258), .Z(n28255) );
  XNOR U37040 ( .A(y[4252]), .B(x[4252]), .Z(n28258) );
  XNOR U37041 ( .A(y[4253]), .B(x[4253]), .Z(n28257) );
  XOR U37042 ( .A(n28231), .B(n28232), .Z(n28250) );
  XNOR U37043 ( .A(n28247), .B(n28248), .Z(n28232) );
  XNOR U37044 ( .A(n28242), .B(n28243), .Z(n28248) );
  XNOR U37045 ( .A(n28244), .B(n28245), .Z(n28243) );
  XNOR U37046 ( .A(y[4249]), .B(x[4249]), .Z(n28245) );
  XNOR U37047 ( .A(y[4250]), .B(x[4250]), .Z(n28244) );
  XNOR U37048 ( .A(y[4248]), .B(x[4248]), .Z(n28242) );
  XNOR U37049 ( .A(n28236), .B(n28237), .Z(n28247) );
  XNOR U37050 ( .A(y[4245]), .B(x[4245]), .Z(n28237) );
  XNOR U37051 ( .A(n28238), .B(n28239), .Z(n28236) );
  XNOR U37052 ( .A(y[4246]), .B(x[4246]), .Z(n28239) );
  XNOR U37053 ( .A(y[4247]), .B(x[4247]), .Z(n28238) );
  XOR U37054 ( .A(n28230), .B(n28229), .Z(n28231) );
  XNOR U37055 ( .A(n28225), .B(n28226), .Z(n28229) );
  XNOR U37056 ( .A(y[4242]), .B(x[4242]), .Z(n28226) );
  XNOR U37057 ( .A(n28227), .B(n28228), .Z(n28225) );
  XNOR U37058 ( .A(y[4243]), .B(x[4243]), .Z(n28228) );
  XNOR U37059 ( .A(y[4244]), .B(x[4244]), .Z(n28227) );
  XNOR U37060 ( .A(n28219), .B(n28220), .Z(n28230) );
  XNOR U37061 ( .A(y[4239]), .B(x[4239]), .Z(n28220) );
  XNOR U37062 ( .A(n28221), .B(n28222), .Z(n28219) );
  XNOR U37063 ( .A(y[4240]), .B(x[4240]), .Z(n28222) );
  XNOR U37064 ( .A(y[4241]), .B(x[4241]), .Z(n28221) );
  NAND U37065 ( .A(n28286), .B(n28287), .Z(N62884) );
  NANDN U37066 ( .A(n28288), .B(n28289), .Z(n28287) );
  OR U37067 ( .A(n28290), .B(n28291), .Z(n28289) );
  NAND U37068 ( .A(n28290), .B(n28291), .Z(n28286) );
  XOR U37069 ( .A(n28290), .B(n28292), .Z(N62883) );
  XNOR U37070 ( .A(n28288), .B(n28291), .Z(n28292) );
  AND U37071 ( .A(n28293), .B(n28294), .Z(n28291) );
  NANDN U37072 ( .A(n28295), .B(n28296), .Z(n28294) );
  NANDN U37073 ( .A(n28297), .B(n28298), .Z(n28296) );
  NANDN U37074 ( .A(n28298), .B(n28297), .Z(n28293) );
  NAND U37075 ( .A(n28299), .B(n28300), .Z(n28288) );
  NANDN U37076 ( .A(n28301), .B(n28302), .Z(n28300) );
  OR U37077 ( .A(n28303), .B(n28304), .Z(n28302) );
  NAND U37078 ( .A(n28304), .B(n28303), .Z(n28299) );
  AND U37079 ( .A(n28305), .B(n28306), .Z(n28290) );
  NANDN U37080 ( .A(n28307), .B(n28308), .Z(n28306) );
  NANDN U37081 ( .A(n28309), .B(n28310), .Z(n28308) );
  NANDN U37082 ( .A(n28310), .B(n28309), .Z(n28305) );
  XOR U37083 ( .A(n28304), .B(n28311), .Z(N62882) );
  XOR U37084 ( .A(n28301), .B(n28303), .Z(n28311) );
  XNOR U37085 ( .A(n28297), .B(n28312), .Z(n28303) );
  XNOR U37086 ( .A(n28295), .B(n28298), .Z(n28312) );
  NAND U37087 ( .A(n28313), .B(n28314), .Z(n28298) );
  NAND U37088 ( .A(n28315), .B(n28316), .Z(n28314) );
  OR U37089 ( .A(n28317), .B(n28318), .Z(n28315) );
  NANDN U37090 ( .A(n28319), .B(n28317), .Z(n28313) );
  IV U37091 ( .A(n28318), .Z(n28319) );
  NAND U37092 ( .A(n28320), .B(n28321), .Z(n28295) );
  NAND U37093 ( .A(n28322), .B(n28323), .Z(n28321) );
  NANDN U37094 ( .A(n28324), .B(n28325), .Z(n28322) );
  NANDN U37095 ( .A(n28325), .B(n28324), .Z(n28320) );
  AND U37096 ( .A(n28326), .B(n28327), .Z(n28297) );
  NAND U37097 ( .A(n28328), .B(n28329), .Z(n28327) );
  OR U37098 ( .A(n28330), .B(n28331), .Z(n28328) );
  NANDN U37099 ( .A(n28332), .B(n28330), .Z(n28326) );
  NAND U37100 ( .A(n28333), .B(n28334), .Z(n28301) );
  NANDN U37101 ( .A(n28335), .B(n28336), .Z(n28334) );
  OR U37102 ( .A(n28337), .B(n28338), .Z(n28336) );
  NANDN U37103 ( .A(n28339), .B(n28337), .Z(n28333) );
  IV U37104 ( .A(n28338), .Z(n28339) );
  XNOR U37105 ( .A(n28309), .B(n28340), .Z(n28304) );
  XNOR U37106 ( .A(n28307), .B(n28310), .Z(n28340) );
  NAND U37107 ( .A(n28341), .B(n28342), .Z(n28310) );
  NAND U37108 ( .A(n28343), .B(n28344), .Z(n28342) );
  OR U37109 ( .A(n28345), .B(n28346), .Z(n28343) );
  NANDN U37110 ( .A(n28347), .B(n28345), .Z(n28341) );
  IV U37111 ( .A(n28346), .Z(n28347) );
  NAND U37112 ( .A(n28348), .B(n28349), .Z(n28307) );
  NAND U37113 ( .A(n28350), .B(n28351), .Z(n28349) );
  NANDN U37114 ( .A(n28352), .B(n28353), .Z(n28350) );
  NANDN U37115 ( .A(n28353), .B(n28352), .Z(n28348) );
  AND U37116 ( .A(n28354), .B(n28355), .Z(n28309) );
  NAND U37117 ( .A(n28356), .B(n28357), .Z(n28355) );
  OR U37118 ( .A(n28358), .B(n28359), .Z(n28356) );
  NANDN U37119 ( .A(n28360), .B(n28358), .Z(n28354) );
  XNOR U37120 ( .A(n28335), .B(n28361), .Z(N62881) );
  XOR U37121 ( .A(n28337), .B(n28338), .Z(n28361) );
  XNOR U37122 ( .A(n28351), .B(n28362), .Z(n28338) );
  XOR U37123 ( .A(n28352), .B(n28353), .Z(n28362) );
  XOR U37124 ( .A(n28358), .B(n28363), .Z(n28353) );
  XOR U37125 ( .A(n28357), .B(n28360), .Z(n28363) );
  IV U37126 ( .A(n28359), .Z(n28360) );
  NAND U37127 ( .A(n28364), .B(n28365), .Z(n28359) );
  OR U37128 ( .A(n28366), .B(n28367), .Z(n28365) );
  OR U37129 ( .A(n28368), .B(n28369), .Z(n28364) );
  NAND U37130 ( .A(n28370), .B(n28371), .Z(n28357) );
  OR U37131 ( .A(n28372), .B(n28373), .Z(n28371) );
  OR U37132 ( .A(n28374), .B(n28375), .Z(n28370) );
  NOR U37133 ( .A(n28376), .B(n28377), .Z(n28358) );
  ANDN U37134 ( .B(n28378), .A(n28379), .Z(n28352) );
  XNOR U37135 ( .A(n28345), .B(n28380), .Z(n28351) );
  XNOR U37136 ( .A(n28344), .B(n28346), .Z(n28380) );
  NAND U37137 ( .A(n28381), .B(n28382), .Z(n28346) );
  OR U37138 ( .A(n28383), .B(n28384), .Z(n28382) );
  OR U37139 ( .A(n28385), .B(n28386), .Z(n28381) );
  NAND U37140 ( .A(n28387), .B(n28388), .Z(n28344) );
  OR U37141 ( .A(n28389), .B(n28390), .Z(n28388) );
  OR U37142 ( .A(n28391), .B(n28392), .Z(n28387) );
  ANDN U37143 ( .B(n28393), .A(n28394), .Z(n28345) );
  IV U37144 ( .A(n28395), .Z(n28393) );
  ANDN U37145 ( .B(n28396), .A(n28397), .Z(n28337) );
  XOR U37146 ( .A(n28323), .B(n28398), .Z(n28335) );
  XOR U37147 ( .A(n28324), .B(n28325), .Z(n28398) );
  XOR U37148 ( .A(n28330), .B(n28399), .Z(n28325) );
  XOR U37149 ( .A(n28329), .B(n28332), .Z(n28399) );
  IV U37150 ( .A(n28331), .Z(n28332) );
  NAND U37151 ( .A(n28400), .B(n28401), .Z(n28331) );
  OR U37152 ( .A(n28402), .B(n28403), .Z(n28401) );
  OR U37153 ( .A(n28404), .B(n28405), .Z(n28400) );
  NAND U37154 ( .A(n28406), .B(n28407), .Z(n28329) );
  OR U37155 ( .A(n28408), .B(n28409), .Z(n28407) );
  OR U37156 ( .A(n28410), .B(n28411), .Z(n28406) );
  NOR U37157 ( .A(n28412), .B(n28413), .Z(n28330) );
  ANDN U37158 ( .B(n28414), .A(n28415), .Z(n28324) );
  IV U37159 ( .A(n28416), .Z(n28414) );
  XNOR U37160 ( .A(n28317), .B(n28417), .Z(n28323) );
  XNOR U37161 ( .A(n28316), .B(n28318), .Z(n28417) );
  NAND U37162 ( .A(n28418), .B(n28419), .Z(n28318) );
  OR U37163 ( .A(n28420), .B(n28421), .Z(n28419) );
  OR U37164 ( .A(n28422), .B(n28423), .Z(n28418) );
  NAND U37165 ( .A(n28424), .B(n28425), .Z(n28316) );
  OR U37166 ( .A(n28426), .B(n28427), .Z(n28425) );
  OR U37167 ( .A(n28428), .B(n28429), .Z(n28424) );
  ANDN U37168 ( .B(n28430), .A(n28431), .Z(n28317) );
  IV U37169 ( .A(n28432), .Z(n28430) );
  XNOR U37170 ( .A(n28397), .B(n28396), .Z(N62880) );
  XOR U37171 ( .A(n28416), .B(n28415), .Z(n28396) );
  XNOR U37172 ( .A(n28431), .B(n28432), .Z(n28415) );
  XNOR U37173 ( .A(n28426), .B(n28427), .Z(n28432) );
  XNOR U37174 ( .A(n28428), .B(n28429), .Z(n28427) );
  XNOR U37175 ( .A(y[4237]), .B(x[4237]), .Z(n28429) );
  XNOR U37176 ( .A(y[4238]), .B(x[4238]), .Z(n28428) );
  XNOR U37177 ( .A(y[4236]), .B(x[4236]), .Z(n28426) );
  XNOR U37178 ( .A(n28420), .B(n28421), .Z(n28431) );
  XNOR U37179 ( .A(y[4233]), .B(x[4233]), .Z(n28421) );
  XNOR U37180 ( .A(n28422), .B(n28423), .Z(n28420) );
  XNOR U37181 ( .A(y[4234]), .B(x[4234]), .Z(n28423) );
  XNOR U37182 ( .A(y[4235]), .B(x[4235]), .Z(n28422) );
  XNOR U37183 ( .A(n28413), .B(n28412), .Z(n28416) );
  XNOR U37184 ( .A(n28408), .B(n28409), .Z(n28412) );
  XNOR U37185 ( .A(y[4230]), .B(x[4230]), .Z(n28409) );
  XNOR U37186 ( .A(n28410), .B(n28411), .Z(n28408) );
  XNOR U37187 ( .A(y[4231]), .B(x[4231]), .Z(n28411) );
  XNOR U37188 ( .A(y[4232]), .B(x[4232]), .Z(n28410) );
  XNOR U37189 ( .A(n28402), .B(n28403), .Z(n28413) );
  XNOR U37190 ( .A(y[4227]), .B(x[4227]), .Z(n28403) );
  XNOR U37191 ( .A(n28404), .B(n28405), .Z(n28402) );
  XNOR U37192 ( .A(y[4228]), .B(x[4228]), .Z(n28405) );
  XNOR U37193 ( .A(y[4229]), .B(x[4229]), .Z(n28404) );
  XOR U37194 ( .A(n28378), .B(n28379), .Z(n28397) );
  XNOR U37195 ( .A(n28394), .B(n28395), .Z(n28379) );
  XNOR U37196 ( .A(n28389), .B(n28390), .Z(n28395) );
  XNOR U37197 ( .A(n28391), .B(n28392), .Z(n28390) );
  XNOR U37198 ( .A(y[4225]), .B(x[4225]), .Z(n28392) );
  XNOR U37199 ( .A(y[4226]), .B(x[4226]), .Z(n28391) );
  XNOR U37200 ( .A(y[4224]), .B(x[4224]), .Z(n28389) );
  XNOR U37201 ( .A(n28383), .B(n28384), .Z(n28394) );
  XNOR U37202 ( .A(y[4221]), .B(x[4221]), .Z(n28384) );
  XNOR U37203 ( .A(n28385), .B(n28386), .Z(n28383) );
  XNOR U37204 ( .A(y[4222]), .B(x[4222]), .Z(n28386) );
  XNOR U37205 ( .A(y[4223]), .B(x[4223]), .Z(n28385) );
  XOR U37206 ( .A(n28377), .B(n28376), .Z(n28378) );
  XNOR U37207 ( .A(n28372), .B(n28373), .Z(n28376) );
  XNOR U37208 ( .A(y[4218]), .B(x[4218]), .Z(n28373) );
  XNOR U37209 ( .A(n28374), .B(n28375), .Z(n28372) );
  XNOR U37210 ( .A(y[4219]), .B(x[4219]), .Z(n28375) );
  XNOR U37211 ( .A(y[4220]), .B(x[4220]), .Z(n28374) );
  XNOR U37212 ( .A(n28366), .B(n28367), .Z(n28377) );
  XNOR U37213 ( .A(y[4215]), .B(x[4215]), .Z(n28367) );
  XNOR U37214 ( .A(n28368), .B(n28369), .Z(n28366) );
  XNOR U37215 ( .A(y[4216]), .B(x[4216]), .Z(n28369) );
  XNOR U37216 ( .A(y[4217]), .B(x[4217]), .Z(n28368) );
  NAND U37217 ( .A(n28433), .B(n28434), .Z(N62871) );
  NANDN U37218 ( .A(n28435), .B(n28436), .Z(n28434) );
  OR U37219 ( .A(n28437), .B(n28438), .Z(n28436) );
  NAND U37220 ( .A(n28437), .B(n28438), .Z(n28433) );
  XOR U37221 ( .A(n28437), .B(n28439), .Z(N62870) );
  XNOR U37222 ( .A(n28435), .B(n28438), .Z(n28439) );
  AND U37223 ( .A(n28440), .B(n28441), .Z(n28438) );
  NANDN U37224 ( .A(n28442), .B(n28443), .Z(n28441) );
  NANDN U37225 ( .A(n28444), .B(n28445), .Z(n28443) );
  NANDN U37226 ( .A(n28445), .B(n28444), .Z(n28440) );
  NAND U37227 ( .A(n28446), .B(n28447), .Z(n28435) );
  NANDN U37228 ( .A(n28448), .B(n28449), .Z(n28447) );
  OR U37229 ( .A(n28450), .B(n28451), .Z(n28449) );
  NAND U37230 ( .A(n28451), .B(n28450), .Z(n28446) );
  AND U37231 ( .A(n28452), .B(n28453), .Z(n28437) );
  NANDN U37232 ( .A(n28454), .B(n28455), .Z(n28453) );
  NANDN U37233 ( .A(n28456), .B(n28457), .Z(n28455) );
  NANDN U37234 ( .A(n28457), .B(n28456), .Z(n28452) );
  XOR U37235 ( .A(n28451), .B(n28458), .Z(N62869) );
  XOR U37236 ( .A(n28448), .B(n28450), .Z(n28458) );
  XNOR U37237 ( .A(n28444), .B(n28459), .Z(n28450) );
  XNOR U37238 ( .A(n28442), .B(n28445), .Z(n28459) );
  NAND U37239 ( .A(n28460), .B(n28461), .Z(n28445) );
  NAND U37240 ( .A(n28462), .B(n28463), .Z(n28461) );
  OR U37241 ( .A(n28464), .B(n28465), .Z(n28462) );
  NANDN U37242 ( .A(n28466), .B(n28464), .Z(n28460) );
  IV U37243 ( .A(n28465), .Z(n28466) );
  NAND U37244 ( .A(n28467), .B(n28468), .Z(n28442) );
  NAND U37245 ( .A(n28469), .B(n28470), .Z(n28468) );
  NANDN U37246 ( .A(n28471), .B(n28472), .Z(n28469) );
  NANDN U37247 ( .A(n28472), .B(n28471), .Z(n28467) );
  AND U37248 ( .A(n28473), .B(n28474), .Z(n28444) );
  NAND U37249 ( .A(n28475), .B(n28476), .Z(n28474) );
  OR U37250 ( .A(n28477), .B(n28478), .Z(n28475) );
  NANDN U37251 ( .A(n28479), .B(n28477), .Z(n28473) );
  NAND U37252 ( .A(n28480), .B(n28481), .Z(n28448) );
  NANDN U37253 ( .A(n28482), .B(n28483), .Z(n28481) );
  OR U37254 ( .A(n28484), .B(n28485), .Z(n28483) );
  NANDN U37255 ( .A(n28486), .B(n28484), .Z(n28480) );
  IV U37256 ( .A(n28485), .Z(n28486) );
  XNOR U37257 ( .A(n28456), .B(n28487), .Z(n28451) );
  XNOR U37258 ( .A(n28454), .B(n28457), .Z(n28487) );
  NAND U37259 ( .A(n28488), .B(n28489), .Z(n28457) );
  NAND U37260 ( .A(n28490), .B(n28491), .Z(n28489) );
  OR U37261 ( .A(n28492), .B(n28493), .Z(n28490) );
  NANDN U37262 ( .A(n28494), .B(n28492), .Z(n28488) );
  IV U37263 ( .A(n28493), .Z(n28494) );
  NAND U37264 ( .A(n28495), .B(n28496), .Z(n28454) );
  NAND U37265 ( .A(n28497), .B(n28498), .Z(n28496) );
  NANDN U37266 ( .A(n28499), .B(n28500), .Z(n28497) );
  NANDN U37267 ( .A(n28500), .B(n28499), .Z(n28495) );
  AND U37268 ( .A(n28501), .B(n28502), .Z(n28456) );
  NAND U37269 ( .A(n28503), .B(n28504), .Z(n28502) );
  OR U37270 ( .A(n28505), .B(n28506), .Z(n28503) );
  NANDN U37271 ( .A(n28507), .B(n28505), .Z(n28501) );
  XNOR U37272 ( .A(n28482), .B(n28508), .Z(N62868) );
  XOR U37273 ( .A(n28484), .B(n28485), .Z(n28508) );
  XNOR U37274 ( .A(n28498), .B(n28509), .Z(n28485) );
  XOR U37275 ( .A(n28499), .B(n28500), .Z(n28509) );
  XOR U37276 ( .A(n28505), .B(n28510), .Z(n28500) );
  XOR U37277 ( .A(n28504), .B(n28507), .Z(n28510) );
  IV U37278 ( .A(n28506), .Z(n28507) );
  NAND U37279 ( .A(n28511), .B(n28512), .Z(n28506) );
  OR U37280 ( .A(n28513), .B(n28514), .Z(n28512) );
  OR U37281 ( .A(n28515), .B(n28516), .Z(n28511) );
  NAND U37282 ( .A(n28517), .B(n28518), .Z(n28504) );
  OR U37283 ( .A(n28519), .B(n28520), .Z(n28518) );
  OR U37284 ( .A(n28521), .B(n28522), .Z(n28517) );
  NOR U37285 ( .A(n28523), .B(n28524), .Z(n28505) );
  ANDN U37286 ( .B(n28525), .A(n28526), .Z(n28499) );
  XNOR U37287 ( .A(n28492), .B(n28527), .Z(n28498) );
  XNOR U37288 ( .A(n28491), .B(n28493), .Z(n28527) );
  NAND U37289 ( .A(n28528), .B(n28529), .Z(n28493) );
  OR U37290 ( .A(n28530), .B(n28531), .Z(n28529) );
  OR U37291 ( .A(n28532), .B(n28533), .Z(n28528) );
  NAND U37292 ( .A(n28534), .B(n28535), .Z(n28491) );
  OR U37293 ( .A(n28536), .B(n28537), .Z(n28535) );
  OR U37294 ( .A(n28538), .B(n28539), .Z(n28534) );
  ANDN U37295 ( .B(n28540), .A(n28541), .Z(n28492) );
  IV U37296 ( .A(n28542), .Z(n28540) );
  ANDN U37297 ( .B(n28543), .A(n28544), .Z(n28484) );
  XOR U37298 ( .A(n28470), .B(n28545), .Z(n28482) );
  XOR U37299 ( .A(n28471), .B(n28472), .Z(n28545) );
  XOR U37300 ( .A(n28477), .B(n28546), .Z(n28472) );
  XOR U37301 ( .A(n28476), .B(n28479), .Z(n28546) );
  IV U37302 ( .A(n28478), .Z(n28479) );
  NAND U37303 ( .A(n28547), .B(n28548), .Z(n28478) );
  OR U37304 ( .A(n28549), .B(n28550), .Z(n28548) );
  OR U37305 ( .A(n28551), .B(n28552), .Z(n28547) );
  NAND U37306 ( .A(n28553), .B(n28554), .Z(n28476) );
  OR U37307 ( .A(n28555), .B(n28556), .Z(n28554) );
  OR U37308 ( .A(n28557), .B(n28558), .Z(n28553) );
  NOR U37309 ( .A(n28559), .B(n28560), .Z(n28477) );
  ANDN U37310 ( .B(n28561), .A(n28562), .Z(n28471) );
  IV U37311 ( .A(n28563), .Z(n28561) );
  XNOR U37312 ( .A(n28464), .B(n28564), .Z(n28470) );
  XNOR U37313 ( .A(n28463), .B(n28465), .Z(n28564) );
  NAND U37314 ( .A(n28565), .B(n28566), .Z(n28465) );
  OR U37315 ( .A(n28567), .B(n28568), .Z(n28566) );
  OR U37316 ( .A(n28569), .B(n28570), .Z(n28565) );
  NAND U37317 ( .A(n28571), .B(n28572), .Z(n28463) );
  OR U37318 ( .A(n28573), .B(n28574), .Z(n28572) );
  OR U37319 ( .A(n28575), .B(n28576), .Z(n28571) );
  ANDN U37320 ( .B(n28577), .A(n28578), .Z(n28464) );
  IV U37321 ( .A(n28579), .Z(n28577) );
  XNOR U37322 ( .A(n28544), .B(n28543), .Z(N62867) );
  XOR U37323 ( .A(n28563), .B(n28562), .Z(n28543) );
  XNOR U37324 ( .A(n28578), .B(n28579), .Z(n28562) );
  XNOR U37325 ( .A(n28573), .B(n28574), .Z(n28579) );
  XNOR U37326 ( .A(n28575), .B(n28576), .Z(n28574) );
  XNOR U37327 ( .A(y[4213]), .B(x[4213]), .Z(n28576) );
  XNOR U37328 ( .A(y[4214]), .B(x[4214]), .Z(n28575) );
  XNOR U37329 ( .A(y[4212]), .B(x[4212]), .Z(n28573) );
  XNOR U37330 ( .A(n28567), .B(n28568), .Z(n28578) );
  XNOR U37331 ( .A(y[4209]), .B(x[4209]), .Z(n28568) );
  XNOR U37332 ( .A(n28569), .B(n28570), .Z(n28567) );
  XNOR U37333 ( .A(y[4210]), .B(x[4210]), .Z(n28570) );
  XNOR U37334 ( .A(y[4211]), .B(x[4211]), .Z(n28569) );
  XNOR U37335 ( .A(n28560), .B(n28559), .Z(n28563) );
  XNOR U37336 ( .A(n28555), .B(n28556), .Z(n28559) );
  XNOR U37337 ( .A(y[4206]), .B(x[4206]), .Z(n28556) );
  XNOR U37338 ( .A(n28557), .B(n28558), .Z(n28555) );
  XNOR U37339 ( .A(y[4207]), .B(x[4207]), .Z(n28558) );
  XNOR U37340 ( .A(y[4208]), .B(x[4208]), .Z(n28557) );
  XNOR U37341 ( .A(n28549), .B(n28550), .Z(n28560) );
  XNOR U37342 ( .A(y[4203]), .B(x[4203]), .Z(n28550) );
  XNOR U37343 ( .A(n28551), .B(n28552), .Z(n28549) );
  XNOR U37344 ( .A(y[4204]), .B(x[4204]), .Z(n28552) );
  XNOR U37345 ( .A(y[4205]), .B(x[4205]), .Z(n28551) );
  XOR U37346 ( .A(n28525), .B(n28526), .Z(n28544) );
  XNOR U37347 ( .A(n28541), .B(n28542), .Z(n28526) );
  XNOR U37348 ( .A(n28536), .B(n28537), .Z(n28542) );
  XNOR U37349 ( .A(n28538), .B(n28539), .Z(n28537) );
  XNOR U37350 ( .A(y[4201]), .B(x[4201]), .Z(n28539) );
  XNOR U37351 ( .A(y[4202]), .B(x[4202]), .Z(n28538) );
  XNOR U37352 ( .A(y[4200]), .B(x[4200]), .Z(n28536) );
  XNOR U37353 ( .A(n28530), .B(n28531), .Z(n28541) );
  XNOR U37354 ( .A(y[4197]), .B(x[4197]), .Z(n28531) );
  XNOR U37355 ( .A(n28532), .B(n28533), .Z(n28530) );
  XNOR U37356 ( .A(y[4198]), .B(x[4198]), .Z(n28533) );
  XNOR U37357 ( .A(y[4199]), .B(x[4199]), .Z(n28532) );
  XOR U37358 ( .A(n28524), .B(n28523), .Z(n28525) );
  XNOR U37359 ( .A(n28519), .B(n28520), .Z(n28523) );
  XNOR U37360 ( .A(y[4194]), .B(x[4194]), .Z(n28520) );
  XNOR U37361 ( .A(n28521), .B(n28522), .Z(n28519) );
  XNOR U37362 ( .A(y[4195]), .B(x[4195]), .Z(n28522) );
  XNOR U37363 ( .A(y[4196]), .B(x[4196]), .Z(n28521) );
  XNOR U37364 ( .A(n28513), .B(n28514), .Z(n28524) );
  XNOR U37365 ( .A(y[4191]), .B(x[4191]), .Z(n28514) );
  XNOR U37366 ( .A(n28515), .B(n28516), .Z(n28513) );
  XNOR U37367 ( .A(y[4192]), .B(x[4192]), .Z(n28516) );
  XNOR U37368 ( .A(y[4193]), .B(x[4193]), .Z(n28515) );
  NAND U37369 ( .A(n28580), .B(n28581), .Z(N62858) );
  NANDN U37370 ( .A(n28582), .B(n28583), .Z(n28581) );
  OR U37371 ( .A(n28584), .B(n28585), .Z(n28583) );
  NAND U37372 ( .A(n28584), .B(n28585), .Z(n28580) );
  XOR U37373 ( .A(n28584), .B(n28586), .Z(N62857) );
  XNOR U37374 ( .A(n28582), .B(n28585), .Z(n28586) );
  AND U37375 ( .A(n28587), .B(n28588), .Z(n28585) );
  NANDN U37376 ( .A(n28589), .B(n28590), .Z(n28588) );
  NANDN U37377 ( .A(n28591), .B(n28592), .Z(n28590) );
  NANDN U37378 ( .A(n28592), .B(n28591), .Z(n28587) );
  NAND U37379 ( .A(n28593), .B(n28594), .Z(n28582) );
  NANDN U37380 ( .A(n28595), .B(n28596), .Z(n28594) );
  OR U37381 ( .A(n28597), .B(n28598), .Z(n28596) );
  NAND U37382 ( .A(n28598), .B(n28597), .Z(n28593) );
  AND U37383 ( .A(n28599), .B(n28600), .Z(n28584) );
  NANDN U37384 ( .A(n28601), .B(n28602), .Z(n28600) );
  NANDN U37385 ( .A(n28603), .B(n28604), .Z(n28602) );
  NANDN U37386 ( .A(n28604), .B(n28603), .Z(n28599) );
  XOR U37387 ( .A(n28598), .B(n28605), .Z(N62856) );
  XOR U37388 ( .A(n28595), .B(n28597), .Z(n28605) );
  XNOR U37389 ( .A(n28591), .B(n28606), .Z(n28597) );
  XNOR U37390 ( .A(n28589), .B(n28592), .Z(n28606) );
  NAND U37391 ( .A(n28607), .B(n28608), .Z(n28592) );
  NAND U37392 ( .A(n28609), .B(n28610), .Z(n28608) );
  OR U37393 ( .A(n28611), .B(n28612), .Z(n28609) );
  NANDN U37394 ( .A(n28613), .B(n28611), .Z(n28607) );
  IV U37395 ( .A(n28612), .Z(n28613) );
  NAND U37396 ( .A(n28614), .B(n28615), .Z(n28589) );
  NAND U37397 ( .A(n28616), .B(n28617), .Z(n28615) );
  NANDN U37398 ( .A(n28618), .B(n28619), .Z(n28616) );
  NANDN U37399 ( .A(n28619), .B(n28618), .Z(n28614) );
  AND U37400 ( .A(n28620), .B(n28621), .Z(n28591) );
  NAND U37401 ( .A(n28622), .B(n28623), .Z(n28621) );
  OR U37402 ( .A(n28624), .B(n28625), .Z(n28622) );
  NANDN U37403 ( .A(n28626), .B(n28624), .Z(n28620) );
  NAND U37404 ( .A(n28627), .B(n28628), .Z(n28595) );
  NANDN U37405 ( .A(n28629), .B(n28630), .Z(n28628) );
  OR U37406 ( .A(n28631), .B(n28632), .Z(n28630) );
  NANDN U37407 ( .A(n28633), .B(n28631), .Z(n28627) );
  IV U37408 ( .A(n28632), .Z(n28633) );
  XNOR U37409 ( .A(n28603), .B(n28634), .Z(n28598) );
  XNOR U37410 ( .A(n28601), .B(n28604), .Z(n28634) );
  NAND U37411 ( .A(n28635), .B(n28636), .Z(n28604) );
  NAND U37412 ( .A(n28637), .B(n28638), .Z(n28636) );
  OR U37413 ( .A(n28639), .B(n28640), .Z(n28637) );
  NANDN U37414 ( .A(n28641), .B(n28639), .Z(n28635) );
  IV U37415 ( .A(n28640), .Z(n28641) );
  NAND U37416 ( .A(n28642), .B(n28643), .Z(n28601) );
  NAND U37417 ( .A(n28644), .B(n28645), .Z(n28643) );
  NANDN U37418 ( .A(n28646), .B(n28647), .Z(n28644) );
  NANDN U37419 ( .A(n28647), .B(n28646), .Z(n28642) );
  AND U37420 ( .A(n28648), .B(n28649), .Z(n28603) );
  NAND U37421 ( .A(n28650), .B(n28651), .Z(n28649) );
  OR U37422 ( .A(n28652), .B(n28653), .Z(n28650) );
  NANDN U37423 ( .A(n28654), .B(n28652), .Z(n28648) );
  XNOR U37424 ( .A(n28629), .B(n28655), .Z(N62855) );
  XOR U37425 ( .A(n28631), .B(n28632), .Z(n28655) );
  XNOR U37426 ( .A(n28645), .B(n28656), .Z(n28632) );
  XOR U37427 ( .A(n28646), .B(n28647), .Z(n28656) );
  XOR U37428 ( .A(n28652), .B(n28657), .Z(n28647) );
  XOR U37429 ( .A(n28651), .B(n28654), .Z(n28657) );
  IV U37430 ( .A(n28653), .Z(n28654) );
  NAND U37431 ( .A(n28658), .B(n28659), .Z(n28653) );
  OR U37432 ( .A(n28660), .B(n28661), .Z(n28659) );
  OR U37433 ( .A(n28662), .B(n28663), .Z(n28658) );
  NAND U37434 ( .A(n28664), .B(n28665), .Z(n28651) );
  OR U37435 ( .A(n28666), .B(n28667), .Z(n28665) );
  OR U37436 ( .A(n28668), .B(n28669), .Z(n28664) );
  NOR U37437 ( .A(n28670), .B(n28671), .Z(n28652) );
  ANDN U37438 ( .B(n28672), .A(n28673), .Z(n28646) );
  XNOR U37439 ( .A(n28639), .B(n28674), .Z(n28645) );
  XNOR U37440 ( .A(n28638), .B(n28640), .Z(n28674) );
  NAND U37441 ( .A(n28675), .B(n28676), .Z(n28640) );
  OR U37442 ( .A(n28677), .B(n28678), .Z(n28676) );
  OR U37443 ( .A(n28679), .B(n28680), .Z(n28675) );
  NAND U37444 ( .A(n28681), .B(n28682), .Z(n28638) );
  OR U37445 ( .A(n28683), .B(n28684), .Z(n28682) );
  OR U37446 ( .A(n28685), .B(n28686), .Z(n28681) );
  ANDN U37447 ( .B(n28687), .A(n28688), .Z(n28639) );
  IV U37448 ( .A(n28689), .Z(n28687) );
  ANDN U37449 ( .B(n28690), .A(n28691), .Z(n28631) );
  XOR U37450 ( .A(n28617), .B(n28692), .Z(n28629) );
  XOR U37451 ( .A(n28618), .B(n28619), .Z(n28692) );
  XOR U37452 ( .A(n28624), .B(n28693), .Z(n28619) );
  XOR U37453 ( .A(n28623), .B(n28626), .Z(n28693) );
  IV U37454 ( .A(n28625), .Z(n28626) );
  NAND U37455 ( .A(n28694), .B(n28695), .Z(n28625) );
  OR U37456 ( .A(n28696), .B(n28697), .Z(n28695) );
  OR U37457 ( .A(n28698), .B(n28699), .Z(n28694) );
  NAND U37458 ( .A(n28700), .B(n28701), .Z(n28623) );
  OR U37459 ( .A(n28702), .B(n28703), .Z(n28701) );
  OR U37460 ( .A(n28704), .B(n28705), .Z(n28700) );
  NOR U37461 ( .A(n28706), .B(n28707), .Z(n28624) );
  ANDN U37462 ( .B(n28708), .A(n28709), .Z(n28618) );
  IV U37463 ( .A(n28710), .Z(n28708) );
  XNOR U37464 ( .A(n28611), .B(n28711), .Z(n28617) );
  XNOR U37465 ( .A(n28610), .B(n28612), .Z(n28711) );
  NAND U37466 ( .A(n28712), .B(n28713), .Z(n28612) );
  OR U37467 ( .A(n28714), .B(n28715), .Z(n28713) );
  OR U37468 ( .A(n28716), .B(n28717), .Z(n28712) );
  NAND U37469 ( .A(n28718), .B(n28719), .Z(n28610) );
  OR U37470 ( .A(n28720), .B(n28721), .Z(n28719) );
  OR U37471 ( .A(n28722), .B(n28723), .Z(n28718) );
  ANDN U37472 ( .B(n28724), .A(n28725), .Z(n28611) );
  IV U37473 ( .A(n28726), .Z(n28724) );
  XNOR U37474 ( .A(n28691), .B(n28690), .Z(N62854) );
  XOR U37475 ( .A(n28710), .B(n28709), .Z(n28690) );
  XNOR U37476 ( .A(n28725), .B(n28726), .Z(n28709) );
  XNOR U37477 ( .A(n28720), .B(n28721), .Z(n28726) );
  XNOR U37478 ( .A(n28722), .B(n28723), .Z(n28721) );
  XNOR U37479 ( .A(y[4189]), .B(x[4189]), .Z(n28723) );
  XNOR U37480 ( .A(y[4190]), .B(x[4190]), .Z(n28722) );
  XNOR U37481 ( .A(y[4188]), .B(x[4188]), .Z(n28720) );
  XNOR U37482 ( .A(n28714), .B(n28715), .Z(n28725) );
  XNOR U37483 ( .A(y[4185]), .B(x[4185]), .Z(n28715) );
  XNOR U37484 ( .A(n28716), .B(n28717), .Z(n28714) );
  XNOR U37485 ( .A(y[4186]), .B(x[4186]), .Z(n28717) );
  XNOR U37486 ( .A(y[4187]), .B(x[4187]), .Z(n28716) );
  XNOR U37487 ( .A(n28707), .B(n28706), .Z(n28710) );
  XNOR U37488 ( .A(n28702), .B(n28703), .Z(n28706) );
  XNOR U37489 ( .A(y[4182]), .B(x[4182]), .Z(n28703) );
  XNOR U37490 ( .A(n28704), .B(n28705), .Z(n28702) );
  XNOR U37491 ( .A(y[4183]), .B(x[4183]), .Z(n28705) );
  XNOR U37492 ( .A(y[4184]), .B(x[4184]), .Z(n28704) );
  XNOR U37493 ( .A(n28696), .B(n28697), .Z(n28707) );
  XNOR U37494 ( .A(y[4179]), .B(x[4179]), .Z(n28697) );
  XNOR U37495 ( .A(n28698), .B(n28699), .Z(n28696) );
  XNOR U37496 ( .A(y[4180]), .B(x[4180]), .Z(n28699) );
  XNOR U37497 ( .A(y[4181]), .B(x[4181]), .Z(n28698) );
  XOR U37498 ( .A(n28672), .B(n28673), .Z(n28691) );
  XNOR U37499 ( .A(n28688), .B(n28689), .Z(n28673) );
  XNOR U37500 ( .A(n28683), .B(n28684), .Z(n28689) );
  XNOR U37501 ( .A(n28685), .B(n28686), .Z(n28684) );
  XNOR U37502 ( .A(y[4177]), .B(x[4177]), .Z(n28686) );
  XNOR U37503 ( .A(y[4178]), .B(x[4178]), .Z(n28685) );
  XNOR U37504 ( .A(y[4176]), .B(x[4176]), .Z(n28683) );
  XNOR U37505 ( .A(n28677), .B(n28678), .Z(n28688) );
  XNOR U37506 ( .A(y[4173]), .B(x[4173]), .Z(n28678) );
  XNOR U37507 ( .A(n28679), .B(n28680), .Z(n28677) );
  XNOR U37508 ( .A(y[4174]), .B(x[4174]), .Z(n28680) );
  XNOR U37509 ( .A(y[4175]), .B(x[4175]), .Z(n28679) );
  XOR U37510 ( .A(n28671), .B(n28670), .Z(n28672) );
  XNOR U37511 ( .A(n28666), .B(n28667), .Z(n28670) );
  XNOR U37512 ( .A(y[4170]), .B(x[4170]), .Z(n28667) );
  XNOR U37513 ( .A(n28668), .B(n28669), .Z(n28666) );
  XNOR U37514 ( .A(y[4171]), .B(x[4171]), .Z(n28669) );
  XNOR U37515 ( .A(y[4172]), .B(x[4172]), .Z(n28668) );
  XNOR U37516 ( .A(n28660), .B(n28661), .Z(n28671) );
  XNOR U37517 ( .A(y[4167]), .B(x[4167]), .Z(n28661) );
  XNOR U37518 ( .A(n28662), .B(n28663), .Z(n28660) );
  XNOR U37519 ( .A(y[4168]), .B(x[4168]), .Z(n28663) );
  XNOR U37520 ( .A(y[4169]), .B(x[4169]), .Z(n28662) );
  NAND U37521 ( .A(n28727), .B(n28728), .Z(N62845) );
  NANDN U37522 ( .A(n28729), .B(n28730), .Z(n28728) );
  OR U37523 ( .A(n28731), .B(n28732), .Z(n28730) );
  NAND U37524 ( .A(n28731), .B(n28732), .Z(n28727) );
  XOR U37525 ( .A(n28731), .B(n28733), .Z(N62844) );
  XNOR U37526 ( .A(n28729), .B(n28732), .Z(n28733) );
  AND U37527 ( .A(n28734), .B(n28735), .Z(n28732) );
  NANDN U37528 ( .A(n28736), .B(n28737), .Z(n28735) );
  NANDN U37529 ( .A(n28738), .B(n28739), .Z(n28737) );
  NANDN U37530 ( .A(n28739), .B(n28738), .Z(n28734) );
  NAND U37531 ( .A(n28740), .B(n28741), .Z(n28729) );
  NANDN U37532 ( .A(n28742), .B(n28743), .Z(n28741) );
  OR U37533 ( .A(n28744), .B(n28745), .Z(n28743) );
  NAND U37534 ( .A(n28745), .B(n28744), .Z(n28740) );
  AND U37535 ( .A(n28746), .B(n28747), .Z(n28731) );
  NANDN U37536 ( .A(n28748), .B(n28749), .Z(n28747) );
  NANDN U37537 ( .A(n28750), .B(n28751), .Z(n28749) );
  NANDN U37538 ( .A(n28751), .B(n28750), .Z(n28746) );
  XOR U37539 ( .A(n28745), .B(n28752), .Z(N62843) );
  XOR U37540 ( .A(n28742), .B(n28744), .Z(n28752) );
  XNOR U37541 ( .A(n28738), .B(n28753), .Z(n28744) );
  XNOR U37542 ( .A(n28736), .B(n28739), .Z(n28753) );
  NAND U37543 ( .A(n28754), .B(n28755), .Z(n28739) );
  NAND U37544 ( .A(n28756), .B(n28757), .Z(n28755) );
  OR U37545 ( .A(n28758), .B(n28759), .Z(n28756) );
  NANDN U37546 ( .A(n28760), .B(n28758), .Z(n28754) );
  IV U37547 ( .A(n28759), .Z(n28760) );
  NAND U37548 ( .A(n28761), .B(n28762), .Z(n28736) );
  NAND U37549 ( .A(n28763), .B(n28764), .Z(n28762) );
  NANDN U37550 ( .A(n28765), .B(n28766), .Z(n28763) );
  NANDN U37551 ( .A(n28766), .B(n28765), .Z(n28761) );
  AND U37552 ( .A(n28767), .B(n28768), .Z(n28738) );
  NAND U37553 ( .A(n28769), .B(n28770), .Z(n28768) );
  OR U37554 ( .A(n28771), .B(n28772), .Z(n28769) );
  NANDN U37555 ( .A(n28773), .B(n28771), .Z(n28767) );
  NAND U37556 ( .A(n28774), .B(n28775), .Z(n28742) );
  NANDN U37557 ( .A(n28776), .B(n28777), .Z(n28775) );
  OR U37558 ( .A(n28778), .B(n28779), .Z(n28777) );
  NANDN U37559 ( .A(n28780), .B(n28778), .Z(n28774) );
  IV U37560 ( .A(n28779), .Z(n28780) );
  XNOR U37561 ( .A(n28750), .B(n28781), .Z(n28745) );
  XNOR U37562 ( .A(n28748), .B(n28751), .Z(n28781) );
  NAND U37563 ( .A(n28782), .B(n28783), .Z(n28751) );
  NAND U37564 ( .A(n28784), .B(n28785), .Z(n28783) );
  OR U37565 ( .A(n28786), .B(n28787), .Z(n28784) );
  NANDN U37566 ( .A(n28788), .B(n28786), .Z(n28782) );
  IV U37567 ( .A(n28787), .Z(n28788) );
  NAND U37568 ( .A(n28789), .B(n28790), .Z(n28748) );
  NAND U37569 ( .A(n28791), .B(n28792), .Z(n28790) );
  NANDN U37570 ( .A(n28793), .B(n28794), .Z(n28791) );
  NANDN U37571 ( .A(n28794), .B(n28793), .Z(n28789) );
  AND U37572 ( .A(n28795), .B(n28796), .Z(n28750) );
  NAND U37573 ( .A(n28797), .B(n28798), .Z(n28796) );
  OR U37574 ( .A(n28799), .B(n28800), .Z(n28797) );
  NANDN U37575 ( .A(n28801), .B(n28799), .Z(n28795) );
  XNOR U37576 ( .A(n28776), .B(n28802), .Z(N62842) );
  XOR U37577 ( .A(n28778), .B(n28779), .Z(n28802) );
  XNOR U37578 ( .A(n28792), .B(n28803), .Z(n28779) );
  XOR U37579 ( .A(n28793), .B(n28794), .Z(n28803) );
  XOR U37580 ( .A(n28799), .B(n28804), .Z(n28794) );
  XOR U37581 ( .A(n28798), .B(n28801), .Z(n28804) );
  IV U37582 ( .A(n28800), .Z(n28801) );
  NAND U37583 ( .A(n28805), .B(n28806), .Z(n28800) );
  OR U37584 ( .A(n28807), .B(n28808), .Z(n28806) );
  OR U37585 ( .A(n28809), .B(n28810), .Z(n28805) );
  NAND U37586 ( .A(n28811), .B(n28812), .Z(n28798) );
  OR U37587 ( .A(n28813), .B(n28814), .Z(n28812) );
  OR U37588 ( .A(n28815), .B(n28816), .Z(n28811) );
  NOR U37589 ( .A(n28817), .B(n28818), .Z(n28799) );
  ANDN U37590 ( .B(n28819), .A(n28820), .Z(n28793) );
  XNOR U37591 ( .A(n28786), .B(n28821), .Z(n28792) );
  XNOR U37592 ( .A(n28785), .B(n28787), .Z(n28821) );
  NAND U37593 ( .A(n28822), .B(n28823), .Z(n28787) );
  OR U37594 ( .A(n28824), .B(n28825), .Z(n28823) );
  OR U37595 ( .A(n28826), .B(n28827), .Z(n28822) );
  NAND U37596 ( .A(n28828), .B(n28829), .Z(n28785) );
  OR U37597 ( .A(n28830), .B(n28831), .Z(n28829) );
  OR U37598 ( .A(n28832), .B(n28833), .Z(n28828) );
  ANDN U37599 ( .B(n28834), .A(n28835), .Z(n28786) );
  IV U37600 ( .A(n28836), .Z(n28834) );
  ANDN U37601 ( .B(n28837), .A(n28838), .Z(n28778) );
  XOR U37602 ( .A(n28764), .B(n28839), .Z(n28776) );
  XOR U37603 ( .A(n28765), .B(n28766), .Z(n28839) );
  XOR U37604 ( .A(n28771), .B(n28840), .Z(n28766) );
  XOR U37605 ( .A(n28770), .B(n28773), .Z(n28840) );
  IV U37606 ( .A(n28772), .Z(n28773) );
  NAND U37607 ( .A(n28841), .B(n28842), .Z(n28772) );
  OR U37608 ( .A(n28843), .B(n28844), .Z(n28842) );
  OR U37609 ( .A(n28845), .B(n28846), .Z(n28841) );
  NAND U37610 ( .A(n28847), .B(n28848), .Z(n28770) );
  OR U37611 ( .A(n28849), .B(n28850), .Z(n28848) );
  OR U37612 ( .A(n28851), .B(n28852), .Z(n28847) );
  NOR U37613 ( .A(n28853), .B(n28854), .Z(n28771) );
  ANDN U37614 ( .B(n28855), .A(n28856), .Z(n28765) );
  IV U37615 ( .A(n28857), .Z(n28855) );
  XNOR U37616 ( .A(n28758), .B(n28858), .Z(n28764) );
  XNOR U37617 ( .A(n28757), .B(n28759), .Z(n28858) );
  NAND U37618 ( .A(n28859), .B(n28860), .Z(n28759) );
  OR U37619 ( .A(n28861), .B(n28862), .Z(n28860) );
  OR U37620 ( .A(n28863), .B(n28864), .Z(n28859) );
  NAND U37621 ( .A(n28865), .B(n28866), .Z(n28757) );
  OR U37622 ( .A(n28867), .B(n28868), .Z(n28866) );
  OR U37623 ( .A(n28869), .B(n28870), .Z(n28865) );
  ANDN U37624 ( .B(n28871), .A(n28872), .Z(n28758) );
  IV U37625 ( .A(n28873), .Z(n28871) );
  XNOR U37626 ( .A(n28838), .B(n28837), .Z(N62841) );
  XOR U37627 ( .A(n28857), .B(n28856), .Z(n28837) );
  XNOR U37628 ( .A(n28872), .B(n28873), .Z(n28856) );
  XNOR U37629 ( .A(n28867), .B(n28868), .Z(n28873) );
  XNOR U37630 ( .A(n28869), .B(n28870), .Z(n28868) );
  XNOR U37631 ( .A(y[4165]), .B(x[4165]), .Z(n28870) );
  XNOR U37632 ( .A(y[4166]), .B(x[4166]), .Z(n28869) );
  XNOR U37633 ( .A(y[4164]), .B(x[4164]), .Z(n28867) );
  XNOR U37634 ( .A(n28861), .B(n28862), .Z(n28872) );
  XNOR U37635 ( .A(y[4161]), .B(x[4161]), .Z(n28862) );
  XNOR U37636 ( .A(n28863), .B(n28864), .Z(n28861) );
  XNOR U37637 ( .A(y[4162]), .B(x[4162]), .Z(n28864) );
  XNOR U37638 ( .A(y[4163]), .B(x[4163]), .Z(n28863) );
  XNOR U37639 ( .A(n28854), .B(n28853), .Z(n28857) );
  XNOR U37640 ( .A(n28849), .B(n28850), .Z(n28853) );
  XNOR U37641 ( .A(y[4158]), .B(x[4158]), .Z(n28850) );
  XNOR U37642 ( .A(n28851), .B(n28852), .Z(n28849) );
  XNOR U37643 ( .A(y[4159]), .B(x[4159]), .Z(n28852) );
  XNOR U37644 ( .A(y[4160]), .B(x[4160]), .Z(n28851) );
  XNOR U37645 ( .A(n28843), .B(n28844), .Z(n28854) );
  XNOR U37646 ( .A(y[4155]), .B(x[4155]), .Z(n28844) );
  XNOR U37647 ( .A(n28845), .B(n28846), .Z(n28843) );
  XNOR U37648 ( .A(y[4156]), .B(x[4156]), .Z(n28846) );
  XNOR U37649 ( .A(y[4157]), .B(x[4157]), .Z(n28845) );
  XOR U37650 ( .A(n28819), .B(n28820), .Z(n28838) );
  XNOR U37651 ( .A(n28835), .B(n28836), .Z(n28820) );
  XNOR U37652 ( .A(n28830), .B(n28831), .Z(n28836) );
  XNOR U37653 ( .A(n28832), .B(n28833), .Z(n28831) );
  XNOR U37654 ( .A(y[4153]), .B(x[4153]), .Z(n28833) );
  XNOR U37655 ( .A(y[4154]), .B(x[4154]), .Z(n28832) );
  XNOR U37656 ( .A(y[4152]), .B(x[4152]), .Z(n28830) );
  XNOR U37657 ( .A(n28824), .B(n28825), .Z(n28835) );
  XNOR U37658 ( .A(y[4149]), .B(x[4149]), .Z(n28825) );
  XNOR U37659 ( .A(n28826), .B(n28827), .Z(n28824) );
  XNOR U37660 ( .A(y[4150]), .B(x[4150]), .Z(n28827) );
  XNOR U37661 ( .A(y[4151]), .B(x[4151]), .Z(n28826) );
  XOR U37662 ( .A(n28818), .B(n28817), .Z(n28819) );
  XNOR U37663 ( .A(n28813), .B(n28814), .Z(n28817) );
  XNOR U37664 ( .A(y[4146]), .B(x[4146]), .Z(n28814) );
  XNOR U37665 ( .A(n28815), .B(n28816), .Z(n28813) );
  XNOR U37666 ( .A(y[4147]), .B(x[4147]), .Z(n28816) );
  XNOR U37667 ( .A(y[4148]), .B(x[4148]), .Z(n28815) );
  XNOR U37668 ( .A(n28807), .B(n28808), .Z(n28818) );
  XNOR U37669 ( .A(y[4143]), .B(x[4143]), .Z(n28808) );
  XNOR U37670 ( .A(n28809), .B(n28810), .Z(n28807) );
  XNOR U37671 ( .A(y[4144]), .B(x[4144]), .Z(n28810) );
  XNOR U37672 ( .A(y[4145]), .B(x[4145]), .Z(n28809) );
  NAND U37673 ( .A(n28874), .B(n28875), .Z(N62832) );
  NANDN U37674 ( .A(n28876), .B(n28877), .Z(n28875) );
  OR U37675 ( .A(n28878), .B(n28879), .Z(n28877) );
  NAND U37676 ( .A(n28878), .B(n28879), .Z(n28874) );
  XOR U37677 ( .A(n28878), .B(n28880), .Z(N62831) );
  XNOR U37678 ( .A(n28876), .B(n28879), .Z(n28880) );
  AND U37679 ( .A(n28881), .B(n28882), .Z(n28879) );
  NANDN U37680 ( .A(n28883), .B(n28884), .Z(n28882) );
  NANDN U37681 ( .A(n28885), .B(n28886), .Z(n28884) );
  NANDN U37682 ( .A(n28886), .B(n28885), .Z(n28881) );
  NAND U37683 ( .A(n28887), .B(n28888), .Z(n28876) );
  NANDN U37684 ( .A(n28889), .B(n28890), .Z(n28888) );
  OR U37685 ( .A(n28891), .B(n28892), .Z(n28890) );
  NAND U37686 ( .A(n28892), .B(n28891), .Z(n28887) );
  AND U37687 ( .A(n28893), .B(n28894), .Z(n28878) );
  NANDN U37688 ( .A(n28895), .B(n28896), .Z(n28894) );
  NANDN U37689 ( .A(n28897), .B(n28898), .Z(n28896) );
  NANDN U37690 ( .A(n28898), .B(n28897), .Z(n28893) );
  XOR U37691 ( .A(n28892), .B(n28899), .Z(N62830) );
  XOR U37692 ( .A(n28889), .B(n28891), .Z(n28899) );
  XNOR U37693 ( .A(n28885), .B(n28900), .Z(n28891) );
  XNOR U37694 ( .A(n28883), .B(n28886), .Z(n28900) );
  NAND U37695 ( .A(n28901), .B(n28902), .Z(n28886) );
  NAND U37696 ( .A(n28903), .B(n28904), .Z(n28902) );
  OR U37697 ( .A(n28905), .B(n28906), .Z(n28903) );
  NANDN U37698 ( .A(n28907), .B(n28905), .Z(n28901) );
  IV U37699 ( .A(n28906), .Z(n28907) );
  NAND U37700 ( .A(n28908), .B(n28909), .Z(n28883) );
  NAND U37701 ( .A(n28910), .B(n28911), .Z(n28909) );
  NANDN U37702 ( .A(n28912), .B(n28913), .Z(n28910) );
  NANDN U37703 ( .A(n28913), .B(n28912), .Z(n28908) );
  AND U37704 ( .A(n28914), .B(n28915), .Z(n28885) );
  NAND U37705 ( .A(n28916), .B(n28917), .Z(n28915) );
  OR U37706 ( .A(n28918), .B(n28919), .Z(n28916) );
  NANDN U37707 ( .A(n28920), .B(n28918), .Z(n28914) );
  NAND U37708 ( .A(n28921), .B(n28922), .Z(n28889) );
  NANDN U37709 ( .A(n28923), .B(n28924), .Z(n28922) );
  OR U37710 ( .A(n28925), .B(n28926), .Z(n28924) );
  NANDN U37711 ( .A(n28927), .B(n28925), .Z(n28921) );
  IV U37712 ( .A(n28926), .Z(n28927) );
  XNOR U37713 ( .A(n28897), .B(n28928), .Z(n28892) );
  XNOR U37714 ( .A(n28895), .B(n28898), .Z(n28928) );
  NAND U37715 ( .A(n28929), .B(n28930), .Z(n28898) );
  NAND U37716 ( .A(n28931), .B(n28932), .Z(n28930) );
  OR U37717 ( .A(n28933), .B(n28934), .Z(n28931) );
  NANDN U37718 ( .A(n28935), .B(n28933), .Z(n28929) );
  IV U37719 ( .A(n28934), .Z(n28935) );
  NAND U37720 ( .A(n28936), .B(n28937), .Z(n28895) );
  NAND U37721 ( .A(n28938), .B(n28939), .Z(n28937) );
  NANDN U37722 ( .A(n28940), .B(n28941), .Z(n28938) );
  NANDN U37723 ( .A(n28941), .B(n28940), .Z(n28936) );
  AND U37724 ( .A(n28942), .B(n28943), .Z(n28897) );
  NAND U37725 ( .A(n28944), .B(n28945), .Z(n28943) );
  OR U37726 ( .A(n28946), .B(n28947), .Z(n28944) );
  NANDN U37727 ( .A(n28948), .B(n28946), .Z(n28942) );
  XNOR U37728 ( .A(n28923), .B(n28949), .Z(N62829) );
  XOR U37729 ( .A(n28925), .B(n28926), .Z(n28949) );
  XNOR U37730 ( .A(n28939), .B(n28950), .Z(n28926) );
  XOR U37731 ( .A(n28940), .B(n28941), .Z(n28950) );
  XOR U37732 ( .A(n28946), .B(n28951), .Z(n28941) );
  XOR U37733 ( .A(n28945), .B(n28948), .Z(n28951) );
  IV U37734 ( .A(n28947), .Z(n28948) );
  NAND U37735 ( .A(n28952), .B(n28953), .Z(n28947) );
  OR U37736 ( .A(n28954), .B(n28955), .Z(n28953) );
  OR U37737 ( .A(n28956), .B(n28957), .Z(n28952) );
  NAND U37738 ( .A(n28958), .B(n28959), .Z(n28945) );
  OR U37739 ( .A(n28960), .B(n28961), .Z(n28959) );
  OR U37740 ( .A(n28962), .B(n28963), .Z(n28958) );
  NOR U37741 ( .A(n28964), .B(n28965), .Z(n28946) );
  ANDN U37742 ( .B(n28966), .A(n28967), .Z(n28940) );
  XNOR U37743 ( .A(n28933), .B(n28968), .Z(n28939) );
  XNOR U37744 ( .A(n28932), .B(n28934), .Z(n28968) );
  NAND U37745 ( .A(n28969), .B(n28970), .Z(n28934) );
  OR U37746 ( .A(n28971), .B(n28972), .Z(n28970) );
  OR U37747 ( .A(n28973), .B(n28974), .Z(n28969) );
  NAND U37748 ( .A(n28975), .B(n28976), .Z(n28932) );
  OR U37749 ( .A(n28977), .B(n28978), .Z(n28976) );
  OR U37750 ( .A(n28979), .B(n28980), .Z(n28975) );
  ANDN U37751 ( .B(n28981), .A(n28982), .Z(n28933) );
  IV U37752 ( .A(n28983), .Z(n28981) );
  ANDN U37753 ( .B(n28984), .A(n28985), .Z(n28925) );
  XOR U37754 ( .A(n28911), .B(n28986), .Z(n28923) );
  XOR U37755 ( .A(n28912), .B(n28913), .Z(n28986) );
  XOR U37756 ( .A(n28918), .B(n28987), .Z(n28913) );
  XOR U37757 ( .A(n28917), .B(n28920), .Z(n28987) );
  IV U37758 ( .A(n28919), .Z(n28920) );
  NAND U37759 ( .A(n28988), .B(n28989), .Z(n28919) );
  OR U37760 ( .A(n28990), .B(n28991), .Z(n28989) );
  OR U37761 ( .A(n28992), .B(n28993), .Z(n28988) );
  NAND U37762 ( .A(n28994), .B(n28995), .Z(n28917) );
  OR U37763 ( .A(n28996), .B(n28997), .Z(n28995) );
  OR U37764 ( .A(n28998), .B(n28999), .Z(n28994) );
  NOR U37765 ( .A(n29000), .B(n29001), .Z(n28918) );
  ANDN U37766 ( .B(n29002), .A(n29003), .Z(n28912) );
  IV U37767 ( .A(n29004), .Z(n29002) );
  XNOR U37768 ( .A(n28905), .B(n29005), .Z(n28911) );
  XNOR U37769 ( .A(n28904), .B(n28906), .Z(n29005) );
  NAND U37770 ( .A(n29006), .B(n29007), .Z(n28906) );
  OR U37771 ( .A(n29008), .B(n29009), .Z(n29007) );
  OR U37772 ( .A(n29010), .B(n29011), .Z(n29006) );
  NAND U37773 ( .A(n29012), .B(n29013), .Z(n28904) );
  OR U37774 ( .A(n29014), .B(n29015), .Z(n29013) );
  OR U37775 ( .A(n29016), .B(n29017), .Z(n29012) );
  ANDN U37776 ( .B(n29018), .A(n29019), .Z(n28905) );
  IV U37777 ( .A(n29020), .Z(n29018) );
  XNOR U37778 ( .A(n28985), .B(n28984), .Z(N62828) );
  XOR U37779 ( .A(n29004), .B(n29003), .Z(n28984) );
  XNOR U37780 ( .A(n29019), .B(n29020), .Z(n29003) );
  XNOR U37781 ( .A(n29014), .B(n29015), .Z(n29020) );
  XNOR U37782 ( .A(n29016), .B(n29017), .Z(n29015) );
  XNOR U37783 ( .A(y[4141]), .B(x[4141]), .Z(n29017) );
  XNOR U37784 ( .A(y[4142]), .B(x[4142]), .Z(n29016) );
  XNOR U37785 ( .A(y[4140]), .B(x[4140]), .Z(n29014) );
  XNOR U37786 ( .A(n29008), .B(n29009), .Z(n29019) );
  XNOR U37787 ( .A(y[4137]), .B(x[4137]), .Z(n29009) );
  XNOR U37788 ( .A(n29010), .B(n29011), .Z(n29008) );
  XNOR U37789 ( .A(y[4138]), .B(x[4138]), .Z(n29011) );
  XNOR U37790 ( .A(y[4139]), .B(x[4139]), .Z(n29010) );
  XNOR U37791 ( .A(n29001), .B(n29000), .Z(n29004) );
  XNOR U37792 ( .A(n28996), .B(n28997), .Z(n29000) );
  XNOR U37793 ( .A(y[4134]), .B(x[4134]), .Z(n28997) );
  XNOR U37794 ( .A(n28998), .B(n28999), .Z(n28996) );
  XNOR U37795 ( .A(y[4135]), .B(x[4135]), .Z(n28999) );
  XNOR U37796 ( .A(y[4136]), .B(x[4136]), .Z(n28998) );
  XNOR U37797 ( .A(n28990), .B(n28991), .Z(n29001) );
  XNOR U37798 ( .A(y[4131]), .B(x[4131]), .Z(n28991) );
  XNOR U37799 ( .A(n28992), .B(n28993), .Z(n28990) );
  XNOR U37800 ( .A(y[4132]), .B(x[4132]), .Z(n28993) );
  XNOR U37801 ( .A(y[4133]), .B(x[4133]), .Z(n28992) );
  XOR U37802 ( .A(n28966), .B(n28967), .Z(n28985) );
  XNOR U37803 ( .A(n28982), .B(n28983), .Z(n28967) );
  XNOR U37804 ( .A(n28977), .B(n28978), .Z(n28983) );
  XNOR U37805 ( .A(n28979), .B(n28980), .Z(n28978) );
  XNOR U37806 ( .A(y[4129]), .B(x[4129]), .Z(n28980) );
  XNOR U37807 ( .A(y[4130]), .B(x[4130]), .Z(n28979) );
  XNOR U37808 ( .A(y[4128]), .B(x[4128]), .Z(n28977) );
  XNOR U37809 ( .A(n28971), .B(n28972), .Z(n28982) );
  XNOR U37810 ( .A(y[4125]), .B(x[4125]), .Z(n28972) );
  XNOR U37811 ( .A(n28973), .B(n28974), .Z(n28971) );
  XNOR U37812 ( .A(y[4126]), .B(x[4126]), .Z(n28974) );
  XNOR U37813 ( .A(y[4127]), .B(x[4127]), .Z(n28973) );
  XOR U37814 ( .A(n28965), .B(n28964), .Z(n28966) );
  XNOR U37815 ( .A(n28960), .B(n28961), .Z(n28964) );
  XNOR U37816 ( .A(y[4122]), .B(x[4122]), .Z(n28961) );
  XNOR U37817 ( .A(n28962), .B(n28963), .Z(n28960) );
  XNOR U37818 ( .A(y[4123]), .B(x[4123]), .Z(n28963) );
  XNOR U37819 ( .A(y[4124]), .B(x[4124]), .Z(n28962) );
  XNOR U37820 ( .A(n28954), .B(n28955), .Z(n28965) );
  XNOR U37821 ( .A(y[4119]), .B(x[4119]), .Z(n28955) );
  XNOR U37822 ( .A(n28956), .B(n28957), .Z(n28954) );
  XNOR U37823 ( .A(y[4120]), .B(x[4120]), .Z(n28957) );
  XNOR U37824 ( .A(y[4121]), .B(x[4121]), .Z(n28956) );
  NAND U37825 ( .A(n29021), .B(n29022), .Z(N62819) );
  NANDN U37826 ( .A(n29023), .B(n29024), .Z(n29022) );
  OR U37827 ( .A(n29025), .B(n29026), .Z(n29024) );
  NAND U37828 ( .A(n29025), .B(n29026), .Z(n29021) );
  XOR U37829 ( .A(n29025), .B(n29027), .Z(N62818) );
  XNOR U37830 ( .A(n29023), .B(n29026), .Z(n29027) );
  AND U37831 ( .A(n29028), .B(n29029), .Z(n29026) );
  NANDN U37832 ( .A(n29030), .B(n29031), .Z(n29029) );
  NANDN U37833 ( .A(n29032), .B(n29033), .Z(n29031) );
  NANDN U37834 ( .A(n29033), .B(n29032), .Z(n29028) );
  NAND U37835 ( .A(n29034), .B(n29035), .Z(n29023) );
  NANDN U37836 ( .A(n29036), .B(n29037), .Z(n29035) );
  OR U37837 ( .A(n29038), .B(n29039), .Z(n29037) );
  NAND U37838 ( .A(n29039), .B(n29038), .Z(n29034) );
  AND U37839 ( .A(n29040), .B(n29041), .Z(n29025) );
  NANDN U37840 ( .A(n29042), .B(n29043), .Z(n29041) );
  NANDN U37841 ( .A(n29044), .B(n29045), .Z(n29043) );
  NANDN U37842 ( .A(n29045), .B(n29044), .Z(n29040) );
  XOR U37843 ( .A(n29039), .B(n29046), .Z(N62817) );
  XOR U37844 ( .A(n29036), .B(n29038), .Z(n29046) );
  XNOR U37845 ( .A(n29032), .B(n29047), .Z(n29038) );
  XNOR U37846 ( .A(n29030), .B(n29033), .Z(n29047) );
  NAND U37847 ( .A(n29048), .B(n29049), .Z(n29033) );
  NAND U37848 ( .A(n29050), .B(n29051), .Z(n29049) );
  OR U37849 ( .A(n29052), .B(n29053), .Z(n29050) );
  NANDN U37850 ( .A(n29054), .B(n29052), .Z(n29048) );
  IV U37851 ( .A(n29053), .Z(n29054) );
  NAND U37852 ( .A(n29055), .B(n29056), .Z(n29030) );
  NAND U37853 ( .A(n29057), .B(n29058), .Z(n29056) );
  NANDN U37854 ( .A(n29059), .B(n29060), .Z(n29057) );
  NANDN U37855 ( .A(n29060), .B(n29059), .Z(n29055) );
  AND U37856 ( .A(n29061), .B(n29062), .Z(n29032) );
  NAND U37857 ( .A(n29063), .B(n29064), .Z(n29062) );
  OR U37858 ( .A(n29065), .B(n29066), .Z(n29063) );
  NANDN U37859 ( .A(n29067), .B(n29065), .Z(n29061) );
  NAND U37860 ( .A(n29068), .B(n29069), .Z(n29036) );
  NANDN U37861 ( .A(n29070), .B(n29071), .Z(n29069) );
  OR U37862 ( .A(n29072), .B(n29073), .Z(n29071) );
  NANDN U37863 ( .A(n29074), .B(n29072), .Z(n29068) );
  IV U37864 ( .A(n29073), .Z(n29074) );
  XNOR U37865 ( .A(n29044), .B(n29075), .Z(n29039) );
  XNOR U37866 ( .A(n29042), .B(n29045), .Z(n29075) );
  NAND U37867 ( .A(n29076), .B(n29077), .Z(n29045) );
  NAND U37868 ( .A(n29078), .B(n29079), .Z(n29077) );
  OR U37869 ( .A(n29080), .B(n29081), .Z(n29078) );
  NANDN U37870 ( .A(n29082), .B(n29080), .Z(n29076) );
  IV U37871 ( .A(n29081), .Z(n29082) );
  NAND U37872 ( .A(n29083), .B(n29084), .Z(n29042) );
  NAND U37873 ( .A(n29085), .B(n29086), .Z(n29084) );
  NANDN U37874 ( .A(n29087), .B(n29088), .Z(n29085) );
  NANDN U37875 ( .A(n29088), .B(n29087), .Z(n29083) );
  AND U37876 ( .A(n29089), .B(n29090), .Z(n29044) );
  NAND U37877 ( .A(n29091), .B(n29092), .Z(n29090) );
  OR U37878 ( .A(n29093), .B(n29094), .Z(n29091) );
  NANDN U37879 ( .A(n29095), .B(n29093), .Z(n29089) );
  XNOR U37880 ( .A(n29070), .B(n29096), .Z(N62816) );
  XOR U37881 ( .A(n29072), .B(n29073), .Z(n29096) );
  XNOR U37882 ( .A(n29086), .B(n29097), .Z(n29073) );
  XOR U37883 ( .A(n29087), .B(n29088), .Z(n29097) );
  XOR U37884 ( .A(n29093), .B(n29098), .Z(n29088) );
  XOR U37885 ( .A(n29092), .B(n29095), .Z(n29098) );
  IV U37886 ( .A(n29094), .Z(n29095) );
  NAND U37887 ( .A(n29099), .B(n29100), .Z(n29094) );
  OR U37888 ( .A(n29101), .B(n29102), .Z(n29100) );
  OR U37889 ( .A(n29103), .B(n29104), .Z(n29099) );
  NAND U37890 ( .A(n29105), .B(n29106), .Z(n29092) );
  OR U37891 ( .A(n29107), .B(n29108), .Z(n29106) );
  OR U37892 ( .A(n29109), .B(n29110), .Z(n29105) );
  NOR U37893 ( .A(n29111), .B(n29112), .Z(n29093) );
  ANDN U37894 ( .B(n29113), .A(n29114), .Z(n29087) );
  XNOR U37895 ( .A(n29080), .B(n29115), .Z(n29086) );
  XNOR U37896 ( .A(n29079), .B(n29081), .Z(n29115) );
  NAND U37897 ( .A(n29116), .B(n29117), .Z(n29081) );
  OR U37898 ( .A(n29118), .B(n29119), .Z(n29117) );
  OR U37899 ( .A(n29120), .B(n29121), .Z(n29116) );
  NAND U37900 ( .A(n29122), .B(n29123), .Z(n29079) );
  OR U37901 ( .A(n29124), .B(n29125), .Z(n29123) );
  OR U37902 ( .A(n29126), .B(n29127), .Z(n29122) );
  ANDN U37903 ( .B(n29128), .A(n29129), .Z(n29080) );
  IV U37904 ( .A(n29130), .Z(n29128) );
  ANDN U37905 ( .B(n29131), .A(n29132), .Z(n29072) );
  XOR U37906 ( .A(n29058), .B(n29133), .Z(n29070) );
  XOR U37907 ( .A(n29059), .B(n29060), .Z(n29133) );
  XOR U37908 ( .A(n29065), .B(n29134), .Z(n29060) );
  XOR U37909 ( .A(n29064), .B(n29067), .Z(n29134) );
  IV U37910 ( .A(n29066), .Z(n29067) );
  NAND U37911 ( .A(n29135), .B(n29136), .Z(n29066) );
  OR U37912 ( .A(n29137), .B(n29138), .Z(n29136) );
  OR U37913 ( .A(n29139), .B(n29140), .Z(n29135) );
  NAND U37914 ( .A(n29141), .B(n29142), .Z(n29064) );
  OR U37915 ( .A(n29143), .B(n29144), .Z(n29142) );
  OR U37916 ( .A(n29145), .B(n29146), .Z(n29141) );
  NOR U37917 ( .A(n29147), .B(n29148), .Z(n29065) );
  ANDN U37918 ( .B(n29149), .A(n29150), .Z(n29059) );
  IV U37919 ( .A(n29151), .Z(n29149) );
  XNOR U37920 ( .A(n29052), .B(n29152), .Z(n29058) );
  XNOR U37921 ( .A(n29051), .B(n29053), .Z(n29152) );
  NAND U37922 ( .A(n29153), .B(n29154), .Z(n29053) );
  OR U37923 ( .A(n29155), .B(n29156), .Z(n29154) );
  OR U37924 ( .A(n29157), .B(n29158), .Z(n29153) );
  NAND U37925 ( .A(n29159), .B(n29160), .Z(n29051) );
  OR U37926 ( .A(n29161), .B(n29162), .Z(n29160) );
  OR U37927 ( .A(n29163), .B(n29164), .Z(n29159) );
  ANDN U37928 ( .B(n29165), .A(n29166), .Z(n29052) );
  IV U37929 ( .A(n29167), .Z(n29165) );
  XNOR U37930 ( .A(n29132), .B(n29131), .Z(N62815) );
  XOR U37931 ( .A(n29151), .B(n29150), .Z(n29131) );
  XNOR U37932 ( .A(n29166), .B(n29167), .Z(n29150) );
  XNOR U37933 ( .A(n29161), .B(n29162), .Z(n29167) );
  XNOR U37934 ( .A(n29163), .B(n29164), .Z(n29162) );
  XNOR U37935 ( .A(y[4117]), .B(x[4117]), .Z(n29164) );
  XNOR U37936 ( .A(y[4118]), .B(x[4118]), .Z(n29163) );
  XNOR U37937 ( .A(y[4116]), .B(x[4116]), .Z(n29161) );
  XNOR U37938 ( .A(n29155), .B(n29156), .Z(n29166) );
  XNOR U37939 ( .A(y[4113]), .B(x[4113]), .Z(n29156) );
  XNOR U37940 ( .A(n29157), .B(n29158), .Z(n29155) );
  XNOR U37941 ( .A(y[4114]), .B(x[4114]), .Z(n29158) );
  XNOR U37942 ( .A(y[4115]), .B(x[4115]), .Z(n29157) );
  XNOR U37943 ( .A(n29148), .B(n29147), .Z(n29151) );
  XNOR U37944 ( .A(n29143), .B(n29144), .Z(n29147) );
  XNOR U37945 ( .A(y[4110]), .B(x[4110]), .Z(n29144) );
  XNOR U37946 ( .A(n29145), .B(n29146), .Z(n29143) );
  XNOR U37947 ( .A(y[4111]), .B(x[4111]), .Z(n29146) );
  XNOR U37948 ( .A(y[4112]), .B(x[4112]), .Z(n29145) );
  XNOR U37949 ( .A(n29137), .B(n29138), .Z(n29148) );
  XNOR U37950 ( .A(y[4107]), .B(x[4107]), .Z(n29138) );
  XNOR U37951 ( .A(n29139), .B(n29140), .Z(n29137) );
  XNOR U37952 ( .A(y[4108]), .B(x[4108]), .Z(n29140) );
  XNOR U37953 ( .A(y[4109]), .B(x[4109]), .Z(n29139) );
  XOR U37954 ( .A(n29113), .B(n29114), .Z(n29132) );
  XNOR U37955 ( .A(n29129), .B(n29130), .Z(n29114) );
  XNOR U37956 ( .A(n29124), .B(n29125), .Z(n29130) );
  XNOR U37957 ( .A(n29126), .B(n29127), .Z(n29125) );
  XNOR U37958 ( .A(y[4105]), .B(x[4105]), .Z(n29127) );
  XNOR U37959 ( .A(y[4106]), .B(x[4106]), .Z(n29126) );
  XNOR U37960 ( .A(y[4104]), .B(x[4104]), .Z(n29124) );
  XNOR U37961 ( .A(n29118), .B(n29119), .Z(n29129) );
  XNOR U37962 ( .A(y[4101]), .B(x[4101]), .Z(n29119) );
  XNOR U37963 ( .A(n29120), .B(n29121), .Z(n29118) );
  XNOR U37964 ( .A(y[4102]), .B(x[4102]), .Z(n29121) );
  XNOR U37965 ( .A(y[4103]), .B(x[4103]), .Z(n29120) );
  XOR U37966 ( .A(n29112), .B(n29111), .Z(n29113) );
  XNOR U37967 ( .A(n29107), .B(n29108), .Z(n29111) );
  XNOR U37968 ( .A(y[4098]), .B(x[4098]), .Z(n29108) );
  XNOR U37969 ( .A(n29109), .B(n29110), .Z(n29107) );
  XNOR U37970 ( .A(y[4099]), .B(x[4099]), .Z(n29110) );
  XNOR U37971 ( .A(y[4100]), .B(x[4100]), .Z(n29109) );
  XNOR U37972 ( .A(n29101), .B(n29102), .Z(n29112) );
  XNOR U37973 ( .A(y[4095]), .B(x[4095]), .Z(n29102) );
  XNOR U37974 ( .A(n29103), .B(n29104), .Z(n29101) );
  XNOR U37975 ( .A(y[4096]), .B(x[4096]), .Z(n29104) );
  XNOR U37976 ( .A(y[4097]), .B(x[4097]), .Z(n29103) );
  NAND U37977 ( .A(n29168), .B(n29169), .Z(N62806) );
  NANDN U37978 ( .A(n29170), .B(n29171), .Z(n29169) );
  OR U37979 ( .A(n29172), .B(n29173), .Z(n29171) );
  NAND U37980 ( .A(n29172), .B(n29173), .Z(n29168) );
  XOR U37981 ( .A(n29172), .B(n29174), .Z(N62805) );
  XNOR U37982 ( .A(n29170), .B(n29173), .Z(n29174) );
  AND U37983 ( .A(n29175), .B(n29176), .Z(n29173) );
  NANDN U37984 ( .A(n29177), .B(n29178), .Z(n29176) );
  NANDN U37985 ( .A(n29179), .B(n29180), .Z(n29178) );
  NANDN U37986 ( .A(n29180), .B(n29179), .Z(n29175) );
  NAND U37987 ( .A(n29181), .B(n29182), .Z(n29170) );
  NANDN U37988 ( .A(n29183), .B(n29184), .Z(n29182) );
  OR U37989 ( .A(n29185), .B(n29186), .Z(n29184) );
  NAND U37990 ( .A(n29186), .B(n29185), .Z(n29181) );
  AND U37991 ( .A(n29187), .B(n29188), .Z(n29172) );
  NANDN U37992 ( .A(n29189), .B(n29190), .Z(n29188) );
  NANDN U37993 ( .A(n29191), .B(n29192), .Z(n29190) );
  NANDN U37994 ( .A(n29192), .B(n29191), .Z(n29187) );
  XOR U37995 ( .A(n29186), .B(n29193), .Z(N62804) );
  XOR U37996 ( .A(n29183), .B(n29185), .Z(n29193) );
  XNOR U37997 ( .A(n29179), .B(n29194), .Z(n29185) );
  XNOR U37998 ( .A(n29177), .B(n29180), .Z(n29194) );
  NAND U37999 ( .A(n29195), .B(n29196), .Z(n29180) );
  NAND U38000 ( .A(n29197), .B(n29198), .Z(n29196) );
  OR U38001 ( .A(n29199), .B(n29200), .Z(n29197) );
  NANDN U38002 ( .A(n29201), .B(n29199), .Z(n29195) );
  IV U38003 ( .A(n29200), .Z(n29201) );
  NAND U38004 ( .A(n29202), .B(n29203), .Z(n29177) );
  NAND U38005 ( .A(n29204), .B(n29205), .Z(n29203) );
  NANDN U38006 ( .A(n29206), .B(n29207), .Z(n29204) );
  NANDN U38007 ( .A(n29207), .B(n29206), .Z(n29202) );
  AND U38008 ( .A(n29208), .B(n29209), .Z(n29179) );
  NAND U38009 ( .A(n29210), .B(n29211), .Z(n29209) );
  OR U38010 ( .A(n29212), .B(n29213), .Z(n29210) );
  NANDN U38011 ( .A(n29214), .B(n29212), .Z(n29208) );
  NAND U38012 ( .A(n29215), .B(n29216), .Z(n29183) );
  NANDN U38013 ( .A(n29217), .B(n29218), .Z(n29216) );
  OR U38014 ( .A(n29219), .B(n29220), .Z(n29218) );
  NANDN U38015 ( .A(n29221), .B(n29219), .Z(n29215) );
  IV U38016 ( .A(n29220), .Z(n29221) );
  XNOR U38017 ( .A(n29191), .B(n29222), .Z(n29186) );
  XNOR U38018 ( .A(n29189), .B(n29192), .Z(n29222) );
  NAND U38019 ( .A(n29223), .B(n29224), .Z(n29192) );
  NAND U38020 ( .A(n29225), .B(n29226), .Z(n29224) );
  OR U38021 ( .A(n29227), .B(n29228), .Z(n29225) );
  NANDN U38022 ( .A(n29229), .B(n29227), .Z(n29223) );
  IV U38023 ( .A(n29228), .Z(n29229) );
  NAND U38024 ( .A(n29230), .B(n29231), .Z(n29189) );
  NAND U38025 ( .A(n29232), .B(n29233), .Z(n29231) );
  NANDN U38026 ( .A(n29234), .B(n29235), .Z(n29232) );
  NANDN U38027 ( .A(n29235), .B(n29234), .Z(n29230) );
  AND U38028 ( .A(n29236), .B(n29237), .Z(n29191) );
  NAND U38029 ( .A(n29238), .B(n29239), .Z(n29237) );
  OR U38030 ( .A(n29240), .B(n29241), .Z(n29238) );
  NANDN U38031 ( .A(n29242), .B(n29240), .Z(n29236) );
  XNOR U38032 ( .A(n29217), .B(n29243), .Z(N62803) );
  XOR U38033 ( .A(n29219), .B(n29220), .Z(n29243) );
  XNOR U38034 ( .A(n29233), .B(n29244), .Z(n29220) );
  XOR U38035 ( .A(n29234), .B(n29235), .Z(n29244) );
  XOR U38036 ( .A(n29240), .B(n29245), .Z(n29235) );
  XOR U38037 ( .A(n29239), .B(n29242), .Z(n29245) );
  IV U38038 ( .A(n29241), .Z(n29242) );
  NAND U38039 ( .A(n29246), .B(n29247), .Z(n29241) );
  OR U38040 ( .A(n29248), .B(n29249), .Z(n29247) );
  OR U38041 ( .A(n29250), .B(n29251), .Z(n29246) );
  NAND U38042 ( .A(n29252), .B(n29253), .Z(n29239) );
  OR U38043 ( .A(n29254), .B(n29255), .Z(n29253) );
  OR U38044 ( .A(n29256), .B(n29257), .Z(n29252) );
  NOR U38045 ( .A(n29258), .B(n29259), .Z(n29240) );
  ANDN U38046 ( .B(n29260), .A(n29261), .Z(n29234) );
  XNOR U38047 ( .A(n29227), .B(n29262), .Z(n29233) );
  XNOR U38048 ( .A(n29226), .B(n29228), .Z(n29262) );
  NAND U38049 ( .A(n29263), .B(n29264), .Z(n29228) );
  OR U38050 ( .A(n29265), .B(n29266), .Z(n29264) );
  OR U38051 ( .A(n29267), .B(n29268), .Z(n29263) );
  NAND U38052 ( .A(n29269), .B(n29270), .Z(n29226) );
  OR U38053 ( .A(n29271), .B(n29272), .Z(n29270) );
  OR U38054 ( .A(n29273), .B(n29274), .Z(n29269) );
  ANDN U38055 ( .B(n29275), .A(n29276), .Z(n29227) );
  IV U38056 ( .A(n29277), .Z(n29275) );
  ANDN U38057 ( .B(n29278), .A(n29279), .Z(n29219) );
  XOR U38058 ( .A(n29205), .B(n29280), .Z(n29217) );
  XOR U38059 ( .A(n29206), .B(n29207), .Z(n29280) );
  XOR U38060 ( .A(n29212), .B(n29281), .Z(n29207) );
  XOR U38061 ( .A(n29211), .B(n29214), .Z(n29281) );
  IV U38062 ( .A(n29213), .Z(n29214) );
  NAND U38063 ( .A(n29282), .B(n29283), .Z(n29213) );
  OR U38064 ( .A(n29284), .B(n29285), .Z(n29283) );
  OR U38065 ( .A(n29286), .B(n29287), .Z(n29282) );
  NAND U38066 ( .A(n29288), .B(n29289), .Z(n29211) );
  OR U38067 ( .A(n29290), .B(n29291), .Z(n29289) );
  OR U38068 ( .A(n29292), .B(n29293), .Z(n29288) );
  NOR U38069 ( .A(n29294), .B(n29295), .Z(n29212) );
  ANDN U38070 ( .B(n29296), .A(n29297), .Z(n29206) );
  IV U38071 ( .A(n29298), .Z(n29296) );
  XNOR U38072 ( .A(n29199), .B(n29299), .Z(n29205) );
  XNOR U38073 ( .A(n29198), .B(n29200), .Z(n29299) );
  NAND U38074 ( .A(n29300), .B(n29301), .Z(n29200) );
  OR U38075 ( .A(n29302), .B(n29303), .Z(n29301) );
  OR U38076 ( .A(n29304), .B(n29305), .Z(n29300) );
  NAND U38077 ( .A(n29306), .B(n29307), .Z(n29198) );
  OR U38078 ( .A(n29308), .B(n29309), .Z(n29307) );
  OR U38079 ( .A(n29310), .B(n29311), .Z(n29306) );
  ANDN U38080 ( .B(n29312), .A(n29313), .Z(n29199) );
  IV U38081 ( .A(n29314), .Z(n29312) );
  XNOR U38082 ( .A(n29279), .B(n29278), .Z(N62802) );
  XOR U38083 ( .A(n29298), .B(n29297), .Z(n29278) );
  XNOR U38084 ( .A(n29313), .B(n29314), .Z(n29297) );
  XNOR U38085 ( .A(n29308), .B(n29309), .Z(n29314) );
  XNOR U38086 ( .A(n29310), .B(n29311), .Z(n29309) );
  XNOR U38087 ( .A(y[4093]), .B(x[4093]), .Z(n29311) );
  XNOR U38088 ( .A(y[4094]), .B(x[4094]), .Z(n29310) );
  XNOR U38089 ( .A(y[4092]), .B(x[4092]), .Z(n29308) );
  XNOR U38090 ( .A(n29302), .B(n29303), .Z(n29313) );
  XNOR U38091 ( .A(y[4089]), .B(x[4089]), .Z(n29303) );
  XNOR U38092 ( .A(n29304), .B(n29305), .Z(n29302) );
  XNOR U38093 ( .A(y[4090]), .B(x[4090]), .Z(n29305) );
  XNOR U38094 ( .A(y[4091]), .B(x[4091]), .Z(n29304) );
  XNOR U38095 ( .A(n29295), .B(n29294), .Z(n29298) );
  XNOR U38096 ( .A(n29290), .B(n29291), .Z(n29294) );
  XNOR U38097 ( .A(y[4086]), .B(x[4086]), .Z(n29291) );
  XNOR U38098 ( .A(n29292), .B(n29293), .Z(n29290) );
  XNOR U38099 ( .A(y[4087]), .B(x[4087]), .Z(n29293) );
  XNOR U38100 ( .A(y[4088]), .B(x[4088]), .Z(n29292) );
  XNOR U38101 ( .A(n29284), .B(n29285), .Z(n29295) );
  XNOR U38102 ( .A(y[4083]), .B(x[4083]), .Z(n29285) );
  XNOR U38103 ( .A(n29286), .B(n29287), .Z(n29284) );
  XNOR U38104 ( .A(y[4084]), .B(x[4084]), .Z(n29287) );
  XNOR U38105 ( .A(y[4085]), .B(x[4085]), .Z(n29286) );
  XOR U38106 ( .A(n29260), .B(n29261), .Z(n29279) );
  XNOR U38107 ( .A(n29276), .B(n29277), .Z(n29261) );
  XNOR U38108 ( .A(n29271), .B(n29272), .Z(n29277) );
  XNOR U38109 ( .A(n29273), .B(n29274), .Z(n29272) );
  XNOR U38110 ( .A(y[4081]), .B(x[4081]), .Z(n29274) );
  XNOR U38111 ( .A(y[4082]), .B(x[4082]), .Z(n29273) );
  XNOR U38112 ( .A(y[4080]), .B(x[4080]), .Z(n29271) );
  XNOR U38113 ( .A(n29265), .B(n29266), .Z(n29276) );
  XNOR U38114 ( .A(y[4077]), .B(x[4077]), .Z(n29266) );
  XNOR U38115 ( .A(n29267), .B(n29268), .Z(n29265) );
  XNOR U38116 ( .A(y[4078]), .B(x[4078]), .Z(n29268) );
  XNOR U38117 ( .A(y[4079]), .B(x[4079]), .Z(n29267) );
  XOR U38118 ( .A(n29259), .B(n29258), .Z(n29260) );
  XNOR U38119 ( .A(n29254), .B(n29255), .Z(n29258) );
  XNOR U38120 ( .A(y[4074]), .B(x[4074]), .Z(n29255) );
  XNOR U38121 ( .A(n29256), .B(n29257), .Z(n29254) );
  XNOR U38122 ( .A(y[4075]), .B(x[4075]), .Z(n29257) );
  XNOR U38123 ( .A(y[4076]), .B(x[4076]), .Z(n29256) );
  XNOR U38124 ( .A(n29248), .B(n29249), .Z(n29259) );
  XNOR U38125 ( .A(y[4071]), .B(x[4071]), .Z(n29249) );
  XNOR U38126 ( .A(n29250), .B(n29251), .Z(n29248) );
  XNOR U38127 ( .A(y[4072]), .B(x[4072]), .Z(n29251) );
  XNOR U38128 ( .A(y[4073]), .B(x[4073]), .Z(n29250) );
  NAND U38129 ( .A(n29315), .B(n29316), .Z(N62793) );
  NANDN U38130 ( .A(n29317), .B(n29318), .Z(n29316) );
  OR U38131 ( .A(n29319), .B(n29320), .Z(n29318) );
  NAND U38132 ( .A(n29319), .B(n29320), .Z(n29315) );
  XOR U38133 ( .A(n29319), .B(n29321), .Z(N62792) );
  XNOR U38134 ( .A(n29317), .B(n29320), .Z(n29321) );
  AND U38135 ( .A(n29322), .B(n29323), .Z(n29320) );
  NANDN U38136 ( .A(n29324), .B(n29325), .Z(n29323) );
  NANDN U38137 ( .A(n29326), .B(n29327), .Z(n29325) );
  NANDN U38138 ( .A(n29327), .B(n29326), .Z(n29322) );
  NAND U38139 ( .A(n29328), .B(n29329), .Z(n29317) );
  NANDN U38140 ( .A(n29330), .B(n29331), .Z(n29329) );
  OR U38141 ( .A(n29332), .B(n29333), .Z(n29331) );
  NAND U38142 ( .A(n29333), .B(n29332), .Z(n29328) );
  AND U38143 ( .A(n29334), .B(n29335), .Z(n29319) );
  NANDN U38144 ( .A(n29336), .B(n29337), .Z(n29335) );
  NANDN U38145 ( .A(n29338), .B(n29339), .Z(n29337) );
  NANDN U38146 ( .A(n29339), .B(n29338), .Z(n29334) );
  XOR U38147 ( .A(n29333), .B(n29340), .Z(N62791) );
  XOR U38148 ( .A(n29330), .B(n29332), .Z(n29340) );
  XNOR U38149 ( .A(n29326), .B(n29341), .Z(n29332) );
  XNOR U38150 ( .A(n29324), .B(n29327), .Z(n29341) );
  NAND U38151 ( .A(n29342), .B(n29343), .Z(n29327) );
  NAND U38152 ( .A(n29344), .B(n29345), .Z(n29343) );
  OR U38153 ( .A(n29346), .B(n29347), .Z(n29344) );
  NANDN U38154 ( .A(n29348), .B(n29346), .Z(n29342) );
  IV U38155 ( .A(n29347), .Z(n29348) );
  NAND U38156 ( .A(n29349), .B(n29350), .Z(n29324) );
  NAND U38157 ( .A(n29351), .B(n29352), .Z(n29350) );
  NANDN U38158 ( .A(n29353), .B(n29354), .Z(n29351) );
  NANDN U38159 ( .A(n29354), .B(n29353), .Z(n29349) );
  AND U38160 ( .A(n29355), .B(n29356), .Z(n29326) );
  NAND U38161 ( .A(n29357), .B(n29358), .Z(n29356) );
  OR U38162 ( .A(n29359), .B(n29360), .Z(n29357) );
  NANDN U38163 ( .A(n29361), .B(n29359), .Z(n29355) );
  NAND U38164 ( .A(n29362), .B(n29363), .Z(n29330) );
  NANDN U38165 ( .A(n29364), .B(n29365), .Z(n29363) );
  OR U38166 ( .A(n29366), .B(n29367), .Z(n29365) );
  NANDN U38167 ( .A(n29368), .B(n29366), .Z(n29362) );
  IV U38168 ( .A(n29367), .Z(n29368) );
  XNOR U38169 ( .A(n29338), .B(n29369), .Z(n29333) );
  XNOR U38170 ( .A(n29336), .B(n29339), .Z(n29369) );
  NAND U38171 ( .A(n29370), .B(n29371), .Z(n29339) );
  NAND U38172 ( .A(n29372), .B(n29373), .Z(n29371) );
  OR U38173 ( .A(n29374), .B(n29375), .Z(n29372) );
  NANDN U38174 ( .A(n29376), .B(n29374), .Z(n29370) );
  IV U38175 ( .A(n29375), .Z(n29376) );
  NAND U38176 ( .A(n29377), .B(n29378), .Z(n29336) );
  NAND U38177 ( .A(n29379), .B(n29380), .Z(n29378) );
  NANDN U38178 ( .A(n29381), .B(n29382), .Z(n29379) );
  NANDN U38179 ( .A(n29382), .B(n29381), .Z(n29377) );
  AND U38180 ( .A(n29383), .B(n29384), .Z(n29338) );
  NAND U38181 ( .A(n29385), .B(n29386), .Z(n29384) );
  OR U38182 ( .A(n29387), .B(n29388), .Z(n29385) );
  NANDN U38183 ( .A(n29389), .B(n29387), .Z(n29383) );
  XNOR U38184 ( .A(n29364), .B(n29390), .Z(N62790) );
  XOR U38185 ( .A(n29366), .B(n29367), .Z(n29390) );
  XNOR U38186 ( .A(n29380), .B(n29391), .Z(n29367) );
  XOR U38187 ( .A(n29381), .B(n29382), .Z(n29391) );
  XOR U38188 ( .A(n29387), .B(n29392), .Z(n29382) );
  XOR U38189 ( .A(n29386), .B(n29389), .Z(n29392) );
  IV U38190 ( .A(n29388), .Z(n29389) );
  NAND U38191 ( .A(n29393), .B(n29394), .Z(n29388) );
  OR U38192 ( .A(n29395), .B(n29396), .Z(n29394) );
  OR U38193 ( .A(n29397), .B(n29398), .Z(n29393) );
  NAND U38194 ( .A(n29399), .B(n29400), .Z(n29386) );
  OR U38195 ( .A(n29401), .B(n29402), .Z(n29400) );
  OR U38196 ( .A(n29403), .B(n29404), .Z(n29399) );
  NOR U38197 ( .A(n29405), .B(n29406), .Z(n29387) );
  ANDN U38198 ( .B(n29407), .A(n29408), .Z(n29381) );
  XNOR U38199 ( .A(n29374), .B(n29409), .Z(n29380) );
  XNOR U38200 ( .A(n29373), .B(n29375), .Z(n29409) );
  NAND U38201 ( .A(n29410), .B(n29411), .Z(n29375) );
  OR U38202 ( .A(n29412), .B(n29413), .Z(n29411) );
  OR U38203 ( .A(n29414), .B(n29415), .Z(n29410) );
  NAND U38204 ( .A(n29416), .B(n29417), .Z(n29373) );
  OR U38205 ( .A(n29418), .B(n29419), .Z(n29417) );
  OR U38206 ( .A(n29420), .B(n29421), .Z(n29416) );
  ANDN U38207 ( .B(n29422), .A(n29423), .Z(n29374) );
  IV U38208 ( .A(n29424), .Z(n29422) );
  ANDN U38209 ( .B(n29425), .A(n29426), .Z(n29366) );
  XOR U38210 ( .A(n29352), .B(n29427), .Z(n29364) );
  XOR U38211 ( .A(n29353), .B(n29354), .Z(n29427) );
  XOR U38212 ( .A(n29359), .B(n29428), .Z(n29354) );
  XOR U38213 ( .A(n29358), .B(n29361), .Z(n29428) );
  IV U38214 ( .A(n29360), .Z(n29361) );
  NAND U38215 ( .A(n29429), .B(n29430), .Z(n29360) );
  OR U38216 ( .A(n29431), .B(n29432), .Z(n29430) );
  OR U38217 ( .A(n29433), .B(n29434), .Z(n29429) );
  NAND U38218 ( .A(n29435), .B(n29436), .Z(n29358) );
  OR U38219 ( .A(n29437), .B(n29438), .Z(n29436) );
  OR U38220 ( .A(n29439), .B(n29440), .Z(n29435) );
  NOR U38221 ( .A(n29441), .B(n29442), .Z(n29359) );
  ANDN U38222 ( .B(n29443), .A(n29444), .Z(n29353) );
  IV U38223 ( .A(n29445), .Z(n29443) );
  XNOR U38224 ( .A(n29346), .B(n29446), .Z(n29352) );
  XNOR U38225 ( .A(n29345), .B(n29347), .Z(n29446) );
  NAND U38226 ( .A(n29447), .B(n29448), .Z(n29347) );
  OR U38227 ( .A(n29449), .B(n29450), .Z(n29448) );
  OR U38228 ( .A(n29451), .B(n29452), .Z(n29447) );
  NAND U38229 ( .A(n29453), .B(n29454), .Z(n29345) );
  OR U38230 ( .A(n29455), .B(n29456), .Z(n29454) );
  OR U38231 ( .A(n29457), .B(n29458), .Z(n29453) );
  ANDN U38232 ( .B(n29459), .A(n29460), .Z(n29346) );
  IV U38233 ( .A(n29461), .Z(n29459) );
  XNOR U38234 ( .A(n29426), .B(n29425), .Z(N62789) );
  XOR U38235 ( .A(n29445), .B(n29444), .Z(n29425) );
  XNOR U38236 ( .A(n29460), .B(n29461), .Z(n29444) );
  XNOR U38237 ( .A(n29455), .B(n29456), .Z(n29461) );
  XNOR U38238 ( .A(n29457), .B(n29458), .Z(n29456) );
  XNOR U38239 ( .A(y[4069]), .B(x[4069]), .Z(n29458) );
  XNOR U38240 ( .A(y[4070]), .B(x[4070]), .Z(n29457) );
  XNOR U38241 ( .A(y[4068]), .B(x[4068]), .Z(n29455) );
  XNOR U38242 ( .A(n29449), .B(n29450), .Z(n29460) );
  XNOR U38243 ( .A(y[4065]), .B(x[4065]), .Z(n29450) );
  XNOR U38244 ( .A(n29451), .B(n29452), .Z(n29449) );
  XNOR U38245 ( .A(y[4066]), .B(x[4066]), .Z(n29452) );
  XNOR U38246 ( .A(y[4067]), .B(x[4067]), .Z(n29451) );
  XNOR U38247 ( .A(n29442), .B(n29441), .Z(n29445) );
  XNOR U38248 ( .A(n29437), .B(n29438), .Z(n29441) );
  XNOR U38249 ( .A(y[4062]), .B(x[4062]), .Z(n29438) );
  XNOR U38250 ( .A(n29439), .B(n29440), .Z(n29437) );
  XNOR U38251 ( .A(y[4063]), .B(x[4063]), .Z(n29440) );
  XNOR U38252 ( .A(y[4064]), .B(x[4064]), .Z(n29439) );
  XNOR U38253 ( .A(n29431), .B(n29432), .Z(n29442) );
  XNOR U38254 ( .A(y[4059]), .B(x[4059]), .Z(n29432) );
  XNOR U38255 ( .A(n29433), .B(n29434), .Z(n29431) );
  XNOR U38256 ( .A(y[4060]), .B(x[4060]), .Z(n29434) );
  XNOR U38257 ( .A(y[4061]), .B(x[4061]), .Z(n29433) );
  XOR U38258 ( .A(n29407), .B(n29408), .Z(n29426) );
  XNOR U38259 ( .A(n29423), .B(n29424), .Z(n29408) );
  XNOR U38260 ( .A(n29418), .B(n29419), .Z(n29424) );
  XNOR U38261 ( .A(n29420), .B(n29421), .Z(n29419) );
  XNOR U38262 ( .A(y[4057]), .B(x[4057]), .Z(n29421) );
  XNOR U38263 ( .A(y[4058]), .B(x[4058]), .Z(n29420) );
  XNOR U38264 ( .A(y[4056]), .B(x[4056]), .Z(n29418) );
  XNOR U38265 ( .A(n29412), .B(n29413), .Z(n29423) );
  XNOR U38266 ( .A(y[4053]), .B(x[4053]), .Z(n29413) );
  XNOR U38267 ( .A(n29414), .B(n29415), .Z(n29412) );
  XNOR U38268 ( .A(y[4054]), .B(x[4054]), .Z(n29415) );
  XNOR U38269 ( .A(y[4055]), .B(x[4055]), .Z(n29414) );
  XOR U38270 ( .A(n29406), .B(n29405), .Z(n29407) );
  XNOR U38271 ( .A(n29401), .B(n29402), .Z(n29405) );
  XNOR U38272 ( .A(y[4050]), .B(x[4050]), .Z(n29402) );
  XNOR U38273 ( .A(n29403), .B(n29404), .Z(n29401) );
  XNOR U38274 ( .A(y[4051]), .B(x[4051]), .Z(n29404) );
  XNOR U38275 ( .A(y[4052]), .B(x[4052]), .Z(n29403) );
  XNOR U38276 ( .A(n29395), .B(n29396), .Z(n29406) );
  XNOR U38277 ( .A(y[4047]), .B(x[4047]), .Z(n29396) );
  XNOR U38278 ( .A(n29397), .B(n29398), .Z(n29395) );
  XNOR U38279 ( .A(y[4048]), .B(x[4048]), .Z(n29398) );
  XNOR U38280 ( .A(y[4049]), .B(x[4049]), .Z(n29397) );
  NAND U38281 ( .A(n29462), .B(n29463), .Z(N62780) );
  NANDN U38282 ( .A(n29464), .B(n29465), .Z(n29463) );
  OR U38283 ( .A(n29466), .B(n29467), .Z(n29465) );
  NAND U38284 ( .A(n29466), .B(n29467), .Z(n29462) );
  XOR U38285 ( .A(n29466), .B(n29468), .Z(N62779) );
  XNOR U38286 ( .A(n29464), .B(n29467), .Z(n29468) );
  AND U38287 ( .A(n29469), .B(n29470), .Z(n29467) );
  NANDN U38288 ( .A(n29471), .B(n29472), .Z(n29470) );
  NANDN U38289 ( .A(n29473), .B(n29474), .Z(n29472) );
  NANDN U38290 ( .A(n29474), .B(n29473), .Z(n29469) );
  NAND U38291 ( .A(n29475), .B(n29476), .Z(n29464) );
  NANDN U38292 ( .A(n29477), .B(n29478), .Z(n29476) );
  OR U38293 ( .A(n29479), .B(n29480), .Z(n29478) );
  NAND U38294 ( .A(n29480), .B(n29479), .Z(n29475) );
  AND U38295 ( .A(n29481), .B(n29482), .Z(n29466) );
  NANDN U38296 ( .A(n29483), .B(n29484), .Z(n29482) );
  NANDN U38297 ( .A(n29485), .B(n29486), .Z(n29484) );
  NANDN U38298 ( .A(n29486), .B(n29485), .Z(n29481) );
  XOR U38299 ( .A(n29480), .B(n29487), .Z(N62778) );
  XOR U38300 ( .A(n29477), .B(n29479), .Z(n29487) );
  XNOR U38301 ( .A(n29473), .B(n29488), .Z(n29479) );
  XNOR U38302 ( .A(n29471), .B(n29474), .Z(n29488) );
  NAND U38303 ( .A(n29489), .B(n29490), .Z(n29474) );
  NAND U38304 ( .A(n29491), .B(n29492), .Z(n29490) );
  OR U38305 ( .A(n29493), .B(n29494), .Z(n29491) );
  NANDN U38306 ( .A(n29495), .B(n29493), .Z(n29489) );
  IV U38307 ( .A(n29494), .Z(n29495) );
  NAND U38308 ( .A(n29496), .B(n29497), .Z(n29471) );
  NAND U38309 ( .A(n29498), .B(n29499), .Z(n29497) );
  NANDN U38310 ( .A(n29500), .B(n29501), .Z(n29498) );
  NANDN U38311 ( .A(n29501), .B(n29500), .Z(n29496) );
  AND U38312 ( .A(n29502), .B(n29503), .Z(n29473) );
  NAND U38313 ( .A(n29504), .B(n29505), .Z(n29503) );
  OR U38314 ( .A(n29506), .B(n29507), .Z(n29504) );
  NANDN U38315 ( .A(n29508), .B(n29506), .Z(n29502) );
  NAND U38316 ( .A(n29509), .B(n29510), .Z(n29477) );
  NANDN U38317 ( .A(n29511), .B(n29512), .Z(n29510) );
  OR U38318 ( .A(n29513), .B(n29514), .Z(n29512) );
  NANDN U38319 ( .A(n29515), .B(n29513), .Z(n29509) );
  IV U38320 ( .A(n29514), .Z(n29515) );
  XNOR U38321 ( .A(n29485), .B(n29516), .Z(n29480) );
  XNOR U38322 ( .A(n29483), .B(n29486), .Z(n29516) );
  NAND U38323 ( .A(n29517), .B(n29518), .Z(n29486) );
  NAND U38324 ( .A(n29519), .B(n29520), .Z(n29518) );
  OR U38325 ( .A(n29521), .B(n29522), .Z(n29519) );
  NANDN U38326 ( .A(n29523), .B(n29521), .Z(n29517) );
  IV U38327 ( .A(n29522), .Z(n29523) );
  NAND U38328 ( .A(n29524), .B(n29525), .Z(n29483) );
  NAND U38329 ( .A(n29526), .B(n29527), .Z(n29525) );
  NANDN U38330 ( .A(n29528), .B(n29529), .Z(n29526) );
  NANDN U38331 ( .A(n29529), .B(n29528), .Z(n29524) );
  AND U38332 ( .A(n29530), .B(n29531), .Z(n29485) );
  NAND U38333 ( .A(n29532), .B(n29533), .Z(n29531) );
  OR U38334 ( .A(n29534), .B(n29535), .Z(n29532) );
  NANDN U38335 ( .A(n29536), .B(n29534), .Z(n29530) );
  XNOR U38336 ( .A(n29511), .B(n29537), .Z(N62777) );
  XOR U38337 ( .A(n29513), .B(n29514), .Z(n29537) );
  XNOR U38338 ( .A(n29527), .B(n29538), .Z(n29514) );
  XOR U38339 ( .A(n29528), .B(n29529), .Z(n29538) );
  XOR U38340 ( .A(n29534), .B(n29539), .Z(n29529) );
  XOR U38341 ( .A(n29533), .B(n29536), .Z(n29539) );
  IV U38342 ( .A(n29535), .Z(n29536) );
  NAND U38343 ( .A(n29540), .B(n29541), .Z(n29535) );
  OR U38344 ( .A(n29542), .B(n29543), .Z(n29541) );
  OR U38345 ( .A(n29544), .B(n29545), .Z(n29540) );
  NAND U38346 ( .A(n29546), .B(n29547), .Z(n29533) );
  OR U38347 ( .A(n29548), .B(n29549), .Z(n29547) );
  OR U38348 ( .A(n29550), .B(n29551), .Z(n29546) );
  NOR U38349 ( .A(n29552), .B(n29553), .Z(n29534) );
  ANDN U38350 ( .B(n29554), .A(n29555), .Z(n29528) );
  XNOR U38351 ( .A(n29521), .B(n29556), .Z(n29527) );
  XNOR U38352 ( .A(n29520), .B(n29522), .Z(n29556) );
  NAND U38353 ( .A(n29557), .B(n29558), .Z(n29522) );
  OR U38354 ( .A(n29559), .B(n29560), .Z(n29558) );
  OR U38355 ( .A(n29561), .B(n29562), .Z(n29557) );
  NAND U38356 ( .A(n29563), .B(n29564), .Z(n29520) );
  OR U38357 ( .A(n29565), .B(n29566), .Z(n29564) );
  OR U38358 ( .A(n29567), .B(n29568), .Z(n29563) );
  ANDN U38359 ( .B(n29569), .A(n29570), .Z(n29521) );
  IV U38360 ( .A(n29571), .Z(n29569) );
  ANDN U38361 ( .B(n29572), .A(n29573), .Z(n29513) );
  XOR U38362 ( .A(n29499), .B(n29574), .Z(n29511) );
  XOR U38363 ( .A(n29500), .B(n29501), .Z(n29574) );
  XOR U38364 ( .A(n29506), .B(n29575), .Z(n29501) );
  XOR U38365 ( .A(n29505), .B(n29508), .Z(n29575) );
  IV U38366 ( .A(n29507), .Z(n29508) );
  NAND U38367 ( .A(n29576), .B(n29577), .Z(n29507) );
  OR U38368 ( .A(n29578), .B(n29579), .Z(n29577) );
  OR U38369 ( .A(n29580), .B(n29581), .Z(n29576) );
  NAND U38370 ( .A(n29582), .B(n29583), .Z(n29505) );
  OR U38371 ( .A(n29584), .B(n29585), .Z(n29583) );
  OR U38372 ( .A(n29586), .B(n29587), .Z(n29582) );
  NOR U38373 ( .A(n29588), .B(n29589), .Z(n29506) );
  ANDN U38374 ( .B(n29590), .A(n29591), .Z(n29500) );
  IV U38375 ( .A(n29592), .Z(n29590) );
  XNOR U38376 ( .A(n29493), .B(n29593), .Z(n29499) );
  XNOR U38377 ( .A(n29492), .B(n29494), .Z(n29593) );
  NAND U38378 ( .A(n29594), .B(n29595), .Z(n29494) );
  OR U38379 ( .A(n29596), .B(n29597), .Z(n29595) );
  OR U38380 ( .A(n29598), .B(n29599), .Z(n29594) );
  NAND U38381 ( .A(n29600), .B(n29601), .Z(n29492) );
  OR U38382 ( .A(n29602), .B(n29603), .Z(n29601) );
  OR U38383 ( .A(n29604), .B(n29605), .Z(n29600) );
  ANDN U38384 ( .B(n29606), .A(n29607), .Z(n29493) );
  IV U38385 ( .A(n29608), .Z(n29606) );
  XNOR U38386 ( .A(n29573), .B(n29572), .Z(N62776) );
  XOR U38387 ( .A(n29592), .B(n29591), .Z(n29572) );
  XNOR U38388 ( .A(n29607), .B(n29608), .Z(n29591) );
  XNOR U38389 ( .A(n29602), .B(n29603), .Z(n29608) );
  XNOR U38390 ( .A(n29604), .B(n29605), .Z(n29603) );
  XNOR U38391 ( .A(y[4045]), .B(x[4045]), .Z(n29605) );
  XNOR U38392 ( .A(y[4046]), .B(x[4046]), .Z(n29604) );
  XNOR U38393 ( .A(y[4044]), .B(x[4044]), .Z(n29602) );
  XNOR U38394 ( .A(n29596), .B(n29597), .Z(n29607) );
  XNOR U38395 ( .A(y[4041]), .B(x[4041]), .Z(n29597) );
  XNOR U38396 ( .A(n29598), .B(n29599), .Z(n29596) );
  XNOR U38397 ( .A(y[4042]), .B(x[4042]), .Z(n29599) );
  XNOR U38398 ( .A(y[4043]), .B(x[4043]), .Z(n29598) );
  XNOR U38399 ( .A(n29589), .B(n29588), .Z(n29592) );
  XNOR U38400 ( .A(n29584), .B(n29585), .Z(n29588) );
  XNOR U38401 ( .A(y[4038]), .B(x[4038]), .Z(n29585) );
  XNOR U38402 ( .A(n29586), .B(n29587), .Z(n29584) );
  XNOR U38403 ( .A(y[4039]), .B(x[4039]), .Z(n29587) );
  XNOR U38404 ( .A(y[4040]), .B(x[4040]), .Z(n29586) );
  XNOR U38405 ( .A(n29578), .B(n29579), .Z(n29589) );
  XNOR U38406 ( .A(y[4035]), .B(x[4035]), .Z(n29579) );
  XNOR U38407 ( .A(n29580), .B(n29581), .Z(n29578) );
  XNOR U38408 ( .A(y[4036]), .B(x[4036]), .Z(n29581) );
  XNOR U38409 ( .A(y[4037]), .B(x[4037]), .Z(n29580) );
  XOR U38410 ( .A(n29554), .B(n29555), .Z(n29573) );
  XNOR U38411 ( .A(n29570), .B(n29571), .Z(n29555) );
  XNOR U38412 ( .A(n29565), .B(n29566), .Z(n29571) );
  XNOR U38413 ( .A(n29567), .B(n29568), .Z(n29566) );
  XNOR U38414 ( .A(y[4033]), .B(x[4033]), .Z(n29568) );
  XNOR U38415 ( .A(y[4034]), .B(x[4034]), .Z(n29567) );
  XNOR U38416 ( .A(y[4032]), .B(x[4032]), .Z(n29565) );
  XNOR U38417 ( .A(n29559), .B(n29560), .Z(n29570) );
  XNOR U38418 ( .A(y[4029]), .B(x[4029]), .Z(n29560) );
  XNOR U38419 ( .A(n29561), .B(n29562), .Z(n29559) );
  XNOR U38420 ( .A(y[4030]), .B(x[4030]), .Z(n29562) );
  XNOR U38421 ( .A(y[4031]), .B(x[4031]), .Z(n29561) );
  XOR U38422 ( .A(n29553), .B(n29552), .Z(n29554) );
  XNOR U38423 ( .A(n29548), .B(n29549), .Z(n29552) );
  XNOR U38424 ( .A(y[4026]), .B(x[4026]), .Z(n29549) );
  XNOR U38425 ( .A(n29550), .B(n29551), .Z(n29548) );
  XNOR U38426 ( .A(y[4027]), .B(x[4027]), .Z(n29551) );
  XNOR U38427 ( .A(y[4028]), .B(x[4028]), .Z(n29550) );
  XNOR U38428 ( .A(n29542), .B(n29543), .Z(n29553) );
  XNOR U38429 ( .A(y[4023]), .B(x[4023]), .Z(n29543) );
  XNOR U38430 ( .A(n29544), .B(n29545), .Z(n29542) );
  XNOR U38431 ( .A(y[4024]), .B(x[4024]), .Z(n29545) );
  XNOR U38432 ( .A(y[4025]), .B(x[4025]), .Z(n29544) );
  NAND U38433 ( .A(n29609), .B(n29610), .Z(N62767) );
  NANDN U38434 ( .A(n29611), .B(n29612), .Z(n29610) );
  OR U38435 ( .A(n29613), .B(n29614), .Z(n29612) );
  NAND U38436 ( .A(n29613), .B(n29614), .Z(n29609) );
  XOR U38437 ( .A(n29613), .B(n29615), .Z(N62766) );
  XNOR U38438 ( .A(n29611), .B(n29614), .Z(n29615) );
  AND U38439 ( .A(n29616), .B(n29617), .Z(n29614) );
  NANDN U38440 ( .A(n29618), .B(n29619), .Z(n29617) );
  NANDN U38441 ( .A(n29620), .B(n29621), .Z(n29619) );
  NANDN U38442 ( .A(n29621), .B(n29620), .Z(n29616) );
  NAND U38443 ( .A(n29622), .B(n29623), .Z(n29611) );
  NANDN U38444 ( .A(n29624), .B(n29625), .Z(n29623) );
  OR U38445 ( .A(n29626), .B(n29627), .Z(n29625) );
  NAND U38446 ( .A(n29627), .B(n29626), .Z(n29622) );
  AND U38447 ( .A(n29628), .B(n29629), .Z(n29613) );
  NANDN U38448 ( .A(n29630), .B(n29631), .Z(n29629) );
  NANDN U38449 ( .A(n29632), .B(n29633), .Z(n29631) );
  NANDN U38450 ( .A(n29633), .B(n29632), .Z(n29628) );
  XOR U38451 ( .A(n29627), .B(n29634), .Z(N62765) );
  XOR U38452 ( .A(n29624), .B(n29626), .Z(n29634) );
  XNOR U38453 ( .A(n29620), .B(n29635), .Z(n29626) );
  XNOR U38454 ( .A(n29618), .B(n29621), .Z(n29635) );
  NAND U38455 ( .A(n29636), .B(n29637), .Z(n29621) );
  NAND U38456 ( .A(n29638), .B(n29639), .Z(n29637) );
  OR U38457 ( .A(n29640), .B(n29641), .Z(n29638) );
  NANDN U38458 ( .A(n29642), .B(n29640), .Z(n29636) );
  IV U38459 ( .A(n29641), .Z(n29642) );
  NAND U38460 ( .A(n29643), .B(n29644), .Z(n29618) );
  NAND U38461 ( .A(n29645), .B(n29646), .Z(n29644) );
  NANDN U38462 ( .A(n29647), .B(n29648), .Z(n29645) );
  NANDN U38463 ( .A(n29648), .B(n29647), .Z(n29643) );
  AND U38464 ( .A(n29649), .B(n29650), .Z(n29620) );
  NAND U38465 ( .A(n29651), .B(n29652), .Z(n29650) );
  OR U38466 ( .A(n29653), .B(n29654), .Z(n29651) );
  NANDN U38467 ( .A(n29655), .B(n29653), .Z(n29649) );
  NAND U38468 ( .A(n29656), .B(n29657), .Z(n29624) );
  NANDN U38469 ( .A(n29658), .B(n29659), .Z(n29657) );
  OR U38470 ( .A(n29660), .B(n29661), .Z(n29659) );
  NANDN U38471 ( .A(n29662), .B(n29660), .Z(n29656) );
  IV U38472 ( .A(n29661), .Z(n29662) );
  XNOR U38473 ( .A(n29632), .B(n29663), .Z(n29627) );
  XNOR U38474 ( .A(n29630), .B(n29633), .Z(n29663) );
  NAND U38475 ( .A(n29664), .B(n29665), .Z(n29633) );
  NAND U38476 ( .A(n29666), .B(n29667), .Z(n29665) );
  OR U38477 ( .A(n29668), .B(n29669), .Z(n29666) );
  NANDN U38478 ( .A(n29670), .B(n29668), .Z(n29664) );
  IV U38479 ( .A(n29669), .Z(n29670) );
  NAND U38480 ( .A(n29671), .B(n29672), .Z(n29630) );
  NAND U38481 ( .A(n29673), .B(n29674), .Z(n29672) );
  NANDN U38482 ( .A(n29675), .B(n29676), .Z(n29673) );
  NANDN U38483 ( .A(n29676), .B(n29675), .Z(n29671) );
  AND U38484 ( .A(n29677), .B(n29678), .Z(n29632) );
  NAND U38485 ( .A(n29679), .B(n29680), .Z(n29678) );
  OR U38486 ( .A(n29681), .B(n29682), .Z(n29679) );
  NANDN U38487 ( .A(n29683), .B(n29681), .Z(n29677) );
  XNOR U38488 ( .A(n29658), .B(n29684), .Z(N62764) );
  XOR U38489 ( .A(n29660), .B(n29661), .Z(n29684) );
  XNOR U38490 ( .A(n29674), .B(n29685), .Z(n29661) );
  XOR U38491 ( .A(n29675), .B(n29676), .Z(n29685) );
  XOR U38492 ( .A(n29681), .B(n29686), .Z(n29676) );
  XOR U38493 ( .A(n29680), .B(n29683), .Z(n29686) );
  IV U38494 ( .A(n29682), .Z(n29683) );
  NAND U38495 ( .A(n29687), .B(n29688), .Z(n29682) );
  OR U38496 ( .A(n29689), .B(n29690), .Z(n29688) );
  OR U38497 ( .A(n29691), .B(n29692), .Z(n29687) );
  NAND U38498 ( .A(n29693), .B(n29694), .Z(n29680) );
  OR U38499 ( .A(n29695), .B(n29696), .Z(n29694) );
  OR U38500 ( .A(n29697), .B(n29698), .Z(n29693) );
  NOR U38501 ( .A(n29699), .B(n29700), .Z(n29681) );
  ANDN U38502 ( .B(n29701), .A(n29702), .Z(n29675) );
  XNOR U38503 ( .A(n29668), .B(n29703), .Z(n29674) );
  XNOR U38504 ( .A(n29667), .B(n29669), .Z(n29703) );
  NAND U38505 ( .A(n29704), .B(n29705), .Z(n29669) );
  OR U38506 ( .A(n29706), .B(n29707), .Z(n29705) );
  OR U38507 ( .A(n29708), .B(n29709), .Z(n29704) );
  NAND U38508 ( .A(n29710), .B(n29711), .Z(n29667) );
  OR U38509 ( .A(n29712), .B(n29713), .Z(n29711) );
  OR U38510 ( .A(n29714), .B(n29715), .Z(n29710) );
  ANDN U38511 ( .B(n29716), .A(n29717), .Z(n29668) );
  IV U38512 ( .A(n29718), .Z(n29716) );
  ANDN U38513 ( .B(n29719), .A(n29720), .Z(n29660) );
  XOR U38514 ( .A(n29646), .B(n29721), .Z(n29658) );
  XOR U38515 ( .A(n29647), .B(n29648), .Z(n29721) );
  XOR U38516 ( .A(n29653), .B(n29722), .Z(n29648) );
  XOR U38517 ( .A(n29652), .B(n29655), .Z(n29722) );
  IV U38518 ( .A(n29654), .Z(n29655) );
  NAND U38519 ( .A(n29723), .B(n29724), .Z(n29654) );
  OR U38520 ( .A(n29725), .B(n29726), .Z(n29724) );
  OR U38521 ( .A(n29727), .B(n29728), .Z(n29723) );
  NAND U38522 ( .A(n29729), .B(n29730), .Z(n29652) );
  OR U38523 ( .A(n29731), .B(n29732), .Z(n29730) );
  OR U38524 ( .A(n29733), .B(n29734), .Z(n29729) );
  NOR U38525 ( .A(n29735), .B(n29736), .Z(n29653) );
  ANDN U38526 ( .B(n29737), .A(n29738), .Z(n29647) );
  IV U38527 ( .A(n29739), .Z(n29737) );
  XNOR U38528 ( .A(n29640), .B(n29740), .Z(n29646) );
  XNOR U38529 ( .A(n29639), .B(n29641), .Z(n29740) );
  NAND U38530 ( .A(n29741), .B(n29742), .Z(n29641) );
  OR U38531 ( .A(n29743), .B(n29744), .Z(n29742) );
  OR U38532 ( .A(n29745), .B(n29746), .Z(n29741) );
  NAND U38533 ( .A(n29747), .B(n29748), .Z(n29639) );
  OR U38534 ( .A(n29749), .B(n29750), .Z(n29748) );
  OR U38535 ( .A(n29751), .B(n29752), .Z(n29747) );
  ANDN U38536 ( .B(n29753), .A(n29754), .Z(n29640) );
  IV U38537 ( .A(n29755), .Z(n29753) );
  XNOR U38538 ( .A(n29720), .B(n29719), .Z(N62763) );
  XOR U38539 ( .A(n29739), .B(n29738), .Z(n29719) );
  XNOR U38540 ( .A(n29754), .B(n29755), .Z(n29738) );
  XNOR U38541 ( .A(n29749), .B(n29750), .Z(n29755) );
  XNOR U38542 ( .A(n29751), .B(n29752), .Z(n29750) );
  XNOR U38543 ( .A(y[4021]), .B(x[4021]), .Z(n29752) );
  XNOR U38544 ( .A(y[4022]), .B(x[4022]), .Z(n29751) );
  XNOR U38545 ( .A(y[4020]), .B(x[4020]), .Z(n29749) );
  XNOR U38546 ( .A(n29743), .B(n29744), .Z(n29754) );
  XNOR U38547 ( .A(y[4017]), .B(x[4017]), .Z(n29744) );
  XNOR U38548 ( .A(n29745), .B(n29746), .Z(n29743) );
  XNOR U38549 ( .A(y[4018]), .B(x[4018]), .Z(n29746) );
  XNOR U38550 ( .A(y[4019]), .B(x[4019]), .Z(n29745) );
  XNOR U38551 ( .A(n29736), .B(n29735), .Z(n29739) );
  XNOR U38552 ( .A(n29731), .B(n29732), .Z(n29735) );
  XNOR U38553 ( .A(y[4014]), .B(x[4014]), .Z(n29732) );
  XNOR U38554 ( .A(n29733), .B(n29734), .Z(n29731) );
  XNOR U38555 ( .A(y[4015]), .B(x[4015]), .Z(n29734) );
  XNOR U38556 ( .A(y[4016]), .B(x[4016]), .Z(n29733) );
  XNOR U38557 ( .A(n29725), .B(n29726), .Z(n29736) );
  XNOR U38558 ( .A(y[4011]), .B(x[4011]), .Z(n29726) );
  XNOR U38559 ( .A(n29727), .B(n29728), .Z(n29725) );
  XNOR U38560 ( .A(y[4012]), .B(x[4012]), .Z(n29728) );
  XNOR U38561 ( .A(y[4013]), .B(x[4013]), .Z(n29727) );
  XOR U38562 ( .A(n29701), .B(n29702), .Z(n29720) );
  XNOR U38563 ( .A(n29717), .B(n29718), .Z(n29702) );
  XNOR U38564 ( .A(n29712), .B(n29713), .Z(n29718) );
  XNOR U38565 ( .A(n29714), .B(n29715), .Z(n29713) );
  XNOR U38566 ( .A(y[4009]), .B(x[4009]), .Z(n29715) );
  XNOR U38567 ( .A(y[4010]), .B(x[4010]), .Z(n29714) );
  XNOR U38568 ( .A(y[4008]), .B(x[4008]), .Z(n29712) );
  XNOR U38569 ( .A(n29706), .B(n29707), .Z(n29717) );
  XNOR U38570 ( .A(y[4005]), .B(x[4005]), .Z(n29707) );
  XNOR U38571 ( .A(n29708), .B(n29709), .Z(n29706) );
  XNOR U38572 ( .A(y[4006]), .B(x[4006]), .Z(n29709) );
  XNOR U38573 ( .A(y[4007]), .B(x[4007]), .Z(n29708) );
  XOR U38574 ( .A(n29700), .B(n29699), .Z(n29701) );
  XNOR U38575 ( .A(n29695), .B(n29696), .Z(n29699) );
  XNOR U38576 ( .A(y[4002]), .B(x[4002]), .Z(n29696) );
  XNOR U38577 ( .A(n29697), .B(n29698), .Z(n29695) );
  XNOR U38578 ( .A(y[4003]), .B(x[4003]), .Z(n29698) );
  XNOR U38579 ( .A(y[4004]), .B(x[4004]), .Z(n29697) );
  XNOR U38580 ( .A(n29689), .B(n29690), .Z(n29700) );
  XNOR U38581 ( .A(y[3999]), .B(x[3999]), .Z(n29690) );
  XNOR U38582 ( .A(n29691), .B(n29692), .Z(n29689) );
  XNOR U38583 ( .A(y[4000]), .B(x[4000]), .Z(n29692) );
  XNOR U38584 ( .A(y[4001]), .B(x[4001]), .Z(n29691) );
  NAND U38585 ( .A(n29756), .B(n29757), .Z(N62754) );
  NANDN U38586 ( .A(n29758), .B(n29759), .Z(n29757) );
  OR U38587 ( .A(n29760), .B(n29761), .Z(n29759) );
  NAND U38588 ( .A(n29760), .B(n29761), .Z(n29756) );
  XOR U38589 ( .A(n29760), .B(n29762), .Z(N62753) );
  XNOR U38590 ( .A(n29758), .B(n29761), .Z(n29762) );
  AND U38591 ( .A(n29763), .B(n29764), .Z(n29761) );
  NANDN U38592 ( .A(n29765), .B(n29766), .Z(n29764) );
  NANDN U38593 ( .A(n29767), .B(n29768), .Z(n29766) );
  NANDN U38594 ( .A(n29768), .B(n29767), .Z(n29763) );
  NAND U38595 ( .A(n29769), .B(n29770), .Z(n29758) );
  NANDN U38596 ( .A(n29771), .B(n29772), .Z(n29770) );
  OR U38597 ( .A(n29773), .B(n29774), .Z(n29772) );
  NAND U38598 ( .A(n29774), .B(n29773), .Z(n29769) );
  AND U38599 ( .A(n29775), .B(n29776), .Z(n29760) );
  NANDN U38600 ( .A(n29777), .B(n29778), .Z(n29776) );
  NANDN U38601 ( .A(n29779), .B(n29780), .Z(n29778) );
  NANDN U38602 ( .A(n29780), .B(n29779), .Z(n29775) );
  XOR U38603 ( .A(n29774), .B(n29781), .Z(N62752) );
  XOR U38604 ( .A(n29771), .B(n29773), .Z(n29781) );
  XNOR U38605 ( .A(n29767), .B(n29782), .Z(n29773) );
  XNOR U38606 ( .A(n29765), .B(n29768), .Z(n29782) );
  NAND U38607 ( .A(n29783), .B(n29784), .Z(n29768) );
  NAND U38608 ( .A(n29785), .B(n29786), .Z(n29784) );
  OR U38609 ( .A(n29787), .B(n29788), .Z(n29785) );
  NANDN U38610 ( .A(n29789), .B(n29787), .Z(n29783) );
  IV U38611 ( .A(n29788), .Z(n29789) );
  NAND U38612 ( .A(n29790), .B(n29791), .Z(n29765) );
  NAND U38613 ( .A(n29792), .B(n29793), .Z(n29791) );
  NANDN U38614 ( .A(n29794), .B(n29795), .Z(n29792) );
  NANDN U38615 ( .A(n29795), .B(n29794), .Z(n29790) );
  AND U38616 ( .A(n29796), .B(n29797), .Z(n29767) );
  NAND U38617 ( .A(n29798), .B(n29799), .Z(n29797) );
  OR U38618 ( .A(n29800), .B(n29801), .Z(n29798) );
  NANDN U38619 ( .A(n29802), .B(n29800), .Z(n29796) );
  NAND U38620 ( .A(n29803), .B(n29804), .Z(n29771) );
  NANDN U38621 ( .A(n29805), .B(n29806), .Z(n29804) );
  OR U38622 ( .A(n29807), .B(n29808), .Z(n29806) );
  NANDN U38623 ( .A(n29809), .B(n29807), .Z(n29803) );
  IV U38624 ( .A(n29808), .Z(n29809) );
  XNOR U38625 ( .A(n29779), .B(n29810), .Z(n29774) );
  XNOR U38626 ( .A(n29777), .B(n29780), .Z(n29810) );
  NAND U38627 ( .A(n29811), .B(n29812), .Z(n29780) );
  NAND U38628 ( .A(n29813), .B(n29814), .Z(n29812) );
  OR U38629 ( .A(n29815), .B(n29816), .Z(n29813) );
  NANDN U38630 ( .A(n29817), .B(n29815), .Z(n29811) );
  IV U38631 ( .A(n29816), .Z(n29817) );
  NAND U38632 ( .A(n29818), .B(n29819), .Z(n29777) );
  NAND U38633 ( .A(n29820), .B(n29821), .Z(n29819) );
  NANDN U38634 ( .A(n29822), .B(n29823), .Z(n29820) );
  NANDN U38635 ( .A(n29823), .B(n29822), .Z(n29818) );
  AND U38636 ( .A(n29824), .B(n29825), .Z(n29779) );
  NAND U38637 ( .A(n29826), .B(n29827), .Z(n29825) );
  OR U38638 ( .A(n29828), .B(n29829), .Z(n29826) );
  NANDN U38639 ( .A(n29830), .B(n29828), .Z(n29824) );
  XNOR U38640 ( .A(n29805), .B(n29831), .Z(N62751) );
  XOR U38641 ( .A(n29807), .B(n29808), .Z(n29831) );
  XNOR U38642 ( .A(n29821), .B(n29832), .Z(n29808) );
  XOR U38643 ( .A(n29822), .B(n29823), .Z(n29832) );
  XOR U38644 ( .A(n29828), .B(n29833), .Z(n29823) );
  XOR U38645 ( .A(n29827), .B(n29830), .Z(n29833) );
  IV U38646 ( .A(n29829), .Z(n29830) );
  NAND U38647 ( .A(n29834), .B(n29835), .Z(n29829) );
  OR U38648 ( .A(n29836), .B(n29837), .Z(n29835) );
  OR U38649 ( .A(n29838), .B(n29839), .Z(n29834) );
  NAND U38650 ( .A(n29840), .B(n29841), .Z(n29827) );
  OR U38651 ( .A(n29842), .B(n29843), .Z(n29841) );
  OR U38652 ( .A(n29844), .B(n29845), .Z(n29840) );
  NOR U38653 ( .A(n29846), .B(n29847), .Z(n29828) );
  ANDN U38654 ( .B(n29848), .A(n29849), .Z(n29822) );
  XNOR U38655 ( .A(n29815), .B(n29850), .Z(n29821) );
  XNOR U38656 ( .A(n29814), .B(n29816), .Z(n29850) );
  NAND U38657 ( .A(n29851), .B(n29852), .Z(n29816) );
  OR U38658 ( .A(n29853), .B(n29854), .Z(n29852) );
  OR U38659 ( .A(n29855), .B(n29856), .Z(n29851) );
  NAND U38660 ( .A(n29857), .B(n29858), .Z(n29814) );
  OR U38661 ( .A(n29859), .B(n29860), .Z(n29858) );
  OR U38662 ( .A(n29861), .B(n29862), .Z(n29857) );
  ANDN U38663 ( .B(n29863), .A(n29864), .Z(n29815) );
  IV U38664 ( .A(n29865), .Z(n29863) );
  ANDN U38665 ( .B(n29866), .A(n29867), .Z(n29807) );
  XOR U38666 ( .A(n29793), .B(n29868), .Z(n29805) );
  XOR U38667 ( .A(n29794), .B(n29795), .Z(n29868) );
  XOR U38668 ( .A(n29800), .B(n29869), .Z(n29795) );
  XOR U38669 ( .A(n29799), .B(n29802), .Z(n29869) );
  IV U38670 ( .A(n29801), .Z(n29802) );
  NAND U38671 ( .A(n29870), .B(n29871), .Z(n29801) );
  OR U38672 ( .A(n29872), .B(n29873), .Z(n29871) );
  OR U38673 ( .A(n29874), .B(n29875), .Z(n29870) );
  NAND U38674 ( .A(n29876), .B(n29877), .Z(n29799) );
  OR U38675 ( .A(n29878), .B(n29879), .Z(n29877) );
  OR U38676 ( .A(n29880), .B(n29881), .Z(n29876) );
  NOR U38677 ( .A(n29882), .B(n29883), .Z(n29800) );
  ANDN U38678 ( .B(n29884), .A(n29885), .Z(n29794) );
  IV U38679 ( .A(n29886), .Z(n29884) );
  XNOR U38680 ( .A(n29787), .B(n29887), .Z(n29793) );
  XNOR U38681 ( .A(n29786), .B(n29788), .Z(n29887) );
  NAND U38682 ( .A(n29888), .B(n29889), .Z(n29788) );
  OR U38683 ( .A(n29890), .B(n29891), .Z(n29889) );
  OR U38684 ( .A(n29892), .B(n29893), .Z(n29888) );
  NAND U38685 ( .A(n29894), .B(n29895), .Z(n29786) );
  OR U38686 ( .A(n29896), .B(n29897), .Z(n29895) );
  OR U38687 ( .A(n29898), .B(n29899), .Z(n29894) );
  ANDN U38688 ( .B(n29900), .A(n29901), .Z(n29787) );
  IV U38689 ( .A(n29902), .Z(n29900) );
  XNOR U38690 ( .A(n29867), .B(n29866), .Z(N62750) );
  XOR U38691 ( .A(n29886), .B(n29885), .Z(n29866) );
  XNOR U38692 ( .A(n29901), .B(n29902), .Z(n29885) );
  XNOR U38693 ( .A(n29896), .B(n29897), .Z(n29902) );
  XNOR U38694 ( .A(n29898), .B(n29899), .Z(n29897) );
  XNOR U38695 ( .A(y[3997]), .B(x[3997]), .Z(n29899) );
  XNOR U38696 ( .A(y[3998]), .B(x[3998]), .Z(n29898) );
  XNOR U38697 ( .A(y[3996]), .B(x[3996]), .Z(n29896) );
  XNOR U38698 ( .A(n29890), .B(n29891), .Z(n29901) );
  XNOR U38699 ( .A(y[3993]), .B(x[3993]), .Z(n29891) );
  XNOR U38700 ( .A(n29892), .B(n29893), .Z(n29890) );
  XNOR U38701 ( .A(y[3994]), .B(x[3994]), .Z(n29893) );
  XNOR U38702 ( .A(y[3995]), .B(x[3995]), .Z(n29892) );
  XNOR U38703 ( .A(n29883), .B(n29882), .Z(n29886) );
  XNOR U38704 ( .A(n29878), .B(n29879), .Z(n29882) );
  XNOR U38705 ( .A(y[3990]), .B(x[3990]), .Z(n29879) );
  XNOR U38706 ( .A(n29880), .B(n29881), .Z(n29878) );
  XNOR U38707 ( .A(y[3991]), .B(x[3991]), .Z(n29881) );
  XNOR U38708 ( .A(y[3992]), .B(x[3992]), .Z(n29880) );
  XNOR U38709 ( .A(n29872), .B(n29873), .Z(n29883) );
  XNOR U38710 ( .A(y[3987]), .B(x[3987]), .Z(n29873) );
  XNOR U38711 ( .A(n29874), .B(n29875), .Z(n29872) );
  XNOR U38712 ( .A(y[3988]), .B(x[3988]), .Z(n29875) );
  XNOR U38713 ( .A(y[3989]), .B(x[3989]), .Z(n29874) );
  XOR U38714 ( .A(n29848), .B(n29849), .Z(n29867) );
  XNOR U38715 ( .A(n29864), .B(n29865), .Z(n29849) );
  XNOR U38716 ( .A(n29859), .B(n29860), .Z(n29865) );
  XNOR U38717 ( .A(n29861), .B(n29862), .Z(n29860) );
  XNOR U38718 ( .A(y[3985]), .B(x[3985]), .Z(n29862) );
  XNOR U38719 ( .A(y[3986]), .B(x[3986]), .Z(n29861) );
  XNOR U38720 ( .A(y[3984]), .B(x[3984]), .Z(n29859) );
  XNOR U38721 ( .A(n29853), .B(n29854), .Z(n29864) );
  XNOR U38722 ( .A(y[3981]), .B(x[3981]), .Z(n29854) );
  XNOR U38723 ( .A(n29855), .B(n29856), .Z(n29853) );
  XNOR U38724 ( .A(y[3982]), .B(x[3982]), .Z(n29856) );
  XNOR U38725 ( .A(y[3983]), .B(x[3983]), .Z(n29855) );
  XOR U38726 ( .A(n29847), .B(n29846), .Z(n29848) );
  XNOR U38727 ( .A(n29842), .B(n29843), .Z(n29846) );
  XNOR U38728 ( .A(y[3978]), .B(x[3978]), .Z(n29843) );
  XNOR U38729 ( .A(n29844), .B(n29845), .Z(n29842) );
  XNOR U38730 ( .A(y[3979]), .B(x[3979]), .Z(n29845) );
  XNOR U38731 ( .A(y[3980]), .B(x[3980]), .Z(n29844) );
  XNOR U38732 ( .A(n29836), .B(n29837), .Z(n29847) );
  XNOR U38733 ( .A(y[3975]), .B(x[3975]), .Z(n29837) );
  XNOR U38734 ( .A(n29838), .B(n29839), .Z(n29836) );
  XNOR U38735 ( .A(y[3976]), .B(x[3976]), .Z(n29839) );
  XNOR U38736 ( .A(y[3977]), .B(x[3977]), .Z(n29838) );
  NAND U38737 ( .A(n29903), .B(n29904), .Z(N62741) );
  NANDN U38738 ( .A(n29905), .B(n29906), .Z(n29904) );
  OR U38739 ( .A(n29907), .B(n29908), .Z(n29906) );
  NAND U38740 ( .A(n29907), .B(n29908), .Z(n29903) );
  XOR U38741 ( .A(n29907), .B(n29909), .Z(N62740) );
  XNOR U38742 ( .A(n29905), .B(n29908), .Z(n29909) );
  AND U38743 ( .A(n29910), .B(n29911), .Z(n29908) );
  NANDN U38744 ( .A(n29912), .B(n29913), .Z(n29911) );
  NANDN U38745 ( .A(n29914), .B(n29915), .Z(n29913) );
  NANDN U38746 ( .A(n29915), .B(n29914), .Z(n29910) );
  NAND U38747 ( .A(n29916), .B(n29917), .Z(n29905) );
  NANDN U38748 ( .A(n29918), .B(n29919), .Z(n29917) );
  OR U38749 ( .A(n29920), .B(n29921), .Z(n29919) );
  NAND U38750 ( .A(n29921), .B(n29920), .Z(n29916) );
  AND U38751 ( .A(n29922), .B(n29923), .Z(n29907) );
  NANDN U38752 ( .A(n29924), .B(n29925), .Z(n29923) );
  NANDN U38753 ( .A(n29926), .B(n29927), .Z(n29925) );
  NANDN U38754 ( .A(n29927), .B(n29926), .Z(n29922) );
  XOR U38755 ( .A(n29921), .B(n29928), .Z(N62739) );
  XOR U38756 ( .A(n29918), .B(n29920), .Z(n29928) );
  XNOR U38757 ( .A(n29914), .B(n29929), .Z(n29920) );
  XNOR U38758 ( .A(n29912), .B(n29915), .Z(n29929) );
  NAND U38759 ( .A(n29930), .B(n29931), .Z(n29915) );
  NAND U38760 ( .A(n29932), .B(n29933), .Z(n29931) );
  OR U38761 ( .A(n29934), .B(n29935), .Z(n29932) );
  NANDN U38762 ( .A(n29936), .B(n29934), .Z(n29930) );
  IV U38763 ( .A(n29935), .Z(n29936) );
  NAND U38764 ( .A(n29937), .B(n29938), .Z(n29912) );
  NAND U38765 ( .A(n29939), .B(n29940), .Z(n29938) );
  NANDN U38766 ( .A(n29941), .B(n29942), .Z(n29939) );
  NANDN U38767 ( .A(n29942), .B(n29941), .Z(n29937) );
  AND U38768 ( .A(n29943), .B(n29944), .Z(n29914) );
  NAND U38769 ( .A(n29945), .B(n29946), .Z(n29944) );
  OR U38770 ( .A(n29947), .B(n29948), .Z(n29945) );
  NANDN U38771 ( .A(n29949), .B(n29947), .Z(n29943) );
  NAND U38772 ( .A(n29950), .B(n29951), .Z(n29918) );
  NANDN U38773 ( .A(n29952), .B(n29953), .Z(n29951) );
  OR U38774 ( .A(n29954), .B(n29955), .Z(n29953) );
  NANDN U38775 ( .A(n29956), .B(n29954), .Z(n29950) );
  IV U38776 ( .A(n29955), .Z(n29956) );
  XNOR U38777 ( .A(n29926), .B(n29957), .Z(n29921) );
  XNOR U38778 ( .A(n29924), .B(n29927), .Z(n29957) );
  NAND U38779 ( .A(n29958), .B(n29959), .Z(n29927) );
  NAND U38780 ( .A(n29960), .B(n29961), .Z(n29959) );
  OR U38781 ( .A(n29962), .B(n29963), .Z(n29960) );
  NANDN U38782 ( .A(n29964), .B(n29962), .Z(n29958) );
  IV U38783 ( .A(n29963), .Z(n29964) );
  NAND U38784 ( .A(n29965), .B(n29966), .Z(n29924) );
  NAND U38785 ( .A(n29967), .B(n29968), .Z(n29966) );
  NANDN U38786 ( .A(n29969), .B(n29970), .Z(n29967) );
  NANDN U38787 ( .A(n29970), .B(n29969), .Z(n29965) );
  AND U38788 ( .A(n29971), .B(n29972), .Z(n29926) );
  NAND U38789 ( .A(n29973), .B(n29974), .Z(n29972) );
  OR U38790 ( .A(n29975), .B(n29976), .Z(n29973) );
  NANDN U38791 ( .A(n29977), .B(n29975), .Z(n29971) );
  XNOR U38792 ( .A(n29952), .B(n29978), .Z(N62738) );
  XOR U38793 ( .A(n29954), .B(n29955), .Z(n29978) );
  XNOR U38794 ( .A(n29968), .B(n29979), .Z(n29955) );
  XOR U38795 ( .A(n29969), .B(n29970), .Z(n29979) );
  XOR U38796 ( .A(n29975), .B(n29980), .Z(n29970) );
  XOR U38797 ( .A(n29974), .B(n29977), .Z(n29980) );
  IV U38798 ( .A(n29976), .Z(n29977) );
  NAND U38799 ( .A(n29981), .B(n29982), .Z(n29976) );
  OR U38800 ( .A(n29983), .B(n29984), .Z(n29982) );
  OR U38801 ( .A(n29985), .B(n29986), .Z(n29981) );
  NAND U38802 ( .A(n29987), .B(n29988), .Z(n29974) );
  OR U38803 ( .A(n29989), .B(n29990), .Z(n29988) );
  OR U38804 ( .A(n29991), .B(n29992), .Z(n29987) );
  NOR U38805 ( .A(n29993), .B(n29994), .Z(n29975) );
  ANDN U38806 ( .B(n29995), .A(n29996), .Z(n29969) );
  XNOR U38807 ( .A(n29962), .B(n29997), .Z(n29968) );
  XNOR U38808 ( .A(n29961), .B(n29963), .Z(n29997) );
  NAND U38809 ( .A(n29998), .B(n29999), .Z(n29963) );
  OR U38810 ( .A(n30000), .B(n30001), .Z(n29999) );
  OR U38811 ( .A(n30002), .B(n30003), .Z(n29998) );
  NAND U38812 ( .A(n30004), .B(n30005), .Z(n29961) );
  OR U38813 ( .A(n30006), .B(n30007), .Z(n30005) );
  OR U38814 ( .A(n30008), .B(n30009), .Z(n30004) );
  ANDN U38815 ( .B(n30010), .A(n30011), .Z(n29962) );
  IV U38816 ( .A(n30012), .Z(n30010) );
  ANDN U38817 ( .B(n30013), .A(n30014), .Z(n29954) );
  XOR U38818 ( .A(n29940), .B(n30015), .Z(n29952) );
  XOR U38819 ( .A(n29941), .B(n29942), .Z(n30015) );
  XOR U38820 ( .A(n29947), .B(n30016), .Z(n29942) );
  XOR U38821 ( .A(n29946), .B(n29949), .Z(n30016) );
  IV U38822 ( .A(n29948), .Z(n29949) );
  NAND U38823 ( .A(n30017), .B(n30018), .Z(n29948) );
  OR U38824 ( .A(n30019), .B(n30020), .Z(n30018) );
  OR U38825 ( .A(n30021), .B(n30022), .Z(n30017) );
  NAND U38826 ( .A(n30023), .B(n30024), .Z(n29946) );
  OR U38827 ( .A(n30025), .B(n30026), .Z(n30024) );
  OR U38828 ( .A(n30027), .B(n30028), .Z(n30023) );
  NOR U38829 ( .A(n30029), .B(n30030), .Z(n29947) );
  ANDN U38830 ( .B(n30031), .A(n30032), .Z(n29941) );
  IV U38831 ( .A(n30033), .Z(n30031) );
  XNOR U38832 ( .A(n29934), .B(n30034), .Z(n29940) );
  XNOR U38833 ( .A(n29933), .B(n29935), .Z(n30034) );
  NAND U38834 ( .A(n30035), .B(n30036), .Z(n29935) );
  OR U38835 ( .A(n30037), .B(n30038), .Z(n30036) );
  OR U38836 ( .A(n30039), .B(n30040), .Z(n30035) );
  NAND U38837 ( .A(n30041), .B(n30042), .Z(n29933) );
  OR U38838 ( .A(n30043), .B(n30044), .Z(n30042) );
  OR U38839 ( .A(n30045), .B(n30046), .Z(n30041) );
  ANDN U38840 ( .B(n30047), .A(n30048), .Z(n29934) );
  IV U38841 ( .A(n30049), .Z(n30047) );
  XNOR U38842 ( .A(n30014), .B(n30013), .Z(N62737) );
  XOR U38843 ( .A(n30033), .B(n30032), .Z(n30013) );
  XNOR U38844 ( .A(n30048), .B(n30049), .Z(n30032) );
  XNOR U38845 ( .A(n30043), .B(n30044), .Z(n30049) );
  XNOR U38846 ( .A(n30045), .B(n30046), .Z(n30044) );
  XNOR U38847 ( .A(y[3973]), .B(x[3973]), .Z(n30046) );
  XNOR U38848 ( .A(y[3974]), .B(x[3974]), .Z(n30045) );
  XNOR U38849 ( .A(y[3972]), .B(x[3972]), .Z(n30043) );
  XNOR U38850 ( .A(n30037), .B(n30038), .Z(n30048) );
  XNOR U38851 ( .A(y[3969]), .B(x[3969]), .Z(n30038) );
  XNOR U38852 ( .A(n30039), .B(n30040), .Z(n30037) );
  XNOR U38853 ( .A(y[3970]), .B(x[3970]), .Z(n30040) );
  XNOR U38854 ( .A(y[3971]), .B(x[3971]), .Z(n30039) );
  XNOR U38855 ( .A(n30030), .B(n30029), .Z(n30033) );
  XNOR U38856 ( .A(n30025), .B(n30026), .Z(n30029) );
  XNOR U38857 ( .A(y[3966]), .B(x[3966]), .Z(n30026) );
  XNOR U38858 ( .A(n30027), .B(n30028), .Z(n30025) );
  XNOR U38859 ( .A(y[3967]), .B(x[3967]), .Z(n30028) );
  XNOR U38860 ( .A(y[3968]), .B(x[3968]), .Z(n30027) );
  XNOR U38861 ( .A(n30019), .B(n30020), .Z(n30030) );
  XNOR U38862 ( .A(y[3963]), .B(x[3963]), .Z(n30020) );
  XNOR U38863 ( .A(n30021), .B(n30022), .Z(n30019) );
  XNOR U38864 ( .A(y[3964]), .B(x[3964]), .Z(n30022) );
  XNOR U38865 ( .A(y[3965]), .B(x[3965]), .Z(n30021) );
  XOR U38866 ( .A(n29995), .B(n29996), .Z(n30014) );
  XNOR U38867 ( .A(n30011), .B(n30012), .Z(n29996) );
  XNOR U38868 ( .A(n30006), .B(n30007), .Z(n30012) );
  XNOR U38869 ( .A(n30008), .B(n30009), .Z(n30007) );
  XNOR U38870 ( .A(y[3961]), .B(x[3961]), .Z(n30009) );
  XNOR U38871 ( .A(y[3962]), .B(x[3962]), .Z(n30008) );
  XNOR U38872 ( .A(y[3960]), .B(x[3960]), .Z(n30006) );
  XNOR U38873 ( .A(n30000), .B(n30001), .Z(n30011) );
  XNOR U38874 ( .A(y[3957]), .B(x[3957]), .Z(n30001) );
  XNOR U38875 ( .A(n30002), .B(n30003), .Z(n30000) );
  XNOR U38876 ( .A(y[3958]), .B(x[3958]), .Z(n30003) );
  XNOR U38877 ( .A(y[3959]), .B(x[3959]), .Z(n30002) );
  XOR U38878 ( .A(n29994), .B(n29993), .Z(n29995) );
  XNOR U38879 ( .A(n29989), .B(n29990), .Z(n29993) );
  XNOR U38880 ( .A(y[3954]), .B(x[3954]), .Z(n29990) );
  XNOR U38881 ( .A(n29991), .B(n29992), .Z(n29989) );
  XNOR U38882 ( .A(y[3955]), .B(x[3955]), .Z(n29992) );
  XNOR U38883 ( .A(y[3956]), .B(x[3956]), .Z(n29991) );
  XNOR U38884 ( .A(n29983), .B(n29984), .Z(n29994) );
  XNOR U38885 ( .A(y[3951]), .B(x[3951]), .Z(n29984) );
  XNOR U38886 ( .A(n29985), .B(n29986), .Z(n29983) );
  XNOR U38887 ( .A(y[3952]), .B(x[3952]), .Z(n29986) );
  XNOR U38888 ( .A(y[3953]), .B(x[3953]), .Z(n29985) );
  NAND U38889 ( .A(n30050), .B(n30051), .Z(N62728) );
  NANDN U38890 ( .A(n30052), .B(n30053), .Z(n30051) );
  OR U38891 ( .A(n30054), .B(n30055), .Z(n30053) );
  NAND U38892 ( .A(n30054), .B(n30055), .Z(n30050) );
  XOR U38893 ( .A(n30054), .B(n30056), .Z(N62727) );
  XNOR U38894 ( .A(n30052), .B(n30055), .Z(n30056) );
  AND U38895 ( .A(n30057), .B(n30058), .Z(n30055) );
  NANDN U38896 ( .A(n30059), .B(n30060), .Z(n30058) );
  NANDN U38897 ( .A(n30061), .B(n30062), .Z(n30060) );
  NANDN U38898 ( .A(n30062), .B(n30061), .Z(n30057) );
  NAND U38899 ( .A(n30063), .B(n30064), .Z(n30052) );
  NANDN U38900 ( .A(n30065), .B(n30066), .Z(n30064) );
  OR U38901 ( .A(n30067), .B(n30068), .Z(n30066) );
  NAND U38902 ( .A(n30068), .B(n30067), .Z(n30063) );
  AND U38903 ( .A(n30069), .B(n30070), .Z(n30054) );
  NANDN U38904 ( .A(n30071), .B(n30072), .Z(n30070) );
  NANDN U38905 ( .A(n30073), .B(n30074), .Z(n30072) );
  NANDN U38906 ( .A(n30074), .B(n30073), .Z(n30069) );
  XOR U38907 ( .A(n30068), .B(n30075), .Z(N62726) );
  XOR U38908 ( .A(n30065), .B(n30067), .Z(n30075) );
  XNOR U38909 ( .A(n30061), .B(n30076), .Z(n30067) );
  XNOR U38910 ( .A(n30059), .B(n30062), .Z(n30076) );
  NAND U38911 ( .A(n30077), .B(n30078), .Z(n30062) );
  NAND U38912 ( .A(n30079), .B(n30080), .Z(n30078) );
  OR U38913 ( .A(n30081), .B(n30082), .Z(n30079) );
  NANDN U38914 ( .A(n30083), .B(n30081), .Z(n30077) );
  IV U38915 ( .A(n30082), .Z(n30083) );
  NAND U38916 ( .A(n30084), .B(n30085), .Z(n30059) );
  NAND U38917 ( .A(n30086), .B(n30087), .Z(n30085) );
  NANDN U38918 ( .A(n30088), .B(n30089), .Z(n30086) );
  NANDN U38919 ( .A(n30089), .B(n30088), .Z(n30084) );
  AND U38920 ( .A(n30090), .B(n30091), .Z(n30061) );
  NAND U38921 ( .A(n30092), .B(n30093), .Z(n30091) );
  OR U38922 ( .A(n30094), .B(n30095), .Z(n30092) );
  NANDN U38923 ( .A(n30096), .B(n30094), .Z(n30090) );
  NAND U38924 ( .A(n30097), .B(n30098), .Z(n30065) );
  NANDN U38925 ( .A(n30099), .B(n30100), .Z(n30098) );
  OR U38926 ( .A(n30101), .B(n30102), .Z(n30100) );
  NANDN U38927 ( .A(n30103), .B(n30101), .Z(n30097) );
  IV U38928 ( .A(n30102), .Z(n30103) );
  XNOR U38929 ( .A(n30073), .B(n30104), .Z(n30068) );
  XNOR U38930 ( .A(n30071), .B(n30074), .Z(n30104) );
  NAND U38931 ( .A(n30105), .B(n30106), .Z(n30074) );
  NAND U38932 ( .A(n30107), .B(n30108), .Z(n30106) );
  OR U38933 ( .A(n30109), .B(n30110), .Z(n30107) );
  NANDN U38934 ( .A(n30111), .B(n30109), .Z(n30105) );
  IV U38935 ( .A(n30110), .Z(n30111) );
  NAND U38936 ( .A(n30112), .B(n30113), .Z(n30071) );
  NAND U38937 ( .A(n30114), .B(n30115), .Z(n30113) );
  NANDN U38938 ( .A(n30116), .B(n30117), .Z(n30114) );
  NANDN U38939 ( .A(n30117), .B(n30116), .Z(n30112) );
  AND U38940 ( .A(n30118), .B(n30119), .Z(n30073) );
  NAND U38941 ( .A(n30120), .B(n30121), .Z(n30119) );
  OR U38942 ( .A(n30122), .B(n30123), .Z(n30120) );
  NANDN U38943 ( .A(n30124), .B(n30122), .Z(n30118) );
  XNOR U38944 ( .A(n30099), .B(n30125), .Z(N62725) );
  XOR U38945 ( .A(n30101), .B(n30102), .Z(n30125) );
  XNOR U38946 ( .A(n30115), .B(n30126), .Z(n30102) );
  XOR U38947 ( .A(n30116), .B(n30117), .Z(n30126) );
  XOR U38948 ( .A(n30122), .B(n30127), .Z(n30117) );
  XOR U38949 ( .A(n30121), .B(n30124), .Z(n30127) );
  IV U38950 ( .A(n30123), .Z(n30124) );
  NAND U38951 ( .A(n30128), .B(n30129), .Z(n30123) );
  OR U38952 ( .A(n30130), .B(n30131), .Z(n30129) );
  OR U38953 ( .A(n30132), .B(n30133), .Z(n30128) );
  NAND U38954 ( .A(n30134), .B(n30135), .Z(n30121) );
  OR U38955 ( .A(n30136), .B(n30137), .Z(n30135) );
  OR U38956 ( .A(n30138), .B(n30139), .Z(n30134) );
  NOR U38957 ( .A(n30140), .B(n30141), .Z(n30122) );
  ANDN U38958 ( .B(n30142), .A(n30143), .Z(n30116) );
  XNOR U38959 ( .A(n30109), .B(n30144), .Z(n30115) );
  XNOR U38960 ( .A(n30108), .B(n30110), .Z(n30144) );
  NAND U38961 ( .A(n30145), .B(n30146), .Z(n30110) );
  OR U38962 ( .A(n30147), .B(n30148), .Z(n30146) );
  OR U38963 ( .A(n30149), .B(n30150), .Z(n30145) );
  NAND U38964 ( .A(n30151), .B(n30152), .Z(n30108) );
  OR U38965 ( .A(n30153), .B(n30154), .Z(n30152) );
  OR U38966 ( .A(n30155), .B(n30156), .Z(n30151) );
  ANDN U38967 ( .B(n30157), .A(n30158), .Z(n30109) );
  IV U38968 ( .A(n30159), .Z(n30157) );
  ANDN U38969 ( .B(n30160), .A(n30161), .Z(n30101) );
  XOR U38970 ( .A(n30087), .B(n30162), .Z(n30099) );
  XOR U38971 ( .A(n30088), .B(n30089), .Z(n30162) );
  XOR U38972 ( .A(n30094), .B(n30163), .Z(n30089) );
  XOR U38973 ( .A(n30093), .B(n30096), .Z(n30163) );
  IV U38974 ( .A(n30095), .Z(n30096) );
  NAND U38975 ( .A(n30164), .B(n30165), .Z(n30095) );
  OR U38976 ( .A(n30166), .B(n30167), .Z(n30165) );
  OR U38977 ( .A(n30168), .B(n30169), .Z(n30164) );
  NAND U38978 ( .A(n30170), .B(n30171), .Z(n30093) );
  OR U38979 ( .A(n30172), .B(n30173), .Z(n30171) );
  OR U38980 ( .A(n30174), .B(n30175), .Z(n30170) );
  NOR U38981 ( .A(n30176), .B(n30177), .Z(n30094) );
  ANDN U38982 ( .B(n30178), .A(n30179), .Z(n30088) );
  IV U38983 ( .A(n30180), .Z(n30178) );
  XNOR U38984 ( .A(n30081), .B(n30181), .Z(n30087) );
  XNOR U38985 ( .A(n30080), .B(n30082), .Z(n30181) );
  NAND U38986 ( .A(n30182), .B(n30183), .Z(n30082) );
  OR U38987 ( .A(n30184), .B(n30185), .Z(n30183) );
  OR U38988 ( .A(n30186), .B(n30187), .Z(n30182) );
  NAND U38989 ( .A(n30188), .B(n30189), .Z(n30080) );
  OR U38990 ( .A(n30190), .B(n30191), .Z(n30189) );
  OR U38991 ( .A(n30192), .B(n30193), .Z(n30188) );
  ANDN U38992 ( .B(n30194), .A(n30195), .Z(n30081) );
  IV U38993 ( .A(n30196), .Z(n30194) );
  XNOR U38994 ( .A(n30161), .B(n30160), .Z(N62724) );
  XOR U38995 ( .A(n30180), .B(n30179), .Z(n30160) );
  XNOR U38996 ( .A(n30195), .B(n30196), .Z(n30179) );
  XNOR U38997 ( .A(n30190), .B(n30191), .Z(n30196) );
  XNOR U38998 ( .A(n30192), .B(n30193), .Z(n30191) );
  XNOR U38999 ( .A(y[3949]), .B(x[3949]), .Z(n30193) );
  XNOR U39000 ( .A(y[3950]), .B(x[3950]), .Z(n30192) );
  XNOR U39001 ( .A(y[3948]), .B(x[3948]), .Z(n30190) );
  XNOR U39002 ( .A(n30184), .B(n30185), .Z(n30195) );
  XNOR U39003 ( .A(y[3945]), .B(x[3945]), .Z(n30185) );
  XNOR U39004 ( .A(n30186), .B(n30187), .Z(n30184) );
  XNOR U39005 ( .A(y[3946]), .B(x[3946]), .Z(n30187) );
  XNOR U39006 ( .A(y[3947]), .B(x[3947]), .Z(n30186) );
  XNOR U39007 ( .A(n30177), .B(n30176), .Z(n30180) );
  XNOR U39008 ( .A(n30172), .B(n30173), .Z(n30176) );
  XNOR U39009 ( .A(y[3942]), .B(x[3942]), .Z(n30173) );
  XNOR U39010 ( .A(n30174), .B(n30175), .Z(n30172) );
  XNOR U39011 ( .A(y[3943]), .B(x[3943]), .Z(n30175) );
  XNOR U39012 ( .A(y[3944]), .B(x[3944]), .Z(n30174) );
  XNOR U39013 ( .A(n30166), .B(n30167), .Z(n30177) );
  XNOR U39014 ( .A(y[3939]), .B(x[3939]), .Z(n30167) );
  XNOR U39015 ( .A(n30168), .B(n30169), .Z(n30166) );
  XNOR U39016 ( .A(y[3940]), .B(x[3940]), .Z(n30169) );
  XNOR U39017 ( .A(y[3941]), .B(x[3941]), .Z(n30168) );
  XOR U39018 ( .A(n30142), .B(n30143), .Z(n30161) );
  XNOR U39019 ( .A(n30158), .B(n30159), .Z(n30143) );
  XNOR U39020 ( .A(n30153), .B(n30154), .Z(n30159) );
  XNOR U39021 ( .A(n30155), .B(n30156), .Z(n30154) );
  XNOR U39022 ( .A(y[3937]), .B(x[3937]), .Z(n30156) );
  XNOR U39023 ( .A(y[3938]), .B(x[3938]), .Z(n30155) );
  XNOR U39024 ( .A(y[3936]), .B(x[3936]), .Z(n30153) );
  XNOR U39025 ( .A(n30147), .B(n30148), .Z(n30158) );
  XNOR U39026 ( .A(y[3933]), .B(x[3933]), .Z(n30148) );
  XNOR U39027 ( .A(n30149), .B(n30150), .Z(n30147) );
  XNOR U39028 ( .A(y[3934]), .B(x[3934]), .Z(n30150) );
  XNOR U39029 ( .A(y[3935]), .B(x[3935]), .Z(n30149) );
  XOR U39030 ( .A(n30141), .B(n30140), .Z(n30142) );
  XNOR U39031 ( .A(n30136), .B(n30137), .Z(n30140) );
  XNOR U39032 ( .A(y[3930]), .B(x[3930]), .Z(n30137) );
  XNOR U39033 ( .A(n30138), .B(n30139), .Z(n30136) );
  XNOR U39034 ( .A(y[3931]), .B(x[3931]), .Z(n30139) );
  XNOR U39035 ( .A(y[3932]), .B(x[3932]), .Z(n30138) );
  XNOR U39036 ( .A(n30130), .B(n30131), .Z(n30141) );
  XNOR U39037 ( .A(y[3927]), .B(x[3927]), .Z(n30131) );
  XNOR U39038 ( .A(n30132), .B(n30133), .Z(n30130) );
  XNOR U39039 ( .A(y[3928]), .B(x[3928]), .Z(n30133) );
  XNOR U39040 ( .A(y[3929]), .B(x[3929]), .Z(n30132) );
  NAND U39041 ( .A(n30197), .B(n30198), .Z(N62715) );
  NANDN U39042 ( .A(n30199), .B(n30200), .Z(n30198) );
  OR U39043 ( .A(n30201), .B(n30202), .Z(n30200) );
  NAND U39044 ( .A(n30201), .B(n30202), .Z(n30197) );
  XOR U39045 ( .A(n30201), .B(n30203), .Z(N62714) );
  XNOR U39046 ( .A(n30199), .B(n30202), .Z(n30203) );
  AND U39047 ( .A(n30204), .B(n30205), .Z(n30202) );
  NANDN U39048 ( .A(n30206), .B(n30207), .Z(n30205) );
  NANDN U39049 ( .A(n30208), .B(n30209), .Z(n30207) );
  NANDN U39050 ( .A(n30209), .B(n30208), .Z(n30204) );
  NAND U39051 ( .A(n30210), .B(n30211), .Z(n30199) );
  NANDN U39052 ( .A(n30212), .B(n30213), .Z(n30211) );
  OR U39053 ( .A(n30214), .B(n30215), .Z(n30213) );
  NAND U39054 ( .A(n30215), .B(n30214), .Z(n30210) );
  AND U39055 ( .A(n30216), .B(n30217), .Z(n30201) );
  NANDN U39056 ( .A(n30218), .B(n30219), .Z(n30217) );
  NANDN U39057 ( .A(n30220), .B(n30221), .Z(n30219) );
  NANDN U39058 ( .A(n30221), .B(n30220), .Z(n30216) );
  XOR U39059 ( .A(n30215), .B(n30222), .Z(N62713) );
  XOR U39060 ( .A(n30212), .B(n30214), .Z(n30222) );
  XNOR U39061 ( .A(n30208), .B(n30223), .Z(n30214) );
  XNOR U39062 ( .A(n30206), .B(n30209), .Z(n30223) );
  NAND U39063 ( .A(n30224), .B(n30225), .Z(n30209) );
  NAND U39064 ( .A(n30226), .B(n30227), .Z(n30225) );
  OR U39065 ( .A(n30228), .B(n30229), .Z(n30226) );
  NANDN U39066 ( .A(n30230), .B(n30228), .Z(n30224) );
  IV U39067 ( .A(n30229), .Z(n30230) );
  NAND U39068 ( .A(n30231), .B(n30232), .Z(n30206) );
  NAND U39069 ( .A(n30233), .B(n30234), .Z(n30232) );
  NANDN U39070 ( .A(n30235), .B(n30236), .Z(n30233) );
  NANDN U39071 ( .A(n30236), .B(n30235), .Z(n30231) );
  AND U39072 ( .A(n30237), .B(n30238), .Z(n30208) );
  NAND U39073 ( .A(n30239), .B(n30240), .Z(n30238) );
  OR U39074 ( .A(n30241), .B(n30242), .Z(n30239) );
  NANDN U39075 ( .A(n30243), .B(n30241), .Z(n30237) );
  NAND U39076 ( .A(n30244), .B(n30245), .Z(n30212) );
  NANDN U39077 ( .A(n30246), .B(n30247), .Z(n30245) );
  OR U39078 ( .A(n30248), .B(n30249), .Z(n30247) );
  NANDN U39079 ( .A(n30250), .B(n30248), .Z(n30244) );
  IV U39080 ( .A(n30249), .Z(n30250) );
  XNOR U39081 ( .A(n30220), .B(n30251), .Z(n30215) );
  XNOR U39082 ( .A(n30218), .B(n30221), .Z(n30251) );
  NAND U39083 ( .A(n30252), .B(n30253), .Z(n30221) );
  NAND U39084 ( .A(n30254), .B(n30255), .Z(n30253) );
  OR U39085 ( .A(n30256), .B(n30257), .Z(n30254) );
  NANDN U39086 ( .A(n30258), .B(n30256), .Z(n30252) );
  IV U39087 ( .A(n30257), .Z(n30258) );
  NAND U39088 ( .A(n30259), .B(n30260), .Z(n30218) );
  NAND U39089 ( .A(n30261), .B(n30262), .Z(n30260) );
  NANDN U39090 ( .A(n30263), .B(n30264), .Z(n30261) );
  NANDN U39091 ( .A(n30264), .B(n30263), .Z(n30259) );
  AND U39092 ( .A(n30265), .B(n30266), .Z(n30220) );
  NAND U39093 ( .A(n30267), .B(n30268), .Z(n30266) );
  OR U39094 ( .A(n30269), .B(n30270), .Z(n30267) );
  NANDN U39095 ( .A(n30271), .B(n30269), .Z(n30265) );
  XNOR U39096 ( .A(n30246), .B(n30272), .Z(N62712) );
  XOR U39097 ( .A(n30248), .B(n30249), .Z(n30272) );
  XNOR U39098 ( .A(n30262), .B(n30273), .Z(n30249) );
  XOR U39099 ( .A(n30263), .B(n30264), .Z(n30273) );
  XOR U39100 ( .A(n30269), .B(n30274), .Z(n30264) );
  XOR U39101 ( .A(n30268), .B(n30271), .Z(n30274) );
  IV U39102 ( .A(n30270), .Z(n30271) );
  NAND U39103 ( .A(n30275), .B(n30276), .Z(n30270) );
  OR U39104 ( .A(n30277), .B(n30278), .Z(n30276) );
  OR U39105 ( .A(n30279), .B(n30280), .Z(n30275) );
  NAND U39106 ( .A(n30281), .B(n30282), .Z(n30268) );
  OR U39107 ( .A(n30283), .B(n30284), .Z(n30282) );
  OR U39108 ( .A(n30285), .B(n30286), .Z(n30281) );
  NOR U39109 ( .A(n30287), .B(n30288), .Z(n30269) );
  ANDN U39110 ( .B(n30289), .A(n30290), .Z(n30263) );
  XNOR U39111 ( .A(n30256), .B(n30291), .Z(n30262) );
  XNOR U39112 ( .A(n30255), .B(n30257), .Z(n30291) );
  NAND U39113 ( .A(n30292), .B(n30293), .Z(n30257) );
  OR U39114 ( .A(n30294), .B(n30295), .Z(n30293) );
  OR U39115 ( .A(n30296), .B(n30297), .Z(n30292) );
  NAND U39116 ( .A(n30298), .B(n30299), .Z(n30255) );
  OR U39117 ( .A(n30300), .B(n30301), .Z(n30299) );
  OR U39118 ( .A(n30302), .B(n30303), .Z(n30298) );
  ANDN U39119 ( .B(n30304), .A(n30305), .Z(n30256) );
  IV U39120 ( .A(n30306), .Z(n30304) );
  ANDN U39121 ( .B(n30307), .A(n30308), .Z(n30248) );
  XOR U39122 ( .A(n30234), .B(n30309), .Z(n30246) );
  XOR U39123 ( .A(n30235), .B(n30236), .Z(n30309) );
  XOR U39124 ( .A(n30241), .B(n30310), .Z(n30236) );
  XOR U39125 ( .A(n30240), .B(n30243), .Z(n30310) );
  IV U39126 ( .A(n30242), .Z(n30243) );
  NAND U39127 ( .A(n30311), .B(n30312), .Z(n30242) );
  OR U39128 ( .A(n30313), .B(n30314), .Z(n30312) );
  OR U39129 ( .A(n30315), .B(n30316), .Z(n30311) );
  NAND U39130 ( .A(n30317), .B(n30318), .Z(n30240) );
  OR U39131 ( .A(n30319), .B(n30320), .Z(n30318) );
  OR U39132 ( .A(n30321), .B(n30322), .Z(n30317) );
  NOR U39133 ( .A(n30323), .B(n30324), .Z(n30241) );
  ANDN U39134 ( .B(n30325), .A(n30326), .Z(n30235) );
  IV U39135 ( .A(n30327), .Z(n30325) );
  XNOR U39136 ( .A(n30228), .B(n30328), .Z(n30234) );
  XNOR U39137 ( .A(n30227), .B(n30229), .Z(n30328) );
  NAND U39138 ( .A(n30329), .B(n30330), .Z(n30229) );
  OR U39139 ( .A(n30331), .B(n30332), .Z(n30330) );
  OR U39140 ( .A(n30333), .B(n30334), .Z(n30329) );
  NAND U39141 ( .A(n30335), .B(n30336), .Z(n30227) );
  OR U39142 ( .A(n30337), .B(n30338), .Z(n30336) );
  OR U39143 ( .A(n30339), .B(n30340), .Z(n30335) );
  ANDN U39144 ( .B(n30341), .A(n30342), .Z(n30228) );
  IV U39145 ( .A(n30343), .Z(n30341) );
  XNOR U39146 ( .A(n30308), .B(n30307), .Z(N62711) );
  XOR U39147 ( .A(n30327), .B(n30326), .Z(n30307) );
  XNOR U39148 ( .A(n30342), .B(n30343), .Z(n30326) );
  XNOR U39149 ( .A(n30337), .B(n30338), .Z(n30343) );
  XNOR U39150 ( .A(n30339), .B(n30340), .Z(n30338) );
  XNOR U39151 ( .A(y[3925]), .B(x[3925]), .Z(n30340) );
  XNOR U39152 ( .A(y[3926]), .B(x[3926]), .Z(n30339) );
  XNOR U39153 ( .A(y[3924]), .B(x[3924]), .Z(n30337) );
  XNOR U39154 ( .A(n30331), .B(n30332), .Z(n30342) );
  XNOR U39155 ( .A(y[3921]), .B(x[3921]), .Z(n30332) );
  XNOR U39156 ( .A(n30333), .B(n30334), .Z(n30331) );
  XNOR U39157 ( .A(y[3922]), .B(x[3922]), .Z(n30334) );
  XNOR U39158 ( .A(y[3923]), .B(x[3923]), .Z(n30333) );
  XNOR U39159 ( .A(n30324), .B(n30323), .Z(n30327) );
  XNOR U39160 ( .A(n30319), .B(n30320), .Z(n30323) );
  XNOR U39161 ( .A(y[3918]), .B(x[3918]), .Z(n30320) );
  XNOR U39162 ( .A(n30321), .B(n30322), .Z(n30319) );
  XNOR U39163 ( .A(y[3919]), .B(x[3919]), .Z(n30322) );
  XNOR U39164 ( .A(y[3920]), .B(x[3920]), .Z(n30321) );
  XNOR U39165 ( .A(n30313), .B(n30314), .Z(n30324) );
  XNOR U39166 ( .A(y[3915]), .B(x[3915]), .Z(n30314) );
  XNOR U39167 ( .A(n30315), .B(n30316), .Z(n30313) );
  XNOR U39168 ( .A(y[3916]), .B(x[3916]), .Z(n30316) );
  XNOR U39169 ( .A(y[3917]), .B(x[3917]), .Z(n30315) );
  XOR U39170 ( .A(n30289), .B(n30290), .Z(n30308) );
  XNOR U39171 ( .A(n30305), .B(n30306), .Z(n30290) );
  XNOR U39172 ( .A(n30300), .B(n30301), .Z(n30306) );
  XNOR U39173 ( .A(n30302), .B(n30303), .Z(n30301) );
  XNOR U39174 ( .A(y[3913]), .B(x[3913]), .Z(n30303) );
  XNOR U39175 ( .A(y[3914]), .B(x[3914]), .Z(n30302) );
  XNOR U39176 ( .A(y[3912]), .B(x[3912]), .Z(n30300) );
  XNOR U39177 ( .A(n30294), .B(n30295), .Z(n30305) );
  XNOR U39178 ( .A(y[3909]), .B(x[3909]), .Z(n30295) );
  XNOR U39179 ( .A(n30296), .B(n30297), .Z(n30294) );
  XNOR U39180 ( .A(y[3910]), .B(x[3910]), .Z(n30297) );
  XNOR U39181 ( .A(y[3911]), .B(x[3911]), .Z(n30296) );
  XOR U39182 ( .A(n30288), .B(n30287), .Z(n30289) );
  XNOR U39183 ( .A(n30283), .B(n30284), .Z(n30287) );
  XNOR U39184 ( .A(y[3906]), .B(x[3906]), .Z(n30284) );
  XNOR U39185 ( .A(n30285), .B(n30286), .Z(n30283) );
  XNOR U39186 ( .A(y[3907]), .B(x[3907]), .Z(n30286) );
  XNOR U39187 ( .A(y[3908]), .B(x[3908]), .Z(n30285) );
  XNOR U39188 ( .A(n30277), .B(n30278), .Z(n30288) );
  XNOR U39189 ( .A(y[3903]), .B(x[3903]), .Z(n30278) );
  XNOR U39190 ( .A(n30279), .B(n30280), .Z(n30277) );
  XNOR U39191 ( .A(y[3904]), .B(x[3904]), .Z(n30280) );
  XNOR U39192 ( .A(y[3905]), .B(x[3905]), .Z(n30279) );
  NAND U39193 ( .A(n30344), .B(n30345), .Z(N62702) );
  NANDN U39194 ( .A(n30346), .B(n30347), .Z(n30345) );
  OR U39195 ( .A(n30348), .B(n30349), .Z(n30347) );
  NAND U39196 ( .A(n30348), .B(n30349), .Z(n30344) );
  XOR U39197 ( .A(n30348), .B(n30350), .Z(N62701) );
  XNOR U39198 ( .A(n30346), .B(n30349), .Z(n30350) );
  AND U39199 ( .A(n30351), .B(n30352), .Z(n30349) );
  NANDN U39200 ( .A(n30353), .B(n30354), .Z(n30352) );
  NANDN U39201 ( .A(n30355), .B(n30356), .Z(n30354) );
  NANDN U39202 ( .A(n30356), .B(n30355), .Z(n30351) );
  NAND U39203 ( .A(n30357), .B(n30358), .Z(n30346) );
  NANDN U39204 ( .A(n30359), .B(n30360), .Z(n30358) );
  OR U39205 ( .A(n30361), .B(n30362), .Z(n30360) );
  NAND U39206 ( .A(n30362), .B(n30361), .Z(n30357) );
  AND U39207 ( .A(n30363), .B(n30364), .Z(n30348) );
  NANDN U39208 ( .A(n30365), .B(n30366), .Z(n30364) );
  NANDN U39209 ( .A(n30367), .B(n30368), .Z(n30366) );
  NANDN U39210 ( .A(n30368), .B(n30367), .Z(n30363) );
  XOR U39211 ( .A(n30362), .B(n30369), .Z(N62700) );
  XOR U39212 ( .A(n30359), .B(n30361), .Z(n30369) );
  XNOR U39213 ( .A(n30355), .B(n30370), .Z(n30361) );
  XNOR U39214 ( .A(n30353), .B(n30356), .Z(n30370) );
  NAND U39215 ( .A(n30371), .B(n30372), .Z(n30356) );
  NAND U39216 ( .A(n30373), .B(n30374), .Z(n30372) );
  OR U39217 ( .A(n30375), .B(n30376), .Z(n30373) );
  NANDN U39218 ( .A(n30377), .B(n30375), .Z(n30371) );
  IV U39219 ( .A(n30376), .Z(n30377) );
  NAND U39220 ( .A(n30378), .B(n30379), .Z(n30353) );
  NAND U39221 ( .A(n30380), .B(n30381), .Z(n30379) );
  NANDN U39222 ( .A(n30382), .B(n30383), .Z(n30380) );
  NANDN U39223 ( .A(n30383), .B(n30382), .Z(n30378) );
  AND U39224 ( .A(n30384), .B(n30385), .Z(n30355) );
  NAND U39225 ( .A(n30386), .B(n30387), .Z(n30385) );
  OR U39226 ( .A(n30388), .B(n30389), .Z(n30386) );
  NANDN U39227 ( .A(n30390), .B(n30388), .Z(n30384) );
  NAND U39228 ( .A(n30391), .B(n30392), .Z(n30359) );
  NANDN U39229 ( .A(n30393), .B(n30394), .Z(n30392) );
  OR U39230 ( .A(n30395), .B(n30396), .Z(n30394) );
  NANDN U39231 ( .A(n30397), .B(n30395), .Z(n30391) );
  IV U39232 ( .A(n30396), .Z(n30397) );
  XNOR U39233 ( .A(n30367), .B(n30398), .Z(n30362) );
  XNOR U39234 ( .A(n30365), .B(n30368), .Z(n30398) );
  NAND U39235 ( .A(n30399), .B(n30400), .Z(n30368) );
  NAND U39236 ( .A(n30401), .B(n30402), .Z(n30400) );
  OR U39237 ( .A(n30403), .B(n30404), .Z(n30401) );
  NANDN U39238 ( .A(n30405), .B(n30403), .Z(n30399) );
  IV U39239 ( .A(n30404), .Z(n30405) );
  NAND U39240 ( .A(n30406), .B(n30407), .Z(n30365) );
  NAND U39241 ( .A(n30408), .B(n30409), .Z(n30407) );
  NANDN U39242 ( .A(n30410), .B(n30411), .Z(n30408) );
  NANDN U39243 ( .A(n30411), .B(n30410), .Z(n30406) );
  AND U39244 ( .A(n30412), .B(n30413), .Z(n30367) );
  NAND U39245 ( .A(n30414), .B(n30415), .Z(n30413) );
  OR U39246 ( .A(n30416), .B(n30417), .Z(n30414) );
  NANDN U39247 ( .A(n30418), .B(n30416), .Z(n30412) );
  XNOR U39248 ( .A(n30393), .B(n30419), .Z(N62699) );
  XOR U39249 ( .A(n30395), .B(n30396), .Z(n30419) );
  XNOR U39250 ( .A(n30409), .B(n30420), .Z(n30396) );
  XOR U39251 ( .A(n30410), .B(n30411), .Z(n30420) );
  XOR U39252 ( .A(n30416), .B(n30421), .Z(n30411) );
  XOR U39253 ( .A(n30415), .B(n30418), .Z(n30421) );
  IV U39254 ( .A(n30417), .Z(n30418) );
  NAND U39255 ( .A(n30422), .B(n30423), .Z(n30417) );
  OR U39256 ( .A(n30424), .B(n30425), .Z(n30423) );
  OR U39257 ( .A(n30426), .B(n30427), .Z(n30422) );
  NAND U39258 ( .A(n30428), .B(n30429), .Z(n30415) );
  OR U39259 ( .A(n30430), .B(n30431), .Z(n30429) );
  OR U39260 ( .A(n30432), .B(n30433), .Z(n30428) );
  NOR U39261 ( .A(n30434), .B(n30435), .Z(n30416) );
  ANDN U39262 ( .B(n30436), .A(n30437), .Z(n30410) );
  XNOR U39263 ( .A(n30403), .B(n30438), .Z(n30409) );
  XNOR U39264 ( .A(n30402), .B(n30404), .Z(n30438) );
  NAND U39265 ( .A(n30439), .B(n30440), .Z(n30404) );
  OR U39266 ( .A(n30441), .B(n30442), .Z(n30440) );
  OR U39267 ( .A(n30443), .B(n30444), .Z(n30439) );
  NAND U39268 ( .A(n30445), .B(n30446), .Z(n30402) );
  OR U39269 ( .A(n30447), .B(n30448), .Z(n30446) );
  OR U39270 ( .A(n30449), .B(n30450), .Z(n30445) );
  ANDN U39271 ( .B(n30451), .A(n30452), .Z(n30403) );
  IV U39272 ( .A(n30453), .Z(n30451) );
  ANDN U39273 ( .B(n30454), .A(n30455), .Z(n30395) );
  XOR U39274 ( .A(n30381), .B(n30456), .Z(n30393) );
  XOR U39275 ( .A(n30382), .B(n30383), .Z(n30456) );
  XOR U39276 ( .A(n30388), .B(n30457), .Z(n30383) );
  XOR U39277 ( .A(n30387), .B(n30390), .Z(n30457) );
  IV U39278 ( .A(n30389), .Z(n30390) );
  NAND U39279 ( .A(n30458), .B(n30459), .Z(n30389) );
  OR U39280 ( .A(n30460), .B(n30461), .Z(n30459) );
  OR U39281 ( .A(n30462), .B(n30463), .Z(n30458) );
  NAND U39282 ( .A(n30464), .B(n30465), .Z(n30387) );
  OR U39283 ( .A(n30466), .B(n30467), .Z(n30465) );
  OR U39284 ( .A(n30468), .B(n30469), .Z(n30464) );
  NOR U39285 ( .A(n30470), .B(n30471), .Z(n30388) );
  ANDN U39286 ( .B(n30472), .A(n30473), .Z(n30382) );
  IV U39287 ( .A(n30474), .Z(n30472) );
  XNOR U39288 ( .A(n30375), .B(n30475), .Z(n30381) );
  XNOR U39289 ( .A(n30374), .B(n30376), .Z(n30475) );
  NAND U39290 ( .A(n30476), .B(n30477), .Z(n30376) );
  OR U39291 ( .A(n30478), .B(n30479), .Z(n30477) );
  OR U39292 ( .A(n30480), .B(n30481), .Z(n30476) );
  NAND U39293 ( .A(n30482), .B(n30483), .Z(n30374) );
  OR U39294 ( .A(n30484), .B(n30485), .Z(n30483) );
  OR U39295 ( .A(n30486), .B(n30487), .Z(n30482) );
  ANDN U39296 ( .B(n30488), .A(n30489), .Z(n30375) );
  IV U39297 ( .A(n30490), .Z(n30488) );
  XNOR U39298 ( .A(n30455), .B(n30454), .Z(N62698) );
  XOR U39299 ( .A(n30474), .B(n30473), .Z(n30454) );
  XNOR U39300 ( .A(n30489), .B(n30490), .Z(n30473) );
  XNOR U39301 ( .A(n30484), .B(n30485), .Z(n30490) );
  XNOR U39302 ( .A(n30486), .B(n30487), .Z(n30485) );
  XNOR U39303 ( .A(y[3901]), .B(x[3901]), .Z(n30487) );
  XNOR U39304 ( .A(y[3902]), .B(x[3902]), .Z(n30486) );
  XNOR U39305 ( .A(y[3900]), .B(x[3900]), .Z(n30484) );
  XNOR U39306 ( .A(n30478), .B(n30479), .Z(n30489) );
  XNOR U39307 ( .A(y[3897]), .B(x[3897]), .Z(n30479) );
  XNOR U39308 ( .A(n30480), .B(n30481), .Z(n30478) );
  XNOR U39309 ( .A(y[3898]), .B(x[3898]), .Z(n30481) );
  XNOR U39310 ( .A(y[3899]), .B(x[3899]), .Z(n30480) );
  XNOR U39311 ( .A(n30471), .B(n30470), .Z(n30474) );
  XNOR U39312 ( .A(n30466), .B(n30467), .Z(n30470) );
  XNOR U39313 ( .A(y[3894]), .B(x[3894]), .Z(n30467) );
  XNOR U39314 ( .A(n30468), .B(n30469), .Z(n30466) );
  XNOR U39315 ( .A(y[3895]), .B(x[3895]), .Z(n30469) );
  XNOR U39316 ( .A(y[3896]), .B(x[3896]), .Z(n30468) );
  XNOR U39317 ( .A(n30460), .B(n30461), .Z(n30471) );
  XNOR U39318 ( .A(y[3891]), .B(x[3891]), .Z(n30461) );
  XNOR U39319 ( .A(n30462), .B(n30463), .Z(n30460) );
  XNOR U39320 ( .A(y[3892]), .B(x[3892]), .Z(n30463) );
  XNOR U39321 ( .A(y[3893]), .B(x[3893]), .Z(n30462) );
  XOR U39322 ( .A(n30436), .B(n30437), .Z(n30455) );
  XNOR U39323 ( .A(n30452), .B(n30453), .Z(n30437) );
  XNOR U39324 ( .A(n30447), .B(n30448), .Z(n30453) );
  XNOR U39325 ( .A(n30449), .B(n30450), .Z(n30448) );
  XNOR U39326 ( .A(y[3889]), .B(x[3889]), .Z(n30450) );
  XNOR U39327 ( .A(y[3890]), .B(x[3890]), .Z(n30449) );
  XNOR U39328 ( .A(y[3888]), .B(x[3888]), .Z(n30447) );
  XNOR U39329 ( .A(n30441), .B(n30442), .Z(n30452) );
  XNOR U39330 ( .A(y[3885]), .B(x[3885]), .Z(n30442) );
  XNOR U39331 ( .A(n30443), .B(n30444), .Z(n30441) );
  XNOR U39332 ( .A(y[3886]), .B(x[3886]), .Z(n30444) );
  XNOR U39333 ( .A(y[3887]), .B(x[3887]), .Z(n30443) );
  XOR U39334 ( .A(n30435), .B(n30434), .Z(n30436) );
  XNOR U39335 ( .A(n30430), .B(n30431), .Z(n30434) );
  XNOR U39336 ( .A(y[3882]), .B(x[3882]), .Z(n30431) );
  XNOR U39337 ( .A(n30432), .B(n30433), .Z(n30430) );
  XNOR U39338 ( .A(y[3883]), .B(x[3883]), .Z(n30433) );
  XNOR U39339 ( .A(y[3884]), .B(x[3884]), .Z(n30432) );
  XNOR U39340 ( .A(n30424), .B(n30425), .Z(n30435) );
  XNOR U39341 ( .A(y[3879]), .B(x[3879]), .Z(n30425) );
  XNOR U39342 ( .A(n30426), .B(n30427), .Z(n30424) );
  XNOR U39343 ( .A(y[3880]), .B(x[3880]), .Z(n30427) );
  XNOR U39344 ( .A(y[3881]), .B(x[3881]), .Z(n30426) );
  NAND U39345 ( .A(n30491), .B(n30492), .Z(N62689) );
  NANDN U39346 ( .A(n30493), .B(n30494), .Z(n30492) );
  OR U39347 ( .A(n30495), .B(n30496), .Z(n30494) );
  NAND U39348 ( .A(n30495), .B(n30496), .Z(n30491) );
  XOR U39349 ( .A(n30495), .B(n30497), .Z(N62688) );
  XNOR U39350 ( .A(n30493), .B(n30496), .Z(n30497) );
  AND U39351 ( .A(n30498), .B(n30499), .Z(n30496) );
  NANDN U39352 ( .A(n30500), .B(n30501), .Z(n30499) );
  NANDN U39353 ( .A(n30502), .B(n30503), .Z(n30501) );
  NANDN U39354 ( .A(n30503), .B(n30502), .Z(n30498) );
  NAND U39355 ( .A(n30504), .B(n30505), .Z(n30493) );
  NANDN U39356 ( .A(n30506), .B(n30507), .Z(n30505) );
  OR U39357 ( .A(n30508), .B(n30509), .Z(n30507) );
  NAND U39358 ( .A(n30509), .B(n30508), .Z(n30504) );
  AND U39359 ( .A(n30510), .B(n30511), .Z(n30495) );
  NANDN U39360 ( .A(n30512), .B(n30513), .Z(n30511) );
  NANDN U39361 ( .A(n30514), .B(n30515), .Z(n30513) );
  NANDN U39362 ( .A(n30515), .B(n30514), .Z(n30510) );
  XOR U39363 ( .A(n30509), .B(n30516), .Z(N62687) );
  XOR U39364 ( .A(n30506), .B(n30508), .Z(n30516) );
  XNOR U39365 ( .A(n30502), .B(n30517), .Z(n30508) );
  XNOR U39366 ( .A(n30500), .B(n30503), .Z(n30517) );
  NAND U39367 ( .A(n30518), .B(n30519), .Z(n30503) );
  NAND U39368 ( .A(n30520), .B(n30521), .Z(n30519) );
  OR U39369 ( .A(n30522), .B(n30523), .Z(n30520) );
  NANDN U39370 ( .A(n30524), .B(n30522), .Z(n30518) );
  IV U39371 ( .A(n30523), .Z(n30524) );
  NAND U39372 ( .A(n30525), .B(n30526), .Z(n30500) );
  NAND U39373 ( .A(n30527), .B(n30528), .Z(n30526) );
  NANDN U39374 ( .A(n30529), .B(n30530), .Z(n30527) );
  NANDN U39375 ( .A(n30530), .B(n30529), .Z(n30525) );
  AND U39376 ( .A(n30531), .B(n30532), .Z(n30502) );
  NAND U39377 ( .A(n30533), .B(n30534), .Z(n30532) );
  OR U39378 ( .A(n30535), .B(n30536), .Z(n30533) );
  NANDN U39379 ( .A(n30537), .B(n30535), .Z(n30531) );
  NAND U39380 ( .A(n30538), .B(n30539), .Z(n30506) );
  NANDN U39381 ( .A(n30540), .B(n30541), .Z(n30539) );
  OR U39382 ( .A(n30542), .B(n30543), .Z(n30541) );
  NANDN U39383 ( .A(n30544), .B(n30542), .Z(n30538) );
  IV U39384 ( .A(n30543), .Z(n30544) );
  XNOR U39385 ( .A(n30514), .B(n30545), .Z(n30509) );
  XNOR U39386 ( .A(n30512), .B(n30515), .Z(n30545) );
  NAND U39387 ( .A(n30546), .B(n30547), .Z(n30515) );
  NAND U39388 ( .A(n30548), .B(n30549), .Z(n30547) );
  OR U39389 ( .A(n30550), .B(n30551), .Z(n30548) );
  NANDN U39390 ( .A(n30552), .B(n30550), .Z(n30546) );
  IV U39391 ( .A(n30551), .Z(n30552) );
  NAND U39392 ( .A(n30553), .B(n30554), .Z(n30512) );
  NAND U39393 ( .A(n30555), .B(n30556), .Z(n30554) );
  NANDN U39394 ( .A(n30557), .B(n30558), .Z(n30555) );
  NANDN U39395 ( .A(n30558), .B(n30557), .Z(n30553) );
  AND U39396 ( .A(n30559), .B(n30560), .Z(n30514) );
  NAND U39397 ( .A(n30561), .B(n30562), .Z(n30560) );
  OR U39398 ( .A(n30563), .B(n30564), .Z(n30561) );
  NANDN U39399 ( .A(n30565), .B(n30563), .Z(n30559) );
  XNOR U39400 ( .A(n30540), .B(n30566), .Z(N62686) );
  XOR U39401 ( .A(n30542), .B(n30543), .Z(n30566) );
  XNOR U39402 ( .A(n30556), .B(n30567), .Z(n30543) );
  XOR U39403 ( .A(n30557), .B(n30558), .Z(n30567) );
  XOR U39404 ( .A(n30563), .B(n30568), .Z(n30558) );
  XOR U39405 ( .A(n30562), .B(n30565), .Z(n30568) );
  IV U39406 ( .A(n30564), .Z(n30565) );
  NAND U39407 ( .A(n30569), .B(n30570), .Z(n30564) );
  OR U39408 ( .A(n30571), .B(n30572), .Z(n30570) );
  OR U39409 ( .A(n30573), .B(n30574), .Z(n30569) );
  NAND U39410 ( .A(n30575), .B(n30576), .Z(n30562) );
  OR U39411 ( .A(n30577), .B(n30578), .Z(n30576) );
  OR U39412 ( .A(n30579), .B(n30580), .Z(n30575) );
  NOR U39413 ( .A(n30581), .B(n30582), .Z(n30563) );
  ANDN U39414 ( .B(n30583), .A(n30584), .Z(n30557) );
  XNOR U39415 ( .A(n30550), .B(n30585), .Z(n30556) );
  XNOR U39416 ( .A(n30549), .B(n30551), .Z(n30585) );
  NAND U39417 ( .A(n30586), .B(n30587), .Z(n30551) );
  OR U39418 ( .A(n30588), .B(n30589), .Z(n30587) );
  OR U39419 ( .A(n30590), .B(n30591), .Z(n30586) );
  NAND U39420 ( .A(n30592), .B(n30593), .Z(n30549) );
  OR U39421 ( .A(n30594), .B(n30595), .Z(n30593) );
  OR U39422 ( .A(n30596), .B(n30597), .Z(n30592) );
  ANDN U39423 ( .B(n30598), .A(n30599), .Z(n30550) );
  IV U39424 ( .A(n30600), .Z(n30598) );
  ANDN U39425 ( .B(n30601), .A(n30602), .Z(n30542) );
  XOR U39426 ( .A(n30528), .B(n30603), .Z(n30540) );
  XOR U39427 ( .A(n30529), .B(n30530), .Z(n30603) );
  XOR U39428 ( .A(n30535), .B(n30604), .Z(n30530) );
  XOR U39429 ( .A(n30534), .B(n30537), .Z(n30604) );
  IV U39430 ( .A(n30536), .Z(n30537) );
  NAND U39431 ( .A(n30605), .B(n30606), .Z(n30536) );
  OR U39432 ( .A(n30607), .B(n30608), .Z(n30606) );
  OR U39433 ( .A(n30609), .B(n30610), .Z(n30605) );
  NAND U39434 ( .A(n30611), .B(n30612), .Z(n30534) );
  OR U39435 ( .A(n30613), .B(n30614), .Z(n30612) );
  OR U39436 ( .A(n30615), .B(n30616), .Z(n30611) );
  NOR U39437 ( .A(n30617), .B(n30618), .Z(n30535) );
  ANDN U39438 ( .B(n30619), .A(n30620), .Z(n30529) );
  IV U39439 ( .A(n30621), .Z(n30619) );
  XNOR U39440 ( .A(n30522), .B(n30622), .Z(n30528) );
  XNOR U39441 ( .A(n30521), .B(n30523), .Z(n30622) );
  NAND U39442 ( .A(n30623), .B(n30624), .Z(n30523) );
  OR U39443 ( .A(n30625), .B(n30626), .Z(n30624) );
  OR U39444 ( .A(n30627), .B(n30628), .Z(n30623) );
  NAND U39445 ( .A(n30629), .B(n30630), .Z(n30521) );
  OR U39446 ( .A(n30631), .B(n30632), .Z(n30630) );
  OR U39447 ( .A(n30633), .B(n30634), .Z(n30629) );
  ANDN U39448 ( .B(n30635), .A(n30636), .Z(n30522) );
  IV U39449 ( .A(n30637), .Z(n30635) );
  XNOR U39450 ( .A(n30602), .B(n30601), .Z(N62685) );
  XOR U39451 ( .A(n30621), .B(n30620), .Z(n30601) );
  XNOR U39452 ( .A(n30636), .B(n30637), .Z(n30620) );
  XNOR U39453 ( .A(n30631), .B(n30632), .Z(n30637) );
  XNOR U39454 ( .A(n30633), .B(n30634), .Z(n30632) );
  XNOR U39455 ( .A(y[3877]), .B(x[3877]), .Z(n30634) );
  XNOR U39456 ( .A(y[3878]), .B(x[3878]), .Z(n30633) );
  XNOR U39457 ( .A(y[3876]), .B(x[3876]), .Z(n30631) );
  XNOR U39458 ( .A(n30625), .B(n30626), .Z(n30636) );
  XNOR U39459 ( .A(y[3873]), .B(x[3873]), .Z(n30626) );
  XNOR U39460 ( .A(n30627), .B(n30628), .Z(n30625) );
  XNOR U39461 ( .A(y[3874]), .B(x[3874]), .Z(n30628) );
  XNOR U39462 ( .A(y[3875]), .B(x[3875]), .Z(n30627) );
  XNOR U39463 ( .A(n30618), .B(n30617), .Z(n30621) );
  XNOR U39464 ( .A(n30613), .B(n30614), .Z(n30617) );
  XNOR U39465 ( .A(y[3870]), .B(x[3870]), .Z(n30614) );
  XNOR U39466 ( .A(n30615), .B(n30616), .Z(n30613) );
  XNOR U39467 ( .A(y[3871]), .B(x[3871]), .Z(n30616) );
  XNOR U39468 ( .A(y[3872]), .B(x[3872]), .Z(n30615) );
  XNOR U39469 ( .A(n30607), .B(n30608), .Z(n30618) );
  XNOR U39470 ( .A(y[3867]), .B(x[3867]), .Z(n30608) );
  XNOR U39471 ( .A(n30609), .B(n30610), .Z(n30607) );
  XNOR U39472 ( .A(y[3868]), .B(x[3868]), .Z(n30610) );
  XNOR U39473 ( .A(y[3869]), .B(x[3869]), .Z(n30609) );
  XOR U39474 ( .A(n30583), .B(n30584), .Z(n30602) );
  XNOR U39475 ( .A(n30599), .B(n30600), .Z(n30584) );
  XNOR U39476 ( .A(n30594), .B(n30595), .Z(n30600) );
  XNOR U39477 ( .A(n30596), .B(n30597), .Z(n30595) );
  XNOR U39478 ( .A(y[3865]), .B(x[3865]), .Z(n30597) );
  XNOR U39479 ( .A(y[3866]), .B(x[3866]), .Z(n30596) );
  XNOR U39480 ( .A(y[3864]), .B(x[3864]), .Z(n30594) );
  XNOR U39481 ( .A(n30588), .B(n30589), .Z(n30599) );
  XNOR U39482 ( .A(y[3861]), .B(x[3861]), .Z(n30589) );
  XNOR U39483 ( .A(n30590), .B(n30591), .Z(n30588) );
  XNOR U39484 ( .A(y[3862]), .B(x[3862]), .Z(n30591) );
  XNOR U39485 ( .A(y[3863]), .B(x[3863]), .Z(n30590) );
  XOR U39486 ( .A(n30582), .B(n30581), .Z(n30583) );
  XNOR U39487 ( .A(n30577), .B(n30578), .Z(n30581) );
  XNOR U39488 ( .A(y[3858]), .B(x[3858]), .Z(n30578) );
  XNOR U39489 ( .A(n30579), .B(n30580), .Z(n30577) );
  XNOR U39490 ( .A(y[3859]), .B(x[3859]), .Z(n30580) );
  XNOR U39491 ( .A(y[3860]), .B(x[3860]), .Z(n30579) );
  XNOR U39492 ( .A(n30571), .B(n30572), .Z(n30582) );
  XNOR U39493 ( .A(y[3855]), .B(x[3855]), .Z(n30572) );
  XNOR U39494 ( .A(n30573), .B(n30574), .Z(n30571) );
  XNOR U39495 ( .A(y[3856]), .B(x[3856]), .Z(n30574) );
  XNOR U39496 ( .A(y[3857]), .B(x[3857]), .Z(n30573) );
  NAND U39497 ( .A(n30638), .B(n30639), .Z(N62676) );
  NANDN U39498 ( .A(n30640), .B(n30641), .Z(n30639) );
  OR U39499 ( .A(n30642), .B(n30643), .Z(n30641) );
  NAND U39500 ( .A(n30642), .B(n30643), .Z(n30638) );
  XOR U39501 ( .A(n30642), .B(n30644), .Z(N62675) );
  XNOR U39502 ( .A(n30640), .B(n30643), .Z(n30644) );
  AND U39503 ( .A(n30645), .B(n30646), .Z(n30643) );
  NANDN U39504 ( .A(n30647), .B(n30648), .Z(n30646) );
  NANDN U39505 ( .A(n30649), .B(n30650), .Z(n30648) );
  NANDN U39506 ( .A(n30650), .B(n30649), .Z(n30645) );
  NAND U39507 ( .A(n30651), .B(n30652), .Z(n30640) );
  NANDN U39508 ( .A(n30653), .B(n30654), .Z(n30652) );
  OR U39509 ( .A(n30655), .B(n30656), .Z(n30654) );
  NAND U39510 ( .A(n30656), .B(n30655), .Z(n30651) );
  AND U39511 ( .A(n30657), .B(n30658), .Z(n30642) );
  NANDN U39512 ( .A(n30659), .B(n30660), .Z(n30658) );
  NANDN U39513 ( .A(n30661), .B(n30662), .Z(n30660) );
  NANDN U39514 ( .A(n30662), .B(n30661), .Z(n30657) );
  XOR U39515 ( .A(n30656), .B(n30663), .Z(N62674) );
  XOR U39516 ( .A(n30653), .B(n30655), .Z(n30663) );
  XNOR U39517 ( .A(n30649), .B(n30664), .Z(n30655) );
  XNOR U39518 ( .A(n30647), .B(n30650), .Z(n30664) );
  NAND U39519 ( .A(n30665), .B(n30666), .Z(n30650) );
  NAND U39520 ( .A(n30667), .B(n30668), .Z(n30666) );
  OR U39521 ( .A(n30669), .B(n30670), .Z(n30667) );
  NANDN U39522 ( .A(n30671), .B(n30669), .Z(n30665) );
  IV U39523 ( .A(n30670), .Z(n30671) );
  NAND U39524 ( .A(n30672), .B(n30673), .Z(n30647) );
  NAND U39525 ( .A(n30674), .B(n30675), .Z(n30673) );
  NANDN U39526 ( .A(n30676), .B(n30677), .Z(n30674) );
  NANDN U39527 ( .A(n30677), .B(n30676), .Z(n30672) );
  AND U39528 ( .A(n30678), .B(n30679), .Z(n30649) );
  NAND U39529 ( .A(n30680), .B(n30681), .Z(n30679) );
  OR U39530 ( .A(n30682), .B(n30683), .Z(n30680) );
  NANDN U39531 ( .A(n30684), .B(n30682), .Z(n30678) );
  NAND U39532 ( .A(n30685), .B(n30686), .Z(n30653) );
  NANDN U39533 ( .A(n30687), .B(n30688), .Z(n30686) );
  OR U39534 ( .A(n30689), .B(n30690), .Z(n30688) );
  NANDN U39535 ( .A(n30691), .B(n30689), .Z(n30685) );
  IV U39536 ( .A(n30690), .Z(n30691) );
  XNOR U39537 ( .A(n30661), .B(n30692), .Z(n30656) );
  XNOR U39538 ( .A(n30659), .B(n30662), .Z(n30692) );
  NAND U39539 ( .A(n30693), .B(n30694), .Z(n30662) );
  NAND U39540 ( .A(n30695), .B(n30696), .Z(n30694) );
  OR U39541 ( .A(n30697), .B(n30698), .Z(n30695) );
  NANDN U39542 ( .A(n30699), .B(n30697), .Z(n30693) );
  IV U39543 ( .A(n30698), .Z(n30699) );
  NAND U39544 ( .A(n30700), .B(n30701), .Z(n30659) );
  NAND U39545 ( .A(n30702), .B(n30703), .Z(n30701) );
  NANDN U39546 ( .A(n30704), .B(n30705), .Z(n30702) );
  NANDN U39547 ( .A(n30705), .B(n30704), .Z(n30700) );
  AND U39548 ( .A(n30706), .B(n30707), .Z(n30661) );
  NAND U39549 ( .A(n30708), .B(n30709), .Z(n30707) );
  OR U39550 ( .A(n30710), .B(n30711), .Z(n30708) );
  NANDN U39551 ( .A(n30712), .B(n30710), .Z(n30706) );
  XNOR U39552 ( .A(n30687), .B(n30713), .Z(N62673) );
  XOR U39553 ( .A(n30689), .B(n30690), .Z(n30713) );
  XNOR U39554 ( .A(n30703), .B(n30714), .Z(n30690) );
  XOR U39555 ( .A(n30704), .B(n30705), .Z(n30714) );
  XOR U39556 ( .A(n30710), .B(n30715), .Z(n30705) );
  XOR U39557 ( .A(n30709), .B(n30712), .Z(n30715) );
  IV U39558 ( .A(n30711), .Z(n30712) );
  NAND U39559 ( .A(n30716), .B(n30717), .Z(n30711) );
  OR U39560 ( .A(n30718), .B(n30719), .Z(n30717) );
  OR U39561 ( .A(n30720), .B(n30721), .Z(n30716) );
  NAND U39562 ( .A(n30722), .B(n30723), .Z(n30709) );
  OR U39563 ( .A(n30724), .B(n30725), .Z(n30723) );
  OR U39564 ( .A(n30726), .B(n30727), .Z(n30722) );
  NOR U39565 ( .A(n30728), .B(n30729), .Z(n30710) );
  ANDN U39566 ( .B(n30730), .A(n30731), .Z(n30704) );
  XNOR U39567 ( .A(n30697), .B(n30732), .Z(n30703) );
  XNOR U39568 ( .A(n30696), .B(n30698), .Z(n30732) );
  NAND U39569 ( .A(n30733), .B(n30734), .Z(n30698) );
  OR U39570 ( .A(n30735), .B(n30736), .Z(n30734) );
  OR U39571 ( .A(n30737), .B(n30738), .Z(n30733) );
  NAND U39572 ( .A(n30739), .B(n30740), .Z(n30696) );
  OR U39573 ( .A(n30741), .B(n30742), .Z(n30740) );
  OR U39574 ( .A(n30743), .B(n30744), .Z(n30739) );
  ANDN U39575 ( .B(n30745), .A(n30746), .Z(n30697) );
  IV U39576 ( .A(n30747), .Z(n30745) );
  ANDN U39577 ( .B(n30748), .A(n30749), .Z(n30689) );
  XOR U39578 ( .A(n30675), .B(n30750), .Z(n30687) );
  XOR U39579 ( .A(n30676), .B(n30677), .Z(n30750) );
  XOR U39580 ( .A(n30682), .B(n30751), .Z(n30677) );
  XOR U39581 ( .A(n30681), .B(n30684), .Z(n30751) );
  IV U39582 ( .A(n30683), .Z(n30684) );
  NAND U39583 ( .A(n30752), .B(n30753), .Z(n30683) );
  OR U39584 ( .A(n30754), .B(n30755), .Z(n30753) );
  OR U39585 ( .A(n30756), .B(n30757), .Z(n30752) );
  NAND U39586 ( .A(n30758), .B(n30759), .Z(n30681) );
  OR U39587 ( .A(n30760), .B(n30761), .Z(n30759) );
  OR U39588 ( .A(n30762), .B(n30763), .Z(n30758) );
  NOR U39589 ( .A(n30764), .B(n30765), .Z(n30682) );
  ANDN U39590 ( .B(n30766), .A(n30767), .Z(n30676) );
  IV U39591 ( .A(n30768), .Z(n30766) );
  XNOR U39592 ( .A(n30669), .B(n30769), .Z(n30675) );
  XNOR U39593 ( .A(n30668), .B(n30670), .Z(n30769) );
  NAND U39594 ( .A(n30770), .B(n30771), .Z(n30670) );
  OR U39595 ( .A(n30772), .B(n30773), .Z(n30771) );
  OR U39596 ( .A(n30774), .B(n30775), .Z(n30770) );
  NAND U39597 ( .A(n30776), .B(n30777), .Z(n30668) );
  OR U39598 ( .A(n30778), .B(n30779), .Z(n30777) );
  OR U39599 ( .A(n30780), .B(n30781), .Z(n30776) );
  ANDN U39600 ( .B(n30782), .A(n30783), .Z(n30669) );
  IV U39601 ( .A(n30784), .Z(n30782) );
  XNOR U39602 ( .A(n30749), .B(n30748), .Z(N62672) );
  XOR U39603 ( .A(n30768), .B(n30767), .Z(n30748) );
  XNOR U39604 ( .A(n30783), .B(n30784), .Z(n30767) );
  XNOR U39605 ( .A(n30778), .B(n30779), .Z(n30784) );
  XNOR U39606 ( .A(n30780), .B(n30781), .Z(n30779) );
  XNOR U39607 ( .A(y[3853]), .B(x[3853]), .Z(n30781) );
  XNOR U39608 ( .A(y[3854]), .B(x[3854]), .Z(n30780) );
  XNOR U39609 ( .A(y[3852]), .B(x[3852]), .Z(n30778) );
  XNOR U39610 ( .A(n30772), .B(n30773), .Z(n30783) );
  XNOR U39611 ( .A(y[3849]), .B(x[3849]), .Z(n30773) );
  XNOR U39612 ( .A(n30774), .B(n30775), .Z(n30772) );
  XNOR U39613 ( .A(y[3850]), .B(x[3850]), .Z(n30775) );
  XNOR U39614 ( .A(y[3851]), .B(x[3851]), .Z(n30774) );
  XNOR U39615 ( .A(n30765), .B(n30764), .Z(n30768) );
  XNOR U39616 ( .A(n30760), .B(n30761), .Z(n30764) );
  XNOR U39617 ( .A(y[3846]), .B(x[3846]), .Z(n30761) );
  XNOR U39618 ( .A(n30762), .B(n30763), .Z(n30760) );
  XNOR U39619 ( .A(y[3847]), .B(x[3847]), .Z(n30763) );
  XNOR U39620 ( .A(y[3848]), .B(x[3848]), .Z(n30762) );
  XNOR U39621 ( .A(n30754), .B(n30755), .Z(n30765) );
  XNOR U39622 ( .A(y[3843]), .B(x[3843]), .Z(n30755) );
  XNOR U39623 ( .A(n30756), .B(n30757), .Z(n30754) );
  XNOR U39624 ( .A(y[3844]), .B(x[3844]), .Z(n30757) );
  XNOR U39625 ( .A(y[3845]), .B(x[3845]), .Z(n30756) );
  XOR U39626 ( .A(n30730), .B(n30731), .Z(n30749) );
  XNOR U39627 ( .A(n30746), .B(n30747), .Z(n30731) );
  XNOR U39628 ( .A(n30741), .B(n30742), .Z(n30747) );
  XNOR U39629 ( .A(n30743), .B(n30744), .Z(n30742) );
  XNOR U39630 ( .A(y[3841]), .B(x[3841]), .Z(n30744) );
  XNOR U39631 ( .A(y[3842]), .B(x[3842]), .Z(n30743) );
  XNOR U39632 ( .A(y[3840]), .B(x[3840]), .Z(n30741) );
  XNOR U39633 ( .A(n30735), .B(n30736), .Z(n30746) );
  XNOR U39634 ( .A(y[3837]), .B(x[3837]), .Z(n30736) );
  XNOR U39635 ( .A(n30737), .B(n30738), .Z(n30735) );
  XNOR U39636 ( .A(y[3838]), .B(x[3838]), .Z(n30738) );
  XNOR U39637 ( .A(y[3839]), .B(x[3839]), .Z(n30737) );
  XOR U39638 ( .A(n30729), .B(n30728), .Z(n30730) );
  XNOR U39639 ( .A(n30724), .B(n30725), .Z(n30728) );
  XNOR U39640 ( .A(y[3834]), .B(x[3834]), .Z(n30725) );
  XNOR U39641 ( .A(n30726), .B(n30727), .Z(n30724) );
  XNOR U39642 ( .A(y[3835]), .B(x[3835]), .Z(n30727) );
  XNOR U39643 ( .A(y[3836]), .B(x[3836]), .Z(n30726) );
  XNOR U39644 ( .A(n30718), .B(n30719), .Z(n30729) );
  XNOR U39645 ( .A(y[3831]), .B(x[3831]), .Z(n30719) );
  XNOR U39646 ( .A(n30720), .B(n30721), .Z(n30718) );
  XNOR U39647 ( .A(y[3832]), .B(x[3832]), .Z(n30721) );
  XNOR U39648 ( .A(y[3833]), .B(x[3833]), .Z(n30720) );
  NAND U39649 ( .A(n30785), .B(n30786), .Z(N62663) );
  NANDN U39650 ( .A(n30787), .B(n30788), .Z(n30786) );
  OR U39651 ( .A(n30789), .B(n30790), .Z(n30788) );
  NAND U39652 ( .A(n30789), .B(n30790), .Z(n30785) );
  XOR U39653 ( .A(n30789), .B(n30791), .Z(N62662) );
  XNOR U39654 ( .A(n30787), .B(n30790), .Z(n30791) );
  AND U39655 ( .A(n30792), .B(n30793), .Z(n30790) );
  NANDN U39656 ( .A(n30794), .B(n30795), .Z(n30793) );
  NANDN U39657 ( .A(n30796), .B(n30797), .Z(n30795) );
  NANDN U39658 ( .A(n30797), .B(n30796), .Z(n30792) );
  NAND U39659 ( .A(n30798), .B(n30799), .Z(n30787) );
  NANDN U39660 ( .A(n30800), .B(n30801), .Z(n30799) );
  OR U39661 ( .A(n30802), .B(n30803), .Z(n30801) );
  NAND U39662 ( .A(n30803), .B(n30802), .Z(n30798) );
  AND U39663 ( .A(n30804), .B(n30805), .Z(n30789) );
  NANDN U39664 ( .A(n30806), .B(n30807), .Z(n30805) );
  NANDN U39665 ( .A(n30808), .B(n30809), .Z(n30807) );
  NANDN U39666 ( .A(n30809), .B(n30808), .Z(n30804) );
  XOR U39667 ( .A(n30803), .B(n30810), .Z(N62661) );
  XOR U39668 ( .A(n30800), .B(n30802), .Z(n30810) );
  XNOR U39669 ( .A(n30796), .B(n30811), .Z(n30802) );
  XNOR U39670 ( .A(n30794), .B(n30797), .Z(n30811) );
  NAND U39671 ( .A(n30812), .B(n30813), .Z(n30797) );
  NAND U39672 ( .A(n30814), .B(n30815), .Z(n30813) );
  OR U39673 ( .A(n30816), .B(n30817), .Z(n30814) );
  NANDN U39674 ( .A(n30818), .B(n30816), .Z(n30812) );
  IV U39675 ( .A(n30817), .Z(n30818) );
  NAND U39676 ( .A(n30819), .B(n30820), .Z(n30794) );
  NAND U39677 ( .A(n30821), .B(n30822), .Z(n30820) );
  NANDN U39678 ( .A(n30823), .B(n30824), .Z(n30821) );
  NANDN U39679 ( .A(n30824), .B(n30823), .Z(n30819) );
  AND U39680 ( .A(n30825), .B(n30826), .Z(n30796) );
  NAND U39681 ( .A(n30827), .B(n30828), .Z(n30826) );
  OR U39682 ( .A(n30829), .B(n30830), .Z(n30827) );
  NANDN U39683 ( .A(n30831), .B(n30829), .Z(n30825) );
  NAND U39684 ( .A(n30832), .B(n30833), .Z(n30800) );
  NANDN U39685 ( .A(n30834), .B(n30835), .Z(n30833) );
  OR U39686 ( .A(n30836), .B(n30837), .Z(n30835) );
  NANDN U39687 ( .A(n30838), .B(n30836), .Z(n30832) );
  IV U39688 ( .A(n30837), .Z(n30838) );
  XNOR U39689 ( .A(n30808), .B(n30839), .Z(n30803) );
  XNOR U39690 ( .A(n30806), .B(n30809), .Z(n30839) );
  NAND U39691 ( .A(n30840), .B(n30841), .Z(n30809) );
  NAND U39692 ( .A(n30842), .B(n30843), .Z(n30841) );
  OR U39693 ( .A(n30844), .B(n30845), .Z(n30842) );
  NANDN U39694 ( .A(n30846), .B(n30844), .Z(n30840) );
  IV U39695 ( .A(n30845), .Z(n30846) );
  NAND U39696 ( .A(n30847), .B(n30848), .Z(n30806) );
  NAND U39697 ( .A(n30849), .B(n30850), .Z(n30848) );
  NANDN U39698 ( .A(n30851), .B(n30852), .Z(n30849) );
  NANDN U39699 ( .A(n30852), .B(n30851), .Z(n30847) );
  AND U39700 ( .A(n30853), .B(n30854), .Z(n30808) );
  NAND U39701 ( .A(n30855), .B(n30856), .Z(n30854) );
  OR U39702 ( .A(n30857), .B(n30858), .Z(n30855) );
  NANDN U39703 ( .A(n30859), .B(n30857), .Z(n30853) );
  XNOR U39704 ( .A(n30834), .B(n30860), .Z(N62660) );
  XOR U39705 ( .A(n30836), .B(n30837), .Z(n30860) );
  XNOR U39706 ( .A(n30850), .B(n30861), .Z(n30837) );
  XOR U39707 ( .A(n30851), .B(n30852), .Z(n30861) );
  XOR U39708 ( .A(n30857), .B(n30862), .Z(n30852) );
  XOR U39709 ( .A(n30856), .B(n30859), .Z(n30862) );
  IV U39710 ( .A(n30858), .Z(n30859) );
  NAND U39711 ( .A(n30863), .B(n30864), .Z(n30858) );
  OR U39712 ( .A(n30865), .B(n30866), .Z(n30864) );
  OR U39713 ( .A(n30867), .B(n30868), .Z(n30863) );
  NAND U39714 ( .A(n30869), .B(n30870), .Z(n30856) );
  OR U39715 ( .A(n30871), .B(n30872), .Z(n30870) );
  OR U39716 ( .A(n30873), .B(n30874), .Z(n30869) );
  NOR U39717 ( .A(n30875), .B(n30876), .Z(n30857) );
  ANDN U39718 ( .B(n30877), .A(n30878), .Z(n30851) );
  XNOR U39719 ( .A(n30844), .B(n30879), .Z(n30850) );
  XNOR U39720 ( .A(n30843), .B(n30845), .Z(n30879) );
  NAND U39721 ( .A(n30880), .B(n30881), .Z(n30845) );
  OR U39722 ( .A(n30882), .B(n30883), .Z(n30881) );
  OR U39723 ( .A(n30884), .B(n30885), .Z(n30880) );
  NAND U39724 ( .A(n30886), .B(n30887), .Z(n30843) );
  OR U39725 ( .A(n30888), .B(n30889), .Z(n30887) );
  OR U39726 ( .A(n30890), .B(n30891), .Z(n30886) );
  ANDN U39727 ( .B(n30892), .A(n30893), .Z(n30844) );
  IV U39728 ( .A(n30894), .Z(n30892) );
  ANDN U39729 ( .B(n30895), .A(n30896), .Z(n30836) );
  XOR U39730 ( .A(n30822), .B(n30897), .Z(n30834) );
  XOR U39731 ( .A(n30823), .B(n30824), .Z(n30897) );
  XOR U39732 ( .A(n30829), .B(n30898), .Z(n30824) );
  XOR U39733 ( .A(n30828), .B(n30831), .Z(n30898) );
  IV U39734 ( .A(n30830), .Z(n30831) );
  NAND U39735 ( .A(n30899), .B(n30900), .Z(n30830) );
  OR U39736 ( .A(n30901), .B(n30902), .Z(n30900) );
  OR U39737 ( .A(n30903), .B(n30904), .Z(n30899) );
  NAND U39738 ( .A(n30905), .B(n30906), .Z(n30828) );
  OR U39739 ( .A(n30907), .B(n30908), .Z(n30906) );
  OR U39740 ( .A(n30909), .B(n30910), .Z(n30905) );
  NOR U39741 ( .A(n30911), .B(n30912), .Z(n30829) );
  ANDN U39742 ( .B(n30913), .A(n30914), .Z(n30823) );
  IV U39743 ( .A(n30915), .Z(n30913) );
  XNOR U39744 ( .A(n30816), .B(n30916), .Z(n30822) );
  XNOR U39745 ( .A(n30815), .B(n30817), .Z(n30916) );
  NAND U39746 ( .A(n30917), .B(n30918), .Z(n30817) );
  OR U39747 ( .A(n30919), .B(n30920), .Z(n30918) );
  OR U39748 ( .A(n30921), .B(n30922), .Z(n30917) );
  NAND U39749 ( .A(n30923), .B(n30924), .Z(n30815) );
  OR U39750 ( .A(n30925), .B(n30926), .Z(n30924) );
  OR U39751 ( .A(n30927), .B(n30928), .Z(n30923) );
  ANDN U39752 ( .B(n30929), .A(n30930), .Z(n30816) );
  IV U39753 ( .A(n30931), .Z(n30929) );
  XNOR U39754 ( .A(n30896), .B(n30895), .Z(N62659) );
  XOR U39755 ( .A(n30915), .B(n30914), .Z(n30895) );
  XNOR U39756 ( .A(n30930), .B(n30931), .Z(n30914) );
  XNOR U39757 ( .A(n30925), .B(n30926), .Z(n30931) );
  XNOR U39758 ( .A(n30927), .B(n30928), .Z(n30926) );
  XNOR U39759 ( .A(y[3829]), .B(x[3829]), .Z(n30928) );
  XNOR U39760 ( .A(y[3830]), .B(x[3830]), .Z(n30927) );
  XNOR U39761 ( .A(y[3828]), .B(x[3828]), .Z(n30925) );
  XNOR U39762 ( .A(n30919), .B(n30920), .Z(n30930) );
  XNOR U39763 ( .A(y[3825]), .B(x[3825]), .Z(n30920) );
  XNOR U39764 ( .A(n30921), .B(n30922), .Z(n30919) );
  XNOR U39765 ( .A(y[3826]), .B(x[3826]), .Z(n30922) );
  XNOR U39766 ( .A(y[3827]), .B(x[3827]), .Z(n30921) );
  XNOR U39767 ( .A(n30912), .B(n30911), .Z(n30915) );
  XNOR U39768 ( .A(n30907), .B(n30908), .Z(n30911) );
  XNOR U39769 ( .A(y[3822]), .B(x[3822]), .Z(n30908) );
  XNOR U39770 ( .A(n30909), .B(n30910), .Z(n30907) );
  XNOR U39771 ( .A(y[3823]), .B(x[3823]), .Z(n30910) );
  XNOR U39772 ( .A(y[3824]), .B(x[3824]), .Z(n30909) );
  XNOR U39773 ( .A(n30901), .B(n30902), .Z(n30912) );
  XNOR U39774 ( .A(y[3819]), .B(x[3819]), .Z(n30902) );
  XNOR U39775 ( .A(n30903), .B(n30904), .Z(n30901) );
  XNOR U39776 ( .A(y[3820]), .B(x[3820]), .Z(n30904) );
  XNOR U39777 ( .A(y[3821]), .B(x[3821]), .Z(n30903) );
  XOR U39778 ( .A(n30877), .B(n30878), .Z(n30896) );
  XNOR U39779 ( .A(n30893), .B(n30894), .Z(n30878) );
  XNOR U39780 ( .A(n30888), .B(n30889), .Z(n30894) );
  XNOR U39781 ( .A(n30890), .B(n30891), .Z(n30889) );
  XNOR U39782 ( .A(y[3817]), .B(x[3817]), .Z(n30891) );
  XNOR U39783 ( .A(y[3818]), .B(x[3818]), .Z(n30890) );
  XNOR U39784 ( .A(y[3816]), .B(x[3816]), .Z(n30888) );
  XNOR U39785 ( .A(n30882), .B(n30883), .Z(n30893) );
  XNOR U39786 ( .A(y[3813]), .B(x[3813]), .Z(n30883) );
  XNOR U39787 ( .A(n30884), .B(n30885), .Z(n30882) );
  XNOR U39788 ( .A(y[3814]), .B(x[3814]), .Z(n30885) );
  XNOR U39789 ( .A(y[3815]), .B(x[3815]), .Z(n30884) );
  XOR U39790 ( .A(n30876), .B(n30875), .Z(n30877) );
  XNOR U39791 ( .A(n30871), .B(n30872), .Z(n30875) );
  XNOR U39792 ( .A(y[3810]), .B(x[3810]), .Z(n30872) );
  XNOR U39793 ( .A(n30873), .B(n30874), .Z(n30871) );
  XNOR U39794 ( .A(y[3811]), .B(x[3811]), .Z(n30874) );
  XNOR U39795 ( .A(y[3812]), .B(x[3812]), .Z(n30873) );
  XNOR U39796 ( .A(n30865), .B(n30866), .Z(n30876) );
  XNOR U39797 ( .A(y[3807]), .B(x[3807]), .Z(n30866) );
  XNOR U39798 ( .A(n30867), .B(n30868), .Z(n30865) );
  XNOR U39799 ( .A(y[3808]), .B(x[3808]), .Z(n30868) );
  XNOR U39800 ( .A(y[3809]), .B(x[3809]), .Z(n30867) );
  NAND U39801 ( .A(n30932), .B(n30933), .Z(N62650) );
  NANDN U39802 ( .A(n30934), .B(n30935), .Z(n30933) );
  OR U39803 ( .A(n30936), .B(n30937), .Z(n30935) );
  NAND U39804 ( .A(n30936), .B(n30937), .Z(n30932) );
  XOR U39805 ( .A(n30936), .B(n30938), .Z(N62649) );
  XNOR U39806 ( .A(n30934), .B(n30937), .Z(n30938) );
  AND U39807 ( .A(n30939), .B(n30940), .Z(n30937) );
  NANDN U39808 ( .A(n30941), .B(n30942), .Z(n30940) );
  NANDN U39809 ( .A(n30943), .B(n30944), .Z(n30942) );
  NANDN U39810 ( .A(n30944), .B(n30943), .Z(n30939) );
  NAND U39811 ( .A(n30945), .B(n30946), .Z(n30934) );
  NANDN U39812 ( .A(n30947), .B(n30948), .Z(n30946) );
  OR U39813 ( .A(n30949), .B(n30950), .Z(n30948) );
  NAND U39814 ( .A(n30950), .B(n30949), .Z(n30945) );
  AND U39815 ( .A(n30951), .B(n30952), .Z(n30936) );
  NANDN U39816 ( .A(n30953), .B(n30954), .Z(n30952) );
  NANDN U39817 ( .A(n30955), .B(n30956), .Z(n30954) );
  NANDN U39818 ( .A(n30956), .B(n30955), .Z(n30951) );
  XOR U39819 ( .A(n30950), .B(n30957), .Z(N62648) );
  XOR U39820 ( .A(n30947), .B(n30949), .Z(n30957) );
  XNOR U39821 ( .A(n30943), .B(n30958), .Z(n30949) );
  XNOR U39822 ( .A(n30941), .B(n30944), .Z(n30958) );
  NAND U39823 ( .A(n30959), .B(n30960), .Z(n30944) );
  NAND U39824 ( .A(n30961), .B(n30962), .Z(n30960) );
  OR U39825 ( .A(n30963), .B(n30964), .Z(n30961) );
  NANDN U39826 ( .A(n30965), .B(n30963), .Z(n30959) );
  IV U39827 ( .A(n30964), .Z(n30965) );
  NAND U39828 ( .A(n30966), .B(n30967), .Z(n30941) );
  NAND U39829 ( .A(n30968), .B(n30969), .Z(n30967) );
  NANDN U39830 ( .A(n30970), .B(n30971), .Z(n30968) );
  NANDN U39831 ( .A(n30971), .B(n30970), .Z(n30966) );
  AND U39832 ( .A(n30972), .B(n30973), .Z(n30943) );
  NAND U39833 ( .A(n30974), .B(n30975), .Z(n30973) );
  OR U39834 ( .A(n30976), .B(n30977), .Z(n30974) );
  NANDN U39835 ( .A(n30978), .B(n30976), .Z(n30972) );
  NAND U39836 ( .A(n30979), .B(n30980), .Z(n30947) );
  NANDN U39837 ( .A(n30981), .B(n30982), .Z(n30980) );
  OR U39838 ( .A(n30983), .B(n30984), .Z(n30982) );
  NANDN U39839 ( .A(n30985), .B(n30983), .Z(n30979) );
  IV U39840 ( .A(n30984), .Z(n30985) );
  XNOR U39841 ( .A(n30955), .B(n30986), .Z(n30950) );
  XNOR U39842 ( .A(n30953), .B(n30956), .Z(n30986) );
  NAND U39843 ( .A(n30987), .B(n30988), .Z(n30956) );
  NAND U39844 ( .A(n30989), .B(n30990), .Z(n30988) );
  OR U39845 ( .A(n30991), .B(n30992), .Z(n30989) );
  NANDN U39846 ( .A(n30993), .B(n30991), .Z(n30987) );
  IV U39847 ( .A(n30992), .Z(n30993) );
  NAND U39848 ( .A(n30994), .B(n30995), .Z(n30953) );
  NAND U39849 ( .A(n30996), .B(n30997), .Z(n30995) );
  NANDN U39850 ( .A(n30998), .B(n30999), .Z(n30996) );
  NANDN U39851 ( .A(n30999), .B(n30998), .Z(n30994) );
  AND U39852 ( .A(n31000), .B(n31001), .Z(n30955) );
  NAND U39853 ( .A(n31002), .B(n31003), .Z(n31001) );
  OR U39854 ( .A(n31004), .B(n31005), .Z(n31002) );
  NANDN U39855 ( .A(n31006), .B(n31004), .Z(n31000) );
  XNOR U39856 ( .A(n30981), .B(n31007), .Z(N62647) );
  XOR U39857 ( .A(n30983), .B(n30984), .Z(n31007) );
  XNOR U39858 ( .A(n30997), .B(n31008), .Z(n30984) );
  XOR U39859 ( .A(n30998), .B(n30999), .Z(n31008) );
  XOR U39860 ( .A(n31004), .B(n31009), .Z(n30999) );
  XOR U39861 ( .A(n31003), .B(n31006), .Z(n31009) );
  IV U39862 ( .A(n31005), .Z(n31006) );
  NAND U39863 ( .A(n31010), .B(n31011), .Z(n31005) );
  OR U39864 ( .A(n31012), .B(n31013), .Z(n31011) );
  OR U39865 ( .A(n31014), .B(n31015), .Z(n31010) );
  NAND U39866 ( .A(n31016), .B(n31017), .Z(n31003) );
  OR U39867 ( .A(n31018), .B(n31019), .Z(n31017) );
  OR U39868 ( .A(n31020), .B(n31021), .Z(n31016) );
  NOR U39869 ( .A(n31022), .B(n31023), .Z(n31004) );
  ANDN U39870 ( .B(n31024), .A(n31025), .Z(n30998) );
  XNOR U39871 ( .A(n30991), .B(n31026), .Z(n30997) );
  XNOR U39872 ( .A(n30990), .B(n30992), .Z(n31026) );
  NAND U39873 ( .A(n31027), .B(n31028), .Z(n30992) );
  OR U39874 ( .A(n31029), .B(n31030), .Z(n31028) );
  OR U39875 ( .A(n31031), .B(n31032), .Z(n31027) );
  NAND U39876 ( .A(n31033), .B(n31034), .Z(n30990) );
  OR U39877 ( .A(n31035), .B(n31036), .Z(n31034) );
  OR U39878 ( .A(n31037), .B(n31038), .Z(n31033) );
  ANDN U39879 ( .B(n31039), .A(n31040), .Z(n30991) );
  IV U39880 ( .A(n31041), .Z(n31039) );
  ANDN U39881 ( .B(n31042), .A(n31043), .Z(n30983) );
  XOR U39882 ( .A(n30969), .B(n31044), .Z(n30981) );
  XOR U39883 ( .A(n30970), .B(n30971), .Z(n31044) );
  XOR U39884 ( .A(n30976), .B(n31045), .Z(n30971) );
  XOR U39885 ( .A(n30975), .B(n30978), .Z(n31045) );
  IV U39886 ( .A(n30977), .Z(n30978) );
  NAND U39887 ( .A(n31046), .B(n31047), .Z(n30977) );
  OR U39888 ( .A(n31048), .B(n31049), .Z(n31047) );
  OR U39889 ( .A(n31050), .B(n31051), .Z(n31046) );
  NAND U39890 ( .A(n31052), .B(n31053), .Z(n30975) );
  OR U39891 ( .A(n31054), .B(n31055), .Z(n31053) );
  OR U39892 ( .A(n31056), .B(n31057), .Z(n31052) );
  NOR U39893 ( .A(n31058), .B(n31059), .Z(n30976) );
  ANDN U39894 ( .B(n31060), .A(n31061), .Z(n30970) );
  IV U39895 ( .A(n31062), .Z(n31060) );
  XNOR U39896 ( .A(n30963), .B(n31063), .Z(n30969) );
  XNOR U39897 ( .A(n30962), .B(n30964), .Z(n31063) );
  NAND U39898 ( .A(n31064), .B(n31065), .Z(n30964) );
  OR U39899 ( .A(n31066), .B(n31067), .Z(n31065) );
  OR U39900 ( .A(n31068), .B(n31069), .Z(n31064) );
  NAND U39901 ( .A(n31070), .B(n31071), .Z(n30962) );
  OR U39902 ( .A(n31072), .B(n31073), .Z(n31071) );
  OR U39903 ( .A(n31074), .B(n31075), .Z(n31070) );
  ANDN U39904 ( .B(n31076), .A(n31077), .Z(n30963) );
  IV U39905 ( .A(n31078), .Z(n31076) );
  XNOR U39906 ( .A(n31043), .B(n31042), .Z(N62646) );
  XOR U39907 ( .A(n31062), .B(n31061), .Z(n31042) );
  XNOR U39908 ( .A(n31077), .B(n31078), .Z(n31061) );
  XNOR U39909 ( .A(n31072), .B(n31073), .Z(n31078) );
  XNOR U39910 ( .A(n31074), .B(n31075), .Z(n31073) );
  XNOR U39911 ( .A(y[3805]), .B(x[3805]), .Z(n31075) );
  XNOR U39912 ( .A(y[3806]), .B(x[3806]), .Z(n31074) );
  XNOR U39913 ( .A(y[3804]), .B(x[3804]), .Z(n31072) );
  XNOR U39914 ( .A(n31066), .B(n31067), .Z(n31077) );
  XNOR U39915 ( .A(y[3801]), .B(x[3801]), .Z(n31067) );
  XNOR U39916 ( .A(n31068), .B(n31069), .Z(n31066) );
  XNOR U39917 ( .A(y[3802]), .B(x[3802]), .Z(n31069) );
  XNOR U39918 ( .A(y[3803]), .B(x[3803]), .Z(n31068) );
  XNOR U39919 ( .A(n31059), .B(n31058), .Z(n31062) );
  XNOR U39920 ( .A(n31054), .B(n31055), .Z(n31058) );
  XNOR U39921 ( .A(y[3798]), .B(x[3798]), .Z(n31055) );
  XNOR U39922 ( .A(n31056), .B(n31057), .Z(n31054) );
  XNOR U39923 ( .A(y[3799]), .B(x[3799]), .Z(n31057) );
  XNOR U39924 ( .A(y[3800]), .B(x[3800]), .Z(n31056) );
  XNOR U39925 ( .A(n31048), .B(n31049), .Z(n31059) );
  XNOR U39926 ( .A(y[3795]), .B(x[3795]), .Z(n31049) );
  XNOR U39927 ( .A(n31050), .B(n31051), .Z(n31048) );
  XNOR U39928 ( .A(y[3796]), .B(x[3796]), .Z(n31051) );
  XNOR U39929 ( .A(y[3797]), .B(x[3797]), .Z(n31050) );
  XOR U39930 ( .A(n31024), .B(n31025), .Z(n31043) );
  XNOR U39931 ( .A(n31040), .B(n31041), .Z(n31025) );
  XNOR U39932 ( .A(n31035), .B(n31036), .Z(n31041) );
  XNOR U39933 ( .A(n31037), .B(n31038), .Z(n31036) );
  XNOR U39934 ( .A(y[3793]), .B(x[3793]), .Z(n31038) );
  XNOR U39935 ( .A(y[3794]), .B(x[3794]), .Z(n31037) );
  XNOR U39936 ( .A(y[3792]), .B(x[3792]), .Z(n31035) );
  XNOR U39937 ( .A(n31029), .B(n31030), .Z(n31040) );
  XNOR U39938 ( .A(y[3789]), .B(x[3789]), .Z(n31030) );
  XNOR U39939 ( .A(n31031), .B(n31032), .Z(n31029) );
  XNOR U39940 ( .A(y[3790]), .B(x[3790]), .Z(n31032) );
  XNOR U39941 ( .A(y[3791]), .B(x[3791]), .Z(n31031) );
  XOR U39942 ( .A(n31023), .B(n31022), .Z(n31024) );
  XNOR U39943 ( .A(n31018), .B(n31019), .Z(n31022) );
  XNOR U39944 ( .A(y[3786]), .B(x[3786]), .Z(n31019) );
  XNOR U39945 ( .A(n31020), .B(n31021), .Z(n31018) );
  XNOR U39946 ( .A(y[3787]), .B(x[3787]), .Z(n31021) );
  XNOR U39947 ( .A(y[3788]), .B(x[3788]), .Z(n31020) );
  XNOR U39948 ( .A(n31012), .B(n31013), .Z(n31023) );
  XNOR U39949 ( .A(y[3783]), .B(x[3783]), .Z(n31013) );
  XNOR U39950 ( .A(n31014), .B(n31015), .Z(n31012) );
  XNOR U39951 ( .A(y[3784]), .B(x[3784]), .Z(n31015) );
  XNOR U39952 ( .A(y[3785]), .B(x[3785]), .Z(n31014) );
  NAND U39953 ( .A(n31079), .B(n31080), .Z(N62637) );
  NANDN U39954 ( .A(n31081), .B(n31082), .Z(n31080) );
  OR U39955 ( .A(n31083), .B(n31084), .Z(n31082) );
  NAND U39956 ( .A(n31083), .B(n31084), .Z(n31079) );
  XOR U39957 ( .A(n31083), .B(n31085), .Z(N62636) );
  XNOR U39958 ( .A(n31081), .B(n31084), .Z(n31085) );
  AND U39959 ( .A(n31086), .B(n31087), .Z(n31084) );
  NANDN U39960 ( .A(n31088), .B(n31089), .Z(n31087) );
  NANDN U39961 ( .A(n31090), .B(n31091), .Z(n31089) );
  NANDN U39962 ( .A(n31091), .B(n31090), .Z(n31086) );
  NAND U39963 ( .A(n31092), .B(n31093), .Z(n31081) );
  NANDN U39964 ( .A(n31094), .B(n31095), .Z(n31093) );
  OR U39965 ( .A(n31096), .B(n31097), .Z(n31095) );
  NAND U39966 ( .A(n31097), .B(n31096), .Z(n31092) );
  AND U39967 ( .A(n31098), .B(n31099), .Z(n31083) );
  NANDN U39968 ( .A(n31100), .B(n31101), .Z(n31099) );
  NANDN U39969 ( .A(n31102), .B(n31103), .Z(n31101) );
  NANDN U39970 ( .A(n31103), .B(n31102), .Z(n31098) );
  XOR U39971 ( .A(n31097), .B(n31104), .Z(N62635) );
  XOR U39972 ( .A(n31094), .B(n31096), .Z(n31104) );
  XNOR U39973 ( .A(n31090), .B(n31105), .Z(n31096) );
  XNOR U39974 ( .A(n31088), .B(n31091), .Z(n31105) );
  NAND U39975 ( .A(n31106), .B(n31107), .Z(n31091) );
  NAND U39976 ( .A(n31108), .B(n31109), .Z(n31107) );
  OR U39977 ( .A(n31110), .B(n31111), .Z(n31108) );
  NANDN U39978 ( .A(n31112), .B(n31110), .Z(n31106) );
  IV U39979 ( .A(n31111), .Z(n31112) );
  NAND U39980 ( .A(n31113), .B(n31114), .Z(n31088) );
  NAND U39981 ( .A(n31115), .B(n31116), .Z(n31114) );
  NANDN U39982 ( .A(n31117), .B(n31118), .Z(n31115) );
  NANDN U39983 ( .A(n31118), .B(n31117), .Z(n31113) );
  AND U39984 ( .A(n31119), .B(n31120), .Z(n31090) );
  NAND U39985 ( .A(n31121), .B(n31122), .Z(n31120) );
  OR U39986 ( .A(n31123), .B(n31124), .Z(n31121) );
  NANDN U39987 ( .A(n31125), .B(n31123), .Z(n31119) );
  NAND U39988 ( .A(n31126), .B(n31127), .Z(n31094) );
  NANDN U39989 ( .A(n31128), .B(n31129), .Z(n31127) );
  OR U39990 ( .A(n31130), .B(n31131), .Z(n31129) );
  NANDN U39991 ( .A(n31132), .B(n31130), .Z(n31126) );
  IV U39992 ( .A(n31131), .Z(n31132) );
  XNOR U39993 ( .A(n31102), .B(n31133), .Z(n31097) );
  XNOR U39994 ( .A(n31100), .B(n31103), .Z(n31133) );
  NAND U39995 ( .A(n31134), .B(n31135), .Z(n31103) );
  NAND U39996 ( .A(n31136), .B(n31137), .Z(n31135) );
  OR U39997 ( .A(n31138), .B(n31139), .Z(n31136) );
  NANDN U39998 ( .A(n31140), .B(n31138), .Z(n31134) );
  IV U39999 ( .A(n31139), .Z(n31140) );
  NAND U40000 ( .A(n31141), .B(n31142), .Z(n31100) );
  NAND U40001 ( .A(n31143), .B(n31144), .Z(n31142) );
  NANDN U40002 ( .A(n31145), .B(n31146), .Z(n31143) );
  NANDN U40003 ( .A(n31146), .B(n31145), .Z(n31141) );
  AND U40004 ( .A(n31147), .B(n31148), .Z(n31102) );
  NAND U40005 ( .A(n31149), .B(n31150), .Z(n31148) );
  OR U40006 ( .A(n31151), .B(n31152), .Z(n31149) );
  NANDN U40007 ( .A(n31153), .B(n31151), .Z(n31147) );
  XNOR U40008 ( .A(n31128), .B(n31154), .Z(N62634) );
  XOR U40009 ( .A(n31130), .B(n31131), .Z(n31154) );
  XNOR U40010 ( .A(n31144), .B(n31155), .Z(n31131) );
  XOR U40011 ( .A(n31145), .B(n31146), .Z(n31155) );
  XOR U40012 ( .A(n31151), .B(n31156), .Z(n31146) );
  XOR U40013 ( .A(n31150), .B(n31153), .Z(n31156) );
  IV U40014 ( .A(n31152), .Z(n31153) );
  NAND U40015 ( .A(n31157), .B(n31158), .Z(n31152) );
  OR U40016 ( .A(n31159), .B(n31160), .Z(n31158) );
  OR U40017 ( .A(n31161), .B(n31162), .Z(n31157) );
  NAND U40018 ( .A(n31163), .B(n31164), .Z(n31150) );
  OR U40019 ( .A(n31165), .B(n31166), .Z(n31164) );
  OR U40020 ( .A(n31167), .B(n31168), .Z(n31163) );
  NOR U40021 ( .A(n31169), .B(n31170), .Z(n31151) );
  ANDN U40022 ( .B(n31171), .A(n31172), .Z(n31145) );
  XNOR U40023 ( .A(n31138), .B(n31173), .Z(n31144) );
  XNOR U40024 ( .A(n31137), .B(n31139), .Z(n31173) );
  NAND U40025 ( .A(n31174), .B(n31175), .Z(n31139) );
  OR U40026 ( .A(n31176), .B(n31177), .Z(n31175) );
  OR U40027 ( .A(n31178), .B(n31179), .Z(n31174) );
  NAND U40028 ( .A(n31180), .B(n31181), .Z(n31137) );
  OR U40029 ( .A(n31182), .B(n31183), .Z(n31181) );
  OR U40030 ( .A(n31184), .B(n31185), .Z(n31180) );
  ANDN U40031 ( .B(n31186), .A(n31187), .Z(n31138) );
  IV U40032 ( .A(n31188), .Z(n31186) );
  ANDN U40033 ( .B(n31189), .A(n31190), .Z(n31130) );
  XOR U40034 ( .A(n31116), .B(n31191), .Z(n31128) );
  XOR U40035 ( .A(n31117), .B(n31118), .Z(n31191) );
  XOR U40036 ( .A(n31123), .B(n31192), .Z(n31118) );
  XOR U40037 ( .A(n31122), .B(n31125), .Z(n31192) );
  IV U40038 ( .A(n31124), .Z(n31125) );
  NAND U40039 ( .A(n31193), .B(n31194), .Z(n31124) );
  OR U40040 ( .A(n31195), .B(n31196), .Z(n31194) );
  OR U40041 ( .A(n31197), .B(n31198), .Z(n31193) );
  NAND U40042 ( .A(n31199), .B(n31200), .Z(n31122) );
  OR U40043 ( .A(n31201), .B(n31202), .Z(n31200) );
  OR U40044 ( .A(n31203), .B(n31204), .Z(n31199) );
  NOR U40045 ( .A(n31205), .B(n31206), .Z(n31123) );
  ANDN U40046 ( .B(n31207), .A(n31208), .Z(n31117) );
  IV U40047 ( .A(n31209), .Z(n31207) );
  XNOR U40048 ( .A(n31110), .B(n31210), .Z(n31116) );
  XNOR U40049 ( .A(n31109), .B(n31111), .Z(n31210) );
  NAND U40050 ( .A(n31211), .B(n31212), .Z(n31111) );
  OR U40051 ( .A(n31213), .B(n31214), .Z(n31212) );
  OR U40052 ( .A(n31215), .B(n31216), .Z(n31211) );
  NAND U40053 ( .A(n31217), .B(n31218), .Z(n31109) );
  OR U40054 ( .A(n31219), .B(n31220), .Z(n31218) );
  OR U40055 ( .A(n31221), .B(n31222), .Z(n31217) );
  ANDN U40056 ( .B(n31223), .A(n31224), .Z(n31110) );
  IV U40057 ( .A(n31225), .Z(n31223) );
  XNOR U40058 ( .A(n31190), .B(n31189), .Z(N62633) );
  XOR U40059 ( .A(n31209), .B(n31208), .Z(n31189) );
  XNOR U40060 ( .A(n31224), .B(n31225), .Z(n31208) );
  XNOR U40061 ( .A(n31219), .B(n31220), .Z(n31225) );
  XNOR U40062 ( .A(n31221), .B(n31222), .Z(n31220) );
  XNOR U40063 ( .A(y[3781]), .B(x[3781]), .Z(n31222) );
  XNOR U40064 ( .A(y[3782]), .B(x[3782]), .Z(n31221) );
  XNOR U40065 ( .A(y[3780]), .B(x[3780]), .Z(n31219) );
  XNOR U40066 ( .A(n31213), .B(n31214), .Z(n31224) );
  XNOR U40067 ( .A(y[3777]), .B(x[3777]), .Z(n31214) );
  XNOR U40068 ( .A(n31215), .B(n31216), .Z(n31213) );
  XNOR U40069 ( .A(y[3778]), .B(x[3778]), .Z(n31216) );
  XNOR U40070 ( .A(y[3779]), .B(x[3779]), .Z(n31215) );
  XNOR U40071 ( .A(n31206), .B(n31205), .Z(n31209) );
  XNOR U40072 ( .A(n31201), .B(n31202), .Z(n31205) );
  XNOR U40073 ( .A(y[3774]), .B(x[3774]), .Z(n31202) );
  XNOR U40074 ( .A(n31203), .B(n31204), .Z(n31201) );
  XNOR U40075 ( .A(y[3775]), .B(x[3775]), .Z(n31204) );
  XNOR U40076 ( .A(y[3776]), .B(x[3776]), .Z(n31203) );
  XNOR U40077 ( .A(n31195), .B(n31196), .Z(n31206) );
  XNOR U40078 ( .A(y[3771]), .B(x[3771]), .Z(n31196) );
  XNOR U40079 ( .A(n31197), .B(n31198), .Z(n31195) );
  XNOR U40080 ( .A(y[3772]), .B(x[3772]), .Z(n31198) );
  XNOR U40081 ( .A(y[3773]), .B(x[3773]), .Z(n31197) );
  XOR U40082 ( .A(n31171), .B(n31172), .Z(n31190) );
  XNOR U40083 ( .A(n31187), .B(n31188), .Z(n31172) );
  XNOR U40084 ( .A(n31182), .B(n31183), .Z(n31188) );
  XNOR U40085 ( .A(n31184), .B(n31185), .Z(n31183) );
  XNOR U40086 ( .A(y[3769]), .B(x[3769]), .Z(n31185) );
  XNOR U40087 ( .A(y[3770]), .B(x[3770]), .Z(n31184) );
  XNOR U40088 ( .A(y[3768]), .B(x[3768]), .Z(n31182) );
  XNOR U40089 ( .A(n31176), .B(n31177), .Z(n31187) );
  XNOR U40090 ( .A(y[3765]), .B(x[3765]), .Z(n31177) );
  XNOR U40091 ( .A(n31178), .B(n31179), .Z(n31176) );
  XNOR U40092 ( .A(y[3766]), .B(x[3766]), .Z(n31179) );
  XNOR U40093 ( .A(y[3767]), .B(x[3767]), .Z(n31178) );
  XOR U40094 ( .A(n31170), .B(n31169), .Z(n31171) );
  XNOR U40095 ( .A(n31165), .B(n31166), .Z(n31169) );
  XNOR U40096 ( .A(y[3762]), .B(x[3762]), .Z(n31166) );
  XNOR U40097 ( .A(n31167), .B(n31168), .Z(n31165) );
  XNOR U40098 ( .A(y[3763]), .B(x[3763]), .Z(n31168) );
  XNOR U40099 ( .A(y[3764]), .B(x[3764]), .Z(n31167) );
  XNOR U40100 ( .A(n31159), .B(n31160), .Z(n31170) );
  XNOR U40101 ( .A(y[3759]), .B(x[3759]), .Z(n31160) );
  XNOR U40102 ( .A(n31161), .B(n31162), .Z(n31159) );
  XNOR U40103 ( .A(y[3760]), .B(x[3760]), .Z(n31162) );
  XNOR U40104 ( .A(y[3761]), .B(x[3761]), .Z(n31161) );
  NAND U40105 ( .A(n31226), .B(n31227), .Z(N62624) );
  NANDN U40106 ( .A(n31228), .B(n31229), .Z(n31227) );
  OR U40107 ( .A(n31230), .B(n31231), .Z(n31229) );
  NAND U40108 ( .A(n31230), .B(n31231), .Z(n31226) );
  XOR U40109 ( .A(n31230), .B(n31232), .Z(N62623) );
  XNOR U40110 ( .A(n31228), .B(n31231), .Z(n31232) );
  AND U40111 ( .A(n31233), .B(n31234), .Z(n31231) );
  NANDN U40112 ( .A(n31235), .B(n31236), .Z(n31234) );
  NANDN U40113 ( .A(n31237), .B(n31238), .Z(n31236) );
  NANDN U40114 ( .A(n31238), .B(n31237), .Z(n31233) );
  NAND U40115 ( .A(n31239), .B(n31240), .Z(n31228) );
  NANDN U40116 ( .A(n31241), .B(n31242), .Z(n31240) );
  OR U40117 ( .A(n31243), .B(n31244), .Z(n31242) );
  NAND U40118 ( .A(n31244), .B(n31243), .Z(n31239) );
  AND U40119 ( .A(n31245), .B(n31246), .Z(n31230) );
  NANDN U40120 ( .A(n31247), .B(n31248), .Z(n31246) );
  NANDN U40121 ( .A(n31249), .B(n31250), .Z(n31248) );
  NANDN U40122 ( .A(n31250), .B(n31249), .Z(n31245) );
  XOR U40123 ( .A(n31244), .B(n31251), .Z(N62622) );
  XOR U40124 ( .A(n31241), .B(n31243), .Z(n31251) );
  XNOR U40125 ( .A(n31237), .B(n31252), .Z(n31243) );
  XNOR U40126 ( .A(n31235), .B(n31238), .Z(n31252) );
  NAND U40127 ( .A(n31253), .B(n31254), .Z(n31238) );
  NAND U40128 ( .A(n31255), .B(n31256), .Z(n31254) );
  OR U40129 ( .A(n31257), .B(n31258), .Z(n31255) );
  NANDN U40130 ( .A(n31259), .B(n31257), .Z(n31253) );
  IV U40131 ( .A(n31258), .Z(n31259) );
  NAND U40132 ( .A(n31260), .B(n31261), .Z(n31235) );
  NAND U40133 ( .A(n31262), .B(n31263), .Z(n31261) );
  NANDN U40134 ( .A(n31264), .B(n31265), .Z(n31262) );
  NANDN U40135 ( .A(n31265), .B(n31264), .Z(n31260) );
  AND U40136 ( .A(n31266), .B(n31267), .Z(n31237) );
  NAND U40137 ( .A(n31268), .B(n31269), .Z(n31267) );
  OR U40138 ( .A(n31270), .B(n31271), .Z(n31268) );
  NANDN U40139 ( .A(n31272), .B(n31270), .Z(n31266) );
  NAND U40140 ( .A(n31273), .B(n31274), .Z(n31241) );
  NANDN U40141 ( .A(n31275), .B(n31276), .Z(n31274) );
  OR U40142 ( .A(n31277), .B(n31278), .Z(n31276) );
  NANDN U40143 ( .A(n31279), .B(n31277), .Z(n31273) );
  IV U40144 ( .A(n31278), .Z(n31279) );
  XNOR U40145 ( .A(n31249), .B(n31280), .Z(n31244) );
  XNOR U40146 ( .A(n31247), .B(n31250), .Z(n31280) );
  NAND U40147 ( .A(n31281), .B(n31282), .Z(n31250) );
  NAND U40148 ( .A(n31283), .B(n31284), .Z(n31282) );
  OR U40149 ( .A(n31285), .B(n31286), .Z(n31283) );
  NANDN U40150 ( .A(n31287), .B(n31285), .Z(n31281) );
  IV U40151 ( .A(n31286), .Z(n31287) );
  NAND U40152 ( .A(n31288), .B(n31289), .Z(n31247) );
  NAND U40153 ( .A(n31290), .B(n31291), .Z(n31289) );
  NANDN U40154 ( .A(n31292), .B(n31293), .Z(n31290) );
  NANDN U40155 ( .A(n31293), .B(n31292), .Z(n31288) );
  AND U40156 ( .A(n31294), .B(n31295), .Z(n31249) );
  NAND U40157 ( .A(n31296), .B(n31297), .Z(n31295) );
  OR U40158 ( .A(n31298), .B(n31299), .Z(n31296) );
  NANDN U40159 ( .A(n31300), .B(n31298), .Z(n31294) );
  XNOR U40160 ( .A(n31275), .B(n31301), .Z(N62621) );
  XOR U40161 ( .A(n31277), .B(n31278), .Z(n31301) );
  XNOR U40162 ( .A(n31291), .B(n31302), .Z(n31278) );
  XOR U40163 ( .A(n31292), .B(n31293), .Z(n31302) );
  XOR U40164 ( .A(n31298), .B(n31303), .Z(n31293) );
  XOR U40165 ( .A(n31297), .B(n31300), .Z(n31303) );
  IV U40166 ( .A(n31299), .Z(n31300) );
  NAND U40167 ( .A(n31304), .B(n31305), .Z(n31299) );
  OR U40168 ( .A(n31306), .B(n31307), .Z(n31305) );
  OR U40169 ( .A(n31308), .B(n31309), .Z(n31304) );
  NAND U40170 ( .A(n31310), .B(n31311), .Z(n31297) );
  OR U40171 ( .A(n31312), .B(n31313), .Z(n31311) );
  OR U40172 ( .A(n31314), .B(n31315), .Z(n31310) );
  NOR U40173 ( .A(n31316), .B(n31317), .Z(n31298) );
  ANDN U40174 ( .B(n31318), .A(n31319), .Z(n31292) );
  XNOR U40175 ( .A(n31285), .B(n31320), .Z(n31291) );
  XNOR U40176 ( .A(n31284), .B(n31286), .Z(n31320) );
  NAND U40177 ( .A(n31321), .B(n31322), .Z(n31286) );
  OR U40178 ( .A(n31323), .B(n31324), .Z(n31322) );
  OR U40179 ( .A(n31325), .B(n31326), .Z(n31321) );
  NAND U40180 ( .A(n31327), .B(n31328), .Z(n31284) );
  OR U40181 ( .A(n31329), .B(n31330), .Z(n31328) );
  OR U40182 ( .A(n31331), .B(n31332), .Z(n31327) );
  ANDN U40183 ( .B(n31333), .A(n31334), .Z(n31285) );
  IV U40184 ( .A(n31335), .Z(n31333) );
  ANDN U40185 ( .B(n31336), .A(n31337), .Z(n31277) );
  XOR U40186 ( .A(n31263), .B(n31338), .Z(n31275) );
  XOR U40187 ( .A(n31264), .B(n31265), .Z(n31338) );
  XOR U40188 ( .A(n31270), .B(n31339), .Z(n31265) );
  XOR U40189 ( .A(n31269), .B(n31272), .Z(n31339) );
  IV U40190 ( .A(n31271), .Z(n31272) );
  NAND U40191 ( .A(n31340), .B(n31341), .Z(n31271) );
  OR U40192 ( .A(n31342), .B(n31343), .Z(n31341) );
  OR U40193 ( .A(n31344), .B(n31345), .Z(n31340) );
  NAND U40194 ( .A(n31346), .B(n31347), .Z(n31269) );
  OR U40195 ( .A(n31348), .B(n31349), .Z(n31347) );
  OR U40196 ( .A(n31350), .B(n31351), .Z(n31346) );
  NOR U40197 ( .A(n31352), .B(n31353), .Z(n31270) );
  ANDN U40198 ( .B(n31354), .A(n31355), .Z(n31264) );
  IV U40199 ( .A(n31356), .Z(n31354) );
  XNOR U40200 ( .A(n31257), .B(n31357), .Z(n31263) );
  XNOR U40201 ( .A(n31256), .B(n31258), .Z(n31357) );
  NAND U40202 ( .A(n31358), .B(n31359), .Z(n31258) );
  OR U40203 ( .A(n31360), .B(n31361), .Z(n31359) );
  OR U40204 ( .A(n31362), .B(n31363), .Z(n31358) );
  NAND U40205 ( .A(n31364), .B(n31365), .Z(n31256) );
  OR U40206 ( .A(n31366), .B(n31367), .Z(n31365) );
  OR U40207 ( .A(n31368), .B(n31369), .Z(n31364) );
  ANDN U40208 ( .B(n31370), .A(n31371), .Z(n31257) );
  IV U40209 ( .A(n31372), .Z(n31370) );
  XNOR U40210 ( .A(n31337), .B(n31336), .Z(N62620) );
  XOR U40211 ( .A(n31356), .B(n31355), .Z(n31336) );
  XNOR U40212 ( .A(n31371), .B(n31372), .Z(n31355) );
  XNOR U40213 ( .A(n31366), .B(n31367), .Z(n31372) );
  XNOR U40214 ( .A(n31368), .B(n31369), .Z(n31367) );
  XNOR U40215 ( .A(y[3757]), .B(x[3757]), .Z(n31369) );
  XNOR U40216 ( .A(y[3758]), .B(x[3758]), .Z(n31368) );
  XNOR U40217 ( .A(y[3756]), .B(x[3756]), .Z(n31366) );
  XNOR U40218 ( .A(n31360), .B(n31361), .Z(n31371) );
  XNOR U40219 ( .A(y[3753]), .B(x[3753]), .Z(n31361) );
  XNOR U40220 ( .A(n31362), .B(n31363), .Z(n31360) );
  XNOR U40221 ( .A(y[3754]), .B(x[3754]), .Z(n31363) );
  XNOR U40222 ( .A(y[3755]), .B(x[3755]), .Z(n31362) );
  XNOR U40223 ( .A(n31353), .B(n31352), .Z(n31356) );
  XNOR U40224 ( .A(n31348), .B(n31349), .Z(n31352) );
  XNOR U40225 ( .A(y[3750]), .B(x[3750]), .Z(n31349) );
  XNOR U40226 ( .A(n31350), .B(n31351), .Z(n31348) );
  XNOR U40227 ( .A(y[3751]), .B(x[3751]), .Z(n31351) );
  XNOR U40228 ( .A(y[3752]), .B(x[3752]), .Z(n31350) );
  XNOR U40229 ( .A(n31342), .B(n31343), .Z(n31353) );
  XNOR U40230 ( .A(y[3747]), .B(x[3747]), .Z(n31343) );
  XNOR U40231 ( .A(n31344), .B(n31345), .Z(n31342) );
  XNOR U40232 ( .A(y[3748]), .B(x[3748]), .Z(n31345) );
  XNOR U40233 ( .A(y[3749]), .B(x[3749]), .Z(n31344) );
  XOR U40234 ( .A(n31318), .B(n31319), .Z(n31337) );
  XNOR U40235 ( .A(n31334), .B(n31335), .Z(n31319) );
  XNOR U40236 ( .A(n31329), .B(n31330), .Z(n31335) );
  XNOR U40237 ( .A(n31331), .B(n31332), .Z(n31330) );
  XNOR U40238 ( .A(y[3745]), .B(x[3745]), .Z(n31332) );
  XNOR U40239 ( .A(y[3746]), .B(x[3746]), .Z(n31331) );
  XNOR U40240 ( .A(y[3744]), .B(x[3744]), .Z(n31329) );
  XNOR U40241 ( .A(n31323), .B(n31324), .Z(n31334) );
  XNOR U40242 ( .A(y[3741]), .B(x[3741]), .Z(n31324) );
  XNOR U40243 ( .A(n31325), .B(n31326), .Z(n31323) );
  XNOR U40244 ( .A(y[3742]), .B(x[3742]), .Z(n31326) );
  XNOR U40245 ( .A(y[3743]), .B(x[3743]), .Z(n31325) );
  XOR U40246 ( .A(n31317), .B(n31316), .Z(n31318) );
  XNOR U40247 ( .A(n31312), .B(n31313), .Z(n31316) );
  XNOR U40248 ( .A(y[3738]), .B(x[3738]), .Z(n31313) );
  XNOR U40249 ( .A(n31314), .B(n31315), .Z(n31312) );
  XNOR U40250 ( .A(y[3739]), .B(x[3739]), .Z(n31315) );
  XNOR U40251 ( .A(y[3740]), .B(x[3740]), .Z(n31314) );
  XNOR U40252 ( .A(n31306), .B(n31307), .Z(n31317) );
  XNOR U40253 ( .A(y[3735]), .B(x[3735]), .Z(n31307) );
  XNOR U40254 ( .A(n31308), .B(n31309), .Z(n31306) );
  XNOR U40255 ( .A(y[3736]), .B(x[3736]), .Z(n31309) );
  XNOR U40256 ( .A(y[3737]), .B(x[3737]), .Z(n31308) );
  NAND U40257 ( .A(n31373), .B(n31374), .Z(N62611) );
  NANDN U40258 ( .A(n31375), .B(n31376), .Z(n31374) );
  OR U40259 ( .A(n31377), .B(n31378), .Z(n31376) );
  NAND U40260 ( .A(n31377), .B(n31378), .Z(n31373) );
  XOR U40261 ( .A(n31377), .B(n31379), .Z(N62610) );
  XNOR U40262 ( .A(n31375), .B(n31378), .Z(n31379) );
  AND U40263 ( .A(n31380), .B(n31381), .Z(n31378) );
  NANDN U40264 ( .A(n31382), .B(n31383), .Z(n31381) );
  NANDN U40265 ( .A(n31384), .B(n31385), .Z(n31383) );
  NANDN U40266 ( .A(n31385), .B(n31384), .Z(n31380) );
  NAND U40267 ( .A(n31386), .B(n31387), .Z(n31375) );
  NANDN U40268 ( .A(n31388), .B(n31389), .Z(n31387) );
  OR U40269 ( .A(n31390), .B(n31391), .Z(n31389) );
  NAND U40270 ( .A(n31391), .B(n31390), .Z(n31386) );
  AND U40271 ( .A(n31392), .B(n31393), .Z(n31377) );
  NANDN U40272 ( .A(n31394), .B(n31395), .Z(n31393) );
  NANDN U40273 ( .A(n31396), .B(n31397), .Z(n31395) );
  NANDN U40274 ( .A(n31397), .B(n31396), .Z(n31392) );
  XOR U40275 ( .A(n31391), .B(n31398), .Z(N62609) );
  XOR U40276 ( .A(n31388), .B(n31390), .Z(n31398) );
  XNOR U40277 ( .A(n31384), .B(n31399), .Z(n31390) );
  XNOR U40278 ( .A(n31382), .B(n31385), .Z(n31399) );
  NAND U40279 ( .A(n31400), .B(n31401), .Z(n31385) );
  NAND U40280 ( .A(n31402), .B(n31403), .Z(n31401) );
  OR U40281 ( .A(n31404), .B(n31405), .Z(n31402) );
  NANDN U40282 ( .A(n31406), .B(n31404), .Z(n31400) );
  IV U40283 ( .A(n31405), .Z(n31406) );
  NAND U40284 ( .A(n31407), .B(n31408), .Z(n31382) );
  NAND U40285 ( .A(n31409), .B(n31410), .Z(n31408) );
  NANDN U40286 ( .A(n31411), .B(n31412), .Z(n31409) );
  NANDN U40287 ( .A(n31412), .B(n31411), .Z(n31407) );
  AND U40288 ( .A(n31413), .B(n31414), .Z(n31384) );
  NAND U40289 ( .A(n31415), .B(n31416), .Z(n31414) );
  OR U40290 ( .A(n31417), .B(n31418), .Z(n31415) );
  NANDN U40291 ( .A(n31419), .B(n31417), .Z(n31413) );
  NAND U40292 ( .A(n31420), .B(n31421), .Z(n31388) );
  NANDN U40293 ( .A(n31422), .B(n31423), .Z(n31421) );
  OR U40294 ( .A(n31424), .B(n31425), .Z(n31423) );
  NANDN U40295 ( .A(n31426), .B(n31424), .Z(n31420) );
  IV U40296 ( .A(n31425), .Z(n31426) );
  XNOR U40297 ( .A(n31396), .B(n31427), .Z(n31391) );
  XNOR U40298 ( .A(n31394), .B(n31397), .Z(n31427) );
  NAND U40299 ( .A(n31428), .B(n31429), .Z(n31397) );
  NAND U40300 ( .A(n31430), .B(n31431), .Z(n31429) );
  OR U40301 ( .A(n31432), .B(n31433), .Z(n31430) );
  NANDN U40302 ( .A(n31434), .B(n31432), .Z(n31428) );
  IV U40303 ( .A(n31433), .Z(n31434) );
  NAND U40304 ( .A(n31435), .B(n31436), .Z(n31394) );
  NAND U40305 ( .A(n31437), .B(n31438), .Z(n31436) );
  NANDN U40306 ( .A(n31439), .B(n31440), .Z(n31437) );
  NANDN U40307 ( .A(n31440), .B(n31439), .Z(n31435) );
  AND U40308 ( .A(n31441), .B(n31442), .Z(n31396) );
  NAND U40309 ( .A(n31443), .B(n31444), .Z(n31442) );
  OR U40310 ( .A(n31445), .B(n31446), .Z(n31443) );
  NANDN U40311 ( .A(n31447), .B(n31445), .Z(n31441) );
  XNOR U40312 ( .A(n31422), .B(n31448), .Z(N62608) );
  XOR U40313 ( .A(n31424), .B(n31425), .Z(n31448) );
  XNOR U40314 ( .A(n31438), .B(n31449), .Z(n31425) );
  XOR U40315 ( .A(n31439), .B(n31440), .Z(n31449) );
  XOR U40316 ( .A(n31445), .B(n31450), .Z(n31440) );
  XOR U40317 ( .A(n31444), .B(n31447), .Z(n31450) );
  IV U40318 ( .A(n31446), .Z(n31447) );
  NAND U40319 ( .A(n31451), .B(n31452), .Z(n31446) );
  OR U40320 ( .A(n31453), .B(n31454), .Z(n31452) );
  OR U40321 ( .A(n31455), .B(n31456), .Z(n31451) );
  NAND U40322 ( .A(n31457), .B(n31458), .Z(n31444) );
  OR U40323 ( .A(n31459), .B(n31460), .Z(n31458) );
  OR U40324 ( .A(n31461), .B(n31462), .Z(n31457) );
  NOR U40325 ( .A(n31463), .B(n31464), .Z(n31445) );
  ANDN U40326 ( .B(n31465), .A(n31466), .Z(n31439) );
  XNOR U40327 ( .A(n31432), .B(n31467), .Z(n31438) );
  XNOR U40328 ( .A(n31431), .B(n31433), .Z(n31467) );
  NAND U40329 ( .A(n31468), .B(n31469), .Z(n31433) );
  OR U40330 ( .A(n31470), .B(n31471), .Z(n31469) );
  OR U40331 ( .A(n31472), .B(n31473), .Z(n31468) );
  NAND U40332 ( .A(n31474), .B(n31475), .Z(n31431) );
  OR U40333 ( .A(n31476), .B(n31477), .Z(n31475) );
  OR U40334 ( .A(n31478), .B(n31479), .Z(n31474) );
  ANDN U40335 ( .B(n31480), .A(n31481), .Z(n31432) );
  IV U40336 ( .A(n31482), .Z(n31480) );
  ANDN U40337 ( .B(n31483), .A(n31484), .Z(n31424) );
  XOR U40338 ( .A(n31410), .B(n31485), .Z(n31422) );
  XOR U40339 ( .A(n31411), .B(n31412), .Z(n31485) );
  XOR U40340 ( .A(n31417), .B(n31486), .Z(n31412) );
  XOR U40341 ( .A(n31416), .B(n31419), .Z(n31486) );
  IV U40342 ( .A(n31418), .Z(n31419) );
  NAND U40343 ( .A(n31487), .B(n31488), .Z(n31418) );
  OR U40344 ( .A(n31489), .B(n31490), .Z(n31488) );
  OR U40345 ( .A(n31491), .B(n31492), .Z(n31487) );
  NAND U40346 ( .A(n31493), .B(n31494), .Z(n31416) );
  OR U40347 ( .A(n31495), .B(n31496), .Z(n31494) );
  OR U40348 ( .A(n31497), .B(n31498), .Z(n31493) );
  NOR U40349 ( .A(n31499), .B(n31500), .Z(n31417) );
  ANDN U40350 ( .B(n31501), .A(n31502), .Z(n31411) );
  IV U40351 ( .A(n31503), .Z(n31501) );
  XNOR U40352 ( .A(n31404), .B(n31504), .Z(n31410) );
  XNOR U40353 ( .A(n31403), .B(n31405), .Z(n31504) );
  NAND U40354 ( .A(n31505), .B(n31506), .Z(n31405) );
  OR U40355 ( .A(n31507), .B(n31508), .Z(n31506) );
  OR U40356 ( .A(n31509), .B(n31510), .Z(n31505) );
  NAND U40357 ( .A(n31511), .B(n31512), .Z(n31403) );
  OR U40358 ( .A(n31513), .B(n31514), .Z(n31512) );
  OR U40359 ( .A(n31515), .B(n31516), .Z(n31511) );
  ANDN U40360 ( .B(n31517), .A(n31518), .Z(n31404) );
  IV U40361 ( .A(n31519), .Z(n31517) );
  XNOR U40362 ( .A(n31484), .B(n31483), .Z(N62607) );
  XOR U40363 ( .A(n31503), .B(n31502), .Z(n31483) );
  XNOR U40364 ( .A(n31518), .B(n31519), .Z(n31502) );
  XNOR U40365 ( .A(n31513), .B(n31514), .Z(n31519) );
  XNOR U40366 ( .A(n31515), .B(n31516), .Z(n31514) );
  XNOR U40367 ( .A(y[3733]), .B(x[3733]), .Z(n31516) );
  XNOR U40368 ( .A(y[3734]), .B(x[3734]), .Z(n31515) );
  XNOR U40369 ( .A(y[3732]), .B(x[3732]), .Z(n31513) );
  XNOR U40370 ( .A(n31507), .B(n31508), .Z(n31518) );
  XNOR U40371 ( .A(y[3729]), .B(x[3729]), .Z(n31508) );
  XNOR U40372 ( .A(n31509), .B(n31510), .Z(n31507) );
  XNOR U40373 ( .A(y[3730]), .B(x[3730]), .Z(n31510) );
  XNOR U40374 ( .A(y[3731]), .B(x[3731]), .Z(n31509) );
  XNOR U40375 ( .A(n31500), .B(n31499), .Z(n31503) );
  XNOR U40376 ( .A(n31495), .B(n31496), .Z(n31499) );
  XNOR U40377 ( .A(y[3726]), .B(x[3726]), .Z(n31496) );
  XNOR U40378 ( .A(n31497), .B(n31498), .Z(n31495) );
  XNOR U40379 ( .A(y[3727]), .B(x[3727]), .Z(n31498) );
  XNOR U40380 ( .A(y[3728]), .B(x[3728]), .Z(n31497) );
  XNOR U40381 ( .A(n31489), .B(n31490), .Z(n31500) );
  XNOR U40382 ( .A(y[3723]), .B(x[3723]), .Z(n31490) );
  XNOR U40383 ( .A(n31491), .B(n31492), .Z(n31489) );
  XNOR U40384 ( .A(y[3724]), .B(x[3724]), .Z(n31492) );
  XNOR U40385 ( .A(y[3725]), .B(x[3725]), .Z(n31491) );
  XOR U40386 ( .A(n31465), .B(n31466), .Z(n31484) );
  XNOR U40387 ( .A(n31481), .B(n31482), .Z(n31466) );
  XNOR U40388 ( .A(n31476), .B(n31477), .Z(n31482) );
  XNOR U40389 ( .A(n31478), .B(n31479), .Z(n31477) );
  XNOR U40390 ( .A(y[3721]), .B(x[3721]), .Z(n31479) );
  XNOR U40391 ( .A(y[3722]), .B(x[3722]), .Z(n31478) );
  XNOR U40392 ( .A(y[3720]), .B(x[3720]), .Z(n31476) );
  XNOR U40393 ( .A(n31470), .B(n31471), .Z(n31481) );
  XNOR U40394 ( .A(y[3717]), .B(x[3717]), .Z(n31471) );
  XNOR U40395 ( .A(n31472), .B(n31473), .Z(n31470) );
  XNOR U40396 ( .A(y[3718]), .B(x[3718]), .Z(n31473) );
  XNOR U40397 ( .A(y[3719]), .B(x[3719]), .Z(n31472) );
  XOR U40398 ( .A(n31464), .B(n31463), .Z(n31465) );
  XNOR U40399 ( .A(n31459), .B(n31460), .Z(n31463) );
  XNOR U40400 ( .A(y[3714]), .B(x[3714]), .Z(n31460) );
  XNOR U40401 ( .A(n31461), .B(n31462), .Z(n31459) );
  XNOR U40402 ( .A(y[3715]), .B(x[3715]), .Z(n31462) );
  XNOR U40403 ( .A(y[3716]), .B(x[3716]), .Z(n31461) );
  XNOR U40404 ( .A(n31453), .B(n31454), .Z(n31464) );
  XNOR U40405 ( .A(y[3711]), .B(x[3711]), .Z(n31454) );
  XNOR U40406 ( .A(n31455), .B(n31456), .Z(n31453) );
  XNOR U40407 ( .A(y[3712]), .B(x[3712]), .Z(n31456) );
  XNOR U40408 ( .A(y[3713]), .B(x[3713]), .Z(n31455) );
  NAND U40409 ( .A(n31520), .B(n31521), .Z(N62598) );
  NANDN U40410 ( .A(n31522), .B(n31523), .Z(n31521) );
  OR U40411 ( .A(n31524), .B(n31525), .Z(n31523) );
  NAND U40412 ( .A(n31524), .B(n31525), .Z(n31520) );
  XOR U40413 ( .A(n31524), .B(n31526), .Z(N62597) );
  XNOR U40414 ( .A(n31522), .B(n31525), .Z(n31526) );
  AND U40415 ( .A(n31527), .B(n31528), .Z(n31525) );
  NANDN U40416 ( .A(n31529), .B(n31530), .Z(n31528) );
  NANDN U40417 ( .A(n31531), .B(n31532), .Z(n31530) );
  NANDN U40418 ( .A(n31532), .B(n31531), .Z(n31527) );
  NAND U40419 ( .A(n31533), .B(n31534), .Z(n31522) );
  NANDN U40420 ( .A(n31535), .B(n31536), .Z(n31534) );
  OR U40421 ( .A(n31537), .B(n31538), .Z(n31536) );
  NAND U40422 ( .A(n31538), .B(n31537), .Z(n31533) );
  AND U40423 ( .A(n31539), .B(n31540), .Z(n31524) );
  NANDN U40424 ( .A(n31541), .B(n31542), .Z(n31540) );
  NANDN U40425 ( .A(n31543), .B(n31544), .Z(n31542) );
  NANDN U40426 ( .A(n31544), .B(n31543), .Z(n31539) );
  XOR U40427 ( .A(n31538), .B(n31545), .Z(N62596) );
  XOR U40428 ( .A(n31535), .B(n31537), .Z(n31545) );
  XNOR U40429 ( .A(n31531), .B(n31546), .Z(n31537) );
  XNOR U40430 ( .A(n31529), .B(n31532), .Z(n31546) );
  NAND U40431 ( .A(n31547), .B(n31548), .Z(n31532) );
  NAND U40432 ( .A(n31549), .B(n31550), .Z(n31548) );
  OR U40433 ( .A(n31551), .B(n31552), .Z(n31549) );
  NANDN U40434 ( .A(n31553), .B(n31551), .Z(n31547) );
  IV U40435 ( .A(n31552), .Z(n31553) );
  NAND U40436 ( .A(n31554), .B(n31555), .Z(n31529) );
  NAND U40437 ( .A(n31556), .B(n31557), .Z(n31555) );
  NANDN U40438 ( .A(n31558), .B(n31559), .Z(n31556) );
  NANDN U40439 ( .A(n31559), .B(n31558), .Z(n31554) );
  AND U40440 ( .A(n31560), .B(n31561), .Z(n31531) );
  NAND U40441 ( .A(n31562), .B(n31563), .Z(n31561) );
  OR U40442 ( .A(n31564), .B(n31565), .Z(n31562) );
  NANDN U40443 ( .A(n31566), .B(n31564), .Z(n31560) );
  NAND U40444 ( .A(n31567), .B(n31568), .Z(n31535) );
  NANDN U40445 ( .A(n31569), .B(n31570), .Z(n31568) );
  OR U40446 ( .A(n31571), .B(n31572), .Z(n31570) );
  NANDN U40447 ( .A(n31573), .B(n31571), .Z(n31567) );
  IV U40448 ( .A(n31572), .Z(n31573) );
  XNOR U40449 ( .A(n31543), .B(n31574), .Z(n31538) );
  XNOR U40450 ( .A(n31541), .B(n31544), .Z(n31574) );
  NAND U40451 ( .A(n31575), .B(n31576), .Z(n31544) );
  NAND U40452 ( .A(n31577), .B(n31578), .Z(n31576) );
  OR U40453 ( .A(n31579), .B(n31580), .Z(n31577) );
  NANDN U40454 ( .A(n31581), .B(n31579), .Z(n31575) );
  IV U40455 ( .A(n31580), .Z(n31581) );
  NAND U40456 ( .A(n31582), .B(n31583), .Z(n31541) );
  NAND U40457 ( .A(n31584), .B(n31585), .Z(n31583) );
  NANDN U40458 ( .A(n31586), .B(n31587), .Z(n31584) );
  NANDN U40459 ( .A(n31587), .B(n31586), .Z(n31582) );
  AND U40460 ( .A(n31588), .B(n31589), .Z(n31543) );
  NAND U40461 ( .A(n31590), .B(n31591), .Z(n31589) );
  OR U40462 ( .A(n31592), .B(n31593), .Z(n31590) );
  NANDN U40463 ( .A(n31594), .B(n31592), .Z(n31588) );
  XNOR U40464 ( .A(n31569), .B(n31595), .Z(N62595) );
  XOR U40465 ( .A(n31571), .B(n31572), .Z(n31595) );
  XNOR U40466 ( .A(n31585), .B(n31596), .Z(n31572) );
  XOR U40467 ( .A(n31586), .B(n31587), .Z(n31596) );
  XOR U40468 ( .A(n31592), .B(n31597), .Z(n31587) );
  XOR U40469 ( .A(n31591), .B(n31594), .Z(n31597) );
  IV U40470 ( .A(n31593), .Z(n31594) );
  NAND U40471 ( .A(n31598), .B(n31599), .Z(n31593) );
  OR U40472 ( .A(n31600), .B(n31601), .Z(n31599) );
  OR U40473 ( .A(n31602), .B(n31603), .Z(n31598) );
  NAND U40474 ( .A(n31604), .B(n31605), .Z(n31591) );
  OR U40475 ( .A(n31606), .B(n31607), .Z(n31605) );
  OR U40476 ( .A(n31608), .B(n31609), .Z(n31604) );
  NOR U40477 ( .A(n31610), .B(n31611), .Z(n31592) );
  ANDN U40478 ( .B(n31612), .A(n31613), .Z(n31586) );
  XNOR U40479 ( .A(n31579), .B(n31614), .Z(n31585) );
  XNOR U40480 ( .A(n31578), .B(n31580), .Z(n31614) );
  NAND U40481 ( .A(n31615), .B(n31616), .Z(n31580) );
  OR U40482 ( .A(n31617), .B(n31618), .Z(n31616) );
  OR U40483 ( .A(n31619), .B(n31620), .Z(n31615) );
  NAND U40484 ( .A(n31621), .B(n31622), .Z(n31578) );
  OR U40485 ( .A(n31623), .B(n31624), .Z(n31622) );
  OR U40486 ( .A(n31625), .B(n31626), .Z(n31621) );
  ANDN U40487 ( .B(n31627), .A(n31628), .Z(n31579) );
  IV U40488 ( .A(n31629), .Z(n31627) );
  ANDN U40489 ( .B(n31630), .A(n31631), .Z(n31571) );
  XOR U40490 ( .A(n31557), .B(n31632), .Z(n31569) );
  XOR U40491 ( .A(n31558), .B(n31559), .Z(n31632) );
  XOR U40492 ( .A(n31564), .B(n31633), .Z(n31559) );
  XOR U40493 ( .A(n31563), .B(n31566), .Z(n31633) );
  IV U40494 ( .A(n31565), .Z(n31566) );
  NAND U40495 ( .A(n31634), .B(n31635), .Z(n31565) );
  OR U40496 ( .A(n31636), .B(n31637), .Z(n31635) );
  OR U40497 ( .A(n31638), .B(n31639), .Z(n31634) );
  NAND U40498 ( .A(n31640), .B(n31641), .Z(n31563) );
  OR U40499 ( .A(n31642), .B(n31643), .Z(n31641) );
  OR U40500 ( .A(n31644), .B(n31645), .Z(n31640) );
  NOR U40501 ( .A(n31646), .B(n31647), .Z(n31564) );
  ANDN U40502 ( .B(n31648), .A(n31649), .Z(n31558) );
  IV U40503 ( .A(n31650), .Z(n31648) );
  XNOR U40504 ( .A(n31551), .B(n31651), .Z(n31557) );
  XNOR U40505 ( .A(n31550), .B(n31552), .Z(n31651) );
  NAND U40506 ( .A(n31652), .B(n31653), .Z(n31552) );
  OR U40507 ( .A(n31654), .B(n31655), .Z(n31653) );
  OR U40508 ( .A(n31656), .B(n31657), .Z(n31652) );
  NAND U40509 ( .A(n31658), .B(n31659), .Z(n31550) );
  OR U40510 ( .A(n31660), .B(n31661), .Z(n31659) );
  OR U40511 ( .A(n31662), .B(n31663), .Z(n31658) );
  ANDN U40512 ( .B(n31664), .A(n31665), .Z(n31551) );
  IV U40513 ( .A(n31666), .Z(n31664) );
  XNOR U40514 ( .A(n31631), .B(n31630), .Z(N62594) );
  XOR U40515 ( .A(n31650), .B(n31649), .Z(n31630) );
  XNOR U40516 ( .A(n31665), .B(n31666), .Z(n31649) );
  XNOR U40517 ( .A(n31660), .B(n31661), .Z(n31666) );
  XNOR U40518 ( .A(n31662), .B(n31663), .Z(n31661) );
  XNOR U40519 ( .A(y[3709]), .B(x[3709]), .Z(n31663) );
  XNOR U40520 ( .A(y[3710]), .B(x[3710]), .Z(n31662) );
  XNOR U40521 ( .A(y[3708]), .B(x[3708]), .Z(n31660) );
  XNOR U40522 ( .A(n31654), .B(n31655), .Z(n31665) );
  XNOR U40523 ( .A(y[3705]), .B(x[3705]), .Z(n31655) );
  XNOR U40524 ( .A(n31656), .B(n31657), .Z(n31654) );
  XNOR U40525 ( .A(y[3706]), .B(x[3706]), .Z(n31657) );
  XNOR U40526 ( .A(y[3707]), .B(x[3707]), .Z(n31656) );
  XNOR U40527 ( .A(n31647), .B(n31646), .Z(n31650) );
  XNOR U40528 ( .A(n31642), .B(n31643), .Z(n31646) );
  XNOR U40529 ( .A(y[3702]), .B(x[3702]), .Z(n31643) );
  XNOR U40530 ( .A(n31644), .B(n31645), .Z(n31642) );
  XNOR U40531 ( .A(y[3703]), .B(x[3703]), .Z(n31645) );
  XNOR U40532 ( .A(y[3704]), .B(x[3704]), .Z(n31644) );
  XNOR U40533 ( .A(n31636), .B(n31637), .Z(n31647) );
  XNOR U40534 ( .A(y[3699]), .B(x[3699]), .Z(n31637) );
  XNOR U40535 ( .A(n31638), .B(n31639), .Z(n31636) );
  XNOR U40536 ( .A(y[3700]), .B(x[3700]), .Z(n31639) );
  XNOR U40537 ( .A(y[3701]), .B(x[3701]), .Z(n31638) );
  XOR U40538 ( .A(n31612), .B(n31613), .Z(n31631) );
  XNOR U40539 ( .A(n31628), .B(n31629), .Z(n31613) );
  XNOR U40540 ( .A(n31623), .B(n31624), .Z(n31629) );
  XNOR U40541 ( .A(n31625), .B(n31626), .Z(n31624) );
  XNOR U40542 ( .A(y[3697]), .B(x[3697]), .Z(n31626) );
  XNOR U40543 ( .A(y[3698]), .B(x[3698]), .Z(n31625) );
  XNOR U40544 ( .A(y[3696]), .B(x[3696]), .Z(n31623) );
  XNOR U40545 ( .A(n31617), .B(n31618), .Z(n31628) );
  XNOR U40546 ( .A(y[3693]), .B(x[3693]), .Z(n31618) );
  XNOR U40547 ( .A(n31619), .B(n31620), .Z(n31617) );
  XNOR U40548 ( .A(y[3694]), .B(x[3694]), .Z(n31620) );
  XNOR U40549 ( .A(y[3695]), .B(x[3695]), .Z(n31619) );
  XOR U40550 ( .A(n31611), .B(n31610), .Z(n31612) );
  XNOR U40551 ( .A(n31606), .B(n31607), .Z(n31610) );
  XNOR U40552 ( .A(y[3690]), .B(x[3690]), .Z(n31607) );
  XNOR U40553 ( .A(n31608), .B(n31609), .Z(n31606) );
  XNOR U40554 ( .A(y[3691]), .B(x[3691]), .Z(n31609) );
  XNOR U40555 ( .A(y[3692]), .B(x[3692]), .Z(n31608) );
  XNOR U40556 ( .A(n31600), .B(n31601), .Z(n31611) );
  XNOR U40557 ( .A(y[3687]), .B(x[3687]), .Z(n31601) );
  XNOR U40558 ( .A(n31602), .B(n31603), .Z(n31600) );
  XNOR U40559 ( .A(y[3688]), .B(x[3688]), .Z(n31603) );
  XNOR U40560 ( .A(y[3689]), .B(x[3689]), .Z(n31602) );
  NAND U40561 ( .A(n31667), .B(n31668), .Z(N62585) );
  NANDN U40562 ( .A(n31669), .B(n31670), .Z(n31668) );
  OR U40563 ( .A(n31671), .B(n31672), .Z(n31670) );
  NAND U40564 ( .A(n31671), .B(n31672), .Z(n31667) );
  XOR U40565 ( .A(n31671), .B(n31673), .Z(N62584) );
  XNOR U40566 ( .A(n31669), .B(n31672), .Z(n31673) );
  AND U40567 ( .A(n31674), .B(n31675), .Z(n31672) );
  NANDN U40568 ( .A(n31676), .B(n31677), .Z(n31675) );
  NANDN U40569 ( .A(n31678), .B(n31679), .Z(n31677) );
  NANDN U40570 ( .A(n31679), .B(n31678), .Z(n31674) );
  NAND U40571 ( .A(n31680), .B(n31681), .Z(n31669) );
  NANDN U40572 ( .A(n31682), .B(n31683), .Z(n31681) );
  OR U40573 ( .A(n31684), .B(n31685), .Z(n31683) );
  NAND U40574 ( .A(n31685), .B(n31684), .Z(n31680) );
  AND U40575 ( .A(n31686), .B(n31687), .Z(n31671) );
  NANDN U40576 ( .A(n31688), .B(n31689), .Z(n31687) );
  NANDN U40577 ( .A(n31690), .B(n31691), .Z(n31689) );
  NANDN U40578 ( .A(n31691), .B(n31690), .Z(n31686) );
  XOR U40579 ( .A(n31685), .B(n31692), .Z(N62583) );
  XOR U40580 ( .A(n31682), .B(n31684), .Z(n31692) );
  XNOR U40581 ( .A(n31678), .B(n31693), .Z(n31684) );
  XNOR U40582 ( .A(n31676), .B(n31679), .Z(n31693) );
  NAND U40583 ( .A(n31694), .B(n31695), .Z(n31679) );
  NAND U40584 ( .A(n31696), .B(n31697), .Z(n31695) );
  OR U40585 ( .A(n31698), .B(n31699), .Z(n31696) );
  NANDN U40586 ( .A(n31700), .B(n31698), .Z(n31694) );
  IV U40587 ( .A(n31699), .Z(n31700) );
  NAND U40588 ( .A(n31701), .B(n31702), .Z(n31676) );
  NAND U40589 ( .A(n31703), .B(n31704), .Z(n31702) );
  NANDN U40590 ( .A(n31705), .B(n31706), .Z(n31703) );
  NANDN U40591 ( .A(n31706), .B(n31705), .Z(n31701) );
  AND U40592 ( .A(n31707), .B(n31708), .Z(n31678) );
  NAND U40593 ( .A(n31709), .B(n31710), .Z(n31708) );
  OR U40594 ( .A(n31711), .B(n31712), .Z(n31709) );
  NANDN U40595 ( .A(n31713), .B(n31711), .Z(n31707) );
  NAND U40596 ( .A(n31714), .B(n31715), .Z(n31682) );
  NANDN U40597 ( .A(n31716), .B(n31717), .Z(n31715) );
  OR U40598 ( .A(n31718), .B(n31719), .Z(n31717) );
  NANDN U40599 ( .A(n31720), .B(n31718), .Z(n31714) );
  IV U40600 ( .A(n31719), .Z(n31720) );
  XNOR U40601 ( .A(n31690), .B(n31721), .Z(n31685) );
  XNOR U40602 ( .A(n31688), .B(n31691), .Z(n31721) );
  NAND U40603 ( .A(n31722), .B(n31723), .Z(n31691) );
  NAND U40604 ( .A(n31724), .B(n31725), .Z(n31723) );
  OR U40605 ( .A(n31726), .B(n31727), .Z(n31724) );
  NANDN U40606 ( .A(n31728), .B(n31726), .Z(n31722) );
  IV U40607 ( .A(n31727), .Z(n31728) );
  NAND U40608 ( .A(n31729), .B(n31730), .Z(n31688) );
  NAND U40609 ( .A(n31731), .B(n31732), .Z(n31730) );
  NANDN U40610 ( .A(n31733), .B(n31734), .Z(n31731) );
  NANDN U40611 ( .A(n31734), .B(n31733), .Z(n31729) );
  AND U40612 ( .A(n31735), .B(n31736), .Z(n31690) );
  NAND U40613 ( .A(n31737), .B(n31738), .Z(n31736) );
  OR U40614 ( .A(n31739), .B(n31740), .Z(n31737) );
  NANDN U40615 ( .A(n31741), .B(n31739), .Z(n31735) );
  XNOR U40616 ( .A(n31716), .B(n31742), .Z(N62582) );
  XOR U40617 ( .A(n31718), .B(n31719), .Z(n31742) );
  XNOR U40618 ( .A(n31732), .B(n31743), .Z(n31719) );
  XOR U40619 ( .A(n31733), .B(n31734), .Z(n31743) );
  XOR U40620 ( .A(n31739), .B(n31744), .Z(n31734) );
  XOR U40621 ( .A(n31738), .B(n31741), .Z(n31744) );
  IV U40622 ( .A(n31740), .Z(n31741) );
  NAND U40623 ( .A(n31745), .B(n31746), .Z(n31740) );
  OR U40624 ( .A(n31747), .B(n31748), .Z(n31746) );
  OR U40625 ( .A(n31749), .B(n31750), .Z(n31745) );
  NAND U40626 ( .A(n31751), .B(n31752), .Z(n31738) );
  OR U40627 ( .A(n31753), .B(n31754), .Z(n31752) );
  OR U40628 ( .A(n31755), .B(n31756), .Z(n31751) );
  NOR U40629 ( .A(n31757), .B(n31758), .Z(n31739) );
  ANDN U40630 ( .B(n31759), .A(n31760), .Z(n31733) );
  XNOR U40631 ( .A(n31726), .B(n31761), .Z(n31732) );
  XNOR U40632 ( .A(n31725), .B(n31727), .Z(n31761) );
  NAND U40633 ( .A(n31762), .B(n31763), .Z(n31727) );
  OR U40634 ( .A(n31764), .B(n31765), .Z(n31763) );
  OR U40635 ( .A(n31766), .B(n31767), .Z(n31762) );
  NAND U40636 ( .A(n31768), .B(n31769), .Z(n31725) );
  OR U40637 ( .A(n31770), .B(n31771), .Z(n31769) );
  OR U40638 ( .A(n31772), .B(n31773), .Z(n31768) );
  ANDN U40639 ( .B(n31774), .A(n31775), .Z(n31726) );
  IV U40640 ( .A(n31776), .Z(n31774) );
  ANDN U40641 ( .B(n31777), .A(n31778), .Z(n31718) );
  XOR U40642 ( .A(n31704), .B(n31779), .Z(n31716) );
  XOR U40643 ( .A(n31705), .B(n31706), .Z(n31779) );
  XOR U40644 ( .A(n31711), .B(n31780), .Z(n31706) );
  XOR U40645 ( .A(n31710), .B(n31713), .Z(n31780) );
  IV U40646 ( .A(n31712), .Z(n31713) );
  NAND U40647 ( .A(n31781), .B(n31782), .Z(n31712) );
  OR U40648 ( .A(n31783), .B(n31784), .Z(n31782) );
  OR U40649 ( .A(n31785), .B(n31786), .Z(n31781) );
  NAND U40650 ( .A(n31787), .B(n31788), .Z(n31710) );
  OR U40651 ( .A(n31789), .B(n31790), .Z(n31788) );
  OR U40652 ( .A(n31791), .B(n31792), .Z(n31787) );
  NOR U40653 ( .A(n31793), .B(n31794), .Z(n31711) );
  ANDN U40654 ( .B(n31795), .A(n31796), .Z(n31705) );
  IV U40655 ( .A(n31797), .Z(n31795) );
  XNOR U40656 ( .A(n31698), .B(n31798), .Z(n31704) );
  XNOR U40657 ( .A(n31697), .B(n31699), .Z(n31798) );
  NAND U40658 ( .A(n31799), .B(n31800), .Z(n31699) );
  OR U40659 ( .A(n31801), .B(n31802), .Z(n31800) );
  OR U40660 ( .A(n31803), .B(n31804), .Z(n31799) );
  NAND U40661 ( .A(n31805), .B(n31806), .Z(n31697) );
  OR U40662 ( .A(n31807), .B(n31808), .Z(n31806) );
  OR U40663 ( .A(n31809), .B(n31810), .Z(n31805) );
  ANDN U40664 ( .B(n31811), .A(n31812), .Z(n31698) );
  IV U40665 ( .A(n31813), .Z(n31811) );
  XNOR U40666 ( .A(n31778), .B(n31777), .Z(N62581) );
  XOR U40667 ( .A(n31797), .B(n31796), .Z(n31777) );
  XNOR U40668 ( .A(n31812), .B(n31813), .Z(n31796) );
  XNOR U40669 ( .A(n31807), .B(n31808), .Z(n31813) );
  XNOR U40670 ( .A(n31809), .B(n31810), .Z(n31808) );
  XNOR U40671 ( .A(y[3685]), .B(x[3685]), .Z(n31810) );
  XNOR U40672 ( .A(y[3686]), .B(x[3686]), .Z(n31809) );
  XNOR U40673 ( .A(y[3684]), .B(x[3684]), .Z(n31807) );
  XNOR U40674 ( .A(n31801), .B(n31802), .Z(n31812) );
  XNOR U40675 ( .A(y[3681]), .B(x[3681]), .Z(n31802) );
  XNOR U40676 ( .A(n31803), .B(n31804), .Z(n31801) );
  XNOR U40677 ( .A(y[3682]), .B(x[3682]), .Z(n31804) );
  XNOR U40678 ( .A(y[3683]), .B(x[3683]), .Z(n31803) );
  XNOR U40679 ( .A(n31794), .B(n31793), .Z(n31797) );
  XNOR U40680 ( .A(n31789), .B(n31790), .Z(n31793) );
  XNOR U40681 ( .A(y[3678]), .B(x[3678]), .Z(n31790) );
  XNOR U40682 ( .A(n31791), .B(n31792), .Z(n31789) );
  XNOR U40683 ( .A(y[3679]), .B(x[3679]), .Z(n31792) );
  XNOR U40684 ( .A(y[3680]), .B(x[3680]), .Z(n31791) );
  XNOR U40685 ( .A(n31783), .B(n31784), .Z(n31794) );
  XNOR U40686 ( .A(y[3675]), .B(x[3675]), .Z(n31784) );
  XNOR U40687 ( .A(n31785), .B(n31786), .Z(n31783) );
  XNOR U40688 ( .A(y[3676]), .B(x[3676]), .Z(n31786) );
  XNOR U40689 ( .A(y[3677]), .B(x[3677]), .Z(n31785) );
  XOR U40690 ( .A(n31759), .B(n31760), .Z(n31778) );
  XNOR U40691 ( .A(n31775), .B(n31776), .Z(n31760) );
  XNOR U40692 ( .A(n31770), .B(n31771), .Z(n31776) );
  XNOR U40693 ( .A(n31772), .B(n31773), .Z(n31771) );
  XNOR U40694 ( .A(y[3673]), .B(x[3673]), .Z(n31773) );
  XNOR U40695 ( .A(y[3674]), .B(x[3674]), .Z(n31772) );
  XNOR U40696 ( .A(y[3672]), .B(x[3672]), .Z(n31770) );
  XNOR U40697 ( .A(n31764), .B(n31765), .Z(n31775) );
  XNOR U40698 ( .A(y[3669]), .B(x[3669]), .Z(n31765) );
  XNOR U40699 ( .A(n31766), .B(n31767), .Z(n31764) );
  XNOR U40700 ( .A(y[3670]), .B(x[3670]), .Z(n31767) );
  XNOR U40701 ( .A(y[3671]), .B(x[3671]), .Z(n31766) );
  XOR U40702 ( .A(n31758), .B(n31757), .Z(n31759) );
  XNOR U40703 ( .A(n31753), .B(n31754), .Z(n31757) );
  XNOR U40704 ( .A(y[3666]), .B(x[3666]), .Z(n31754) );
  XNOR U40705 ( .A(n31755), .B(n31756), .Z(n31753) );
  XNOR U40706 ( .A(y[3667]), .B(x[3667]), .Z(n31756) );
  XNOR U40707 ( .A(y[3668]), .B(x[3668]), .Z(n31755) );
  XNOR U40708 ( .A(n31747), .B(n31748), .Z(n31758) );
  XNOR U40709 ( .A(y[3663]), .B(x[3663]), .Z(n31748) );
  XNOR U40710 ( .A(n31749), .B(n31750), .Z(n31747) );
  XNOR U40711 ( .A(y[3664]), .B(x[3664]), .Z(n31750) );
  XNOR U40712 ( .A(y[3665]), .B(x[3665]), .Z(n31749) );
  NAND U40713 ( .A(n31814), .B(n31815), .Z(N62572) );
  NANDN U40714 ( .A(n31816), .B(n31817), .Z(n31815) );
  OR U40715 ( .A(n31818), .B(n31819), .Z(n31817) );
  NAND U40716 ( .A(n31818), .B(n31819), .Z(n31814) );
  XOR U40717 ( .A(n31818), .B(n31820), .Z(N62571) );
  XNOR U40718 ( .A(n31816), .B(n31819), .Z(n31820) );
  AND U40719 ( .A(n31821), .B(n31822), .Z(n31819) );
  NANDN U40720 ( .A(n31823), .B(n31824), .Z(n31822) );
  NANDN U40721 ( .A(n31825), .B(n31826), .Z(n31824) );
  NANDN U40722 ( .A(n31826), .B(n31825), .Z(n31821) );
  NAND U40723 ( .A(n31827), .B(n31828), .Z(n31816) );
  NANDN U40724 ( .A(n31829), .B(n31830), .Z(n31828) );
  OR U40725 ( .A(n31831), .B(n31832), .Z(n31830) );
  NAND U40726 ( .A(n31832), .B(n31831), .Z(n31827) );
  AND U40727 ( .A(n31833), .B(n31834), .Z(n31818) );
  NANDN U40728 ( .A(n31835), .B(n31836), .Z(n31834) );
  NANDN U40729 ( .A(n31837), .B(n31838), .Z(n31836) );
  NANDN U40730 ( .A(n31838), .B(n31837), .Z(n31833) );
  XOR U40731 ( .A(n31832), .B(n31839), .Z(N62570) );
  XOR U40732 ( .A(n31829), .B(n31831), .Z(n31839) );
  XNOR U40733 ( .A(n31825), .B(n31840), .Z(n31831) );
  XNOR U40734 ( .A(n31823), .B(n31826), .Z(n31840) );
  NAND U40735 ( .A(n31841), .B(n31842), .Z(n31826) );
  NAND U40736 ( .A(n31843), .B(n31844), .Z(n31842) );
  OR U40737 ( .A(n31845), .B(n31846), .Z(n31843) );
  NANDN U40738 ( .A(n31847), .B(n31845), .Z(n31841) );
  IV U40739 ( .A(n31846), .Z(n31847) );
  NAND U40740 ( .A(n31848), .B(n31849), .Z(n31823) );
  NAND U40741 ( .A(n31850), .B(n31851), .Z(n31849) );
  NANDN U40742 ( .A(n31852), .B(n31853), .Z(n31850) );
  NANDN U40743 ( .A(n31853), .B(n31852), .Z(n31848) );
  AND U40744 ( .A(n31854), .B(n31855), .Z(n31825) );
  NAND U40745 ( .A(n31856), .B(n31857), .Z(n31855) );
  OR U40746 ( .A(n31858), .B(n31859), .Z(n31856) );
  NANDN U40747 ( .A(n31860), .B(n31858), .Z(n31854) );
  NAND U40748 ( .A(n31861), .B(n31862), .Z(n31829) );
  NANDN U40749 ( .A(n31863), .B(n31864), .Z(n31862) );
  OR U40750 ( .A(n31865), .B(n31866), .Z(n31864) );
  NANDN U40751 ( .A(n31867), .B(n31865), .Z(n31861) );
  IV U40752 ( .A(n31866), .Z(n31867) );
  XNOR U40753 ( .A(n31837), .B(n31868), .Z(n31832) );
  XNOR U40754 ( .A(n31835), .B(n31838), .Z(n31868) );
  NAND U40755 ( .A(n31869), .B(n31870), .Z(n31838) );
  NAND U40756 ( .A(n31871), .B(n31872), .Z(n31870) );
  OR U40757 ( .A(n31873), .B(n31874), .Z(n31871) );
  NANDN U40758 ( .A(n31875), .B(n31873), .Z(n31869) );
  IV U40759 ( .A(n31874), .Z(n31875) );
  NAND U40760 ( .A(n31876), .B(n31877), .Z(n31835) );
  NAND U40761 ( .A(n31878), .B(n31879), .Z(n31877) );
  NANDN U40762 ( .A(n31880), .B(n31881), .Z(n31878) );
  NANDN U40763 ( .A(n31881), .B(n31880), .Z(n31876) );
  AND U40764 ( .A(n31882), .B(n31883), .Z(n31837) );
  NAND U40765 ( .A(n31884), .B(n31885), .Z(n31883) );
  OR U40766 ( .A(n31886), .B(n31887), .Z(n31884) );
  NANDN U40767 ( .A(n31888), .B(n31886), .Z(n31882) );
  XNOR U40768 ( .A(n31863), .B(n31889), .Z(N62569) );
  XOR U40769 ( .A(n31865), .B(n31866), .Z(n31889) );
  XNOR U40770 ( .A(n31879), .B(n31890), .Z(n31866) );
  XOR U40771 ( .A(n31880), .B(n31881), .Z(n31890) );
  XOR U40772 ( .A(n31886), .B(n31891), .Z(n31881) );
  XOR U40773 ( .A(n31885), .B(n31888), .Z(n31891) );
  IV U40774 ( .A(n31887), .Z(n31888) );
  NAND U40775 ( .A(n31892), .B(n31893), .Z(n31887) );
  OR U40776 ( .A(n31894), .B(n31895), .Z(n31893) );
  OR U40777 ( .A(n31896), .B(n31897), .Z(n31892) );
  NAND U40778 ( .A(n31898), .B(n31899), .Z(n31885) );
  OR U40779 ( .A(n31900), .B(n31901), .Z(n31899) );
  OR U40780 ( .A(n31902), .B(n31903), .Z(n31898) );
  NOR U40781 ( .A(n31904), .B(n31905), .Z(n31886) );
  ANDN U40782 ( .B(n31906), .A(n31907), .Z(n31880) );
  XNOR U40783 ( .A(n31873), .B(n31908), .Z(n31879) );
  XNOR U40784 ( .A(n31872), .B(n31874), .Z(n31908) );
  NAND U40785 ( .A(n31909), .B(n31910), .Z(n31874) );
  OR U40786 ( .A(n31911), .B(n31912), .Z(n31910) );
  OR U40787 ( .A(n31913), .B(n31914), .Z(n31909) );
  NAND U40788 ( .A(n31915), .B(n31916), .Z(n31872) );
  OR U40789 ( .A(n31917), .B(n31918), .Z(n31916) );
  OR U40790 ( .A(n31919), .B(n31920), .Z(n31915) );
  ANDN U40791 ( .B(n31921), .A(n31922), .Z(n31873) );
  IV U40792 ( .A(n31923), .Z(n31921) );
  ANDN U40793 ( .B(n31924), .A(n31925), .Z(n31865) );
  XOR U40794 ( .A(n31851), .B(n31926), .Z(n31863) );
  XOR U40795 ( .A(n31852), .B(n31853), .Z(n31926) );
  XOR U40796 ( .A(n31858), .B(n31927), .Z(n31853) );
  XOR U40797 ( .A(n31857), .B(n31860), .Z(n31927) );
  IV U40798 ( .A(n31859), .Z(n31860) );
  NAND U40799 ( .A(n31928), .B(n31929), .Z(n31859) );
  OR U40800 ( .A(n31930), .B(n31931), .Z(n31929) );
  OR U40801 ( .A(n31932), .B(n31933), .Z(n31928) );
  NAND U40802 ( .A(n31934), .B(n31935), .Z(n31857) );
  OR U40803 ( .A(n31936), .B(n31937), .Z(n31935) );
  OR U40804 ( .A(n31938), .B(n31939), .Z(n31934) );
  NOR U40805 ( .A(n31940), .B(n31941), .Z(n31858) );
  ANDN U40806 ( .B(n31942), .A(n31943), .Z(n31852) );
  IV U40807 ( .A(n31944), .Z(n31942) );
  XNOR U40808 ( .A(n31845), .B(n31945), .Z(n31851) );
  XNOR U40809 ( .A(n31844), .B(n31846), .Z(n31945) );
  NAND U40810 ( .A(n31946), .B(n31947), .Z(n31846) );
  OR U40811 ( .A(n31948), .B(n31949), .Z(n31947) );
  OR U40812 ( .A(n31950), .B(n31951), .Z(n31946) );
  NAND U40813 ( .A(n31952), .B(n31953), .Z(n31844) );
  OR U40814 ( .A(n31954), .B(n31955), .Z(n31953) );
  OR U40815 ( .A(n31956), .B(n31957), .Z(n31952) );
  ANDN U40816 ( .B(n31958), .A(n31959), .Z(n31845) );
  IV U40817 ( .A(n31960), .Z(n31958) );
  XNOR U40818 ( .A(n31925), .B(n31924), .Z(N62568) );
  XOR U40819 ( .A(n31944), .B(n31943), .Z(n31924) );
  XNOR U40820 ( .A(n31959), .B(n31960), .Z(n31943) );
  XNOR U40821 ( .A(n31954), .B(n31955), .Z(n31960) );
  XNOR U40822 ( .A(n31956), .B(n31957), .Z(n31955) );
  XNOR U40823 ( .A(y[3661]), .B(x[3661]), .Z(n31957) );
  XNOR U40824 ( .A(y[3662]), .B(x[3662]), .Z(n31956) );
  XNOR U40825 ( .A(y[3660]), .B(x[3660]), .Z(n31954) );
  XNOR U40826 ( .A(n31948), .B(n31949), .Z(n31959) );
  XNOR U40827 ( .A(y[3657]), .B(x[3657]), .Z(n31949) );
  XNOR U40828 ( .A(n31950), .B(n31951), .Z(n31948) );
  XNOR U40829 ( .A(y[3658]), .B(x[3658]), .Z(n31951) );
  XNOR U40830 ( .A(y[3659]), .B(x[3659]), .Z(n31950) );
  XNOR U40831 ( .A(n31941), .B(n31940), .Z(n31944) );
  XNOR U40832 ( .A(n31936), .B(n31937), .Z(n31940) );
  XNOR U40833 ( .A(y[3654]), .B(x[3654]), .Z(n31937) );
  XNOR U40834 ( .A(n31938), .B(n31939), .Z(n31936) );
  XNOR U40835 ( .A(y[3655]), .B(x[3655]), .Z(n31939) );
  XNOR U40836 ( .A(y[3656]), .B(x[3656]), .Z(n31938) );
  XNOR U40837 ( .A(n31930), .B(n31931), .Z(n31941) );
  XNOR U40838 ( .A(y[3651]), .B(x[3651]), .Z(n31931) );
  XNOR U40839 ( .A(n31932), .B(n31933), .Z(n31930) );
  XNOR U40840 ( .A(y[3652]), .B(x[3652]), .Z(n31933) );
  XNOR U40841 ( .A(y[3653]), .B(x[3653]), .Z(n31932) );
  XOR U40842 ( .A(n31906), .B(n31907), .Z(n31925) );
  XNOR U40843 ( .A(n31922), .B(n31923), .Z(n31907) );
  XNOR U40844 ( .A(n31917), .B(n31918), .Z(n31923) );
  XNOR U40845 ( .A(n31919), .B(n31920), .Z(n31918) );
  XNOR U40846 ( .A(y[3649]), .B(x[3649]), .Z(n31920) );
  XNOR U40847 ( .A(y[3650]), .B(x[3650]), .Z(n31919) );
  XNOR U40848 ( .A(y[3648]), .B(x[3648]), .Z(n31917) );
  XNOR U40849 ( .A(n31911), .B(n31912), .Z(n31922) );
  XNOR U40850 ( .A(y[3645]), .B(x[3645]), .Z(n31912) );
  XNOR U40851 ( .A(n31913), .B(n31914), .Z(n31911) );
  XNOR U40852 ( .A(y[3646]), .B(x[3646]), .Z(n31914) );
  XNOR U40853 ( .A(y[3647]), .B(x[3647]), .Z(n31913) );
  XOR U40854 ( .A(n31905), .B(n31904), .Z(n31906) );
  XNOR U40855 ( .A(n31900), .B(n31901), .Z(n31904) );
  XNOR U40856 ( .A(y[3642]), .B(x[3642]), .Z(n31901) );
  XNOR U40857 ( .A(n31902), .B(n31903), .Z(n31900) );
  XNOR U40858 ( .A(y[3643]), .B(x[3643]), .Z(n31903) );
  XNOR U40859 ( .A(y[3644]), .B(x[3644]), .Z(n31902) );
  XNOR U40860 ( .A(n31894), .B(n31895), .Z(n31905) );
  XNOR U40861 ( .A(y[3639]), .B(x[3639]), .Z(n31895) );
  XNOR U40862 ( .A(n31896), .B(n31897), .Z(n31894) );
  XNOR U40863 ( .A(y[3640]), .B(x[3640]), .Z(n31897) );
  XNOR U40864 ( .A(y[3641]), .B(x[3641]), .Z(n31896) );
  NAND U40865 ( .A(n31961), .B(n31962), .Z(N62559) );
  NANDN U40866 ( .A(n31963), .B(n31964), .Z(n31962) );
  OR U40867 ( .A(n31965), .B(n31966), .Z(n31964) );
  NAND U40868 ( .A(n31965), .B(n31966), .Z(n31961) );
  XOR U40869 ( .A(n31965), .B(n31967), .Z(N62558) );
  XNOR U40870 ( .A(n31963), .B(n31966), .Z(n31967) );
  AND U40871 ( .A(n31968), .B(n31969), .Z(n31966) );
  NANDN U40872 ( .A(n31970), .B(n31971), .Z(n31969) );
  NANDN U40873 ( .A(n31972), .B(n31973), .Z(n31971) );
  NANDN U40874 ( .A(n31973), .B(n31972), .Z(n31968) );
  NAND U40875 ( .A(n31974), .B(n31975), .Z(n31963) );
  NANDN U40876 ( .A(n31976), .B(n31977), .Z(n31975) );
  OR U40877 ( .A(n31978), .B(n31979), .Z(n31977) );
  NAND U40878 ( .A(n31979), .B(n31978), .Z(n31974) );
  AND U40879 ( .A(n31980), .B(n31981), .Z(n31965) );
  NANDN U40880 ( .A(n31982), .B(n31983), .Z(n31981) );
  NANDN U40881 ( .A(n31984), .B(n31985), .Z(n31983) );
  NANDN U40882 ( .A(n31985), .B(n31984), .Z(n31980) );
  XOR U40883 ( .A(n31979), .B(n31986), .Z(N62557) );
  XOR U40884 ( .A(n31976), .B(n31978), .Z(n31986) );
  XNOR U40885 ( .A(n31972), .B(n31987), .Z(n31978) );
  XNOR U40886 ( .A(n31970), .B(n31973), .Z(n31987) );
  NAND U40887 ( .A(n31988), .B(n31989), .Z(n31973) );
  NAND U40888 ( .A(n31990), .B(n31991), .Z(n31989) );
  OR U40889 ( .A(n31992), .B(n31993), .Z(n31990) );
  NANDN U40890 ( .A(n31994), .B(n31992), .Z(n31988) );
  IV U40891 ( .A(n31993), .Z(n31994) );
  NAND U40892 ( .A(n31995), .B(n31996), .Z(n31970) );
  NAND U40893 ( .A(n31997), .B(n31998), .Z(n31996) );
  NANDN U40894 ( .A(n31999), .B(n32000), .Z(n31997) );
  NANDN U40895 ( .A(n32000), .B(n31999), .Z(n31995) );
  AND U40896 ( .A(n32001), .B(n32002), .Z(n31972) );
  NAND U40897 ( .A(n32003), .B(n32004), .Z(n32002) );
  OR U40898 ( .A(n32005), .B(n32006), .Z(n32003) );
  NANDN U40899 ( .A(n32007), .B(n32005), .Z(n32001) );
  NAND U40900 ( .A(n32008), .B(n32009), .Z(n31976) );
  NANDN U40901 ( .A(n32010), .B(n32011), .Z(n32009) );
  OR U40902 ( .A(n32012), .B(n32013), .Z(n32011) );
  NANDN U40903 ( .A(n32014), .B(n32012), .Z(n32008) );
  IV U40904 ( .A(n32013), .Z(n32014) );
  XNOR U40905 ( .A(n31984), .B(n32015), .Z(n31979) );
  XNOR U40906 ( .A(n31982), .B(n31985), .Z(n32015) );
  NAND U40907 ( .A(n32016), .B(n32017), .Z(n31985) );
  NAND U40908 ( .A(n32018), .B(n32019), .Z(n32017) );
  OR U40909 ( .A(n32020), .B(n32021), .Z(n32018) );
  NANDN U40910 ( .A(n32022), .B(n32020), .Z(n32016) );
  IV U40911 ( .A(n32021), .Z(n32022) );
  NAND U40912 ( .A(n32023), .B(n32024), .Z(n31982) );
  NAND U40913 ( .A(n32025), .B(n32026), .Z(n32024) );
  NANDN U40914 ( .A(n32027), .B(n32028), .Z(n32025) );
  NANDN U40915 ( .A(n32028), .B(n32027), .Z(n32023) );
  AND U40916 ( .A(n32029), .B(n32030), .Z(n31984) );
  NAND U40917 ( .A(n32031), .B(n32032), .Z(n32030) );
  OR U40918 ( .A(n32033), .B(n32034), .Z(n32031) );
  NANDN U40919 ( .A(n32035), .B(n32033), .Z(n32029) );
  XNOR U40920 ( .A(n32010), .B(n32036), .Z(N62556) );
  XOR U40921 ( .A(n32012), .B(n32013), .Z(n32036) );
  XNOR U40922 ( .A(n32026), .B(n32037), .Z(n32013) );
  XOR U40923 ( .A(n32027), .B(n32028), .Z(n32037) );
  XOR U40924 ( .A(n32033), .B(n32038), .Z(n32028) );
  XOR U40925 ( .A(n32032), .B(n32035), .Z(n32038) );
  IV U40926 ( .A(n32034), .Z(n32035) );
  NAND U40927 ( .A(n32039), .B(n32040), .Z(n32034) );
  OR U40928 ( .A(n32041), .B(n32042), .Z(n32040) );
  OR U40929 ( .A(n32043), .B(n32044), .Z(n32039) );
  NAND U40930 ( .A(n32045), .B(n32046), .Z(n32032) );
  OR U40931 ( .A(n32047), .B(n32048), .Z(n32046) );
  OR U40932 ( .A(n32049), .B(n32050), .Z(n32045) );
  NOR U40933 ( .A(n32051), .B(n32052), .Z(n32033) );
  ANDN U40934 ( .B(n32053), .A(n32054), .Z(n32027) );
  XNOR U40935 ( .A(n32020), .B(n32055), .Z(n32026) );
  XNOR U40936 ( .A(n32019), .B(n32021), .Z(n32055) );
  NAND U40937 ( .A(n32056), .B(n32057), .Z(n32021) );
  OR U40938 ( .A(n32058), .B(n32059), .Z(n32057) );
  OR U40939 ( .A(n32060), .B(n32061), .Z(n32056) );
  NAND U40940 ( .A(n32062), .B(n32063), .Z(n32019) );
  OR U40941 ( .A(n32064), .B(n32065), .Z(n32063) );
  OR U40942 ( .A(n32066), .B(n32067), .Z(n32062) );
  ANDN U40943 ( .B(n32068), .A(n32069), .Z(n32020) );
  IV U40944 ( .A(n32070), .Z(n32068) );
  ANDN U40945 ( .B(n32071), .A(n32072), .Z(n32012) );
  XOR U40946 ( .A(n31998), .B(n32073), .Z(n32010) );
  XOR U40947 ( .A(n31999), .B(n32000), .Z(n32073) );
  XOR U40948 ( .A(n32005), .B(n32074), .Z(n32000) );
  XOR U40949 ( .A(n32004), .B(n32007), .Z(n32074) );
  IV U40950 ( .A(n32006), .Z(n32007) );
  NAND U40951 ( .A(n32075), .B(n32076), .Z(n32006) );
  OR U40952 ( .A(n32077), .B(n32078), .Z(n32076) );
  OR U40953 ( .A(n32079), .B(n32080), .Z(n32075) );
  NAND U40954 ( .A(n32081), .B(n32082), .Z(n32004) );
  OR U40955 ( .A(n32083), .B(n32084), .Z(n32082) );
  OR U40956 ( .A(n32085), .B(n32086), .Z(n32081) );
  NOR U40957 ( .A(n32087), .B(n32088), .Z(n32005) );
  ANDN U40958 ( .B(n32089), .A(n32090), .Z(n31999) );
  IV U40959 ( .A(n32091), .Z(n32089) );
  XNOR U40960 ( .A(n31992), .B(n32092), .Z(n31998) );
  XNOR U40961 ( .A(n31991), .B(n31993), .Z(n32092) );
  NAND U40962 ( .A(n32093), .B(n32094), .Z(n31993) );
  OR U40963 ( .A(n32095), .B(n32096), .Z(n32094) );
  OR U40964 ( .A(n32097), .B(n32098), .Z(n32093) );
  NAND U40965 ( .A(n32099), .B(n32100), .Z(n31991) );
  OR U40966 ( .A(n32101), .B(n32102), .Z(n32100) );
  OR U40967 ( .A(n32103), .B(n32104), .Z(n32099) );
  ANDN U40968 ( .B(n32105), .A(n32106), .Z(n31992) );
  IV U40969 ( .A(n32107), .Z(n32105) );
  XNOR U40970 ( .A(n32072), .B(n32071), .Z(N62555) );
  XOR U40971 ( .A(n32091), .B(n32090), .Z(n32071) );
  XNOR U40972 ( .A(n32106), .B(n32107), .Z(n32090) );
  XNOR U40973 ( .A(n32101), .B(n32102), .Z(n32107) );
  XNOR U40974 ( .A(n32103), .B(n32104), .Z(n32102) );
  XNOR U40975 ( .A(y[3637]), .B(x[3637]), .Z(n32104) );
  XNOR U40976 ( .A(y[3638]), .B(x[3638]), .Z(n32103) );
  XNOR U40977 ( .A(y[3636]), .B(x[3636]), .Z(n32101) );
  XNOR U40978 ( .A(n32095), .B(n32096), .Z(n32106) );
  XNOR U40979 ( .A(y[3633]), .B(x[3633]), .Z(n32096) );
  XNOR U40980 ( .A(n32097), .B(n32098), .Z(n32095) );
  XNOR U40981 ( .A(y[3634]), .B(x[3634]), .Z(n32098) );
  XNOR U40982 ( .A(y[3635]), .B(x[3635]), .Z(n32097) );
  XNOR U40983 ( .A(n32088), .B(n32087), .Z(n32091) );
  XNOR U40984 ( .A(n32083), .B(n32084), .Z(n32087) );
  XNOR U40985 ( .A(y[3630]), .B(x[3630]), .Z(n32084) );
  XNOR U40986 ( .A(n32085), .B(n32086), .Z(n32083) );
  XNOR U40987 ( .A(y[3631]), .B(x[3631]), .Z(n32086) );
  XNOR U40988 ( .A(y[3632]), .B(x[3632]), .Z(n32085) );
  XNOR U40989 ( .A(n32077), .B(n32078), .Z(n32088) );
  XNOR U40990 ( .A(y[3627]), .B(x[3627]), .Z(n32078) );
  XNOR U40991 ( .A(n32079), .B(n32080), .Z(n32077) );
  XNOR U40992 ( .A(y[3628]), .B(x[3628]), .Z(n32080) );
  XNOR U40993 ( .A(y[3629]), .B(x[3629]), .Z(n32079) );
  XOR U40994 ( .A(n32053), .B(n32054), .Z(n32072) );
  XNOR U40995 ( .A(n32069), .B(n32070), .Z(n32054) );
  XNOR U40996 ( .A(n32064), .B(n32065), .Z(n32070) );
  XNOR U40997 ( .A(n32066), .B(n32067), .Z(n32065) );
  XNOR U40998 ( .A(y[3625]), .B(x[3625]), .Z(n32067) );
  XNOR U40999 ( .A(y[3626]), .B(x[3626]), .Z(n32066) );
  XNOR U41000 ( .A(y[3624]), .B(x[3624]), .Z(n32064) );
  XNOR U41001 ( .A(n32058), .B(n32059), .Z(n32069) );
  XNOR U41002 ( .A(y[3621]), .B(x[3621]), .Z(n32059) );
  XNOR U41003 ( .A(n32060), .B(n32061), .Z(n32058) );
  XNOR U41004 ( .A(y[3622]), .B(x[3622]), .Z(n32061) );
  XNOR U41005 ( .A(y[3623]), .B(x[3623]), .Z(n32060) );
  XOR U41006 ( .A(n32052), .B(n32051), .Z(n32053) );
  XNOR U41007 ( .A(n32047), .B(n32048), .Z(n32051) );
  XNOR U41008 ( .A(y[3618]), .B(x[3618]), .Z(n32048) );
  XNOR U41009 ( .A(n32049), .B(n32050), .Z(n32047) );
  XNOR U41010 ( .A(y[3619]), .B(x[3619]), .Z(n32050) );
  XNOR U41011 ( .A(y[3620]), .B(x[3620]), .Z(n32049) );
  XNOR U41012 ( .A(n32041), .B(n32042), .Z(n32052) );
  XNOR U41013 ( .A(y[3615]), .B(x[3615]), .Z(n32042) );
  XNOR U41014 ( .A(n32043), .B(n32044), .Z(n32041) );
  XNOR U41015 ( .A(y[3616]), .B(x[3616]), .Z(n32044) );
  XNOR U41016 ( .A(y[3617]), .B(x[3617]), .Z(n32043) );
  NAND U41017 ( .A(n32108), .B(n32109), .Z(N62546) );
  NANDN U41018 ( .A(n32110), .B(n32111), .Z(n32109) );
  OR U41019 ( .A(n32112), .B(n32113), .Z(n32111) );
  NAND U41020 ( .A(n32112), .B(n32113), .Z(n32108) );
  XOR U41021 ( .A(n32112), .B(n32114), .Z(N62545) );
  XNOR U41022 ( .A(n32110), .B(n32113), .Z(n32114) );
  AND U41023 ( .A(n32115), .B(n32116), .Z(n32113) );
  NANDN U41024 ( .A(n32117), .B(n32118), .Z(n32116) );
  NANDN U41025 ( .A(n32119), .B(n32120), .Z(n32118) );
  NANDN U41026 ( .A(n32120), .B(n32119), .Z(n32115) );
  NAND U41027 ( .A(n32121), .B(n32122), .Z(n32110) );
  NANDN U41028 ( .A(n32123), .B(n32124), .Z(n32122) );
  OR U41029 ( .A(n32125), .B(n32126), .Z(n32124) );
  NAND U41030 ( .A(n32126), .B(n32125), .Z(n32121) );
  AND U41031 ( .A(n32127), .B(n32128), .Z(n32112) );
  NANDN U41032 ( .A(n32129), .B(n32130), .Z(n32128) );
  NANDN U41033 ( .A(n32131), .B(n32132), .Z(n32130) );
  NANDN U41034 ( .A(n32132), .B(n32131), .Z(n32127) );
  XOR U41035 ( .A(n32126), .B(n32133), .Z(N62544) );
  XOR U41036 ( .A(n32123), .B(n32125), .Z(n32133) );
  XNOR U41037 ( .A(n32119), .B(n32134), .Z(n32125) );
  XNOR U41038 ( .A(n32117), .B(n32120), .Z(n32134) );
  NAND U41039 ( .A(n32135), .B(n32136), .Z(n32120) );
  NAND U41040 ( .A(n32137), .B(n32138), .Z(n32136) );
  OR U41041 ( .A(n32139), .B(n32140), .Z(n32137) );
  NANDN U41042 ( .A(n32141), .B(n32139), .Z(n32135) );
  IV U41043 ( .A(n32140), .Z(n32141) );
  NAND U41044 ( .A(n32142), .B(n32143), .Z(n32117) );
  NAND U41045 ( .A(n32144), .B(n32145), .Z(n32143) );
  NANDN U41046 ( .A(n32146), .B(n32147), .Z(n32144) );
  NANDN U41047 ( .A(n32147), .B(n32146), .Z(n32142) );
  AND U41048 ( .A(n32148), .B(n32149), .Z(n32119) );
  NAND U41049 ( .A(n32150), .B(n32151), .Z(n32149) );
  OR U41050 ( .A(n32152), .B(n32153), .Z(n32150) );
  NANDN U41051 ( .A(n32154), .B(n32152), .Z(n32148) );
  NAND U41052 ( .A(n32155), .B(n32156), .Z(n32123) );
  NANDN U41053 ( .A(n32157), .B(n32158), .Z(n32156) );
  OR U41054 ( .A(n32159), .B(n32160), .Z(n32158) );
  NANDN U41055 ( .A(n32161), .B(n32159), .Z(n32155) );
  IV U41056 ( .A(n32160), .Z(n32161) );
  XNOR U41057 ( .A(n32131), .B(n32162), .Z(n32126) );
  XNOR U41058 ( .A(n32129), .B(n32132), .Z(n32162) );
  NAND U41059 ( .A(n32163), .B(n32164), .Z(n32132) );
  NAND U41060 ( .A(n32165), .B(n32166), .Z(n32164) );
  OR U41061 ( .A(n32167), .B(n32168), .Z(n32165) );
  NANDN U41062 ( .A(n32169), .B(n32167), .Z(n32163) );
  IV U41063 ( .A(n32168), .Z(n32169) );
  NAND U41064 ( .A(n32170), .B(n32171), .Z(n32129) );
  NAND U41065 ( .A(n32172), .B(n32173), .Z(n32171) );
  NANDN U41066 ( .A(n32174), .B(n32175), .Z(n32172) );
  NANDN U41067 ( .A(n32175), .B(n32174), .Z(n32170) );
  AND U41068 ( .A(n32176), .B(n32177), .Z(n32131) );
  NAND U41069 ( .A(n32178), .B(n32179), .Z(n32177) );
  OR U41070 ( .A(n32180), .B(n32181), .Z(n32178) );
  NANDN U41071 ( .A(n32182), .B(n32180), .Z(n32176) );
  XNOR U41072 ( .A(n32157), .B(n32183), .Z(N62543) );
  XOR U41073 ( .A(n32159), .B(n32160), .Z(n32183) );
  XNOR U41074 ( .A(n32173), .B(n32184), .Z(n32160) );
  XOR U41075 ( .A(n32174), .B(n32175), .Z(n32184) );
  XOR U41076 ( .A(n32180), .B(n32185), .Z(n32175) );
  XOR U41077 ( .A(n32179), .B(n32182), .Z(n32185) );
  IV U41078 ( .A(n32181), .Z(n32182) );
  NAND U41079 ( .A(n32186), .B(n32187), .Z(n32181) );
  OR U41080 ( .A(n32188), .B(n32189), .Z(n32187) );
  OR U41081 ( .A(n32190), .B(n32191), .Z(n32186) );
  NAND U41082 ( .A(n32192), .B(n32193), .Z(n32179) );
  OR U41083 ( .A(n32194), .B(n32195), .Z(n32193) );
  OR U41084 ( .A(n32196), .B(n32197), .Z(n32192) );
  NOR U41085 ( .A(n32198), .B(n32199), .Z(n32180) );
  ANDN U41086 ( .B(n32200), .A(n32201), .Z(n32174) );
  XNOR U41087 ( .A(n32167), .B(n32202), .Z(n32173) );
  XNOR U41088 ( .A(n32166), .B(n32168), .Z(n32202) );
  NAND U41089 ( .A(n32203), .B(n32204), .Z(n32168) );
  OR U41090 ( .A(n32205), .B(n32206), .Z(n32204) );
  OR U41091 ( .A(n32207), .B(n32208), .Z(n32203) );
  NAND U41092 ( .A(n32209), .B(n32210), .Z(n32166) );
  OR U41093 ( .A(n32211), .B(n32212), .Z(n32210) );
  OR U41094 ( .A(n32213), .B(n32214), .Z(n32209) );
  ANDN U41095 ( .B(n32215), .A(n32216), .Z(n32167) );
  IV U41096 ( .A(n32217), .Z(n32215) );
  ANDN U41097 ( .B(n32218), .A(n32219), .Z(n32159) );
  XOR U41098 ( .A(n32145), .B(n32220), .Z(n32157) );
  XOR U41099 ( .A(n32146), .B(n32147), .Z(n32220) );
  XOR U41100 ( .A(n32152), .B(n32221), .Z(n32147) );
  XOR U41101 ( .A(n32151), .B(n32154), .Z(n32221) );
  IV U41102 ( .A(n32153), .Z(n32154) );
  NAND U41103 ( .A(n32222), .B(n32223), .Z(n32153) );
  OR U41104 ( .A(n32224), .B(n32225), .Z(n32223) );
  OR U41105 ( .A(n32226), .B(n32227), .Z(n32222) );
  NAND U41106 ( .A(n32228), .B(n32229), .Z(n32151) );
  OR U41107 ( .A(n32230), .B(n32231), .Z(n32229) );
  OR U41108 ( .A(n32232), .B(n32233), .Z(n32228) );
  NOR U41109 ( .A(n32234), .B(n32235), .Z(n32152) );
  ANDN U41110 ( .B(n32236), .A(n32237), .Z(n32146) );
  IV U41111 ( .A(n32238), .Z(n32236) );
  XNOR U41112 ( .A(n32139), .B(n32239), .Z(n32145) );
  XNOR U41113 ( .A(n32138), .B(n32140), .Z(n32239) );
  NAND U41114 ( .A(n32240), .B(n32241), .Z(n32140) );
  OR U41115 ( .A(n32242), .B(n32243), .Z(n32241) );
  OR U41116 ( .A(n32244), .B(n32245), .Z(n32240) );
  NAND U41117 ( .A(n32246), .B(n32247), .Z(n32138) );
  OR U41118 ( .A(n32248), .B(n32249), .Z(n32247) );
  OR U41119 ( .A(n32250), .B(n32251), .Z(n32246) );
  ANDN U41120 ( .B(n32252), .A(n32253), .Z(n32139) );
  IV U41121 ( .A(n32254), .Z(n32252) );
  XNOR U41122 ( .A(n32219), .B(n32218), .Z(N62542) );
  XOR U41123 ( .A(n32238), .B(n32237), .Z(n32218) );
  XNOR U41124 ( .A(n32253), .B(n32254), .Z(n32237) );
  XNOR U41125 ( .A(n32248), .B(n32249), .Z(n32254) );
  XNOR U41126 ( .A(n32250), .B(n32251), .Z(n32249) );
  XNOR U41127 ( .A(y[3613]), .B(x[3613]), .Z(n32251) );
  XNOR U41128 ( .A(y[3614]), .B(x[3614]), .Z(n32250) );
  XNOR U41129 ( .A(y[3612]), .B(x[3612]), .Z(n32248) );
  XNOR U41130 ( .A(n32242), .B(n32243), .Z(n32253) );
  XNOR U41131 ( .A(y[3609]), .B(x[3609]), .Z(n32243) );
  XNOR U41132 ( .A(n32244), .B(n32245), .Z(n32242) );
  XNOR U41133 ( .A(y[3610]), .B(x[3610]), .Z(n32245) );
  XNOR U41134 ( .A(y[3611]), .B(x[3611]), .Z(n32244) );
  XNOR U41135 ( .A(n32235), .B(n32234), .Z(n32238) );
  XNOR U41136 ( .A(n32230), .B(n32231), .Z(n32234) );
  XNOR U41137 ( .A(y[3606]), .B(x[3606]), .Z(n32231) );
  XNOR U41138 ( .A(n32232), .B(n32233), .Z(n32230) );
  XNOR U41139 ( .A(y[3607]), .B(x[3607]), .Z(n32233) );
  XNOR U41140 ( .A(y[3608]), .B(x[3608]), .Z(n32232) );
  XNOR U41141 ( .A(n32224), .B(n32225), .Z(n32235) );
  XNOR U41142 ( .A(y[3603]), .B(x[3603]), .Z(n32225) );
  XNOR U41143 ( .A(n32226), .B(n32227), .Z(n32224) );
  XNOR U41144 ( .A(y[3604]), .B(x[3604]), .Z(n32227) );
  XNOR U41145 ( .A(y[3605]), .B(x[3605]), .Z(n32226) );
  XOR U41146 ( .A(n32200), .B(n32201), .Z(n32219) );
  XNOR U41147 ( .A(n32216), .B(n32217), .Z(n32201) );
  XNOR U41148 ( .A(n32211), .B(n32212), .Z(n32217) );
  XNOR U41149 ( .A(n32213), .B(n32214), .Z(n32212) );
  XNOR U41150 ( .A(y[3601]), .B(x[3601]), .Z(n32214) );
  XNOR U41151 ( .A(y[3602]), .B(x[3602]), .Z(n32213) );
  XNOR U41152 ( .A(y[3600]), .B(x[3600]), .Z(n32211) );
  XNOR U41153 ( .A(n32205), .B(n32206), .Z(n32216) );
  XNOR U41154 ( .A(y[3597]), .B(x[3597]), .Z(n32206) );
  XNOR U41155 ( .A(n32207), .B(n32208), .Z(n32205) );
  XNOR U41156 ( .A(y[3598]), .B(x[3598]), .Z(n32208) );
  XNOR U41157 ( .A(y[3599]), .B(x[3599]), .Z(n32207) );
  XOR U41158 ( .A(n32199), .B(n32198), .Z(n32200) );
  XNOR U41159 ( .A(n32194), .B(n32195), .Z(n32198) );
  XNOR U41160 ( .A(y[3594]), .B(x[3594]), .Z(n32195) );
  XNOR U41161 ( .A(n32196), .B(n32197), .Z(n32194) );
  XNOR U41162 ( .A(y[3595]), .B(x[3595]), .Z(n32197) );
  XNOR U41163 ( .A(y[3596]), .B(x[3596]), .Z(n32196) );
  XNOR U41164 ( .A(n32188), .B(n32189), .Z(n32199) );
  XNOR U41165 ( .A(y[3591]), .B(x[3591]), .Z(n32189) );
  XNOR U41166 ( .A(n32190), .B(n32191), .Z(n32188) );
  XNOR U41167 ( .A(y[3592]), .B(x[3592]), .Z(n32191) );
  XNOR U41168 ( .A(y[3593]), .B(x[3593]), .Z(n32190) );
  NAND U41169 ( .A(n32255), .B(n32256), .Z(N62533) );
  NANDN U41170 ( .A(n32257), .B(n32258), .Z(n32256) );
  OR U41171 ( .A(n32259), .B(n32260), .Z(n32258) );
  NAND U41172 ( .A(n32259), .B(n32260), .Z(n32255) );
  XOR U41173 ( .A(n32259), .B(n32261), .Z(N62532) );
  XNOR U41174 ( .A(n32257), .B(n32260), .Z(n32261) );
  AND U41175 ( .A(n32262), .B(n32263), .Z(n32260) );
  NANDN U41176 ( .A(n32264), .B(n32265), .Z(n32263) );
  NANDN U41177 ( .A(n32266), .B(n32267), .Z(n32265) );
  NANDN U41178 ( .A(n32267), .B(n32266), .Z(n32262) );
  NAND U41179 ( .A(n32268), .B(n32269), .Z(n32257) );
  NANDN U41180 ( .A(n32270), .B(n32271), .Z(n32269) );
  OR U41181 ( .A(n32272), .B(n32273), .Z(n32271) );
  NAND U41182 ( .A(n32273), .B(n32272), .Z(n32268) );
  AND U41183 ( .A(n32274), .B(n32275), .Z(n32259) );
  NANDN U41184 ( .A(n32276), .B(n32277), .Z(n32275) );
  NANDN U41185 ( .A(n32278), .B(n32279), .Z(n32277) );
  NANDN U41186 ( .A(n32279), .B(n32278), .Z(n32274) );
  XOR U41187 ( .A(n32273), .B(n32280), .Z(N62531) );
  XOR U41188 ( .A(n32270), .B(n32272), .Z(n32280) );
  XNOR U41189 ( .A(n32266), .B(n32281), .Z(n32272) );
  XNOR U41190 ( .A(n32264), .B(n32267), .Z(n32281) );
  NAND U41191 ( .A(n32282), .B(n32283), .Z(n32267) );
  NAND U41192 ( .A(n32284), .B(n32285), .Z(n32283) );
  OR U41193 ( .A(n32286), .B(n32287), .Z(n32284) );
  NANDN U41194 ( .A(n32288), .B(n32286), .Z(n32282) );
  IV U41195 ( .A(n32287), .Z(n32288) );
  NAND U41196 ( .A(n32289), .B(n32290), .Z(n32264) );
  NAND U41197 ( .A(n32291), .B(n32292), .Z(n32290) );
  NANDN U41198 ( .A(n32293), .B(n32294), .Z(n32291) );
  NANDN U41199 ( .A(n32294), .B(n32293), .Z(n32289) );
  AND U41200 ( .A(n32295), .B(n32296), .Z(n32266) );
  NAND U41201 ( .A(n32297), .B(n32298), .Z(n32296) );
  OR U41202 ( .A(n32299), .B(n32300), .Z(n32297) );
  NANDN U41203 ( .A(n32301), .B(n32299), .Z(n32295) );
  NAND U41204 ( .A(n32302), .B(n32303), .Z(n32270) );
  NANDN U41205 ( .A(n32304), .B(n32305), .Z(n32303) );
  OR U41206 ( .A(n32306), .B(n32307), .Z(n32305) );
  NANDN U41207 ( .A(n32308), .B(n32306), .Z(n32302) );
  IV U41208 ( .A(n32307), .Z(n32308) );
  XNOR U41209 ( .A(n32278), .B(n32309), .Z(n32273) );
  XNOR U41210 ( .A(n32276), .B(n32279), .Z(n32309) );
  NAND U41211 ( .A(n32310), .B(n32311), .Z(n32279) );
  NAND U41212 ( .A(n32312), .B(n32313), .Z(n32311) );
  OR U41213 ( .A(n32314), .B(n32315), .Z(n32312) );
  NANDN U41214 ( .A(n32316), .B(n32314), .Z(n32310) );
  IV U41215 ( .A(n32315), .Z(n32316) );
  NAND U41216 ( .A(n32317), .B(n32318), .Z(n32276) );
  NAND U41217 ( .A(n32319), .B(n32320), .Z(n32318) );
  NANDN U41218 ( .A(n32321), .B(n32322), .Z(n32319) );
  NANDN U41219 ( .A(n32322), .B(n32321), .Z(n32317) );
  AND U41220 ( .A(n32323), .B(n32324), .Z(n32278) );
  NAND U41221 ( .A(n32325), .B(n32326), .Z(n32324) );
  OR U41222 ( .A(n32327), .B(n32328), .Z(n32325) );
  NANDN U41223 ( .A(n32329), .B(n32327), .Z(n32323) );
  XNOR U41224 ( .A(n32304), .B(n32330), .Z(N62530) );
  XOR U41225 ( .A(n32306), .B(n32307), .Z(n32330) );
  XNOR U41226 ( .A(n32320), .B(n32331), .Z(n32307) );
  XOR U41227 ( .A(n32321), .B(n32322), .Z(n32331) );
  XOR U41228 ( .A(n32327), .B(n32332), .Z(n32322) );
  XOR U41229 ( .A(n32326), .B(n32329), .Z(n32332) );
  IV U41230 ( .A(n32328), .Z(n32329) );
  NAND U41231 ( .A(n32333), .B(n32334), .Z(n32328) );
  OR U41232 ( .A(n32335), .B(n32336), .Z(n32334) );
  OR U41233 ( .A(n32337), .B(n32338), .Z(n32333) );
  NAND U41234 ( .A(n32339), .B(n32340), .Z(n32326) );
  OR U41235 ( .A(n32341), .B(n32342), .Z(n32340) );
  OR U41236 ( .A(n32343), .B(n32344), .Z(n32339) );
  NOR U41237 ( .A(n32345), .B(n32346), .Z(n32327) );
  ANDN U41238 ( .B(n32347), .A(n32348), .Z(n32321) );
  XNOR U41239 ( .A(n32314), .B(n32349), .Z(n32320) );
  XNOR U41240 ( .A(n32313), .B(n32315), .Z(n32349) );
  NAND U41241 ( .A(n32350), .B(n32351), .Z(n32315) );
  OR U41242 ( .A(n32352), .B(n32353), .Z(n32351) );
  OR U41243 ( .A(n32354), .B(n32355), .Z(n32350) );
  NAND U41244 ( .A(n32356), .B(n32357), .Z(n32313) );
  OR U41245 ( .A(n32358), .B(n32359), .Z(n32357) );
  OR U41246 ( .A(n32360), .B(n32361), .Z(n32356) );
  ANDN U41247 ( .B(n32362), .A(n32363), .Z(n32314) );
  IV U41248 ( .A(n32364), .Z(n32362) );
  ANDN U41249 ( .B(n32365), .A(n32366), .Z(n32306) );
  XOR U41250 ( .A(n32292), .B(n32367), .Z(n32304) );
  XOR U41251 ( .A(n32293), .B(n32294), .Z(n32367) );
  XOR U41252 ( .A(n32299), .B(n32368), .Z(n32294) );
  XOR U41253 ( .A(n32298), .B(n32301), .Z(n32368) );
  IV U41254 ( .A(n32300), .Z(n32301) );
  NAND U41255 ( .A(n32369), .B(n32370), .Z(n32300) );
  OR U41256 ( .A(n32371), .B(n32372), .Z(n32370) );
  OR U41257 ( .A(n32373), .B(n32374), .Z(n32369) );
  NAND U41258 ( .A(n32375), .B(n32376), .Z(n32298) );
  OR U41259 ( .A(n32377), .B(n32378), .Z(n32376) );
  OR U41260 ( .A(n32379), .B(n32380), .Z(n32375) );
  NOR U41261 ( .A(n32381), .B(n32382), .Z(n32299) );
  ANDN U41262 ( .B(n32383), .A(n32384), .Z(n32293) );
  IV U41263 ( .A(n32385), .Z(n32383) );
  XNOR U41264 ( .A(n32286), .B(n32386), .Z(n32292) );
  XNOR U41265 ( .A(n32285), .B(n32287), .Z(n32386) );
  NAND U41266 ( .A(n32387), .B(n32388), .Z(n32287) );
  OR U41267 ( .A(n32389), .B(n32390), .Z(n32388) );
  OR U41268 ( .A(n32391), .B(n32392), .Z(n32387) );
  NAND U41269 ( .A(n32393), .B(n32394), .Z(n32285) );
  OR U41270 ( .A(n32395), .B(n32396), .Z(n32394) );
  OR U41271 ( .A(n32397), .B(n32398), .Z(n32393) );
  ANDN U41272 ( .B(n32399), .A(n32400), .Z(n32286) );
  IV U41273 ( .A(n32401), .Z(n32399) );
  XNOR U41274 ( .A(n32366), .B(n32365), .Z(N62529) );
  XOR U41275 ( .A(n32385), .B(n32384), .Z(n32365) );
  XNOR U41276 ( .A(n32400), .B(n32401), .Z(n32384) );
  XNOR U41277 ( .A(n32395), .B(n32396), .Z(n32401) );
  XNOR U41278 ( .A(n32397), .B(n32398), .Z(n32396) );
  XNOR U41279 ( .A(y[3589]), .B(x[3589]), .Z(n32398) );
  XNOR U41280 ( .A(y[3590]), .B(x[3590]), .Z(n32397) );
  XNOR U41281 ( .A(y[3588]), .B(x[3588]), .Z(n32395) );
  XNOR U41282 ( .A(n32389), .B(n32390), .Z(n32400) );
  XNOR U41283 ( .A(y[3585]), .B(x[3585]), .Z(n32390) );
  XNOR U41284 ( .A(n32391), .B(n32392), .Z(n32389) );
  XNOR U41285 ( .A(y[3586]), .B(x[3586]), .Z(n32392) );
  XNOR U41286 ( .A(y[3587]), .B(x[3587]), .Z(n32391) );
  XNOR U41287 ( .A(n32382), .B(n32381), .Z(n32385) );
  XNOR U41288 ( .A(n32377), .B(n32378), .Z(n32381) );
  XNOR U41289 ( .A(y[3582]), .B(x[3582]), .Z(n32378) );
  XNOR U41290 ( .A(n32379), .B(n32380), .Z(n32377) );
  XNOR U41291 ( .A(y[3583]), .B(x[3583]), .Z(n32380) );
  XNOR U41292 ( .A(y[3584]), .B(x[3584]), .Z(n32379) );
  XNOR U41293 ( .A(n32371), .B(n32372), .Z(n32382) );
  XNOR U41294 ( .A(y[3579]), .B(x[3579]), .Z(n32372) );
  XNOR U41295 ( .A(n32373), .B(n32374), .Z(n32371) );
  XNOR U41296 ( .A(y[3580]), .B(x[3580]), .Z(n32374) );
  XNOR U41297 ( .A(y[3581]), .B(x[3581]), .Z(n32373) );
  XOR U41298 ( .A(n32347), .B(n32348), .Z(n32366) );
  XNOR U41299 ( .A(n32363), .B(n32364), .Z(n32348) );
  XNOR U41300 ( .A(n32358), .B(n32359), .Z(n32364) );
  XNOR U41301 ( .A(n32360), .B(n32361), .Z(n32359) );
  XNOR U41302 ( .A(y[3577]), .B(x[3577]), .Z(n32361) );
  XNOR U41303 ( .A(y[3578]), .B(x[3578]), .Z(n32360) );
  XNOR U41304 ( .A(y[3576]), .B(x[3576]), .Z(n32358) );
  XNOR U41305 ( .A(n32352), .B(n32353), .Z(n32363) );
  XNOR U41306 ( .A(y[3573]), .B(x[3573]), .Z(n32353) );
  XNOR U41307 ( .A(n32354), .B(n32355), .Z(n32352) );
  XNOR U41308 ( .A(y[3574]), .B(x[3574]), .Z(n32355) );
  XNOR U41309 ( .A(y[3575]), .B(x[3575]), .Z(n32354) );
  XOR U41310 ( .A(n32346), .B(n32345), .Z(n32347) );
  XNOR U41311 ( .A(n32341), .B(n32342), .Z(n32345) );
  XNOR U41312 ( .A(y[3570]), .B(x[3570]), .Z(n32342) );
  XNOR U41313 ( .A(n32343), .B(n32344), .Z(n32341) );
  XNOR U41314 ( .A(y[3571]), .B(x[3571]), .Z(n32344) );
  XNOR U41315 ( .A(y[3572]), .B(x[3572]), .Z(n32343) );
  XNOR U41316 ( .A(n32335), .B(n32336), .Z(n32346) );
  XNOR U41317 ( .A(y[3567]), .B(x[3567]), .Z(n32336) );
  XNOR U41318 ( .A(n32337), .B(n32338), .Z(n32335) );
  XNOR U41319 ( .A(y[3568]), .B(x[3568]), .Z(n32338) );
  XNOR U41320 ( .A(y[3569]), .B(x[3569]), .Z(n32337) );
  NAND U41321 ( .A(n32402), .B(n32403), .Z(N62520) );
  NANDN U41322 ( .A(n32404), .B(n32405), .Z(n32403) );
  OR U41323 ( .A(n32406), .B(n32407), .Z(n32405) );
  NAND U41324 ( .A(n32406), .B(n32407), .Z(n32402) );
  XOR U41325 ( .A(n32406), .B(n32408), .Z(N62519) );
  XNOR U41326 ( .A(n32404), .B(n32407), .Z(n32408) );
  AND U41327 ( .A(n32409), .B(n32410), .Z(n32407) );
  NANDN U41328 ( .A(n32411), .B(n32412), .Z(n32410) );
  NANDN U41329 ( .A(n32413), .B(n32414), .Z(n32412) );
  NANDN U41330 ( .A(n32414), .B(n32413), .Z(n32409) );
  NAND U41331 ( .A(n32415), .B(n32416), .Z(n32404) );
  NANDN U41332 ( .A(n32417), .B(n32418), .Z(n32416) );
  OR U41333 ( .A(n32419), .B(n32420), .Z(n32418) );
  NAND U41334 ( .A(n32420), .B(n32419), .Z(n32415) );
  AND U41335 ( .A(n32421), .B(n32422), .Z(n32406) );
  NANDN U41336 ( .A(n32423), .B(n32424), .Z(n32422) );
  NANDN U41337 ( .A(n32425), .B(n32426), .Z(n32424) );
  NANDN U41338 ( .A(n32426), .B(n32425), .Z(n32421) );
  XOR U41339 ( .A(n32420), .B(n32427), .Z(N62518) );
  XOR U41340 ( .A(n32417), .B(n32419), .Z(n32427) );
  XNOR U41341 ( .A(n32413), .B(n32428), .Z(n32419) );
  XNOR U41342 ( .A(n32411), .B(n32414), .Z(n32428) );
  NAND U41343 ( .A(n32429), .B(n32430), .Z(n32414) );
  NAND U41344 ( .A(n32431), .B(n32432), .Z(n32430) );
  OR U41345 ( .A(n32433), .B(n32434), .Z(n32431) );
  NANDN U41346 ( .A(n32435), .B(n32433), .Z(n32429) );
  IV U41347 ( .A(n32434), .Z(n32435) );
  NAND U41348 ( .A(n32436), .B(n32437), .Z(n32411) );
  NAND U41349 ( .A(n32438), .B(n32439), .Z(n32437) );
  NANDN U41350 ( .A(n32440), .B(n32441), .Z(n32438) );
  NANDN U41351 ( .A(n32441), .B(n32440), .Z(n32436) );
  AND U41352 ( .A(n32442), .B(n32443), .Z(n32413) );
  NAND U41353 ( .A(n32444), .B(n32445), .Z(n32443) );
  OR U41354 ( .A(n32446), .B(n32447), .Z(n32444) );
  NANDN U41355 ( .A(n32448), .B(n32446), .Z(n32442) );
  NAND U41356 ( .A(n32449), .B(n32450), .Z(n32417) );
  NANDN U41357 ( .A(n32451), .B(n32452), .Z(n32450) );
  OR U41358 ( .A(n32453), .B(n32454), .Z(n32452) );
  NANDN U41359 ( .A(n32455), .B(n32453), .Z(n32449) );
  IV U41360 ( .A(n32454), .Z(n32455) );
  XNOR U41361 ( .A(n32425), .B(n32456), .Z(n32420) );
  XNOR U41362 ( .A(n32423), .B(n32426), .Z(n32456) );
  NAND U41363 ( .A(n32457), .B(n32458), .Z(n32426) );
  NAND U41364 ( .A(n32459), .B(n32460), .Z(n32458) );
  OR U41365 ( .A(n32461), .B(n32462), .Z(n32459) );
  NANDN U41366 ( .A(n32463), .B(n32461), .Z(n32457) );
  IV U41367 ( .A(n32462), .Z(n32463) );
  NAND U41368 ( .A(n32464), .B(n32465), .Z(n32423) );
  NAND U41369 ( .A(n32466), .B(n32467), .Z(n32465) );
  NANDN U41370 ( .A(n32468), .B(n32469), .Z(n32466) );
  NANDN U41371 ( .A(n32469), .B(n32468), .Z(n32464) );
  AND U41372 ( .A(n32470), .B(n32471), .Z(n32425) );
  NAND U41373 ( .A(n32472), .B(n32473), .Z(n32471) );
  OR U41374 ( .A(n32474), .B(n32475), .Z(n32472) );
  NANDN U41375 ( .A(n32476), .B(n32474), .Z(n32470) );
  XNOR U41376 ( .A(n32451), .B(n32477), .Z(N62517) );
  XOR U41377 ( .A(n32453), .B(n32454), .Z(n32477) );
  XNOR U41378 ( .A(n32467), .B(n32478), .Z(n32454) );
  XOR U41379 ( .A(n32468), .B(n32469), .Z(n32478) );
  XOR U41380 ( .A(n32474), .B(n32479), .Z(n32469) );
  XOR U41381 ( .A(n32473), .B(n32476), .Z(n32479) );
  IV U41382 ( .A(n32475), .Z(n32476) );
  NAND U41383 ( .A(n32480), .B(n32481), .Z(n32475) );
  OR U41384 ( .A(n32482), .B(n32483), .Z(n32481) );
  OR U41385 ( .A(n32484), .B(n32485), .Z(n32480) );
  NAND U41386 ( .A(n32486), .B(n32487), .Z(n32473) );
  OR U41387 ( .A(n32488), .B(n32489), .Z(n32487) );
  OR U41388 ( .A(n32490), .B(n32491), .Z(n32486) );
  NOR U41389 ( .A(n32492), .B(n32493), .Z(n32474) );
  ANDN U41390 ( .B(n32494), .A(n32495), .Z(n32468) );
  XNOR U41391 ( .A(n32461), .B(n32496), .Z(n32467) );
  XNOR U41392 ( .A(n32460), .B(n32462), .Z(n32496) );
  NAND U41393 ( .A(n32497), .B(n32498), .Z(n32462) );
  OR U41394 ( .A(n32499), .B(n32500), .Z(n32498) );
  OR U41395 ( .A(n32501), .B(n32502), .Z(n32497) );
  NAND U41396 ( .A(n32503), .B(n32504), .Z(n32460) );
  OR U41397 ( .A(n32505), .B(n32506), .Z(n32504) );
  OR U41398 ( .A(n32507), .B(n32508), .Z(n32503) );
  ANDN U41399 ( .B(n32509), .A(n32510), .Z(n32461) );
  IV U41400 ( .A(n32511), .Z(n32509) );
  ANDN U41401 ( .B(n32512), .A(n32513), .Z(n32453) );
  XOR U41402 ( .A(n32439), .B(n32514), .Z(n32451) );
  XOR U41403 ( .A(n32440), .B(n32441), .Z(n32514) );
  XOR U41404 ( .A(n32446), .B(n32515), .Z(n32441) );
  XOR U41405 ( .A(n32445), .B(n32448), .Z(n32515) );
  IV U41406 ( .A(n32447), .Z(n32448) );
  NAND U41407 ( .A(n32516), .B(n32517), .Z(n32447) );
  OR U41408 ( .A(n32518), .B(n32519), .Z(n32517) );
  OR U41409 ( .A(n32520), .B(n32521), .Z(n32516) );
  NAND U41410 ( .A(n32522), .B(n32523), .Z(n32445) );
  OR U41411 ( .A(n32524), .B(n32525), .Z(n32523) );
  OR U41412 ( .A(n32526), .B(n32527), .Z(n32522) );
  NOR U41413 ( .A(n32528), .B(n32529), .Z(n32446) );
  ANDN U41414 ( .B(n32530), .A(n32531), .Z(n32440) );
  IV U41415 ( .A(n32532), .Z(n32530) );
  XNOR U41416 ( .A(n32433), .B(n32533), .Z(n32439) );
  XNOR U41417 ( .A(n32432), .B(n32434), .Z(n32533) );
  NAND U41418 ( .A(n32534), .B(n32535), .Z(n32434) );
  OR U41419 ( .A(n32536), .B(n32537), .Z(n32535) );
  OR U41420 ( .A(n32538), .B(n32539), .Z(n32534) );
  NAND U41421 ( .A(n32540), .B(n32541), .Z(n32432) );
  OR U41422 ( .A(n32542), .B(n32543), .Z(n32541) );
  OR U41423 ( .A(n32544), .B(n32545), .Z(n32540) );
  ANDN U41424 ( .B(n32546), .A(n32547), .Z(n32433) );
  IV U41425 ( .A(n32548), .Z(n32546) );
  XNOR U41426 ( .A(n32513), .B(n32512), .Z(N62516) );
  XOR U41427 ( .A(n32532), .B(n32531), .Z(n32512) );
  XNOR U41428 ( .A(n32547), .B(n32548), .Z(n32531) );
  XNOR U41429 ( .A(n32542), .B(n32543), .Z(n32548) );
  XNOR U41430 ( .A(n32544), .B(n32545), .Z(n32543) );
  XNOR U41431 ( .A(y[3565]), .B(x[3565]), .Z(n32545) );
  XNOR U41432 ( .A(y[3566]), .B(x[3566]), .Z(n32544) );
  XNOR U41433 ( .A(y[3564]), .B(x[3564]), .Z(n32542) );
  XNOR U41434 ( .A(n32536), .B(n32537), .Z(n32547) );
  XNOR U41435 ( .A(y[3561]), .B(x[3561]), .Z(n32537) );
  XNOR U41436 ( .A(n32538), .B(n32539), .Z(n32536) );
  XNOR U41437 ( .A(y[3562]), .B(x[3562]), .Z(n32539) );
  XNOR U41438 ( .A(y[3563]), .B(x[3563]), .Z(n32538) );
  XNOR U41439 ( .A(n32529), .B(n32528), .Z(n32532) );
  XNOR U41440 ( .A(n32524), .B(n32525), .Z(n32528) );
  XNOR U41441 ( .A(y[3558]), .B(x[3558]), .Z(n32525) );
  XNOR U41442 ( .A(n32526), .B(n32527), .Z(n32524) );
  XNOR U41443 ( .A(y[3559]), .B(x[3559]), .Z(n32527) );
  XNOR U41444 ( .A(y[3560]), .B(x[3560]), .Z(n32526) );
  XNOR U41445 ( .A(n32518), .B(n32519), .Z(n32529) );
  XNOR U41446 ( .A(y[3555]), .B(x[3555]), .Z(n32519) );
  XNOR U41447 ( .A(n32520), .B(n32521), .Z(n32518) );
  XNOR U41448 ( .A(y[3556]), .B(x[3556]), .Z(n32521) );
  XNOR U41449 ( .A(y[3557]), .B(x[3557]), .Z(n32520) );
  XOR U41450 ( .A(n32494), .B(n32495), .Z(n32513) );
  XNOR U41451 ( .A(n32510), .B(n32511), .Z(n32495) );
  XNOR U41452 ( .A(n32505), .B(n32506), .Z(n32511) );
  XNOR U41453 ( .A(n32507), .B(n32508), .Z(n32506) );
  XNOR U41454 ( .A(y[3553]), .B(x[3553]), .Z(n32508) );
  XNOR U41455 ( .A(y[3554]), .B(x[3554]), .Z(n32507) );
  XNOR U41456 ( .A(y[3552]), .B(x[3552]), .Z(n32505) );
  XNOR U41457 ( .A(n32499), .B(n32500), .Z(n32510) );
  XNOR U41458 ( .A(y[3549]), .B(x[3549]), .Z(n32500) );
  XNOR U41459 ( .A(n32501), .B(n32502), .Z(n32499) );
  XNOR U41460 ( .A(y[3550]), .B(x[3550]), .Z(n32502) );
  XNOR U41461 ( .A(y[3551]), .B(x[3551]), .Z(n32501) );
  XOR U41462 ( .A(n32493), .B(n32492), .Z(n32494) );
  XNOR U41463 ( .A(n32488), .B(n32489), .Z(n32492) );
  XNOR U41464 ( .A(y[3546]), .B(x[3546]), .Z(n32489) );
  XNOR U41465 ( .A(n32490), .B(n32491), .Z(n32488) );
  XNOR U41466 ( .A(y[3547]), .B(x[3547]), .Z(n32491) );
  XNOR U41467 ( .A(y[3548]), .B(x[3548]), .Z(n32490) );
  XNOR U41468 ( .A(n32482), .B(n32483), .Z(n32493) );
  XNOR U41469 ( .A(y[3543]), .B(x[3543]), .Z(n32483) );
  XNOR U41470 ( .A(n32484), .B(n32485), .Z(n32482) );
  XNOR U41471 ( .A(y[3544]), .B(x[3544]), .Z(n32485) );
  XNOR U41472 ( .A(y[3545]), .B(x[3545]), .Z(n32484) );
  NAND U41473 ( .A(n32549), .B(n32550), .Z(N62507) );
  NANDN U41474 ( .A(n32551), .B(n32552), .Z(n32550) );
  OR U41475 ( .A(n32553), .B(n32554), .Z(n32552) );
  NAND U41476 ( .A(n32553), .B(n32554), .Z(n32549) );
  XOR U41477 ( .A(n32553), .B(n32555), .Z(N62506) );
  XNOR U41478 ( .A(n32551), .B(n32554), .Z(n32555) );
  AND U41479 ( .A(n32556), .B(n32557), .Z(n32554) );
  NANDN U41480 ( .A(n32558), .B(n32559), .Z(n32557) );
  NANDN U41481 ( .A(n32560), .B(n32561), .Z(n32559) );
  NANDN U41482 ( .A(n32561), .B(n32560), .Z(n32556) );
  NAND U41483 ( .A(n32562), .B(n32563), .Z(n32551) );
  NANDN U41484 ( .A(n32564), .B(n32565), .Z(n32563) );
  OR U41485 ( .A(n32566), .B(n32567), .Z(n32565) );
  NAND U41486 ( .A(n32567), .B(n32566), .Z(n32562) );
  AND U41487 ( .A(n32568), .B(n32569), .Z(n32553) );
  NANDN U41488 ( .A(n32570), .B(n32571), .Z(n32569) );
  NANDN U41489 ( .A(n32572), .B(n32573), .Z(n32571) );
  NANDN U41490 ( .A(n32573), .B(n32572), .Z(n32568) );
  XOR U41491 ( .A(n32567), .B(n32574), .Z(N62505) );
  XOR U41492 ( .A(n32564), .B(n32566), .Z(n32574) );
  XNOR U41493 ( .A(n32560), .B(n32575), .Z(n32566) );
  XNOR U41494 ( .A(n32558), .B(n32561), .Z(n32575) );
  NAND U41495 ( .A(n32576), .B(n32577), .Z(n32561) );
  NAND U41496 ( .A(n32578), .B(n32579), .Z(n32577) );
  OR U41497 ( .A(n32580), .B(n32581), .Z(n32578) );
  NANDN U41498 ( .A(n32582), .B(n32580), .Z(n32576) );
  IV U41499 ( .A(n32581), .Z(n32582) );
  NAND U41500 ( .A(n32583), .B(n32584), .Z(n32558) );
  NAND U41501 ( .A(n32585), .B(n32586), .Z(n32584) );
  NANDN U41502 ( .A(n32587), .B(n32588), .Z(n32585) );
  NANDN U41503 ( .A(n32588), .B(n32587), .Z(n32583) );
  AND U41504 ( .A(n32589), .B(n32590), .Z(n32560) );
  NAND U41505 ( .A(n32591), .B(n32592), .Z(n32590) );
  OR U41506 ( .A(n32593), .B(n32594), .Z(n32591) );
  NANDN U41507 ( .A(n32595), .B(n32593), .Z(n32589) );
  NAND U41508 ( .A(n32596), .B(n32597), .Z(n32564) );
  NANDN U41509 ( .A(n32598), .B(n32599), .Z(n32597) );
  OR U41510 ( .A(n32600), .B(n32601), .Z(n32599) );
  NANDN U41511 ( .A(n32602), .B(n32600), .Z(n32596) );
  IV U41512 ( .A(n32601), .Z(n32602) );
  XNOR U41513 ( .A(n32572), .B(n32603), .Z(n32567) );
  XNOR U41514 ( .A(n32570), .B(n32573), .Z(n32603) );
  NAND U41515 ( .A(n32604), .B(n32605), .Z(n32573) );
  NAND U41516 ( .A(n32606), .B(n32607), .Z(n32605) );
  OR U41517 ( .A(n32608), .B(n32609), .Z(n32606) );
  NANDN U41518 ( .A(n32610), .B(n32608), .Z(n32604) );
  IV U41519 ( .A(n32609), .Z(n32610) );
  NAND U41520 ( .A(n32611), .B(n32612), .Z(n32570) );
  NAND U41521 ( .A(n32613), .B(n32614), .Z(n32612) );
  NANDN U41522 ( .A(n32615), .B(n32616), .Z(n32613) );
  NANDN U41523 ( .A(n32616), .B(n32615), .Z(n32611) );
  AND U41524 ( .A(n32617), .B(n32618), .Z(n32572) );
  NAND U41525 ( .A(n32619), .B(n32620), .Z(n32618) );
  OR U41526 ( .A(n32621), .B(n32622), .Z(n32619) );
  NANDN U41527 ( .A(n32623), .B(n32621), .Z(n32617) );
  XNOR U41528 ( .A(n32598), .B(n32624), .Z(N62504) );
  XOR U41529 ( .A(n32600), .B(n32601), .Z(n32624) );
  XNOR U41530 ( .A(n32614), .B(n32625), .Z(n32601) );
  XOR U41531 ( .A(n32615), .B(n32616), .Z(n32625) );
  XOR U41532 ( .A(n32621), .B(n32626), .Z(n32616) );
  XOR U41533 ( .A(n32620), .B(n32623), .Z(n32626) );
  IV U41534 ( .A(n32622), .Z(n32623) );
  NAND U41535 ( .A(n32627), .B(n32628), .Z(n32622) );
  OR U41536 ( .A(n32629), .B(n32630), .Z(n32628) );
  OR U41537 ( .A(n32631), .B(n32632), .Z(n32627) );
  NAND U41538 ( .A(n32633), .B(n32634), .Z(n32620) );
  OR U41539 ( .A(n32635), .B(n32636), .Z(n32634) );
  OR U41540 ( .A(n32637), .B(n32638), .Z(n32633) );
  NOR U41541 ( .A(n32639), .B(n32640), .Z(n32621) );
  ANDN U41542 ( .B(n32641), .A(n32642), .Z(n32615) );
  XNOR U41543 ( .A(n32608), .B(n32643), .Z(n32614) );
  XNOR U41544 ( .A(n32607), .B(n32609), .Z(n32643) );
  NAND U41545 ( .A(n32644), .B(n32645), .Z(n32609) );
  OR U41546 ( .A(n32646), .B(n32647), .Z(n32645) );
  OR U41547 ( .A(n32648), .B(n32649), .Z(n32644) );
  NAND U41548 ( .A(n32650), .B(n32651), .Z(n32607) );
  OR U41549 ( .A(n32652), .B(n32653), .Z(n32651) );
  OR U41550 ( .A(n32654), .B(n32655), .Z(n32650) );
  ANDN U41551 ( .B(n32656), .A(n32657), .Z(n32608) );
  IV U41552 ( .A(n32658), .Z(n32656) );
  ANDN U41553 ( .B(n32659), .A(n32660), .Z(n32600) );
  XOR U41554 ( .A(n32586), .B(n32661), .Z(n32598) );
  XOR U41555 ( .A(n32587), .B(n32588), .Z(n32661) );
  XOR U41556 ( .A(n32593), .B(n32662), .Z(n32588) );
  XOR U41557 ( .A(n32592), .B(n32595), .Z(n32662) );
  IV U41558 ( .A(n32594), .Z(n32595) );
  NAND U41559 ( .A(n32663), .B(n32664), .Z(n32594) );
  OR U41560 ( .A(n32665), .B(n32666), .Z(n32664) );
  OR U41561 ( .A(n32667), .B(n32668), .Z(n32663) );
  NAND U41562 ( .A(n32669), .B(n32670), .Z(n32592) );
  OR U41563 ( .A(n32671), .B(n32672), .Z(n32670) );
  OR U41564 ( .A(n32673), .B(n32674), .Z(n32669) );
  NOR U41565 ( .A(n32675), .B(n32676), .Z(n32593) );
  ANDN U41566 ( .B(n32677), .A(n32678), .Z(n32587) );
  IV U41567 ( .A(n32679), .Z(n32677) );
  XNOR U41568 ( .A(n32580), .B(n32680), .Z(n32586) );
  XNOR U41569 ( .A(n32579), .B(n32581), .Z(n32680) );
  NAND U41570 ( .A(n32681), .B(n32682), .Z(n32581) );
  OR U41571 ( .A(n32683), .B(n32684), .Z(n32682) );
  OR U41572 ( .A(n32685), .B(n32686), .Z(n32681) );
  NAND U41573 ( .A(n32687), .B(n32688), .Z(n32579) );
  OR U41574 ( .A(n32689), .B(n32690), .Z(n32688) );
  OR U41575 ( .A(n32691), .B(n32692), .Z(n32687) );
  ANDN U41576 ( .B(n32693), .A(n32694), .Z(n32580) );
  IV U41577 ( .A(n32695), .Z(n32693) );
  XNOR U41578 ( .A(n32660), .B(n32659), .Z(N62503) );
  XOR U41579 ( .A(n32679), .B(n32678), .Z(n32659) );
  XNOR U41580 ( .A(n32694), .B(n32695), .Z(n32678) );
  XNOR U41581 ( .A(n32689), .B(n32690), .Z(n32695) );
  XNOR U41582 ( .A(n32691), .B(n32692), .Z(n32690) );
  XNOR U41583 ( .A(y[3541]), .B(x[3541]), .Z(n32692) );
  XNOR U41584 ( .A(y[3542]), .B(x[3542]), .Z(n32691) );
  XNOR U41585 ( .A(y[3540]), .B(x[3540]), .Z(n32689) );
  XNOR U41586 ( .A(n32683), .B(n32684), .Z(n32694) );
  XNOR U41587 ( .A(y[3537]), .B(x[3537]), .Z(n32684) );
  XNOR U41588 ( .A(n32685), .B(n32686), .Z(n32683) );
  XNOR U41589 ( .A(y[3538]), .B(x[3538]), .Z(n32686) );
  XNOR U41590 ( .A(y[3539]), .B(x[3539]), .Z(n32685) );
  XNOR U41591 ( .A(n32676), .B(n32675), .Z(n32679) );
  XNOR U41592 ( .A(n32671), .B(n32672), .Z(n32675) );
  XNOR U41593 ( .A(y[3534]), .B(x[3534]), .Z(n32672) );
  XNOR U41594 ( .A(n32673), .B(n32674), .Z(n32671) );
  XNOR U41595 ( .A(y[3535]), .B(x[3535]), .Z(n32674) );
  XNOR U41596 ( .A(y[3536]), .B(x[3536]), .Z(n32673) );
  XNOR U41597 ( .A(n32665), .B(n32666), .Z(n32676) );
  XNOR U41598 ( .A(y[3531]), .B(x[3531]), .Z(n32666) );
  XNOR U41599 ( .A(n32667), .B(n32668), .Z(n32665) );
  XNOR U41600 ( .A(y[3532]), .B(x[3532]), .Z(n32668) );
  XNOR U41601 ( .A(y[3533]), .B(x[3533]), .Z(n32667) );
  XOR U41602 ( .A(n32641), .B(n32642), .Z(n32660) );
  XNOR U41603 ( .A(n32657), .B(n32658), .Z(n32642) );
  XNOR U41604 ( .A(n32652), .B(n32653), .Z(n32658) );
  XNOR U41605 ( .A(n32654), .B(n32655), .Z(n32653) );
  XNOR U41606 ( .A(y[3529]), .B(x[3529]), .Z(n32655) );
  XNOR U41607 ( .A(y[3530]), .B(x[3530]), .Z(n32654) );
  XNOR U41608 ( .A(y[3528]), .B(x[3528]), .Z(n32652) );
  XNOR U41609 ( .A(n32646), .B(n32647), .Z(n32657) );
  XNOR U41610 ( .A(y[3525]), .B(x[3525]), .Z(n32647) );
  XNOR U41611 ( .A(n32648), .B(n32649), .Z(n32646) );
  XNOR U41612 ( .A(y[3526]), .B(x[3526]), .Z(n32649) );
  XNOR U41613 ( .A(y[3527]), .B(x[3527]), .Z(n32648) );
  XOR U41614 ( .A(n32640), .B(n32639), .Z(n32641) );
  XNOR U41615 ( .A(n32635), .B(n32636), .Z(n32639) );
  XNOR U41616 ( .A(y[3522]), .B(x[3522]), .Z(n32636) );
  XNOR U41617 ( .A(n32637), .B(n32638), .Z(n32635) );
  XNOR U41618 ( .A(y[3523]), .B(x[3523]), .Z(n32638) );
  XNOR U41619 ( .A(y[3524]), .B(x[3524]), .Z(n32637) );
  XNOR U41620 ( .A(n32629), .B(n32630), .Z(n32640) );
  XNOR U41621 ( .A(y[3519]), .B(x[3519]), .Z(n32630) );
  XNOR U41622 ( .A(n32631), .B(n32632), .Z(n32629) );
  XNOR U41623 ( .A(y[3520]), .B(x[3520]), .Z(n32632) );
  XNOR U41624 ( .A(y[3521]), .B(x[3521]), .Z(n32631) );
  NAND U41625 ( .A(n32696), .B(n32697), .Z(N62494) );
  NANDN U41626 ( .A(n32698), .B(n32699), .Z(n32697) );
  OR U41627 ( .A(n32700), .B(n32701), .Z(n32699) );
  NAND U41628 ( .A(n32700), .B(n32701), .Z(n32696) );
  XOR U41629 ( .A(n32700), .B(n32702), .Z(N62493) );
  XNOR U41630 ( .A(n32698), .B(n32701), .Z(n32702) );
  AND U41631 ( .A(n32703), .B(n32704), .Z(n32701) );
  NANDN U41632 ( .A(n32705), .B(n32706), .Z(n32704) );
  NANDN U41633 ( .A(n32707), .B(n32708), .Z(n32706) );
  NANDN U41634 ( .A(n32708), .B(n32707), .Z(n32703) );
  NAND U41635 ( .A(n32709), .B(n32710), .Z(n32698) );
  NANDN U41636 ( .A(n32711), .B(n32712), .Z(n32710) );
  OR U41637 ( .A(n32713), .B(n32714), .Z(n32712) );
  NAND U41638 ( .A(n32714), .B(n32713), .Z(n32709) );
  AND U41639 ( .A(n32715), .B(n32716), .Z(n32700) );
  NANDN U41640 ( .A(n32717), .B(n32718), .Z(n32716) );
  NANDN U41641 ( .A(n32719), .B(n32720), .Z(n32718) );
  NANDN U41642 ( .A(n32720), .B(n32719), .Z(n32715) );
  XOR U41643 ( .A(n32714), .B(n32721), .Z(N62492) );
  XOR U41644 ( .A(n32711), .B(n32713), .Z(n32721) );
  XNOR U41645 ( .A(n32707), .B(n32722), .Z(n32713) );
  XNOR U41646 ( .A(n32705), .B(n32708), .Z(n32722) );
  NAND U41647 ( .A(n32723), .B(n32724), .Z(n32708) );
  NAND U41648 ( .A(n32725), .B(n32726), .Z(n32724) );
  OR U41649 ( .A(n32727), .B(n32728), .Z(n32725) );
  NANDN U41650 ( .A(n32729), .B(n32727), .Z(n32723) );
  IV U41651 ( .A(n32728), .Z(n32729) );
  NAND U41652 ( .A(n32730), .B(n32731), .Z(n32705) );
  NAND U41653 ( .A(n32732), .B(n32733), .Z(n32731) );
  NANDN U41654 ( .A(n32734), .B(n32735), .Z(n32732) );
  NANDN U41655 ( .A(n32735), .B(n32734), .Z(n32730) );
  AND U41656 ( .A(n32736), .B(n32737), .Z(n32707) );
  NAND U41657 ( .A(n32738), .B(n32739), .Z(n32737) );
  OR U41658 ( .A(n32740), .B(n32741), .Z(n32738) );
  NANDN U41659 ( .A(n32742), .B(n32740), .Z(n32736) );
  NAND U41660 ( .A(n32743), .B(n32744), .Z(n32711) );
  NANDN U41661 ( .A(n32745), .B(n32746), .Z(n32744) );
  OR U41662 ( .A(n32747), .B(n32748), .Z(n32746) );
  NANDN U41663 ( .A(n32749), .B(n32747), .Z(n32743) );
  IV U41664 ( .A(n32748), .Z(n32749) );
  XNOR U41665 ( .A(n32719), .B(n32750), .Z(n32714) );
  XNOR U41666 ( .A(n32717), .B(n32720), .Z(n32750) );
  NAND U41667 ( .A(n32751), .B(n32752), .Z(n32720) );
  NAND U41668 ( .A(n32753), .B(n32754), .Z(n32752) );
  OR U41669 ( .A(n32755), .B(n32756), .Z(n32753) );
  NANDN U41670 ( .A(n32757), .B(n32755), .Z(n32751) );
  IV U41671 ( .A(n32756), .Z(n32757) );
  NAND U41672 ( .A(n32758), .B(n32759), .Z(n32717) );
  NAND U41673 ( .A(n32760), .B(n32761), .Z(n32759) );
  NANDN U41674 ( .A(n32762), .B(n32763), .Z(n32760) );
  NANDN U41675 ( .A(n32763), .B(n32762), .Z(n32758) );
  AND U41676 ( .A(n32764), .B(n32765), .Z(n32719) );
  NAND U41677 ( .A(n32766), .B(n32767), .Z(n32765) );
  OR U41678 ( .A(n32768), .B(n32769), .Z(n32766) );
  NANDN U41679 ( .A(n32770), .B(n32768), .Z(n32764) );
  XNOR U41680 ( .A(n32745), .B(n32771), .Z(N62491) );
  XOR U41681 ( .A(n32747), .B(n32748), .Z(n32771) );
  XNOR U41682 ( .A(n32761), .B(n32772), .Z(n32748) );
  XOR U41683 ( .A(n32762), .B(n32763), .Z(n32772) );
  XOR U41684 ( .A(n32768), .B(n32773), .Z(n32763) );
  XOR U41685 ( .A(n32767), .B(n32770), .Z(n32773) );
  IV U41686 ( .A(n32769), .Z(n32770) );
  NAND U41687 ( .A(n32774), .B(n32775), .Z(n32769) );
  OR U41688 ( .A(n32776), .B(n32777), .Z(n32775) );
  OR U41689 ( .A(n32778), .B(n32779), .Z(n32774) );
  NAND U41690 ( .A(n32780), .B(n32781), .Z(n32767) );
  OR U41691 ( .A(n32782), .B(n32783), .Z(n32781) );
  OR U41692 ( .A(n32784), .B(n32785), .Z(n32780) );
  NOR U41693 ( .A(n32786), .B(n32787), .Z(n32768) );
  ANDN U41694 ( .B(n32788), .A(n32789), .Z(n32762) );
  XNOR U41695 ( .A(n32755), .B(n32790), .Z(n32761) );
  XNOR U41696 ( .A(n32754), .B(n32756), .Z(n32790) );
  NAND U41697 ( .A(n32791), .B(n32792), .Z(n32756) );
  OR U41698 ( .A(n32793), .B(n32794), .Z(n32792) );
  OR U41699 ( .A(n32795), .B(n32796), .Z(n32791) );
  NAND U41700 ( .A(n32797), .B(n32798), .Z(n32754) );
  OR U41701 ( .A(n32799), .B(n32800), .Z(n32798) );
  OR U41702 ( .A(n32801), .B(n32802), .Z(n32797) );
  ANDN U41703 ( .B(n32803), .A(n32804), .Z(n32755) );
  IV U41704 ( .A(n32805), .Z(n32803) );
  ANDN U41705 ( .B(n32806), .A(n32807), .Z(n32747) );
  XOR U41706 ( .A(n32733), .B(n32808), .Z(n32745) );
  XOR U41707 ( .A(n32734), .B(n32735), .Z(n32808) );
  XOR U41708 ( .A(n32740), .B(n32809), .Z(n32735) );
  XOR U41709 ( .A(n32739), .B(n32742), .Z(n32809) );
  IV U41710 ( .A(n32741), .Z(n32742) );
  NAND U41711 ( .A(n32810), .B(n32811), .Z(n32741) );
  OR U41712 ( .A(n32812), .B(n32813), .Z(n32811) );
  OR U41713 ( .A(n32814), .B(n32815), .Z(n32810) );
  NAND U41714 ( .A(n32816), .B(n32817), .Z(n32739) );
  OR U41715 ( .A(n32818), .B(n32819), .Z(n32817) );
  OR U41716 ( .A(n32820), .B(n32821), .Z(n32816) );
  NOR U41717 ( .A(n32822), .B(n32823), .Z(n32740) );
  ANDN U41718 ( .B(n32824), .A(n32825), .Z(n32734) );
  IV U41719 ( .A(n32826), .Z(n32824) );
  XNOR U41720 ( .A(n32727), .B(n32827), .Z(n32733) );
  XNOR U41721 ( .A(n32726), .B(n32728), .Z(n32827) );
  NAND U41722 ( .A(n32828), .B(n32829), .Z(n32728) );
  OR U41723 ( .A(n32830), .B(n32831), .Z(n32829) );
  OR U41724 ( .A(n32832), .B(n32833), .Z(n32828) );
  NAND U41725 ( .A(n32834), .B(n32835), .Z(n32726) );
  OR U41726 ( .A(n32836), .B(n32837), .Z(n32835) );
  OR U41727 ( .A(n32838), .B(n32839), .Z(n32834) );
  ANDN U41728 ( .B(n32840), .A(n32841), .Z(n32727) );
  IV U41729 ( .A(n32842), .Z(n32840) );
  XNOR U41730 ( .A(n32807), .B(n32806), .Z(N62490) );
  XOR U41731 ( .A(n32826), .B(n32825), .Z(n32806) );
  XNOR U41732 ( .A(n32841), .B(n32842), .Z(n32825) );
  XNOR U41733 ( .A(n32836), .B(n32837), .Z(n32842) );
  XNOR U41734 ( .A(n32838), .B(n32839), .Z(n32837) );
  XNOR U41735 ( .A(y[3517]), .B(x[3517]), .Z(n32839) );
  XNOR U41736 ( .A(y[3518]), .B(x[3518]), .Z(n32838) );
  XNOR U41737 ( .A(y[3516]), .B(x[3516]), .Z(n32836) );
  XNOR U41738 ( .A(n32830), .B(n32831), .Z(n32841) );
  XNOR U41739 ( .A(y[3513]), .B(x[3513]), .Z(n32831) );
  XNOR U41740 ( .A(n32832), .B(n32833), .Z(n32830) );
  XNOR U41741 ( .A(y[3514]), .B(x[3514]), .Z(n32833) );
  XNOR U41742 ( .A(y[3515]), .B(x[3515]), .Z(n32832) );
  XNOR U41743 ( .A(n32823), .B(n32822), .Z(n32826) );
  XNOR U41744 ( .A(n32818), .B(n32819), .Z(n32822) );
  XNOR U41745 ( .A(y[3510]), .B(x[3510]), .Z(n32819) );
  XNOR U41746 ( .A(n32820), .B(n32821), .Z(n32818) );
  XNOR U41747 ( .A(y[3511]), .B(x[3511]), .Z(n32821) );
  XNOR U41748 ( .A(y[3512]), .B(x[3512]), .Z(n32820) );
  XNOR U41749 ( .A(n32812), .B(n32813), .Z(n32823) );
  XNOR U41750 ( .A(y[3507]), .B(x[3507]), .Z(n32813) );
  XNOR U41751 ( .A(n32814), .B(n32815), .Z(n32812) );
  XNOR U41752 ( .A(y[3508]), .B(x[3508]), .Z(n32815) );
  XNOR U41753 ( .A(y[3509]), .B(x[3509]), .Z(n32814) );
  XOR U41754 ( .A(n32788), .B(n32789), .Z(n32807) );
  XNOR U41755 ( .A(n32804), .B(n32805), .Z(n32789) );
  XNOR U41756 ( .A(n32799), .B(n32800), .Z(n32805) );
  XNOR U41757 ( .A(n32801), .B(n32802), .Z(n32800) );
  XNOR U41758 ( .A(y[3505]), .B(x[3505]), .Z(n32802) );
  XNOR U41759 ( .A(y[3506]), .B(x[3506]), .Z(n32801) );
  XNOR U41760 ( .A(y[3504]), .B(x[3504]), .Z(n32799) );
  XNOR U41761 ( .A(n32793), .B(n32794), .Z(n32804) );
  XNOR U41762 ( .A(y[3501]), .B(x[3501]), .Z(n32794) );
  XNOR U41763 ( .A(n32795), .B(n32796), .Z(n32793) );
  XNOR U41764 ( .A(y[3502]), .B(x[3502]), .Z(n32796) );
  XNOR U41765 ( .A(y[3503]), .B(x[3503]), .Z(n32795) );
  XOR U41766 ( .A(n32787), .B(n32786), .Z(n32788) );
  XNOR U41767 ( .A(n32782), .B(n32783), .Z(n32786) );
  XNOR U41768 ( .A(y[3498]), .B(x[3498]), .Z(n32783) );
  XNOR U41769 ( .A(n32784), .B(n32785), .Z(n32782) );
  XNOR U41770 ( .A(y[3499]), .B(x[3499]), .Z(n32785) );
  XNOR U41771 ( .A(y[3500]), .B(x[3500]), .Z(n32784) );
  XNOR U41772 ( .A(n32776), .B(n32777), .Z(n32787) );
  XNOR U41773 ( .A(y[3495]), .B(x[3495]), .Z(n32777) );
  XNOR U41774 ( .A(n32778), .B(n32779), .Z(n32776) );
  XNOR U41775 ( .A(y[3496]), .B(x[3496]), .Z(n32779) );
  XNOR U41776 ( .A(y[3497]), .B(x[3497]), .Z(n32778) );
  NAND U41777 ( .A(n32843), .B(n32844), .Z(N62481) );
  NANDN U41778 ( .A(n32845), .B(n32846), .Z(n32844) );
  OR U41779 ( .A(n32847), .B(n32848), .Z(n32846) );
  NAND U41780 ( .A(n32847), .B(n32848), .Z(n32843) );
  XOR U41781 ( .A(n32847), .B(n32849), .Z(N62480) );
  XNOR U41782 ( .A(n32845), .B(n32848), .Z(n32849) );
  AND U41783 ( .A(n32850), .B(n32851), .Z(n32848) );
  NANDN U41784 ( .A(n32852), .B(n32853), .Z(n32851) );
  NANDN U41785 ( .A(n32854), .B(n32855), .Z(n32853) );
  NANDN U41786 ( .A(n32855), .B(n32854), .Z(n32850) );
  NAND U41787 ( .A(n32856), .B(n32857), .Z(n32845) );
  NANDN U41788 ( .A(n32858), .B(n32859), .Z(n32857) );
  OR U41789 ( .A(n32860), .B(n32861), .Z(n32859) );
  NAND U41790 ( .A(n32861), .B(n32860), .Z(n32856) );
  AND U41791 ( .A(n32862), .B(n32863), .Z(n32847) );
  NANDN U41792 ( .A(n32864), .B(n32865), .Z(n32863) );
  NANDN U41793 ( .A(n32866), .B(n32867), .Z(n32865) );
  NANDN U41794 ( .A(n32867), .B(n32866), .Z(n32862) );
  XOR U41795 ( .A(n32861), .B(n32868), .Z(N62479) );
  XOR U41796 ( .A(n32858), .B(n32860), .Z(n32868) );
  XNOR U41797 ( .A(n32854), .B(n32869), .Z(n32860) );
  XNOR U41798 ( .A(n32852), .B(n32855), .Z(n32869) );
  NAND U41799 ( .A(n32870), .B(n32871), .Z(n32855) );
  NAND U41800 ( .A(n32872), .B(n32873), .Z(n32871) );
  OR U41801 ( .A(n32874), .B(n32875), .Z(n32872) );
  NANDN U41802 ( .A(n32876), .B(n32874), .Z(n32870) );
  IV U41803 ( .A(n32875), .Z(n32876) );
  NAND U41804 ( .A(n32877), .B(n32878), .Z(n32852) );
  NAND U41805 ( .A(n32879), .B(n32880), .Z(n32878) );
  NANDN U41806 ( .A(n32881), .B(n32882), .Z(n32879) );
  NANDN U41807 ( .A(n32882), .B(n32881), .Z(n32877) );
  AND U41808 ( .A(n32883), .B(n32884), .Z(n32854) );
  NAND U41809 ( .A(n32885), .B(n32886), .Z(n32884) );
  OR U41810 ( .A(n32887), .B(n32888), .Z(n32885) );
  NANDN U41811 ( .A(n32889), .B(n32887), .Z(n32883) );
  NAND U41812 ( .A(n32890), .B(n32891), .Z(n32858) );
  NANDN U41813 ( .A(n32892), .B(n32893), .Z(n32891) );
  OR U41814 ( .A(n32894), .B(n32895), .Z(n32893) );
  NANDN U41815 ( .A(n32896), .B(n32894), .Z(n32890) );
  IV U41816 ( .A(n32895), .Z(n32896) );
  XNOR U41817 ( .A(n32866), .B(n32897), .Z(n32861) );
  XNOR U41818 ( .A(n32864), .B(n32867), .Z(n32897) );
  NAND U41819 ( .A(n32898), .B(n32899), .Z(n32867) );
  NAND U41820 ( .A(n32900), .B(n32901), .Z(n32899) );
  OR U41821 ( .A(n32902), .B(n32903), .Z(n32900) );
  NANDN U41822 ( .A(n32904), .B(n32902), .Z(n32898) );
  IV U41823 ( .A(n32903), .Z(n32904) );
  NAND U41824 ( .A(n32905), .B(n32906), .Z(n32864) );
  NAND U41825 ( .A(n32907), .B(n32908), .Z(n32906) );
  NANDN U41826 ( .A(n32909), .B(n32910), .Z(n32907) );
  NANDN U41827 ( .A(n32910), .B(n32909), .Z(n32905) );
  AND U41828 ( .A(n32911), .B(n32912), .Z(n32866) );
  NAND U41829 ( .A(n32913), .B(n32914), .Z(n32912) );
  OR U41830 ( .A(n32915), .B(n32916), .Z(n32913) );
  NANDN U41831 ( .A(n32917), .B(n32915), .Z(n32911) );
  XNOR U41832 ( .A(n32892), .B(n32918), .Z(N62478) );
  XOR U41833 ( .A(n32894), .B(n32895), .Z(n32918) );
  XNOR U41834 ( .A(n32908), .B(n32919), .Z(n32895) );
  XOR U41835 ( .A(n32909), .B(n32910), .Z(n32919) );
  XOR U41836 ( .A(n32915), .B(n32920), .Z(n32910) );
  XOR U41837 ( .A(n32914), .B(n32917), .Z(n32920) );
  IV U41838 ( .A(n32916), .Z(n32917) );
  NAND U41839 ( .A(n32921), .B(n32922), .Z(n32916) );
  OR U41840 ( .A(n32923), .B(n32924), .Z(n32922) );
  OR U41841 ( .A(n32925), .B(n32926), .Z(n32921) );
  NAND U41842 ( .A(n32927), .B(n32928), .Z(n32914) );
  OR U41843 ( .A(n32929), .B(n32930), .Z(n32928) );
  OR U41844 ( .A(n32931), .B(n32932), .Z(n32927) );
  NOR U41845 ( .A(n32933), .B(n32934), .Z(n32915) );
  ANDN U41846 ( .B(n32935), .A(n32936), .Z(n32909) );
  XNOR U41847 ( .A(n32902), .B(n32937), .Z(n32908) );
  XNOR U41848 ( .A(n32901), .B(n32903), .Z(n32937) );
  NAND U41849 ( .A(n32938), .B(n32939), .Z(n32903) );
  OR U41850 ( .A(n32940), .B(n32941), .Z(n32939) );
  OR U41851 ( .A(n32942), .B(n32943), .Z(n32938) );
  NAND U41852 ( .A(n32944), .B(n32945), .Z(n32901) );
  OR U41853 ( .A(n32946), .B(n32947), .Z(n32945) );
  OR U41854 ( .A(n32948), .B(n32949), .Z(n32944) );
  ANDN U41855 ( .B(n32950), .A(n32951), .Z(n32902) );
  IV U41856 ( .A(n32952), .Z(n32950) );
  ANDN U41857 ( .B(n32953), .A(n32954), .Z(n32894) );
  XOR U41858 ( .A(n32880), .B(n32955), .Z(n32892) );
  XOR U41859 ( .A(n32881), .B(n32882), .Z(n32955) );
  XOR U41860 ( .A(n32887), .B(n32956), .Z(n32882) );
  XOR U41861 ( .A(n32886), .B(n32889), .Z(n32956) );
  IV U41862 ( .A(n32888), .Z(n32889) );
  NAND U41863 ( .A(n32957), .B(n32958), .Z(n32888) );
  OR U41864 ( .A(n32959), .B(n32960), .Z(n32958) );
  OR U41865 ( .A(n32961), .B(n32962), .Z(n32957) );
  NAND U41866 ( .A(n32963), .B(n32964), .Z(n32886) );
  OR U41867 ( .A(n32965), .B(n32966), .Z(n32964) );
  OR U41868 ( .A(n32967), .B(n32968), .Z(n32963) );
  NOR U41869 ( .A(n32969), .B(n32970), .Z(n32887) );
  ANDN U41870 ( .B(n32971), .A(n32972), .Z(n32881) );
  IV U41871 ( .A(n32973), .Z(n32971) );
  XNOR U41872 ( .A(n32874), .B(n32974), .Z(n32880) );
  XNOR U41873 ( .A(n32873), .B(n32875), .Z(n32974) );
  NAND U41874 ( .A(n32975), .B(n32976), .Z(n32875) );
  OR U41875 ( .A(n32977), .B(n32978), .Z(n32976) );
  OR U41876 ( .A(n32979), .B(n32980), .Z(n32975) );
  NAND U41877 ( .A(n32981), .B(n32982), .Z(n32873) );
  OR U41878 ( .A(n32983), .B(n32984), .Z(n32982) );
  OR U41879 ( .A(n32985), .B(n32986), .Z(n32981) );
  ANDN U41880 ( .B(n32987), .A(n32988), .Z(n32874) );
  IV U41881 ( .A(n32989), .Z(n32987) );
  XNOR U41882 ( .A(n32954), .B(n32953), .Z(N62477) );
  XOR U41883 ( .A(n32973), .B(n32972), .Z(n32953) );
  XNOR U41884 ( .A(n32988), .B(n32989), .Z(n32972) );
  XNOR U41885 ( .A(n32983), .B(n32984), .Z(n32989) );
  XNOR U41886 ( .A(n32985), .B(n32986), .Z(n32984) );
  XNOR U41887 ( .A(y[3493]), .B(x[3493]), .Z(n32986) );
  XNOR U41888 ( .A(y[3494]), .B(x[3494]), .Z(n32985) );
  XNOR U41889 ( .A(y[3492]), .B(x[3492]), .Z(n32983) );
  XNOR U41890 ( .A(n32977), .B(n32978), .Z(n32988) );
  XNOR U41891 ( .A(y[3489]), .B(x[3489]), .Z(n32978) );
  XNOR U41892 ( .A(n32979), .B(n32980), .Z(n32977) );
  XNOR U41893 ( .A(y[3490]), .B(x[3490]), .Z(n32980) );
  XNOR U41894 ( .A(y[3491]), .B(x[3491]), .Z(n32979) );
  XNOR U41895 ( .A(n32970), .B(n32969), .Z(n32973) );
  XNOR U41896 ( .A(n32965), .B(n32966), .Z(n32969) );
  XNOR U41897 ( .A(y[3486]), .B(x[3486]), .Z(n32966) );
  XNOR U41898 ( .A(n32967), .B(n32968), .Z(n32965) );
  XNOR U41899 ( .A(y[3487]), .B(x[3487]), .Z(n32968) );
  XNOR U41900 ( .A(y[3488]), .B(x[3488]), .Z(n32967) );
  XNOR U41901 ( .A(n32959), .B(n32960), .Z(n32970) );
  XNOR U41902 ( .A(y[3483]), .B(x[3483]), .Z(n32960) );
  XNOR U41903 ( .A(n32961), .B(n32962), .Z(n32959) );
  XNOR U41904 ( .A(y[3484]), .B(x[3484]), .Z(n32962) );
  XNOR U41905 ( .A(y[3485]), .B(x[3485]), .Z(n32961) );
  XOR U41906 ( .A(n32935), .B(n32936), .Z(n32954) );
  XNOR U41907 ( .A(n32951), .B(n32952), .Z(n32936) );
  XNOR U41908 ( .A(n32946), .B(n32947), .Z(n32952) );
  XNOR U41909 ( .A(n32948), .B(n32949), .Z(n32947) );
  XNOR U41910 ( .A(y[3481]), .B(x[3481]), .Z(n32949) );
  XNOR U41911 ( .A(y[3482]), .B(x[3482]), .Z(n32948) );
  XNOR U41912 ( .A(y[3480]), .B(x[3480]), .Z(n32946) );
  XNOR U41913 ( .A(n32940), .B(n32941), .Z(n32951) );
  XNOR U41914 ( .A(y[3477]), .B(x[3477]), .Z(n32941) );
  XNOR U41915 ( .A(n32942), .B(n32943), .Z(n32940) );
  XNOR U41916 ( .A(y[3478]), .B(x[3478]), .Z(n32943) );
  XNOR U41917 ( .A(y[3479]), .B(x[3479]), .Z(n32942) );
  XOR U41918 ( .A(n32934), .B(n32933), .Z(n32935) );
  XNOR U41919 ( .A(n32929), .B(n32930), .Z(n32933) );
  XNOR U41920 ( .A(y[3474]), .B(x[3474]), .Z(n32930) );
  XNOR U41921 ( .A(n32931), .B(n32932), .Z(n32929) );
  XNOR U41922 ( .A(y[3475]), .B(x[3475]), .Z(n32932) );
  XNOR U41923 ( .A(y[3476]), .B(x[3476]), .Z(n32931) );
  XNOR U41924 ( .A(n32923), .B(n32924), .Z(n32934) );
  XNOR U41925 ( .A(y[3471]), .B(x[3471]), .Z(n32924) );
  XNOR U41926 ( .A(n32925), .B(n32926), .Z(n32923) );
  XNOR U41927 ( .A(y[3472]), .B(x[3472]), .Z(n32926) );
  XNOR U41928 ( .A(y[3473]), .B(x[3473]), .Z(n32925) );
  NAND U41929 ( .A(n32990), .B(n32991), .Z(N62468) );
  NANDN U41930 ( .A(n32992), .B(n32993), .Z(n32991) );
  OR U41931 ( .A(n32994), .B(n32995), .Z(n32993) );
  NAND U41932 ( .A(n32994), .B(n32995), .Z(n32990) );
  XOR U41933 ( .A(n32994), .B(n32996), .Z(N62467) );
  XNOR U41934 ( .A(n32992), .B(n32995), .Z(n32996) );
  AND U41935 ( .A(n32997), .B(n32998), .Z(n32995) );
  NANDN U41936 ( .A(n32999), .B(n33000), .Z(n32998) );
  NANDN U41937 ( .A(n33001), .B(n33002), .Z(n33000) );
  NANDN U41938 ( .A(n33002), .B(n33001), .Z(n32997) );
  NAND U41939 ( .A(n33003), .B(n33004), .Z(n32992) );
  NANDN U41940 ( .A(n33005), .B(n33006), .Z(n33004) );
  OR U41941 ( .A(n33007), .B(n33008), .Z(n33006) );
  NAND U41942 ( .A(n33008), .B(n33007), .Z(n33003) );
  AND U41943 ( .A(n33009), .B(n33010), .Z(n32994) );
  NANDN U41944 ( .A(n33011), .B(n33012), .Z(n33010) );
  NANDN U41945 ( .A(n33013), .B(n33014), .Z(n33012) );
  NANDN U41946 ( .A(n33014), .B(n33013), .Z(n33009) );
  XOR U41947 ( .A(n33008), .B(n33015), .Z(N62466) );
  XOR U41948 ( .A(n33005), .B(n33007), .Z(n33015) );
  XNOR U41949 ( .A(n33001), .B(n33016), .Z(n33007) );
  XNOR U41950 ( .A(n32999), .B(n33002), .Z(n33016) );
  NAND U41951 ( .A(n33017), .B(n33018), .Z(n33002) );
  NAND U41952 ( .A(n33019), .B(n33020), .Z(n33018) );
  OR U41953 ( .A(n33021), .B(n33022), .Z(n33019) );
  NANDN U41954 ( .A(n33023), .B(n33021), .Z(n33017) );
  IV U41955 ( .A(n33022), .Z(n33023) );
  NAND U41956 ( .A(n33024), .B(n33025), .Z(n32999) );
  NAND U41957 ( .A(n33026), .B(n33027), .Z(n33025) );
  NANDN U41958 ( .A(n33028), .B(n33029), .Z(n33026) );
  NANDN U41959 ( .A(n33029), .B(n33028), .Z(n33024) );
  AND U41960 ( .A(n33030), .B(n33031), .Z(n33001) );
  NAND U41961 ( .A(n33032), .B(n33033), .Z(n33031) );
  OR U41962 ( .A(n33034), .B(n33035), .Z(n33032) );
  NANDN U41963 ( .A(n33036), .B(n33034), .Z(n33030) );
  NAND U41964 ( .A(n33037), .B(n33038), .Z(n33005) );
  NANDN U41965 ( .A(n33039), .B(n33040), .Z(n33038) );
  OR U41966 ( .A(n33041), .B(n33042), .Z(n33040) );
  NANDN U41967 ( .A(n33043), .B(n33041), .Z(n33037) );
  IV U41968 ( .A(n33042), .Z(n33043) );
  XNOR U41969 ( .A(n33013), .B(n33044), .Z(n33008) );
  XNOR U41970 ( .A(n33011), .B(n33014), .Z(n33044) );
  NAND U41971 ( .A(n33045), .B(n33046), .Z(n33014) );
  NAND U41972 ( .A(n33047), .B(n33048), .Z(n33046) );
  OR U41973 ( .A(n33049), .B(n33050), .Z(n33047) );
  NANDN U41974 ( .A(n33051), .B(n33049), .Z(n33045) );
  IV U41975 ( .A(n33050), .Z(n33051) );
  NAND U41976 ( .A(n33052), .B(n33053), .Z(n33011) );
  NAND U41977 ( .A(n33054), .B(n33055), .Z(n33053) );
  NANDN U41978 ( .A(n33056), .B(n33057), .Z(n33054) );
  NANDN U41979 ( .A(n33057), .B(n33056), .Z(n33052) );
  AND U41980 ( .A(n33058), .B(n33059), .Z(n33013) );
  NAND U41981 ( .A(n33060), .B(n33061), .Z(n33059) );
  OR U41982 ( .A(n33062), .B(n33063), .Z(n33060) );
  NANDN U41983 ( .A(n33064), .B(n33062), .Z(n33058) );
  XNOR U41984 ( .A(n33039), .B(n33065), .Z(N62465) );
  XOR U41985 ( .A(n33041), .B(n33042), .Z(n33065) );
  XNOR U41986 ( .A(n33055), .B(n33066), .Z(n33042) );
  XOR U41987 ( .A(n33056), .B(n33057), .Z(n33066) );
  XOR U41988 ( .A(n33062), .B(n33067), .Z(n33057) );
  XOR U41989 ( .A(n33061), .B(n33064), .Z(n33067) );
  IV U41990 ( .A(n33063), .Z(n33064) );
  NAND U41991 ( .A(n33068), .B(n33069), .Z(n33063) );
  OR U41992 ( .A(n33070), .B(n33071), .Z(n33069) );
  OR U41993 ( .A(n33072), .B(n33073), .Z(n33068) );
  NAND U41994 ( .A(n33074), .B(n33075), .Z(n33061) );
  OR U41995 ( .A(n33076), .B(n33077), .Z(n33075) );
  OR U41996 ( .A(n33078), .B(n33079), .Z(n33074) );
  NOR U41997 ( .A(n33080), .B(n33081), .Z(n33062) );
  ANDN U41998 ( .B(n33082), .A(n33083), .Z(n33056) );
  XNOR U41999 ( .A(n33049), .B(n33084), .Z(n33055) );
  XNOR U42000 ( .A(n33048), .B(n33050), .Z(n33084) );
  NAND U42001 ( .A(n33085), .B(n33086), .Z(n33050) );
  OR U42002 ( .A(n33087), .B(n33088), .Z(n33086) );
  OR U42003 ( .A(n33089), .B(n33090), .Z(n33085) );
  NAND U42004 ( .A(n33091), .B(n33092), .Z(n33048) );
  OR U42005 ( .A(n33093), .B(n33094), .Z(n33092) );
  OR U42006 ( .A(n33095), .B(n33096), .Z(n33091) );
  ANDN U42007 ( .B(n33097), .A(n33098), .Z(n33049) );
  IV U42008 ( .A(n33099), .Z(n33097) );
  ANDN U42009 ( .B(n33100), .A(n33101), .Z(n33041) );
  XOR U42010 ( .A(n33027), .B(n33102), .Z(n33039) );
  XOR U42011 ( .A(n33028), .B(n33029), .Z(n33102) );
  XOR U42012 ( .A(n33034), .B(n33103), .Z(n33029) );
  XOR U42013 ( .A(n33033), .B(n33036), .Z(n33103) );
  IV U42014 ( .A(n33035), .Z(n33036) );
  NAND U42015 ( .A(n33104), .B(n33105), .Z(n33035) );
  OR U42016 ( .A(n33106), .B(n33107), .Z(n33105) );
  OR U42017 ( .A(n33108), .B(n33109), .Z(n33104) );
  NAND U42018 ( .A(n33110), .B(n33111), .Z(n33033) );
  OR U42019 ( .A(n33112), .B(n33113), .Z(n33111) );
  OR U42020 ( .A(n33114), .B(n33115), .Z(n33110) );
  NOR U42021 ( .A(n33116), .B(n33117), .Z(n33034) );
  ANDN U42022 ( .B(n33118), .A(n33119), .Z(n33028) );
  IV U42023 ( .A(n33120), .Z(n33118) );
  XNOR U42024 ( .A(n33021), .B(n33121), .Z(n33027) );
  XNOR U42025 ( .A(n33020), .B(n33022), .Z(n33121) );
  NAND U42026 ( .A(n33122), .B(n33123), .Z(n33022) );
  OR U42027 ( .A(n33124), .B(n33125), .Z(n33123) );
  OR U42028 ( .A(n33126), .B(n33127), .Z(n33122) );
  NAND U42029 ( .A(n33128), .B(n33129), .Z(n33020) );
  OR U42030 ( .A(n33130), .B(n33131), .Z(n33129) );
  OR U42031 ( .A(n33132), .B(n33133), .Z(n33128) );
  ANDN U42032 ( .B(n33134), .A(n33135), .Z(n33021) );
  IV U42033 ( .A(n33136), .Z(n33134) );
  XNOR U42034 ( .A(n33101), .B(n33100), .Z(N62464) );
  XOR U42035 ( .A(n33120), .B(n33119), .Z(n33100) );
  XNOR U42036 ( .A(n33135), .B(n33136), .Z(n33119) );
  XNOR U42037 ( .A(n33130), .B(n33131), .Z(n33136) );
  XNOR U42038 ( .A(n33132), .B(n33133), .Z(n33131) );
  XNOR U42039 ( .A(y[3469]), .B(x[3469]), .Z(n33133) );
  XNOR U42040 ( .A(y[3470]), .B(x[3470]), .Z(n33132) );
  XNOR U42041 ( .A(y[3468]), .B(x[3468]), .Z(n33130) );
  XNOR U42042 ( .A(n33124), .B(n33125), .Z(n33135) );
  XNOR U42043 ( .A(y[3465]), .B(x[3465]), .Z(n33125) );
  XNOR U42044 ( .A(n33126), .B(n33127), .Z(n33124) );
  XNOR U42045 ( .A(y[3466]), .B(x[3466]), .Z(n33127) );
  XNOR U42046 ( .A(y[3467]), .B(x[3467]), .Z(n33126) );
  XNOR U42047 ( .A(n33117), .B(n33116), .Z(n33120) );
  XNOR U42048 ( .A(n33112), .B(n33113), .Z(n33116) );
  XNOR U42049 ( .A(y[3462]), .B(x[3462]), .Z(n33113) );
  XNOR U42050 ( .A(n33114), .B(n33115), .Z(n33112) );
  XNOR U42051 ( .A(y[3463]), .B(x[3463]), .Z(n33115) );
  XNOR U42052 ( .A(y[3464]), .B(x[3464]), .Z(n33114) );
  XNOR U42053 ( .A(n33106), .B(n33107), .Z(n33117) );
  XNOR U42054 ( .A(y[3459]), .B(x[3459]), .Z(n33107) );
  XNOR U42055 ( .A(n33108), .B(n33109), .Z(n33106) );
  XNOR U42056 ( .A(y[3460]), .B(x[3460]), .Z(n33109) );
  XNOR U42057 ( .A(y[3461]), .B(x[3461]), .Z(n33108) );
  XOR U42058 ( .A(n33082), .B(n33083), .Z(n33101) );
  XNOR U42059 ( .A(n33098), .B(n33099), .Z(n33083) );
  XNOR U42060 ( .A(n33093), .B(n33094), .Z(n33099) );
  XNOR U42061 ( .A(n33095), .B(n33096), .Z(n33094) );
  XNOR U42062 ( .A(y[3457]), .B(x[3457]), .Z(n33096) );
  XNOR U42063 ( .A(y[3458]), .B(x[3458]), .Z(n33095) );
  XNOR U42064 ( .A(y[3456]), .B(x[3456]), .Z(n33093) );
  XNOR U42065 ( .A(n33087), .B(n33088), .Z(n33098) );
  XNOR U42066 ( .A(y[3453]), .B(x[3453]), .Z(n33088) );
  XNOR U42067 ( .A(n33089), .B(n33090), .Z(n33087) );
  XNOR U42068 ( .A(y[3454]), .B(x[3454]), .Z(n33090) );
  XNOR U42069 ( .A(y[3455]), .B(x[3455]), .Z(n33089) );
  XOR U42070 ( .A(n33081), .B(n33080), .Z(n33082) );
  XNOR U42071 ( .A(n33076), .B(n33077), .Z(n33080) );
  XNOR U42072 ( .A(y[3450]), .B(x[3450]), .Z(n33077) );
  XNOR U42073 ( .A(n33078), .B(n33079), .Z(n33076) );
  XNOR U42074 ( .A(y[3451]), .B(x[3451]), .Z(n33079) );
  XNOR U42075 ( .A(y[3452]), .B(x[3452]), .Z(n33078) );
  XNOR U42076 ( .A(n33070), .B(n33071), .Z(n33081) );
  XNOR U42077 ( .A(y[3447]), .B(x[3447]), .Z(n33071) );
  XNOR U42078 ( .A(n33072), .B(n33073), .Z(n33070) );
  XNOR U42079 ( .A(y[3448]), .B(x[3448]), .Z(n33073) );
  XNOR U42080 ( .A(y[3449]), .B(x[3449]), .Z(n33072) );
  NAND U42081 ( .A(n33137), .B(n33138), .Z(N62455) );
  NANDN U42082 ( .A(n33139), .B(n33140), .Z(n33138) );
  OR U42083 ( .A(n33141), .B(n33142), .Z(n33140) );
  NAND U42084 ( .A(n33141), .B(n33142), .Z(n33137) );
  XOR U42085 ( .A(n33141), .B(n33143), .Z(N62454) );
  XNOR U42086 ( .A(n33139), .B(n33142), .Z(n33143) );
  AND U42087 ( .A(n33144), .B(n33145), .Z(n33142) );
  NANDN U42088 ( .A(n33146), .B(n33147), .Z(n33145) );
  NANDN U42089 ( .A(n33148), .B(n33149), .Z(n33147) );
  NANDN U42090 ( .A(n33149), .B(n33148), .Z(n33144) );
  NAND U42091 ( .A(n33150), .B(n33151), .Z(n33139) );
  NANDN U42092 ( .A(n33152), .B(n33153), .Z(n33151) );
  OR U42093 ( .A(n33154), .B(n33155), .Z(n33153) );
  NAND U42094 ( .A(n33155), .B(n33154), .Z(n33150) );
  AND U42095 ( .A(n33156), .B(n33157), .Z(n33141) );
  NANDN U42096 ( .A(n33158), .B(n33159), .Z(n33157) );
  NANDN U42097 ( .A(n33160), .B(n33161), .Z(n33159) );
  NANDN U42098 ( .A(n33161), .B(n33160), .Z(n33156) );
  XOR U42099 ( .A(n33155), .B(n33162), .Z(N62453) );
  XOR U42100 ( .A(n33152), .B(n33154), .Z(n33162) );
  XNOR U42101 ( .A(n33148), .B(n33163), .Z(n33154) );
  XNOR U42102 ( .A(n33146), .B(n33149), .Z(n33163) );
  NAND U42103 ( .A(n33164), .B(n33165), .Z(n33149) );
  NAND U42104 ( .A(n33166), .B(n33167), .Z(n33165) );
  OR U42105 ( .A(n33168), .B(n33169), .Z(n33166) );
  NANDN U42106 ( .A(n33170), .B(n33168), .Z(n33164) );
  IV U42107 ( .A(n33169), .Z(n33170) );
  NAND U42108 ( .A(n33171), .B(n33172), .Z(n33146) );
  NAND U42109 ( .A(n33173), .B(n33174), .Z(n33172) );
  NANDN U42110 ( .A(n33175), .B(n33176), .Z(n33173) );
  NANDN U42111 ( .A(n33176), .B(n33175), .Z(n33171) );
  AND U42112 ( .A(n33177), .B(n33178), .Z(n33148) );
  NAND U42113 ( .A(n33179), .B(n33180), .Z(n33178) );
  OR U42114 ( .A(n33181), .B(n33182), .Z(n33179) );
  NANDN U42115 ( .A(n33183), .B(n33181), .Z(n33177) );
  NAND U42116 ( .A(n33184), .B(n33185), .Z(n33152) );
  NANDN U42117 ( .A(n33186), .B(n33187), .Z(n33185) );
  OR U42118 ( .A(n33188), .B(n33189), .Z(n33187) );
  NANDN U42119 ( .A(n33190), .B(n33188), .Z(n33184) );
  IV U42120 ( .A(n33189), .Z(n33190) );
  XNOR U42121 ( .A(n33160), .B(n33191), .Z(n33155) );
  XNOR U42122 ( .A(n33158), .B(n33161), .Z(n33191) );
  NAND U42123 ( .A(n33192), .B(n33193), .Z(n33161) );
  NAND U42124 ( .A(n33194), .B(n33195), .Z(n33193) );
  OR U42125 ( .A(n33196), .B(n33197), .Z(n33194) );
  NANDN U42126 ( .A(n33198), .B(n33196), .Z(n33192) );
  IV U42127 ( .A(n33197), .Z(n33198) );
  NAND U42128 ( .A(n33199), .B(n33200), .Z(n33158) );
  NAND U42129 ( .A(n33201), .B(n33202), .Z(n33200) );
  NANDN U42130 ( .A(n33203), .B(n33204), .Z(n33201) );
  NANDN U42131 ( .A(n33204), .B(n33203), .Z(n33199) );
  AND U42132 ( .A(n33205), .B(n33206), .Z(n33160) );
  NAND U42133 ( .A(n33207), .B(n33208), .Z(n33206) );
  OR U42134 ( .A(n33209), .B(n33210), .Z(n33207) );
  NANDN U42135 ( .A(n33211), .B(n33209), .Z(n33205) );
  XNOR U42136 ( .A(n33186), .B(n33212), .Z(N62452) );
  XOR U42137 ( .A(n33188), .B(n33189), .Z(n33212) );
  XNOR U42138 ( .A(n33202), .B(n33213), .Z(n33189) );
  XOR U42139 ( .A(n33203), .B(n33204), .Z(n33213) );
  XOR U42140 ( .A(n33209), .B(n33214), .Z(n33204) );
  XOR U42141 ( .A(n33208), .B(n33211), .Z(n33214) );
  IV U42142 ( .A(n33210), .Z(n33211) );
  NAND U42143 ( .A(n33215), .B(n33216), .Z(n33210) );
  OR U42144 ( .A(n33217), .B(n33218), .Z(n33216) );
  OR U42145 ( .A(n33219), .B(n33220), .Z(n33215) );
  NAND U42146 ( .A(n33221), .B(n33222), .Z(n33208) );
  OR U42147 ( .A(n33223), .B(n33224), .Z(n33222) );
  OR U42148 ( .A(n33225), .B(n33226), .Z(n33221) );
  NOR U42149 ( .A(n33227), .B(n33228), .Z(n33209) );
  ANDN U42150 ( .B(n33229), .A(n33230), .Z(n33203) );
  XNOR U42151 ( .A(n33196), .B(n33231), .Z(n33202) );
  XNOR U42152 ( .A(n33195), .B(n33197), .Z(n33231) );
  NAND U42153 ( .A(n33232), .B(n33233), .Z(n33197) );
  OR U42154 ( .A(n33234), .B(n33235), .Z(n33233) );
  OR U42155 ( .A(n33236), .B(n33237), .Z(n33232) );
  NAND U42156 ( .A(n33238), .B(n33239), .Z(n33195) );
  OR U42157 ( .A(n33240), .B(n33241), .Z(n33239) );
  OR U42158 ( .A(n33242), .B(n33243), .Z(n33238) );
  ANDN U42159 ( .B(n33244), .A(n33245), .Z(n33196) );
  IV U42160 ( .A(n33246), .Z(n33244) );
  ANDN U42161 ( .B(n33247), .A(n33248), .Z(n33188) );
  XOR U42162 ( .A(n33174), .B(n33249), .Z(n33186) );
  XOR U42163 ( .A(n33175), .B(n33176), .Z(n33249) );
  XOR U42164 ( .A(n33181), .B(n33250), .Z(n33176) );
  XOR U42165 ( .A(n33180), .B(n33183), .Z(n33250) );
  IV U42166 ( .A(n33182), .Z(n33183) );
  NAND U42167 ( .A(n33251), .B(n33252), .Z(n33182) );
  OR U42168 ( .A(n33253), .B(n33254), .Z(n33252) );
  OR U42169 ( .A(n33255), .B(n33256), .Z(n33251) );
  NAND U42170 ( .A(n33257), .B(n33258), .Z(n33180) );
  OR U42171 ( .A(n33259), .B(n33260), .Z(n33258) );
  OR U42172 ( .A(n33261), .B(n33262), .Z(n33257) );
  NOR U42173 ( .A(n33263), .B(n33264), .Z(n33181) );
  ANDN U42174 ( .B(n33265), .A(n33266), .Z(n33175) );
  IV U42175 ( .A(n33267), .Z(n33265) );
  XNOR U42176 ( .A(n33168), .B(n33268), .Z(n33174) );
  XNOR U42177 ( .A(n33167), .B(n33169), .Z(n33268) );
  NAND U42178 ( .A(n33269), .B(n33270), .Z(n33169) );
  OR U42179 ( .A(n33271), .B(n33272), .Z(n33270) );
  OR U42180 ( .A(n33273), .B(n33274), .Z(n33269) );
  NAND U42181 ( .A(n33275), .B(n33276), .Z(n33167) );
  OR U42182 ( .A(n33277), .B(n33278), .Z(n33276) );
  OR U42183 ( .A(n33279), .B(n33280), .Z(n33275) );
  ANDN U42184 ( .B(n33281), .A(n33282), .Z(n33168) );
  IV U42185 ( .A(n33283), .Z(n33281) );
  XNOR U42186 ( .A(n33248), .B(n33247), .Z(N62451) );
  XOR U42187 ( .A(n33267), .B(n33266), .Z(n33247) );
  XNOR U42188 ( .A(n33282), .B(n33283), .Z(n33266) );
  XNOR U42189 ( .A(n33277), .B(n33278), .Z(n33283) );
  XNOR U42190 ( .A(n33279), .B(n33280), .Z(n33278) );
  XNOR U42191 ( .A(y[3445]), .B(x[3445]), .Z(n33280) );
  XNOR U42192 ( .A(y[3446]), .B(x[3446]), .Z(n33279) );
  XNOR U42193 ( .A(y[3444]), .B(x[3444]), .Z(n33277) );
  XNOR U42194 ( .A(n33271), .B(n33272), .Z(n33282) );
  XNOR U42195 ( .A(y[3441]), .B(x[3441]), .Z(n33272) );
  XNOR U42196 ( .A(n33273), .B(n33274), .Z(n33271) );
  XNOR U42197 ( .A(y[3442]), .B(x[3442]), .Z(n33274) );
  XNOR U42198 ( .A(y[3443]), .B(x[3443]), .Z(n33273) );
  XNOR U42199 ( .A(n33264), .B(n33263), .Z(n33267) );
  XNOR U42200 ( .A(n33259), .B(n33260), .Z(n33263) );
  XNOR U42201 ( .A(y[3438]), .B(x[3438]), .Z(n33260) );
  XNOR U42202 ( .A(n33261), .B(n33262), .Z(n33259) );
  XNOR U42203 ( .A(y[3439]), .B(x[3439]), .Z(n33262) );
  XNOR U42204 ( .A(y[3440]), .B(x[3440]), .Z(n33261) );
  XNOR U42205 ( .A(n33253), .B(n33254), .Z(n33264) );
  XNOR U42206 ( .A(y[3435]), .B(x[3435]), .Z(n33254) );
  XNOR U42207 ( .A(n33255), .B(n33256), .Z(n33253) );
  XNOR U42208 ( .A(y[3436]), .B(x[3436]), .Z(n33256) );
  XNOR U42209 ( .A(y[3437]), .B(x[3437]), .Z(n33255) );
  XOR U42210 ( .A(n33229), .B(n33230), .Z(n33248) );
  XNOR U42211 ( .A(n33245), .B(n33246), .Z(n33230) );
  XNOR U42212 ( .A(n33240), .B(n33241), .Z(n33246) );
  XNOR U42213 ( .A(n33242), .B(n33243), .Z(n33241) );
  XNOR U42214 ( .A(y[3433]), .B(x[3433]), .Z(n33243) );
  XNOR U42215 ( .A(y[3434]), .B(x[3434]), .Z(n33242) );
  XNOR U42216 ( .A(y[3432]), .B(x[3432]), .Z(n33240) );
  XNOR U42217 ( .A(n33234), .B(n33235), .Z(n33245) );
  XNOR U42218 ( .A(y[3429]), .B(x[3429]), .Z(n33235) );
  XNOR U42219 ( .A(n33236), .B(n33237), .Z(n33234) );
  XNOR U42220 ( .A(y[3430]), .B(x[3430]), .Z(n33237) );
  XNOR U42221 ( .A(y[3431]), .B(x[3431]), .Z(n33236) );
  XOR U42222 ( .A(n33228), .B(n33227), .Z(n33229) );
  XNOR U42223 ( .A(n33223), .B(n33224), .Z(n33227) );
  XNOR U42224 ( .A(y[3426]), .B(x[3426]), .Z(n33224) );
  XNOR U42225 ( .A(n33225), .B(n33226), .Z(n33223) );
  XNOR U42226 ( .A(y[3427]), .B(x[3427]), .Z(n33226) );
  XNOR U42227 ( .A(y[3428]), .B(x[3428]), .Z(n33225) );
  XNOR U42228 ( .A(n33217), .B(n33218), .Z(n33228) );
  XNOR U42229 ( .A(y[3423]), .B(x[3423]), .Z(n33218) );
  XNOR U42230 ( .A(n33219), .B(n33220), .Z(n33217) );
  XNOR U42231 ( .A(y[3424]), .B(x[3424]), .Z(n33220) );
  XNOR U42232 ( .A(y[3425]), .B(x[3425]), .Z(n33219) );
  NAND U42233 ( .A(n33284), .B(n33285), .Z(N62442) );
  NANDN U42234 ( .A(n33286), .B(n33287), .Z(n33285) );
  OR U42235 ( .A(n33288), .B(n33289), .Z(n33287) );
  NAND U42236 ( .A(n33288), .B(n33289), .Z(n33284) );
  XOR U42237 ( .A(n33288), .B(n33290), .Z(N62441) );
  XNOR U42238 ( .A(n33286), .B(n33289), .Z(n33290) );
  AND U42239 ( .A(n33291), .B(n33292), .Z(n33289) );
  NANDN U42240 ( .A(n33293), .B(n33294), .Z(n33292) );
  NANDN U42241 ( .A(n33295), .B(n33296), .Z(n33294) );
  NANDN U42242 ( .A(n33296), .B(n33295), .Z(n33291) );
  NAND U42243 ( .A(n33297), .B(n33298), .Z(n33286) );
  NANDN U42244 ( .A(n33299), .B(n33300), .Z(n33298) );
  OR U42245 ( .A(n33301), .B(n33302), .Z(n33300) );
  NAND U42246 ( .A(n33302), .B(n33301), .Z(n33297) );
  AND U42247 ( .A(n33303), .B(n33304), .Z(n33288) );
  NANDN U42248 ( .A(n33305), .B(n33306), .Z(n33304) );
  NANDN U42249 ( .A(n33307), .B(n33308), .Z(n33306) );
  NANDN U42250 ( .A(n33308), .B(n33307), .Z(n33303) );
  XOR U42251 ( .A(n33302), .B(n33309), .Z(N62440) );
  XOR U42252 ( .A(n33299), .B(n33301), .Z(n33309) );
  XNOR U42253 ( .A(n33295), .B(n33310), .Z(n33301) );
  XNOR U42254 ( .A(n33293), .B(n33296), .Z(n33310) );
  NAND U42255 ( .A(n33311), .B(n33312), .Z(n33296) );
  NAND U42256 ( .A(n33313), .B(n33314), .Z(n33312) );
  OR U42257 ( .A(n33315), .B(n33316), .Z(n33313) );
  NANDN U42258 ( .A(n33317), .B(n33315), .Z(n33311) );
  IV U42259 ( .A(n33316), .Z(n33317) );
  NAND U42260 ( .A(n33318), .B(n33319), .Z(n33293) );
  NAND U42261 ( .A(n33320), .B(n33321), .Z(n33319) );
  NANDN U42262 ( .A(n33322), .B(n33323), .Z(n33320) );
  NANDN U42263 ( .A(n33323), .B(n33322), .Z(n33318) );
  AND U42264 ( .A(n33324), .B(n33325), .Z(n33295) );
  NAND U42265 ( .A(n33326), .B(n33327), .Z(n33325) );
  OR U42266 ( .A(n33328), .B(n33329), .Z(n33326) );
  NANDN U42267 ( .A(n33330), .B(n33328), .Z(n33324) );
  NAND U42268 ( .A(n33331), .B(n33332), .Z(n33299) );
  NANDN U42269 ( .A(n33333), .B(n33334), .Z(n33332) );
  OR U42270 ( .A(n33335), .B(n33336), .Z(n33334) );
  NANDN U42271 ( .A(n33337), .B(n33335), .Z(n33331) );
  IV U42272 ( .A(n33336), .Z(n33337) );
  XNOR U42273 ( .A(n33307), .B(n33338), .Z(n33302) );
  XNOR U42274 ( .A(n33305), .B(n33308), .Z(n33338) );
  NAND U42275 ( .A(n33339), .B(n33340), .Z(n33308) );
  NAND U42276 ( .A(n33341), .B(n33342), .Z(n33340) );
  OR U42277 ( .A(n33343), .B(n33344), .Z(n33341) );
  NANDN U42278 ( .A(n33345), .B(n33343), .Z(n33339) );
  IV U42279 ( .A(n33344), .Z(n33345) );
  NAND U42280 ( .A(n33346), .B(n33347), .Z(n33305) );
  NAND U42281 ( .A(n33348), .B(n33349), .Z(n33347) );
  NANDN U42282 ( .A(n33350), .B(n33351), .Z(n33348) );
  NANDN U42283 ( .A(n33351), .B(n33350), .Z(n33346) );
  AND U42284 ( .A(n33352), .B(n33353), .Z(n33307) );
  NAND U42285 ( .A(n33354), .B(n33355), .Z(n33353) );
  OR U42286 ( .A(n33356), .B(n33357), .Z(n33354) );
  NANDN U42287 ( .A(n33358), .B(n33356), .Z(n33352) );
  XNOR U42288 ( .A(n33333), .B(n33359), .Z(N62439) );
  XOR U42289 ( .A(n33335), .B(n33336), .Z(n33359) );
  XNOR U42290 ( .A(n33349), .B(n33360), .Z(n33336) );
  XOR U42291 ( .A(n33350), .B(n33351), .Z(n33360) );
  XOR U42292 ( .A(n33356), .B(n33361), .Z(n33351) );
  XOR U42293 ( .A(n33355), .B(n33358), .Z(n33361) );
  IV U42294 ( .A(n33357), .Z(n33358) );
  NAND U42295 ( .A(n33362), .B(n33363), .Z(n33357) );
  OR U42296 ( .A(n33364), .B(n33365), .Z(n33363) );
  OR U42297 ( .A(n33366), .B(n33367), .Z(n33362) );
  NAND U42298 ( .A(n33368), .B(n33369), .Z(n33355) );
  OR U42299 ( .A(n33370), .B(n33371), .Z(n33369) );
  OR U42300 ( .A(n33372), .B(n33373), .Z(n33368) );
  NOR U42301 ( .A(n33374), .B(n33375), .Z(n33356) );
  ANDN U42302 ( .B(n33376), .A(n33377), .Z(n33350) );
  XNOR U42303 ( .A(n33343), .B(n33378), .Z(n33349) );
  XNOR U42304 ( .A(n33342), .B(n33344), .Z(n33378) );
  NAND U42305 ( .A(n33379), .B(n33380), .Z(n33344) );
  OR U42306 ( .A(n33381), .B(n33382), .Z(n33380) );
  OR U42307 ( .A(n33383), .B(n33384), .Z(n33379) );
  NAND U42308 ( .A(n33385), .B(n33386), .Z(n33342) );
  OR U42309 ( .A(n33387), .B(n33388), .Z(n33386) );
  OR U42310 ( .A(n33389), .B(n33390), .Z(n33385) );
  ANDN U42311 ( .B(n33391), .A(n33392), .Z(n33343) );
  IV U42312 ( .A(n33393), .Z(n33391) );
  ANDN U42313 ( .B(n33394), .A(n33395), .Z(n33335) );
  XOR U42314 ( .A(n33321), .B(n33396), .Z(n33333) );
  XOR U42315 ( .A(n33322), .B(n33323), .Z(n33396) );
  XOR U42316 ( .A(n33328), .B(n33397), .Z(n33323) );
  XOR U42317 ( .A(n33327), .B(n33330), .Z(n33397) );
  IV U42318 ( .A(n33329), .Z(n33330) );
  NAND U42319 ( .A(n33398), .B(n33399), .Z(n33329) );
  OR U42320 ( .A(n33400), .B(n33401), .Z(n33399) );
  OR U42321 ( .A(n33402), .B(n33403), .Z(n33398) );
  NAND U42322 ( .A(n33404), .B(n33405), .Z(n33327) );
  OR U42323 ( .A(n33406), .B(n33407), .Z(n33405) );
  OR U42324 ( .A(n33408), .B(n33409), .Z(n33404) );
  NOR U42325 ( .A(n33410), .B(n33411), .Z(n33328) );
  ANDN U42326 ( .B(n33412), .A(n33413), .Z(n33322) );
  IV U42327 ( .A(n33414), .Z(n33412) );
  XNOR U42328 ( .A(n33315), .B(n33415), .Z(n33321) );
  XNOR U42329 ( .A(n33314), .B(n33316), .Z(n33415) );
  NAND U42330 ( .A(n33416), .B(n33417), .Z(n33316) );
  OR U42331 ( .A(n33418), .B(n33419), .Z(n33417) );
  OR U42332 ( .A(n33420), .B(n33421), .Z(n33416) );
  NAND U42333 ( .A(n33422), .B(n33423), .Z(n33314) );
  OR U42334 ( .A(n33424), .B(n33425), .Z(n33423) );
  OR U42335 ( .A(n33426), .B(n33427), .Z(n33422) );
  ANDN U42336 ( .B(n33428), .A(n33429), .Z(n33315) );
  IV U42337 ( .A(n33430), .Z(n33428) );
  XNOR U42338 ( .A(n33395), .B(n33394), .Z(N62438) );
  XOR U42339 ( .A(n33414), .B(n33413), .Z(n33394) );
  XNOR U42340 ( .A(n33429), .B(n33430), .Z(n33413) );
  XNOR U42341 ( .A(n33424), .B(n33425), .Z(n33430) );
  XNOR U42342 ( .A(n33426), .B(n33427), .Z(n33425) );
  XNOR U42343 ( .A(y[3421]), .B(x[3421]), .Z(n33427) );
  XNOR U42344 ( .A(y[3422]), .B(x[3422]), .Z(n33426) );
  XNOR U42345 ( .A(y[3420]), .B(x[3420]), .Z(n33424) );
  XNOR U42346 ( .A(n33418), .B(n33419), .Z(n33429) );
  XNOR U42347 ( .A(y[3417]), .B(x[3417]), .Z(n33419) );
  XNOR U42348 ( .A(n33420), .B(n33421), .Z(n33418) );
  XNOR U42349 ( .A(y[3418]), .B(x[3418]), .Z(n33421) );
  XNOR U42350 ( .A(y[3419]), .B(x[3419]), .Z(n33420) );
  XNOR U42351 ( .A(n33411), .B(n33410), .Z(n33414) );
  XNOR U42352 ( .A(n33406), .B(n33407), .Z(n33410) );
  XNOR U42353 ( .A(y[3414]), .B(x[3414]), .Z(n33407) );
  XNOR U42354 ( .A(n33408), .B(n33409), .Z(n33406) );
  XNOR U42355 ( .A(y[3415]), .B(x[3415]), .Z(n33409) );
  XNOR U42356 ( .A(y[3416]), .B(x[3416]), .Z(n33408) );
  XNOR U42357 ( .A(n33400), .B(n33401), .Z(n33411) );
  XNOR U42358 ( .A(y[3411]), .B(x[3411]), .Z(n33401) );
  XNOR U42359 ( .A(n33402), .B(n33403), .Z(n33400) );
  XNOR U42360 ( .A(y[3412]), .B(x[3412]), .Z(n33403) );
  XNOR U42361 ( .A(y[3413]), .B(x[3413]), .Z(n33402) );
  XOR U42362 ( .A(n33376), .B(n33377), .Z(n33395) );
  XNOR U42363 ( .A(n33392), .B(n33393), .Z(n33377) );
  XNOR U42364 ( .A(n33387), .B(n33388), .Z(n33393) );
  XNOR U42365 ( .A(n33389), .B(n33390), .Z(n33388) );
  XNOR U42366 ( .A(y[3409]), .B(x[3409]), .Z(n33390) );
  XNOR U42367 ( .A(y[3410]), .B(x[3410]), .Z(n33389) );
  XNOR U42368 ( .A(y[3408]), .B(x[3408]), .Z(n33387) );
  XNOR U42369 ( .A(n33381), .B(n33382), .Z(n33392) );
  XNOR U42370 ( .A(y[3405]), .B(x[3405]), .Z(n33382) );
  XNOR U42371 ( .A(n33383), .B(n33384), .Z(n33381) );
  XNOR U42372 ( .A(y[3406]), .B(x[3406]), .Z(n33384) );
  XNOR U42373 ( .A(y[3407]), .B(x[3407]), .Z(n33383) );
  XOR U42374 ( .A(n33375), .B(n33374), .Z(n33376) );
  XNOR U42375 ( .A(n33370), .B(n33371), .Z(n33374) );
  XNOR U42376 ( .A(y[3402]), .B(x[3402]), .Z(n33371) );
  XNOR U42377 ( .A(n33372), .B(n33373), .Z(n33370) );
  XNOR U42378 ( .A(y[3403]), .B(x[3403]), .Z(n33373) );
  XNOR U42379 ( .A(y[3404]), .B(x[3404]), .Z(n33372) );
  XNOR U42380 ( .A(n33364), .B(n33365), .Z(n33375) );
  XNOR U42381 ( .A(y[3399]), .B(x[3399]), .Z(n33365) );
  XNOR U42382 ( .A(n33366), .B(n33367), .Z(n33364) );
  XNOR U42383 ( .A(y[3400]), .B(x[3400]), .Z(n33367) );
  XNOR U42384 ( .A(y[3401]), .B(x[3401]), .Z(n33366) );
  NAND U42385 ( .A(n33431), .B(n33432), .Z(N62429) );
  NANDN U42386 ( .A(n33433), .B(n33434), .Z(n33432) );
  OR U42387 ( .A(n33435), .B(n33436), .Z(n33434) );
  NAND U42388 ( .A(n33435), .B(n33436), .Z(n33431) );
  XOR U42389 ( .A(n33435), .B(n33437), .Z(N62428) );
  XNOR U42390 ( .A(n33433), .B(n33436), .Z(n33437) );
  AND U42391 ( .A(n33438), .B(n33439), .Z(n33436) );
  NANDN U42392 ( .A(n33440), .B(n33441), .Z(n33439) );
  NANDN U42393 ( .A(n33442), .B(n33443), .Z(n33441) );
  NANDN U42394 ( .A(n33443), .B(n33442), .Z(n33438) );
  NAND U42395 ( .A(n33444), .B(n33445), .Z(n33433) );
  NANDN U42396 ( .A(n33446), .B(n33447), .Z(n33445) );
  OR U42397 ( .A(n33448), .B(n33449), .Z(n33447) );
  NAND U42398 ( .A(n33449), .B(n33448), .Z(n33444) );
  AND U42399 ( .A(n33450), .B(n33451), .Z(n33435) );
  NANDN U42400 ( .A(n33452), .B(n33453), .Z(n33451) );
  NANDN U42401 ( .A(n33454), .B(n33455), .Z(n33453) );
  NANDN U42402 ( .A(n33455), .B(n33454), .Z(n33450) );
  XOR U42403 ( .A(n33449), .B(n33456), .Z(N62427) );
  XOR U42404 ( .A(n33446), .B(n33448), .Z(n33456) );
  XNOR U42405 ( .A(n33442), .B(n33457), .Z(n33448) );
  XNOR U42406 ( .A(n33440), .B(n33443), .Z(n33457) );
  NAND U42407 ( .A(n33458), .B(n33459), .Z(n33443) );
  NAND U42408 ( .A(n33460), .B(n33461), .Z(n33459) );
  OR U42409 ( .A(n33462), .B(n33463), .Z(n33460) );
  NANDN U42410 ( .A(n33464), .B(n33462), .Z(n33458) );
  IV U42411 ( .A(n33463), .Z(n33464) );
  NAND U42412 ( .A(n33465), .B(n33466), .Z(n33440) );
  NAND U42413 ( .A(n33467), .B(n33468), .Z(n33466) );
  NANDN U42414 ( .A(n33469), .B(n33470), .Z(n33467) );
  NANDN U42415 ( .A(n33470), .B(n33469), .Z(n33465) );
  AND U42416 ( .A(n33471), .B(n33472), .Z(n33442) );
  NAND U42417 ( .A(n33473), .B(n33474), .Z(n33472) );
  OR U42418 ( .A(n33475), .B(n33476), .Z(n33473) );
  NANDN U42419 ( .A(n33477), .B(n33475), .Z(n33471) );
  NAND U42420 ( .A(n33478), .B(n33479), .Z(n33446) );
  NANDN U42421 ( .A(n33480), .B(n33481), .Z(n33479) );
  OR U42422 ( .A(n33482), .B(n33483), .Z(n33481) );
  NANDN U42423 ( .A(n33484), .B(n33482), .Z(n33478) );
  IV U42424 ( .A(n33483), .Z(n33484) );
  XNOR U42425 ( .A(n33454), .B(n33485), .Z(n33449) );
  XNOR U42426 ( .A(n33452), .B(n33455), .Z(n33485) );
  NAND U42427 ( .A(n33486), .B(n33487), .Z(n33455) );
  NAND U42428 ( .A(n33488), .B(n33489), .Z(n33487) );
  OR U42429 ( .A(n33490), .B(n33491), .Z(n33488) );
  NANDN U42430 ( .A(n33492), .B(n33490), .Z(n33486) );
  IV U42431 ( .A(n33491), .Z(n33492) );
  NAND U42432 ( .A(n33493), .B(n33494), .Z(n33452) );
  NAND U42433 ( .A(n33495), .B(n33496), .Z(n33494) );
  NANDN U42434 ( .A(n33497), .B(n33498), .Z(n33495) );
  NANDN U42435 ( .A(n33498), .B(n33497), .Z(n33493) );
  AND U42436 ( .A(n33499), .B(n33500), .Z(n33454) );
  NAND U42437 ( .A(n33501), .B(n33502), .Z(n33500) );
  OR U42438 ( .A(n33503), .B(n33504), .Z(n33501) );
  NANDN U42439 ( .A(n33505), .B(n33503), .Z(n33499) );
  XNOR U42440 ( .A(n33480), .B(n33506), .Z(N62426) );
  XOR U42441 ( .A(n33482), .B(n33483), .Z(n33506) );
  XNOR U42442 ( .A(n33496), .B(n33507), .Z(n33483) );
  XOR U42443 ( .A(n33497), .B(n33498), .Z(n33507) );
  XOR U42444 ( .A(n33503), .B(n33508), .Z(n33498) );
  XOR U42445 ( .A(n33502), .B(n33505), .Z(n33508) );
  IV U42446 ( .A(n33504), .Z(n33505) );
  NAND U42447 ( .A(n33509), .B(n33510), .Z(n33504) );
  OR U42448 ( .A(n33511), .B(n33512), .Z(n33510) );
  OR U42449 ( .A(n33513), .B(n33514), .Z(n33509) );
  NAND U42450 ( .A(n33515), .B(n33516), .Z(n33502) );
  OR U42451 ( .A(n33517), .B(n33518), .Z(n33516) );
  OR U42452 ( .A(n33519), .B(n33520), .Z(n33515) );
  NOR U42453 ( .A(n33521), .B(n33522), .Z(n33503) );
  ANDN U42454 ( .B(n33523), .A(n33524), .Z(n33497) );
  XNOR U42455 ( .A(n33490), .B(n33525), .Z(n33496) );
  XNOR U42456 ( .A(n33489), .B(n33491), .Z(n33525) );
  NAND U42457 ( .A(n33526), .B(n33527), .Z(n33491) );
  OR U42458 ( .A(n33528), .B(n33529), .Z(n33527) );
  OR U42459 ( .A(n33530), .B(n33531), .Z(n33526) );
  NAND U42460 ( .A(n33532), .B(n33533), .Z(n33489) );
  OR U42461 ( .A(n33534), .B(n33535), .Z(n33533) );
  OR U42462 ( .A(n33536), .B(n33537), .Z(n33532) );
  ANDN U42463 ( .B(n33538), .A(n33539), .Z(n33490) );
  IV U42464 ( .A(n33540), .Z(n33538) );
  ANDN U42465 ( .B(n33541), .A(n33542), .Z(n33482) );
  XOR U42466 ( .A(n33468), .B(n33543), .Z(n33480) );
  XOR U42467 ( .A(n33469), .B(n33470), .Z(n33543) );
  XOR U42468 ( .A(n33475), .B(n33544), .Z(n33470) );
  XOR U42469 ( .A(n33474), .B(n33477), .Z(n33544) );
  IV U42470 ( .A(n33476), .Z(n33477) );
  NAND U42471 ( .A(n33545), .B(n33546), .Z(n33476) );
  OR U42472 ( .A(n33547), .B(n33548), .Z(n33546) );
  OR U42473 ( .A(n33549), .B(n33550), .Z(n33545) );
  NAND U42474 ( .A(n33551), .B(n33552), .Z(n33474) );
  OR U42475 ( .A(n33553), .B(n33554), .Z(n33552) );
  OR U42476 ( .A(n33555), .B(n33556), .Z(n33551) );
  NOR U42477 ( .A(n33557), .B(n33558), .Z(n33475) );
  ANDN U42478 ( .B(n33559), .A(n33560), .Z(n33469) );
  IV U42479 ( .A(n33561), .Z(n33559) );
  XNOR U42480 ( .A(n33462), .B(n33562), .Z(n33468) );
  XNOR U42481 ( .A(n33461), .B(n33463), .Z(n33562) );
  NAND U42482 ( .A(n33563), .B(n33564), .Z(n33463) );
  OR U42483 ( .A(n33565), .B(n33566), .Z(n33564) );
  OR U42484 ( .A(n33567), .B(n33568), .Z(n33563) );
  NAND U42485 ( .A(n33569), .B(n33570), .Z(n33461) );
  OR U42486 ( .A(n33571), .B(n33572), .Z(n33570) );
  OR U42487 ( .A(n33573), .B(n33574), .Z(n33569) );
  ANDN U42488 ( .B(n33575), .A(n33576), .Z(n33462) );
  IV U42489 ( .A(n33577), .Z(n33575) );
  XNOR U42490 ( .A(n33542), .B(n33541), .Z(N62425) );
  XOR U42491 ( .A(n33561), .B(n33560), .Z(n33541) );
  XNOR U42492 ( .A(n33576), .B(n33577), .Z(n33560) );
  XNOR U42493 ( .A(n33571), .B(n33572), .Z(n33577) );
  XNOR U42494 ( .A(n33573), .B(n33574), .Z(n33572) );
  XNOR U42495 ( .A(y[3397]), .B(x[3397]), .Z(n33574) );
  XNOR U42496 ( .A(y[3398]), .B(x[3398]), .Z(n33573) );
  XNOR U42497 ( .A(y[3396]), .B(x[3396]), .Z(n33571) );
  XNOR U42498 ( .A(n33565), .B(n33566), .Z(n33576) );
  XNOR U42499 ( .A(y[3393]), .B(x[3393]), .Z(n33566) );
  XNOR U42500 ( .A(n33567), .B(n33568), .Z(n33565) );
  XNOR U42501 ( .A(y[3394]), .B(x[3394]), .Z(n33568) );
  XNOR U42502 ( .A(y[3395]), .B(x[3395]), .Z(n33567) );
  XNOR U42503 ( .A(n33558), .B(n33557), .Z(n33561) );
  XNOR U42504 ( .A(n33553), .B(n33554), .Z(n33557) );
  XNOR U42505 ( .A(y[3390]), .B(x[3390]), .Z(n33554) );
  XNOR U42506 ( .A(n33555), .B(n33556), .Z(n33553) );
  XNOR U42507 ( .A(y[3391]), .B(x[3391]), .Z(n33556) );
  XNOR U42508 ( .A(y[3392]), .B(x[3392]), .Z(n33555) );
  XNOR U42509 ( .A(n33547), .B(n33548), .Z(n33558) );
  XNOR U42510 ( .A(y[3387]), .B(x[3387]), .Z(n33548) );
  XNOR U42511 ( .A(n33549), .B(n33550), .Z(n33547) );
  XNOR U42512 ( .A(y[3388]), .B(x[3388]), .Z(n33550) );
  XNOR U42513 ( .A(y[3389]), .B(x[3389]), .Z(n33549) );
  XOR U42514 ( .A(n33523), .B(n33524), .Z(n33542) );
  XNOR U42515 ( .A(n33539), .B(n33540), .Z(n33524) );
  XNOR U42516 ( .A(n33534), .B(n33535), .Z(n33540) );
  XNOR U42517 ( .A(n33536), .B(n33537), .Z(n33535) );
  XNOR U42518 ( .A(y[3385]), .B(x[3385]), .Z(n33537) );
  XNOR U42519 ( .A(y[3386]), .B(x[3386]), .Z(n33536) );
  XNOR U42520 ( .A(y[3384]), .B(x[3384]), .Z(n33534) );
  XNOR U42521 ( .A(n33528), .B(n33529), .Z(n33539) );
  XNOR U42522 ( .A(y[3381]), .B(x[3381]), .Z(n33529) );
  XNOR U42523 ( .A(n33530), .B(n33531), .Z(n33528) );
  XNOR U42524 ( .A(y[3382]), .B(x[3382]), .Z(n33531) );
  XNOR U42525 ( .A(y[3383]), .B(x[3383]), .Z(n33530) );
  XOR U42526 ( .A(n33522), .B(n33521), .Z(n33523) );
  XNOR U42527 ( .A(n33517), .B(n33518), .Z(n33521) );
  XNOR U42528 ( .A(y[3378]), .B(x[3378]), .Z(n33518) );
  XNOR U42529 ( .A(n33519), .B(n33520), .Z(n33517) );
  XNOR U42530 ( .A(y[3379]), .B(x[3379]), .Z(n33520) );
  XNOR U42531 ( .A(y[3380]), .B(x[3380]), .Z(n33519) );
  XNOR U42532 ( .A(n33511), .B(n33512), .Z(n33522) );
  XNOR U42533 ( .A(y[3375]), .B(x[3375]), .Z(n33512) );
  XNOR U42534 ( .A(n33513), .B(n33514), .Z(n33511) );
  XNOR U42535 ( .A(y[3376]), .B(x[3376]), .Z(n33514) );
  XNOR U42536 ( .A(y[3377]), .B(x[3377]), .Z(n33513) );
  NAND U42537 ( .A(n33578), .B(n33579), .Z(N62416) );
  NANDN U42538 ( .A(n33580), .B(n33581), .Z(n33579) );
  OR U42539 ( .A(n33582), .B(n33583), .Z(n33581) );
  NAND U42540 ( .A(n33582), .B(n33583), .Z(n33578) );
  XOR U42541 ( .A(n33582), .B(n33584), .Z(N62415) );
  XNOR U42542 ( .A(n33580), .B(n33583), .Z(n33584) );
  AND U42543 ( .A(n33585), .B(n33586), .Z(n33583) );
  NANDN U42544 ( .A(n33587), .B(n33588), .Z(n33586) );
  NANDN U42545 ( .A(n33589), .B(n33590), .Z(n33588) );
  NANDN U42546 ( .A(n33590), .B(n33589), .Z(n33585) );
  NAND U42547 ( .A(n33591), .B(n33592), .Z(n33580) );
  NANDN U42548 ( .A(n33593), .B(n33594), .Z(n33592) );
  OR U42549 ( .A(n33595), .B(n33596), .Z(n33594) );
  NAND U42550 ( .A(n33596), .B(n33595), .Z(n33591) );
  AND U42551 ( .A(n33597), .B(n33598), .Z(n33582) );
  NANDN U42552 ( .A(n33599), .B(n33600), .Z(n33598) );
  NANDN U42553 ( .A(n33601), .B(n33602), .Z(n33600) );
  NANDN U42554 ( .A(n33602), .B(n33601), .Z(n33597) );
  XOR U42555 ( .A(n33596), .B(n33603), .Z(N62414) );
  XOR U42556 ( .A(n33593), .B(n33595), .Z(n33603) );
  XNOR U42557 ( .A(n33589), .B(n33604), .Z(n33595) );
  XNOR U42558 ( .A(n33587), .B(n33590), .Z(n33604) );
  NAND U42559 ( .A(n33605), .B(n33606), .Z(n33590) );
  NAND U42560 ( .A(n33607), .B(n33608), .Z(n33606) );
  OR U42561 ( .A(n33609), .B(n33610), .Z(n33607) );
  NANDN U42562 ( .A(n33611), .B(n33609), .Z(n33605) );
  IV U42563 ( .A(n33610), .Z(n33611) );
  NAND U42564 ( .A(n33612), .B(n33613), .Z(n33587) );
  NAND U42565 ( .A(n33614), .B(n33615), .Z(n33613) );
  NANDN U42566 ( .A(n33616), .B(n33617), .Z(n33614) );
  NANDN U42567 ( .A(n33617), .B(n33616), .Z(n33612) );
  AND U42568 ( .A(n33618), .B(n33619), .Z(n33589) );
  NAND U42569 ( .A(n33620), .B(n33621), .Z(n33619) );
  OR U42570 ( .A(n33622), .B(n33623), .Z(n33620) );
  NANDN U42571 ( .A(n33624), .B(n33622), .Z(n33618) );
  NAND U42572 ( .A(n33625), .B(n33626), .Z(n33593) );
  NANDN U42573 ( .A(n33627), .B(n33628), .Z(n33626) );
  OR U42574 ( .A(n33629), .B(n33630), .Z(n33628) );
  NANDN U42575 ( .A(n33631), .B(n33629), .Z(n33625) );
  IV U42576 ( .A(n33630), .Z(n33631) );
  XNOR U42577 ( .A(n33601), .B(n33632), .Z(n33596) );
  XNOR U42578 ( .A(n33599), .B(n33602), .Z(n33632) );
  NAND U42579 ( .A(n33633), .B(n33634), .Z(n33602) );
  NAND U42580 ( .A(n33635), .B(n33636), .Z(n33634) );
  OR U42581 ( .A(n33637), .B(n33638), .Z(n33635) );
  NANDN U42582 ( .A(n33639), .B(n33637), .Z(n33633) );
  IV U42583 ( .A(n33638), .Z(n33639) );
  NAND U42584 ( .A(n33640), .B(n33641), .Z(n33599) );
  NAND U42585 ( .A(n33642), .B(n33643), .Z(n33641) );
  NANDN U42586 ( .A(n33644), .B(n33645), .Z(n33642) );
  NANDN U42587 ( .A(n33645), .B(n33644), .Z(n33640) );
  AND U42588 ( .A(n33646), .B(n33647), .Z(n33601) );
  NAND U42589 ( .A(n33648), .B(n33649), .Z(n33647) );
  OR U42590 ( .A(n33650), .B(n33651), .Z(n33648) );
  NANDN U42591 ( .A(n33652), .B(n33650), .Z(n33646) );
  XNOR U42592 ( .A(n33627), .B(n33653), .Z(N62413) );
  XOR U42593 ( .A(n33629), .B(n33630), .Z(n33653) );
  XNOR U42594 ( .A(n33643), .B(n33654), .Z(n33630) );
  XOR U42595 ( .A(n33644), .B(n33645), .Z(n33654) );
  XOR U42596 ( .A(n33650), .B(n33655), .Z(n33645) );
  XOR U42597 ( .A(n33649), .B(n33652), .Z(n33655) );
  IV U42598 ( .A(n33651), .Z(n33652) );
  NAND U42599 ( .A(n33656), .B(n33657), .Z(n33651) );
  OR U42600 ( .A(n33658), .B(n33659), .Z(n33657) );
  OR U42601 ( .A(n33660), .B(n33661), .Z(n33656) );
  NAND U42602 ( .A(n33662), .B(n33663), .Z(n33649) );
  OR U42603 ( .A(n33664), .B(n33665), .Z(n33663) );
  OR U42604 ( .A(n33666), .B(n33667), .Z(n33662) );
  NOR U42605 ( .A(n33668), .B(n33669), .Z(n33650) );
  ANDN U42606 ( .B(n33670), .A(n33671), .Z(n33644) );
  XNOR U42607 ( .A(n33637), .B(n33672), .Z(n33643) );
  XNOR U42608 ( .A(n33636), .B(n33638), .Z(n33672) );
  NAND U42609 ( .A(n33673), .B(n33674), .Z(n33638) );
  OR U42610 ( .A(n33675), .B(n33676), .Z(n33674) );
  OR U42611 ( .A(n33677), .B(n33678), .Z(n33673) );
  NAND U42612 ( .A(n33679), .B(n33680), .Z(n33636) );
  OR U42613 ( .A(n33681), .B(n33682), .Z(n33680) );
  OR U42614 ( .A(n33683), .B(n33684), .Z(n33679) );
  ANDN U42615 ( .B(n33685), .A(n33686), .Z(n33637) );
  IV U42616 ( .A(n33687), .Z(n33685) );
  ANDN U42617 ( .B(n33688), .A(n33689), .Z(n33629) );
  XOR U42618 ( .A(n33615), .B(n33690), .Z(n33627) );
  XOR U42619 ( .A(n33616), .B(n33617), .Z(n33690) );
  XOR U42620 ( .A(n33622), .B(n33691), .Z(n33617) );
  XOR U42621 ( .A(n33621), .B(n33624), .Z(n33691) );
  IV U42622 ( .A(n33623), .Z(n33624) );
  NAND U42623 ( .A(n33692), .B(n33693), .Z(n33623) );
  OR U42624 ( .A(n33694), .B(n33695), .Z(n33693) );
  OR U42625 ( .A(n33696), .B(n33697), .Z(n33692) );
  NAND U42626 ( .A(n33698), .B(n33699), .Z(n33621) );
  OR U42627 ( .A(n33700), .B(n33701), .Z(n33699) );
  OR U42628 ( .A(n33702), .B(n33703), .Z(n33698) );
  NOR U42629 ( .A(n33704), .B(n33705), .Z(n33622) );
  ANDN U42630 ( .B(n33706), .A(n33707), .Z(n33616) );
  IV U42631 ( .A(n33708), .Z(n33706) );
  XNOR U42632 ( .A(n33609), .B(n33709), .Z(n33615) );
  XNOR U42633 ( .A(n33608), .B(n33610), .Z(n33709) );
  NAND U42634 ( .A(n33710), .B(n33711), .Z(n33610) );
  OR U42635 ( .A(n33712), .B(n33713), .Z(n33711) );
  OR U42636 ( .A(n33714), .B(n33715), .Z(n33710) );
  NAND U42637 ( .A(n33716), .B(n33717), .Z(n33608) );
  OR U42638 ( .A(n33718), .B(n33719), .Z(n33717) );
  OR U42639 ( .A(n33720), .B(n33721), .Z(n33716) );
  ANDN U42640 ( .B(n33722), .A(n33723), .Z(n33609) );
  IV U42641 ( .A(n33724), .Z(n33722) );
  XNOR U42642 ( .A(n33689), .B(n33688), .Z(N62412) );
  XOR U42643 ( .A(n33708), .B(n33707), .Z(n33688) );
  XNOR U42644 ( .A(n33723), .B(n33724), .Z(n33707) );
  XNOR U42645 ( .A(n33718), .B(n33719), .Z(n33724) );
  XNOR U42646 ( .A(n33720), .B(n33721), .Z(n33719) );
  XNOR U42647 ( .A(y[3373]), .B(x[3373]), .Z(n33721) );
  XNOR U42648 ( .A(y[3374]), .B(x[3374]), .Z(n33720) );
  XNOR U42649 ( .A(y[3372]), .B(x[3372]), .Z(n33718) );
  XNOR U42650 ( .A(n33712), .B(n33713), .Z(n33723) );
  XNOR U42651 ( .A(y[3369]), .B(x[3369]), .Z(n33713) );
  XNOR U42652 ( .A(n33714), .B(n33715), .Z(n33712) );
  XNOR U42653 ( .A(y[3370]), .B(x[3370]), .Z(n33715) );
  XNOR U42654 ( .A(y[3371]), .B(x[3371]), .Z(n33714) );
  XNOR U42655 ( .A(n33705), .B(n33704), .Z(n33708) );
  XNOR U42656 ( .A(n33700), .B(n33701), .Z(n33704) );
  XNOR U42657 ( .A(y[3366]), .B(x[3366]), .Z(n33701) );
  XNOR U42658 ( .A(n33702), .B(n33703), .Z(n33700) );
  XNOR U42659 ( .A(y[3367]), .B(x[3367]), .Z(n33703) );
  XNOR U42660 ( .A(y[3368]), .B(x[3368]), .Z(n33702) );
  XNOR U42661 ( .A(n33694), .B(n33695), .Z(n33705) );
  XNOR U42662 ( .A(y[3363]), .B(x[3363]), .Z(n33695) );
  XNOR U42663 ( .A(n33696), .B(n33697), .Z(n33694) );
  XNOR U42664 ( .A(y[3364]), .B(x[3364]), .Z(n33697) );
  XNOR U42665 ( .A(y[3365]), .B(x[3365]), .Z(n33696) );
  XOR U42666 ( .A(n33670), .B(n33671), .Z(n33689) );
  XNOR U42667 ( .A(n33686), .B(n33687), .Z(n33671) );
  XNOR U42668 ( .A(n33681), .B(n33682), .Z(n33687) );
  XNOR U42669 ( .A(n33683), .B(n33684), .Z(n33682) );
  XNOR U42670 ( .A(y[3361]), .B(x[3361]), .Z(n33684) );
  XNOR U42671 ( .A(y[3362]), .B(x[3362]), .Z(n33683) );
  XNOR U42672 ( .A(y[3360]), .B(x[3360]), .Z(n33681) );
  XNOR U42673 ( .A(n33675), .B(n33676), .Z(n33686) );
  XNOR U42674 ( .A(y[3357]), .B(x[3357]), .Z(n33676) );
  XNOR U42675 ( .A(n33677), .B(n33678), .Z(n33675) );
  XNOR U42676 ( .A(y[3358]), .B(x[3358]), .Z(n33678) );
  XNOR U42677 ( .A(y[3359]), .B(x[3359]), .Z(n33677) );
  XOR U42678 ( .A(n33669), .B(n33668), .Z(n33670) );
  XNOR U42679 ( .A(n33664), .B(n33665), .Z(n33668) );
  XNOR U42680 ( .A(y[3354]), .B(x[3354]), .Z(n33665) );
  XNOR U42681 ( .A(n33666), .B(n33667), .Z(n33664) );
  XNOR U42682 ( .A(y[3355]), .B(x[3355]), .Z(n33667) );
  XNOR U42683 ( .A(y[3356]), .B(x[3356]), .Z(n33666) );
  XNOR U42684 ( .A(n33658), .B(n33659), .Z(n33669) );
  XNOR U42685 ( .A(y[3351]), .B(x[3351]), .Z(n33659) );
  XNOR U42686 ( .A(n33660), .B(n33661), .Z(n33658) );
  XNOR U42687 ( .A(y[3352]), .B(x[3352]), .Z(n33661) );
  XNOR U42688 ( .A(y[3353]), .B(x[3353]), .Z(n33660) );
  NAND U42689 ( .A(n33725), .B(n33726), .Z(N62403) );
  NANDN U42690 ( .A(n33727), .B(n33728), .Z(n33726) );
  OR U42691 ( .A(n33729), .B(n33730), .Z(n33728) );
  NAND U42692 ( .A(n33729), .B(n33730), .Z(n33725) );
  XOR U42693 ( .A(n33729), .B(n33731), .Z(N62402) );
  XNOR U42694 ( .A(n33727), .B(n33730), .Z(n33731) );
  AND U42695 ( .A(n33732), .B(n33733), .Z(n33730) );
  NANDN U42696 ( .A(n33734), .B(n33735), .Z(n33733) );
  NANDN U42697 ( .A(n33736), .B(n33737), .Z(n33735) );
  NANDN U42698 ( .A(n33737), .B(n33736), .Z(n33732) );
  NAND U42699 ( .A(n33738), .B(n33739), .Z(n33727) );
  NANDN U42700 ( .A(n33740), .B(n33741), .Z(n33739) );
  OR U42701 ( .A(n33742), .B(n33743), .Z(n33741) );
  NAND U42702 ( .A(n33743), .B(n33742), .Z(n33738) );
  AND U42703 ( .A(n33744), .B(n33745), .Z(n33729) );
  NANDN U42704 ( .A(n33746), .B(n33747), .Z(n33745) );
  NANDN U42705 ( .A(n33748), .B(n33749), .Z(n33747) );
  NANDN U42706 ( .A(n33749), .B(n33748), .Z(n33744) );
  XOR U42707 ( .A(n33743), .B(n33750), .Z(N62401) );
  XOR U42708 ( .A(n33740), .B(n33742), .Z(n33750) );
  XNOR U42709 ( .A(n33736), .B(n33751), .Z(n33742) );
  XNOR U42710 ( .A(n33734), .B(n33737), .Z(n33751) );
  NAND U42711 ( .A(n33752), .B(n33753), .Z(n33737) );
  NAND U42712 ( .A(n33754), .B(n33755), .Z(n33753) );
  OR U42713 ( .A(n33756), .B(n33757), .Z(n33754) );
  NANDN U42714 ( .A(n33758), .B(n33756), .Z(n33752) );
  IV U42715 ( .A(n33757), .Z(n33758) );
  NAND U42716 ( .A(n33759), .B(n33760), .Z(n33734) );
  NAND U42717 ( .A(n33761), .B(n33762), .Z(n33760) );
  NANDN U42718 ( .A(n33763), .B(n33764), .Z(n33761) );
  NANDN U42719 ( .A(n33764), .B(n33763), .Z(n33759) );
  AND U42720 ( .A(n33765), .B(n33766), .Z(n33736) );
  NAND U42721 ( .A(n33767), .B(n33768), .Z(n33766) );
  OR U42722 ( .A(n33769), .B(n33770), .Z(n33767) );
  NANDN U42723 ( .A(n33771), .B(n33769), .Z(n33765) );
  NAND U42724 ( .A(n33772), .B(n33773), .Z(n33740) );
  NANDN U42725 ( .A(n33774), .B(n33775), .Z(n33773) );
  OR U42726 ( .A(n33776), .B(n33777), .Z(n33775) );
  NANDN U42727 ( .A(n33778), .B(n33776), .Z(n33772) );
  IV U42728 ( .A(n33777), .Z(n33778) );
  XNOR U42729 ( .A(n33748), .B(n33779), .Z(n33743) );
  XNOR U42730 ( .A(n33746), .B(n33749), .Z(n33779) );
  NAND U42731 ( .A(n33780), .B(n33781), .Z(n33749) );
  NAND U42732 ( .A(n33782), .B(n33783), .Z(n33781) );
  OR U42733 ( .A(n33784), .B(n33785), .Z(n33782) );
  NANDN U42734 ( .A(n33786), .B(n33784), .Z(n33780) );
  IV U42735 ( .A(n33785), .Z(n33786) );
  NAND U42736 ( .A(n33787), .B(n33788), .Z(n33746) );
  NAND U42737 ( .A(n33789), .B(n33790), .Z(n33788) );
  NANDN U42738 ( .A(n33791), .B(n33792), .Z(n33789) );
  NANDN U42739 ( .A(n33792), .B(n33791), .Z(n33787) );
  AND U42740 ( .A(n33793), .B(n33794), .Z(n33748) );
  NAND U42741 ( .A(n33795), .B(n33796), .Z(n33794) );
  OR U42742 ( .A(n33797), .B(n33798), .Z(n33795) );
  NANDN U42743 ( .A(n33799), .B(n33797), .Z(n33793) );
  XNOR U42744 ( .A(n33774), .B(n33800), .Z(N62400) );
  XOR U42745 ( .A(n33776), .B(n33777), .Z(n33800) );
  XNOR U42746 ( .A(n33790), .B(n33801), .Z(n33777) );
  XOR U42747 ( .A(n33791), .B(n33792), .Z(n33801) );
  XOR U42748 ( .A(n33797), .B(n33802), .Z(n33792) );
  XOR U42749 ( .A(n33796), .B(n33799), .Z(n33802) );
  IV U42750 ( .A(n33798), .Z(n33799) );
  NAND U42751 ( .A(n33803), .B(n33804), .Z(n33798) );
  OR U42752 ( .A(n33805), .B(n33806), .Z(n33804) );
  OR U42753 ( .A(n33807), .B(n33808), .Z(n33803) );
  NAND U42754 ( .A(n33809), .B(n33810), .Z(n33796) );
  OR U42755 ( .A(n33811), .B(n33812), .Z(n33810) );
  OR U42756 ( .A(n33813), .B(n33814), .Z(n33809) );
  NOR U42757 ( .A(n33815), .B(n33816), .Z(n33797) );
  ANDN U42758 ( .B(n33817), .A(n33818), .Z(n33791) );
  XNOR U42759 ( .A(n33784), .B(n33819), .Z(n33790) );
  XNOR U42760 ( .A(n33783), .B(n33785), .Z(n33819) );
  NAND U42761 ( .A(n33820), .B(n33821), .Z(n33785) );
  OR U42762 ( .A(n33822), .B(n33823), .Z(n33821) );
  OR U42763 ( .A(n33824), .B(n33825), .Z(n33820) );
  NAND U42764 ( .A(n33826), .B(n33827), .Z(n33783) );
  OR U42765 ( .A(n33828), .B(n33829), .Z(n33827) );
  OR U42766 ( .A(n33830), .B(n33831), .Z(n33826) );
  ANDN U42767 ( .B(n33832), .A(n33833), .Z(n33784) );
  IV U42768 ( .A(n33834), .Z(n33832) );
  ANDN U42769 ( .B(n33835), .A(n33836), .Z(n33776) );
  XOR U42770 ( .A(n33762), .B(n33837), .Z(n33774) );
  XOR U42771 ( .A(n33763), .B(n33764), .Z(n33837) );
  XOR U42772 ( .A(n33769), .B(n33838), .Z(n33764) );
  XOR U42773 ( .A(n33768), .B(n33771), .Z(n33838) );
  IV U42774 ( .A(n33770), .Z(n33771) );
  NAND U42775 ( .A(n33839), .B(n33840), .Z(n33770) );
  OR U42776 ( .A(n33841), .B(n33842), .Z(n33840) );
  OR U42777 ( .A(n33843), .B(n33844), .Z(n33839) );
  NAND U42778 ( .A(n33845), .B(n33846), .Z(n33768) );
  OR U42779 ( .A(n33847), .B(n33848), .Z(n33846) );
  OR U42780 ( .A(n33849), .B(n33850), .Z(n33845) );
  NOR U42781 ( .A(n33851), .B(n33852), .Z(n33769) );
  ANDN U42782 ( .B(n33853), .A(n33854), .Z(n33763) );
  IV U42783 ( .A(n33855), .Z(n33853) );
  XNOR U42784 ( .A(n33756), .B(n33856), .Z(n33762) );
  XNOR U42785 ( .A(n33755), .B(n33757), .Z(n33856) );
  NAND U42786 ( .A(n33857), .B(n33858), .Z(n33757) );
  OR U42787 ( .A(n33859), .B(n33860), .Z(n33858) );
  OR U42788 ( .A(n33861), .B(n33862), .Z(n33857) );
  NAND U42789 ( .A(n33863), .B(n33864), .Z(n33755) );
  OR U42790 ( .A(n33865), .B(n33866), .Z(n33864) );
  OR U42791 ( .A(n33867), .B(n33868), .Z(n33863) );
  ANDN U42792 ( .B(n33869), .A(n33870), .Z(n33756) );
  IV U42793 ( .A(n33871), .Z(n33869) );
  XNOR U42794 ( .A(n33836), .B(n33835), .Z(N62399) );
  XOR U42795 ( .A(n33855), .B(n33854), .Z(n33835) );
  XNOR U42796 ( .A(n33870), .B(n33871), .Z(n33854) );
  XNOR U42797 ( .A(n33865), .B(n33866), .Z(n33871) );
  XNOR U42798 ( .A(n33867), .B(n33868), .Z(n33866) );
  XNOR U42799 ( .A(y[3349]), .B(x[3349]), .Z(n33868) );
  XNOR U42800 ( .A(y[3350]), .B(x[3350]), .Z(n33867) );
  XNOR U42801 ( .A(y[3348]), .B(x[3348]), .Z(n33865) );
  XNOR U42802 ( .A(n33859), .B(n33860), .Z(n33870) );
  XNOR U42803 ( .A(y[3345]), .B(x[3345]), .Z(n33860) );
  XNOR U42804 ( .A(n33861), .B(n33862), .Z(n33859) );
  XNOR U42805 ( .A(y[3346]), .B(x[3346]), .Z(n33862) );
  XNOR U42806 ( .A(y[3347]), .B(x[3347]), .Z(n33861) );
  XNOR U42807 ( .A(n33852), .B(n33851), .Z(n33855) );
  XNOR U42808 ( .A(n33847), .B(n33848), .Z(n33851) );
  XNOR U42809 ( .A(y[3342]), .B(x[3342]), .Z(n33848) );
  XNOR U42810 ( .A(n33849), .B(n33850), .Z(n33847) );
  XNOR U42811 ( .A(y[3343]), .B(x[3343]), .Z(n33850) );
  XNOR U42812 ( .A(y[3344]), .B(x[3344]), .Z(n33849) );
  XNOR U42813 ( .A(n33841), .B(n33842), .Z(n33852) );
  XNOR U42814 ( .A(y[3339]), .B(x[3339]), .Z(n33842) );
  XNOR U42815 ( .A(n33843), .B(n33844), .Z(n33841) );
  XNOR U42816 ( .A(y[3340]), .B(x[3340]), .Z(n33844) );
  XNOR U42817 ( .A(y[3341]), .B(x[3341]), .Z(n33843) );
  XOR U42818 ( .A(n33817), .B(n33818), .Z(n33836) );
  XNOR U42819 ( .A(n33833), .B(n33834), .Z(n33818) );
  XNOR U42820 ( .A(n33828), .B(n33829), .Z(n33834) );
  XNOR U42821 ( .A(n33830), .B(n33831), .Z(n33829) );
  XNOR U42822 ( .A(y[3337]), .B(x[3337]), .Z(n33831) );
  XNOR U42823 ( .A(y[3338]), .B(x[3338]), .Z(n33830) );
  XNOR U42824 ( .A(y[3336]), .B(x[3336]), .Z(n33828) );
  XNOR U42825 ( .A(n33822), .B(n33823), .Z(n33833) );
  XNOR U42826 ( .A(y[3333]), .B(x[3333]), .Z(n33823) );
  XNOR U42827 ( .A(n33824), .B(n33825), .Z(n33822) );
  XNOR U42828 ( .A(y[3334]), .B(x[3334]), .Z(n33825) );
  XNOR U42829 ( .A(y[3335]), .B(x[3335]), .Z(n33824) );
  XOR U42830 ( .A(n33816), .B(n33815), .Z(n33817) );
  XNOR U42831 ( .A(n33811), .B(n33812), .Z(n33815) );
  XNOR U42832 ( .A(y[3330]), .B(x[3330]), .Z(n33812) );
  XNOR U42833 ( .A(n33813), .B(n33814), .Z(n33811) );
  XNOR U42834 ( .A(y[3331]), .B(x[3331]), .Z(n33814) );
  XNOR U42835 ( .A(y[3332]), .B(x[3332]), .Z(n33813) );
  XNOR U42836 ( .A(n33805), .B(n33806), .Z(n33816) );
  XNOR U42837 ( .A(y[3327]), .B(x[3327]), .Z(n33806) );
  XNOR U42838 ( .A(n33807), .B(n33808), .Z(n33805) );
  XNOR U42839 ( .A(y[3328]), .B(x[3328]), .Z(n33808) );
  XNOR U42840 ( .A(y[3329]), .B(x[3329]), .Z(n33807) );
  NAND U42841 ( .A(n33872), .B(n33873), .Z(N62390) );
  NANDN U42842 ( .A(n33874), .B(n33875), .Z(n33873) );
  OR U42843 ( .A(n33876), .B(n33877), .Z(n33875) );
  NAND U42844 ( .A(n33876), .B(n33877), .Z(n33872) );
  XOR U42845 ( .A(n33876), .B(n33878), .Z(N62389) );
  XNOR U42846 ( .A(n33874), .B(n33877), .Z(n33878) );
  AND U42847 ( .A(n33879), .B(n33880), .Z(n33877) );
  NANDN U42848 ( .A(n33881), .B(n33882), .Z(n33880) );
  NANDN U42849 ( .A(n33883), .B(n33884), .Z(n33882) );
  NANDN U42850 ( .A(n33884), .B(n33883), .Z(n33879) );
  NAND U42851 ( .A(n33885), .B(n33886), .Z(n33874) );
  NANDN U42852 ( .A(n33887), .B(n33888), .Z(n33886) );
  OR U42853 ( .A(n33889), .B(n33890), .Z(n33888) );
  NAND U42854 ( .A(n33890), .B(n33889), .Z(n33885) );
  AND U42855 ( .A(n33891), .B(n33892), .Z(n33876) );
  NANDN U42856 ( .A(n33893), .B(n33894), .Z(n33892) );
  NANDN U42857 ( .A(n33895), .B(n33896), .Z(n33894) );
  NANDN U42858 ( .A(n33896), .B(n33895), .Z(n33891) );
  XOR U42859 ( .A(n33890), .B(n33897), .Z(N62388) );
  XOR U42860 ( .A(n33887), .B(n33889), .Z(n33897) );
  XNOR U42861 ( .A(n33883), .B(n33898), .Z(n33889) );
  XNOR U42862 ( .A(n33881), .B(n33884), .Z(n33898) );
  NAND U42863 ( .A(n33899), .B(n33900), .Z(n33884) );
  NAND U42864 ( .A(n33901), .B(n33902), .Z(n33900) );
  OR U42865 ( .A(n33903), .B(n33904), .Z(n33901) );
  NANDN U42866 ( .A(n33905), .B(n33903), .Z(n33899) );
  IV U42867 ( .A(n33904), .Z(n33905) );
  NAND U42868 ( .A(n33906), .B(n33907), .Z(n33881) );
  NAND U42869 ( .A(n33908), .B(n33909), .Z(n33907) );
  NANDN U42870 ( .A(n33910), .B(n33911), .Z(n33908) );
  NANDN U42871 ( .A(n33911), .B(n33910), .Z(n33906) );
  AND U42872 ( .A(n33912), .B(n33913), .Z(n33883) );
  NAND U42873 ( .A(n33914), .B(n33915), .Z(n33913) );
  OR U42874 ( .A(n33916), .B(n33917), .Z(n33914) );
  NANDN U42875 ( .A(n33918), .B(n33916), .Z(n33912) );
  NAND U42876 ( .A(n33919), .B(n33920), .Z(n33887) );
  NANDN U42877 ( .A(n33921), .B(n33922), .Z(n33920) );
  OR U42878 ( .A(n33923), .B(n33924), .Z(n33922) );
  NANDN U42879 ( .A(n33925), .B(n33923), .Z(n33919) );
  IV U42880 ( .A(n33924), .Z(n33925) );
  XNOR U42881 ( .A(n33895), .B(n33926), .Z(n33890) );
  XNOR U42882 ( .A(n33893), .B(n33896), .Z(n33926) );
  NAND U42883 ( .A(n33927), .B(n33928), .Z(n33896) );
  NAND U42884 ( .A(n33929), .B(n33930), .Z(n33928) );
  OR U42885 ( .A(n33931), .B(n33932), .Z(n33929) );
  NANDN U42886 ( .A(n33933), .B(n33931), .Z(n33927) );
  IV U42887 ( .A(n33932), .Z(n33933) );
  NAND U42888 ( .A(n33934), .B(n33935), .Z(n33893) );
  NAND U42889 ( .A(n33936), .B(n33937), .Z(n33935) );
  NANDN U42890 ( .A(n33938), .B(n33939), .Z(n33936) );
  NANDN U42891 ( .A(n33939), .B(n33938), .Z(n33934) );
  AND U42892 ( .A(n33940), .B(n33941), .Z(n33895) );
  NAND U42893 ( .A(n33942), .B(n33943), .Z(n33941) );
  OR U42894 ( .A(n33944), .B(n33945), .Z(n33942) );
  NANDN U42895 ( .A(n33946), .B(n33944), .Z(n33940) );
  XNOR U42896 ( .A(n33921), .B(n33947), .Z(N62387) );
  XOR U42897 ( .A(n33923), .B(n33924), .Z(n33947) );
  XNOR U42898 ( .A(n33937), .B(n33948), .Z(n33924) );
  XOR U42899 ( .A(n33938), .B(n33939), .Z(n33948) );
  XOR U42900 ( .A(n33944), .B(n33949), .Z(n33939) );
  XOR U42901 ( .A(n33943), .B(n33946), .Z(n33949) );
  IV U42902 ( .A(n33945), .Z(n33946) );
  NAND U42903 ( .A(n33950), .B(n33951), .Z(n33945) );
  OR U42904 ( .A(n33952), .B(n33953), .Z(n33951) );
  OR U42905 ( .A(n33954), .B(n33955), .Z(n33950) );
  NAND U42906 ( .A(n33956), .B(n33957), .Z(n33943) );
  OR U42907 ( .A(n33958), .B(n33959), .Z(n33957) );
  OR U42908 ( .A(n33960), .B(n33961), .Z(n33956) );
  NOR U42909 ( .A(n33962), .B(n33963), .Z(n33944) );
  ANDN U42910 ( .B(n33964), .A(n33965), .Z(n33938) );
  XNOR U42911 ( .A(n33931), .B(n33966), .Z(n33937) );
  XNOR U42912 ( .A(n33930), .B(n33932), .Z(n33966) );
  NAND U42913 ( .A(n33967), .B(n33968), .Z(n33932) );
  OR U42914 ( .A(n33969), .B(n33970), .Z(n33968) );
  OR U42915 ( .A(n33971), .B(n33972), .Z(n33967) );
  NAND U42916 ( .A(n33973), .B(n33974), .Z(n33930) );
  OR U42917 ( .A(n33975), .B(n33976), .Z(n33974) );
  OR U42918 ( .A(n33977), .B(n33978), .Z(n33973) );
  ANDN U42919 ( .B(n33979), .A(n33980), .Z(n33931) );
  IV U42920 ( .A(n33981), .Z(n33979) );
  ANDN U42921 ( .B(n33982), .A(n33983), .Z(n33923) );
  XOR U42922 ( .A(n33909), .B(n33984), .Z(n33921) );
  XOR U42923 ( .A(n33910), .B(n33911), .Z(n33984) );
  XOR U42924 ( .A(n33916), .B(n33985), .Z(n33911) );
  XOR U42925 ( .A(n33915), .B(n33918), .Z(n33985) );
  IV U42926 ( .A(n33917), .Z(n33918) );
  NAND U42927 ( .A(n33986), .B(n33987), .Z(n33917) );
  OR U42928 ( .A(n33988), .B(n33989), .Z(n33987) );
  OR U42929 ( .A(n33990), .B(n33991), .Z(n33986) );
  NAND U42930 ( .A(n33992), .B(n33993), .Z(n33915) );
  OR U42931 ( .A(n33994), .B(n33995), .Z(n33993) );
  OR U42932 ( .A(n33996), .B(n33997), .Z(n33992) );
  NOR U42933 ( .A(n33998), .B(n33999), .Z(n33916) );
  ANDN U42934 ( .B(n34000), .A(n34001), .Z(n33910) );
  IV U42935 ( .A(n34002), .Z(n34000) );
  XNOR U42936 ( .A(n33903), .B(n34003), .Z(n33909) );
  XNOR U42937 ( .A(n33902), .B(n33904), .Z(n34003) );
  NAND U42938 ( .A(n34004), .B(n34005), .Z(n33904) );
  OR U42939 ( .A(n34006), .B(n34007), .Z(n34005) );
  OR U42940 ( .A(n34008), .B(n34009), .Z(n34004) );
  NAND U42941 ( .A(n34010), .B(n34011), .Z(n33902) );
  OR U42942 ( .A(n34012), .B(n34013), .Z(n34011) );
  OR U42943 ( .A(n34014), .B(n34015), .Z(n34010) );
  ANDN U42944 ( .B(n34016), .A(n34017), .Z(n33903) );
  IV U42945 ( .A(n34018), .Z(n34016) );
  XNOR U42946 ( .A(n33983), .B(n33982), .Z(N62386) );
  XOR U42947 ( .A(n34002), .B(n34001), .Z(n33982) );
  XNOR U42948 ( .A(n34017), .B(n34018), .Z(n34001) );
  XNOR U42949 ( .A(n34012), .B(n34013), .Z(n34018) );
  XNOR U42950 ( .A(n34014), .B(n34015), .Z(n34013) );
  XNOR U42951 ( .A(y[3325]), .B(x[3325]), .Z(n34015) );
  XNOR U42952 ( .A(y[3326]), .B(x[3326]), .Z(n34014) );
  XNOR U42953 ( .A(y[3324]), .B(x[3324]), .Z(n34012) );
  XNOR U42954 ( .A(n34006), .B(n34007), .Z(n34017) );
  XNOR U42955 ( .A(y[3321]), .B(x[3321]), .Z(n34007) );
  XNOR U42956 ( .A(n34008), .B(n34009), .Z(n34006) );
  XNOR U42957 ( .A(y[3322]), .B(x[3322]), .Z(n34009) );
  XNOR U42958 ( .A(y[3323]), .B(x[3323]), .Z(n34008) );
  XNOR U42959 ( .A(n33999), .B(n33998), .Z(n34002) );
  XNOR U42960 ( .A(n33994), .B(n33995), .Z(n33998) );
  XNOR U42961 ( .A(y[3318]), .B(x[3318]), .Z(n33995) );
  XNOR U42962 ( .A(n33996), .B(n33997), .Z(n33994) );
  XNOR U42963 ( .A(y[3319]), .B(x[3319]), .Z(n33997) );
  XNOR U42964 ( .A(y[3320]), .B(x[3320]), .Z(n33996) );
  XNOR U42965 ( .A(n33988), .B(n33989), .Z(n33999) );
  XNOR U42966 ( .A(y[3315]), .B(x[3315]), .Z(n33989) );
  XNOR U42967 ( .A(n33990), .B(n33991), .Z(n33988) );
  XNOR U42968 ( .A(y[3316]), .B(x[3316]), .Z(n33991) );
  XNOR U42969 ( .A(y[3317]), .B(x[3317]), .Z(n33990) );
  XOR U42970 ( .A(n33964), .B(n33965), .Z(n33983) );
  XNOR U42971 ( .A(n33980), .B(n33981), .Z(n33965) );
  XNOR U42972 ( .A(n33975), .B(n33976), .Z(n33981) );
  XNOR U42973 ( .A(n33977), .B(n33978), .Z(n33976) );
  XNOR U42974 ( .A(y[3313]), .B(x[3313]), .Z(n33978) );
  XNOR U42975 ( .A(y[3314]), .B(x[3314]), .Z(n33977) );
  XNOR U42976 ( .A(y[3312]), .B(x[3312]), .Z(n33975) );
  XNOR U42977 ( .A(n33969), .B(n33970), .Z(n33980) );
  XNOR U42978 ( .A(y[3309]), .B(x[3309]), .Z(n33970) );
  XNOR U42979 ( .A(n33971), .B(n33972), .Z(n33969) );
  XNOR U42980 ( .A(y[3310]), .B(x[3310]), .Z(n33972) );
  XNOR U42981 ( .A(y[3311]), .B(x[3311]), .Z(n33971) );
  XOR U42982 ( .A(n33963), .B(n33962), .Z(n33964) );
  XNOR U42983 ( .A(n33958), .B(n33959), .Z(n33962) );
  XNOR U42984 ( .A(y[3306]), .B(x[3306]), .Z(n33959) );
  XNOR U42985 ( .A(n33960), .B(n33961), .Z(n33958) );
  XNOR U42986 ( .A(y[3307]), .B(x[3307]), .Z(n33961) );
  XNOR U42987 ( .A(y[3308]), .B(x[3308]), .Z(n33960) );
  XNOR U42988 ( .A(n33952), .B(n33953), .Z(n33963) );
  XNOR U42989 ( .A(y[3303]), .B(x[3303]), .Z(n33953) );
  XNOR U42990 ( .A(n33954), .B(n33955), .Z(n33952) );
  XNOR U42991 ( .A(y[3304]), .B(x[3304]), .Z(n33955) );
  XNOR U42992 ( .A(y[3305]), .B(x[3305]), .Z(n33954) );
  NAND U42993 ( .A(n34019), .B(n34020), .Z(N62377) );
  NANDN U42994 ( .A(n34021), .B(n34022), .Z(n34020) );
  OR U42995 ( .A(n34023), .B(n34024), .Z(n34022) );
  NAND U42996 ( .A(n34023), .B(n34024), .Z(n34019) );
  XOR U42997 ( .A(n34023), .B(n34025), .Z(N62376) );
  XNOR U42998 ( .A(n34021), .B(n34024), .Z(n34025) );
  AND U42999 ( .A(n34026), .B(n34027), .Z(n34024) );
  NANDN U43000 ( .A(n34028), .B(n34029), .Z(n34027) );
  NANDN U43001 ( .A(n34030), .B(n34031), .Z(n34029) );
  NANDN U43002 ( .A(n34031), .B(n34030), .Z(n34026) );
  NAND U43003 ( .A(n34032), .B(n34033), .Z(n34021) );
  NANDN U43004 ( .A(n34034), .B(n34035), .Z(n34033) );
  OR U43005 ( .A(n34036), .B(n34037), .Z(n34035) );
  NAND U43006 ( .A(n34037), .B(n34036), .Z(n34032) );
  AND U43007 ( .A(n34038), .B(n34039), .Z(n34023) );
  NANDN U43008 ( .A(n34040), .B(n34041), .Z(n34039) );
  NANDN U43009 ( .A(n34042), .B(n34043), .Z(n34041) );
  NANDN U43010 ( .A(n34043), .B(n34042), .Z(n34038) );
  XOR U43011 ( .A(n34037), .B(n34044), .Z(N62375) );
  XOR U43012 ( .A(n34034), .B(n34036), .Z(n34044) );
  XNOR U43013 ( .A(n34030), .B(n34045), .Z(n34036) );
  XNOR U43014 ( .A(n34028), .B(n34031), .Z(n34045) );
  NAND U43015 ( .A(n34046), .B(n34047), .Z(n34031) );
  NAND U43016 ( .A(n34048), .B(n34049), .Z(n34047) );
  OR U43017 ( .A(n34050), .B(n34051), .Z(n34048) );
  NANDN U43018 ( .A(n34052), .B(n34050), .Z(n34046) );
  IV U43019 ( .A(n34051), .Z(n34052) );
  NAND U43020 ( .A(n34053), .B(n34054), .Z(n34028) );
  NAND U43021 ( .A(n34055), .B(n34056), .Z(n34054) );
  NANDN U43022 ( .A(n34057), .B(n34058), .Z(n34055) );
  NANDN U43023 ( .A(n34058), .B(n34057), .Z(n34053) );
  AND U43024 ( .A(n34059), .B(n34060), .Z(n34030) );
  NAND U43025 ( .A(n34061), .B(n34062), .Z(n34060) );
  OR U43026 ( .A(n34063), .B(n34064), .Z(n34061) );
  NANDN U43027 ( .A(n34065), .B(n34063), .Z(n34059) );
  NAND U43028 ( .A(n34066), .B(n34067), .Z(n34034) );
  NANDN U43029 ( .A(n34068), .B(n34069), .Z(n34067) );
  OR U43030 ( .A(n34070), .B(n34071), .Z(n34069) );
  NANDN U43031 ( .A(n34072), .B(n34070), .Z(n34066) );
  IV U43032 ( .A(n34071), .Z(n34072) );
  XNOR U43033 ( .A(n34042), .B(n34073), .Z(n34037) );
  XNOR U43034 ( .A(n34040), .B(n34043), .Z(n34073) );
  NAND U43035 ( .A(n34074), .B(n34075), .Z(n34043) );
  NAND U43036 ( .A(n34076), .B(n34077), .Z(n34075) );
  OR U43037 ( .A(n34078), .B(n34079), .Z(n34076) );
  NANDN U43038 ( .A(n34080), .B(n34078), .Z(n34074) );
  IV U43039 ( .A(n34079), .Z(n34080) );
  NAND U43040 ( .A(n34081), .B(n34082), .Z(n34040) );
  NAND U43041 ( .A(n34083), .B(n34084), .Z(n34082) );
  NANDN U43042 ( .A(n34085), .B(n34086), .Z(n34083) );
  NANDN U43043 ( .A(n34086), .B(n34085), .Z(n34081) );
  AND U43044 ( .A(n34087), .B(n34088), .Z(n34042) );
  NAND U43045 ( .A(n34089), .B(n34090), .Z(n34088) );
  OR U43046 ( .A(n34091), .B(n34092), .Z(n34089) );
  NANDN U43047 ( .A(n34093), .B(n34091), .Z(n34087) );
  XNOR U43048 ( .A(n34068), .B(n34094), .Z(N62374) );
  XOR U43049 ( .A(n34070), .B(n34071), .Z(n34094) );
  XNOR U43050 ( .A(n34084), .B(n34095), .Z(n34071) );
  XOR U43051 ( .A(n34085), .B(n34086), .Z(n34095) );
  XOR U43052 ( .A(n34091), .B(n34096), .Z(n34086) );
  XOR U43053 ( .A(n34090), .B(n34093), .Z(n34096) );
  IV U43054 ( .A(n34092), .Z(n34093) );
  NAND U43055 ( .A(n34097), .B(n34098), .Z(n34092) );
  OR U43056 ( .A(n34099), .B(n34100), .Z(n34098) );
  OR U43057 ( .A(n34101), .B(n34102), .Z(n34097) );
  NAND U43058 ( .A(n34103), .B(n34104), .Z(n34090) );
  OR U43059 ( .A(n34105), .B(n34106), .Z(n34104) );
  OR U43060 ( .A(n34107), .B(n34108), .Z(n34103) );
  NOR U43061 ( .A(n34109), .B(n34110), .Z(n34091) );
  ANDN U43062 ( .B(n34111), .A(n34112), .Z(n34085) );
  XNOR U43063 ( .A(n34078), .B(n34113), .Z(n34084) );
  XNOR U43064 ( .A(n34077), .B(n34079), .Z(n34113) );
  NAND U43065 ( .A(n34114), .B(n34115), .Z(n34079) );
  OR U43066 ( .A(n34116), .B(n34117), .Z(n34115) );
  OR U43067 ( .A(n34118), .B(n34119), .Z(n34114) );
  NAND U43068 ( .A(n34120), .B(n34121), .Z(n34077) );
  OR U43069 ( .A(n34122), .B(n34123), .Z(n34121) );
  OR U43070 ( .A(n34124), .B(n34125), .Z(n34120) );
  ANDN U43071 ( .B(n34126), .A(n34127), .Z(n34078) );
  IV U43072 ( .A(n34128), .Z(n34126) );
  ANDN U43073 ( .B(n34129), .A(n34130), .Z(n34070) );
  XOR U43074 ( .A(n34056), .B(n34131), .Z(n34068) );
  XOR U43075 ( .A(n34057), .B(n34058), .Z(n34131) );
  XOR U43076 ( .A(n34063), .B(n34132), .Z(n34058) );
  XOR U43077 ( .A(n34062), .B(n34065), .Z(n34132) );
  IV U43078 ( .A(n34064), .Z(n34065) );
  NAND U43079 ( .A(n34133), .B(n34134), .Z(n34064) );
  OR U43080 ( .A(n34135), .B(n34136), .Z(n34134) );
  OR U43081 ( .A(n34137), .B(n34138), .Z(n34133) );
  NAND U43082 ( .A(n34139), .B(n34140), .Z(n34062) );
  OR U43083 ( .A(n34141), .B(n34142), .Z(n34140) );
  OR U43084 ( .A(n34143), .B(n34144), .Z(n34139) );
  NOR U43085 ( .A(n34145), .B(n34146), .Z(n34063) );
  ANDN U43086 ( .B(n34147), .A(n34148), .Z(n34057) );
  IV U43087 ( .A(n34149), .Z(n34147) );
  XNOR U43088 ( .A(n34050), .B(n34150), .Z(n34056) );
  XNOR U43089 ( .A(n34049), .B(n34051), .Z(n34150) );
  NAND U43090 ( .A(n34151), .B(n34152), .Z(n34051) );
  OR U43091 ( .A(n34153), .B(n34154), .Z(n34152) );
  OR U43092 ( .A(n34155), .B(n34156), .Z(n34151) );
  NAND U43093 ( .A(n34157), .B(n34158), .Z(n34049) );
  OR U43094 ( .A(n34159), .B(n34160), .Z(n34158) );
  OR U43095 ( .A(n34161), .B(n34162), .Z(n34157) );
  ANDN U43096 ( .B(n34163), .A(n34164), .Z(n34050) );
  IV U43097 ( .A(n34165), .Z(n34163) );
  XNOR U43098 ( .A(n34130), .B(n34129), .Z(N62373) );
  XOR U43099 ( .A(n34149), .B(n34148), .Z(n34129) );
  XNOR U43100 ( .A(n34164), .B(n34165), .Z(n34148) );
  XNOR U43101 ( .A(n34159), .B(n34160), .Z(n34165) );
  XNOR U43102 ( .A(n34161), .B(n34162), .Z(n34160) );
  XNOR U43103 ( .A(y[3301]), .B(x[3301]), .Z(n34162) );
  XNOR U43104 ( .A(y[3302]), .B(x[3302]), .Z(n34161) );
  XNOR U43105 ( .A(y[3300]), .B(x[3300]), .Z(n34159) );
  XNOR U43106 ( .A(n34153), .B(n34154), .Z(n34164) );
  XNOR U43107 ( .A(y[3297]), .B(x[3297]), .Z(n34154) );
  XNOR U43108 ( .A(n34155), .B(n34156), .Z(n34153) );
  XNOR U43109 ( .A(y[3298]), .B(x[3298]), .Z(n34156) );
  XNOR U43110 ( .A(y[3299]), .B(x[3299]), .Z(n34155) );
  XNOR U43111 ( .A(n34146), .B(n34145), .Z(n34149) );
  XNOR U43112 ( .A(n34141), .B(n34142), .Z(n34145) );
  XNOR U43113 ( .A(y[3294]), .B(x[3294]), .Z(n34142) );
  XNOR U43114 ( .A(n34143), .B(n34144), .Z(n34141) );
  XNOR U43115 ( .A(y[3295]), .B(x[3295]), .Z(n34144) );
  XNOR U43116 ( .A(y[3296]), .B(x[3296]), .Z(n34143) );
  XNOR U43117 ( .A(n34135), .B(n34136), .Z(n34146) );
  XNOR U43118 ( .A(y[3291]), .B(x[3291]), .Z(n34136) );
  XNOR U43119 ( .A(n34137), .B(n34138), .Z(n34135) );
  XNOR U43120 ( .A(y[3292]), .B(x[3292]), .Z(n34138) );
  XNOR U43121 ( .A(y[3293]), .B(x[3293]), .Z(n34137) );
  XOR U43122 ( .A(n34111), .B(n34112), .Z(n34130) );
  XNOR U43123 ( .A(n34127), .B(n34128), .Z(n34112) );
  XNOR U43124 ( .A(n34122), .B(n34123), .Z(n34128) );
  XNOR U43125 ( .A(n34124), .B(n34125), .Z(n34123) );
  XNOR U43126 ( .A(y[3289]), .B(x[3289]), .Z(n34125) );
  XNOR U43127 ( .A(y[3290]), .B(x[3290]), .Z(n34124) );
  XNOR U43128 ( .A(y[3288]), .B(x[3288]), .Z(n34122) );
  XNOR U43129 ( .A(n34116), .B(n34117), .Z(n34127) );
  XNOR U43130 ( .A(y[3285]), .B(x[3285]), .Z(n34117) );
  XNOR U43131 ( .A(n34118), .B(n34119), .Z(n34116) );
  XNOR U43132 ( .A(y[3286]), .B(x[3286]), .Z(n34119) );
  XNOR U43133 ( .A(y[3287]), .B(x[3287]), .Z(n34118) );
  XOR U43134 ( .A(n34110), .B(n34109), .Z(n34111) );
  XNOR U43135 ( .A(n34105), .B(n34106), .Z(n34109) );
  XNOR U43136 ( .A(y[3282]), .B(x[3282]), .Z(n34106) );
  XNOR U43137 ( .A(n34107), .B(n34108), .Z(n34105) );
  XNOR U43138 ( .A(y[3283]), .B(x[3283]), .Z(n34108) );
  XNOR U43139 ( .A(y[3284]), .B(x[3284]), .Z(n34107) );
  XNOR U43140 ( .A(n34099), .B(n34100), .Z(n34110) );
  XNOR U43141 ( .A(y[3279]), .B(x[3279]), .Z(n34100) );
  XNOR U43142 ( .A(n34101), .B(n34102), .Z(n34099) );
  XNOR U43143 ( .A(y[3280]), .B(x[3280]), .Z(n34102) );
  XNOR U43144 ( .A(y[3281]), .B(x[3281]), .Z(n34101) );
  NAND U43145 ( .A(n34166), .B(n34167), .Z(N62364) );
  NANDN U43146 ( .A(n34168), .B(n34169), .Z(n34167) );
  OR U43147 ( .A(n34170), .B(n34171), .Z(n34169) );
  NAND U43148 ( .A(n34170), .B(n34171), .Z(n34166) );
  XOR U43149 ( .A(n34170), .B(n34172), .Z(N62363) );
  XNOR U43150 ( .A(n34168), .B(n34171), .Z(n34172) );
  AND U43151 ( .A(n34173), .B(n34174), .Z(n34171) );
  NANDN U43152 ( .A(n34175), .B(n34176), .Z(n34174) );
  NANDN U43153 ( .A(n34177), .B(n34178), .Z(n34176) );
  NANDN U43154 ( .A(n34178), .B(n34177), .Z(n34173) );
  NAND U43155 ( .A(n34179), .B(n34180), .Z(n34168) );
  NANDN U43156 ( .A(n34181), .B(n34182), .Z(n34180) );
  OR U43157 ( .A(n34183), .B(n34184), .Z(n34182) );
  NAND U43158 ( .A(n34184), .B(n34183), .Z(n34179) );
  AND U43159 ( .A(n34185), .B(n34186), .Z(n34170) );
  NANDN U43160 ( .A(n34187), .B(n34188), .Z(n34186) );
  NANDN U43161 ( .A(n34189), .B(n34190), .Z(n34188) );
  NANDN U43162 ( .A(n34190), .B(n34189), .Z(n34185) );
  XOR U43163 ( .A(n34184), .B(n34191), .Z(N62362) );
  XOR U43164 ( .A(n34181), .B(n34183), .Z(n34191) );
  XNOR U43165 ( .A(n34177), .B(n34192), .Z(n34183) );
  XNOR U43166 ( .A(n34175), .B(n34178), .Z(n34192) );
  NAND U43167 ( .A(n34193), .B(n34194), .Z(n34178) );
  NAND U43168 ( .A(n34195), .B(n34196), .Z(n34194) );
  OR U43169 ( .A(n34197), .B(n34198), .Z(n34195) );
  NANDN U43170 ( .A(n34199), .B(n34197), .Z(n34193) );
  IV U43171 ( .A(n34198), .Z(n34199) );
  NAND U43172 ( .A(n34200), .B(n34201), .Z(n34175) );
  NAND U43173 ( .A(n34202), .B(n34203), .Z(n34201) );
  NANDN U43174 ( .A(n34204), .B(n34205), .Z(n34202) );
  NANDN U43175 ( .A(n34205), .B(n34204), .Z(n34200) );
  AND U43176 ( .A(n34206), .B(n34207), .Z(n34177) );
  NAND U43177 ( .A(n34208), .B(n34209), .Z(n34207) );
  OR U43178 ( .A(n34210), .B(n34211), .Z(n34208) );
  NANDN U43179 ( .A(n34212), .B(n34210), .Z(n34206) );
  NAND U43180 ( .A(n34213), .B(n34214), .Z(n34181) );
  NANDN U43181 ( .A(n34215), .B(n34216), .Z(n34214) );
  OR U43182 ( .A(n34217), .B(n34218), .Z(n34216) );
  NANDN U43183 ( .A(n34219), .B(n34217), .Z(n34213) );
  IV U43184 ( .A(n34218), .Z(n34219) );
  XNOR U43185 ( .A(n34189), .B(n34220), .Z(n34184) );
  XNOR U43186 ( .A(n34187), .B(n34190), .Z(n34220) );
  NAND U43187 ( .A(n34221), .B(n34222), .Z(n34190) );
  NAND U43188 ( .A(n34223), .B(n34224), .Z(n34222) );
  OR U43189 ( .A(n34225), .B(n34226), .Z(n34223) );
  NANDN U43190 ( .A(n34227), .B(n34225), .Z(n34221) );
  IV U43191 ( .A(n34226), .Z(n34227) );
  NAND U43192 ( .A(n34228), .B(n34229), .Z(n34187) );
  NAND U43193 ( .A(n34230), .B(n34231), .Z(n34229) );
  NANDN U43194 ( .A(n34232), .B(n34233), .Z(n34230) );
  NANDN U43195 ( .A(n34233), .B(n34232), .Z(n34228) );
  AND U43196 ( .A(n34234), .B(n34235), .Z(n34189) );
  NAND U43197 ( .A(n34236), .B(n34237), .Z(n34235) );
  OR U43198 ( .A(n34238), .B(n34239), .Z(n34236) );
  NANDN U43199 ( .A(n34240), .B(n34238), .Z(n34234) );
  XNOR U43200 ( .A(n34215), .B(n34241), .Z(N62361) );
  XOR U43201 ( .A(n34217), .B(n34218), .Z(n34241) );
  XNOR U43202 ( .A(n34231), .B(n34242), .Z(n34218) );
  XOR U43203 ( .A(n34232), .B(n34233), .Z(n34242) );
  XOR U43204 ( .A(n34238), .B(n34243), .Z(n34233) );
  XOR U43205 ( .A(n34237), .B(n34240), .Z(n34243) );
  IV U43206 ( .A(n34239), .Z(n34240) );
  NAND U43207 ( .A(n34244), .B(n34245), .Z(n34239) );
  OR U43208 ( .A(n34246), .B(n34247), .Z(n34245) );
  OR U43209 ( .A(n34248), .B(n34249), .Z(n34244) );
  NAND U43210 ( .A(n34250), .B(n34251), .Z(n34237) );
  OR U43211 ( .A(n34252), .B(n34253), .Z(n34251) );
  OR U43212 ( .A(n34254), .B(n34255), .Z(n34250) );
  NOR U43213 ( .A(n34256), .B(n34257), .Z(n34238) );
  ANDN U43214 ( .B(n34258), .A(n34259), .Z(n34232) );
  XNOR U43215 ( .A(n34225), .B(n34260), .Z(n34231) );
  XNOR U43216 ( .A(n34224), .B(n34226), .Z(n34260) );
  NAND U43217 ( .A(n34261), .B(n34262), .Z(n34226) );
  OR U43218 ( .A(n34263), .B(n34264), .Z(n34262) );
  OR U43219 ( .A(n34265), .B(n34266), .Z(n34261) );
  NAND U43220 ( .A(n34267), .B(n34268), .Z(n34224) );
  OR U43221 ( .A(n34269), .B(n34270), .Z(n34268) );
  OR U43222 ( .A(n34271), .B(n34272), .Z(n34267) );
  ANDN U43223 ( .B(n34273), .A(n34274), .Z(n34225) );
  IV U43224 ( .A(n34275), .Z(n34273) );
  ANDN U43225 ( .B(n34276), .A(n34277), .Z(n34217) );
  XOR U43226 ( .A(n34203), .B(n34278), .Z(n34215) );
  XOR U43227 ( .A(n34204), .B(n34205), .Z(n34278) );
  XOR U43228 ( .A(n34210), .B(n34279), .Z(n34205) );
  XOR U43229 ( .A(n34209), .B(n34212), .Z(n34279) );
  IV U43230 ( .A(n34211), .Z(n34212) );
  NAND U43231 ( .A(n34280), .B(n34281), .Z(n34211) );
  OR U43232 ( .A(n34282), .B(n34283), .Z(n34281) );
  OR U43233 ( .A(n34284), .B(n34285), .Z(n34280) );
  NAND U43234 ( .A(n34286), .B(n34287), .Z(n34209) );
  OR U43235 ( .A(n34288), .B(n34289), .Z(n34287) );
  OR U43236 ( .A(n34290), .B(n34291), .Z(n34286) );
  NOR U43237 ( .A(n34292), .B(n34293), .Z(n34210) );
  ANDN U43238 ( .B(n34294), .A(n34295), .Z(n34204) );
  IV U43239 ( .A(n34296), .Z(n34294) );
  XNOR U43240 ( .A(n34197), .B(n34297), .Z(n34203) );
  XNOR U43241 ( .A(n34196), .B(n34198), .Z(n34297) );
  NAND U43242 ( .A(n34298), .B(n34299), .Z(n34198) );
  OR U43243 ( .A(n34300), .B(n34301), .Z(n34299) );
  OR U43244 ( .A(n34302), .B(n34303), .Z(n34298) );
  NAND U43245 ( .A(n34304), .B(n34305), .Z(n34196) );
  OR U43246 ( .A(n34306), .B(n34307), .Z(n34305) );
  OR U43247 ( .A(n34308), .B(n34309), .Z(n34304) );
  ANDN U43248 ( .B(n34310), .A(n34311), .Z(n34197) );
  IV U43249 ( .A(n34312), .Z(n34310) );
  XNOR U43250 ( .A(n34277), .B(n34276), .Z(N62360) );
  XOR U43251 ( .A(n34296), .B(n34295), .Z(n34276) );
  XNOR U43252 ( .A(n34311), .B(n34312), .Z(n34295) );
  XNOR U43253 ( .A(n34306), .B(n34307), .Z(n34312) );
  XNOR U43254 ( .A(n34308), .B(n34309), .Z(n34307) );
  XNOR U43255 ( .A(y[3277]), .B(x[3277]), .Z(n34309) );
  XNOR U43256 ( .A(y[3278]), .B(x[3278]), .Z(n34308) );
  XNOR U43257 ( .A(y[3276]), .B(x[3276]), .Z(n34306) );
  XNOR U43258 ( .A(n34300), .B(n34301), .Z(n34311) );
  XNOR U43259 ( .A(y[3273]), .B(x[3273]), .Z(n34301) );
  XNOR U43260 ( .A(n34302), .B(n34303), .Z(n34300) );
  XNOR U43261 ( .A(y[3274]), .B(x[3274]), .Z(n34303) );
  XNOR U43262 ( .A(y[3275]), .B(x[3275]), .Z(n34302) );
  XNOR U43263 ( .A(n34293), .B(n34292), .Z(n34296) );
  XNOR U43264 ( .A(n34288), .B(n34289), .Z(n34292) );
  XNOR U43265 ( .A(y[3270]), .B(x[3270]), .Z(n34289) );
  XNOR U43266 ( .A(n34290), .B(n34291), .Z(n34288) );
  XNOR U43267 ( .A(y[3271]), .B(x[3271]), .Z(n34291) );
  XNOR U43268 ( .A(y[3272]), .B(x[3272]), .Z(n34290) );
  XNOR U43269 ( .A(n34282), .B(n34283), .Z(n34293) );
  XNOR U43270 ( .A(y[3267]), .B(x[3267]), .Z(n34283) );
  XNOR U43271 ( .A(n34284), .B(n34285), .Z(n34282) );
  XNOR U43272 ( .A(y[3268]), .B(x[3268]), .Z(n34285) );
  XNOR U43273 ( .A(y[3269]), .B(x[3269]), .Z(n34284) );
  XOR U43274 ( .A(n34258), .B(n34259), .Z(n34277) );
  XNOR U43275 ( .A(n34274), .B(n34275), .Z(n34259) );
  XNOR U43276 ( .A(n34269), .B(n34270), .Z(n34275) );
  XNOR U43277 ( .A(n34271), .B(n34272), .Z(n34270) );
  XNOR U43278 ( .A(y[3265]), .B(x[3265]), .Z(n34272) );
  XNOR U43279 ( .A(y[3266]), .B(x[3266]), .Z(n34271) );
  XNOR U43280 ( .A(y[3264]), .B(x[3264]), .Z(n34269) );
  XNOR U43281 ( .A(n34263), .B(n34264), .Z(n34274) );
  XNOR U43282 ( .A(y[3261]), .B(x[3261]), .Z(n34264) );
  XNOR U43283 ( .A(n34265), .B(n34266), .Z(n34263) );
  XNOR U43284 ( .A(y[3262]), .B(x[3262]), .Z(n34266) );
  XNOR U43285 ( .A(y[3263]), .B(x[3263]), .Z(n34265) );
  XOR U43286 ( .A(n34257), .B(n34256), .Z(n34258) );
  XNOR U43287 ( .A(n34252), .B(n34253), .Z(n34256) );
  XNOR U43288 ( .A(y[3258]), .B(x[3258]), .Z(n34253) );
  XNOR U43289 ( .A(n34254), .B(n34255), .Z(n34252) );
  XNOR U43290 ( .A(y[3259]), .B(x[3259]), .Z(n34255) );
  XNOR U43291 ( .A(y[3260]), .B(x[3260]), .Z(n34254) );
  XNOR U43292 ( .A(n34246), .B(n34247), .Z(n34257) );
  XNOR U43293 ( .A(y[3255]), .B(x[3255]), .Z(n34247) );
  XNOR U43294 ( .A(n34248), .B(n34249), .Z(n34246) );
  XNOR U43295 ( .A(y[3256]), .B(x[3256]), .Z(n34249) );
  XNOR U43296 ( .A(y[3257]), .B(x[3257]), .Z(n34248) );
  NAND U43297 ( .A(n34313), .B(n34314), .Z(N62351) );
  NANDN U43298 ( .A(n34315), .B(n34316), .Z(n34314) );
  OR U43299 ( .A(n34317), .B(n34318), .Z(n34316) );
  NAND U43300 ( .A(n34317), .B(n34318), .Z(n34313) );
  XOR U43301 ( .A(n34317), .B(n34319), .Z(N62350) );
  XNOR U43302 ( .A(n34315), .B(n34318), .Z(n34319) );
  AND U43303 ( .A(n34320), .B(n34321), .Z(n34318) );
  NANDN U43304 ( .A(n34322), .B(n34323), .Z(n34321) );
  NANDN U43305 ( .A(n34324), .B(n34325), .Z(n34323) );
  NANDN U43306 ( .A(n34325), .B(n34324), .Z(n34320) );
  NAND U43307 ( .A(n34326), .B(n34327), .Z(n34315) );
  NANDN U43308 ( .A(n34328), .B(n34329), .Z(n34327) );
  OR U43309 ( .A(n34330), .B(n34331), .Z(n34329) );
  NAND U43310 ( .A(n34331), .B(n34330), .Z(n34326) );
  AND U43311 ( .A(n34332), .B(n34333), .Z(n34317) );
  NANDN U43312 ( .A(n34334), .B(n34335), .Z(n34333) );
  NANDN U43313 ( .A(n34336), .B(n34337), .Z(n34335) );
  NANDN U43314 ( .A(n34337), .B(n34336), .Z(n34332) );
  XOR U43315 ( .A(n34331), .B(n34338), .Z(N62349) );
  XOR U43316 ( .A(n34328), .B(n34330), .Z(n34338) );
  XNOR U43317 ( .A(n34324), .B(n34339), .Z(n34330) );
  XNOR U43318 ( .A(n34322), .B(n34325), .Z(n34339) );
  NAND U43319 ( .A(n34340), .B(n34341), .Z(n34325) );
  NAND U43320 ( .A(n34342), .B(n34343), .Z(n34341) );
  OR U43321 ( .A(n34344), .B(n34345), .Z(n34342) );
  NANDN U43322 ( .A(n34346), .B(n34344), .Z(n34340) );
  IV U43323 ( .A(n34345), .Z(n34346) );
  NAND U43324 ( .A(n34347), .B(n34348), .Z(n34322) );
  NAND U43325 ( .A(n34349), .B(n34350), .Z(n34348) );
  NANDN U43326 ( .A(n34351), .B(n34352), .Z(n34349) );
  NANDN U43327 ( .A(n34352), .B(n34351), .Z(n34347) );
  AND U43328 ( .A(n34353), .B(n34354), .Z(n34324) );
  NAND U43329 ( .A(n34355), .B(n34356), .Z(n34354) );
  OR U43330 ( .A(n34357), .B(n34358), .Z(n34355) );
  NANDN U43331 ( .A(n34359), .B(n34357), .Z(n34353) );
  NAND U43332 ( .A(n34360), .B(n34361), .Z(n34328) );
  NANDN U43333 ( .A(n34362), .B(n34363), .Z(n34361) );
  OR U43334 ( .A(n34364), .B(n34365), .Z(n34363) );
  NANDN U43335 ( .A(n34366), .B(n34364), .Z(n34360) );
  IV U43336 ( .A(n34365), .Z(n34366) );
  XNOR U43337 ( .A(n34336), .B(n34367), .Z(n34331) );
  XNOR U43338 ( .A(n34334), .B(n34337), .Z(n34367) );
  NAND U43339 ( .A(n34368), .B(n34369), .Z(n34337) );
  NAND U43340 ( .A(n34370), .B(n34371), .Z(n34369) );
  OR U43341 ( .A(n34372), .B(n34373), .Z(n34370) );
  NANDN U43342 ( .A(n34374), .B(n34372), .Z(n34368) );
  IV U43343 ( .A(n34373), .Z(n34374) );
  NAND U43344 ( .A(n34375), .B(n34376), .Z(n34334) );
  NAND U43345 ( .A(n34377), .B(n34378), .Z(n34376) );
  NANDN U43346 ( .A(n34379), .B(n34380), .Z(n34377) );
  NANDN U43347 ( .A(n34380), .B(n34379), .Z(n34375) );
  AND U43348 ( .A(n34381), .B(n34382), .Z(n34336) );
  NAND U43349 ( .A(n34383), .B(n34384), .Z(n34382) );
  OR U43350 ( .A(n34385), .B(n34386), .Z(n34383) );
  NANDN U43351 ( .A(n34387), .B(n34385), .Z(n34381) );
  XNOR U43352 ( .A(n34362), .B(n34388), .Z(N62348) );
  XOR U43353 ( .A(n34364), .B(n34365), .Z(n34388) );
  XNOR U43354 ( .A(n34378), .B(n34389), .Z(n34365) );
  XOR U43355 ( .A(n34379), .B(n34380), .Z(n34389) );
  XOR U43356 ( .A(n34385), .B(n34390), .Z(n34380) );
  XOR U43357 ( .A(n34384), .B(n34387), .Z(n34390) );
  IV U43358 ( .A(n34386), .Z(n34387) );
  NAND U43359 ( .A(n34391), .B(n34392), .Z(n34386) );
  OR U43360 ( .A(n34393), .B(n34394), .Z(n34392) );
  OR U43361 ( .A(n34395), .B(n34396), .Z(n34391) );
  NAND U43362 ( .A(n34397), .B(n34398), .Z(n34384) );
  OR U43363 ( .A(n34399), .B(n34400), .Z(n34398) );
  OR U43364 ( .A(n34401), .B(n34402), .Z(n34397) );
  NOR U43365 ( .A(n34403), .B(n34404), .Z(n34385) );
  ANDN U43366 ( .B(n34405), .A(n34406), .Z(n34379) );
  XNOR U43367 ( .A(n34372), .B(n34407), .Z(n34378) );
  XNOR U43368 ( .A(n34371), .B(n34373), .Z(n34407) );
  NAND U43369 ( .A(n34408), .B(n34409), .Z(n34373) );
  OR U43370 ( .A(n34410), .B(n34411), .Z(n34409) );
  OR U43371 ( .A(n34412), .B(n34413), .Z(n34408) );
  NAND U43372 ( .A(n34414), .B(n34415), .Z(n34371) );
  OR U43373 ( .A(n34416), .B(n34417), .Z(n34415) );
  OR U43374 ( .A(n34418), .B(n34419), .Z(n34414) );
  ANDN U43375 ( .B(n34420), .A(n34421), .Z(n34372) );
  IV U43376 ( .A(n34422), .Z(n34420) );
  ANDN U43377 ( .B(n34423), .A(n34424), .Z(n34364) );
  XOR U43378 ( .A(n34350), .B(n34425), .Z(n34362) );
  XOR U43379 ( .A(n34351), .B(n34352), .Z(n34425) );
  XOR U43380 ( .A(n34357), .B(n34426), .Z(n34352) );
  XOR U43381 ( .A(n34356), .B(n34359), .Z(n34426) );
  IV U43382 ( .A(n34358), .Z(n34359) );
  NAND U43383 ( .A(n34427), .B(n34428), .Z(n34358) );
  OR U43384 ( .A(n34429), .B(n34430), .Z(n34428) );
  OR U43385 ( .A(n34431), .B(n34432), .Z(n34427) );
  NAND U43386 ( .A(n34433), .B(n34434), .Z(n34356) );
  OR U43387 ( .A(n34435), .B(n34436), .Z(n34434) );
  OR U43388 ( .A(n34437), .B(n34438), .Z(n34433) );
  NOR U43389 ( .A(n34439), .B(n34440), .Z(n34357) );
  ANDN U43390 ( .B(n34441), .A(n34442), .Z(n34351) );
  IV U43391 ( .A(n34443), .Z(n34441) );
  XNOR U43392 ( .A(n34344), .B(n34444), .Z(n34350) );
  XNOR U43393 ( .A(n34343), .B(n34345), .Z(n34444) );
  NAND U43394 ( .A(n34445), .B(n34446), .Z(n34345) );
  OR U43395 ( .A(n34447), .B(n34448), .Z(n34446) );
  OR U43396 ( .A(n34449), .B(n34450), .Z(n34445) );
  NAND U43397 ( .A(n34451), .B(n34452), .Z(n34343) );
  OR U43398 ( .A(n34453), .B(n34454), .Z(n34452) );
  OR U43399 ( .A(n34455), .B(n34456), .Z(n34451) );
  ANDN U43400 ( .B(n34457), .A(n34458), .Z(n34344) );
  IV U43401 ( .A(n34459), .Z(n34457) );
  XNOR U43402 ( .A(n34424), .B(n34423), .Z(N62347) );
  XOR U43403 ( .A(n34443), .B(n34442), .Z(n34423) );
  XNOR U43404 ( .A(n34458), .B(n34459), .Z(n34442) );
  XNOR U43405 ( .A(n34453), .B(n34454), .Z(n34459) );
  XNOR U43406 ( .A(n34455), .B(n34456), .Z(n34454) );
  XNOR U43407 ( .A(y[3253]), .B(x[3253]), .Z(n34456) );
  XNOR U43408 ( .A(y[3254]), .B(x[3254]), .Z(n34455) );
  XNOR U43409 ( .A(y[3252]), .B(x[3252]), .Z(n34453) );
  XNOR U43410 ( .A(n34447), .B(n34448), .Z(n34458) );
  XNOR U43411 ( .A(y[3249]), .B(x[3249]), .Z(n34448) );
  XNOR U43412 ( .A(n34449), .B(n34450), .Z(n34447) );
  XNOR U43413 ( .A(y[3250]), .B(x[3250]), .Z(n34450) );
  XNOR U43414 ( .A(y[3251]), .B(x[3251]), .Z(n34449) );
  XNOR U43415 ( .A(n34440), .B(n34439), .Z(n34443) );
  XNOR U43416 ( .A(n34435), .B(n34436), .Z(n34439) );
  XNOR U43417 ( .A(y[3246]), .B(x[3246]), .Z(n34436) );
  XNOR U43418 ( .A(n34437), .B(n34438), .Z(n34435) );
  XNOR U43419 ( .A(y[3247]), .B(x[3247]), .Z(n34438) );
  XNOR U43420 ( .A(y[3248]), .B(x[3248]), .Z(n34437) );
  XNOR U43421 ( .A(n34429), .B(n34430), .Z(n34440) );
  XNOR U43422 ( .A(y[3243]), .B(x[3243]), .Z(n34430) );
  XNOR U43423 ( .A(n34431), .B(n34432), .Z(n34429) );
  XNOR U43424 ( .A(y[3244]), .B(x[3244]), .Z(n34432) );
  XNOR U43425 ( .A(y[3245]), .B(x[3245]), .Z(n34431) );
  XOR U43426 ( .A(n34405), .B(n34406), .Z(n34424) );
  XNOR U43427 ( .A(n34421), .B(n34422), .Z(n34406) );
  XNOR U43428 ( .A(n34416), .B(n34417), .Z(n34422) );
  XNOR U43429 ( .A(n34418), .B(n34419), .Z(n34417) );
  XNOR U43430 ( .A(y[3241]), .B(x[3241]), .Z(n34419) );
  XNOR U43431 ( .A(y[3242]), .B(x[3242]), .Z(n34418) );
  XNOR U43432 ( .A(y[3240]), .B(x[3240]), .Z(n34416) );
  XNOR U43433 ( .A(n34410), .B(n34411), .Z(n34421) );
  XNOR U43434 ( .A(y[3237]), .B(x[3237]), .Z(n34411) );
  XNOR U43435 ( .A(n34412), .B(n34413), .Z(n34410) );
  XNOR U43436 ( .A(y[3238]), .B(x[3238]), .Z(n34413) );
  XNOR U43437 ( .A(y[3239]), .B(x[3239]), .Z(n34412) );
  XOR U43438 ( .A(n34404), .B(n34403), .Z(n34405) );
  XNOR U43439 ( .A(n34399), .B(n34400), .Z(n34403) );
  XNOR U43440 ( .A(y[3234]), .B(x[3234]), .Z(n34400) );
  XNOR U43441 ( .A(n34401), .B(n34402), .Z(n34399) );
  XNOR U43442 ( .A(y[3235]), .B(x[3235]), .Z(n34402) );
  XNOR U43443 ( .A(y[3236]), .B(x[3236]), .Z(n34401) );
  XNOR U43444 ( .A(n34393), .B(n34394), .Z(n34404) );
  XNOR U43445 ( .A(y[3231]), .B(x[3231]), .Z(n34394) );
  XNOR U43446 ( .A(n34395), .B(n34396), .Z(n34393) );
  XNOR U43447 ( .A(y[3232]), .B(x[3232]), .Z(n34396) );
  XNOR U43448 ( .A(y[3233]), .B(x[3233]), .Z(n34395) );
  NAND U43449 ( .A(n34460), .B(n34461), .Z(N62338) );
  NANDN U43450 ( .A(n34462), .B(n34463), .Z(n34461) );
  OR U43451 ( .A(n34464), .B(n34465), .Z(n34463) );
  NAND U43452 ( .A(n34464), .B(n34465), .Z(n34460) );
  XOR U43453 ( .A(n34464), .B(n34466), .Z(N62337) );
  XNOR U43454 ( .A(n34462), .B(n34465), .Z(n34466) );
  AND U43455 ( .A(n34467), .B(n34468), .Z(n34465) );
  NANDN U43456 ( .A(n34469), .B(n34470), .Z(n34468) );
  NANDN U43457 ( .A(n34471), .B(n34472), .Z(n34470) );
  NANDN U43458 ( .A(n34472), .B(n34471), .Z(n34467) );
  NAND U43459 ( .A(n34473), .B(n34474), .Z(n34462) );
  NANDN U43460 ( .A(n34475), .B(n34476), .Z(n34474) );
  OR U43461 ( .A(n34477), .B(n34478), .Z(n34476) );
  NAND U43462 ( .A(n34478), .B(n34477), .Z(n34473) );
  AND U43463 ( .A(n34479), .B(n34480), .Z(n34464) );
  NANDN U43464 ( .A(n34481), .B(n34482), .Z(n34480) );
  NANDN U43465 ( .A(n34483), .B(n34484), .Z(n34482) );
  NANDN U43466 ( .A(n34484), .B(n34483), .Z(n34479) );
  XOR U43467 ( .A(n34478), .B(n34485), .Z(N62336) );
  XOR U43468 ( .A(n34475), .B(n34477), .Z(n34485) );
  XNOR U43469 ( .A(n34471), .B(n34486), .Z(n34477) );
  XNOR U43470 ( .A(n34469), .B(n34472), .Z(n34486) );
  NAND U43471 ( .A(n34487), .B(n34488), .Z(n34472) );
  NAND U43472 ( .A(n34489), .B(n34490), .Z(n34488) );
  OR U43473 ( .A(n34491), .B(n34492), .Z(n34489) );
  NANDN U43474 ( .A(n34493), .B(n34491), .Z(n34487) );
  IV U43475 ( .A(n34492), .Z(n34493) );
  NAND U43476 ( .A(n34494), .B(n34495), .Z(n34469) );
  NAND U43477 ( .A(n34496), .B(n34497), .Z(n34495) );
  NANDN U43478 ( .A(n34498), .B(n34499), .Z(n34496) );
  NANDN U43479 ( .A(n34499), .B(n34498), .Z(n34494) );
  AND U43480 ( .A(n34500), .B(n34501), .Z(n34471) );
  NAND U43481 ( .A(n34502), .B(n34503), .Z(n34501) );
  OR U43482 ( .A(n34504), .B(n34505), .Z(n34502) );
  NANDN U43483 ( .A(n34506), .B(n34504), .Z(n34500) );
  NAND U43484 ( .A(n34507), .B(n34508), .Z(n34475) );
  NANDN U43485 ( .A(n34509), .B(n34510), .Z(n34508) );
  OR U43486 ( .A(n34511), .B(n34512), .Z(n34510) );
  NANDN U43487 ( .A(n34513), .B(n34511), .Z(n34507) );
  IV U43488 ( .A(n34512), .Z(n34513) );
  XNOR U43489 ( .A(n34483), .B(n34514), .Z(n34478) );
  XNOR U43490 ( .A(n34481), .B(n34484), .Z(n34514) );
  NAND U43491 ( .A(n34515), .B(n34516), .Z(n34484) );
  NAND U43492 ( .A(n34517), .B(n34518), .Z(n34516) );
  OR U43493 ( .A(n34519), .B(n34520), .Z(n34517) );
  NANDN U43494 ( .A(n34521), .B(n34519), .Z(n34515) );
  IV U43495 ( .A(n34520), .Z(n34521) );
  NAND U43496 ( .A(n34522), .B(n34523), .Z(n34481) );
  NAND U43497 ( .A(n34524), .B(n34525), .Z(n34523) );
  NANDN U43498 ( .A(n34526), .B(n34527), .Z(n34524) );
  NANDN U43499 ( .A(n34527), .B(n34526), .Z(n34522) );
  AND U43500 ( .A(n34528), .B(n34529), .Z(n34483) );
  NAND U43501 ( .A(n34530), .B(n34531), .Z(n34529) );
  OR U43502 ( .A(n34532), .B(n34533), .Z(n34530) );
  NANDN U43503 ( .A(n34534), .B(n34532), .Z(n34528) );
  XNOR U43504 ( .A(n34509), .B(n34535), .Z(N62335) );
  XOR U43505 ( .A(n34511), .B(n34512), .Z(n34535) );
  XNOR U43506 ( .A(n34525), .B(n34536), .Z(n34512) );
  XOR U43507 ( .A(n34526), .B(n34527), .Z(n34536) );
  XOR U43508 ( .A(n34532), .B(n34537), .Z(n34527) );
  XOR U43509 ( .A(n34531), .B(n34534), .Z(n34537) );
  IV U43510 ( .A(n34533), .Z(n34534) );
  NAND U43511 ( .A(n34538), .B(n34539), .Z(n34533) );
  OR U43512 ( .A(n34540), .B(n34541), .Z(n34539) );
  OR U43513 ( .A(n34542), .B(n34543), .Z(n34538) );
  NAND U43514 ( .A(n34544), .B(n34545), .Z(n34531) );
  OR U43515 ( .A(n34546), .B(n34547), .Z(n34545) );
  OR U43516 ( .A(n34548), .B(n34549), .Z(n34544) );
  NOR U43517 ( .A(n34550), .B(n34551), .Z(n34532) );
  ANDN U43518 ( .B(n34552), .A(n34553), .Z(n34526) );
  XNOR U43519 ( .A(n34519), .B(n34554), .Z(n34525) );
  XNOR U43520 ( .A(n34518), .B(n34520), .Z(n34554) );
  NAND U43521 ( .A(n34555), .B(n34556), .Z(n34520) );
  OR U43522 ( .A(n34557), .B(n34558), .Z(n34556) );
  OR U43523 ( .A(n34559), .B(n34560), .Z(n34555) );
  NAND U43524 ( .A(n34561), .B(n34562), .Z(n34518) );
  OR U43525 ( .A(n34563), .B(n34564), .Z(n34562) );
  OR U43526 ( .A(n34565), .B(n34566), .Z(n34561) );
  ANDN U43527 ( .B(n34567), .A(n34568), .Z(n34519) );
  IV U43528 ( .A(n34569), .Z(n34567) );
  ANDN U43529 ( .B(n34570), .A(n34571), .Z(n34511) );
  XOR U43530 ( .A(n34497), .B(n34572), .Z(n34509) );
  XOR U43531 ( .A(n34498), .B(n34499), .Z(n34572) );
  XOR U43532 ( .A(n34504), .B(n34573), .Z(n34499) );
  XOR U43533 ( .A(n34503), .B(n34506), .Z(n34573) );
  IV U43534 ( .A(n34505), .Z(n34506) );
  NAND U43535 ( .A(n34574), .B(n34575), .Z(n34505) );
  OR U43536 ( .A(n34576), .B(n34577), .Z(n34575) );
  OR U43537 ( .A(n34578), .B(n34579), .Z(n34574) );
  NAND U43538 ( .A(n34580), .B(n34581), .Z(n34503) );
  OR U43539 ( .A(n34582), .B(n34583), .Z(n34581) );
  OR U43540 ( .A(n34584), .B(n34585), .Z(n34580) );
  NOR U43541 ( .A(n34586), .B(n34587), .Z(n34504) );
  ANDN U43542 ( .B(n34588), .A(n34589), .Z(n34498) );
  IV U43543 ( .A(n34590), .Z(n34588) );
  XNOR U43544 ( .A(n34491), .B(n34591), .Z(n34497) );
  XNOR U43545 ( .A(n34490), .B(n34492), .Z(n34591) );
  NAND U43546 ( .A(n34592), .B(n34593), .Z(n34492) );
  OR U43547 ( .A(n34594), .B(n34595), .Z(n34593) );
  OR U43548 ( .A(n34596), .B(n34597), .Z(n34592) );
  NAND U43549 ( .A(n34598), .B(n34599), .Z(n34490) );
  OR U43550 ( .A(n34600), .B(n34601), .Z(n34599) );
  OR U43551 ( .A(n34602), .B(n34603), .Z(n34598) );
  ANDN U43552 ( .B(n34604), .A(n34605), .Z(n34491) );
  IV U43553 ( .A(n34606), .Z(n34604) );
  XNOR U43554 ( .A(n34571), .B(n34570), .Z(N62334) );
  XOR U43555 ( .A(n34590), .B(n34589), .Z(n34570) );
  XNOR U43556 ( .A(n34605), .B(n34606), .Z(n34589) );
  XNOR U43557 ( .A(n34600), .B(n34601), .Z(n34606) );
  XNOR U43558 ( .A(n34602), .B(n34603), .Z(n34601) );
  XNOR U43559 ( .A(y[3229]), .B(x[3229]), .Z(n34603) );
  XNOR U43560 ( .A(y[3230]), .B(x[3230]), .Z(n34602) );
  XNOR U43561 ( .A(y[3228]), .B(x[3228]), .Z(n34600) );
  XNOR U43562 ( .A(n34594), .B(n34595), .Z(n34605) );
  XNOR U43563 ( .A(y[3225]), .B(x[3225]), .Z(n34595) );
  XNOR U43564 ( .A(n34596), .B(n34597), .Z(n34594) );
  XNOR U43565 ( .A(y[3226]), .B(x[3226]), .Z(n34597) );
  XNOR U43566 ( .A(y[3227]), .B(x[3227]), .Z(n34596) );
  XNOR U43567 ( .A(n34587), .B(n34586), .Z(n34590) );
  XNOR U43568 ( .A(n34582), .B(n34583), .Z(n34586) );
  XNOR U43569 ( .A(y[3222]), .B(x[3222]), .Z(n34583) );
  XNOR U43570 ( .A(n34584), .B(n34585), .Z(n34582) );
  XNOR U43571 ( .A(y[3223]), .B(x[3223]), .Z(n34585) );
  XNOR U43572 ( .A(y[3224]), .B(x[3224]), .Z(n34584) );
  XNOR U43573 ( .A(n34576), .B(n34577), .Z(n34587) );
  XNOR U43574 ( .A(y[3219]), .B(x[3219]), .Z(n34577) );
  XNOR U43575 ( .A(n34578), .B(n34579), .Z(n34576) );
  XNOR U43576 ( .A(y[3220]), .B(x[3220]), .Z(n34579) );
  XNOR U43577 ( .A(y[3221]), .B(x[3221]), .Z(n34578) );
  XOR U43578 ( .A(n34552), .B(n34553), .Z(n34571) );
  XNOR U43579 ( .A(n34568), .B(n34569), .Z(n34553) );
  XNOR U43580 ( .A(n34563), .B(n34564), .Z(n34569) );
  XNOR U43581 ( .A(n34565), .B(n34566), .Z(n34564) );
  XNOR U43582 ( .A(y[3217]), .B(x[3217]), .Z(n34566) );
  XNOR U43583 ( .A(y[3218]), .B(x[3218]), .Z(n34565) );
  XNOR U43584 ( .A(y[3216]), .B(x[3216]), .Z(n34563) );
  XNOR U43585 ( .A(n34557), .B(n34558), .Z(n34568) );
  XNOR U43586 ( .A(y[3213]), .B(x[3213]), .Z(n34558) );
  XNOR U43587 ( .A(n34559), .B(n34560), .Z(n34557) );
  XNOR U43588 ( .A(y[3214]), .B(x[3214]), .Z(n34560) );
  XNOR U43589 ( .A(y[3215]), .B(x[3215]), .Z(n34559) );
  XOR U43590 ( .A(n34551), .B(n34550), .Z(n34552) );
  XNOR U43591 ( .A(n34546), .B(n34547), .Z(n34550) );
  XNOR U43592 ( .A(y[3210]), .B(x[3210]), .Z(n34547) );
  XNOR U43593 ( .A(n34548), .B(n34549), .Z(n34546) );
  XNOR U43594 ( .A(y[3211]), .B(x[3211]), .Z(n34549) );
  XNOR U43595 ( .A(y[3212]), .B(x[3212]), .Z(n34548) );
  XNOR U43596 ( .A(n34540), .B(n34541), .Z(n34551) );
  XNOR U43597 ( .A(y[3207]), .B(x[3207]), .Z(n34541) );
  XNOR U43598 ( .A(n34542), .B(n34543), .Z(n34540) );
  XNOR U43599 ( .A(y[3208]), .B(x[3208]), .Z(n34543) );
  XNOR U43600 ( .A(y[3209]), .B(x[3209]), .Z(n34542) );
  NAND U43601 ( .A(n34607), .B(n34608), .Z(N62325) );
  NANDN U43602 ( .A(n34609), .B(n34610), .Z(n34608) );
  OR U43603 ( .A(n34611), .B(n34612), .Z(n34610) );
  NAND U43604 ( .A(n34611), .B(n34612), .Z(n34607) );
  XOR U43605 ( .A(n34611), .B(n34613), .Z(N62324) );
  XNOR U43606 ( .A(n34609), .B(n34612), .Z(n34613) );
  AND U43607 ( .A(n34614), .B(n34615), .Z(n34612) );
  NANDN U43608 ( .A(n34616), .B(n34617), .Z(n34615) );
  NANDN U43609 ( .A(n34618), .B(n34619), .Z(n34617) );
  NANDN U43610 ( .A(n34619), .B(n34618), .Z(n34614) );
  NAND U43611 ( .A(n34620), .B(n34621), .Z(n34609) );
  NANDN U43612 ( .A(n34622), .B(n34623), .Z(n34621) );
  OR U43613 ( .A(n34624), .B(n34625), .Z(n34623) );
  NAND U43614 ( .A(n34625), .B(n34624), .Z(n34620) );
  AND U43615 ( .A(n34626), .B(n34627), .Z(n34611) );
  NANDN U43616 ( .A(n34628), .B(n34629), .Z(n34627) );
  NANDN U43617 ( .A(n34630), .B(n34631), .Z(n34629) );
  NANDN U43618 ( .A(n34631), .B(n34630), .Z(n34626) );
  XOR U43619 ( .A(n34625), .B(n34632), .Z(N62323) );
  XOR U43620 ( .A(n34622), .B(n34624), .Z(n34632) );
  XNOR U43621 ( .A(n34618), .B(n34633), .Z(n34624) );
  XNOR U43622 ( .A(n34616), .B(n34619), .Z(n34633) );
  NAND U43623 ( .A(n34634), .B(n34635), .Z(n34619) );
  NAND U43624 ( .A(n34636), .B(n34637), .Z(n34635) );
  OR U43625 ( .A(n34638), .B(n34639), .Z(n34636) );
  NANDN U43626 ( .A(n34640), .B(n34638), .Z(n34634) );
  IV U43627 ( .A(n34639), .Z(n34640) );
  NAND U43628 ( .A(n34641), .B(n34642), .Z(n34616) );
  NAND U43629 ( .A(n34643), .B(n34644), .Z(n34642) );
  NANDN U43630 ( .A(n34645), .B(n34646), .Z(n34643) );
  NANDN U43631 ( .A(n34646), .B(n34645), .Z(n34641) );
  AND U43632 ( .A(n34647), .B(n34648), .Z(n34618) );
  NAND U43633 ( .A(n34649), .B(n34650), .Z(n34648) );
  OR U43634 ( .A(n34651), .B(n34652), .Z(n34649) );
  NANDN U43635 ( .A(n34653), .B(n34651), .Z(n34647) );
  NAND U43636 ( .A(n34654), .B(n34655), .Z(n34622) );
  NANDN U43637 ( .A(n34656), .B(n34657), .Z(n34655) );
  OR U43638 ( .A(n34658), .B(n34659), .Z(n34657) );
  NANDN U43639 ( .A(n34660), .B(n34658), .Z(n34654) );
  IV U43640 ( .A(n34659), .Z(n34660) );
  XNOR U43641 ( .A(n34630), .B(n34661), .Z(n34625) );
  XNOR U43642 ( .A(n34628), .B(n34631), .Z(n34661) );
  NAND U43643 ( .A(n34662), .B(n34663), .Z(n34631) );
  NAND U43644 ( .A(n34664), .B(n34665), .Z(n34663) );
  OR U43645 ( .A(n34666), .B(n34667), .Z(n34664) );
  NANDN U43646 ( .A(n34668), .B(n34666), .Z(n34662) );
  IV U43647 ( .A(n34667), .Z(n34668) );
  NAND U43648 ( .A(n34669), .B(n34670), .Z(n34628) );
  NAND U43649 ( .A(n34671), .B(n34672), .Z(n34670) );
  NANDN U43650 ( .A(n34673), .B(n34674), .Z(n34671) );
  NANDN U43651 ( .A(n34674), .B(n34673), .Z(n34669) );
  AND U43652 ( .A(n34675), .B(n34676), .Z(n34630) );
  NAND U43653 ( .A(n34677), .B(n34678), .Z(n34676) );
  OR U43654 ( .A(n34679), .B(n34680), .Z(n34677) );
  NANDN U43655 ( .A(n34681), .B(n34679), .Z(n34675) );
  XNOR U43656 ( .A(n34656), .B(n34682), .Z(N62322) );
  XOR U43657 ( .A(n34658), .B(n34659), .Z(n34682) );
  XNOR U43658 ( .A(n34672), .B(n34683), .Z(n34659) );
  XOR U43659 ( .A(n34673), .B(n34674), .Z(n34683) );
  XOR U43660 ( .A(n34679), .B(n34684), .Z(n34674) );
  XOR U43661 ( .A(n34678), .B(n34681), .Z(n34684) );
  IV U43662 ( .A(n34680), .Z(n34681) );
  NAND U43663 ( .A(n34685), .B(n34686), .Z(n34680) );
  OR U43664 ( .A(n34687), .B(n34688), .Z(n34686) );
  OR U43665 ( .A(n34689), .B(n34690), .Z(n34685) );
  NAND U43666 ( .A(n34691), .B(n34692), .Z(n34678) );
  OR U43667 ( .A(n34693), .B(n34694), .Z(n34692) );
  OR U43668 ( .A(n34695), .B(n34696), .Z(n34691) );
  NOR U43669 ( .A(n34697), .B(n34698), .Z(n34679) );
  ANDN U43670 ( .B(n34699), .A(n34700), .Z(n34673) );
  XNOR U43671 ( .A(n34666), .B(n34701), .Z(n34672) );
  XNOR U43672 ( .A(n34665), .B(n34667), .Z(n34701) );
  NAND U43673 ( .A(n34702), .B(n34703), .Z(n34667) );
  OR U43674 ( .A(n34704), .B(n34705), .Z(n34703) );
  OR U43675 ( .A(n34706), .B(n34707), .Z(n34702) );
  NAND U43676 ( .A(n34708), .B(n34709), .Z(n34665) );
  OR U43677 ( .A(n34710), .B(n34711), .Z(n34709) );
  OR U43678 ( .A(n34712), .B(n34713), .Z(n34708) );
  ANDN U43679 ( .B(n34714), .A(n34715), .Z(n34666) );
  IV U43680 ( .A(n34716), .Z(n34714) );
  ANDN U43681 ( .B(n34717), .A(n34718), .Z(n34658) );
  XOR U43682 ( .A(n34644), .B(n34719), .Z(n34656) );
  XOR U43683 ( .A(n34645), .B(n34646), .Z(n34719) );
  XOR U43684 ( .A(n34651), .B(n34720), .Z(n34646) );
  XOR U43685 ( .A(n34650), .B(n34653), .Z(n34720) );
  IV U43686 ( .A(n34652), .Z(n34653) );
  NAND U43687 ( .A(n34721), .B(n34722), .Z(n34652) );
  OR U43688 ( .A(n34723), .B(n34724), .Z(n34722) );
  OR U43689 ( .A(n34725), .B(n34726), .Z(n34721) );
  NAND U43690 ( .A(n34727), .B(n34728), .Z(n34650) );
  OR U43691 ( .A(n34729), .B(n34730), .Z(n34728) );
  OR U43692 ( .A(n34731), .B(n34732), .Z(n34727) );
  NOR U43693 ( .A(n34733), .B(n34734), .Z(n34651) );
  ANDN U43694 ( .B(n34735), .A(n34736), .Z(n34645) );
  IV U43695 ( .A(n34737), .Z(n34735) );
  XNOR U43696 ( .A(n34638), .B(n34738), .Z(n34644) );
  XNOR U43697 ( .A(n34637), .B(n34639), .Z(n34738) );
  NAND U43698 ( .A(n34739), .B(n34740), .Z(n34639) );
  OR U43699 ( .A(n34741), .B(n34742), .Z(n34740) );
  OR U43700 ( .A(n34743), .B(n34744), .Z(n34739) );
  NAND U43701 ( .A(n34745), .B(n34746), .Z(n34637) );
  OR U43702 ( .A(n34747), .B(n34748), .Z(n34746) );
  OR U43703 ( .A(n34749), .B(n34750), .Z(n34745) );
  ANDN U43704 ( .B(n34751), .A(n34752), .Z(n34638) );
  IV U43705 ( .A(n34753), .Z(n34751) );
  XNOR U43706 ( .A(n34718), .B(n34717), .Z(N62321) );
  XOR U43707 ( .A(n34737), .B(n34736), .Z(n34717) );
  XNOR U43708 ( .A(n34752), .B(n34753), .Z(n34736) );
  XNOR U43709 ( .A(n34747), .B(n34748), .Z(n34753) );
  XNOR U43710 ( .A(n34749), .B(n34750), .Z(n34748) );
  XNOR U43711 ( .A(y[3205]), .B(x[3205]), .Z(n34750) );
  XNOR U43712 ( .A(y[3206]), .B(x[3206]), .Z(n34749) );
  XNOR U43713 ( .A(y[3204]), .B(x[3204]), .Z(n34747) );
  XNOR U43714 ( .A(n34741), .B(n34742), .Z(n34752) );
  XNOR U43715 ( .A(y[3201]), .B(x[3201]), .Z(n34742) );
  XNOR U43716 ( .A(n34743), .B(n34744), .Z(n34741) );
  XNOR U43717 ( .A(y[3202]), .B(x[3202]), .Z(n34744) );
  XNOR U43718 ( .A(y[3203]), .B(x[3203]), .Z(n34743) );
  XNOR U43719 ( .A(n34734), .B(n34733), .Z(n34737) );
  XNOR U43720 ( .A(n34729), .B(n34730), .Z(n34733) );
  XNOR U43721 ( .A(y[3198]), .B(x[3198]), .Z(n34730) );
  XNOR U43722 ( .A(n34731), .B(n34732), .Z(n34729) );
  XNOR U43723 ( .A(y[3199]), .B(x[3199]), .Z(n34732) );
  XNOR U43724 ( .A(y[3200]), .B(x[3200]), .Z(n34731) );
  XNOR U43725 ( .A(n34723), .B(n34724), .Z(n34734) );
  XNOR U43726 ( .A(y[3195]), .B(x[3195]), .Z(n34724) );
  XNOR U43727 ( .A(n34725), .B(n34726), .Z(n34723) );
  XNOR U43728 ( .A(y[3196]), .B(x[3196]), .Z(n34726) );
  XNOR U43729 ( .A(y[3197]), .B(x[3197]), .Z(n34725) );
  XOR U43730 ( .A(n34699), .B(n34700), .Z(n34718) );
  XNOR U43731 ( .A(n34715), .B(n34716), .Z(n34700) );
  XNOR U43732 ( .A(n34710), .B(n34711), .Z(n34716) );
  XNOR U43733 ( .A(n34712), .B(n34713), .Z(n34711) );
  XNOR U43734 ( .A(y[3193]), .B(x[3193]), .Z(n34713) );
  XNOR U43735 ( .A(y[3194]), .B(x[3194]), .Z(n34712) );
  XNOR U43736 ( .A(y[3192]), .B(x[3192]), .Z(n34710) );
  XNOR U43737 ( .A(n34704), .B(n34705), .Z(n34715) );
  XNOR U43738 ( .A(y[3189]), .B(x[3189]), .Z(n34705) );
  XNOR U43739 ( .A(n34706), .B(n34707), .Z(n34704) );
  XNOR U43740 ( .A(y[3190]), .B(x[3190]), .Z(n34707) );
  XNOR U43741 ( .A(y[3191]), .B(x[3191]), .Z(n34706) );
  XOR U43742 ( .A(n34698), .B(n34697), .Z(n34699) );
  XNOR U43743 ( .A(n34693), .B(n34694), .Z(n34697) );
  XNOR U43744 ( .A(y[3186]), .B(x[3186]), .Z(n34694) );
  XNOR U43745 ( .A(n34695), .B(n34696), .Z(n34693) );
  XNOR U43746 ( .A(y[3187]), .B(x[3187]), .Z(n34696) );
  XNOR U43747 ( .A(y[3188]), .B(x[3188]), .Z(n34695) );
  XNOR U43748 ( .A(n34687), .B(n34688), .Z(n34698) );
  XNOR U43749 ( .A(y[3183]), .B(x[3183]), .Z(n34688) );
  XNOR U43750 ( .A(n34689), .B(n34690), .Z(n34687) );
  XNOR U43751 ( .A(y[3184]), .B(x[3184]), .Z(n34690) );
  XNOR U43752 ( .A(y[3185]), .B(x[3185]), .Z(n34689) );
  NAND U43753 ( .A(n34754), .B(n34755), .Z(N62312) );
  NANDN U43754 ( .A(n34756), .B(n34757), .Z(n34755) );
  OR U43755 ( .A(n34758), .B(n34759), .Z(n34757) );
  NAND U43756 ( .A(n34758), .B(n34759), .Z(n34754) );
  XOR U43757 ( .A(n34758), .B(n34760), .Z(N62311) );
  XNOR U43758 ( .A(n34756), .B(n34759), .Z(n34760) );
  AND U43759 ( .A(n34761), .B(n34762), .Z(n34759) );
  NANDN U43760 ( .A(n34763), .B(n34764), .Z(n34762) );
  NANDN U43761 ( .A(n34765), .B(n34766), .Z(n34764) );
  NANDN U43762 ( .A(n34766), .B(n34765), .Z(n34761) );
  NAND U43763 ( .A(n34767), .B(n34768), .Z(n34756) );
  NANDN U43764 ( .A(n34769), .B(n34770), .Z(n34768) );
  OR U43765 ( .A(n34771), .B(n34772), .Z(n34770) );
  NAND U43766 ( .A(n34772), .B(n34771), .Z(n34767) );
  AND U43767 ( .A(n34773), .B(n34774), .Z(n34758) );
  NANDN U43768 ( .A(n34775), .B(n34776), .Z(n34774) );
  NANDN U43769 ( .A(n34777), .B(n34778), .Z(n34776) );
  NANDN U43770 ( .A(n34778), .B(n34777), .Z(n34773) );
  XOR U43771 ( .A(n34772), .B(n34779), .Z(N62310) );
  XOR U43772 ( .A(n34769), .B(n34771), .Z(n34779) );
  XNOR U43773 ( .A(n34765), .B(n34780), .Z(n34771) );
  XNOR U43774 ( .A(n34763), .B(n34766), .Z(n34780) );
  NAND U43775 ( .A(n34781), .B(n34782), .Z(n34766) );
  NAND U43776 ( .A(n34783), .B(n34784), .Z(n34782) );
  OR U43777 ( .A(n34785), .B(n34786), .Z(n34783) );
  NANDN U43778 ( .A(n34787), .B(n34785), .Z(n34781) );
  IV U43779 ( .A(n34786), .Z(n34787) );
  NAND U43780 ( .A(n34788), .B(n34789), .Z(n34763) );
  NAND U43781 ( .A(n34790), .B(n34791), .Z(n34789) );
  NANDN U43782 ( .A(n34792), .B(n34793), .Z(n34790) );
  NANDN U43783 ( .A(n34793), .B(n34792), .Z(n34788) );
  AND U43784 ( .A(n34794), .B(n34795), .Z(n34765) );
  NAND U43785 ( .A(n34796), .B(n34797), .Z(n34795) );
  OR U43786 ( .A(n34798), .B(n34799), .Z(n34796) );
  NANDN U43787 ( .A(n34800), .B(n34798), .Z(n34794) );
  NAND U43788 ( .A(n34801), .B(n34802), .Z(n34769) );
  NANDN U43789 ( .A(n34803), .B(n34804), .Z(n34802) );
  OR U43790 ( .A(n34805), .B(n34806), .Z(n34804) );
  NANDN U43791 ( .A(n34807), .B(n34805), .Z(n34801) );
  IV U43792 ( .A(n34806), .Z(n34807) );
  XNOR U43793 ( .A(n34777), .B(n34808), .Z(n34772) );
  XNOR U43794 ( .A(n34775), .B(n34778), .Z(n34808) );
  NAND U43795 ( .A(n34809), .B(n34810), .Z(n34778) );
  NAND U43796 ( .A(n34811), .B(n34812), .Z(n34810) );
  OR U43797 ( .A(n34813), .B(n34814), .Z(n34811) );
  NANDN U43798 ( .A(n34815), .B(n34813), .Z(n34809) );
  IV U43799 ( .A(n34814), .Z(n34815) );
  NAND U43800 ( .A(n34816), .B(n34817), .Z(n34775) );
  NAND U43801 ( .A(n34818), .B(n34819), .Z(n34817) );
  NANDN U43802 ( .A(n34820), .B(n34821), .Z(n34818) );
  NANDN U43803 ( .A(n34821), .B(n34820), .Z(n34816) );
  AND U43804 ( .A(n34822), .B(n34823), .Z(n34777) );
  NAND U43805 ( .A(n34824), .B(n34825), .Z(n34823) );
  OR U43806 ( .A(n34826), .B(n34827), .Z(n34824) );
  NANDN U43807 ( .A(n34828), .B(n34826), .Z(n34822) );
  XNOR U43808 ( .A(n34803), .B(n34829), .Z(N62309) );
  XOR U43809 ( .A(n34805), .B(n34806), .Z(n34829) );
  XNOR U43810 ( .A(n34819), .B(n34830), .Z(n34806) );
  XOR U43811 ( .A(n34820), .B(n34821), .Z(n34830) );
  XOR U43812 ( .A(n34826), .B(n34831), .Z(n34821) );
  XOR U43813 ( .A(n34825), .B(n34828), .Z(n34831) );
  IV U43814 ( .A(n34827), .Z(n34828) );
  NAND U43815 ( .A(n34832), .B(n34833), .Z(n34827) );
  OR U43816 ( .A(n34834), .B(n34835), .Z(n34833) );
  OR U43817 ( .A(n34836), .B(n34837), .Z(n34832) );
  NAND U43818 ( .A(n34838), .B(n34839), .Z(n34825) );
  OR U43819 ( .A(n34840), .B(n34841), .Z(n34839) );
  OR U43820 ( .A(n34842), .B(n34843), .Z(n34838) );
  NOR U43821 ( .A(n34844), .B(n34845), .Z(n34826) );
  ANDN U43822 ( .B(n34846), .A(n34847), .Z(n34820) );
  XNOR U43823 ( .A(n34813), .B(n34848), .Z(n34819) );
  XNOR U43824 ( .A(n34812), .B(n34814), .Z(n34848) );
  NAND U43825 ( .A(n34849), .B(n34850), .Z(n34814) );
  OR U43826 ( .A(n34851), .B(n34852), .Z(n34850) );
  OR U43827 ( .A(n34853), .B(n34854), .Z(n34849) );
  NAND U43828 ( .A(n34855), .B(n34856), .Z(n34812) );
  OR U43829 ( .A(n34857), .B(n34858), .Z(n34856) );
  OR U43830 ( .A(n34859), .B(n34860), .Z(n34855) );
  ANDN U43831 ( .B(n34861), .A(n34862), .Z(n34813) );
  IV U43832 ( .A(n34863), .Z(n34861) );
  ANDN U43833 ( .B(n34864), .A(n34865), .Z(n34805) );
  XOR U43834 ( .A(n34791), .B(n34866), .Z(n34803) );
  XOR U43835 ( .A(n34792), .B(n34793), .Z(n34866) );
  XOR U43836 ( .A(n34798), .B(n34867), .Z(n34793) );
  XOR U43837 ( .A(n34797), .B(n34800), .Z(n34867) );
  IV U43838 ( .A(n34799), .Z(n34800) );
  NAND U43839 ( .A(n34868), .B(n34869), .Z(n34799) );
  OR U43840 ( .A(n34870), .B(n34871), .Z(n34869) );
  OR U43841 ( .A(n34872), .B(n34873), .Z(n34868) );
  NAND U43842 ( .A(n34874), .B(n34875), .Z(n34797) );
  OR U43843 ( .A(n34876), .B(n34877), .Z(n34875) );
  OR U43844 ( .A(n34878), .B(n34879), .Z(n34874) );
  NOR U43845 ( .A(n34880), .B(n34881), .Z(n34798) );
  ANDN U43846 ( .B(n34882), .A(n34883), .Z(n34792) );
  IV U43847 ( .A(n34884), .Z(n34882) );
  XNOR U43848 ( .A(n34785), .B(n34885), .Z(n34791) );
  XNOR U43849 ( .A(n34784), .B(n34786), .Z(n34885) );
  NAND U43850 ( .A(n34886), .B(n34887), .Z(n34786) );
  OR U43851 ( .A(n34888), .B(n34889), .Z(n34887) );
  OR U43852 ( .A(n34890), .B(n34891), .Z(n34886) );
  NAND U43853 ( .A(n34892), .B(n34893), .Z(n34784) );
  OR U43854 ( .A(n34894), .B(n34895), .Z(n34893) );
  OR U43855 ( .A(n34896), .B(n34897), .Z(n34892) );
  ANDN U43856 ( .B(n34898), .A(n34899), .Z(n34785) );
  IV U43857 ( .A(n34900), .Z(n34898) );
  XNOR U43858 ( .A(n34865), .B(n34864), .Z(N62308) );
  XOR U43859 ( .A(n34884), .B(n34883), .Z(n34864) );
  XNOR U43860 ( .A(n34899), .B(n34900), .Z(n34883) );
  XNOR U43861 ( .A(n34894), .B(n34895), .Z(n34900) );
  XNOR U43862 ( .A(n34896), .B(n34897), .Z(n34895) );
  XNOR U43863 ( .A(y[3181]), .B(x[3181]), .Z(n34897) );
  XNOR U43864 ( .A(y[3182]), .B(x[3182]), .Z(n34896) );
  XNOR U43865 ( .A(y[3180]), .B(x[3180]), .Z(n34894) );
  XNOR U43866 ( .A(n34888), .B(n34889), .Z(n34899) );
  XNOR U43867 ( .A(y[3177]), .B(x[3177]), .Z(n34889) );
  XNOR U43868 ( .A(n34890), .B(n34891), .Z(n34888) );
  XNOR U43869 ( .A(y[3178]), .B(x[3178]), .Z(n34891) );
  XNOR U43870 ( .A(y[3179]), .B(x[3179]), .Z(n34890) );
  XNOR U43871 ( .A(n34881), .B(n34880), .Z(n34884) );
  XNOR U43872 ( .A(n34876), .B(n34877), .Z(n34880) );
  XNOR U43873 ( .A(y[3174]), .B(x[3174]), .Z(n34877) );
  XNOR U43874 ( .A(n34878), .B(n34879), .Z(n34876) );
  XNOR U43875 ( .A(y[3175]), .B(x[3175]), .Z(n34879) );
  XNOR U43876 ( .A(y[3176]), .B(x[3176]), .Z(n34878) );
  XNOR U43877 ( .A(n34870), .B(n34871), .Z(n34881) );
  XNOR U43878 ( .A(y[3171]), .B(x[3171]), .Z(n34871) );
  XNOR U43879 ( .A(n34872), .B(n34873), .Z(n34870) );
  XNOR U43880 ( .A(y[3172]), .B(x[3172]), .Z(n34873) );
  XNOR U43881 ( .A(y[3173]), .B(x[3173]), .Z(n34872) );
  XOR U43882 ( .A(n34846), .B(n34847), .Z(n34865) );
  XNOR U43883 ( .A(n34862), .B(n34863), .Z(n34847) );
  XNOR U43884 ( .A(n34857), .B(n34858), .Z(n34863) );
  XNOR U43885 ( .A(n34859), .B(n34860), .Z(n34858) );
  XNOR U43886 ( .A(y[3169]), .B(x[3169]), .Z(n34860) );
  XNOR U43887 ( .A(y[3170]), .B(x[3170]), .Z(n34859) );
  XNOR U43888 ( .A(y[3168]), .B(x[3168]), .Z(n34857) );
  XNOR U43889 ( .A(n34851), .B(n34852), .Z(n34862) );
  XNOR U43890 ( .A(y[3165]), .B(x[3165]), .Z(n34852) );
  XNOR U43891 ( .A(n34853), .B(n34854), .Z(n34851) );
  XNOR U43892 ( .A(y[3166]), .B(x[3166]), .Z(n34854) );
  XNOR U43893 ( .A(y[3167]), .B(x[3167]), .Z(n34853) );
  XOR U43894 ( .A(n34845), .B(n34844), .Z(n34846) );
  XNOR U43895 ( .A(n34840), .B(n34841), .Z(n34844) );
  XNOR U43896 ( .A(y[3162]), .B(x[3162]), .Z(n34841) );
  XNOR U43897 ( .A(n34842), .B(n34843), .Z(n34840) );
  XNOR U43898 ( .A(y[3163]), .B(x[3163]), .Z(n34843) );
  XNOR U43899 ( .A(y[3164]), .B(x[3164]), .Z(n34842) );
  XNOR U43900 ( .A(n34834), .B(n34835), .Z(n34845) );
  XNOR U43901 ( .A(y[3159]), .B(x[3159]), .Z(n34835) );
  XNOR U43902 ( .A(n34836), .B(n34837), .Z(n34834) );
  XNOR U43903 ( .A(y[3160]), .B(x[3160]), .Z(n34837) );
  XNOR U43904 ( .A(y[3161]), .B(x[3161]), .Z(n34836) );
  NAND U43905 ( .A(n34901), .B(n34902), .Z(N62299) );
  NANDN U43906 ( .A(n34903), .B(n34904), .Z(n34902) );
  OR U43907 ( .A(n34905), .B(n34906), .Z(n34904) );
  NAND U43908 ( .A(n34905), .B(n34906), .Z(n34901) );
  XOR U43909 ( .A(n34905), .B(n34907), .Z(N62298) );
  XNOR U43910 ( .A(n34903), .B(n34906), .Z(n34907) );
  AND U43911 ( .A(n34908), .B(n34909), .Z(n34906) );
  NANDN U43912 ( .A(n34910), .B(n34911), .Z(n34909) );
  NANDN U43913 ( .A(n34912), .B(n34913), .Z(n34911) );
  NANDN U43914 ( .A(n34913), .B(n34912), .Z(n34908) );
  NAND U43915 ( .A(n34914), .B(n34915), .Z(n34903) );
  NANDN U43916 ( .A(n34916), .B(n34917), .Z(n34915) );
  OR U43917 ( .A(n34918), .B(n34919), .Z(n34917) );
  NAND U43918 ( .A(n34919), .B(n34918), .Z(n34914) );
  AND U43919 ( .A(n34920), .B(n34921), .Z(n34905) );
  NANDN U43920 ( .A(n34922), .B(n34923), .Z(n34921) );
  NANDN U43921 ( .A(n34924), .B(n34925), .Z(n34923) );
  NANDN U43922 ( .A(n34925), .B(n34924), .Z(n34920) );
  XOR U43923 ( .A(n34919), .B(n34926), .Z(N62297) );
  XOR U43924 ( .A(n34916), .B(n34918), .Z(n34926) );
  XNOR U43925 ( .A(n34912), .B(n34927), .Z(n34918) );
  XNOR U43926 ( .A(n34910), .B(n34913), .Z(n34927) );
  NAND U43927 ( .A(n34928), .B(n34929), .Z(n34913) );
  NAND U43928 ( .A(n34930), .B(n34931), .Z(n34929) );
  OR U43929 ( .A(n34932), .B(n34933), .Z(n34930) );
  NANDN U43930 ( .A(n34934), .B(n34932), .Z(n34928) );
  IV U43931 ( .A(n34933), .Z(n34934) );
  NAND U43932 ( .A(n34935), .B(n34936), .Z(n34910) );
  NAND U43933 ( .A(n34937), .B(n34938), .Z(n34936) );
  NANDN U43934 ( .A(n34939), .B(n34940), .Z(n34937) );
  NANDN U43935 ( .A(n34940), .B(n34939), .Z(n34935) );
  AND U43936 ( .A(n34941), .B(n34942), .Z(n34912) );
  NAND U43937 ( .A(n34943), .B(n34944), .Z(n34942) );
  OR U43938 ( .A(n34945), .B(n34946), .Z(n34943) );
  NANDN U43939 ( .A(n34947), .B(n34945), .Z(n34941) );
  NAND U43940 ( .A(n34948), .B(n34949), .Z(n34916) );
  NANDN U43941 ( .A(n34950), .B(n34951), .Z(n34949) );
  OR U43942 ( .A(n34952), .B(n34953), .Z(n34951) );
  NANDN U43943 ( .A(n34954), .B(n34952), .Z(n34948) );
  IV U43944 ( .A(n34953), .Z(n34954) );
  XNOR U43945 ( .A(n34924), .B(n34955), .Z(n34919) );
  XNOR U43946 ( .A(n34922), .B(n34925), .Z(n34955) );
  NAND U43947 ( .A(n34956), .B(n34957), .Z(n34925) );
  NAND U43948 ( .A(n34958), .B(n34959), .Z(n34957) );
  OR U43949 ( .A(n34960), .B(n34961), .Z(n34958) );
  NANDN U43950 ( .A(n34962), .B(n34960), .Z(n34956) );
  IV U43951 ( .A(n34961), .Z(n34962) );
  NAND U43952 ( .A(n34963), .B(n34964), .Z(n34922) );
  NAND U43953 ( .A(n34965), .B(n34966), .Z(n34964) );
  NANDN U43954 ( .A(n34967), .B(n34968), .Z(n34965) );
  NANDN U43955 ( .A(n34968), .B(n34967), .Z(n34963) );
  AND U43956 ( .A(n34969), .B(n34970), .Z(n34924) );
  NAND U43957 ( .A(n34971), .B(n34972), .Z(n34970) );
  OR U43958 ( .A(n34973), .B(n34974), .Z(n34971) );
  NANDN U43959 ( .A(n34975), .B(n34973), .Z(n34969) );
  XNOR U43960 ( .A(n34950), .B(n34976), .Z(N62296) );
  XOR U43961 ( .A(n34952), .B(n34953), .Z(n34976) );
  XNOR U43962 ( .A(n34966), .B(n34977), .Z(n34953) );
  XOR U43963 ( .A(n34967), .B(n34968), .Z(n34977) );
  XOR U43964 ( .A(n34973), .B(n34978), .Z(n34968) );
  XOR U43965 ( .A(n34972), .B(n34975), .Z(n34978) );
  IV U43966 ( .A(n34974), .Z(n34975) );
  NAND U43967 ( .A(n34979), .B(n34980), .Z(n34974) );
  OR U43968 ( .A(n34981), .B(n34982), .Z(n34980) );
  OR U43969 ( .A(n34983), .B(n34984), .Z(n34979) );
  NAND U43970 ( .A(n34985), .B(n34986), .Z(n34972) );
  OR U43971 ( .A(n34987), .B(n34988), .Z(n34986) );
  OR U43972 ( .A(n34989), .B(n34990), .Z(n34985) );
  NOR U43973 ( .A(n34991), .B(n34992), .Z(n34973) );
  ANDN U43974 ( .B(n34993), .A(n34994), .Z(n34967) );
  XNOR U43975 ( .A(n34960), .B(n34995), .Z(n34966) );
  XNOR U43976 ( .A(n34959), .B(n34961), .Z(n34995) );
  NAND U43977 ( .A(n34996), .B(n34997), .Z(n34961) );
  OR U43978 ( .A(n34998), .B(n34999), .Z(n34997) );
  OR U43979 ( .A(n35000), .B(n35001), .Z(n34996) );
  NAND U43980 ( .A(n35002), .B(n35003), .Z(n34959) );
  OR U43981 ( .A(n35004), .B(n35005), .Z(n35003) );
  OR U43982 ( .A(n35006), .B(n35007), .Z(n35002) );
  ANDN U43983 ( .B(n35008), .A(n35009), .Z(n34960) );
  IV U43984 ( .A(n35010), .Z(n35008) );
  ANDN U43985 ( .B(n35011), .A(n35012), .Z(n34952) );
  XOR U43986 ( .A(n34938), .B(n35013), .Z(n34950) );
  XOR U43987 ( .A(n34939), .B(n34940), .Z(n35013) );
  XOR U43988 ( .A(n34945), .B(n35014), .Z(n34940) );
  XOR U43989 ( .A(n34944), .B(n34947), .Z(n35014) );
  IV U43990 ( .A(n34946), .Z(n34947) );
  NAND U43991 ( .A(n35015), .B(n35016), .Z(n34946) );
  OR U43992 ( .A(n35017), .B(n35018), .Z(n35016) );
  OR U43993 ( .A(n35019), .B(n35020), .Z(n35015) );
  NAND U43994 ( .A(n35021), .B(n35022), .Z(n34944) );
  OR U43995 ( .A(n35023), .B(n35024), .Z(n35022) );
  OR U43996 ( .A(n35025), .B(n35026), .Z(n35021) );
  NOR U43997 ( .A(n35027), .B(n35028), .Z(n34945) );
  ANDN U43998 ( .B(n35029), .A(n35030), .Z(n34939) );
  IV U43999 ( .A(n35031), .Z(n35029) );
  XNOR U44000 ( .A(n34932), .B(n35032), .Z(n34938) );
  XNOR U44001 ( .A(n34931), .B(n34933), .Z(n35032) );
  NAND U44002 ( .A(n35033), .B(n35034), .Z(n34933) );
  OR U44003 ( .A(n35035), .B(n35036), .Z(n35034) );
  OR U44004 ( .A(n35037), .B(n35038), .Z(n35033) );
  NAND U44005 ( .A(n35039), .B(n35040), .Z(n34931) );
  OR U44006 ( .A(n35041), .B(n35042), .Z(n35040) );
  OR U44007 ( .A(n35043), .B(n35044), .Z(n35039) );
  ANDN U44008 ( .B(n35045), .A(n35046), .Z(n34932) );
  IV U44009 ( .A(n35047), .Z(n35045) );
  XNOR U44010 ( .A(n35012), .B(n35011), .Z(N62295) );
  XOR U44011 ( .A(n35031), .B(n35030), .Z(n35011) );
  XNOR U44012 ( .A(n35046), .B(n35047), .Z(n35030) );
  XNOR U44013 ( .A(n35041), .B(n35042), .Z(n35047) );
  XNOR U44014 ( .A(n35043), .B(n35044), .Z(n35042) );
  XNOR U44015 ( .A(y[3157]), .B(x[3157]), .Z(n35044) );
  XNOR U44016 ( .A(y[3158]), .B(x[3158]), .Z(n35043) );
  XNOR U44017 ( .A(y[3156]), .B(x[3156]), .Z(n35041) );
  XNOR U44018 ( .A(n35035), .B(n35036), .Z(n35046) );
  XNOR U44019 ( .A(y[3153]), .B(x[3153]), .Z(n35036) );
  XNOR U44020 ( .A(n35037), .B(n35038), .Z(n35035) );
  XNOR U44021 ( .A(y[3154]), .B(x[3154]), .Z(n35038) );
  XNOR U44022 ( .A(y[3155]), .B(x[3155]), .Z(n35037) );
  XNOR U44023 ( .A(n35028), .B(n35027), .Z(n35031) );
  XNOR U44024 ( .A(n35023), .B(n35024), .Z(n35027) );
  XNOR U44025 ( .A(y[3150]), .B(x[3150]), .Z(n35024) );
  XNOR U44026 ( .A(n35025), .B(n35026), .Z(n35023) );
  XNOR U44027 ( .A(y[3151]), .B(x[3151]), .Z(n35026) );
  XNOR U44028 ( .A(y[3152]), .B(x[3152]), .Z(n35025) );
  XNOR U44029 ( .A(n35017), .B(n35018), .Z(n35028) );
  XNOR U44030 ( .A(y[3147]), .B(x[3147]), .Z(n35018) );
  XNOR U44031 ( .A(n35019), .B(n35020), .Z(n35017) );
  XNOR U44032 ( .A(y[3148]), .B(x[3148]), .Z(n35020) );
  XNOR U44033 ( .A(y[3149]), .B(x[3149]), .Z(n35019) );
  XOR U44034 ( .A(n34993), .B(n34994), .Z(n35012) );
  XNOR U44035 ( .A(n35009), .B(n35010), .Z(n34994) );
  XNOR U44036 ( .A(n35004), .B(n35005), .Z(n35010) );
  XNOR U44037 ( .A(n35006), .B(n35007), .Z(n35005) );
  XNOR U44038 ( .A(y[3145]), .B(x[3145]), .Z(n35007) );
  XNOR U44039 ( .A(y[3146]), .B(x[3146]), .Z(n35006) );
  XNOR U44040 ( .A(y[3144]), .B(x[3144]), .Z(n35004) );
  XNOR U44041 ( .A(n34998), .B(n34999), .Z(n35009) );
  XNOR U44042 ( .A(y[3141]), .B(x[3141]), .Z(n34999) );
  XNOR U44043 ( .A(n35000), .B(n35001), .Z(n34998) );
  XNOR U44044 ( .A(y[3142]), .B(x[3142]), .Z(n35001) );
  XNOR U44045 ( .A(y[3143]), .B(x[3143]), .Z(n35000) );
  XOR U44046 ( .A(n34992), .B(n34991), .Z(n34993) );
  XNOR U44047 ( .A(n34987), .B(n34988), .Z(n34991) );
  XNOR U44048 ( .A(y[3138]), .B(x[3138]), .Z(n34988) );
  XNOR U44049 ( .A(n34989), .B(n34990), .Z(n34987) );
  XNOR U44050 ( .A(y[3139]), .B(x[3139]), .Z(n34990) );
  XNOR U44051 ( .A(y[3140]), .B(x[3140]), .Z(n34989) );
  XNOR U44052 ( .A(n34981), .B(n34982), .Z(n34992) );
  XNOR U44053 ( .A(y[3135]), .B(x[3135]), .Z(n34982) );
  XNOR U44054 ( .A(n34983), .B(n34984), .Z(n34981) );
  XNOR U44055 ( .A(y[3136]), .B(x[3136]), .Z(n34984) );
  XNOR U44056 ( .A(y[3137]), .B(x[3137]), .Z(n34983) );
  NAND U44057 ( .A(n35048), .B(n35049), .Z(N62286) );
  NANDN U44058 ( .A(n35050), .B(n35051), .Z(n35049) );
  OR U44059 ( .A(n35052), .B(n35053), .Z(n35051) );
  NAND U44060 ( .A(n35052), .B(n35053), .Z(n35048) );
  XOR U44061 ( .A(n35052), .B(n35054), .Z(N62285) );
  XNOR U44062 ( .A(n35050), .B(n35053), .Z(n35054) );
  AND U44063 ( .A(n35055), .B(n35056), .Z(n35053) );
  NANDN U44064 ( .A(n35057), .B(n35058), .Z(n35056) );
  NANDN U44065 ( .A(n35059), .B(n35060), .Z(n35058) );
  NANDN U44066 ( .A(n35060), .B(n35059), .Z(n35055) );
  NAND U44067 ( .A(n35061), .B(n35062), .Z(n35050) );
  NANDN U44068 ( .A(n35063), .B(n35064), .Z(n35062) );
  OR U44069 ( .A(n35065), .B(n35066), .Z(n35064) );
  NAND U44070 ( .A(n35066), .B(n35065), .Z(n35061) );
  AND U44071 ( .A(n35067), .B(n35068), .Z(n35052) );
  NANDN U44072 ( .A(n35069), .B(n35070), .Z(n35068) );
  NANDN U44073 ( .A(n35071), .B(n35072), .Z(n35070) );
  NANDN U44074 ( .A(n35072), .B(n35071), .Z(n35067) );
  XOR U44075 ( .A(n35066), .B(n35073), .Z(N62284) );
  XOR U44076 ( .A(n35063), .B(n35065), .Z(n35073) );
  XNOR U44077 ( .A(n35059), .B(n35074), .Z(n35065) );
  XNOR U44078 ( .A(n35057), .B(n35060), .Z(n35074) );
  NAND U44079 ( .A(n35075), .B(n35076), .Z(n35060) );
  NAND U44080 ( .A(n35077), .B(n35078), .Z(n35076) );
  OR U44081 ( .A(n35079), .B(n35080), .Z(n35077) );
  NANDN U44082 ( .A(n35081), .B(n35079), .Z(n35075) );
  IV U44083 ( .A(n35080), .Z(n35081) );
  NAND U44084 ( .A(n35082), .B(n35083), .Z(n35057) );
  NAND U44085 ( .A(n35084), .B(n35085), .Z(n35083) );
  NANDN U44086 ( .A(n35086), .B(n35087), .Z(n35084) );
  NANDN U44087 ( .A(n35087), .B(n35086), .Z(n35082) );
  AND U44088 ( .A(n35088), .B(n35089), .Z(n35059) );
  NAND U44089 ( .A(n35090), .B(n35091), .Z(n35089) );
  OR U44090 ( .A(n35092), .B(n35093), .Z(n35090) );
  NANDN U44091 ( .A(n35094), .B(n35092), .Z(n35088) );
  NAND U44092 ( .A(n35095), .B(n35096), .Z(n35063) );
  NANDN U44093 ( .A(n35097), .B(n35098), .Z(n35096) );
  OR U44094 ( .A(n35099), .B(n35100), .Z(n35098) );
  NANDN U44095 ( .A(n35101), .B(n35099), .Z(n35095) );
  IV U44096 ( .A(n35100), .Z(n35101) );
  XNOR U44097 ( .A(n35071), .B(n35102), .Z(n35066) );
  XNOR U44098 ( .A(n35069), .B(n35072), .Z(n35102) );
  NAND U44099 ( .A(n35103), .B(n35104), .Z(n35072) );
  NAND U44100 ( .A(n35105), .B(n35106), .Z(n35104) );
  OR U44101 ( .A(n35107), .B(n35108), .Z(n35105) );
  NANDN U44102 ( .A(n35109), .B(n35107), .Z(n35103) );
  IV U44103 ( .A(n35108), .Z(n35109) );
  NAND U44104 ( .A(n35110), .B(n35111), .Z(n35069) );
  NAND U44105 ( .A(n35112), .B(n35113), .Z(n35111) );
  NANDN U44106 ( .A(n35114), .B(n35115), .Z(n35112) );
  NANDN U44107 ( .A(n35115), .B(n35114), .Z(n35110) );
  AND U44108 ( .A(n35116), .B(n35117), .Z(n35071) );
  NAND U44109 ( .A(n35118), .B(n35119), .Z(n35117) );
  OR U44110 ( .A(n35120), .B(n35121), .Z(n35118) );
  NANDN U44111 ( .A(n35122), .B(n35120), .Z(n35116) );
  XNOR U44112 ( .A(n35097), .B(n35123), .Z(N62283) );
  XOR U44113 ( .A(n35099), .B(n35100), .Z(n35123) );
  XNOR U44114 ( .A(n35113), .B(n35124), .Z(n35100) );
  XOR U44115 ( .A(n35114), .B(n35115), .Z(n35124) );
  XOR U44116 ( .A(n35120), .B(n35125), .Z(n35115) );
  XOR U44117 ( .A(n35119), .B(n35122), .Z(n35125) );
  IV U44118 ( .A(n35121), .Z(n35122) );
  NAND U44119 ( .A(n35126), .B(n35127), .Z(n35121) );
  OR U44120 ( .A(n35128), .B(n35129), .Z(n35127) );
  OR U44121 ( .A(n35130), .B(n35131), .Z(n35126) );
  NAND U44122 ( .A(n35132), .B(n35133), .Z(n35119) );
  OR U44123 ( .A(n35134), .B(n35135), .Z(n35133) );
  OR U44124 ( .A(n35136), .B(n35137), .Z(n35132) );
  NOR U44125 ( .A(n35138), .B(n35139), .Z(n35120) );
  ANDN U44126 ( .B(n35140), .A(n35141), .Z(n35114) );
  XNOR U44127 ( .A(n35107), .B(n35142), .Z(n35113) );
  XNOR U44128 ( .A(n35106), .B(n35108), .Z(n35142) );
  NAND U44129 ( .A(n35143), .B(n35144), .Z(n35108) );
  OR U44130 ( .A(n35145), .B(n35146), .Z(n35144) );
  OR U44131 ( .A(n35147), .B(n35148), .Z(n35143) );
  NAND U44132 ( .A(n35149), .B(n35150), .Z(n35106) );
  OR U44133 ( .A(n35151), .B(n35152), .Z(n35150) );
  OR U44134 ( .A(n35153), .B(n35154), .Z(n35149) );
  ANDN U44135 ( .B(n35155), .A(n35156), .Z(n35107) );
  IV U44136 ( .A(n35157), .Z(n35155) );
  ANDN U44137 ( .B(n35158), .A(n35159), .Z(n35099) );
  XOR U44138 ( .A(n35085), .B(n35160), .Z(n35097) );
  XOR U44139 ( .A(n35086), .B(n35087), .Z(n35160) );
  XOR U44140 ( .A(n35092), .B(n35161), .Z(n35087) );
  XOR U44141 ( .A(n35091), .B(n35094), .Z(n35161) );
  IV U44142 ( .A(n35093), .Z(n35094) );
  NAND U44143 ( .A(n35162), .B(n35163), .Z(n35093) );
  OR U44144 ( .A(n35164), .B(n35165), .Z(n35163) );
  OR U44145 ( .A(n35166), .B(n35167), .Z(n35162) );
  NAND U44146 ( .A(n35168), .B(n35169), .Z(n35091) );
  OR U44147 ( .A(n35170), .B(n35171), .Z(n35169) );
  OR U44148 ( .A(n35172), .B(n35173), .Z(n35168) );
  NOR U44149 ( .A(n35174), .B(n35175), .Z(n35092) );
  ANDN U44150 ( .B(n35176), .A(n35177), .Z(n35086) );
  IV U44151 ( .A(n35178), .Z(n35176) );
  XNOR U44152 ( .A(n35079), .B(n35179), .Z(n35085) );
  XNOR U44153 ( .A(n35078), .B(n35080), .Z(n35179) );
  NAND U44154 ( .A(n35180), .B(n35181), .Z(n35080) );
  OR U44155 ( .A(n35182), .B(n35183), .Z(n35181) );
  OR U44156 ( .A(n35184), .B(n35185), .Z(n35180) );
  NAND U44157 ( .A(n35186), .B(n35187), .Z(n35078) );
  OR U44158 ( .A(n35188), .B(n35189), .Z(n35187) );
  OR U44159 ( .A(n35190), .B(n35191), .Z(n35186) );
  ANDN U44160 ( .B(n35192), .A(n35193), .Z(n35079) );
  IV U44161 ( .A(n35194), .Z(n35192) );
  XNOR U44162 ( .A(n35159), .B(n35158), .Z(N62282) );
  XOR U44163 ( .A(n35178), .B(n35177), .Z(n35158) );
  XNOR U44164 ( .A(n35193), .B(n35194), .Z(n35177) );
  XNOR U44165 ( .A(n35188), .B(n35189), .Z(n35194) );
  XNOR U44166 ( .A(n35190), .B(n35191), .Z(n35189) );
  XNOR U44167 ( .A(y[3133]), .B(x[3133]), .Z(n35191) );
  XNOR U44168 ( .A(y[3134]), .B(x[3134]), .Z(n35190) );
  XNOR U44169 ( .A(y[3132]), .B(x[3132]), .Z(n35188) );
  XNOR U44170 ( .A(n35182), .B(n35183), .Z(n35193) );
  XNOR U44171 ( .A(y[3129]), .B(x[3129]), .Z(n35183) );
  XNOR U44172 ( .A(n35184), .B(n35185), .Z(n35182) );
  XNOR U44173 ( .A(y[3130]), .B(x[3130]), .Z(n35185) );
  XNOR U44174 ( .A(y[3131]), .B(x[3131]), .Z(n35184) );
  XNOR U44175 ( .A(n35175), .B(n35174), .Z(n35178) );
  XNOR U44176 ( .A(n35170), .B(n35171), .Z(n35174) );
  XNOR U44177 ( .A(y[3126]), .B(x[3126]), .Z(n35171) );
  XNOR U44178 ( .A(n35172), .B(n35173), .Z(n35170) );
  XNOR U44179 ( .A(y[3127]), .B(x[3127]), .Z(n35173) );
  XNOR U44180 ( .A(y[3128]), .B(x[3128]), .Z(n35172) );
  XNOR U44181 ( .A(n35164), .B(n35165), .Z(n35175) );
  XNOR U44182 ( .A(y[3123]), .B(x[3123]), .Z(n35165) );
  XNOR U44183 ( .A(n35166), .B(n35167), .Z(n35164) );
  XNOR U44184 ( .A(y[3124]), .B(x[3124]), .Z(n35167) );
  XNOR U44185 ( .A(y[3125]), .B(x[3125]), .Z(n35166) );
  XOR U44186 ( .A(n35140), .B(n35141), .Z(n35159) );
  XNOR U44187 ( .A(n35156), .B(n35157), .Z(n35141) );
  XNOR U44188 ( .A(n35151), .B(n35152), .Z(n35157) );
  XNOR U44189 ( .A(n35153), .B(n35154), .Z(n35152) );
  XNOR U44190 ( .A(y[3121]), .B(x[3121]), .Z(n35154) );
  XNOR U44191 ( .A(y[3122]), .B(x[3122]), .Z(n35153) );
  XNOR U44192 ( .A(y[3120]), .B(x[3120]), .Z(n35151) );
  XNOR U44193 ( .A(n35145), .B(n35146), .Z(n35156) );
  XNOR U44194 ( .A(y[3117]), .B(x[3117]), .Z(n35146) );
  XNOR U44195 ( .A(n35147), .B(n35148), .Z(n35145) );
  XNOR U44196 ( .A(y[3118]), .B(x[3118]), .Z(n35148) );
  XNOR U44197 ( .A(y[3119]), .B(x[3119]), .Z(n35147) );
  XOR U44198 ( .A(n35139), .B(n35138), .Z(n35140) );
  XNOR U44199 ( .A(n35134), .B(n35135), .Z(n35138) );
  XNOR U44200 ( .A(y[3114]), .B(x[3114]), .Z(n35135) );
  XNOR U44201 ( .A(n35136), .B(n35137), .Z(n35134) );
  XNOR U44202 ( .A(y[3115]), .B(x[3115]), .Z(n35137) );
  XNOR U44203 ( .A(y[3116]), .B(x[3116]), .Z(n35136) );
  XNOR U44204 ( .A(n35128), .B(n35129), .Z(n35139) );
  XNOR U44205 ( .A(y[3111]), .B(x[3111]), .Z(n35129) );
  XNOR U44206 ( .A(n35130), .B(n35131), .Z(n35128) );
  XNOR U44207 ( .A(y[3112]), .B(x[3112]), .Z(n35131) );
  XNOR U44208 ( .A(y[3113]), .B(x[3113]), .Z(n35130) );
  NAND U44209 ( .A(n35195), .B(n35196), .Z(N62273) );
  NANDN U44210 ( .A(n35197), .B(n35198), .Z(n35196) );
  OR U44211 ( .A(n35199), .B(n35200), .Z(n35198) );
  NAND U44212 ( .A(n35199), .B(n35200), .Z(n35195) );
  XOR U44213 ( .A(n35199), .B(n35201), .Z(N62272) );
  XNOR U44214 ( .A(n35197), .B(n35200), .Z(n35201) );
  AND U44215 ( .A(n35202), .B(n35203), .Z(n35200) );
  NANDN U44216 ( .A(n35204), .B(n35205), .Z(n35203) );
  NANDN U44217 ( .A(n35206), .B(n35207), .Z(n35205) );
  NANDN U44218 ( .A(n35207), .B(n35206), .Z(n35202) );
  NAND U44219 ( .A(n35208), .B(n35209), .Z(n35197) );
  NANDN U44220 ( .A(n35210), .B(n35211), .Z(n35209) );
  OR U44221 ( .A(n35212), .B(n35213), .Z(n35211) );
  NAND U44222 ( .A(n35213), .B(n35212), .Z(n35208) );
  AND U44223 ( .A(n35214), .B(n35215), .Z(n35199) );
  NANDN U44224 ( .A(n35216), .B(n35217), .Z(n35215) );
  NANDN U44225 ( .A(n35218), .B(n35219), .Z(n35217) );
  NANDN U44226 ( .A(n35219), .B(n35218), .Z(n35214) );
  XOR U44227 ( .A(n35213), .B(n35220), .Z(N62271) );
  XOR U44228 ( .A(n35210), .B(n35212), .Z(n35220) );
  XNOR U44229 ( .A(n35206), .B(n35221), .Z(n35212) );
  XNOR U44230 ( .A(n35204), .B(n35207), .Z(n35221) );
  NAND U44231 ( .A(n35222), .B(n35223), .Z(n35207) );
  NAND U44232 ( .A(n35224), .B(n35225), .Z(n35223) );
  OR U44233 ( .A(n35226), .B(n35227), .Z(n35224) );
  NANDN U44234 ( .A(n35228), .B(n35226), .Z(n35222) );
  IV U44235 ( .A(n35227), .Z(n35228) );
  NAND U44236 ( .A(n35229), .B(n35230), .Z(n35204) );
  NAND U44237 ( .A(n35231), .B(n35232), .Z(n35230) );
  NANDN U44238 ( .A(n35233), .B(n35234), .Z(n35231) );
  NANDN U44239 ( .A(n35234), .B(n35233), .Z(n35229) );
  AND U44240 ( .A(n35235), .B(n35236), .Z(n35206) );
  NAND U44241 ( .A(n35237), .B(n35238), .Z(n35236) );
  OR U44242 ( .A(n35239), .B(n35240), .Z(n35237) );
  NANDN U44243 ( .A(n35241), .B(n35239), .Z(n35235) );
  NAND U44244 ( .A(n35242), .B(n35243), .Z(n35210) );
  NANDN U44245 ( .A(n35244), .B(n35245), .Z(n35243) );
  OR U44246 ( .A(n35246), .B(n35247), .Z(n35245) );
  NANDN U44247 ( .A(n35248), .B(n35246), .Z(n35242) );
  IV U44248 ( .A(n35247), .Z(n35248) );
  XNOR U44249 ( .A(n35218), .B(n35249), .Z(n35213) );
  XNOR U44250 ( .A(n35216), .B(n35219), .Z(n35249) );
  NAND U44251 ( .A(n35250), .B(n35251), .Z(n35219) );
  NAND U44252 ( .A(n35252), .B(n35253), .Z(n35251) );
  OR U44253 ( .A(n35254), .B(n35255), .Z(n35252) );
  NANDN U44254 ( .A(n35256), .B(n35254), .Z(n35250) );
  IV U44255 ( .A(n35255), .Z(n35256) );
  NAND U44256 ( .A(n35257), .B(n35258), .Z(n35216) );
  NAND U44257 ( .A(n35259), .B(n35260), .Z(n35258) );
  NANDN U44258 ( .A(n35261), .B(n35262), .Z(n35259) );
  NANDN U44259 ( .A(n35262), .B(n35261), .Z(n35257) );
  AND U44260 ( .A(n35263), .B(n35264), .Z(n35218) );
  NAND U44261 ( .A(n35265), .B(n35266), .Z(n35264) );
  OR U44262 ( .A(n35267), .B(n35268), .Z(n35265) );
  NANDN U44263 ( .A(n35269), .B(n35267), .Z(n35263) );
  XNOR U44264 ( .A(n35244), .B(n35270), .Z(N62270) );
  XOR U44265 ( .A(n35246), .B(n35247), .Z(n35270) );
  XNOR U44266 ( .A(n35260), .B(n35271), .Z(n35247) );
  XOR U44267 ( .A(n35261), .B(n35262), .Z(n35271) );
  XOR U44268 ( .A(n35267), .B(n35272), .Z(n35262) );
  XOR U44269 ( .A(n35266), .B(n35269), .Z(n35272) );
  IV U44270 ( .A(n35268), .Z(n35269) );
  NAND U44271 ( .A(n35273), .B(n35274), .Z(n35268) );
  OR U44272 ( .A(n35275), .B(n35276), .Z(n35274) );
  OR U44273 ( .A(n35277), .B(n35278), .Z(n35273) );
  NAND U44274 ( .A(n35279), .B(n35280), .Z(n35266) );
  OR U44275 ( .A(n35281), .B(n35282), .Z(n35280) );
  OR U44276 ( .A(n35283), .B(n35284), .Z(n35279) );
  NOR U44277 ( .A(n35285), .B(n35286), .Z(n35267) );
  ANDN U44278 ( .B(n35287), .A(n35288), .Z(n35261) );
  XNOR U44279 ( .A(n35254), .B(n35289), .Z(n35260) );
  XNOR U44280 ( .A(n35253), .B(n35255), .Z(n35289) );
  NAND U44281 ( .A(n35290), .B(n35291), .Z(n35255) );
  OR U44282 ( .A(n35292), .B(n35293), .Z(n35291) );
  OR U44283 ( .A(n35294), .B(n35295), .Z(n35290) );
  NAND U44284 ( .A(n35296), .B(n35297), .Z(n35253) );
  OR U44285 ( .A(n35298), .B(n35299), .Z(n35297) );
  OR U44286 ( .A(n35300), .B(n35301), .Z(n35296) );
  ANDN U44287 ( .B(n35302), .A(n35303), .Z(n35254) );
  IV U44288 ( .A(n35304), .Z(n35302) );
  ANDN U44289 ( .B(n35305), .A(n35306), .Z(n35246) );
  XOR U44290 ( .A(n35232), .B(n35307), .Z(n35244) );
  XOR U44291 ( .A(n35233), .B(n35234), .Z(n35307) );
  XOR U44292 ( .A(n35239), .B(n35308), .Z(n35234) );
  XOR U44293 ( .A(n35238), .B(n35241), .Z(n35308) );
  IV U44294 ( .A(n35240), .Z(n35241) );
  NAND U44295 ( .A(n35309), .B(n35310), .Z(n35240) );
  OR U44296 ( .A(n35311), .B(n35312), .Z(n35310) );
  OR U44297 ( .A(n35313), .B(n35314), .Z(n35309) );
  NAND U44298 ( .A(n35315), .B(n35316), .Z(n35238) );
  OR U44299 ( .A(n35317), .B(n35318), .Z(n35316) );
  OR U44300 ( .A(n35319), .B(n35320), .Z(n35315) );
  NOR U44301 ( .A(n35321), .B(n35322), .Z(n35239) );
  ANDN U44302 ( .B(n35323), .A(n35324), .Z(n35233) );
  IV U44303 ( .A(n35325), .Z(n35323) );
  XNOR U44304 ( .A(n35226), .B(n35326), .Z(n35232) );
  XNOR U44305 ( .A(n35225), .B(n35227), .Z(n35326) );
  NAND U44306 ( .A(n35327), .B(n35328), .Z(n35227) );
  OR U44307 ( .A(n35329), .B(n35330), .Z(n35328) );
  OR U44308 ( .A(n35331), .B(n35332), .Z(n35327) );
  NAND U44309 ( .A(n35333), .B(n35334), .Z(n35225) );
  OR U44310 ( .A(n35335), .B(n35336), .Z(n35334) );
  OR U44311 ( .A(n35337), .B(n35338), .Z(n35333) );
  ANDN U44312 ( .B(n35339), .A(n35340), .Z(n35226) );
  IV U44313 ( .A(n35341), .Z(n35339) );
  XNOR U44314 ( .A(n35306), .B(n35305), .Z(N62269) );
  XOR U44315 ( .A(n35325), .B(n35324), .Z(n35305) );
  XNOR U44316 ( .A(n35340), .B(n35341), .Z(n35324) );
  XNOR U44317 ( .A(n35335), .B(n35336), .Z(n35341) );
  XNOR U44318 ( .A(n35337), .B(n35338), .Z(n35336) );
  XNOR U44319 ( .A(y[3109]), .B(x[3109]), .Z(n35338) );
  XNOR U44320 ( .A(y[3110]), .B(x[3110]), .Z(n35337) );
  XNOR U44321 ( .A(y[3108]), .B(x[3108]), .Z(n35335) );
  XNOR U44322 ( .A(n35329), .B(n35330), .Z(n35340) );
  XNOR U44323 ( .A(y[3105]), .B(x[3105]), .Z(n35330) );
  XNOR U44324 ( .A(n35331), .B(n35332), .Z(n35329) );
  XNOR U44325 ( .A(y[3106]), .B(x[3106]), .Z(n35332) );
  XNOR U44326 ( .A(y[3107]), .B(x[3107]), .Z(n35331) );
  XNOR U44327 ( .A(n35322), .B(n35321), .Z(n35325) );
  XNOR U44328 ( .A(n35317), .B(n35318), .Z(n35321) );
  XNOR U44329 ( .A(y[3102]), .B(x[3102]), .Z(n35318) );
  XNOR U44330 ( .A(n35319), .B(n35320), .Z(n35317) );
  XNOR U44331 ( .A(y[3103]), .B(x[3103]), .Z(n35320) );
  XNOR U44332 ( .A(y[3104]), .B(x[3104]), .Z(n35319) );
  XNOR U44333 ( .A(n35311), .B(n35312), .Z(n35322) );
  XNOR U44334 ( .A(y[3099]), .B(x[3099]), .Z(n35312) );
  XNOR U44335 ( .A(n35313), .B(n35314), .Z(n35311) );
  XNOR U44336 ( .A(y[3100]), .B(x[3100]), .Z(n35314) );
  XNOR U44337 ( .A(y[3101]), .B(x[3101]), .Z(n35313) );
  XOR U44338 ( .A(n35287), .B(n35288), .Z(n35306) );
  XNOR U44339 ( .A(n35303), .B(n35304), .Z(n35288) );
  XNOR U44340 ( .A(n35298), .B(n35299), .Z(n35304) );
  XNOR U44341 ( .A(n35300), .B(n35301), .Z(n35299) );
  XNOR U44342 ( .A(y[3097]), .B(x[3097]), .Z(n35301) );
  XNOR U44343 ( .A(y[3098]), .B(x[3098]), .Z(n35300) );
  XNOR U44344 ( .A(y[3096]), .B(x[3096]), .Z(n35298) );
  XNOR U44345 ( .A(n35292), .B(n35293), .Z(n35303) );
  XNOR U44346 ( .A(y[3093]), .B(x[3093]), .Z(n35293) );
  XNOR U44347 ( .A(n35294), .B(n35295), .Z(n35292) );
  XNOR U44348 ( .A(y[3094]), .B(x[3094]), .Z(n35295) );
  XNOR U44349 ( .A(y[3095]), .B(x[3095]), .Z(n35294) );
  XOR U44350 ( .A(n35286), .B(n35285), .Z(n35287) );
  XNOR U44351 ( .A(n35281), .B(n35282), .Z(n35285) );
  XNOR U44352 ( .A(y[3090]), .B(x[3090]), .Z(n35282) );
  XNOR U44353 ( .A(n35283), .B(n35284), .Z(n35281) );
  XNOR U44354 ( .A(y[3091]), .B(x[3091]), .Z(n35284) );
  XNOR U44355 ( .A(y[3092]), .B(x[3092]), .Z(n35283) );
  XNOR U44356 ( .A(n35275), .B(n35276), .Z(n35286) );
  XNOR U44357 ( .A(y[3087]), .B(x[3087]), .Z(n35276) );
  XNOR U44358 ( .A(n35277), .B(n35278), .Z(n35275) );
  XNOR U44359 ( .A(y[3088]), .B(x[3088]), .Z(n35278) );
  XNOR U44360 ( .A(y[3089]), .B(x[3089]), .Z(n35277) );
  NAND U44361 ( .A(n35342), .B(n35343), .Z(N62260) );
  NANDN U44362 ( .A(n35344), .B(n35345), .Z(n35343) );
  OR U44363 ( .A(n35346), .B(n35347), .Z(n35345) );
  NAND U44364 ( .A(n35346), .B(n35347), .Z(n35342) );
  XOR U44365 ( .A(n35346), .B(n35348), .Z(N62259) );
  XNOR U44366 ( .A(n35344), .B(n35347), .Z(n35348) );
  AND U44367 ( .A(n35349), .B(n35350), .Z(n35347) );
  NANDN U44368 ( .A(n35351), .B(n35352), .Z(n35350) );
  NANDN U44369 ( .A(n35353), .B(n35354), .Z(n35352) );
  NANDN U44370 ( .A(n35354), .B(n35353), .Z(n35349) );
  NAND U44371 ( .A(n35355), .B(n35356), .Z(n35344) );
  NANDN U44372 ( .A(n35357), .B(n35358), .Z(n35356) );
  OR U44373 ( .A(n35359), .B(n35360), .Z(n35358) );
  NAND U44374 ( .A(n35360), .B(n35359), .Z(n35355) );
  AND U44375 ( .A(n35361), .B(n35362), .Z(n35346) );
  NANDN U44376 ( .A(n35363), .B(n35364), .Z(n35362) );
  NANDN U44377 ( .A(n35365), .B(n35366), .Z(n35364) );
  NANDN U44378 ( .A(n35366), .B(n35365), .Z(n35361) );
  XOR U44379 ( .A(n35360), .B(n35367), .Z(N62258) );
  XOR U44380 ( .A(n35357), .B(n35359), .Z(n35367) );
  XNOR U44381 ( .A(n35353), .B(n35368), .Z(n35359) );
  XNOR U44382 ( .A(n35351), .B(n35354), .Z(n35368) );
  NAND U44383 ( .A(n35369), .B(n35370), .Z(n35354) );
  NAND U44384 ( .A(n35371), .B(n35372), .Z(n35370) );
  OR U44385 ( .A(n35373), .B(n35374), .Z(n35371) );
  NANDN U44386 ( .A(n35375), .B(n35373), .Z(n35369) );
  IV U44387 ( .A(n35374), .Z(n35375) );
  NAND U44388 ( .A(n35376), .B(n35377), .Z(n35351) );
  NAND U44389 ( .A(n35378), .B(n35379), .Z(n35377) );
  NANDN U44390 ( .A(n35380), .B(n35381), .Z(n35378) );
  NANDN U44391 ( .A(n35381), .B(n35380), .Z(n35376) );
  AND U44392 ( .A(n35382), .B(n35383), .Z(n35353) );
  NAND U44393 ( .A(n35384), .B(n35385), .Z(n35383) );
  OR U44394 ( .A(n35386), .B(n35387), .Z(n35384) );
  NANDN U44395 ( .A(n35388), .B(n35386), .Z(n35382) );
  NAND U44396 ( .A(n35389), .B(n35390), .Z(n35357) );
  NANDN U44397 ( .A(n35391), .B(n35392), .Z(n35390) );
  OR U44398 ( .A(n35393), .B(n35394), .Z(n35392) );
  NANDN U44399 ( .A(n35395), .B(n35393), .Z(n35389) );
  IV U44400 ( .A(n35394), .Z(n35395) );
  XNOR U44401 ( .A(n35365), .B(n35396), .Z(n35360) );
  XNOR U44402 ( .A(n35363), .B(n35366), .Z(n35396) );
  NAND U44403 ( .A(n35397), .B(n35398), .Z(n35366) );
  NAND U44404 ( .A(n35399), .B(n35400), .Z(n35398) );
  OR U44405 ( .A(n35401), .B(n35402), .Z(n35399) );
  NANDN U44406 ( .A(n35403), .B(n35401), .Z(n35397) );
  IV U44407 ( .A(n35402), .Z(n35403) );
  NAND U44408 ( .A(n35404), .B(n35405), .Z(n35363) );
  NAND U44409 ( .A(n35406), .B(n35407), .Z(n35405) );
  NANDN U44410 ( .A(n35408), .B(n35409), .Z(n35406) );
  NANDN U44411 ( .A(n35409), .B(n35408), .Z(n35404) );
  AND U44412 ( .A(n35410), .B(n35411), .Z(n35365) );
  NAND U44413 ( .A(n35412), .B(n35413), .Z(n35411) );
  OR U44414 ( .A(n35414), .B(n35415), .Z(n35412) );
  NANDN U44415 ( .A(n35416), .B(n35414), .Z(n35410) );
  XNOR U44416 ( .A(n35391), .B(n35417), .Z(N62257) );
  XOR U44417 ( .A(n35393), .B(n35394), .Z(n35417) );
  XNOR U44418 ( .A(n35407), .B(n35418), .Z(n35394) );
  XOR U44419 ( .A(n35408), .B(n35409), .Z(n35418) );
  XOR U44420 ( .A(n35414), .B(n35419), .Z(n35409) );
  XOR U44421 ( .A(n35413), .B(n35416), .Z(n35419) );
  IV U44422 ( .A(n35415), .Z(n35416) );
  NAND U44423 ( .A(n35420), .B(n35421), .Z(n35415) );
  OR U44424 ( .A(n35422), .B(n35423), .Z(n35421) );
  OR U44425 ( .A(n35424), .B(n35425), .Z(n35420) );
  NAND U44426 ( .A(n35426), .B(n35427), .Z(n35413) );
  OR U44427 ( .A(n35428), .B(n35429), .Z(n35427) );
  OR U44428 ( .A(n35430), .B(n35431), .Z(n35426) );
  NOR U44429 ( .A(n35432), .B(n35433), .Z(n35414) );
  ANDN U44430 ( .B(n35434), .A(n35435), .Z(n35408) );
  XNOR U44431 ( .A(n35401), .B(n35436), .Z(n35407) );
  XNOR U44432 ( .A(n35400), .B(n35402), .Z(n35436) );
  NAND U44433 ( .A(n35437), .B(n35438), .Z(n35402) );
  OR U44434 ( .A(n35439), .B(n35440), .Z(n35438) );
  OR U44435 ( .A(n35441), .B(n35442), .Z(n35437) );
  NAND U44436 ( .A(n35443), .B(n35444), .Z(n35400) );
  OR U44437 ( .A(n35445), .B(n35446), .Z(n35444) );
  OR U44438 ( .A(n35447), .B(n35448), .Z(n35443) );
  ANDN U44439 ( .B(n35449), .A(n35450), .Z(n35401) );
  IV U44440 ( .A(n35451), .Z(n35449) );
  ANDN U44441 ( .B(n35452), .A(n35453), .Z(n35393) );
  XOR U44442 ( .A(n35379), .B(n35454), .Z(n35391) );
  XOR U44443 ( .A(n35380), .B(n35381), .Z(n35454) );
  XOR U44444 ( .A(n35386), .B(n35455), .Z(n35381) );
  XOR U44445 ( .A(n35385), .B(n35388), .Z(n35455) );
  IV U44446 ( .A(n35387), .Z(n35388) );
  NAND U44447 ( .A(n35456), .B(n35457), .Z(n35387) );
  OR U44448 ( .A(n35458), .B(n35459), .Z(n35457) );
  OR U44449 ( .A(n35460), .B(n35461), .Z(n35456) );
  NAND U44450 ( .A(n35462), .B(n35463), .Z(n35385) );
  OR U44451 ( .A(n35464), .B(n35465), .Z(n35463) );
  OR U44452 ( .A(n35466), .B(n35467), .Z(n35462) );
  NOR U44453 ( .A(n35468), .B(n35469), .Z(n35386) );
  ANDN U44454 ( .B(n35470), .A(n35471), .Z(n35380) );
  IV U44455 ( .A(n35472), .Z(n35470) );
  XNOR U44456 ( .A(n35373), .B(n35473), .Z(n35379) );
  XNOR U44457 ( .A(n35372), .B(n35374), .Z(n35473) );
  NAND U44458 ( .A(n35474), .B(n35475), .Z(n35374) );
  OR U44459 ( .A(n35476), .B(n35477), .Z(n35475) );
  OR U44460 ( .A(n35478), .B(n35479), .Z(n35474) );
  NAND U44461 ( .A(n35480), .B(n35481), .Z(n35372) );
  OR U44462 ( .A(n35482), .B(n35483), .Z(n35481) );
  OR U44463 ( .A(n35484), .B(n35485), .Z(n35480) );
  ANDN U44464 ( .B(n35486), .A(n35487), .Z(n35373) );
  IV U44465 ( .A(n35488), .Z(n35486) );
  XNOR U44466 ( .A(n35453), .B(n35452), .Z(N62256) );
  XOR U44467 ( .A(n35472), .B(n35471), .Z(n35452) );
  XNOR U44468 ( .A(n35487), .B(n35488), .Z(n35471) );
  XNOR U44469 ( .A(n35482), .B(n35483), .Z(n35488) );
  XNOR U44470 ( .A(n35484), .B(n35485), .Z(n35483) );
  XNOR U44471 ( .A(y[3085]), .B(x[3085]), .Z(n35485) );
  XNOR U44472 ( .A(y[3086]), .B(x[3086]), .Z(n35484) );
  XNOR U44473 ( .A(y[3084]), .B(x[3084]), .Z(n35482) );
  XNOR U44474 ( .A(n35476), .B(n35477), .Z(n35487) );
  XNOR U44475 ( .A(y[3081]), .B(x[3081]), .Z(n35477) );
  XNOR U44476 ( .A(n35478), .B(n35479), .Z(n35476) );
  XNOR U44477 ( .A(y[3082]), .B(x[3082]), .Z(n35479) );
  XNOR U44478 ( .A(y[3083]), .B(x[3083]), .Z(n35478) );
  XNOR U44479 ( .A(n35469), .B(n35468), .Z(n35472) );
  XNOR U44480 ( .A(n35464), .B(n35465), .Z(n35468) );
  XNOR U44481 ( .A(y[3078]), .B(x[3078]), .Z(n35465) );
  XNOR U44482 ( .A(n35466), .B(n35467), .Z(n35464) );
  XNOR U44483 ( .A(y[3079]), .B(x[3079]), .Z(n35467) );
  XNOR U44484 ( .A(y[3080]), .B(x[3080]), .Z(n35466) );
  XNOR U44485 ( .A(n35458), .B(n35459), .Z(n35469) );
  XNOR U44486 ( .A(y[3075]), .B(x[3075]), .Z(n35459) );
  XNOR U44487 ( .A(n35460), .B(n35461), .Z(n35458) );
  XNOR U44488 ( .A(y[3076]), .B(x[3076]), .Z(n35461) );
  XNOR U44489 ( .A(y[3077]), .B(x[3077]), .Z(n35460) );
  XOR U44490 ( .A(n35434), .B(n35435), .Z(n35453) );
  XNOR U44491 ( .A(n35450), .B(n35451), .Z(n35435) );
  XNOR U44492 ( .A(n35445), .B(n35446), .Z(n35451) );
  XNOR U44493 ( .A(n35447), .B(n35448), .Z(n35446) );
  XNOR U44494 ( .A(y[3073]), .B(x[3073]), .Z(n35448) );
  XNOR U44495 ( .A(y[3074]), .B(x[3074]), .Z(n35447) );
  XNOR U44496 ( .A(y[3072]), .B(x[3072]), .Z(n35445) );
  XNOR U44497 ( .A(n35439), .B(n35440), .Z(n35450) );
  XNOR U44498 ( .A(y[3069]), .B(x[3069]), .Z(n35440) );
  XNOR U44499 ( .A(n35441), .B(n35442), .Z(n35439) );
  XNOR U44500 ( .A(y[3070]), .B(x[3070]), .Z(n35442) );
  XNOR U44501 ( .A(y[3071]), .B(x[3071]), .Z(n35441) );
  XOR U44502 ( .A(n35433), .B(n35432), .Z(n35434) );
  XNOR U44503 ( .A(n35428), .B(n35429), .Z(n35432) );
  XNOR U44504 ( .A(y[3066]), .B(x[3066]), .Z(n35429) );
  XNOR U44505 ( .A(n35430), .B(n35431), .Z(n35428) );
  XNOR U44506 ( .A(y[3067]), .B(x[3067]), .Z(n35431) );
  XNOR U44507 ( .A(y[3068]), .B(x[3068]), .Z(n35430) );
  XNOR U44508 ( .A(n35422), .B(n35423), .Z(n35433) );
  XNOR U44509 ( .A(y[3063]), .B(x[3063]), .Z(n35423) );
  XNOR U44510 ( .A(n35424), .B(n35425), .Z(n35422) );
  XNOR U44511 ( .A(y[3064]), .B(x[3064]), .Z(n35425) );
  XNOR U44512 ( .A(y[3065]), .B(x[3065]), .Z(n35424) );
  NAND U44513 ( .A(n35489), .B(n35490), .Z(N62247) );
  NANDN U44514 ( .A(n35491), .B(n35492), .Z(n35490) );
  OR U44515 ( .A(n35493), .B(n35494), .Z(n35492) );
  NAND U44516 ( .A(n35493), .B(n35494), .Z(n35489) );
  XOR U44517 ( .A(n35493), .B(n35495), .Z(N62246) );
  XNOR U44518 ( .A(n35491), .B(n35494), .Z(n35495) );
  AND U44519 ( .A(n35496), .B(n35497), .Z(n35494) );
  NANDN U44520 ( .A(n35498), .B(n35499), .Z(n35497) );
  NANDN U44521 ( .A(n35500), .B(n35501), .Z(n35499) );
  NANDN U44522 ( .A(n35501), .B(n35500), .Z(n35496) );
  NAND U44523 ( .A(n35502), .B(n35503), .Z(n35491) );
  NANDN U44524 ( .A(n35504), .B(n35505), .Z(n35503) );
  OR U44525 ( .A(n35506), .B(n35507), .Z(n35505) );
  NAND U44526 ( .A(n35507), .B(n35506), .Z(n35502) );
  AND U44527 ( .A(n35508), .B(n35509), .Z(n35493) );
  NANDN U44528 ( .A(n35510), .B(n35511), .Z(n35509) );
  NANDN U44529 ( .A(n35512), .B(n35513), .Z(n35511) );
  NANDN U44530 ( .A(n35513), .B(n35512), .Z(n35508) );
  XOR U44531 ( .A(n35507), .B(n35514), .Z(N62245) );
  XOR U44532 ( .A(n35504), .B(n35506), .Z(n35514) );
  XNOR U44533 ( .A(n35500), .B(n35515), .Z(n35506) );
  XNOR U44534 ( .A(n35498), .B(n35501), .Z(n35515) );
  NAND U44535 ( .A(n35516), .B(n35517), .Z(n35501) );
  NAND U44536 ( .A(n35518), .B(n35519), .Z(n35517) );
  OR U44537 ( .A(n35520), .B(n35521), .Z(n35518) );
  NANDN U44538 ( .A(n35522), .B(n35520), .Z(n35516) );
  IV U44539 ( .A(n35521), .Z(n35522) );
  NAND U44540 ( .A(n35523), .B(n35524), .Z(n35498) );
  NAND U44541 ( .A(n35525), .B(n35526), .Z(n35524) );
  NANDN U44542 ( .A(n35527), .B(n35528), .Z(n35525) );
  NANDN U44543 ( .A(n35528), .B(n35527), .Z(n35523) );
  AND U44544 ( .A(n35529), .B(n35530), .Z(n35500) );
  NAND U44545 ( .A(n35531), .B(n35532), .Z(n35530) );
  OR U44546 ( .A(n35533), .B(n35534), .Z(n35531) );
  NANDN U44547 ( .A(n35535), .B(n35533), .Z(n35529) );
  NAND U44548 ( .A(n35536), .B(n35537), .Z(n35504) );
  NANDN U44549 ( .A(n35538), .B(n35539), .Z(n35537) );
  OR U44550 ( .A(n35540), .B(n35541), .Z(n35539) );
  NANDN U44551 ( .A(n35542), .B(n35540), .Z(n35536) );
  IV U44552 ( .A(n35541), .Z(n35542) );
  XNOR U44553 ( .A(n35512), .B(n35543), .Z(n35507) );
  XNOR U44554 ( .A(n35510), .B(n35513), .Z(n35543) );
  NAND U44555 ( .A(n35544), .B(n35545), .Z(n35513) );
  NAND U44556 ( .A(n35546), .B(n35547), .Z(n35545) );
  OR U44557 ( .A(n35548), .B(n35549), .Z(n35546) );
  NANDN U44558 ( .A(n35550), .B(n35548), .Z(n35544) );
  IV U44559 ( .A(n35549), .Z(n35550) );
  NAND U44560 ( .A(n35551), .B(n35552), .Z(n35510) );
  NAND U44561 ( .A(n35553), .B(n35554), .Z(n35552) );
  NANDN U44562 ( .A(n35555), .B(n35556), .Z(n35553) );
  NANDN U44563 ( .A(n35556), .B(n35555), .Z(n35551) );
  AND U44564 ( .A(n35557), .B(n35558), .Z(n35512) );
  NAND U44565 ( .A(n35559), .B(n35560), .Z(n35558) );
  OR U44566 ( .A(n35561), .B(n35562), .Z(n35559) );
  NANDN U44567 ( .A(n35563), .B(n35561), .Z(n35557) );
  XNOR U44568 ( .A(n35538), .B(n35564), .Z(N62244) );
  XOR U44569 ( .A(n35540), .B(n35541), .Z(n35564) );
  XNOR U44570 ( .A(n35554), .B(n35565), .Z(n35541) );
  XOR U44571 ( .A(n35555), .B(n35556), .Z(n35565) );
  XOR U44572 ( .A(n35561), .B(n35566), .Z(n35556) );
  XOR U44573 ( .A(n35560), .B(n35563), .Z(n35566) );
  IV U44574 ( .A(n35562), .Z(n35563) );
  NAND U44575 ( .A(n35567), .B(n35568), .Z(n35562) );
  OR U44576 ( .A(n35569), .B(n35570), .Z(n35568) );
  OR U44577 ( .A(n35571), .B(n35572), .Z(n35567) );
  NAND U44578 ( .A(n35573), .B(n35574), .Z(n35560) );
  OR U44579 ( .A(n35575), .B(n35576), .Z(n35574) );
  OR U44580 ( .A(n35577), .B(n35578), .Z(n35573) );
  NOR U44581 ( .A(n35579), .B(n35580), .Z(n35561) );
  ANDN U44582 ( .B(n35581), .A(n35582), .Z(n35555) );
  XNOR U44583 ( .A(n35548), .B(n35583), .Z(n35554) );
  XNOR U44584 ( .A(n35547), .B(n35549), .Z(n35583) );
  NAND U44585 ( .A(n35584), .B(n35585), .Z(n35549) );
  OR U44586 ( .A(n35586), .B(n35587), .Z(n35585) );
  OR U44587 ( .A(n35588), .B(n35589), .Z(n35584) );
  NAND U44588 ( .A(n35590), .B(n35591), .Z(n35547) );
  OR U44589 ( .A(n35592), .B(n35593), .Z(n35591) );
  OR U44590 ( .A(n35594), .B(n35595), .Z(n35590) );
  ANDN U44591 ( .B(n35596), .A(n35597), .Z(n35548) );
  IV U44592 ( .A(n35598), .Z(n35596) );
  ANDN U44593 ( .B(n35599), .A(n35600), .Z(n35540) );
  XOR U44594 ( .A(n35526), .B(n35601), .Z(n35538) );
  XOR U44595 ( .A(n35527), .B(n35528), .Z(n35601) );
  XOR U44596 ( .A(n35533), .B(n35602), .Z(n35528) );
  XOR U44597 ( .A(n35532), .B(n35535), .Z(n35602) );
  IV U44598 ( .A(n35534), .Z(n35535) );
  NAND U44599 ( .A(n35603), .B(n35604), .Z(n35534) );
  OR U44600 ( .A(n35605), .B(n35606), .Z(n35604) );
  OR U44601 ( .A(n35607), .B(n35608), .Z(n35603) );
  NAND U44602 ( .A(n35609), .B(n35610), .Z(n35532) );
  OR U44603 ( .A(n35611), .B(n35612), .Z(n35610) );
  OR U44604 ( .A(n35613), .B(n35614), .Z(n35609) );
  NOR U44605 ( .A(n35615), .B(n35616), .Z(n35533) );
  ANDN U44606 ( .B(n35617), .A(n35618), .Z(n35527) );
  IV U44607 ( .A(n35619), .Z(n35617) );
  XNOR U44608 ( .A(n35520), .B(n35620), .Z(n35526) );
  XNOR U44609 ( .A(n35519), .B(n35521), .Z(n35620) );
  NAND U44610 ( .A(n35621), .B(n35622), .Z(n35521) );
  OR U44611 ( .A(n35623), .B(n35624), .Z(n35622) );
  OR U44612 ( .A(n35625), .B(n35626), .Z(n35621) );
  NAND U44613 ( .A(n35627), .B(n35628), .Z(n35519) );
  OR U44614 ( .A(n35629), .B(n35630), .Z(n35628) );
  OR U44615 ( .A(n35631), .B(n35632), .Z(n35627) );
  ANDN U44616 ( .B(n35633), .A(n35634), .Z(n35520) );
  IV U44617 ( .A(n35635), .Z(n35633) );
  XNOR U44618 ( .A(n35600), .B(n35599), .Z(N62243) );
  XOR U44619 ( .A(n35619), .B(n35618), .Z(n35599) );
  XNOR U44620 ( .A(n35634), .B(n35635), .Z(n35618) );
  XNOR U44621 ( .A(n35629), .B(n35630), .Z(n35635) );
  XNOR U44622 ( .A(n35631), .B(n35632), .Z(n35630) );
  XNOR U44623 ( .A(y[3061]), .B(x[3061]), .Z(n35632) );
  XNOR U44624 ( .A(y[3062]), .B(x[3062]), .Z(n35631) );
  XNOR U44625 ( .A(y[3060]), .B(x[3060]), .Z(n35629) );
  XNOR U44626 ( .A(n35623), .B(n35624), .Z(n35634) );
  XNOR U44627 ( .A(y[3057]), .B(x[3057]), .Z(n35624) );
  XNOR U44628 ( .A(n35625), .B(n35626), .Z(n35623) );
  XNOR U44629 ( .A(y[3058]), .B(x[3058]), .Z(n35626) );
  XNOR U44630 ( .A(y[3059]), .B(x[3059]), .Z(n35625) );
  XNOR U44631 ( .A(n35616), .B(n35615), .Z(n35619) );
  XNOR U44632 ( .A(n35611), .B(n35612), .Z(n35615) );
  XNOR U44633 ( .A(y[3054]), .B(x[3054]), .Z(n35612) );
  XNOR U44634 ( .A(n35613), .B(n35614), .Z(n35611) );
  XNOR U44635 ( .A(y[3055]), .B(x[3055]), .Z(n35614) );
  XNOR U44636 ( .A(y[3056]), .B(x[3056]), .Z(n35613) );
  XNOR U44637 ( .A(n35605), .B(n35606), .Z(n35616) );
  XNOR U44638 ( .A(y[3051]), .B(x[3051]), .Z(n35606) );
  XNOR U44639 ( .A(n35607), .B(n35608), .Z(n35605) );
  XNOR U44640 ( .A(y[3052]), .B(x[3052]), .Z(n35608) );
  XNOR U44641 ( .A(y[3053]), .B(x[3053]), .Z(n35607) );
  XOR U44642 ( .A(n35581), .B(n35582), .Z(n35600) );
  XNOR U44643 ( .A(n35597), .B(n35598), .Z(n35582) );
  XNOR U44644 ( .A(n35592), .B(n35593), .Z(n35598) );
  XNOR U44645 ( .A(n35594), .B(n35595), .Z(n35593) );
  XNOR U44646 ( .A(y[3049]), .B(x[3049]), .Z(n35595) );
  XNOR U44647 ( .A(y[3050]), .B(x[3050]), .Z(n35594) );
  XNOR U44648 ( .A(y[3048]), .B(x[3048]), .Z(n35592) );
  XNOR U44649 ( .A(n35586), .B(n35587), .Z(n35597) );
  XNOR U44650 ( .A(y[3045]), .B(x[3045]), .Z(n35587) );
  XNOR U44651 ( .A(n35588), .B(n35589), .Z(n35586) );
  XNOR U44652 ( .A(y[3046]), .B(x[3046]), .Z(n35589) );
  XNOR U44653 ( .A(y[3047]), .B(x[3047]), .Z(n35588) );
  XOR U44654 ( .A(n35580), .B(n35579), .Z(n35581) );
  XNOR U44655 ( .A(n35575), .B(n35576), .Z(n35579) );
  XNOR U44656 ( .A(y[3042]), .B(x[3042]), .Z(n35576) );
  XNOR U44657 ( .A(n35577), .B(n35578), .Z(n35575) );
  XNOR U44658 ( .A(y[3043]), .B(x[3043]), .Z(n35578) );
  XNOR U44659 ( .A(y[3044]), .B(x[3044]), .Z(n35577) );
  XNOR U44660 ( .A(n35569), .B(n35570), .Z(n35580) );
  XNOR U44661 ( .A(y[3039]), .B(x[3039]), .Z(n35570) );
  XNOR U44662 ( .A(n35571), .B(n35572), .Z(n35569) );
  XNOR U44663 ( .A(y[3040]), .B(x[3040]), .Z(n35572) );
  XNOR U44664 ( .A(y[3041]), .B(x[3041]), .Z(n35571) );
  NAND U44665 ( .A(n35636), .B(n35637), .Z(N62234) );
  NANDN U44666 ( .A(n35638), .B(n35639), .Z(n35637) );
  OR U44667 ( .A(n35640), .B(n35641), .Z(n35639) );
  NAND U44668 ( .A(n35640), .B(n35641), .Z(n35636) );
  XOR U44669 ( .A(n35640), .B(n35642), .Z(N62233) );
  XNOR U44670 ( .A(n35638), .B(n35641), .Z(n35642) );
  AND U44671 ( .A(n35643), .B(n35644), .Z(n35641) );
  NANDN U44672 ( .A(n35645), .B(n35646), .Z(n35644) );
  NANDN U44673 ( .A(n35647), .B(n35648), .Z(n35646) );
  NANDN U44674 ( .A(n35648), .B(n35647), .Z(n35643) );
  NAND U44675 ( .A(n35649), .B(n35650), .Z(n35638) );
  NANDN U44676 ( .A(n35651), .B(n35652), .Z(n35650) );
  OR U44677 ( .A(n35653), .B(n35654), .Z(n35652) );
  NAND U44678 ( .A(n35654), .B(n35653), .Z(n35649) );
  AND U44679 ( .A(n35655), .B(n35656), .Z(n35640) );
  NANDN U44680 ( .A(n35657), .B(n35658), .Z(n35656) );
  NANDN U44681 ( .A(n35659), .B(n35660), .Z(n35658) );
  NANDN U44682 ( .A(n35660), .B(n35659), .Z(n35655) );
  XOR U44683 ( .A(n35654), .B(n35661), .Z(N62232) );
  XOR U44684 ( .A(n35651), .B(n35653), .Z(n35661) );
  XNOR U44685 ( .A(n35647), .B(n35662), .Z(n35653) );
  XNOR U44686 ( .A(n35645), .B(n35648), .Z(n35662) );
  NAND U44687 ( .A(n35663), .B(n35664), .Z(n35648) );
  NAND U44688 ( .A(n35665), .B(n35666), .Z(n35664) );
  OR U44689 ( .A(n35667), .B(n35668), .Z(n35665) );
  NANDN U44690 ( .A(n35669), .B(n35667), .Z(n35663) );
  IV U44691 ( .A(n35668), .Z(n35669) );
  NAND U44692 ( .A(n35670), .B(n35671), .Z(n35645) );
  NAND U44693 ( .A(n35672), .B(n35673), .Z(n35671) );
  NANDN U44694 ( .A(n35674), .B(n35675), .Z(n35672) );
  NANDN U44695 ( .A(n35675), .B(n35674), .Z(n35670) );
  AND U44696 ( .A(n35676), .B(n35677), .Z(n35647) );
  NAND U44697 ( .A(n35678), .B(n35679), .Z(n35677) );
  OR U44698 ( .A(n35680), .B(n35681), .Z(n35678) );
  NANDN U44699 ( .A(n35682), .B(n35680), .Z(n35676) );
  NAND U44700 ( .A(n35683), .B(n35684), .Z(n35651) );
  NANDN U44701 ( .A(n35685), .B(n35686), .Z(n35684) );
  OR U44702 ( .A(n35687), .B(n35688), .Z(n35686) );
  NANDN U44703 ( .A(n35689), .B(n35687), .Z(n35683) );
  IV U44704 ( .A(n35688), .Z(n35689) );
  XNOR U44705 ( .A(n35659), .B(n35690), .Z(n35654) );
  XNOR U44706 ( .A(n35657), .B(n35660), .Z(n35690) );
  NAND U44707 ( .A(n35691), .B(n35692), .Z(n35660) );
  NAND U44708 ( .A(n35693), .B(n35694), .Z(n35692) );
  OR U44709 ( .A(n35695), .B(n35696), .Z(n35693) );
  NANDN U44710 ( .A(n35697), .B(n35695), .Z(n35691) );
  IV U44711 ( .A(n35696), .Z(n35697) );
  NAND U44712 ( .A(n35698), .B(n35699), .Z(n35657) );
  NAND U44713 ( .A(n35700), .B(n35701), .Z(n35699) );
  NANDN U44714 ( .A(n35702), .B(n35703), .Z(n35700) );
  NANDN U44715 ( .A(n35703), .B(n35702), .Z(n35698) );
  AND U44716 ( .A(n35704), .B(n35705), .Z(n35659) );
  NAND U44717 ( .A(n35706), .B(n35707), .Z(n35705) );
  OR U44718 ( .A(n35708), .B(n35709), .Z(n35706) );
  NANDN U44719 ( .A(n35710), .B(n35708), .Z(n35704) );
  XNOR U44720 ( .A(n35685), .B(n35711), .Z(N62231) );
  XOR U44721 ( .A(n35687), .B(n35688), .Z(n35711) );
  XNOR U44722 ( .A(n35701), .B(n35712), .Z(n35688) );
  XOR U44723 ( .A(n35702), .B(n35703), .Z(n35712) );
  XOR U44724 ( .A(n35708), .B(n35713), .Z(n35703) );
  XOR U44725 ( .A(n35707), .B(n35710), .Z(n35713) );
  IV U44726 ( .A(n35709), .Z(n35710) );
  NAND U44727 ( .A(n35714), .B(n35715), .Z(n35709) );
  OR U44728 ( .A(n35716), .B(n35717), .Z(n35715) );
  OR U44729 ( .A(n35718), .B(n35719), .Z(n35714) );
  NAND U44730 ( .A(n35720), .B(n35721), .Z(n35707) );
  OR U44731 ( .A(n35722), .B(n35723), .Z(n35721) );
  OR U44732 ( .A(n35724), .B(n35725), .Z(n35720) );
  NOR U44733 ( .A(n35726), .B(n35727), .Z(n35708) );
  ANDN U44734 ( .B(n35728), .A(n35729), .Z(n35702) );
  XNOR U44735 ( .A(n35695), .B(n35730), .Z(n35701) );
  XNOR U44736 ( .A(n35694), .B(n35696), .Z(n35730) );
  NAND U44737 ( .A(n35731), .B(n35732), .Z(n35696) );
  OR U44738 ( .A(n35733), .B(n35734), .Z(n35732) );
  OR U44739 ( .A(n35735), .B(n35736), .Z(n35731) );
  NAND U44740 ( .A(n35737), .B(n35738), .Z(n35694) );
  OR U44741 ( .A(n35739), .B(n35740), .Z(n35738) );
  OR U44742 ( .A(n35741), .B(n35742), .Z(n35737) );
  ANDN U44743 ( .B(n35743), .A(n35744), .Z(n35695) );
  IV U44744 ( .A(n35745), .Z(n35743) );
  ANDN U44745 ( .B(n35746), .A(n35747), .Z(n35687) );
  XOR U44746 ( .A(n35673), .B(n35748), .Z(n35685) );
  XOR U44747 ( .A(n35674), .B(n35675), .Z(n35748) );
  XOR U44748 ( .A(n35680), .B(n35749), .Z(n35675) );
  XOR U44749 ( .A(n35679), .B(n35682), .Z(n35749) );
  IV U44750 ( .A(n35681), .Z(n35682) );
  NAND U44751 ( .A(n35750), .B(n35751), .Z(n35681) );
  OR U44752 ( .A(n35752), .B(n35753), .Z(n35751) );
  OR U44753 ( .A(n35754), .B(n35755), .Z(n35750) );
  NAND U44754 ( .A(n35756), .B(n35757), .Z(n35679) );
  OR U44755 ( .A(n35758), .B(n35759), .Z(n35757) );
  OR U44756 ( .A(n35760), .B(n35761), .Z(n35756) );
  NOR U44757 ( .A(n35762), .B(n35763), .Z(n35680) );
  ANDN U44758 ( .B(n35764), .A(n35765), .Z(n35674) );
  IV U44759 ( .A(n35766), .Z(n35764) );
  XNOR U44760 ( .A(n35667), .B(n35767), .Z(n35673) );
  XNOR U44761 ( .A(n35666), .B(n35668), .Z(n35767) );
  NAND U44762 ( .A(n35768), .B(n35769), .Z(n35668) );
  OR U44763 ( .A(n35770), .B(n35771), .Z(n35769) );
  OR U44764 ( .A(n35772), .B(n35773), .Z(n35768) );
  NAND U44765 ( .A(n35774), .B(n35775), .Z(n35666) );
  OR U44766 ( .A(n35776), .B(n35777), .Z(n35775) );
  OR U44767 ( .A(n35778), .B(n35779), .Z(n35774) );
  ANDN U44768 ( .B(n35780), .A(n35781), .Z(n35667) );
  IV U44769 ( .A(n35782), .Z(n35780) );
  XNOR U44770 ( .A(n35747), .B(n35746), .Z(N62230) );
  XOR U44771 ( .A(n35766), .B(n35765), .Z(n35746) );
  XNOR U44772 ( .A(n35781), .B(n35782), .Z(n35765) );
  XNOR U44773 ( .A(n35776), .B(n35777), .Z(n35782) );
  XNOR U44774 ( .A(n35778), .B(n35779), .Z(n35777) );
  XNOR U44775 ( .A(y[3037]), .B(x[3037]), .Z(n35779) );
  XNOR U44776 ( .A(y[3038]), .B(x[3038]), .Z(n35778) );
  XNOR U44777 ( .A(y[3036]), .B(x[3036]), .Z(n35776) );
  XNOR U44778 ( .A(n35770), .B(n35771), .Z(n35781) );
  XNOR U44779 ( .A(y[3033]), .B(x[3033]), .Z(n35771) );
  XNOR U44780 ( .A(n35772), .B(n35773), .Z(n35770) );
  XNOR U44781 ( .A(y[3034]), .B(x[3034]), .Z(n35773) );
  XNOR U44782 ( .A(y[3035]), .B(x[3035]), .Z(n35772) );
  XNOR U44783 ( .A(n35763), .B(n35762), .Z(n35766) );
  XNOR U44784 ( .A(n35758), .B(n35759), .Z(n35762) );
  XNOR U44785 ( .A(y[3030]), .B(x[3030]), .Z(n35759) );
  XNOR U44786 ( .A(n35760), .B(n35761), .Z(n35758) );
  XNOR U44787 ( .A(y[3031]), .B(x[3031]), .Z(n35761) );
  XNOR U44788 ( .A(y[3032]), .B(x[3032]), .Z(n35760) );
  XNOR U44789 ( .A(n35752), .B(n35753), .Z(n35763) );
  XNOR U44790 ( .A(y[3027]), .B(x[3027]), .Z(n35753) );
  XNOR U44791 ( .A(n35754), .B(n35755), .Z(n35752) );
  XNOR U44792 ( .A(y[3028]), .B(x[3028]), .Z(n35755) );
  XNOR U44793 ( .A(y[3029]), .B(x[3029]), .Z(n35754) );
  XOR U44794 ( .A(n35728), .B(n35729), .Z(n35747) );
  XNOR U44795 ( .A(n35744), .B(n35745), .Z(n35729) );
  XNOR U44796 ( .A(n35739), .B(n35740), .Z(n35745) );
  XNOR U44797 ( .A(n35741), .B(n35742), .Z(n35740) );
  XNOR U44798 ( .A(y[3025]), .B(x[3025]), .Z(n35742) );
  XNOR U44799 ( .A(y[3026]), .B(x[3026]), .Z(n35741) );
  XNOR U44800 ( .A(y[3024]), .B(x[3024]), .Z(n35739) );
  XNOR U44801 ( .A(n35733), .B(n35734), .Z(n35744) );
  XNOR U44802 ( .A(y[3021]), .B(x[3021]), .Z(n35734) );
  XNOR U44803 ( .A(n35735), .B(n35736), .Z(n35733) );
  XNOR U44804 ( .A(y[3022]), .B(x[3022]), .Z(n35736) );
  XNOR U44805 ( .A(y[3023]), .B(x[3023]), .Z(n35735) );
  XOR U44806 ( .A(n35727), .B(n35726), .Z(n35728) );
  XNOR U44807 ( .A(n35722), .B(n35723), .Z(n35726) );
  XNOR U44808 ( .A(y[3018]), .B(x[3018]), .Z(n35723) );
  XNOR U44809 ( .A(n35724), .B(n35725), .Z(n35722) );
  XNOR U44810 ( .A(y[3019]), .B(x[3019]), .Z(n35725) );
  XNOR U44811 ( .A(y[3020]), .B(x[3020]), .Z(n35724) );
  XNOR U44812 ( .A(n35716), .B(n35717), .Z(n35727) );
  XNOR U44813 ( .A(y[3015]), .B(x[3015]), .Z(n35717) );
  XNOR U44814 ( .A(n35718), .B(n35719), .Z(n35716) );
  XNOR U44815 ( .A(y[3016]), .B(x[3016]), .Z(n35719) );
  XNOR U44816 ( .A(y[3017]), .B(x[3017]), .Z(n35718) );
  NAND U44817 ( .A(n35783), .B(n35784), .Z(N62221) );
  NANDN U44818 ( .A(n35785), .B(n35786), .Z(n35784) );
  OR U44819 ( .A(n35787), .B(n35788), .Z(n35786) );
  NAND U44820 ( .A(n35787), .B(n35788), .Z(n35783) );
  XOR U44821 ( .A(n35787), .B(n35789), .Z(N62220) );
  XNOR U44822 ( .A(n35785), .B(n35788), .Z(n35789) );
  AND U44823 ( .A(n35790), .B(n35791), .Z(n35788) );
  NANDN U44824 ( .A(n35792), .B(n35793), .Z(n35791) );
  NANDN U44825 ( .A(n35794), .B(n35795), .Z(n35793) );
  NANDN U44826 ( .A(n35795), .B(n35794), .Z(n35790) );
  NAND U44827 ( .A(n35796), .B(n35797), .Z(n35785) );
  NANDN U44828 ( .A(n35798), .B(n35799), .Z(n35797) );
  OR U44829 ( .A(n35800), .B(n35801), .Z(n35799) );
  NAND U44830 ( .A(n35801), .B(n35800), .Z(n35796) );
  AND U44831 ( .A(n35802), .B(n35803), .Z(n35787) );
  NANDN U44832 ( .A(n35804), .B(n35805), .Z(n35803) );
  NANDN U44833 ( .A(n35806), .B(n35807), .Z(n35805) );
  NANDN U44834 ( .A(n35807), .B(n35806), .Z(n35802) );
  XOR U44835 ( .A(n35801), .B(n35808), .Z(N62219) );
  XOR U44836 ( .A(n35798), .B(n35800), .Z(n35808) );
  XNOR U44837 ( .A(n35794), .B(n35809), .Z(n35800) );
  XNOR U44838 ( .A(n35792), .B(n35795), .Z(n35809) );
  NAND U44839 ( .A(n35810), .B(n35811), .Z(n35795) );
  NAND U44840 ( .A(n35812), .B(n35813), .Z(n35811) );
  OR U44841 ( .A(n35814), .B(n35815), .Z(n35812) );
  NANDN U44842 ( .A(n35816), .B(n35814), .Z(n35810) );
  IV U44843 ( .A(n35815), .Z(n35816) );
  NAND U44844 ( .A(n35817), .B(n35818), .Z(n35792) );
  NAND U44845 ( .A(n35819), .B(n35820), .Z(n35818) );
  NANDN U44846 ( .A(n35821), .B(n35822), .Z(n35819) );
  NANDN U44847 ( .A(n35822), .B(n35821), .Z(n35817) );
  AND U44848 ( .A(n35823), .B(n35824), .Z(n35794) );
  NAND U44849 ( .A(n35825), .B(n35826), .Z(n35824) );
  OR U44850 ( .A(n35827), .B(n35828), .Z(n35825) );
  NANDN U44851 ( .A(n35829), .B(n35827), .Z(n35823) );
  NAND U44852 ( .A(n35830), .B(n35831), .Z(n35798) );
  NANDN U44853 ( .A(n35832), .B(n35833), .Z(n35831) );
  OR U44854 ( .A(n35834), .B(n35835), .Z(n35833) );
  NANDN U44855 ( .A(n35836), .B(n35834), .Z(n35830) );
  IV U44856 ( .A(n35835), .Z(n35836) );
  XNOR U44857 ( .A(n35806), .B(n35837), .Z(n35801) );
  XNOR U44858 ( .A(n35804), .B(n35807), .Z(n35837) );
  NAND U44859 ( .A(n35838), .B(n35839), .Z(n35807) );
  NAND U44860 ( .A(n35840), .B(n35841), .Z(n35839) );
  OR U44861 ( .A(n35842), .B(n35843), .Z(n35840) );
  NANDN U44862 ( .A(n35844), .B(n35842), .Z(n35838) );
  IV U44863 ( .A(n35843), .Z(n35844) );
  NAND U44864 ( .A(n35845), .B(n35846), .Z(n35804) );
  NAND U44865 ( .A(n35847), .B(n35848), .Z(n35846) );
  NANDN U44866 ( .A(n35849), .B(n35850), .Z(n35847) );
  NANDN U44867 ( .A(n35850), .B(n35849), .Z(n35845) );
  AND U44868 ( .A(n35851), .B(n35852), .Z(n35806) );
  NAND U44869 ( .A(n35853), .B(n35854), .Z(n35852) );
  OR U44870 ( .A(n35855), .B(n35856), .Z(n35853) );
  NANDN U44871 ( .A(n35857), .B(n35855), .Z(n35851) );
  XNOR U44872 ( .A(n35832), .B(n35858), .Z(N62218) );
  XOR U44873 ( .A(n35834), .B(n35835), .Z(n35858) );
  XNOR U44874 ( .A(n35848), .B(n35859), .Z(n35835) );
  XOR U44875 ( .A(n35849), .B(n35850), .Z(n35859) );
  XOR U44876 ( .A(n35855), .B(n35860), .Z(n35850) );
  XOR U44877 ( .A(n35854), .B(n35857), .Z(n35860) );
  IV U44878 ( .A(n35856), .Z(n35857) );
  NAND U44879 ( .A(n35861), .B(n35862), .Z(n35856) );
  OR U44880 ( .A(n35863), .B(n35864), .Z(n35862) );
  OR U44881 ( .A(n35865), .B(n35866), .Z(n35861) );
  NAND U44882 ( .A(n35867), .B(n35868), .Z(n35854) );
  OR U44883 ( .A(n35869), .B(n35870), .Z(n35868) );
  OR U44884 ( .A(n35871), .B(n35872), .Z(n35867) );
  NOR U44885 ( .A(n35873), .B(n35874), .Z(n35855) );
  ANDN U44886 ( .B(n35875), .A(n35876), .Z(n35849) );
  XNOR U44887 ( .A(n35842), .B(n35877), .Z(n35848) );
  XNOR U44888 ( .A(n35841), .B(n35843), .Z(n35877) );
  NAND U44889 ( .A(n35878), .B(n35879), .Z(n35843) );
  OR U44890 ( .A(n35880), .B(n35881), .Z(n35879) );
  OR U44891 ( .A(n35882), .B(n35883), .Z(n35878) );
  NAND U44892 ( .A(n35884), .B(n35885), .Z(n35841) );
  OR U44893 ( .A(n35886), .B(n35887), .Z(n35885) );
  OR U44894 ( .A(n35888), .B(n35889), .Z(n35884) );
  ANDN U44895 ( .B(n35890), .A(n35891), .Z(n35842) );
  IV U44896 ( .A(n35892), .Z(n35890) );
  ANDN U44897 ( .B(n35893), .A(n35894), .Z(n35834) );
  XOR U44898 ( .A(n35820), .B(n35895), .Z(n35832) );
  XOR U44899 ( .A(n35821), .B(n35822), .Z(n35895) );
  XOR U44900 ( .A(n35827), .B(n35896), .Z(n35822) );
  XOR U44901 ( .A(n35826), .B(n35829), .Z(n35896) );
  IV U44902 ( .A(n35828), .Z(n35829) );
  NAND U44903 ( .A(n35897), .B(n35898), .Z(n35828) );
  OR U44904 ( .A(n35899), .B(n35900), .Z(n35898) );
  OR U44905 ( .A(n35901), .B(n35902), .Z(n35897) );
  NAND U44906 ( .A(n35903), .B(n35904), .Z(n35826) );
  OR U44907 ( .A(n35905), .B(n35906), .Z(n35904) );
  OR U44908 ( .A(n35907), .B(n35908), .Z(n35903) );
  NOR U44909 ( .A(n35909), .B(n35910), .Z(n35827) );
  ANDN U44910 ( .B(n35911), .A(n35912), .Z(n35821) );
  IV U44911 ( .A(n35913), .Z(n35911) );
  XNOR U44912 ( .A(n35814), .B(n35914), .Z(n35820) );
  XNOR U44913 ( .A(n35813), .B(n35815), .Z(n35914) );
  NAND U44914 ( .A(n35915), .B(n35916), .Z(n35815) );
  OR U44915 ( .A(n35917), .B(n35918), .Z(n35916) );
  OR U44916 ( .A(n35919), .B(n35920), .Z(n35915) );
  NAND U44917 ( .A(n35921), .B(n35922), .Z(n35813) );
  OR U44918 ( .A(n35923), .B(n35924), .Z(n35922) );
  OR U44919 ( .A(n35925), .B(n35926), .Z(n35921) );
  ANDN U44920 ( .B(n35927), .A(n35928), .Z(n35814) );
  IV U44921 ( .A(n35929), .Z(n35927) );
  XNOR U44922 ( .A(n35894), .B(n35893), .Z(N62217) );
  XOR U44923 ( .A(n35913), .B(n35912), .Z(n35893) );
  XNOR U44924 ( .A(n35928), .B(n35929), .Z(n35912) );
  XNOR U44925 ( .A(n35923), .B(n35924), .Z(n35929) );
  XNOR U44926 ( .A(n35925), .B(n35926), .Z(n35924) );
  XNOR U44927 ( .A(y[3013]), .B(x[3013]), .Z(n35926) );
  XNOR U44928 ( .A(y[3014]), .B(x[3014]), .Z(n35925) );
  XNOR U44929 ( .A(y[3012]), .B(x[3012]), .Z(n35923) );
  XNOR U44930 ( .A(n35917), .B(n35918), .Z(n35928) );
  XNOR U44931 ( .A(y[3009]), .B(x[3009]), .Z(n35918) );
  XNOR U44932 ( .A(n35919), .B(n35920), .Z(n35917) );
  XNOR U44933 ( .A(y[3010]), .B(x[3010]), .Z(n35920) );
  XNOR U44934 ( .A(y[3011]), .B(x[3011]), .Z(n35919) );
  XNOR U44935 ( .A(n35910), .B(n35909), .Z(n35913) );
  XNOR U44936 ( .A(n35905), .B(n35906), .Z(n35909) );
  XNOR U44937 ( .A(y[3006]), .B(x[3006]), .Z(n35906) );
  XNOR U44938 ( .A(n35907), .B(n35908), .Z(n35905) );
  XNOR U44939 ( .A(y[3007]), .B(x[3007]), .Z(n35908) );
  XNOR U44940 ( .A(y[3008]), .B(x[3008]), .Z(n35907) );
  XNOR U44941 ( .A(n35899), .B(n35900), .Z(n35910) );
  XNOR U44942 ( .A(y[3003]), .B(x[3003]), .Z(n35900) );
  XNOR U44943 ( .A(n35901), .B(n35902), .Z(n35899) );
  XNOR U44944 ( .A(y[3004]), .B(x[3004]), .Z(n35902) );
  XNOR U44945 ( .A(y[3005]), .B(x[3005]), .Z(n35901) );
  XOR U44946 ( .A(n35875), .B(n35876), .Z(n35894) );
  XNOR U44947 ( .A(n35891), .B(n35892), .Z(n35876) );
  XNOR U44948 ( .A(n35886), .B(n35887), .Z(n35892) );
  XNOR U44949 ( .A(n35888), .B(n35889), .Z(n35887) );
  XNOR U44950 ( .A(y[3001]), .B(x[3001]), .Z(n35889) );
  XNOR U44951 ( .A(y[3002]), .B(x[3002]), .Z(n35888) );
  XNOR U44952 ( .A(y[3000]), .B(x[3000]), .Z(n35886) );
  XNOR U44953 ( .A(n35880), .B(n35881), .Z(n35891) );
  XNOR U44954 ( .A(y[2997]), .B(x[2997]), .Z(n35881) );
  XNOR U44955 ( .A(n35882), .B(n35883), .Z(n35880) );
  XNOR U44956 ( .A(y[2998]), .B(x[2998]), .Z(n35883) );
  XNOR U44957 ( .A(y[2999]), .B(x[2999]), .Z(n35882) );
  XOR U44958 ( .A(n35874), .B(n35873), .Z(n35875) );
  XNOR U44959 ( .A(n35869), .B(n35870), .Z(n35873) );
  XNOR U44960 ( .A(y[2994]), .B(x[2994]), .Z(n35870) );
  XNOR U44961 ( .A(n35871), .B(n35872), .Z(n35869) );
  XNOR U44962 ( .A(y[2995]), .B(x[2995]), .Z(n35872) );
  XNOR U44963 ( .A(y[2996]), .B(x[2996]), .Z(n35871) );
  XNOR U44964 ( .A(n35863), .B(n35864), .Z(n35874) );
  XNOR U44965 ( .A(y[2991]), .B(x[2991]), .Z(n35864) );
  XNOR U44966 ( .A(n35865), .B(n35866), .Z(n35863) );
  XNOR U44967 ( .A(y[2992]), .B(x[2992]), .Z(n35866) );
  XNOR U44968 ( .A(y[2993]), .B(x[2993]), .Z(n35865) );
  NAND U44969 ( .A(n35930), .B(n35931), .Z(N62208) );
  NANDN U44970 ( .A(n35932), .B(n35933), .Z(n35931) );
  OR U44971 ( .A(n35934), .B(n35935), .Z(n35933) );
  NAND U44972 ( .A(n35934), .B(n35935), .Z(n35930) );
  XOR U44973 ( .A(n35934), .B(n35936), .Z(N62207) );
  XNOR U44974 ( .A(n35932), .B(n35935), .Z(n35936) );
  AND U44975 ( .A(n35937), .B(n35938), .Z(n35935) );
  NANDN U44976 ( .A(n35939), .B(n35940), .Z(n35938) );
  NANDN U44977 ( .A(n35941), .B(n35942), .Z(n35940) );
  NANDN U44978 ( .A(n35942), .B(n35941), .Z(n35937) );
  NAND U44979 ( .A(n35943), .B(n35944), .Z(n35932) );
  NANDN U44980 ( .A(n35945), .B(n35946), .Z(n35944) );
  OR U44981 ( .A(n35947), .B(n35948), .Z(n35946) );
  NAND U44982 ( .A(n35948), .B(n35947), .Z(n35943) );
  AND U44983 ( .A(n35949), .B(n35950), .Z(n35934) );
  NANDN U44984 ( .A(n35951), .B(n35952), .Z(n35950) );
  NANDN U44985 ( .A(n35953), .B(n35954), .Z(n35952) );
  NANDN U44986 ( .A(n35954), .B(n35953), .Z(n35949) );
  XOR U44987 ( .A(n35948), .B(n35955), .Z(N62206) );
  XOR U44988 ( .A(n35945), .B(n35947), .Z(n35955) );
  XNOR U44989 ( .A(n35941), .B(n35956), .Z(n35947) );
  XNOR U44990 ( .A(n35939), .B(n35942), .Z(n35956) );
  NAND U44991 ( .A(n35957), .B(n35958), .Z(n35942) );
  NAND U44992 ( .A(n35959), .B(n35960), .Z(n35958) );
  OR U44993 ( .A(n35961), .B(n35962), .Z(n35959) );
  NANDN U44994 ( .A(n35963), .B(n35961), .Z(n35957) );
  IV U44995 ( .A(n35962), .Z(n35963) );
  NAND U44996 ( .A(n35964), .B(n35965), .Z(n35939) );
  NAND U44997 ( .A(n35966), .B(n35967), .Z(n35965) );
  NANDN U44998 ( .A(n35968), .B(n35969), .Z(n35966) );
  NANDN U44999 ( .A(n35969), .B(n35968), .Z(n35964) );
  AND U45000 ( .A(n35970), .B(n35971), .Z(n35941) );
  NAND U45001 ( .A(n35972), .B(n35973), .Z(n35971) );
  OR U45002 ( .A(n35974), .B(n35975), .Z(n35972) );
  NANDN U45003 ( .A(n35976), .B(n35974), .Z(n35970) );
  NAND U45004 ( .A(n35977), .B(n35978), .Z(n35945) );
  NANDN U45005 ( .A(n35979), .B(n35980), .Z(n35978) );
  OR U45006 ( .A(n35981), .B(n35982), .Z(n35980) );
  NANDN U45007 ( .A(n35983), .B(n35981), .Z(n35977) );
  IV U45008 ( .A(n35982), .Z(n35983) );
  XNOR U45009 ( .A(n35953), .B(n35984), .Z(n35948) );
  XNOR U45010 ( .A(n35951), .B(n35954), .Z(n35984) );
  NAND U45011 ( .A(n35985), .B(n35986), .Z(n35954) );
  NAND U45012 ( .A(n35987), .B(n35988), .Z(n35986) );
  OR U45013 ( .A(n35989), .B(n35990), .Z(n35987) );
  NANDN U45014 ( .A(n35991), .B(n35989), .Z(n35985) );
  IV U45015 ( .A(n35990), .Z(n35991) );
  NAND U45016 ( .A(n35992), .B(n35993), .Z(n35951) );
  NAND U45017 ( .A(n35994), .B(n35995), .Z(n35993) );
  NANDN U45018 ( .A(n35996), .B(n35997), .Z(n35994) );
  NANDN U45019 ( .A(n35997), .B(n35996), .Z(n35992) );
  AND U45020 ( .A(n35998), .B(n35999), .Z(n35953) );
  NAND U45021 ( .A(n36000), .B(n36001), .Z(n35999) );
  OR U45022 ( .A(n36002), .B(n36003), .Z(n36000) );
  NANDN U45023 ( .A(n36004), .B(n36002), .Z(n35998) );
  XNOR U45024 ( .A(n35979), .B(n36005), .Z(N62205) );
  XOR U45025 ( .A(n35981), .B(n35982), .Z(n36005) );
  XNOR U45026 ( .A(n35995), .B(n36006), .Z(n35982) );
  XOR U45027 ( .A(n35996), .B(n35997), .Z(n36006) );
  XOR U45028 ( .A(n36002), .B(n36007), .Z(n35997) );
  XOR U45029 ( .A(n36001), .B(n36004), .Z(n36007) );
  IV U45030 ( .A(n36003), .Z(n36004) );
  NAND U45031 ( .A(n36008), .B(n36009), .Z(n36003) );
  OR U45032 ( .A(n36010), .B(n36011), .Z(n36009) );
  OR U45033 ( .A(n36012), .B(n36013), .Z(n36008) );
  NAND U45034 ( .A(n36014), .B(n36015), .Z(n36001) );
  OR U45035 ( .A(n36016), .B(n36017), .Z(n36015) );
  OR U45036 ( .A(n36018), .B(n36019), .Z(n36014) );
  NOR U45037 ( .A(n36020), .B(n36021), .Z(n36002) );
  ANDN U45038 ( .B(n36022), .A(n36023), .Z(n35996) );
  XNOR U45039 ( .A(n35989), .B(n36024), .Z(n35995) );
  XNOR U45040 ( .A(n35988), .B(n35990), .Z(n36024) );
  NAND U45041 ( .A(n36025), .B(n36026), .Z(n35990) );
  OR U45042 ( .A(n36027), .B(n36028), .Z(n36026) );
  OR U45043 ( .A(n36029), .B(n36030), .Z(n36025) );
  NAND U45044 ( .A(n36031), .B(n36032), .Z(n35988) );
  OR U45045 ( .A(n36033), .B(n36034), .Z(n36032) );
  OR U45046 ( .A(n36035), .B(n36036), .Z(n36031) );
  ANDN U45047 ( .B(n36037), .A(n36038), .Z(n35989) );
  IV U45048 ( .A(n36039), .Z(n36037) );
  ANDN U45049 ( .B(n36040), .A(n36041), .Z(n35981) );
  XOR U45050 ( .A(n35967), .B(n36042), .Z(n35979) );
  XOR U45051 ( .A(n35968), .B(n35969), .Z(n36042) );
  XOR U45052 ( .A(n35974), .B(n36043), .Z(n35969) );
  XOR U45053 ( .A(n35973), .B(n35976), .Z(n36043) );
  IV U45054 ( .A(n35975), .Z(n35976) );
  NAND U45055 ( .A(n36044), .B(n36045), .Z(n35975) );
  OR U45056 ( .A(n36046), .B(n36047), .Z(n36045) );
  OR U45057 ( .A(n36048), .B(n36049), .Z(n36044) );
  NAND U45058 ( .A(n36050), .B(n36051), .Z(n35973) );
  OR U45059 ( .A(n36052), .B(n36053), .Z(n36051) );
  OR U45060 ( .A(n36054), .B(n36055), .Z(n36050) );
  NOR U45061 ( .A(n36056), .B(n36057), .Z(n35974) );
  ANDN U45062 ( .B(n36058), .A(n36059), .Z(n35968) );
  IV U45063 ( .A(n36060), .Z(n36058) );
  XNOR U45064 ( .A(n35961), .B(n36061), .Z(n35967) );
  XNOR U45065 ( .A(n35960), .B(n35962), .Z(n36061) );
  NAND U45066 ( .A(n36062), .B(n36063), .Z(n35962) );
  OR U45067 ( .A(n36064), .B(n36065), .Z(n36063) );
  OR U45068 ( .A(n36066), .B(n36067), .Z(n36062) );
  NAND U45069 ( .A(n36068), .B(n36069), .Z(n35960) );
  OR U45070 ( .A(n36070), .B(n36071), .Z(n36069) );
  OR U45071 ( .A(n36072), .B(n36073), .Z(n36068) );
  ANDN U45072 ( .B(n36074), .A(n36075), .Z(n35961) );
  IV U45073 ( .A(n36076), .Z(n36074) );
  XNOR U45074 ( .A(n36041), .B(n36040), .Z(N62204) );
  XOR U45075 ( .A(n36060), .B(n36059), .Z(n36040) );
  XNOR U45076 ( .A(n36075), .B(n36076), .Z(n36059) );
  XNOR U45077 ( .A(n36070), .B(n36071), .Z(n36076) );
  XNOR U45078 ( .A(n36072), .B(n36073), .Z(n36071) );
  XNOR U45079 ( .A(y[2989]), .B(x[2989]), .Z(n36073) );
  XNOR U45080 ( .A(y[2990]), .B(x[2990]), .Z(n36072) );
  XNOR U45081 ( .A(y[2988]), .B(x[2988]), .Z(n36070) );
  XNOR U45082 ( .A(n36064), .B(n36065), .Z(n36075) );
  XNOR U45083 ( .A(y[2985]), .B(x[2985]), .Z(n36065) );
  XNOR U45084 ( .A(n36066), .B(n36067), .Z(n36064) );
  XNOR U45085 ( .A(y[2986]), .B(x[2986]), .Z(n36067) );
  XNOR U45086 ( .A(y[2987]), .B(x[2987]), .Z(n36066) );
  XNOR U45087 ( .A(n36057), .B(n36056), .Z(n36060) );
  XNOR U45088 ( .A(n36052), .B(n36053), .Z(n36056) );
  XNOR U45089 ( .A(y[2982]), .B(x[2982]), .Z(n36053) );
  XNOR U45090 ( .A(n36054), .B(n36055), .Z(n36052) );
  XNOR U45091 ( .A(y[2983]), .B(x[2983]), .Z(n36055) );
  XNOR U45092 ( .A(y[2984]), .B(x[2984]), .Z(n36054) );
  XNOR U45093 ( .A(n36046), .B(n36047), .Z(n36057) );
  XNOR U45094 ( .A(y[2979]), .B(x[2979]), .Z(n36047) );
  XNOR U45095 ( .A(n36048), .B(n36049), .Z(n36046) );
  XNOR U45096 ( .A(y[2980]), .B(x[2980]), .Z(n36049) );
  XNOR U45097 ( .A(y[2981]), .B(x[2981]), .Z(n36048) );
  XOR U45098 ( .A(n36022), .B(n36023), .Z(n36041) );
  XNOR U45099 ( .A(n36038), .B(n36039), .Z(n36023) );
  XNOR U45100 ( .A(n36033), .B(n36034), .Z(n36039) );
  XNOR U45101 ( .A(n36035), .B(n36036), .Z(n36034) );
  XNOR U45102 ( .A(y[2977]), .B(x[2977]), .Z(n36036) );
  XNOR U45103 ( .A(y[2978]), .B(x[2978]), .Z(n36035) );
  XNOR U45104 ( .A(y[2976]), .B(x[2976]), .Z(n36033) );
  XNOR U45105 ( .A(n36027), .B(n36028), .Z(n36038) );
  XNOR U45106 ( .A(y[2973]), .B(x[2973]), .Z(n36028) );
  XNOR U45107 ( .A(n36029), .B(n36030), .Z(n36027) );
  XNOR U45108 ( .A(y[2974]), .B(x[2974]), .Z(n36030) );
  XNOR U45109 ( .A(y[2975]), .B(x[2975]), .Z(n36029) );
  XOR U45110 ( .A(n36021), .B(n36020), .Z(n36022) );
  XNOR U45111 ( .A(n36016), .B(n36017), .Z(n36020) );
  XNOR U45112 ( .A(y[2970]), .B(x[2970]), .Z(n36017) );
  XNOR U45113 ( .A(n36018), .B(n36019), .Z(n36016) );
  XNOR U45114 ( .A(y[2971]), .B(x[2971]), .Z(n36019) );
  XNOR U45115 ( .A(y[2972]), .B(x[2972]), .Z(n36018) );
  XNOR U45116 ( .A(n36010), .B(n36011), .Z(n36021) );
  XNOR U45117 ( .A(y[2967]), .B(x[2967]), .Z(n36011) );
  XNOR U45118 ( .A(n36012), .B(n36013), .Z(n36010) );
  XNOR U45119 ( .A(y[2968]), .B(x[2968]), .Z(n36013) );
  XNOR U45120 ( .A(y[2969]), .B(x[2969]), .Z(n36012) );
  NAND U45121 ( .A(n36077), .B(n36078), .Z(N62195) );
  NANDN U45122 ( .A(n36079), .B(n36080), .Z(n36078) );
  OR U45123 ( .A(n36081), .B(n36082), .Z(n36080) );
  NAND U45124 ( .A(n36081), .B(n36082), .Z(n36077) );
  XOR U45125 ( .A(n36081), .B(n36083), .Z(N62194) );
  XNOR U45126 ( .A(n36079), .B(n36082), .Z(n36083) );
  AND U45127 ( .A(n36084), .B(n36085), .Z(n36082) );
  NANDN U45128 ( .A(n36086), .B(n36087), .Z(n36085) );
  NANDN U45129 ( .A(n36088), .B(n36089), .Z(n36087) );
  NANDN U45130 ( .A(n36089), .B(n36088), .Z(n36084) );
  NAND U45131 ( .A(n36090), .B(n36091), .Z(n36079) );
  NANDN U45132 ( .A(n36092), .B(n36093), .Z(n36091) );
  OR U45133 ( .A(n36094), .B(n36095), .Z(n36093) );
  NAND U45134 ( .A(n36095), .B(n36094), .Z(n36090) );
  AND U45135 ( .A(n36096), .B(n36097), .Z(n36081) );
  NANDN U45136 ( .A(n36098), .B(n36099), .Z(n36097) );
  NANDN U45137 ( .A(n36100), .B(n36101), .Z(n36099) );
  NANDN U45138 ( .A(n36101), .B(n36100), .Z(n36096) );
  XOR U45139 ( .A(n36095), .B(n36102), .Z(N62193) );
  XOR U45140 ( .A(n36092), .B(n36094), .Z(n36102) );
  XNOR U45141 ( .A(n36088), .B(n36103), .Z(n36094) );
  XNOR U45142 ( .A(n36086), .B(n36089), .Z(n36103) );
  NAND U45143 ( .A(n36104), .B(n36105), .Z(n36089) );
  NAND U45144 ( .A(n36106), .B(n36107), .Z(n36105) );
  OR U45145 ( .A(n36108), .B(n36109), .Z(n36106) );
  NANDN U45146 ( .A(n36110), .B(n36108), .Z(n36104) );
  IV U45147 ( .A(n36109), .Z(n36110) );
  NAND U45148 ( .A(n36111), .B(n36112), .Z(n36086) );
  NAND U45149 ( .A(n36113), .B(n36114), .Z(n36112) );
  NANDN U45150 ( .A(n36115), .B(n36116), .Z(n36113) );
  NANDN U45151 ( .A(n36116), .B(n36115), .Z(n36111) );
  AND U45152 ( .A(n36117), .B(n36118), .Z(n36088) );
  NAND U45153 ( .A(n36119), .B(n36120), .Z(n36118) );
  OR U45154 ( .A(n36121), .B(n36122), .Z(n36119) );
  NANDN U45155 ( .A(n36123), .B(n36121), .Z(n36117) );
  NAND U45156 ( .A(n36124), .B(n36125), .Z(n36092) );
  NANDN U45157 ( .A(n36126), .B(n36127), .Z(n36125) );
  OR U45158 ( .A(n36128), .B(n36129), .Z(n36127) );
  NANDN U45159 ( .A(n36130), .B(n36128), .Z(n36124) );
  IV U45160 ( .A(n36129), .Z(n36130) );
  XNOR U45161 ( .A(n36100), .B(n36131), .Z(n36095) );
  XNOR U45162 ( .A(n36098), .B(n36101), .Z(n36131) );
  NAND U45163 ( .A(n36132), .B(n36133), .Z(n36101) );
  NAND U45164 ( .A(n36134), .B(n36135), .Z(n36133) );
  OR U45165 ( .A(n36136), .B(n36137), .Z(n36134) );
  NANDN U45166 ( .A(n36138), .B(n36136), .Z(n36132) );
  IV U45167 ( .A(n36137), .Z(n36138) );
  NAND U45168 ( .A(n36139), .B(n36140), .Z(n36098) );
  NAND U45169 ( .A(n36141), .B(n36142), .Z(n36140) );
  NANDN U45170 ( .A(n36143), .B(n36144), .Z(n36141) );
  NANDN U45171 ( .A(n36144), .B(n36143), .Z(n36139) );
  AND U45172 ( .A(n36145), .B(n36146), .Z(n36100) );
  NAND U45173 ( .A(n36147), .B(n36148), .Z(n36146) );
  OR U45174 ( .A(n36149), .B(n36150), .Z(n36147) );
  NANDN U45175 ( .A(n36151), .B(n36149), .Z(n36145) );
  XNOR U45176 ( .A(n36126), .B(n36152), .Z(N62192) );
  XOR U45177 ( .A(n36128), .B(n36129), .Z(n36152) );
  XNOR U45178 ( .A(n36142), .B(n36153), .Z(n36129) );
  XOR U45179 ( .A(n36143), .B(n36144), .Z(n36153) );
  XOR U45180 ( .A(n36149), .B(n36154), .Z(n36144) );
  XOR U45181 ( .A(n36148), .B(n36151), .Z(n36154) );
  IV U45182 ( .A(n36150), .Z(n36151) );
  NAND U45183 ( .A(n36155), .B(n36156), .Z(n36150) );
  OR U45184 ( .A(n36157), .B(n36158), .Z(n36156) );
  OR U45185 ( .A(n36159), .B(n36160), .Z(n36155) );
  NAND U45186 ( .A(n36161), .B(n36162), .Z(n36148) );
  OR U45187 ( .A(n36163), .B(n36164), .Z(n36162) );
  OR U45188 ( .A(n36165), .B(n36166), .Z(n36161) );
  NOR U45189 ( .A(n36167), .B(n36168), .Z(n36149) );
  ANDN U45190 ( .B(n36169), .A(n36170), .Z(n36143) );
  XNOR U45191 ( .A(n36136), .B(n36171), .Z(n36142) );
  XNOR U45192 ( .A(n36135), .B(n36137), .Z(n36171) );
  NAND U45193 ( .A(n36172), .B(n36173), .Z(n36137) );
  OR U45194 ( .A(n36174), .B(n36175), .Z(n36173) );
  OR U45195 ( .A(n36176), .B(n36177), .Z(n36172) );
  NAND U45196 ( .A(n36178), .B(n36179), .Z(n36135) );
  OR U45197 ( .A(n36180), .B(n36181), .Z(n36179) );
  OR U45198 ( .A(n36182), .B(n36183), .Z(n36178) );
  ANDN U45199 ( .B(n36184), .A(n36185), .Z(n36136) );
  IV U45200 ( .A(n36186), .Z(n36184) );
  ANDN U45201 ( .B(n36187), .A(n36188), .Z(n36128) );
  XOR U45202 ( .A(n36114), .B(n36189), .Z(n36126) );
  XOR U45203 ( .A(n36115), .B(n36116), .Z(n36189) );
  XOR U45204 ( .A(n36121), .B(n36190), .Z(n36116) );
  XOR U45205 ( .A(n36120), .B(n36123), .Z(n36190) );
  IV U45206 ( .A(n36122), .Z(n36123) );
  NAND U45207 ( .A(n36191), .B(n36192), .Z(n36122) );
  OR U45208 ( .A(n36193), .B(n36194), .Z(n36192) );
  OR U45209 ( .A(n36195), .B(n36196), .Z(n36191) );
  NAND U45210 ( .A(n36197), .B(n36198), .Z(n36120) );
  OR U45211 ( .A(n36199), .B(n36200), .Z(n36198) );
  OR U45212 ( .A(n36201), .B(n36202), .Z(n36197) );
  NOR U45213 ( .A(n36203), .B(n36204), .Z(n36121) );
  ANDN U45214 ( .B(n36205), .A(n36206), .Z(n36115) );
  IV U45215 ( .A(n36207), .Z(n36205) );
  XNOR U45216 ( .A(n36108), .B(n36208), .Z(n36114) );
  XNOR U45217 ( .A(n36107), .B(n36109), .Z(n36208) );
  NAND U45218 ( .A(n36209), .B(n36210), .Z(n36109) );
  OR U45219 ( .A(n36211), .B(n36212), .Z(n36210) );
  OR U45220 ( .A(n36213), .B(n36214), .Z(n36209) );
  NAND U45221 ( .A(n36215), .B(n36216), .Z(n36107) );
  OR U45222 ( .A(n36217), .B(n36218), .Z(n36216) );
  OR U45223 ( .A(n36219), .B(n36220), .Z(n36215) );
  ANDN U45224 ( .B(n36221), .A(n36222), .Z(n36108) );
  IV U45225 ( .A(n36223), .Z(n36221) );
  XNOR U45226 ( .A(n36188), .B(n36187), .Z(N62191) );
  XOR U45227 ( .A(n36207), .B(n36206), .Z(n36187) );
  XNOR U45228 ( .A(n36222), .B(n36223), .Z(n36206) );
  XNOR U45229 ( .A(n36217), .B(n36218), .Z(n36223) );
  XNOR U45230 ( .A(n36219), .B(n36220), .Z(n36218) );
  XNOR U45231 ( .A(y[2965]), .B(x[2965]), .Z(n36220) );
  XNOR U45232 ( .A(y[2966]), .B(x[2966]), .Z(n36219) );
  XNOR U45233 ( .A(y[2964]), .B(x[2964]), .Z(n36217) );
  XNOR U45234 ( .A(n36211), .B(n36212), .Z(n36222) );
  XNOR U45235 ( .A(y[2961]), .B(x[2961]), .Z(n36212) );
  XNOR U45236 ( .A(n36213), .B(n36214), .Z(n36211) );
  XNOR U45237 ( .A(y[2962]), .B(x[2962]), .Z(n36214) );
  XNOR U45238 ( .A(y[2963]), .B(x[2963]), .Z(n36213) );
  XNOR U45239 ( .A(n36204), .B(n36203), .Z(n36207) );
  XNOR U45240 ( .A(n36199), .B(n36200), .Z(n36203) );
  XNOR U45241 ( .A(y[2958]), .B(x[2958]), .Z(n36200) );
  XNOR U45242 ( .A(n36201), .B(n36202), .Z(n36199) );
  XNOR U45243 ( .A(y[2959]), .B(x[2959]), .Z(n36202) );
  XNOR U45244 ( .A(y[2960]), .B(x[2960]), .Z(n36201) );
  XNOR U45245 ( .A(n36193), .B(n36194), .Z(n36204) );
  XNOR U45246 ( .A(y[2955]), .B(x[2955]), .Z(n36194) );
  XNOR U45247 ( .A(n36195), .B(n36196), .Z(n36193) );
  XNOR U45248 ( .A(y[2956]), .B(x[2956]), .Z(n36196) );
  XNOR U45249 ( .A(y[2957]), .B(x[2957]), .Z(n36195) );
  XOR U45250 ( .A(n36169), .B(n36170), .Z(n36188) );
  XNOR U45251 ( .A(n36185), .B(n36186), .Z(n36170) );
  XNOR U45252 ( .A(n36180), .B(n36181), .Z(n36186) );
  XNOR U45253 ( .A(n36182), .B(n36183), .Z(n36181) );
  XNOR U45254 ( .A(y[2953]), .B(x[2953]), .Z(n36183) );
  XNOR U45255 ( .A(y[2954]), .B(x[2954]), .Z(n36182) );
  XNOR U45256 ( .A(y[2952]), .B(x[2952]), .Z(n36180) );
  XNOR U45257 ( .A(n36174), .B(n36175), .Z(n36185) );
  XNOR U45258 ( .A(y[2949]), .B(x[2949]), .Z(n36175) );
  XNOR U45259 ( .A(n36176), .B(n36177), .Z(n36174) );
  XNOR U45260 ( .A(y[2950]), .B(x[2950]), .Z(n36177) );
  XNOR U45261 ( .A(y[2951]), .B(x[2951]), .Z(n36176) );
  XOR U45262 ( .A(n36168), .B(n36167), .Z(n36169) );
  XNOR U45263 ( .A(n36163), .B(n36164), .Z(n36167) );
  XNOR U45264 ( .A(y[2946]), .B(x[2946]), .Z(n36164) );
  XNOR U45265 ( .A(n36165), .B(n36166), .Z(n36163) );
  XNOR U45266 ( .A(y[2947]), .B(x[2947]), .Z(n36166) );
  XNOR U45267 ( .A(y[2948]), .B(x[2948]), .Z(n36165) );
  XNOR U45268 ( .A(n36157), .B(n36158), .Z(n36168) );
  XNOR U45269 ( .A(y[2943]), .B(x[2943]), .Z(n36158) );
  XNOR U45270 ( .A(n36159), .B(n36160), .Z(n36157) );
  XNOR U45271 ( .A(y[2944]), .B(x[2944]), .Z(n36160) );
  XNOR U45272 ( .A(y[2945]), .B(x[2945]), .Z(n36159) );
  NAND U45273 ( .A(n36224), .B(n36225), .Z(N62182) );
  NANDN U45274 ( .A(n36226), .B(n36227), .Z(n36225) );
  OR U45275 ( .A(n36228), .B(n36229), .Z(n36227) );
  NAND U45276 ( .A(n36228), .B(n36229), .Z(n36224) );
  XOR U45277 ( .A(n36228), .B(n36230), .Z(N62181) );
  XNOR U45278 ( .A(n36226), .B(n36229), .Z(n36230) );
  AND U45279 ( .A(n36231), .B(n36232), .Z(n36229) );
  NANDN U45280 ( .A(n36233), .B(n36234), .Z(n36232) );
  NANDN U45281 ( .A(n36235), .B(n36236), .Z(n36234) );
  NANDN U45282 ( .A(n36236), .B(n36235), .Z(n36231) );
  NAND U45283 ( .A(n36237), .B(n36238), .Z(n36226) );
  NANDN U45284 ( .A(n36239), .B(n36240), .Z(n36238) );
  OR U45285 ( .A(n36241), .B(n36242), .Z(n36240) );
  NAND U45286 ( .A(n36242), .B(n36241), .Z(n36237) );
  AND U45287 ( .A(n36243), .B(n36244), .Z(n36228) );
  NANDN U45288 ( .A(n36245), .B(n36246), .Z(n36244) );
  NANDN U45289 ( .A(n36247), .B(n36248), .Z(n36246) );
  NANDN U45290 ( .A(n36248), .B(n36247), .Z(n36243) );
  XOR U45291 ( .A(n36242), .B(n36249), .Z(N62180) );
  XOR U45292 ( .A(n36239), .B(n36241), .Z(n36249) );
  XNOR U45293 ( .A(n36235), .B(n36250), .Z(n36241) );
  XNOR U45294 ( .A(n36233), .B(n36236), .Z(n36250) );
  NAND U45295 ( .A(n36251), .B(n36252), .Z(n36236) );
  NAND U45296 ( .A(n36253), .B(n36254), .Z(n36252) );
  OR U45297 ( .A(n36255), .B(n36256), .Z(n36253) );
  NANDN U45298 ( .A(n36257), .B(n36255), .Z(n36251) );
  IV U45299 ( .A(n36256), .Z(n36257) );
  NAND U45300 ( .A(n36258), .B(n36259), .Z(n36233) );
  NAND U45301 ( .A(n36260), .B(n36261), .Z(n36259) );
  NANDN U45302 ( .A(n36262), .B(n36263), .Z(n36260) );
  NANDN U45303 ( .A(n36263), .B(n36262), .Z(n36258) );
  AND U45304 ( .A(n36264), .B(n36265), .Z(n36235) );
  NAND U45305 ( .A(n36266), .B(n36267), .Z(n36265) );
  OR U45306 ( .A(n36268), .B(n36269), .Z(n36266) );
  NANDN U45307 ( .A(n36270), .B(n36268), .Z(n36264) );
  NAND U45308 ( .A(n36271), .B(n36272), .Z(n36239) );
  NANDN U45309 ( .A(n36273), .B(n36274), .Z(n36272) );
  OR U45310 ( .A(n36275), .B(n36276), .Z(n36274) );
  NANDN U45311 ( .A(n36277), .B(n36275), .Z(n36271) );
  IV U45312 ( .A(n36276), .Z(n36277) );
  XNOR U45313 ( .A(n36247), .B(n36278), .Z(n36242) );
  XNOR U45314 ( .A(n36245), .B(n36248), .Z(n36278) );
  NAND U45315 ( .A(n36279), .B(n36280), .Z(n36248) );
  NAND U45316 ( .A(n36281), .B(n36282), .Z(n36280) );
  OR U45317 ( .A(n36283), .B(n36284), .Z(n36281) );
  NANDN U45318 ( .A(n36285), .B(n36283), .Z(n36279) );
  IV U45319 ( .A(n36284), .Z(n36285) );
  NAND U45320 ( .A(n36286), .B(n36287), .Z(n36245) );
  NAND U45321 ( .A(n36288), .B(n36289), .Z(n36287) );
  NANDN U45322 ( .A(n36290), .B(n36291), .Z(n36288) );
  NANDN U45323 ( .A(n36291), .B(n36290), .Z(n36286) );
  AND U45324 ( .A(n36292), .B(n36293), .Z(n36247) );
  NAND U45325 ( .A(n36294), .B(n36295), .Z(n36293) );
  OR U45326 ( .A(n36296), .B(n36297), .Z(n36294) );
  NANDN U45327 ( .A(n36298), .B(n36296), .Z(n36292) );
  XNOR U45328 ( .A(n36273), .B(n36299), .Z(N62179) );
  XOR U45329 ( .A(n36275), .B(n36276), .Z(n36299) );
  XNOR U45330 ( .A(n36289), .B(n36300), .Z(n36276) );
  XOR U45331 ( .A(n36290), .B(n36291), .Z(n36300) );
  XOR U45332 ( .A(n36296), .B(n36301), .Z(n36291) );
  XOR U45333 ( .A(n36295), .B(n36298), .Z(n36301) );
  IV U45334 ( .A(n36297), .Z(n36298) );
  NAND U45335 ( .A(n36302), .B(n36303), .Z(n36297) );
  OR U45336 ( .A(n36304), .B(n36305), .Z(n36303) );
  OR U45337 ( .A(n36306), .B(n36307), .Z(n36302) );
  NAND U45338 ( .A(n36308), .B(n36309), .Z(n36295) );
  OR U45339 ( .A(n36310), .B(n36311), .Z(n36309) );
  OR U45340 ( .A(n36312), .B(n36313), .Z(n36308) );
  NOR U45341 ( .A(n36314), .B(n36315), .Z(n36296) );
  ANDN U45342 ( .B(n36316), .A(n36317), .Z(n36290) );
  XNOR U45343 ( .A(n36283), .B(n36318), .Z(n36289) );
  XNOR U45344 ( .A(n36282), .B(n36284), .Z(n36318) );
  NAND U45345 ( .A(n36319), .B(n36320), .Z(n36284) );
  OR U45346 ( .A(n36321), .B(n36322), .Z(n36320) );
  OR U45347 ( .A(n36323), .B(n36324), .Z(n36319) );
  NAND U45348 ( .A(n36325), .B(n36326), .Z(n36282) );
  OR U45349 ( .A(n36327), .B(n36328), .Z(n36326) );
  OR U45350 ( .A(n36329), .B(n36330), .Z(n36325) );
  ANDN U45351 ( .B(n36331), .A(n36332), .Z(n36283) );
  IV U45352 ( .A(n36333), .Z(n36331) );
  ANDN U45353 ( .B(n36334), .A(n36335), .Z(n36275) );
  XOR U45354 ( .A(n36261), .B(n36336), .Z(n36273) );
  XOR U45355 ( .A(n36262), .B(n36263), .Z(n36336) );
  XOR U45356 ( .A(n36268), .B(n36337), .Z(n36263) );
  XOR U45357 ( .A(n36267), .B(n36270), .Z(n36337) );
  IV U45358 ( .A(n36269), .Z(n36270) );
  NAND U45359 ( .A(n36338), .B(n36339), .Z(n36269) );
  OR U45360 ( .A(n36340), .B(n36341), .Z(n36339) );
  OR U45361 ( .A(n36342), .B(n36343), .Z(n36338) );
  NAND U45362 ( .A(n36344), .B(n36345), .Z(n36267) );
  OR U45363 ( .A(n36346), .B(n36347), .Z(n36345) );
  OR U45364 ( .A(n36348), .B(n36349), .Z(n36344) );
  NOR U45365 ( .A(n36350), .B(n36351), .Z(n36268) );
  ANDN U45366 ( .B(n36352), .A(n36353), .Z(n36262) );
  IV U45367 ( .A(n36354), .Z(n36352) );
  XNOR U45368 ( .A(n36255), .B(n36355), .Z(n36261) );
  XNOR U45369 ( .A(n36254), .B(n36256), .Z(n36355) );
  NAND U45370 ( .A(n36356), .B(n36357), .Z(n36256) );
  OR U45371 ( .A(n36358), .B(n36359), .Z(n36357) );
  OR U45372 ( .A(n36360), .B(n36361), .Z(n36356) );
  NAND U45373 ( .A(n36362), .B(n36363), .Z(n36254) );
  OR U45374 ( .A(n36364), .B(n36365), .Z(n36363) );
  OR U45375 ( .A(n36366), .B(n36367), .Z(n36362) );
  ANDN U45376 ( .B(n36368), .A(n36369), .Z(n36255) );
  IV U45377 ( .A(n36370), .Z(n36368) );
  XNOR U45378 ( .A(n36335), .B(n36334), .Z(N62178) );
  XOR U45379 ( .A(n36354), .B(n36353), .Z(n36334) );
  XNOR U45380 ( .A(n36369), .B(n36370), .Z(n36353) );
  XNOR U45381 ( .A(n36364), .B(n36365), .Z(n36370) );
  XNOR U45382 ( .A(n36366), .B(n36367), .Z(n36365) );
  XNOR U45383 ( .A(y[2941]), .B(x[2941]), .Z(n36367) );
  XNOR U45384 ( .A(y[2942]), .B(x[2942]), .Z(n36366) );
  XNOR U45385 ( .A(y[2940]), .B(x[2940]), .Z(n36364) );
  XNOR U45386 ( .A(n36358), .B(n36359), .Z(n36369) );
  XNOR U45387 ( .A(y[2937]), .B(x[2937]), .Z(n36359) );
  XNOR U45388 ( .A(n36360), .B(n36361), .Z(n36358) );
  XNOR U45389 ( .A(y[2938]), .B(x[2938]), .Z(n36361) );
  XNOR U45390 ( .A(y[2939]), .B(x[2939]), .Z(n36360) );
  XNOR U45391 ( .A(n36351), .B(n36350), .Z(n36354) );
  XNOR U45392 ( .A(n36346), .B(n36347), .Z(n36350) );
  XNOR U45393 ( .A(y[2934]), .B(x[2934]), .Z(n36347) );
  XNOR U45394 ( .A(n36348), .B(n36349), .Z(n36346) );
  XNOR U45395 ( .A(y[2935]), .B(x[2935]), .Z(n36349) );
  XNOR U45396 ( .A(y[2936]), .B(x[2936]), .Z(n36348) );
  XNOR U45397 ( .A(n36340), .B(n36341), .Z(n36351) );
  XNOR U45398 ( .A(y[2931]), .B(x[2931]), .Z(n36341) );
  XNOR U45399 ( .A(n36342), .B(n36343), .Z(n36340) );
  XNOR U45400 ( .A(y[2932]), .B(x[2932]), .Z(n36343) );
  XNOR U45401 ( .A(y[2933]), .B(x[2933]), .Z(n36342) );
  XOR U45402 ( .A(n36316), .B(n36317), .Z(n36335) );
  XNOR U45403 ( .A(n36332), .B(n36333), .Z(n36317) );
  XNOR U45404 ( .A(n36327), .B(n36328), .Z(n36333) );
  XNOR U45405 ( .A(n36329), .B(n36330), .Z(n36328) );
  XNOR U45406 ( .A(y[2929]), .B(x[2929]), .Z(n36330) );
  XNOR U45407 ( .A(y[2930]), .B(x[2930]), .Z(n36329) );
  XNOR U45408 ( .A(y[2928]), .B(x[2928]), .Z(n36327) );
  XNOR U45409 ( .A(n36321), .B(n36322), .Z(n36332) );
  XNOR U45410 ( .A(y[2925]), .B(x[2925]), .Z(n36322) );
  XNOR U45411 ( .A(n36323), .B(n36324), .Z(n36321) );
  XNOR U45412 ( .A(y[2926]), .B(x[2926]), .Z(n36324) );
  XNOR U45413 ( .A(y[2927]), .B(x[2927]), .Z(n36323) );
  XOR U45414 ( .A(n36315), .B(n36314), .Z(n36316) );
  XNOR U45415 ( .A(n36310), .B(n36311), .Z(n36314) );
  XNOR U45416 ( .A(y[2922]), .B(x[2922]), .Z(n36311) );
  XNOR U45417 ( .A(n36312), .B(n36313), .Z(n36310) );
  XNOR U45418 ( .A(y[2923]), .B(x[2923]), .Z(n36313) );
  XNOR U45419 ( .A(y[2924]), .B(x[2924]), .Z(n36312) );
  XNOR U45420 ( .A(n36304), .B(n36305), .Z(n36315) );
  XNOR U45421 ( .A(y[2919]), .B(x[2919]), .Z(n36305) );
  XNOR U45422 ( .A(n36306), .B(n36307), .Z(n36304) );
  XNOR U45423 ( .A(y[2920]), .B(x[2920]), .Z(n36307) );
  XNOR U45424 ( .A(y[2921]), .B(x[2921]), .Z(n36306) );
  NAND U45425 ( .A(n36371), .B(n36372), .Z(N62169) );
  NANDN U45426 ( .A(n36373), .B(n36374), .Z(n36372) );
  OR U45427 ( .A(n36375), .B(n36376), .Z(n36374) );
  NAND U45428 ( .A(n36375), .B(n36376), .Z(n36371) );
  XOR U45429 ( .A(n36375), .B(n36377), .Z(N62168) );
  XNOR U45430 ( .A(n36373), .B(n36376), .Z(n36377) );
  AND U45431 ( .A(n36378), .B(n36379), .Z(n36376) );
  NANDN U45432 ( .A(n36380), .B(n36381), .Z(n36379) );
  NANDN U45433 ( .A(n36382), .B(n36383), .Z(n36381) );
  NANDN U45434 ( .A(n36383), .B(n36382), .Z(n36378) );
  NAND U45435 ( .A(n36384), .B(n36385), .Z(n36373) );
  NANDN U45436 ( .A(n36386), .B(n36387), .Z(n36385) );
  OR U45437 ( .A(n36388), .B(n36389), .Z(n36387) );
  NAND U45438 ( .A(n36389), .B(n36388), .Z(n36384) );
  AND U45439 ( .A(n36390), .B(n36391), .Z(n36375) );
  NANDN U45440 ( .A(n36392), .B(n36393), .Z(n36391) );
  NANDN U45441 ( .A(n36394), .B(n36395), .Z(n36393) );
  NANDN U45442 ( .A(n36395), .B(n36394), .Z(n36390) );
  XOR U45443 ( .A(n36389), .B(n36396), .Z(N62167) );
  XOR U45444 ( .A(n36386), .B(n36388), .Z(n36396) );
  XNOR U45445 ( .A(n36382), .B(n36397), .Z(n36388) );
  XNOR U45446 ( .A(n36380), .B(n36383), .Z(n36397) );
  NAND U45447 ( .A(n36398), .B(n36399), .Z(n36383) );
  NAND U45448 ( .A(n36400), .B(n36401), .Z(n36399) );
  OR U45449 ( .A(n36402), .B(n36403), .Z(n36400) );
  NANDN U45450 ( .A(n36404), .B(n36402), .Z(n36398) );
  IV U45451 ( .A(n36403), .Z(n36404) );
  NAND U45452 ( .A(n36405), .B(n36406), .Z(n36380) );
  NAND U45453 ( .A(n36407), .B(n36408), .Z(n36406) );
  NANDN U45454 ( .A(n36409), .B(n36410), .Z(n36407) );
  NANDN U45455 ( .A(n36410), .B(n36409), .Z(n36405) );
  AND U45456 ( .A(n36411), .B(n36412), .Z(n36382) );
  NAND U45457 ( .A(n36413), .B(n36414), .Z(n36412) );
  OR U45458 ( .A(n36415), .B(n36416), .Z(n36413) );
  NANDN U45459 ( .A(n36417), .B(n36415), .Z(n36411) );
  NAND U45460 ( .A(n36418), .B(n36419), .Z(n36386) );
  NANDN U45461 ( .A(n36420), .B(n36421), .Z(n36419) );
  OR U45462 ( .A(n36422), .B(n36423), .Z(n36421) );
  NANDN U45463 ( .A(n36424), .B(n36422), .Z(n36418) );
  IV U45464 ( .A(n36423), .Z(n36424) );
  XNOR U45465 ( .A(n36394), .B(n36425), .Z(n36389) );
  XNOR U45466 ( .A(n36392), .B(n36395), .Z(n36425) );
  NAND U45467 ( .A(n36426), .B(n36427), .Z(n36395) );
  NAND U45468 ( .A(n36428), .B(n36429), .Z(n36427) );
  OR U45469 ( .A(n36430), .B(n36431), .Z(n36428) );
  NANDN U45470 ( .A(n36432), .B(n36430), .Z(n36426) );
  IV U45471 ( .A(n36431), .Z(n36432) );
  NAND U45472 ( .A(n36433), .B(n36434), .Z(n36392) );
  NAND U45473 ( .A(n36435), .B(n36436), .Z(n36434) );
  NANDN U45474 ( .A(n36437), .B(n36438), .Z(n36435) );
  NANDN U45475 ( .A(n36438), .B(n36437), .Z(n36433) );
  AND U45476 ( .A(n36439), .B(n36440), .Z(n36394) );
  NAND U45477 ( .A(n36441), .B(n36442), .Z(n36440) );
  OR U45478 ( .A(n36443), .B(n36444), .Z(n36441) );
  NANDN U45479 ( .A(n36445), .B(n36443), .Z(n36439) );
  XNOR U45480 ( .A(n36420), .B(n36446), .Z(N62166) );
  XOR U45481 ( .A(n36422), .B(n36423), .Z(n36446) );
  XNOR U45482 ( .A(n36436), .B(n36447), .Z(n36423) );
  XOR U45483 ( .A(n36437), .B(n36438), .Z(n36447) );
  XOR U45484 ( .A(n36443), .B(n36448), .Z(n36438) );
  XOR U45485 ( .A(n36442), .B(n36445), .Z(n36448) );
  IV U45486 ( .A(n36444), .Z(n36445) );
  NAND U45487 ( .A(n36449), .B(n36450), .Z(n36444) );
  OR U45488 ( .A(n36451), .B(n36452), .Z(n36450) );
  OR U45489 ( .A(n36453), .B(n36454), .Z(n36449) );
  NAND U45490 ( .A(n36455), .B(n36456), .Z(n36442) );
  OR U45491 ( .A(n36457), .B(n36458), .Z(n36456) );
  OR U45492 ( .A(n36459), .B(n36460), .Z(n36455) );
  NOR U45493 ( .A(n36461), .B(n36462), .Z(n36443) );
  ANDN U45494 ( .B(n36463), .A(n36464), .Z(n36437) );
  XNOR U45495 ( .A(n36430), .B(n36465), .Z(n36436) );
  XNOR U45496 ( .A(n36429), .B(n36431), .Z(n36465) );
  NAND U45497 ( .A(n36466), .B(n36467), .Z(n36431) );
  OR U45498 ( .A(n36468), .B(n36469), .Z(n36467) );
  OR U45499 ( .A(n36470), .B(n36471), .Z(n36466) );
  NAND U45500 ( .A(n36472), .B(n36473), .Z(n36429) );
  OR U45501 ( .A(n36474), .B(n36475), .Z(n36473) );
  OR U45502 ( .A(n36476), .B(n36477), .Z(n36472) );
  ANDN U45503 ( .B(n36478), .A(n36479), .Z(n36430) );
  IV U45504 ( .A(n36480), .Z(n36478) );
  ANDN U45505 ( .B(n36481), .A(n36482), .Z(n36422) );
  XOR U45506 ( .A(n36408), .B(n36483), .Z(n36420) );
  XOR U45507 ( .A(n36409), .B(n36410), .Z(n36483) );
  XOR U45508 ( .A(n36415), .B(n36484), .Z(n36410) );
  XOR U45509 ( .A(n36414), .B(n36417), .Z(n36484) );
  IV U45510 ( .A(n36416), .Z(n36417) );
  NAND U45511 ( .A(n36485), .B(n36486), .Z(n36416) );
  OR U45512 ( .A(n36487), .B(n36488), .Z(n36486) );
  OR U45513 ( .A(n36489), .B(n36490), .Z(n36485) );
  NAND U45514 ( .A(n36491), .B(n36492), .Z(n36414) );
  OR U45515 ( .A(n36493), .B(n36494), .Z(n36492) );
  OR U45516 ( .A(n36495), .B(n36496), .Z(n36491) );
  NOR U45517 ( .A(n36497), .B(n36498), .Z(n36415) );
  ANDN U45518 ( .B(n36499), .A(n36500), .Z(n36409) );
  IV U45519 ( .A(n36501), .Z(n36499) );
  XNOR U45520 ( .A(n36402), .B(n36502), .Z(n36408) );
  XNOR U45521 ( .A(n36401), .B(n36403), .Z(n36502) );
  NAND U45522 ( .A(n36503), .B(n36504), .Z(n36403) );
  OR U45523 ( .A(n36505), .B(n36506), .Z(n36504) );
  OR U45524 ( .A(n36507), .B(n36508), .Z(n36503) );
  NAND U45525 ( .A(n36509), .B(n36510), .Z(n36401) );
  OR U45526 ( .A(n36511), .B(n36512), .Z(n36510) );
  OR U45527 ( .A(n36513), .B(n36514), .Z(n36509) );
  ANDN U45528 ( .B(n36515), .A(n36516), .Z(n36402) );
  IV U45529 ( .A(n36517), .Z(n36515) );
  XNOR U45530 ( .A(n36482), .B(n36481), .Z(N62165) );
  XOR U45531 ( .A(n36501), .B(n36500), .Z(n36481) );
  XNOR U45532 ( .A(n36516), .B(n36517), .Z(n36500) );
  XNOR U45533 ( .A(n36511), .B(n36512), .Z(n36517) );
  XNOR U45534 ( .A(n36513), .B(n36514), .Z(n36512) );
  XNOR U45535 ( .A(y[2917]), .B(x[2917]), .Z(n36514) );
  XNOR U45536 ( .A(y[2918]), .B(x[2918]), .Z(n36513) );
  XNOR U45537 ( .A(y[2916]), .B(x[2916]), .Z(n36511) );
  XNOR U45538 ( .A(n36505), .B(n36506), .Z(n36516) );
  XNOR U45539 ( .A(y[2913]), .B(x[2913]), .Z(n36506) );
  XNOR U45540 ( .A(n36507), .B(n36508), .Z(n36505) );
  XNOR U45541 ( .A(y[2914]), .B(x[2914]), .Z(n36508) );
  XNOR U45542 ( .A(y[2915]), .B(x[2915]), .Z(n36507) );
  XNOR U45543 ( .A(n36498), .B(n36497), .Z(n36501) );
  XNOR U45544 ( .A(n36493), .B(n36494), .Z(n36497) );
  XNOR U45545 ( .A(y[2910]), .B(x[2910]), .Z(n36494) );
  XNOR U45546 ( .A(n36495), .B(n36496), .Z(n36493) );
  XNOR U45547 ( .A(y[2911]), .B(x[2911]), .Z(n36496) );
  XNOR U45548 ( .A(y[2912]), .B(x[2912]), .Z(n36495) );
  XNOR U45549 ( .A(n36487), .B(n36488), .Z(n36498) );
  XNOR U45550 ( .A(y[2907]), .B(x[2907]), .Z(n36488) );
  XNOR U45551 ( .A(n36489), .B(n36490), .Z(n36487) );
  XNOR U45552 ( .A(y[2908]), .B(x[2908]), .Z(n36490) );
  XNOR U45553 ( .A(y[2909]), .B(x[2909]), .Z(n36489) );
  XOR U45554 ( .A(n36463), .B(n36464), .Z(n36482) );
  XNOR U45555 ( .A(n36479), .B(n36480), .Z(n36464) );
  XNOR U45556 ( .A(n36474), .B(n36475), .Z(n36480) );
  XNOR U45557 ( .A(n36476), .B(n36477), .Z(n36475) );
  XNOR U45558 ( .A(y[2905]), .B(x[2905]), .Z(n36477) );
  XNOR U45559 ( .A(y[2906]), .B(x[2906]), .Z(n36476) );
  XNOR U45560 ( .A(y[2904]), .B(x[2904]), .Z(n36474) );
  XNOR U45561 ( .A(n36468), .B(n36469), .Z(n36479) );
  XNOR U45562 ( .A(y[2901]), .B(x[2901]), .Z(n36469) );
  XNOR U45563 ( .A(n36470), .B(n36471), .Z(n36468) );
  XNOR U45564 ( .A(y[2902]), .B(x[2902]), .Z(n36471) );
  XNOR U45565 ( .A(y[2903]), .B(x[2903]), .Z(n36470) );
  XOR U45566 ( .A(n36462), .B(n36461), .Z(n36463) );
  XNOR U45567 ( .A(n36457), .B(n36458), .Z(n36461) );
  XNOR U45568 ( .A(y[2898]), .B(x[2898]), .Z(n36458) );
  XNOR U45569 ( .A(n36459), .B(n36460), .Z(n36457) );
  XNOR U45570 ( .A(y[2899]), .B(x[2899]), .Z(n36460) );
  XNOR U45571 ( .A(y[2900]), .B(x[2900]), .Z(n36459) );
  XNOR U45572 ( .A(n36451), .B(n36452), .Z(n36462) );
  XNOR U45573 ( .A(y[2895]), .B(x[2895]), .Z(n36452) );
  XNOR U45574 ( .A(n36453), .B(n36454), .Z(n36451) );
  XNOR U45575 ( .A(y[2896]), .B(x[2896]), .Z(n36454) );
  XNOR U45576 ( .A(y[2897]), .B(x[2897]), .Z(n36453) );
  NAND U45577 ( .A(n36518), .B(n36519), .Z(N62156) );
  NANDN U45578 ( .A(n36520), .B(n36521), .Z(n36519) );
  OR U45579 ( .A(n36522), .B(n36523), .Z(n36521) );
  NAND U45580 ( .A(n36522), .B(n36523), .Z(n36518) );
  XOR U45581 ( .A(n36522), .B(n36524), .Z(N62155) );
  XNOR U45582 ( .A(n36520), .B(n36523), .Z(n36524) );
  AND U45583 ( .A(n36525), .B(n36526), .Z(n36523) );
  NANDN U45584 ( .A(n36527), .B(n36528), .Z(n36526) );
  NANDN U45585 ( .A(n36529), .B(n36530), .Z(n36528) );
  NANDN U45586 ( .A(n36530), .B(n36529), .Z(n36525) );
  NAND U45587 ( .A(n36531), .B(n36532), .Z(n36520) );
  NANDN U45588 ( .A(n36533), .B(n36534), .Z(n36532) );
  OR U45589 ( .A(n36535), .B(n36536), .Z(n36534) );
  NAND U45590 ( .A(n36536), .B(n36535), .Z(n36531) );
  AND U45591 ( .A(n36537), .B(n36538), .Z(n36522) );
  NANDN U45592 ( .A(n36539), .B(n36540), .Z(n36538) );
  NANDN U45593 ( .A(n36541), .B(n36542), .Z(n36540) );
  NANDN U45594 ( .A(n36542), .B(n36541), .Z(n36537) );
  XOR U45595 ( .A(n36536), .B(n36543), .Z(N62154) );
  XOR U45596 ( .A(n36533), .B(n36535), .Z(n36543) );
  XNOR U45597 ( .A(n36529), .B(n36544), .Z(n36535) );
  XNOR U45598 ( .A(n36527), .B(n36530), .Z(n36544) );
  NAND U45599 ( .A(n36545), .B(n36546), .Z(n36530) );
  NAND U45600 ( .A(n36547), .B(n36548), .Z(n36546) );
  OR U45601 ( .A(n36549), .B(n36550), .Z(n36547) );
  NANDN U45602 ( .A(n36551), .B(n36549), .Z(n36545) );
  IV U45603 ( .A(n36550), .Z(n36551) );
  NAND U45604 ( .A(n36552), .B(n36553), .Z(n36527) );
  NAND U45605 ( .A(n36554), .B(n36555), .Z(n36553) );
  NANDN U45606 ( .A(n36556), .B(n36557), .Z(n36554) );
  NANDN U45607 ( .A(n36557), .B(n36556), .Z(n36552) );
  AND U45608 ( .A(n36558), .B(n36559), .Z(n36529) );
  NAND U45609 ( .A(n36560), .B(n36561), .Z(n36559) );
  OR U45610 ( .A(n36562), .B(n36563), .Z(n36560) );
  NANDN U45611 ( .A(n36564), .B(n36562), .Z(n36558) );
  NAND U45612 ( .A(n36565), .B(n36566), .Z(n36533) );
  NANDN U45613 ( .A(n36567), .B(n36568), .Z(n36566) );
  OR U45614 ( .A(n36569), .B(n36570), .Z(n36568) );
  NANDN U45615 ( .A(n36571), .B(n36569), .Z(n36565) );
  IV U45616 ( .A(n36570), .Z(n36571) );
  XNOR U45617 ( .A(n36541), .B(n36572), .Z(n36536) );
  XNOR U45618 ( .A(n36539), .B(n36542), .Z(n36572) );
  NAND U45619 ( .A(n36573), .B(n36574), .Z(n36542) );
  NAND U45620 ( .A(n36575), .B(n36576), .Z(n36574) );
  OR U45621 ( .A(n36577), .B(n36578), .Z(n36575) );
  NANDN U45622 ( .A(n36579), .B(n36577), .Z(n36573) );
  IV U45623 ( .A(n36578), .Z(n36579) );
  NAND U45624 ( .A(n36580), .B(n36581), .Z(n36539) );
  NAND U45625 ( .A(n36582), .B(n36583), .Z(n36581) );
  NANDN U45626 ( .A(n36584), .B(n36585), .Z(n36582) );
  NANDN U45627 ( .A(n36585), .B(n36584), .Z(n36580) );
  AND U45628 ( .A(n36586), .B(n36587), .Z(n36541) );
  NAND U45629 ( .A(n36588), .B(n36589), .Z(n36587) );
  OR U45630 ( .A(n36590), .B(n36591), .Z(n36588) );
  NANDN U45631 ( .A(n36592), .B(n36590), .Z(n36586) );
  XNOR U45632 ( .A(n36567), .B(n36593), .Z(N62153) );
  XOR U45633 ( .A(n36569), .B(n36570), .Z(n36593) );
  XNOR U45634 ( .A(n36583), .B(n36594), .Z(n36570) );
  XOR U45635 ( .A(n36584), .B(n36585), .Z(n36594) );
  XOR U45636 ( .A(n36590), .B(n36595), .Z(n36585) );
  XOR U45637 ( .A(n36589), .B(n36592), .Z(n36595) );
  IV U45638 ( .A(n36591), .Z(n36592) );
  NAND U45639 ( .A(n36596), .B(n36597), .Z(n36591) );
  OR U45640 ( .A(n36598), .B(n36599), .Z(n36597) );
  OR U45641 ( .A(n36600), .B(n36601), .Z(n36596) );
  NAND U45642 ( .A(n36602), .B(n36603), .Z(n36589) );
  OR U45643 ( .A(n36604), .B(n36605), .Z(n36603) );
  OR U45644 ( .A(n36606), .B(n36607), .Z(n36602) );
  NOR U45645 ( .A(n36608), .B(n36609), .Z(n36590) );
  ANDN U45646 ( .B(n36610), .A(n36611), .Z(n36584) );
  XNOR U45647 ( .A(n36577), .B(n36612), .Z(n36583) );
  XNOR U45648 ( .A(n36576), .B(n36578), .Z(n36612) );
  NAND U45649 ( .A(n36613), .B(n36614), .Z(n36578) );
  OR U45650 ( .A(n36615), .B(n36616), .Z(n36614) );
  OR U45651 ( .A(n36617), .B(n36618), .Z(n36613) );
  NAND U45652 ( .A(n36619), .B(n36620), .Z(n36576) );
  OR U45653 ( .A(n36621), .B(n36622), .Z(n36620) );
  OR U45654 ( .A(n36623), .B(n36624), .Z(n36619) );
  ANDN U45655 ( .B(n36625), .A(n36626), .Z(n36577) );
  IV U45656 ( .A(n36627), .Z(n36625) );
  ANDN U45657 ( .B(n36628), .A(n36629), .Z(n36569) );
  XOR U45658 ( .A(n36555), .B(n36630), .Z(n36567) );
  XOR U45659 ( .A(n36556), .B(n36557), .Z(n36630) );
  XOR U45660 ( .A(n36562), .B(n36631), .Z(n36557) );
  XOR U45661 ( .A(n36561), .B(n36564), .Z(n36631) );
  IV U45662 ( .A(n36563), .Z(n36564) );
  NAND U45663 ( .A(n36632), .B(n36633), .Z(n36563) );
  OR U45664 ( .A(n36634), .B(n36635), .Z(n36633) );
  OR U45665 ( .A(n36636), .B(n36637), .Z(n36632) );
  NAND U45666 ( .A(n36638), .B(n36639), .Z(n36561) );
  OR U45667 ( .A(n36640), .B(n36641), .Z(n36639) );
  OR U45668 ( .A(n36642), .B(n36643), .Z(n36638) );
  NOR U45669 ( .A(n36644), .B(n36645), .Z(n36562) );
  ANDN U45670 ( .B(n36646), .A(n36647), .Z(n36556) );
  IV U45671 ( .A(n36648), .Z(n36646) );
  XNOR U45672 ( .A(n36549), .B(n36649), .Z(n36555) );
  XNOR U45673 ( .A(n36548), .B(n36550), .Z(n36649) );
  NAND U45674 ( .A(n36650), .B(n36651), .Z(n36550) );
  OR U45675 ( .A(n36652), .B(n36653), .Z(n36651) );
  OR U45676 ( .A(n36654), .B(n36655), .Z(n36650) );
  NAND U45677 ( .A(n36656), .B(n36657), .Z(n36548) );
  OR U45678 ( .A(n36658), .B(n36659), .Z(n36657) );
  OR U45679 ( .A(n36660), .B(n36661), .Z(n36656) );
  ANDN U45680 ( .B(n36662), .A(n36663), .Z(n36549) );
  IV U45681 ( .A(n36664), .Z(n36662) );
  XNOR U45682 ( .A(n36629), .B(n36628), .Z(N62152) );
  XOR U45683 ( .A(n36648), .B(n36647), .Z(n36628) );
  XNOR U45684 ( .A(n36663), .B(n36664), .Z(n36647) );
  XNOR U45685 ( .A(n36658), .B(n36659), .Z(n36664) );
  XNOR U45686 ( .A(n36660), .B(n36661), .Z(n36659) );
  XNOR U45687 ( .A(y[2893]), .B(x[2893]), .Z(n36661) );
  XNOR U45688 ( .A(y[2894]), .B(x[2894]), .Z(n36660) );
  XNOR U45689 ( .A(y[2892]), .B(x[2892]), .Z(n36658) );
  XNOR U45690 ( .A(n36652), .B(n36653), .Z(n36663) );
  XNOR U45691 ( .A(y[2889]), .B(x[2889]), .Z(n36653) );
  XNOR U45692 ( .A(n36654), .B(n36655), .Z(n36652) );
  XNOR U45693 ( .A(y[2890]), .B(x[2890]), .Z(n36655) );
  XNOR U45694 ( .A(y[2891]), .B(x[2891]), .Z(n36654) );
  XNOR U45695 ( .A(n36645), .B(n36644), .Z(n36648) );
  XNOR U45696 ( .A(n36640), .B(n36641), .Z(n36644) );
  XNOR U45697 ( .A(y[2886]), .B(x[2886]), .Z(n36641) );
  XNOR U45698 ( .A(n36642), .B(n36643), .Z(n36640) );
  XNOR U45699 ( .A(y[2887]), .B(x[2887]), .Z(n36643) );
  XNOR U45700 ( .A(y[2888]), .B(x[2888]), .Z(n36642) );
  XNOR U45701 ( .A(n36634), .B(n36635), .Z(n36645) );
  XNOR U45702 ( .A(y[2883]), .B(x[2883]), .Z(n36635) );
  XNOR U45703 ( .A(n36636), .B(n36637), .Z(n36634) );
  XNOR U45704 ( .A(y[2884]), .B(x[2884]), .Z(n36637) );
  XNOR U45705 ( .A(y[2885]), .B(x[2885]), .Z(n36636) );
  XOR U45706 ( .A(n36610), .B(n36611), .Z(n36629) );
  XNOR U45707 ( .A(n36626), .B(n36627), .Z(n36611) );
  XNOR U45708 ( .A(n36621), .B(n36622), .Z(n36627) );
  XNOR U45709 ( .A(n36623), .B(n36624), .Z(n36622) );
  XNOR U45710 ( .A(y[2881]), .B(x[2881]), .Z(n36624) );
  XNOR U45711 ( .A(y[2882]), .B(x[2882]), .Z(n36623) );
  XNOR U45712 ( .A(y[2880]), .B(x[2880]), .Z(n36621) );
  XNOR U45713 ( .A(n36615), .B(n36616), .Z(n36626) );
  XNOR U45714 ( .A(y[2877]), .B(x[2877]), .Z(n36616) );
  XNOR U45715 ( .A(n36617), .B(n36618), .Z(n36615) );
  XNOR U45716 ( .A(y[2878]), .B(x[2878]), .Z(n36618) );
  XNOR U45717 ( .A(y[2879]), .B(x[2879]), .Z(n36617) );
  XOR U45718 ( .A(n36609), .B(n36608), .Z(n36610) );
  XNOR U45719 ( .A(n36604), .B(n36605), .Z(n36608) );
  XNOR U45720 ( .A(y[2874]), .B(x[2874]), .Z(n36605) );
  XNOR U45721 ( .A(n36606), .B(n36607), .Z(n36604) );
  XNOR U45722 ( .A(y[2875]), .B(x[2875]), .Z(n36607) );
  XNOR U45723 ( .A(y[2876]), .B(x[2876]), .Z(n36606) );
  XNOR U45724 ( .A(n36598), .B(n36599), .Z(n36609) );
  XNOR U45725 ( .A(y[2871]), .B(x[2871]), .Z(n36599) );
  XNOR U45726 ( .A(n36600), .B(n36601), .Z(n36598) );
  XNOR U45727 ( .A(y[2872]), .B(x[2872]), .Z(n36601) );
  XNOR U45728 ( .A(y[2873]), .B(x[2873]), .Z(n36600) );
  NAND U45729 ( .A(n36665), .B(n36666), .Z(N62143) );
  NANDN U45730 ( .A(n36667), .B(n36668), .Z(n36666) );
  OR U45731 ( .A(n36669), .B(n36670), .Z(n36668) );
  NAND U45732 ( .A(n36669), .B(n36670), .Z(n36665) );
  XOR U45733 ( .A(n36669), .B(n36671), .Z(N62142) );
  XNOR U45734 ( .A(n36667), .B(n36670), .Z(n36671) );
  AND U45735 ( .A(n36672), .B(n36673), .Z(n36670) );
  NANDN U45736 ( .A(n36674), .B(n36675), .Z(n36673) );
  NANDN U45737 ( .A(n36676), .B(n36677), .Z(n36675) );
  NANDN U45738 ( .A(n36677), .B(n36676), .Z(n36672) );
  NAND U45739 ( .A(n36678), .B(n36679), .Z(n36667) );
  NANDN U45740 ( .A(n36680), .B(n36681), .Z(n36679) );
  OR U45741 ( .A(n36682), .B(n36683), .Z(n36681) );
  NAND U45742 ( .A(n36683), .B(n36682), .Z(n36678) );
  AND U45743 ( .A(n36684), .B(n36685), .Z(n36669) );
  NANDN U45744 ( .A(n36686), .B(n36687), .Z(n36685) );
  NANDN U45745 ( .A(n36688), .B(n36689), .Z(n36687) );
  NANDN U45746 ( .A(n36689), .B(n36688), .Z(n36684) );
  XOR U45747 ( .A(n36683), .B(n36690), .Z(N62141) );
  XOR U45748 ( .A(n36680), .B(n36682), .Z(n36690) );
  XNOR U45749 ( .A(n36676), .B(n36691), .Z(n36682) );
  XNOR U45750 ( .A(n36674), .B(n36677), .Z(n36691) );
  NAND U45751 ( .A(n36692), .B(n36693), .Z(n36677) );
  NAND U45752 ( .A(n36694), .B(n36695), .Z(n36693) );
  OR U45753 ( .A(n36696), .B(n36697), .Z(n36694) );
  NANDN U45754 ( .A(n36698), .B(n36696), .Z(n36692) );
  IV U45755 ( .A(n36697), .Z(n36698) );
  NAND U45756 ( .A(n36699), .B(n36700), .Z(n36674) );
  NAND U45757 ( .A(n36701), .B(n36702), .Z(n36700) );
  NANDN U45758 ( .A(n36703), .B(n36704), .Z(n36701) );
  NANDN U45759 ( .A(n36704), .B(n36703), .Z(n36699) );
  AND U45760 ( .A(n36705), .B(n36706), .Z(n36676) );
  NAND U45761 ( .A(n36707), .B(n36708), .Z(n36706) );
  OR U45762 ( .A(n36709), .B(n36710), .Z(n36707) );
  NANDN U45763 ( .A(n36711), .B(n36709), .Z(n36705) );
  NAND U45764 ( .A(n36712), .B(n36713), .Z(n36680) );
  NANDN U45765 ( .A(n36714), .B(n36715), .Z(n36713) );
  OR U45766 ( .A(n36716), .B(n36717), .Z(n36715) );
  NANDN U45767 ( .A(n36718), .B(n36716), .Z(n36712) );
  IV U45768 ( .A(n36717), .Z(n36718) );
  XNOR U45769 ( .A(n36688), .B(n36719), .Z(n36683) );
  XNOR U45770 ( .A(n36686), .B(n36689), .Z(n36719) );
  NAND U45771 ( .A(n36720), .B(n36721), .Z(n36689) );
  NAND U45772 ( .A(n36722), .B(n36723), .Z(n36721) );
  OR U45773 ( .A(n36724), .B(n36725), .Z(n36722) );
  NANDN U45774 ( .A(n36726), .B(n36724), .Z(n36720) );
  IV U45775 ( .A(n36725), .Z(n36726) );
  NAND U45776 ( .A(n36727), .B(n36728), .Z(n36686) );
  NAND U45777 ( .A(n36729), .B(n36730), .Z(n36728) );
  NANDN U45778 ( .A(n36731), .B(n36732), .Z(n36729) );
  NANDN U45779 ( .A(n36732), .B(n36731), .Z(n36727) );
  AND U45780 ( .A(n36733), .B(n36734), .Z(n36688) );
  NAND U45781 ( .A(n36735), .B(n36736), .Z(n36734) );
  OR U45782 ( .A(n36737), .B(n36738), .Z(n36735) );
  NANDN U45783 ( .A(n36739), .B(n36737), .Z(n36733) );
  XNOR U45784 ( .A(n36714), .B(n36740), .Z(N62140) );
  XOR U45785 ( .A(n36716), .B(n36717), .Z(n36740) );
  XNOR U45786 ( .A(n36730), .B(n36741), .Z(n36717) );
  XOR U45787 ( .A(n36731), .B(n36732), .Z(n36741) );
  XOR U45788 ( .A(n36737), .B(n36742), .Z(n36732) );
  XOR U45789 ( .A(n36736), .B(n36739), .Z(n36742) );
  IV U45790 ( .A(n36738), .Z(n36739) );
  NAND U45791 ( .A(n36743), .B(n36744), .Z(n36738) );
  OR U45792 ( .A(n36745), .B(n36746), .Z(n36744) );
  OR U45793 ( .A(n36747), .B(n36748), .Z(n36743) );
  NAND U45794 ( .A(n36749), .B(n36750), .Z(n36736) );
  OR U45795 ( .A(n36751), .B(n36752), .Z(n36750) );
  OR U45796 ( .A(n36753), .B(n36754), .Z(n36749) );
  NOR U45797 ( .A(n36755), .B(n36756), .Z(n36737) );
  ANDN U45798 ( .B(n36757), .A(n36758), .Z(n36731) );
  XNOR U45799 ( .A(n36724), .B(n36759), .Z(n36730) );
  XNOR U45800 ( .A(n36723), .B(n36725), .Z(n36759) );
  NAND U45801 ( .A(n36760), .B(n36761), .Z(n36725) );
  OR U45802 ( .A(n36762), .B(n36763), .Z(n36761) );
  OR U45803 ( .A(n36764), .B(n36765), .Z(n36760) );
  NAND U45804 ( .A(n36766), .B(n36767), .Z(n36723) );
  OR U45805 ( .A(n36768), .B(n36769), .Z(n36767) );
  OR U45806 ( .A(n36770), .B(n36771), .Z(n36766) );
  ANDN U45807 ( .B(n36772), .A(n36773), .Z(n36724) );
  IV U45808 ( .A(n36774), .Z(n36772) );
  ANDN U45809 ( .B(n36775), .A(n36776), .Z(n36716) );
  XOR U45810 ( .A(n36702), .B(n36777), .Z(n36714) );
  XOR U45811 ( .A(n36703), .B(n36704), .Z(n36777) );
  XOR U45812 ( .A(n36709), .B(n36778), .Z(n36704) );
  XOR U45813 ( .A(n36708), .B(n36711), .Z(n36778) );
  IV U45814 ( .A(n36710), .Z(n36711) );
  NAND U45815 ( .A(n36779), .B(n36780), .Z(n36710) );
  OR U45816 ( .A(n36781), .B(n36782), .Z(n36780) );
  OR U45817 ( .A(n36783), .B(n36784), .Z(n36779) );
  NAND U45818 ( .A(n36785), .B(n36786), .Z(n36708) );
  OR U45819 ( .A(n36787), .B(n36788), .Z(n36786) );
  OR U45820 ( .A(n36789), .B(n36790), .Z(n36785) );
  NOR U45821 ( .A(n36791), .B(n36792), .Z(n36709) );
  ANDN U45822 ( .B(n36793), .A(n36794), .Z(n36703) );
  IV U45823 ( .A(n36795), .Z(n36793) );
  XNOR U45824 ( .A(n36696), .B(n36796), .Z(n36702) );
  XNOR U45825 ( .A(n36695), .B(n36697), .Z(n36796) );
  NAND U45826 ( .A(n36797), .B(n36798), .Z(n36697) );
  OR U45827 ( .A(n36799), .B(n36800), .Z(n36798) );
  OR U45828 ( .A(n36801), .B(n36802), .Z(n36797) );
  NAND U45829 ( .A(n36803), .B(n36804), .Z(n36695) );
  OR U45830 ( .A(n36805), .B(n36806), .Z(n36804) );
  OR U45831 ( .A(n36807), .B(n36808), .Z(n36803) );
  ANDN U45832 ( .B(n36809), .A(n36810), .Z(n36696) );
  IV U45833 ( .A(n36811), .Z(n36809) );
  XNOR U45834 ( .A(n36776), .B(n36775), .Z(N62139) );
  XOR U45835 ( .A(n36795), .B(n36794), .Z(n36775) );
  XNOR U45836 ( .A(n36810), .B(n36811), .Z(n36794) );
  XNOR U45837 ( .A(n36805), .B(n36806), .Z(n36811) );
  XNOR U45838 ( .A(n36807), .B(n36808), .Z(n36806) );
  XNOR U45839 ( .A(y[2869]), .B(x[2869]), .Z(n36808) );
  XNOR U45840 ( .A(y[2870]), .B(x[2870]), .Z(n36807) );
  XNOR U45841 ( .A(y[2868]), .B(x[2868]), .Z(n36805) );
  XNOR U45842 ( .A(n36799), .B(n36800), .Z(n36810) );
  XNOR U45843 ( .A(y[2865]), .B(x[2865]), .Z(n36800) );
  XNOR U45844 ( .A(n36801), .B(n36802), .Z(n36799) );
  XNOR U45845 ( .A(y[2866]), .B(x[2866]), .Z(n36802) );
  XNOR U45846 ( .A(y[2867]), .B(x[2867]), .Z(n36801) );
  XNOR U45847 ( .A(n36792), .B(n36791), .Z(n36795) );
  XNOR U45848 ( .A(n36787), .B(n36788), .Z(n36791) );
  XNOR U45849 ( .A(y[2862]), .B(x[2862]), .Z(n36788) );
  XNOR U45850 ( .A(n36789), .B(n36790), .Z(n36787) );
  XNOR U45851 ( .A(y[2863]), .B(x[2863]), .Z(n36790) );
  XNOR U45852 ( .A(y[2864]), .B(x[2864]), .Z(n36789) );
  XNOR U45853 ( .A(n36781), .B(n36782), .Z(n36792) );
  XNOR U45854 ( .A(y[2859]), .B(x[2859]), .Z(n36782) );
  XNOR U45855 ( .A(n36783), .B(n36784), .Z(n36781) );
  XNOR U45856 ( .A(y[2860]), .B(x[2860]), .Z(n36784) );
  XNOR U45857 ( .A(y[2861]), .B(x[2861]), .Z(n36783) );
  XOR U45858 ( .A(n36757), .B(n36758), .Z(n36776) );
  XNOR U45859 ( .A(n36773), .B(n36774), .Z(n36758) );
  XNOR U45860 ( .A(n36768), .B(n36769), .Z(n36774) );
  XNOR U45861 ( .A(n36770), .B(n36771), .Z(n36769) );
  XNOR U45862 ( .A(y[2857]), .B(x[2857]), .Z(n36771) );
  XNOR U45863 ( .A(y[2858]), .B(x[2858]), .Z(n36770) );
  XNOR U45864 ( .A(y[2856]), .B(x[2856]), .Z(n36768) );
  XNOR U45865 ( .A(n36762), .B(n36763), .Z(n36773) );
  XNOR U45866 ( .A(y[2853]), .B(x[2853]), .Z(n36763) );
  XNOR U45867 ( .A(n36764), .B(n36765), .Z(n36762) );
  XNOR U45868 ( .A(y[2854]), .B(x[2854]), .Z(n36765) );
  XNOR U45869 ( .A(y[2855]), .B(x[2855]), .Z(n36764) );
  XOR U45870 ( .A(n36756), .B(n36755), .Z(n36757) );
  XNOR U45871 ( .A(n36751), .B(n36752), .Z(n36755) );
  XNOR U45872 ( .A(y[2850]), .B(x[2850]), .Z(n36752) );
  XNOR U45873 ( .A(n36753), .B(n36754), .Z(n36751) );
  XNOR U45874 ( .A(y[2851]), .B(x[2851]), .Z(n36754) );
  XNOR U45875 ( .A(y[2852]), .B(x[2852]), .Z(n36753) );
  XNOR U45876 ( .A(n36745), .B(n36746), .Z(n36756) );
  XNOR U45877 ( .A(y[2847]), .B(x[2847]), .Z(n36746) );
  XNOR U45878 ( .A(n36747), .B(n36748), .Z(n36745) );
  XNOR U45879 ( .A(y[2848]), .B(x[2848]), .Z(n36748) );
  XNOR U45880 ( .A(y[2849]), .B(x[2849]), .Z(n36747) );
  NAND U45881 ( .A(n36812), .B(n36813), .Z(N62130) );
  NANDN U45882 ( .A(n36814), .B(n36815), .Z(n36813) );
  OR U45883 ( .A(n36816), .B(n36817), .Z(n36815) );
  NAND U45884 ( .A(n36816), .B(n36817), .Z(n36812) );
  XOR U45885 ( .A(n36816), .B(n36818), .Z(N62129) );
  XNOR U45886 ( .A(n36814), .B(n36817), .Z(n36818) );
  AND U45887 ( .A(n36819), .B(n36820), .Z(n36817) );
  NANDN U45888 ( .A(n36821), .B(n36822), .Z(n36820) );
  NANDN U45889 ( .A(n36823), .B(n36824), .Z(n36822) );
  NANDN U45890 ( .A(n36824), .B(n36823), .Z(n36819) );
  NAND U45891 ( .A(n36825), .B(n36826), .Z(n36814) );
  NANDN U45892 ( .A(n36827), .B(n36828), .Z(n36826) );
  OR U45893 ( .A(n36829), .B(n36830), .Z(n36828) );
  NAND U45894 ( .A(n36830), .B(n36829), .Z(n36825) );
  AND U45895 ( .A(n36831), .B(n36832), .Z(n36816) );
  NANDN U45896 ( .A(n36833), .B(n36834), .Z(n36832) );
  NANDN U45897 ( .A(n36835), .B(n36836), .Z(n36834) );
  NANDN U45898 ( .A(n36836), .B(n36835), .Z(n36831) );
  XOR U45899 ( .A(n36830), .B(n36837), .Z(N62128) );
  XOR U45900 ( .A(n36827), .B(n36829), .Z(n36837) );
  XNOR U45901 ( .A(n36823), .B(n36838), .Z(n36829) );
  XNOR U45902 ( .A(n36821), .B(n36824), .Z(n36838) );
  NAND U45903 ( .A(n36839), .B(n36840), .Z(n36824) );
  NAND U45904 ( .A(n36841), .B(n36842), .Z(n36840) );
  OR U45905 ( .A(n36843), .B(n36844), .Z(n36841) );
  NANDN U45906 ( .A(n36845), .B(n36843), .Z(n36839) );
  IV U45907 ( .A(n36844), .Z(n36845) );
  NAND U45908 ( .A(n36846), .B(n36847), .Z(n36821) );
  NAND U45909 ( .A(n36848), .B(n36849), .Z(n36847) );
  NANDN U45910 ( .A(n36850), .B(n36851), .Z(n36848) );
  NANDN U45911 ( .A(n36851), .B(n36850), .Z(n36846) );
  AND U45912 ( .A(n36852), .B(n36853), .Z(n36823) );
  NAND U45913 ( .A(n36854), .B(n36855), .Z(n36853) );
  OR U45914 ( .A(n36856), .B(n36857), .Z(n36854) );
  NANDN U45915 ( .A(n36858), .B(n36856), .Z(n36852) );
  NAND U45916 ( .A(n36859), .B(n36860), .Z(n36827) );
  NANDN U45917 ( .A(n36861), .B(n36862), .Z(n36860) );
  OR U45918 ( .A(n36863), .B(n36864), .Z(n36862) );
  NANDN U45919 ( .A(n36865), .B(n36863), .Z(n36859) );
  IV U45920 ( .A(n36864), .Z(n36865) );
  XNOR U45921 ( .A(n36835), .B(n36866), .Z(n36830) );
  XNOR U45922 ( .A(n36833), .B(n36836), .Z(n36866) );
  NAND U45923 ( .A(n36867), .B(n36868), .Z(n36836) );
  NAND U45924 ( .A(n36869), .B(n36870), .Z(n36868) );
  OR U45925 ( .A(n36871), .B(n36872), .Z(n36869) );
  NANDN U45926 ( .A(n36873), .B(n36871), .Z(n36867) );
  IV U45927 ( .A(n36872), .Z(n36873) );
  NAND U45928 ( .A(n36874), .B(n36875), .Z(n36833) );
  NAND U45929 ( .A(n36876), .B(n36877), .Z(n36875) );
  NANDN U45930 ( .A(n36878), .B(n36879), .Z(n36876) );
  NANDN U45931 ( .A(n36879), .B(n36878), .Z(n36874) );
  AND U45932 ( .A(n36880), .B(n36881), .Z(n36835) );
  NAND U45933 ( .A(n36882), .B(n36883), .Z(n36881) );
  OR U45934 ( .A(n36884), .B(n36885), .Z(n36882) );
  NANDN U45935 ( .A(n36886), .B(n36884), .Z(n36880) );
  XNOR U45936 ( .A(n36861), .B(n36887), .Z(N62127) );
  XOR U45937 ( .A(n36863), .B(n36864), .Z(n36887) );
  XNOR U45938 ( .A(n36877), .B(n36888), .Z(n36864) );
  XOR U45939 ( .A(n36878), .B(n36879), .Z(n36888) );
  XOR U45940 ( .A(n36884), .B(n36889), .Z(n36879) );
  XOR U45941 ( .A(n36883), .B(n36886), .Z(n36889) );
  IV U45942 ( .A(n36885), .Z(n36886) );
  NAND U45943 ( .A(n36890), .B(n36891), .Z(n36885) );
  OR U45944 ( .A(n36892), .B(n36893), .Z(n36891) );
  OR U45945 ( .A(n36894), .B(n36895), .Z(n36890) );
  NAND U45946 ( .A(n36896), .B(n36897), .Z(n36883) );
  OR U45947 ( .A(n36898), .B(n36899), .Z(n36897) );
  OR U45948 ( .A(n36900), .B(n36901), .Z(n36896) );
  NOR U45949 ( .A(n36902), .B(n36903), .Z(n36884) );
  ANDN U45950 ( .B(n36904), .A(n36905), .Z(n36878) );
  XNOR U45951 ( .A(n36871), .B(n36906), .Z(n36877) );
  XNOR U45952 ( .A(n36870), .B(n36872), .Z(n36906) );
  NAND U45953 ( .A(n36907), .B(n36908), .Z(n36872) );
  OR U45954 ( .A(n36909), .B(n36910), .Z(n36908) );
  OR U45955 ( .A(n36911), .B(n36912), .Z(n36907) );
  NAND U45956 ( .A(n36913), .B(n36914), .Z(n36870) );
  OR U45957 ( .A(n36915), .B(n36916), .Z(n36914) );
  OR U45958 ( .A(n36917), .B(n36918), .Z(n36913) );
  ANDN U45959 ( .B(n36919), .A(n36920), .Z(n36871) );
  IV U45960 ( .A(n36921), .Z(n36919) );
  ANDN U45961 ( .B(n36922), .A(n36923), .Z(n36863) );
  XOR U45962 ( .A(n36849), .B(n36924), .Z(n36861) );
  XOR U45963 ( .A(n36850), .B(n36851), .Z(n36924) );
  XOR U45964 ( .A(n36856), .B(n36925), .Z(n36851) );
  XOR U45965 ( .A(n36855), .B(n36858), .Z(n36925) );
  IV U45966 ( .A(n36857), .Z(n36858) );
  NAND U45967 ( .A(n36926), .B(n36927), .Z(n36857) );
  OR U45968 ( .A(n36928), .B(n36929), .Z(n36927) );
  OR U45969 ( .A(n36930), .B(n36931), .Z(n36926) );
  NAND U45970 ( .A(n36932), .B(n36933), .Z(n36855) );
  OR U45971 ( .A(n36934), .B(n36935), .Z(n36933) );
  OR U45972 ( .A(n36936), .B(n36937), .Z(n36932) );
  NOR U45973 ( .A(n36938), .B(n36939), .Z(n36856) );
  ANDN U45974 ( .B(n36940), .A(n36941), .Z(n36850) );
  IV U45975 ( .A(n36942), .Z(n36940) );
  XNOR U45976 ( .A(n36843), .B(n36943), .Z(n36849) );
  XNOR U45977 ( .A(n36842), .B(n36844), .Z(n36943) );
  NAND U45978 ( .A(n36944), .B(n36945), .Z(n36844) );
  OR U45979 ( .A(n36946), .B(n36947), .Z(n36945) );
  OR U45980 ( .A(n36948), .B(n36949), .Z(n36944) );
  NAND U45981 ( .A(n36950), .B(n36951), .Z(n36842) );
  OR U45982 ( .A(n36952), .B(n36953), .Z(n36951) );
  OR U45983 ( .A(n36954), .B(n36955), .Z(n36950) );
  ANDN U45984 ( .B(n36956), .A(n36957), .Z(n36843) );
  IV U45985 ( .A(n36958), .Z(n36956) );
  XNOR U45986 ( .A(n36923), .B(n36922), .Z(N62126) );
  XOR U45987 ( .A(n36942), .B(n36941), .Z(n36922) );
  XNOR U45988 ( .A(n36957), .B(n36958), .Z(n36941) );
  XNOR U45989 ( .A(n36952), .B(n36953), .Z(n36958) );
  XNOR U45990 ( .A(n36954), .B(n36955), .Z(n36953) );
  XNOR U45991 ( .A(y[2845]), .B(x[2845]), .Z(n36955) );
  XNOR U45992 ( .A(y[2846]), .B(x[2846]), .Z(n36954) );
  XNOR U45993 ( .A(y[2844]), .B(x[2844]), .Z(n36952) );
  XNOR U45994 ( .A(n36946), .B(n36947), .Z(n36957) );
  XNOR U45995 ( .A(y[2841]), .B(x[2841]), .Z(n36947) );
  XNOR U45996 ( .A(n36948), .B(n36949), .Z(n36946) );
  XNOR U45997 ( .A(y[2842]), .B(x[2842]), .Z(n36949) );
  XNOR U45998 ( .A(y[2843]), .B(x[2843]), .Z(n36948) );
  XNOR U45999 ( .A(n36939), .B(n36938), .Z(n36942) );
  XNOR U46000 ( .A(n36934), .B(n36935), .Z(n36938) );
  XNOR U46001 ( .A(y[2838]), .B(x[2838]), .Z(n36935) );
  XNOR U46002 ( .A(n36936), .B(n36937), .Z(n36934) );
  XNOR U46003 ( .A(y[2839]), .B(x[2839]), .Z(n36937) );
  XNOR U46004 ( .A(y[2840]), .B(x[2840]), .Z(n36936) );
  XNOR U46005 ( .A(n36928), .B(n36929), .Z(n36939) );
  XNOR U46006 ( .A(y[2835]), .B(x[2835]), .Z(n36929) );
  XNOR U46007 ( .A(n36930), .B(n36931), .Z(n36928) );
  XNOR U46008 ( .A(y[2836]), .B(x[2836]), .Z(n36931) );
  XNOR U46009 ( .A(y[2837]), .B(x[2837]), .Z(n36930) );
  XOR U46010 ( .A(n36904), .B(n36905), .Z(n36923) );
  XNOR U46011 ( .A(n36920), .B(n36921), .Z(n36905) );
  XNOR U46012 ( .A(n36915), .B(n36916), .Z(n36921) );
  XNOR U46013 ( .A(n36917), .B(n36918), .Z(n36916) );
  XNOR U46014 ( .A(y[2833]), .B(x[2833]), .Z(n36918) );
  XNOR U46015 ( .A(y[2834]), .B(x[2834]), .Z(n36917) );
  XNOR U46016 ( .A(y[2832]), .B(x[2832]), .Z(n36915) );
  XNOR U46017 ( .A(n36909), .B(n36910), .Z(n36920) );
  XNOR U46018 ( .A(y[2829]), .B(x[2829]), .Z(n36910) );
  XNOR U46019 ( .A(n36911), .B(n36912), .Z(n36909) );
  XNOR U46020 ( .A(y[2830]), .B(x[2830]), .Z(n36912) );
  XNOR U46021 ( .A(y[2831]), .B(x[2831]), .Z(n36911) );
  XOR U46022 ( .A(n36903), .B(n36902), .Z(n36904) );
  XNOR U46023 ( .A(n36898), .B(n36899), .Z(n36902) );
  XNOR U46024 ( .A(y[2826]), .B(x[2826]), .Z(n36899) );
  XNOR U46025 ( .A(n36900), .B(n36901), .Z(n36898) );
  XNOR U46026 ( .A(y[2827]), .B(x[2827]), .Z(n36901) );
  XNOR U46027 ( .A(y[2828]), .B(x[2828]), .Z(n36900) );
  XNOR U46028 ( .A(n36892), .B(n36893), .Z(n36903) );
  XNOR U46029 ( .A(y[2823]), .B(x[2823]), .Z(n36893) );
  XNOR U46030 ( .A(n36894), .B(n36895), .Z(n36892) );
  XNOR U46031 ( .A(y[2824]), .B(x[2824]), .Z(n36895) );
  XNOR U46032 ( .A(y[2825]), .B(x[2825]), .Z(n36894) );
  NAND U46033 ( .A(n36959), .B(n36960), .Z(N62117) );
  NANDN U46034 ( .A(n36961), .B(n36962), .Z(n36960) );
  OR U46035 ( .A(n36963), .B(n36964), .Z(n36962) );
  NAND U46036 ( .A(n36963), .B(n36964), .Z(n36959) );
  XOR U46037 ( .A(n36963), .B(n36965), .Z(N62116) );
  XNOR U46038 ( .A(n36961), .B(n36964), .Z(n36965) );
  AND U46039 ( .A(n36966), .B(n36967), .Z(n36964) );
  NANDN U46040 ( .A(n36968), .B(n36969), .Z(n36967) );
  NANDN U46041 ( .A(n36970), .B(n36971), .Z(n36969) );
  NANDN U46042 ( .A(n36971), .B(n36970), .Z(n36966) );
  NAND U46043 ( .A(n36972), .B(n36973), .Z(n36961) );
  NANDN U46044 ( .A(n36974), .B(n36975), .Z(n36973) );
  OR U46045 ( .A(n36976), .B(n36977), .Z(n36975) );
  NAND U46046 ( .A(n36977), .B(n36976), .Z(n36972) );
  AND U46047 ( .A(n36978), .B(n36979), .Z(n36963) );
  NANDN U46048 ( .A(n36980), .B(n36981), .Z(n36979) );
  NANDN U46049 ( .A(n36982), .B(n36983), .Z(n36981) );
  NANDN U46050 ( .A(n36983), .B(n36982), .Z(n36978) );
  XOR U46051 ( .A(n36977), .B(n36984), .Z(N62115) );
  XOR U46052 ( .A(n36974), .B(n36976), .Z(n36984) );
  XNOR U46053 ( .A(n36970), .B(n36985), .Z(n36976) );
  XNOR U46054 ( .A(n36968), .B(n36971), .Z(n36985) );
  NAND U46055 ( .A(n36986), .B(n36987), .Z(n36971) );
  NAND U46056 ( .A(n36988), .B(n36989), .Z(n36987) );
  OR U46057 ( .A(n36990), .B(n36991), .Z(n36988) );
  NANDN U46058 ( .A(n36992), .B(n36990), .Z(n36986) );
  IV U46059 ( .A(n36991), .Z(n36992) );
  NAND U46060 ( .A(n36993), .B(n36994), .Z(n36968) );
  NAND U46061 ( .A(n36995), .B(n36996), .Z(n36994) );
  NANDN U46062 ( .A(n36997), .B(n36998), .Z(n36995) );
  NANDN U46063 ( .A(n36998), .B(n36997), .Z(n36993) );
  AND U46064 ( .A(n36999), .B(n37000), .Z(n36970) );
  NAND U46065 ( .A(n37001), .B(n37002), .Z(n37000) );
  OR U46066 ( .A(n37003), .B(n37004), .Z(n37001) );
  NANDN U46067 ( .A(n37005), .B(n37003), .Z(n36999) );
  NAND U46068 ( .A(n37006), .B(n37007), .Z(n36974) );
  NANDN U46069 ( .A(n37008), .B(n37009), .Z(n37007) );
  OR U46070 ( .A(n37010), .B(n37011), .Z(n37009) );
  NANDN U46071 ( .A(n37012), .B(n37010), .Z(n37006) );
  IV U46072 ( .A(n37011), .Z(n37012) );
  XNOR U46073 ( .A(n36982), .B(n37013), .Z(n36977) );
  XNOR U46074 ( .A(n36980), .B(n36983), .Z(n37013) );
  NAND U46075 ( .A(n37014), .B(n37015), .Z(n36983) );
  NAND U46076 ( .A(n37016), .B(n37017), .Z(n37015) );
  OR U46077 ( .A(n37018), .B(n37019), .Z(n37016) );
  NANDN U46078 ( .A(n37020), .B(n37018), .Z(n37014) );
  IV U46079 ( .A(n37019), .Z(n37020) );
  NAND U46080 ( .A(n37021), .B(n37022), .Z(n36980) );
  NAND U46081 ( .A(n37023), .B(n37024), .Z(n37022) );
  NANDN U46082 ( .A(n37025), .B(n37026), .Z(n37023) );
  NANDN U46083 ( .A(n37026), .B(n37025), .Z(n37021) );
  AND U46084 ( .A(n37027), .B(n37028), .Z(n36982) );
  NAND U46085 ( .A(n37029), .B(n37030), .Z(n37028) );
  OR U46086 ( .A(n37031), .B(n37032), .Z(n37029) );
  NANDN U46087 ( .A(n37033), .B(n37031), .Z(n37027) );
  XNOR U46088 ( .A(n37008), .B(n37034), .Z(N62114) );
  XOR U46089 ( .A(n37010), .B(n37011), .Z(n37034) );
  XNOR U46090 ( .A(n37024), .B(n37035), .Z(n37011) );
  XOR U46091 ( .A(n37025), .B(n37026), .Z(n37035) );
  XOR U46092 ( .A(n37031), .B(n37036), .Z(n37026) );
  XOR U46093 ( .A(n37030), .B(n37033), .Z(n37036) );
  IV U46094 ( .A(n37032), .Z(n37033) );
  NAND U46095 ( .A(n37037), .B(n37038), .Z(n37032) );
  OR U46096 ( .A(n37039), .B(n37040), .Z(n37038) );
  OR U46097 ( .A(n37041), .B(n37042), .Z(n37037) );
  NAND U46098 ( .A(n37043), .B(n37044), .Z(n37030) );
  OR U46099 ( .A(n37045), .B(n37046), .Z(n37044) );
  OR U46100 ( .A(n37047), .B(n37048), .Z(n37043) );
  NOR U46101 ( .A(n37049), .B(n37050), .Z(n37031) );
  ANDN U46102 ( .B(n37051), .A(n37052), .Z(n37025) );
  XNOR U46103 ( .A(n37018), .B(n37053), .Z(n37024) );
  XNOR U46104 ( .A(n37017), .B(n37019), .Z(n37053) );
  NAND U46105 ( .A(n37054), .B(n37055), .Z(n37019) );
  OR U46106 ( .A(n37056), .B(n37057), .Z(n37055) );
  OR U46107 ( .A(n37058), .B(n37059), .Z(n37054) );
  NAND U46108 ( .A(n37060), .B(n37061), .Z(n37017) );
  OR U46109 ( .A(n37062), .B(n37063), .Z(n37061) );
  OR U46110 ( .A(n37064), .B(n37065), .Z(n37060) );
  ANDN U46111 ( .B(n37066), .A(n37067), .Z(n37018) );
  IV U46112 ( .A(n37068), .Z(n37066) );
  ANDN U46113 ( .B(n37069), .A(n37070), .Z(n37010) );
  XOR U46114 ( .A(n36996), .B(n37071), .Z(n37008) );
  XOR U46115 ( .A(n36997), .B(n36998), .Z(n37071) );
  XOR U46116 ( .A(n37003), .B(n37072), .Z(n36998) );
  XOR U46117 ( .A(n37002), .B(n37005), .Z(n37072) );
  IV U46118 ( .A(n37004), .Z(n37005) );
  NAND U46119 ( .A(n37073), .B(n37074), .Z(n37004) );
  OR U46120 ( .A(n37075), .B(n37076), .Z(n37074) );
  OR U46121 ( .A(n37077), .B(n37078), .Z(n37073) );
  NAND U46122 ( .A(n37079), .B(n37080), .Z(n37002) );
  OR U46123 ( .A(n37081), .B(n37082), .Z(n37080) );
  OR U46124 ( .A(n37083), .B(n37084), .Z(n37079) );
  NOR U46125 ( .A(n37085), .B(n37086), .Z(n37003) );
  ANDN U46126 ( .B(n37087), .A(n37088), .Z(n36997) );
  IV U46127 ( .A(n37089), .Z(n37087) );
  XNOR U46128 ( .A(n36990), .B(n37090), .Z(n36996) );
  XNOR U46129 ( .A(n36989), .B(n36991), .Z(n37090) );
  NAND U46130 ( .A(n37091), .B(n37092), .Z(n36991) );
  OR U46131 ( .A(n37093), .B(n37094), .Z(n37092) );
  OR U46132 ( .A(n37095), .B(n37096), .Z(n37091) );
  NAND U46133 ( .A(n37097), .B(n37098), .Z(n36989) );
  OR U46134 ( .A(n37099), .B(n37100), .Z(n37098) );
  OR U46135 ( .A(n37101), .B(n37102), .Z(n37097) );
  ANDN U46136 ( .B(n37103), .A(n37104), .Z(n36990) );
  IV U46137 ( .A(n37105), .Z(n37103) );
  XNOR U46138 ( .A(n37070), .B(n37069), .Z(N62113) );
  XOR U46139 ( .A(n37089), .B(n37088), .Z(n37069) );
  XNOR U46140 ( .A(n37104), .B(n37105), .Z(n37088) );
  XNOR U46141 ( .A(n37099), .B(n37100), .Z(n37105) );
  XNOR U46142 ( .A(n37101), .B(n37102), .Z(n37100) );
  XNOR U46143 ( .A(y[2821]), .B(x[2821]), .Z(n37102) );
  XNOR U46144 ( .A(y[2822]), .B(x[2822]), .Z(n37101) );
  XNOR U46145 ( .A(y[2820]), .B(x[2820]), .Z(n37099) );
  XNOR U46146 ( .A(n37093), .B(n37094), .Z(n37104) );
  XNOR U46147 ( .A(y[2817]), .B(x[2817]), .Z(n37094) );
  XNOR U46148 ( .A(n37095), .B(n37096), .Z(n37093) );
  XNOR U46149 ( .A(y[2818]), .B(x[2818]), .Z(n37096) );
  XNOR U46150 ( .A(y[2819]), .B(x[2819]), .Z(n37095) );
  XNOR U46151 ( .A(n37086), .B(n37085), .Z(n37089) );
  XNOR U46152 ( .A(n37081), .B(n37082), .Z(n37085) );
  XNOR U46153 ( .A(y[2814]), .B(x[2814]), .Z(n37082) );
  XNOR U46154 ( .A(n37083), .B(n37084), .Z(n37081) );
  XNOR U46155 ( .A(y[2815]), .B(x[2815]), .Z(n37084) );
  XNOR U46156 ( .A(y[2816]), .B(x[2816]), .Z(n37083) );
  XNOR U46157 ( .A(n37075), .B(n37076), .Z(n37086) );
  XNOR U46158 ( .A(y[2811]), .B(x[2811]), .Z(n37076) );
  XNOR U46159 ( .A(n37077), .B(n37078), .Z(n37075) );
  XNOR U46160 ( .A(y[2812]), .B(x[2812]), .Z(n37078) );
  XNOR U46161 ( .A(y[2813]), .B(x[2813]), .Z(n37077) );
  XOR U46162 ( .A(n37051), .B(n37052), .Z(n37070) );
  XNOR U46163 ( .A(n37067), .B(n37068), .Z(n37052) );
  XNOR U46164 ( .A(n37062), .B(n37063), .Z(n37068) );
  XNOR U46165 ( .A(n37064), .B(n37065), .Z(n37063) );
  XNOR U46166 ( .A(y[2809]), .B(x[2809]), .Z(n37065) );
  XNOR U46167 ( .A(y[2810]), .B(x[2810]), .Z(n37064) );
  XNOR U46168 ( .A(y[2808]), .B(x[2808]), .Z(n37062) );
  XNOR U46169 ( .A(n37056), .B(n37057), .Z(n37067) );
  XNOR U46170 ( .A(y[2805]), .B(x[2805]), .Z(n37057) );
  XNOR U46171 ( .A(n37058), .B(n37059), .Z(n37056) );
  XNOR U46172 ( .A(y[2806]), .B(x[2806]), .Z(n37059) );
  XNOR U46173 ( .A(y[2807]), .B(x[2807]), .Z(n37058) );
  XOR U46174 ( .A(n37050), .B(n37049), .Z(n37051) );
  XNOR U46175 ( .A(n37045), .B(n37046), .Z(n37049) );
  XNOR U46176 ( .A(y[2802]), .B(x[2802]), .Z(n37046) );
  XNOR U46177 ( .A(n37047), .B(n37048), .Z(n37045) );
  XNOR U46178 ( .A(y[2803]), .B(x[2803]), .Z(n37048) );
  XNOR U46179 ( .A(y[2804]), .B(x[2804]), .Z(n37047) );
  XNOR U46180 ( .A(n37039), .B(n37040), .Z(n37050) );
  XNOR U46181 ( .A(y[2799]), .B(x[2799]), .Z(n37040) );
  XNOR U46182 ( .A(n37041), .B(n37042), .Z(n37039) );
  XNOR U46183 ( .A(y[2800]), .B(x[2800]), .Z(n37042) );
  XNOR U46184 ( .A(y[2801]), .B(x[2801]), .Z(n37041) );
  NAND U46185 ( .A(n37106), .B(n37107), .Z(N62104) );
  NANDN U46186 ( .A(n37108), .B(n37109), .Z(n37107) );
  OR U46187 ( .A(n37110), .B(n37111), .Z(n37109) );
  NAND U46188 ( .A(n37110), .B(n37111), .Z(n37106) );
  XOR U46189 ( .A(n37110), .B(n37112), .Z(N62103) );
  XNOR U46190 ( .A(n37108), .B(n37111), .Z(n37112) );
  AND U46191 ( .A(n37113), .B(n37114), .Z(n37111) );
  NANDN U46192 ( .A(n37115), .B(n37116), .Z(n37114) );
  NANDN U46193 ( .A(n37117), .B(n37118), .Z(n37116) );
  NANDN U46194 ( .A(n37118), .B(n37117), .Z(n37113) );
  NAND U46195 ( .A(n37119), .B(n37120), .Z(n37108) );
  NANDN U46196 ( .A(n37121), .B(n37122), .Z(n37120) );
  OR U46197 ( .A(n37123), .B(n37124), .Z(n37122) );
  NAND U46198 ( .A(n37124), .B(n37123), .Z(n37119) );
  AND U46199 ( .A(n37125), .B(n37126), .Z(n37110) );
  NANDN U46200 ( .A(n37127), .B(n37128), .Z(n37126) );
  NANDN U46201 ( .A(n37129), .B(n37130), .Z(n37128) );
  NANDN U46202 ( .A(n37130), .B(n37129), .Z(n37125) );
  XOR U46203 ( .A(n37124), .B(n37131), .Z(N62102) );
  XOR U46204 ( .A(n37121), .B(n37123), .Z(n37131) );
  XNOR U46205 ( .A(n37117), .B(n37132), .Z(n37123) );
  XNOR U46206 ( .A(n37115), .B(n37118), .Z(n37132) );
  NAND U46207 ( .A(n37133), .B(n37134), .Z(n37118) );
  NAND U46208 ( .A(n37135), .B(n37136), .Z(n37134) );
  OR U46209 ( .A(n37137), .B(n37138), .Z(n37135) );
  NANDN U46210 ( .A(n37139), .B(n37137), .Z(n37133) );
  IV U46211 ( .A(n37138), .Z(n37139) );
  NAND U46212 ( .A(n37140), .B(n37141), .Z(n37115) );
  NAND U46213 ( .A(n37142), .B(n37143), .Z(n37141) );
  NANDN U46214 ( .A(n37144), .B(n37145), .Z(n37142) );
  NANDN U46215 ( .A(n37145), .B(n37144), .Z(n37140) );
  AND U46216 ( .A(n37146), .B(n37147), .Z(n37117) );
  NAND U46217 ( .A(n37148), .B(n37149), .Z(n37147) );
  OR U46218 ( .A(n37150), .B(n37151), .Z(n37148) );
  NANDN U46219 ( .A(n37152), .B(n37150), .Z(n37146) );
  NAND U46220 ( .A(n37153), .B(n37154), .Z(n37121) );
  NANDN U46221 ( .A(n37155), .B(n37156), .Z(n37154) );
  OR U46222 ( .A(n37157), .B(n37158), .Z(n37156) );
  NANDN U46223 ( .A(n37159), .B(n37157), .Z(n37153) );
  IV U46224 ( .A(n37158), .Z(n37159) );
  XNOR U46225 ( .A(n37129), .B(n37160), .Z(n37124) );
  XNOR U46226 ( .A(n37127), .B(n37130), .Z(n37160) );
  NAND U46227 ( .A(n37161), .B(n37162), .Z(n37130) );
  NAND U46228 ( .A(n37163), .B(n37164), .Z(n37162) );
  OR U46229 ( .A(n37165), .B(n37166), .Z(n37163) );
  NANDN U46230 ( .A(n37167), .B(n37165), .Z(n37161) );
  IV U46231 ( .A(n37166), .Z(n37167) );
  NAND U46232 ( .A(n37168), .B(n37169), .Z(n37127) );
  NAND U46233 ( .A(n37170), .B(n37171), .Z(n37169) );
  NANDN U46234 ( .A(n37172), .B(n37173), .Z(n37170) );
  NANDN U46235 ( .A(n37173), .B(n37172), .Z(n37168) );
  AND U46236 ( .A(n37174), .B(n37175), .Z(n37129) );
  NAND U46237 ( .A(n37176), .B(n37177), .Z(n37175) );
  OR U46238 ( .A(n37178), .B(n37179), .Z(n37176) );
  NANDN U46239 ( .A(n37180), .B(n37178), .Z(n37174) );
  XNOR U46240 ( .A(n37155), .B(n37181), .Z(N62101) );
  XOR U46241 ( .A(n37157), .B(n37158), .Z(n37181) );
  XNOR U46242 ( .A(n37171), .B(n37182), .Z(n37158) );
  XOR U46243 ( .A(n37172), .B(n37173), .Z(n37182) );
  XOR U46244 ( .A(n37178), .B(n37183), .Z(n37173) );
  XOR U46245 ( .A(n37177), .B(n37180), .Z(n37183) );
  IV U46246 ( .A(n37179), .Z(n37180) );
  NAND U46247 ( .A(n37184), .B(n37185), .Z(n37179) );
  OR U46248 ( .A(n37186), .B(n37187), .Z(n37185) );
  OR U46249 ( .A(n37188), .B(n37189), .Z(n37184) );
  NAND U46250 ( .A(n37190), .B(n37191), .Z(n37177) );
  OR U46251 ( .A(n37192), .B(n37193), .Z(n37191) );
  OR U46252 ( .A(n37194), .B(n37195), .Z(n37190) );
  NOR U46253 ( .A(n37196), .B(n37197), .Z(n37178) );
  ANDN U46254 ( .B(n37198), .A(n37199), .Z(n37172) );
  XNOR U46255 ( .A(n37165), .B(n37200), .Z(n37171) );
  XNOR U46256 ( .A(n37164), .B(n37166), .Z(n37200) );
  NAND U46257 ( .A(n37201), .B(n37202), .Z(n37166) );
  OR U46258 ( .A(n37203), .B(n37204), .Z(n37202) );
  OR U46259 ( .A(n37205), .B(n37206), .Z(n37201) );
  NAND U46260 ( .A(n37207), .B(n37208), .Z(n37164) );
  OR U46261 ( .A(n37209), .B(n37210), .Z(n37208) );
  OR U46262 ( .A(n37211), .B(n37212), .Z(n37207) );
  ANDN U46263 ( .B(n37213), .A(n37214), .Z(n37165) );
  IV U46264 ( .A(n37215), .Z(n37213) );
  ANDN U46265 ( .B(n37216), .A(n37217), .Z(n37157) );
  XOR U46266 ( .A(n37143), .B(n37218), .Z(n37155) );
  XOR U46267 ( .A(n37144), .B(n37145), .Z(n37218) );
  XOR U46268 ( .A(n37150), .B(n37219), .Z(n37145) );
  XOR U46269 ( .A(n37149), .B(n37152), .Z(n37219) );
  IV U46270 ( .A(n37151), .Z(n37152) );
  NAND U46271 ( .A(n37220), .B(n37221), .Z(n37151) );
  OR U46272 ( .A(n37222), .B(n37223), .Z(n37221) );
  OR U46273 ( .A(n37224), .B(n37225), .Z(n37220) );
  NAND U46274 ( .A(n37226), .B(n37227), .Z(n37149) );
  OR U46275 ( .A(n37228), .B(n37229), .Z(n37227) );
  OR U46276 ( .A(n37230), .B(n37231), .Z(n37226) );
  NOR U46277 ( .A(n37232), .B(n37233), .Z(n37150) );
  ANDN U46278 ( .B(n37234), .A(n37235), .Z(n37144) );
  IV U46279 ( .A(n37236), .Z(n37234) );
  XNOR U46280 ( .A(n37137), .B(n37237), .Z(n37143) );
  XNOR U46281 ( .A(n37136), .B(n37138), .Z(n37237) );
  NAND U46282 ( .A(n37238), .B(n37239), .Z(n37138) );
  OR U46283 ( .A(n37240), .B(n37241), .Z(n37239) );
  OR U46284 ( .A(n37242), .B(n37243), .Z(n37238) );
  NAND U46285 ( .A(n37244), .B(n37245), .Z(n37136) );
  OR U46286 ( .A(n37246), .B(n37247), .Z(n37245) );
  OR U46287 ( .A(n37248), .B(n37249), .Z(n37244) );
  ANDN U46288 ( .B(n37250), .A(n37251), .Z(n37137) );
  IV U46289 ( .A(n37252), .Z(n37250) );
  XNOR U46290 ( .A(n37217), .B(n37216), .Z(N62100) );
  XOR U46291 ( .A(n37236), .B(n37235), .Z(n37216) );
  XNOR U46292 ( .A(n37251), .B(n37252), .Z(n37235) );
  XNOR U46293 ( .A(n37246), .B(n37247), .Z(n37252) );
  XNOR U46294 ( .A(n37248), .B(n37249), .Z(n37247) );
  XNOR U46295 ( .A(y[2797]), .B(x[2797]), .Z(n37249) );
  XNOR U46296 ( .A(y[2798]), .B(x[2798]), .Z(n37248) );
  XNOR U46297 ( .A(y[2796]), .B(x[2796]), .Z(n37246) );
  XNOR U46298 ( .A(n37240), .B(n37241), .Z(n37251) );
  XNOR U46299 ( .A(y[2793]), .B(x[2793]), .Z(n37241) );
  XNOR U46300 ( .A(n37242), .B(n37243), .Z(n37240) );
  XNOR U46301 ( .A(y[2794]), .B(x[2794]), .Z(n37243) );
  XNOR U46302 ( .A(y[2795]), .B(x[2795]), .Z(n37242) );
  XNOR U46303 ( .A(n37233), .B(n37232), .Z(n37236) );
  XNOR U46304 ( .A(n37228), .B(n37229), .Z(n37232) );
  XNOR U46305 ( .A(y[2790]), .B(x[2790]), .Z(n37229) );
  XNOR U46306 ( .A(n37230), .B(n37231), .Z(n37228) );
  XNOR U46307 ( .A(y[2791]), .B(x[2791]), .Z(n37231) );
  XNOR U46308 ( .A(y[2792]), .B(x[2792]), .Z(n37230) );
  XNOR U46309 ( .A(n37222), .B(n37223), .Z(n37233) );
  XNOR U46310 ( .A(y[2787]), .B(x[2787]), .Z(n37223) );
  XNOR U46311 ( .A(n37224), .B(n37225), .Z(n37222) );
  XNOR U46312 ( .A(y[2788]), .B(x[2788]), .Z(n37225) );
  XNOR U46313 ( .A(y[2789]), .B(x[2789]), .Z(n37224) );
  XOR U46314 ( .A(n37198), .B(n37199), .Z(n37217) );
  XNOR U46315 ( .A(n37214), .B(n37215), .Z(n37199) );
  XNOR U46316 ( .A(n37209), .B(n37210), .Z(n37215) );
  XNOR U46317 ( .A(n37211), .B(n37212), .Z(n37210) );
  XNOR U46318 ( .A(y[2785]), .B(x[2785]), .Z(n37212) );
  XNOR U46319 ( .A(y[2786]), .B(x[2786]), .Z(n37211) );
  XNOR U46320 ( .A(y[2784]), .B(x[2784]), .Z(n37209) );
  XNOR U46321 ( .A(n37203), .B(n37204), .Z(n37214) );
  XNOR U46322 ( .A(y[2781]), .B(x[2781]), .Z(n37204) );
  XNOR U46323 ( .A(n37205), .B(n37206), .Z(n37203) );
  XNOR U46324 ( .A(y[2782]), .B(x[2782]), .Z(n37206) );
  XNOR U46325 ( .A(y[2783]), .B(x[2783]), .Z(n37205) );
  XOR U46326 ( .A(n37197), .B(n37196), .Z(n37198) );
  XNOR U46327 ( .A(n37192), .B(n37193), .Z(n37196) );
  XNOR U46328 ( .A(y[2778]), .B(x[2778]), .Z(n37193) );
  XNOR U46329 ( .A(n37194), .B(n37195), .Z(n37192) );
  XNOR U46330 ( .A(y[2779]), .B(x[2779]), .Z(n37195) );
  XNOR U46331 ( .A(y[2780]), .B(x[2780]), .Z(n37194) );
  XNOR U46332 ( .A(n37186), .B(n37187), .Z(n37197) );
  XNOR U46333 ( .A(y[2775]), .B(x[2775]), .Z(n37187) );
  XNOR U46334 ( .A(n37188), .B(n37189), .Z(n37186) );
  XNOR U46335 ( .A(y[2776]), .B(x[2776]), .Z(n37189) );
  XNOR U46336 ( .A(y[2777]), .B(x[2777]), .Z(n37188) );
  NAND U46337 ( .A(n37253), .B(n37254), .Z(N62091) );
  NANDN U46338 ( .A(n37255), .B(n37256), .Z(n37254) );
  OR U46339 ( .A(n37257), .B(n37258), .Z(n37256) );
  NAND U46340 ( .A(n37257), .B(n37258), .Z(n37253) );
  XOR U46341 ( .A(n37257), .B(n37259), .Z(N62090) );
  XNOR U46342 ( .A(n37255), .B(n37258), .Z(n37259) );
  AND U46343 ( .A(n37260), .B(n37261), .Z(n37258) );
  NANDN U46344 ( .A(n37262), .B(n37263), .Z(n37261) );
  NANDN U46345 ( .A(n37264), .B(n37265), .Z(n37263) );
  NANDN U46346 ( .A(n37265), .B(n37264), .Z(n37260) );
  NAND U46347 ( .A(n37266), .B(n37267), .Z(n37255) );
  NANDN U46348 ( .A(n37268), .B(n37269), .Z(n37267) );
  OR U46349 ( .A(n37270), .B(n37271), .Z(n37269) );
  NAND U46350 ( .A(n37271), .B(n37270), .Z(n37266) );
  AND U46351 ( .A(n37272), .B(n37273), .Z(n37257) );
  NANDN U46352 ( .A(n37274), .B(n37275), .Z(n37273) );
  NANDN U46353 ( .A(n37276), .B(n37277), .Z(n37275) );
  NANDN U46354 ( .A(n37277), .B(n37276), .Z(n37272) );
  XOR U46355 ( .A(n37271), .B(n37278), .Z(N62089) );
  XOR U46356 ( .A(n37268), .B(n37270), .Z(n37278) );
  XNOR U46357 ( .A(n37264), .B(n37279), .Z(n37270) );
  XNOR U46358 ( .A(n37262), .B(n37265), .Z(n37279) );
  NAND U46359 ( .A(n37280), .B(n37281), .Z(n37265) );
  NAND U46360 ( .A(n37282), .B(n37283), .Z(n37281) );
  OR U46361 ( .A(n37284), .B(n37285), .Z(n37282) );
  NANDN U46362 ( .A(n37286), .B(n37284), .Z(n37280) );
  IV U46363 ( .A(n37285), .Z(n37286) );
  NAND U46364 ( .A(n37287), .B(n37288), .Z(n37262) );
  NAND U46365 ( .A(n37289), .B(n37290), .Z(n37288) );
  NANDN U46366 ( .A(n37291), .B(n37292), .Z(n37289) );
  NANDN U46367 ( .A(n37292), .B(n37291), .Z(n37287) );
  AND U46368 ( .A(n37293), .B(n37294), .Z(n37264) );
  NAND U46369 ( .A(n37295), .B(n37296), .Z(n37294) );
  OR U46370 ( .A(n37297), .B(n37298), .Z(n37295) );
  NANDN U46371 ( .A(n37299), .B(n37297), .Z(n37293) );
  NAND U46372 ( .A(n37300), .B(n37301), .Z(n37268) );
  NANDN U46373 ( .A(n37302), .B(n37303), .Z(n37301) );
  OR U46374 ( .A(n37304), .B(n37305), .Z(n37303) );
  NANDN U46375 ( .A(n37306), .B(n37304), .Z(n37300) );
  IV U46376 ( .A(n37305), .Z(n37306) );
  XNOR U46377 ( .A(n37276), .B(n37307), .Z(n37271) );
  XNOR U46378 ( .A(n37274), .B(n37277), .Z(n37307) );
  NAND U46379 ( .A(n37308), .B(n37309), .Z(n37277) );
  NAND U46380 ( .A(n37310), .B(n37311), .Z(n37309) );
  OR U46381 ( .A(n37312), .B(n37313), .Z(n37310) );
  NANDN U46382 ( .A(n37314), .B(n37312), .Z(n37308) );
  IV U46383 ( .A(n37313), .Z(n37314) );
  NAND U46384 ( .A(n37315), .B(n37316), .Z(n37274) );
  NAND U46385 ( .A(n37317), .B(n37318), .Z(n37316) );
  NANDN U46386 ( .A(n37319), .B(n37320), .Z(n37317) );
  NANDN U46387 ( .A(n37320), .B(n37319), .Z(n37315) );
  AND U46388 ( .A(n37321), .B(n37322), .Z(n37276) );
  NAND U46389 ( .A(n37323), .B(n37324), .Z(n37322) );
  OR U46390 ( .A(n37325), .B(n37326), .Z(n37323) );
  NANDN U46391 ( .A(n37327), .B(n37325), .Z(n37321) );
  XNOR U46392 ( .A(n37302), .B(n37328), .Z(N62088) );
  XOR U46393 ( .A(n37304), .B(n37305), .Z(n37328) );
  XNOR U46394 ( .A(n37318), .B(n37329), .Z(n37305) );
  XOR U46395 ( .A(n37319), .B(n37320), .Z(n37329) );
  XOR U46396 ( .A(n37325), .B(n37330), .Z(n37320) );
  XOR U46397 ( .A(n37324), .B(n37327), .Z(n37330) );
  IV U46398 ( .A(n37326), .Z(n37327) );
  NAND U46399 ( .A(n37331), .B(n37332), .Z(n37326) );
  OR U46400 ( .A(n37333), .B(n37334), .Z(n37332) );
  OR U46401 ( .A(n37335), .B(n37336), .Z(n37331) );
  NAND U46402 ( .A(n37337), .B(n37338), .Z(n37324) );
  OR U46403 ( .A(n37339), .B(n37340), .Z(n37338) );
  OR U46404 ( .A(n37341), .B(n37342), .Z(n37337) );
  NOR U46405 ( .A(n37343), .B(n37344), .Z(n37325) );
  ANDN U46406 ( .B(n37345), .A(n37346), .Z(n37319) );
  XNOR U46407 ( .A(n37312), .B(n37347), .Z(n37318) );
  XNOR U46408 ( .A(n37311), .B(n37313), .Z(n37347) );
  NAND U46409 ( .A(n37348), .B(n37349), .Z(n37313) );
  OR U46410 ( .A(n37350), .B(n37351), .Z(n37349) );
  OR U46411 ( .A(n37352), .B(n37353), .Z(n37348) );
  NAND U46412 ( .A(n37354), .B(n37355), .Z(n37311) );
  OR U46413 ( .A(n37356), .B(n37357), .Z(n37355) );
  OR U46414 ( .A(n37358), .B(n37359), .Z(n37354) );
  ANDN U46415 ( .B(n37360), .A(n37361), .Z(n37312) );
  IV U46416 ( .A(n37362), .Z(n37360) );
  ANDN U46417 ( .B(n37363), .A(n37364), .Z(n37304) );
  XOR U46418 ( .A(n37290), .B(n37365), .Z(n37302) );
  XOR U46419 ( .A(n37291), .B(n37292), .Z(n37365) );
  XOR U46420 ( .A(n37297), .B(n37366), .Z(n37292) );
  XOR U46421 ( .A(n37296), .B(n37299), .Z(n37366) );
  IV U46422 ( .A(n37298), .Z(n37299) );
  NAND U46423 ( .A(n37367), .B(n37368), .Z(n37298) );
  OR U46424 ( .A(n37369), .B(n37370), .Z(n37368) );
  OR U46425 ( .A(n37371), .B(n37372), .Z(n37367) );
  NAND U46426 ( .A(n37373), .B(n37374), .Z(n37296) );
  OR U46427 ( .A(n37375), .B(n37376), .Z(n37374) );
  OR U46428 ( .A(n37377), .B(n37378), .Z(n37373) );
  NOR U46429 ( .A(n37379), .B(n37380), .Z(n37297) );
  ANDN U46430 ( .B(n37381), .A(n37382), .Z(n37291) );
  IV U46431 ( .A(n37383), .Z(n37381) );
  XNOR U46432 ( .A(n37284), .B(n37384), .Z(n37290) );
  XNOR U46433 ( .A(n37283), .B(n37285), .Z(n37384) );
  NAND U46434 ( .A(n37385), .B(n37386), .Z(n37285) );
  OR U46435 ( .A(n37387), .B(n37388), .Z(n37386) );
  OR U46436 ( .A(n37389), .B(n37390), .Z(n37385) );
  NAND U46437 ( .A(n37391), .B(n37392), .Z(n37283) );
  OR U46438 ( .A(n37393), .B(n37394), .Z(n37392) );
  OR U46439 ( .A(n37395), .B(n37396), .Z(n37391) );
  ANDN U46440 ( .B(n37397), .A(n37398), .Z(n37284) );
  IV U46441 ( .A(n37399), .Z(n37397) );
  XNOR U46442 ( .A(n37364), .B(n37363), .Z(N62087) );
  XOR U46443 ( .A(n37383), .B(n37382), .Z(n37363) );
  XNOR U46444 ( .A(n37398), .B(n37399), .Z(n37382) );
  XNOR U46445 ( .A(n37393), .B(n37394), .Z(n37399) );
  XNOR U46446 ( .A(n37395), .B(n37396), .Z(n37394) );
  XNOR U46447 ( .A(y[2773]), .B(x[2773]), .Z(n37396) );
  XNOR U46448 ( .A(y[2774]), .B(x[2774]), .Z(n37395) );
  XNOR U46449 ( .A(y[2772]), .B(x[2772]), .Z(n37393) );
  XNOR U46450 ( .A(n37387), .B(n37388), .Z(n37398) );
  XNOR U46451 ( .A(y[2769]), .B(x[2769]), .Z(n37388) );
  XNOR U46452 ( .A(n37389), .B(n37390), .Z(n37387) );
  XNOR U46453 ( .A(y[2770]), .B(x[2770]), .Z(n37390) );
  XNOR U46454 ( .A(y[2771]), .B(x[2771]), .Z(n37389) );
  XNOR U46455 ( .A(n37380), .B(n37379), .Z(n37383) );
  XNOR U46456 ( .A(n37375), .B(n37376), .Z(n37379) );
  XNOR U46457 ( .A(y[2766]), .B(x[2766]), .Z(n37376) );
  XNOR U46458 ( .A(n37377), .B(n37378), .Z(n37375) );
  XNOR U46459 ( .A(y[2767]), .B(x[2767]), .Z(n37378) );
  XNOR U46460 ( .A(y[2768]), .B(x[2768]), .Z(n37377) );
  XNOR U46461 ( .A(n37369), .B(n37370), .Z(n37380) );
  XNOR U46462 ( .A(y[2763]), .B(x[2763]), .Z(n37370) );
  XNOR U46463 ( .A(n37371), .B(n37372), .Z(n37369) );
  XNOR U46464 ( .A(y[2764]), .B(x[2764]), .Z(n37372) );
  XNOR U46465 ( .A(y[2765]), .B(x[2765]), .Z(n37371) );
  XOR U46466 ( .A(n37345), .B(n37346), .Z(n37364) );
  XNOR U46467 ( .A(n37361), .B(n37362), .Z(n37346) );
  XNOR U46468 ( .A(n37356), .B(n37357), .Z(n37362) );
  XNOR U46469 ( .A(n37358), .B(n37359), .Z(n37357) );
  XNOR U46470 ( .A(y[2761]), .B(x[2761]), .Z(n37359) );
  XNOR U46471 ( .A(y[2762]), .B(x[2762]), .Z(n37358) );
  XNOR U46472 ( .A(y[2760]), .B(x[2760]), .Z(n37356) );
  XNOR U46473 ( .A(n37350), .B(n37351), .Z(n37361) );
  XNOR U46474 ( .A(y[2757]), .B(x[2757]), .Z(n37351) );
  XNOR U46475 ( .A(n37352), .B(n37353), .Z(n37350) );
  XNOR U46476 ( .A(y[2758]), .B(x[2758]), .Z(n37353) );
  XNOR U46477 ( .A(y[2759]), .B(x[2759]), .Z(n37352) );
  XOR U46478 ( .A(n37344), .B(n37343), .Z(n37345) );
  XNOR U46479 ( .A(n37339), .B(n37340), .Z(n37343) );
  XNOR U46480 ( .A(y[2754]), .B(x[2754]), .Z(n37340) );
  XNOR U46481 ( .A(n37341), .B(n37342), .Z(n37339) );
  XNOR U46482 ( .A(y[2755]), .B(x[2755]), .Z(n37342) );
  XNOR U46483 ( .A(y[2756]), .B(x[2756]), .Z(n37341) );
  XNOR U46484 ( .A(n37333), .B(n37334), .Z(n37344) );
  XNOR U46485 ( .A(y[2751]), .B(x[2751]), .Z(n37334) );
  XNOR U46486 ( .A(n37335), .B(n37336), .Z(n37333) );
  XNOR U46487 ( .A(y[2752]), .B(x[2752]), .Z(n37336) );
  XNOR U46488 ( .A(y[2753]), .B(x[2753]), .Z(n37335) );
  NAND U46489 ( .A(n37400), .B(n37401), .Z(N62078) );
  NANDN U46490 ( .A(n37402), .B(n37403), .Z(n37401) );
  OR U46491 ( .A(n37404), .B(n37405), .Z(n37403) );
  NAND U46492 ( .A(n37404), .B(n37405), .Z(n37400) );
  XOR U46493 ( .A(n37404), .B(n37406), .Z(N62077) );
  XNOR U46494 ( .A(n37402), .B(n37405), .Z(n37406) );
  AND U46495 ( .A(n37407), .B(n37408), .Z(n37405) );
  NANDN U46496 ( .A(n37409), .B(n37410), .Z(n37408) );
  NANDN U46497 ( .A(n37411), .B(n37412), .Z(n37410) );
  NANDN U46498 ( .A(n37412), .B(n37411), .Z(n37407) );
  NAND U46499 ( .A(n37413), .B(n37414), .Z(n37402) );
  NANDN U46500 ( .A(n37415), .B(n37416), .Z(n37414) );
  OR U46501 ( .A(n37417), .B(n37418), .Z(n37416) );
  NAND U46502 ( .A(n37418), .B(n37417), .Z(n37413) );
  AND U46503 ( .A(n37419), .B(n37420), .Z(n37404) );
  NANDN U46504 ( .A(n37421), .B(n37422), .Z(n37420) );
  NANDN U46505 ( .A(n37423), .B(n37424), .Z(n37422) );
  NANDN U46506 ( .A(n37424), .B(n37423), .Z(n37419) );
  XOR U46507 ( .A(n37418), .B(n37425), .Z(N62076) );
  XOR U46508 ( .A(n37415), .B(n37417), .Z(n37425) );
  XNOR U46509 ( .A(n37411), .B(n37426), .Z(n37417) );
  XNOR U46510 ( .A(n37409), .B(n37412), .Z(n37426) );
  NAND U46511 ( .A(n37427), .B(n37428), .Z(n37412) );
  NAND U46512 ( .A(n37429), .B(n37430), .Z(n37428) );
  OR U46513 ( .A(n37431), .B(n37432), .Z(n37429) );
  NANDN U46514 ( .A(n37433), .B(n37431), .Z(n37427) );
  IV U46515 ( .A(n37432), .Z(n37433) );
  NAND U46516 ( .A(n37434), .B(n37435), .Z(n37409) );
  NAND U46517 ( .A(n37436), .B(n37437), .Z(n37435) );
  NANDN U46518 ( .A(n37438), .B(n37439), .Z(n37436) );
  NANDN U46519 ( .A(n37439), .B(n37438), .Z(n37434) );
  AND U46520 ( .A(n37440), .B(n37441), .Z(n37411) );
  NAND U46521 ( .A(n37442), .B(n37443), .Z(n37441) );
  OR U46522 ( .A(n37444), .B(n37445), .Z(n37442) );
  NANDN U46523 ( .A(n37446), .B(n37444), .Z(n37440) );
  NAND U46524 ( .A(n37447), .B(n37448), .Z(n37415) );
  NANDN U46525 ( .A(n37449), .B(n37450), .Z(n37448) );
  OR U46526 ( .A(n37451), .B(n37452), .Z(n37450) );
  NANDN U46527 ( .A(n37453), .B(n37451), .Z(n37447) );
  IV U46528 ( .A(n37452), .Z(n37453) );
  XNOR U46529 ( .A(n37423), .B(n37454), .Z(n37418) );
  XNOR U46530 ( .A(n37421), .B(n37424), .Z(n37454) );
  NAND U46531 ( .A(n37455), .B(n37456), .Z(n37424) );
  NAND U46532 ( .A(n37457), .B(n37458), .Z(n37456) );
  OR U46533 ( .A(n37459), .B(n37460), .Z(n37457) );
  NANDN U46534 ( .A(n37461), .B(n37459), .Z(n37455) );
  IV U46535 ( .A(n37460), .Z(n37461) );
  NAND U46536 ( .A(n37462), .B(n37463), .Z(n37421) );
  NAND U46537 ( .A(n37464), .B(n37465), .Z(n37463) );
  NANDN U46538 ( .A(n37466), .B(n37467), .Z(n37464) );
  NANDN U46539 ( .A(n37467), .B(n37466), .Z(n37462) );
  AND U46540 ( .A(n37468), .B(n37469), .Z(n37423) );
  NAND U46541 ( .A(n37470), .B(n37471), .Z(n37469) );
  OR U46542 ( .A(n37472), .B(n37473), .Z(n37470) );
  NANDN U46543 ( .A(n37474), .B(n37472), .Z(n37468) );
  XNOR U46544 ( .A(n37449), .B(n37475), .Z(N62075) );
  XOR U46545 ( .A(n37451), .B(n37452), .Z(n37475) );
  XNOR U46546 ( .A(n37465), .B(n37476), .Z(n37452) );
  XOR U46547 ( .A(n37466), .B(n37467), .Z(n37476) );
  XOR U46548 ( .A(n37472), .B(n37477), .Z(n37467) );
  XOR U46549 ( .A(n37471), .B(n37474), .Z(n37477) );
  IV U46550 ( .A(n37473), .Z(n37474) );
  NAND U46551 ( .A(n37478), .B(n37479), .Z(n37473) );
  OR U46552 ( .A(n37480), .B(n37481), .Z(n37479) );
  OR U46553 ( .A(n37482), .B(n37483), .Z(n37478) );
  NAND U46554 ( .A(n37484), .B(n37485), .Z(n37471) );
  OR U46555 ( .A(n37486), .B(n37487), .Z(n37485) );
  OR U46556 ( .A(n37488), .B(n37489), .Z(n37484) );
  NOR U46557 ( .A(n37490), .B(n37491), .Z(n37472) );
  ANDN U46558 ( .B(n37492), .A(n37493), .Z(n37466) );
  XNOR U46559 ( .A(n37459), .B(n37494), .Z(n37465) );
  XNOR U46560 ( .A(n37458), .B(n37460), .Z(n37494) );
  NAND U46561 ( .A(n37495), .B(n37496), .Z(n37460) );
  OR U46562 ( .A(n37497), .B(n37498), .Z(n37496) );
  OR U46563 ( .A(n37499), .B(n37500), .Z(n37495) );
  NAND U46564 ( .A(n37501), .B(n37502), .Z(n37458) );
  OR U46565 ( .A(n37503), .B(n37504), .Z(n37502) );
  OR U46566 ( .A(n37505), .B(n37506), .Z(n37501) );
  ANDN U46567 ( .B(n37507), .A(n37508), .Z(n37459) );
  IV U46568 ( .A(n37509), .Z(n37507) );
  ANDN U46569 ( .B(n37510), .A(n37511), .Z(n37451) );
  XOR U46570 ( .A(n37437), .B(n37512), .Z(n37449) );
  XOR U46571 ( .A(n37438), .B(n37439), .Z(n37512) );
  XOR U46572 ( .A(n37444), .B(n37513), .Z(n37439) );
  XOR U46573 ( .A(n37443), .B(n37446), .Z(n37513) );
  IV U46574 ( .A(n37445), .Z(n37446) );
  NAND U46575 ( .A(n37514), .B(n37515), .Z(n37445) );
  OR U46576 ( .A(n37516), .B(n37517), .Z(n37515) );
  OR U46577 ( .A(n37518), .B(n37519), .Z(n37514) );
  NAND U46578 ( .A(n37520), .B(n37521), .Z(n37443) );
  OR U46579 ( .A(n37522), .B(n37523), .Z(n37521) );
  OR U46580 ( .A(n37524), .B(n37525), .Z(n37520) );
  NOR U46581 ( .A(n37526), .B(n37527), .Z(n37444) );
  ANDN U46582 ( .B(n37528), .A(n37529), .Z(n37438) );
  IV U46583 ( .A(n37530), .Z(n37528) );
  XNOR U46584 ( .A(n37431), .B(n37531), .Z(n37437) );
  XNOR U46585 ( .A(n37430), .B(n37432), .Z(n37531) );
  NAND U46586 ( .A(n37532), .B(n37533), .Z(n37432) );
  OR U46587 ( .A(n37534), .B(n37535), .Z(n37533) );
  OR U46588 ( .A(n37536), .B(n37537), .Z(n37532) );
  NAND U46589 ( .A(n37538), .B(n37539), .Z(n37430) );
  OR U46590 ( .A(n37540), .B(n37541), .Z(n37539) );
  OR U46591 ( .A(n37542), .B(n37543), .Z(n37538) );
  ANDN U46592 ( .B(n37544), .A(n37545), .Z(n37431) );
  IV U46593 ( .A(n37546), .Z(n37544) );
  XNOR U46594 ( .A(n37511), .B(n37510), .Z(N62074) );
  XOR U46595 ( .A(n37530), .B(n37529), .Z(n37510) );
  XNOR U46596 ( .A(n37545), .B(n37546), .Z(n37529) );
  XNOR U46597 ( .A(n37540), .B(n37541), .Z(n37546) );
  XNOR U46598 ( .A(n37542), .B(n37543), .Z(n37541) );
  XNOR U46599 ( .A(y[2749]), .B(x[2749]), .Z(n37543) );
  XNOR U46600 ( .A(y[2750]), .B(x[2750]), .Z(n37542) );
  XNOR U46601 ( .A(y[2748]), .B(x[2748]), .Z(n37540) );
  XNOR U46602 ( .A(n37534), .B(n37535), .Z(n37545) );
  XNOR U46603 ( .A(y[2745]), .B(x[2745]), .Z(n37535) );
  XNOR U46604 ( .A(n37536), .B(n37537), .Z(n37534) );
  XNOR U46605 ( .A(y[2746]), .B(x[2746]), .Z(n37537) );
  XNOR U46606 ( .A(y[2747]), .B(x[2747]), .Z(n37536) );
  XNOR U46607 ( .A(n37527), .B(n37526), .Z(n37530) );
  XNOR U46608 ( .A(n37522), .B(n37523), .Z(n37526) );
  XNOR U46609 ( .A(y[2742]), .B(x[2742]), .Z(n37523) );
  XNOR U46610 ( .A(n37524), .B(n37525), .Z(n37522) );
  XNOR U46611 ( .A(y[2743]), .B(x[2743]), .Z(n37525) );
  XNOR U46612 ( .A(y[2744]), .B(x[2744]), .Z(n37524) );
  XNOR U46613 ( .A(n37516), .B(n37517), .Z(n37527) );
  XNOR U46614 ( .A(y[2739]), .B(x[2739]), .Z(n37517) );
  XNOR U46615 ( .A(n37518), .B(n37519), .Z(n37516) );
  XNOR U46616 ( .A(y[2740]), .B(x[2740]), .Z(n37519) );
  XNOR U46617 ( .A(y[2741]), .B(x[2741]), .Z(n37518) );
  XOR U46618 ( .A(n37492), .B(n37493), .Z(n37511) );
  XNOR U46619 ( .A(n37508), .B(n37509), .Z(n37493) );
  XNOR U46620 ( .A(n37503), .B(n37504), .Z(n37509) );
  XNOR U46621 ( .A(n37505), .B(n37506), .Z(n37504) );
  XNOR U46622 ( .A(y[2737]), .B(x[2737]), .Z(n37506) );
  XNOR U46623 ( .A(y[2738]), .B(x[2738]), .Z(n37505) );
  XNOR U46624 ( .A(y[2736]), .B(x[2736]), .Z(n37503) );
  XNOR U46625 ( .A(n37497), .B(n37498), .Z(n37508) );
  XNOR U46626 ( .A(y[2733]), .B(x[2733]), .Z(n37498) );
  XNOR U46627 ( .A(n37499), .B(n37500), .Z(n37497) );
  XNOR U46628 ( .A(y[2734]), .B(x[2734]), .Z(n37500) );
  XNOR U46629 ( .A(y[2735]), .B(x[2735]), .Z(n37499) );
  XOR U46630 ( .A(n37491), .B(n37490), .Z(n37492) );
  XNOR U46631 ( .A(n37486), .B(n37487), .Z(n37490) );
  XNOR U46632 ( .A(y[2730]), .B(x[2730]), .Z(n37487) );
  XNOR U46633 ( .A(n37488), .B(n37489), .Z(n37486) );
  XNOR U46634 ( .A(y[2731]), .B(x[2731]), .Z(n37489) );
  XNOR U46635 ( .A(y[2732]), .B(x[2732]), .Z(n37488) );
  XNOR U46636 ( .A(n37480), .B(n37481), .Z(n37491) );
  XNOR U46637 ( .A(y[2727]), .B(x[2727]), .Z(n37481) );
  XNOR U46638 ( .A(n37482), .B(n37483), .Z(n37480) );
  XNOR U46639 ( .A(y[2728]), .B(x[2728]), .Z(n37483) );
  XNOR U46640 ( .A(y[2729]), .B(x[2729]), .Z(n37482) );
  NAND U46641 ( .A(n37547), .B(n37548), .Z(N62065) );
  NANDN U46642 ( .A(n37549), .B(n37550), .Z(n37548) );
  OR U46643 ( .A(n37551), .B(n37552), .Z(n37550) );
  NAND U46644 ( .A(n37551), .B(n37552), .Z(n37547) );
  XOR U46645 ( .A(n37551), .B(n37553), .Z(N62064) );
  XNOR U46646 ( .A(n37549), .B(n37552), .Z(n37553) );
  AND U46647 ( .A(n37554), .B(n37555), .Z(n37552) );
  NANDN U46648 ( .A(n37556), .B(n37557), .Z(n37555) );
  NANDN U46649 ( .A(n37558), .B(n37559), .Z(n37557) );
  NANDN U46650 ( .A(n37559), .B(n37558), .Z(n37554) );
  NAND U46651 ( .A(n37560), .B(n37561), .Z(n37549) );
  NANDN U46652 ( .A(n37562), .B(n37563), .Z(n37561) );
  OR U46653 ( .A(n37564), .B(n37565), .Z(n37563) );
  NAND U46654 ( .A(n37565), .B(n37564), .Z(n37560) );
  AND U46655 ( .A(n37566), .B(n37567), .Z(n37551) );
  NANDN U46656 ( .A(n37568), .B(n37569), .Z(n37567) );
  NANDN U46657 ( .A(n37570), .B(n37571), .Z(n37569) );
  NANDN U46658 ( .A(n37571), .B(n37570), .Z(n37566) );
  XOR U46659 ( .A(n37565), .B(n37572), .Z(N62063) );
  XOR U46660 ( .A(n37562), .B(n37564), .Z(n37572) );
  XNOR U46661 ( .A(n37558), .B(n37573), .Z(n37564) );
  XNOR U46662 ( .A(n37556), .B(n37559), .Z(n37573) );
  NAND U46663 ( .A(n37574), .B(n37575), .Z(n37559) );
  NAND U46664 ( .A(n37576), .B(n37577), .Z(n37575) );
  OR U46665 ( .A(n37578), .B(n37579), .Z(n37576) );
  NANDN U46666 ( .A(n37580), .B(n37578), .Z(n37574) );
  IV U46667 ( .A(n37579), .Z(n37580) );
  NAND U46668 ( .A(n37581), .B(n37582), .Z(n37556) );
  NAND U46669 ( .A(n37583), .B(n37584), .Z(n37582) );
  NANDN U46670 ( .A(n37585), .B(n37586), .Z(n37583) );
  NANDN U46671 ( .A(n37586), .B(n37585), .Z(n37581) );
  AND U46672 ( .A(n37587), .B(n37588), .Z(n37558) );
  NAND U46673 ( .A(n37589), .B(n37590), .Z(n37588) );
  OR U46674 ( .A(n37591), .B(n37592), .Z(n37589) );
  NANDN U46675 ( .A(n37593), .B(n37591), .Z(n37587) );
  NAND U46676 ( .A(n37594), .B(n37595), .Z(n37562) );
  NANDN U46677 ( .A(n37596), .B(n37597), .Z(n37595) );
  OR U46678 ( .A(n37598), .B(n37599), .Z(n37597) );
  NANDN U46679 ( .A(n37600), .B(n37598), .Z(n37594) );
  IV U46680 ( .A(n37599), .Z(n37600) );
  XNOR U46681 ( .A(n37570), .B(n37601), .Z(n37565) );
  XNOR U46682 ( .A(n37568), .B(n37571), .Z(n37601) );
  NAND U46683 ( .A(n37602), .B(n37603), .Z(n37571) );
  NAND U46684 ( .A(n37604), .B(n37605), .Z(n37603) );
  OR U46685 ( .A(n37606), .B(n37607), .Z(n37604) );
  NANDN U46686 ( .A(n37608), .B(n37606), .Z(n37602) );
  IV U46687 ( .A(n37607), .Z(n37608) );
  NAND U46688 ( .A(n37609), .B(n37610), .Z(n37568) );
  NAND U46689 ( .A(n37611), .B(n37612), .Z(n37610) );
  NANDN U46690 ( .A(n37613), .B(n37614), .Z(n37611) );
  NANDN U46691 ( .A(n37614), .B(n37613), .Z(n37609) );
  AND U46692 ( .A(n37615), .B(n37616), .Z(n37570) );
  NAND U46693 ( .A(n37617), .B(n37618), .Z(n37616) );
  OR U46694 ( .A(n37619), .B(n37620), .Z(n37617) );
  NANDN U46695 ( .A(n37621), .B(n37619), .Z(n37615) );
  XNOR U46696 ( .A(n37596), .B(n37622), .Z(N62062) );
  XOR U46697 ( .A(n37598), .B(n37599), .Z(n37622) );
  XNOR U46698 ( .A(n37612), .B(n37623), .Z(n37599) );
  XOR U46699 ( .A(n37613), .B(n37614), .Z(n37623) );
  XOR U46700 ( .A(n37619), .B(n37624), .Z(n37614) );
  XOR U46701 ( .A(n37618), .B(n37621), .Z(n37624) );
  IV U46702 ( .A(n37620), .Z(n37621) );
  NAND U46703 ( .A(n37625), .B(n37626), .Z(n37620) );
  OR U46704 ( .A(n37627), .B(n37628), .Z(n37626) );
  OR U46705 ( .A(n37629), .B(n37630), .Z(n37625) );
  NAND U46706 ( .A(n37631), .B(n37632), .Z(n37618) );
  OR U46707 ( .A(n37633), .B(n37634), .Z(n37632) );
  OR U46708 ( .A(n37635), .B(n37636), .Z(n37631) );
  NOR U46709 ( .A(n37637), .B(n37638), .Z(n37619) );
  ANDN U46710 ( .B(n37639), .A(n37640), .Z(n37613) );
  XNOR U46711 ( .A(n37606), .B(n37641), .Z(n37612) );
  XNOR U46712 ( .A(n37605), .B(n37607), .Z(n37641) );
  NAND U46713 ( .A(n37642), .B(n37643), .Z(n37607) );
  OR U46714 ( .A(n37644), .B(n37645), .Z(n37643) );
  OR U46715 ( .A(n37646), .B(n37647), .Z(n37642) );
  NAND U46716 ( .A(n37648), .B(n37649), .Z(n37605) );
  OR U46717 ( .A(n37650), .B(n37651), .Z(n37649) );
  OR U46718 ( .A(n37652), .B(n37653), .Z(n37648) );
  ANDN U46719 ( .B(n37654), .A(n37655), .Z(n37606) );
  IV U46720 ( .A(n37656), .Z(n37654) );
  ANDN U46721 ( .B(n37657), .A(n37658), .Z(n37598) );
  XOR U46722 ( .A(n37584), .B(n37659), .Z(n37596) );
  XOR U46723 ( .A(n37585), .B(n37586), .Z(n37659) );
  XOR U46724 ( .A(n37591), .B(n37660), .Z(n37586) );
  XOR U46725 ( .A(n37590), .B(n37593), .Z(n37660) );
  IV U46726 ( .A(n37592), .Z(n37593) );
  NAND U46727 ( .A(n37661), .B(n37662), .Z(n37592) );
  OR U46728 ( .A(n37663), .B(n37664), .Z(n37662) );
  OR U46729 ( .A(n37665), .B(n37666), .Z(n37661) );
  NAND U46730 ( .A(n37667), .B(n37668), .Z(n37590) );
  OR U46731 ( .A(n37669), .B(n37670), .Z(n37668) );
  OR U46732 ( .A(n37671), .B(n37672), .Z(n37667) );
  NOR U46733 ( .A(n37673), .B(n37674), .Z(n37591) );
  ANDN U46734 ( .B(n37675), .A(n37676), .Z(n37585) );
  IV U46735 ( .A(n37677), .Z(n37675) );
  XNOR U46736 ( .A(n37578), .B(n37678), .Z(n37584) );
  XNOR U46737 ( .A(n37577), .B(n37579), .Z(n37678) );
  NAND U46738 ( .A(n37679), .B(n37680), .Z(n37579) );
  OR U46739 ( .A(n37681), .B(n37682), .Z(n37680) );
  OR U46740 ( .A(n37683), .B(n37684), .Z(n37679) );
  NAND U46741 ( .A(n37685), .B(n37686), .Z(n37577) );
  OR U46742 ( .A(n37687), .B(n37688), .Z(n37686) );
  OR U46743 ( .A(n37689), .B(n37690), .Z(n37685) );
  ANDN U46744 ( .B(n37691), .A(n37692), .Z(n37578) );
  IV U46745 ( .A(n37693), .Z(n37691) );
  XNOR U46746 ( .A(n37658), .B(n37657), .Z(N62061) );
  XOR U46747 ( .A(n37677), .B(n37676), .Z(n37657) );
  XNOR U46748 ( .A(n37692), .B(n37693), .Z(n37676) );
  XNOR U46749 ( .A(n37687), .B(n37688), .Z(n37693) );
  XNOR U46750 ( .A(n37689), .B(n37690), .Z(n37688) );
  XNOR U46751 ( .A(y[2725]), .B(x[2725]), .Z(n37690) );
  XNOR U46752 ( .A(y[2726]), .B(x[2726]), .Z(n37689) );
  XNOR U46753 ( .A(y[2724]), .B(x[2724]), .Z(n37687) );
  XNOR U46754 ( .A(n37681), .B(n37682), .Z(n37692) );
  XNOR U46755 ( .A(y[2721]), .B(x[2721]), .Z(n37682) );
  XNOR U46756 ( .A(n37683), .B(n37684), .Z(n37681) );
  XNOR U46757 ( .A(y[2722]), .B(x[2722]), .Z(n37684) );
  XNOR U46758 ( .A(y[2723]), .B(x[2723]), .Z(n37683) );
  XNOR U46759 ( .A(n37674), .B(n37673), .Z(n37677) );
  XNOR U46760 ( .A(n37669), .B(n37670), .Z(n37673) );
  XNOR U46761 ( .A(y[2718]), .B(x[2718]), .Z(n37670) );
  XNOR U46762 ( .A(n37671), .B(n37672), .Z(n37669) );
  XNOR U46763 ( .A(y[2719]), .B(x[2719]), .Z(n37672) );
  XNOR U46764 ( .A(y[2720]), .B(x[2720]), .Z(n37671) );
  XNOR U46765 ( .A(n37663), .B(n37664), .Z(n37674) );
  XNOR U46766 ( .A(y[2715]), .B(x[2715]), .Z(n37664) );
  XNOR U46767 ( .A(n37665), .B(n37666), .Z(n37663) );
  XNOR U46768 ( .A(y[2716]), .B(x[2716]), .Z(n37666) );
  XNOR U46769 ( .A(y[2717]), .B(x[2717]), .Z(n37665) );
  XOR U46770 ( .A(n37639), .B(n37640), .Z(n37658) );
  XNOR U46771 ( .A(n37655), .B(n37656), .Z(n37640) );
  XNOR U46772 ( .A(n37650), .B(n37651), .Z(n37656) );
  XNOR U46773 ( .A(n37652), .B(n37653), .Z(n37651) );
  XNOR U46774 ( .A(y[2713]), .B(x[2713]), .Z(n37653) );
  XNOR U46775 ( .A(y[2714]), .B(x[2714]), .Z(n37652) );
  XNOR U46776 ( .A(y[2712]), .B(x[2712]), .Z(n37650) );
  XNOR U46777 ( .A(n37644), .B(n37645), .Z(n37655) );
  XNOR U46778 ( .A(y[2709]), .B(x[2709]), .Z(n37645) );
  XNOR U46779 ( .A(n37646), .B(n37647), .Z(n37644) );
  XNOR U46780 ( .A(y[2710]), .B(x[2710]), .Z(n37647) );
  XNOR U46781 ( .A(y[2711]), .B(x[2711]), .Z(n37646) );
  XOR U46782 ( .A(n37638), .B(n37637), .Z(n37639) );
  XNOR U46783 ( .A(n37633), .B(n37634), .Z(n37637) );
  XNOR U46784 ( .A(y[2706]), .B(x[2706]), .Z(n37634) );
  XNOR U46785 ( .A(n37635), .B(n37636), .Z(n37633) );
  XNOR U46786 ( .A(y[2707]), .B(x[2707]), .Z(n37636) );
  XNOR U46787 ( .A(y[2708]), .B(x[2708]), .Z(n37635) );
  XNOR U46788 ( .A(n37627), .B(n37628), .Z(n37638) );
  XNOR U46789 ( .A(y[2703]), .B(x[2703]), .Z(n37628) );
  XNOR U46790 ( .A(n37629), .B(n37630), .Z(n37627) );
  XNOR U46791 ( .A(y[2704]), .B(x[2704]), .Z(n37630) );
  XNOR U46792 ( .A(y[2705]), .B(x[2705]), .Z(n37629) );
  NAND U46793 ( .A(n37694), .B(n37695), .Z(N62052) );
  NANDN U46794 ( .A(n37696), .B(n37697), .Z(n37695) );
  OR U46795 ( .A(n37698), .B(n37699), .Z(n37697) );
  NAND U46796 ( .A(n37698), .B(n37699), .Z(n37694) );
  XOR U46797 ( .A(n37698), .B(n37700), .Z(N62051) );
  XNOR U46798 ( .A(n37696), .B(n37699), .Z(n37700) );
  AND U46799 ( .A(n37701), .B(n37702), .Z(n37699) );
  NANDN U46800 ( .A(n37703), .B(n37704), .Z(n37702) );
  NANDN U46801 ( .A(n37705), .B(n37706), .Z(n37704) );
  NANDN U46802 ( .A(n37706), .B(n37705), .Z(n37701) );
  NAND U46803 ( .A(n37707), .B(n37708), .Z(n37696) );
  NANDN U46804 ( .A(n37709), .B(n37710), .Z(n37708) );
  OR U46805 ( .A(n37711), .B(n37712), .Z(n37710) );
  NAND U46806 ( .A(n37712), .B(n37711), .Z(n37707) );
  AND U46807 ( .A(n37713), .B(n37714), .Z(n37698) );
  NANDN U46808 ( .A(n37715), .B(n37716), .Z(n37714) );
  NANDN U46809 ( .A(n37717), .B(n37718), .Z(n37716) );
  NANDN U46810 ( .A(n37718), .B(n37717), .Z(n37713) );
  XOR U46811 ( .A(n37712), .B(n37719), .Z(N62050) );
  XOR U46812 ( .A(n37709), .B(n37711), .Z(n37719) );
  XNOR U46813 ( .A(n37705), .B(n37720), .Z(n37711) );
  XNOR U46814 ( .A(n37703), .B(n37706), .Z(n37720) );
  NAND U46815 ( .A(n37721), .B(n37722), .Z(n37706) );
  NAND U46816 ( .A(n37723), .B(n37724), .Z(n37722) );
  OR U46817 ( .A(n37725), .B(n37726), .Z(n37723) );
  NANDN U46818 ( .A(n37727), .B(n37725), .Z(n37721) );
  IV U46819 ( .A(n37726), .Z(n37727) );
  NAND U46820 ( .A(n37728), .B(n37729), .Z(n37703) );
  NAND U46821 ( .A(n37730), .B(n37731), .Z(n37729) );
  NANDN U46822 ( .A(n37732), .B(n37733), .Z(n37730) );
  NANDN U46823 ( .A(n37733), .B(n37732), .Z(n37728) );
  AND U46824 ( .A(n37734), .B(n37735), .Z(n37705) );
  NAND U46825 ( .A(n37736), .B(n37737), .Z(n37735) );
  OR U46826 ( .A(n37738), .B(n37739), .Z(n37736) );
  NANDN U46827 ( .A(n37740), .B(n37738), .Z(n37734) );
  NAND U46828 ( .A(n37741), .B(n37742), .Z(n37709) );
  NANDN U46829 ( .A(n37743), .B(n37744), .Z(n37742) );
  OR U46830 ( .A(n37745), .B(n37746), .Z(n37744) );
  NANDN U46831 ( .A(n37747), .B(n37745), .Z(n37741) );
  IV U46832 ( .A(n37746), .Z(n37747) );
  XNOR U46833 ( .A(n37717), .B(n37748), .Z(n37712) );
  XNOR U46834 ( .A(n37715), .B(n37718), .Z(n37748) );
  NAND U46835 ( .A(n37749), .B(n37750), .Z(n37718) );
  NAND U46836 ( .A(n37751), .B(n37752), .Z(n37750) );
  OR U46837 ( .A(n37753), .B(n37754), .Z(n37751) );
  NANDN U46838 ( .A(n37755), .B(n37753), .Z(n37749) );
  IV U46839 ( .A(n37754), .Z(n37755) );
  NAND U46840 ( .A(n37756), .B(n37757), .Z(n37715) );
  NAND U46841 ( .A(n37758), .B(n37759), .Z(n37757) );
  NANDN U46842 ( .A(n37760), .B(n37761), .Z(n37758) );
  NANDN U46843 ( .A(n37761), .B(n37760), .Z(n37756) );
  AND U46844 ( .A(n37762), .B(n37763), .Z(n37717) );
  NAND U46845 ( .A(n37764), .B(n37765), .Z(n37763) );
  OR U46846 ( .A(n37766), .B(n37767), .Z(n37764) );
  NANDN U46847 ( .A(n37768), .B(n37766), .Z(n37762) );
  XNOR U46848 ( .A(n37743), .B(n37769), .Z(N62049) );
  XOR U46849 ( .A(n37745), .B(n37746), .Z(n37769) );
  XNOR U46850 ( .A(n37759), .B(n37770), .Z(n37746) );
  XOR U46851 ( .A(n37760), .B(n37761), .Z(n37770) );
  XOR U46852 ( .A(n37766), .B(n37771), .Z(n37761) );
  XOR U46853 ( .A(n37765), .B(n37768), .Z(n37771) );
  IV U46854 ( .A(n37767), .Z(n37768) );
  NAND U46855 ( .A(n37772), .B(n37773), .Z(n37767) );
  OR U46856 ( .A(n37774), .B(n37775), .Z(n37773) );
  OR U46857 ( .A(n37776), .B(n37777), .Z(n37772) );
  NAND U46858 ( .A(n37778), .B(n37779), .Z(n37765) );
  OR U46859 ( .A(n37780), .B(n37781), .Z(n37779) );
  OR U46860 ( .A(n37782), .B(n37783), .Z(n37778) );
  NOR U46861 ( .A(n37784), .B(n37785), .Z(n37766) );
  ANDN U46862 ( .B(n37786), .A(n37787), .Z(n37760) );
  XNOR U46863 ( .A(n37753), .B(n37788), .Z(n37759) );
  XNOR U46864 ( .A(n37752), .B(n37754), .Z(n37788) );
  NAND U46865 ( .A(n37789), .B(n37790), .Z(n37754) );
  OR U46866 ( .A(n37791), .B(n37792), .Z(n37790) );
  OR U46867 ( .A(n37793), .B(n37794), .Z(n37789) );
  NAND U46868 ( .A(n37795), .B(n37796), .Z(n37752) );
  OR U46869 ( .A(n37797), .B(n37798), .Z(n37796) );
  OR U46870 ( .A(n37799), .B(n37800), .Z(n37795) );
  ANDN U46871 ( .B(n37801), .A(n37802), .Z(n37753) );
  IV U46872 ( .A(n37803), .Z(n37801) );
  ANDN U46873 ( .B(n37804), .A(n37805), .Z(n37745) );
  XOR U46874 ( .A(n37731), .B(n37806), .Z(n37743) );
  XOR U46875 ( .A(n37732), .B(n37733), .Z(n37806) );
  XOR U46876 ( .A(n37738), .B(n37807), .Z(n37733) );
  XOR U46877 ( .A(n37737), .B(n37740), .Z(n37807) );
  IV U46878 ( .A(n37739), .Z(n37740) );
  NAND U46879 ( .A(n37808), .B(n37809), .Z(n37739) );
  OR U46880 ( .A(n37810), .B(n37811), .Z(n37809) );
  OR U46881 ( .A(n37812), .B(n37813), .Z(n37808) );
  NAND U46882 ( .A(n37814), .B(n37815), .Z(n37737) );
  OR U46883 ( .A(n37816), .B(n37817), .Z(n37815) );
  OR U46884 ( .A(n37818), .B(n37819), .Z(n37814) );
  NOR U46885 ( .A(n37820), .B(n37821), .Z(n37738) );
  ANDN U46886 ( .B(n37822), .A(n37823), .Z(n37732) );
  IV U46887 ( .A(n37824), .Z(n37822) );
  XNOR U46888 ( .A(n37725), .B(n37825), .Z(n37731) );
  XNOR U46889 ( .A(n37724), .B(n37726), .Z(n37825) );
  NAND U46890 ( .A(n37826), .B(n37827), .Z(n37726) );
  OR U46891 ( .A(n37828), .B(n37829), .Z(n37827) );
  OR U46892 ( .A(n37830), .B(n37831), .Z(n37826) );
  NAND U46893 ( .A(n37832), .B(n37833), .Z(n37724) );
  OR U46894 ( .A(n37834), .B(n37835), .Z(n37833) );
  OR U46895 ( .A(n37836), .B(n37837), .Z(n37832) );
  ANDN U46896 ( .B(n37838), .A(n37839), .Z(n37725) );
  IV U46897 ( .A(n37840), .Z(n37838) );
  XNOR U46898 ( .A(n37805), .B(n37804), .Z(N62048) );
  XOR U46899 ( .A(n37824), .B(n37823), .Z(n37804) );
  XNOR U46900 ( .A(n37839), .B(n37840), .Z(n37823) );
  XNOR U46901 ( .A(n37834), .B(n37835), .Z(n37840) );
  XNOR U46902 ( .A(n37836), .B(n37837), .Z(n37835) );
  XNOR U46903 ( .A(y[2701]), .B(x[2701]), .Z(n37837) );
  XNOR U46904 ( .A(y[2702]), .B(x[2702]), .Z(n37836) );
  XNOR U46905 ( .A(y[2700]), .B(x[2700]), .Z(n37834) );
  XNOR U46906 ( .A(n37828), .B(n37829), .Z(n37839) );
  XNOR U46907 ( .A(y[2697]), .B(x[2697]), .Z(n37829) );
  XNOR U46908 ( .A(n37830), .B(n37831), .Z(n37828) );
  XNOR U46909 ( .A(y[2698]), .B(x[2698]), .Z(n37831) );
  XNOR U46910 ( .A(y[2699]), .B(x[2699]), .Z(n37830) );
  XNOR U46911 ( .A(n37821), .B(n37820), .Z(n37824) );
  XNOR U46912 ( .A(n37816), .B(n37817), .Z(n37820) );
  XNOR U46913 ( .A(y[2694]), .B(x[2694]), .Z(n37817) );
  XNOR U46914 ( .A(n37818), .B(n37819), .Z(n37816) );
  XNOR U46915 ( .A(y[2695]), .B(x[2695]), .Z(n37819) );
  XNOR U46916 ( .A(y[2696]), .B(x[2696]), .Z(n37818) );
  XNOR U46917 ( .A(n37810), .B(n37811), .Z(n37821) );
  XNOR U46918 ( .A(y[2691]), .B(x[2691]), .Z(n37811) );
  XNOR U46919 ( .A(n37812), .B(n37813), .Z(n37810) );
  XNOR U46920 ( .A(y[2692]), .B(x[2692]), .Z(n37813) );
  XNOR U46921 ( .A(y[2693]), .B(x[2693]), .Z(n37812) );
  XOR U46922 ( .A(n37786), .B(n37787), .Z(n37805) );
  XNOR U46923 ( .A(n37802), .B(n37803), .Z(n37787) );
  XNOR U46924 ( .A(n37797), .B(n37798), .Z(n37803) );
  XNOR U46925 ( .A(n37799), .B(n37800), .Z(n37798) );
  XNOR U46926 ( .A(y[2689]), .B(x[2689]), .Z(n37800) );
  XNOR U46927 ( .A(y[2690]), .B(x[2690]), .Z(n37799) );
  XNOR U46928 ( .A(y[2688]), .B(x[2688]), .Z(n37797) );
  XNOR U46929 ( .A(n37791), .B(n37792), .Z(n37802) );
  XNOR U46930 ( .A(y[2685]), .B(x[2685]), .Z(n37792) );
  XNOR U46931 ( .A(n37793), .B(n37794), .Z(n37791) );
  XNOR U46932 ( .A(y[2686]), .B(x[2686]), .Z(n37794) );
  XNOR U46933 ( .A(y[2687]), .B(x[2687]), .Z(n37793) );
  XOR U46934 ( .A(n37785), .B(n37784), .Z(n37786) );
  XNOR U46935 ( .A(n37780), .B(n37781), .Z(n37784) );
  XNOR U46936 ( .A(y[2682]), .B(x[2682]), .Z(n37781) );
  XNOR U46937 ( .A(n37782), .B(n37783), .Z(n37780) );
  XNOR U46938 ( .A(y[2683]), .B(x[2683]), .Z(n37783) );
  XNOR U46939 ( .A(y[2684]), .B(x[2684]), .Z(n37782) );
  XNOR U46940 ( .A(n37774), .B(n37775), .Z(n37785) );
  XNOR U46941 ( .A(y[2679]), .B(x[2679]), .Z(n37775) );
  XNOR U46942 ( .A(n37776), .B(n37777), .Z(n37774) );
  XNOR U46943 ( .A(y[2680]), .B(x[2680]), .Z(n37777) );
  XNOR U46944 ( .A(y[2681]), .B(x[2681]), .Z(n37776) );
  NAND U46945 ( .A(n37841), .B(n37842), .Z(N62039) );
  NANDN U46946 ( .A(n37843), .B(n37844), .Z(n37842) );
  OR U46947 ( .A(n37845), .B(n37846), .Z(n37844) );
  NAND U46948 ( .A(n37845), .B(n37846), .Z(n37841) );
  XOR U46949 ( .A(n37845), .B(n37847), .Z(N62038) );
  XNOR U46950 ( .A(n37843), .B(n37846), .Z(n37847) );
  AND U46951 ( .A(n37848), .B(n37849), .Z(n37846) );
  NANDN U46952 ( .A(n37850), .B(n37851), .Z(n37849) );
  NANDN U46953 ( .A(n37852), .B(n37853), .Z(n37851) );
  NANDN U46954 ( .A(n37853), .B(n37852), .Z(n37848) );
  NAND U46955 ( .A(n37854), .B(n37855), .Z(n37843) );
  NANDN U46956 ( .A(n37856), .B(n37857), .Z(n37855) );
  OR U46957 ( .A(n37858), .B(n37859), .Z(n37857) );
  NAND U46958 ( .A(n37859), .B(n37858), .Z(n37854) );
  AND U46959 ( .A(n37860), .B(n37861), .Z(n37845) );
  NANDN U46960 ( .A(n37862), .B(n37863), .Z(n37861) );
  NANDN U46961 ( .A(n37864), .B(n37865), .Z(n37863) );
  NANDN U46962 ( .A(n37865), .B(n37864), .Z(n37860) );
  XOR U46963 ( .A(n37859), .B(n37866), .Z(N62037) );
  XOR U46964 ( .A(n37856), .B(n37858), .Z(n37866) );
  XNOR U46965 ( .A(n37852), .B(n37867), .Z(n37858) );
  XNOR U46966 ( .A(n37850), .B(n37853), .Z(n37867) );
  NAND U46967 ( .A(n37868), .B(n37869), .Z(n37853) );
  NAND U46968 ( .A(n37870), .B(n37871), .Z(n37869) );
  OR U46969 ( .A(n37872), .B(n37873), .Z(n37870) );
  NANDN U46970 ( .A(n37874), .B(n37872), .Z(n37868) );
  IV U46971 ( .A(n37873), .Z(n37874) );
  NAND U46972 ( .A(n37875), .B(n37876), .Z(n37850) );
  NAND U46973 ( .A(n37877), .B(n37878), .Z(n37876) );
  NANDN U46974 ( .A(n37879), .B(n37880), .Z(n37877) );
  NANDN U46975 ( .A(n37880), .B(n37879), .Z(n37875) );
  AND U46976 ( .A(n37881), .B(n37882), .Z(n37852) );
  NAND U46977 ( .A(n37883), .B(n37884), .Z(n37882) );
  OR U46978 ( .A(n37885), .B(n37886), .Z(n37883) );
  NANDN U46979 ( .A(n37887), .B(n37885), .Z(n37881) );
  NAND U46980 ( .A(n37888), .B(n37889), .Z(n37856) );
  NANDN U46981 ( .A(n37890), .B(n37891), .Z(n37889) );
  OR U46982 ( .A(n37892), .B(n37893), .Z(n37891) );
  NANDN U46983 ( .A(n37894), .B(n37892), .Z(n37888) );
  IV U46984 ( .A(n37893), .Z(n37894) );
  XNOR U46985 ( .A(n37864), .B(n37895), .Z(n37859) );
  XNOR U46986 ( .A(n37862), .B(n37865), .Z(n37895) );
  NAND U46987 ( .A(n37896), .B(n37897), .Z(n37865) );
  NAND U46988 ( .A(n37898), .B(n37899), .Z(n37897) );
  OR U46989 ( .A(n37900), .B(n37901), .Z(n37898) );
  NANDN U46990 ( .A(n37902), .B(n37900), .Z(n37896) );
  IV U46991 ( .A(n37901), .Z(n37902) );
  NAND U46992 ( .A(n37903), .B(n37904), .Z(n37862) );
  NAND U46993 ( .A(n37905), .B(n37906), .Z(n37904) );
  NANDN U46994 ( .A(n37907), .B(n37908), .Z(n37905) );
  NANDN U46995 ( .A(n37908), .B(n37907), .Z(n37903) );
  AND U46996 ( .A(n37909), .B(n37910), .Z(n37864) );
  NAND U46997 ( .A(n37911), .B(n37912), .Z(n37910) );
  OR U46998 ( .A(n37913), .B(n37914), .Z(n37911) );
  NANDN U46999 ( .A(n37915), .B(n37913), .Z(n37909) );
  XNOR U47000 ( .A(n37890), .B(n37916), .Z(N62036) );
  XOR U47001 ( .A(n37892), .B(n37893), .Z(n37916) );
  XNOR U47002 ( .A(n37906), .B(n37917), .Z(n37893) );
  XOR U47003 ( .A(n37907), .B(n37908), .Z(n37917) );
  XOR U47004 ( .A(n37913), .B(n37918), .Z(n37908) );
  XOR U47005 ( .A(n37912), .B(n37915), .Z(n37918) );
  IV U47006 ( .A(n37914), .Z(n37915) );
  NAND U47007 ( .A(n37919), .B(n37920), .Z(n37914) );
  OR U47008 ( .A(n37921), .B(n37922), .Z(n37920) );
  OR U47009 ( .A(n37923), .B(n37924), .Z(n37919) );
  NAND U47010 ( .A(n37925), .B(n37926), .Z(n37912) );
  OR U47011 ( .A(n37927), .B(n37928), .Z(n37926) );
  OR U47012 ( .A(n37929), .B(n37930), .Z(n37925) );
  NOR U47013 ( .A(n37931), .B(n37932), .Z(n37913) );
  ANDN U47014 ( .B(n37933), .A(n37934), .Z(n37907) );
  XNOR U47015 ( .A(n37900), .B(n37935), .Z(n37906) );
  XNOR U47016 ( .A(n37899), .B(n37901), .Z(n37935) );
  NAND U47017 ( .A(n37936), .B(n37937), .Z(n37901) );
  OR U47018 ( .A(n37938), .B(n37939), .Z(n37937) );
  OR U47019 ( .A(n37940), .B(n37941), .Z(n37936) );
  NAND U47020 ( .A(n37942), .B(n37943), .Z(n37899) );
  OR U47021 ( .A(n37944), .B(n37945), .Z(n37943) );
  OR U47022 ( .A(n37946), .B(n37947), .Z(n37942) );
  ANDN U47023 ( .B(n37948), .A(n37949), .Z(n37900) );
  IV U47024 ( .A(n37950), .Z(n37948) );
  ANDN U47025 ( .B(n37951), .A(n37952), .Z(n37892) );
  XOR U47026 ( .A(n37878), .B(n37953), .Z(n37890) );
  XOR U47027 ( .A(n37879), .B(n37880), .Z(n37953) );
  XOR U47028 ( .A(n37885), .B(n37954), .Z(n37880) );
  XOR U47029 ( .A(n37884), .B(n37887), .Z(n37954) );
  IV U47030 ( .A(n37886), .Z(n37887) );
  NAND U47031 ( .A(n37955), .B(n37956), .Z(n37886) );
  OR U47032 ( .A(n37957), .B(n37958), .Z(n37956) );
  OR U47033 ( .A(n37959), .B(n37960), .Z(n37955) );
  NAND U47034 ( .A(n37961), .B(n37962), .Z(n37884) );
  OR U47035 ( .A(n37963), .B(n37964), .Z(n37962) );
  OR U47036 ( .A(n37965), .B(n37966), .Z(n37961) );
  NOR U47037 ( .A(n37967), .B(n37968), .Z(n37885) );
  ANDN U47038 ( .B(n37969), .A(n37970), .Z(n37879) );
  IV U47039 ( .A(n37971), .Z(n37969) );
  XNOR U47040 ( .A(n37872), .B(n37972), .Z(n37878) );
  XNOR U47041 ( .A(n37871), .B(n37873), .Z(n37972) );
  NAND U47042 ( .A(n37973), .B(n37974), .Z(n37873) );
  OR U47043 ( .A(n37975), .B(n37976), .Z(n37974) );
  OR U47044 ( .A(n37977), .B(n37978), .Z(n37973) );
  NAND U47045 ( .A(n37979), .B(n37980), .Z(n37871) );
  OR U47046 ( .A(n37981), .B(n37982), .Z(n37980) );
  OR U47047 ( .A(n37983), .B(n37984), .Z(n37979) );
  ANDN U47048 ( .B(n37985), .A(n37986), .Z(n37872) );
  IV U47049 ( .A(n37987), .Z(n37985) );
  XNOR U47050 ( .A(n37952), .B(n37951), .Z(N62035) );
  XOR U47051 ( .A(n37971), .B(n37970), .Z(n37951) );
  XNOR U47052 ( .A(n37986), .B(n37987), .Z(n37970) );
  XNOR U47053 ( .A(n37981), .B(n37982), .Z(n37987) );
  XNOR U47054 ( .A(n37983), .B(n37984), .Z(n37982) );
  XNOR U47055 ( .A(y[2677]), .B(x[2677]), .Z(n37984) );
  XNOR U47056 ( .A(y[2678]), .B(x[2678]), .Z(n37983) );
  XNOR U47057 ( .A(y[2676]), .B(x[2676]), .Z(n37981) );
  XNOR U47058 ( .A(n37975), .B(n37976), .Z(n37986) );
  XNOR U47059 ( .A(y[2673]), .B(x[2673]), .Z(n37976) );
  XNOR U47060 ( .A(n37977), .B(n37978), .Z(n37975) );
  XNOR U47061 ( .A(y[2674]), .B(x[2674]), .Z(n37978) );
  XNOR U47062 ( .A(y[2675]), .B(x[2675]), .Z(n37977) );
  XNOR U47063 ( .A(n37968), .B(n37967), .Z(n37971) );
  XNOR U47064 ( .A(n37963), .B(n37964), .Z(n37967) );
  XNOR U47065 ( .A(y[2670]), .B(x[2670]), .Z(n37964) );
  XNOR U47066 ( .A(n37965), .B(n37966), .Z(n37963) );
  XNOR U47067 ( .A(y[2671]), .B(x[2671]), .Z(n37966) );
  XNOR U47068 ( .A(y[2672]), .B(x[2672]), .Z(n37965) );
  XNOR U47069 ( .A(n37957), .B(n37958), .Z(n37968) );
  XNOR U47070 ( .A(y[2667]), .B(x[2667]), .Z(n37958) );
  XNOR U47071 ( .A(n37959), .B(n37960), .Z(n37957) );
  XNOR U47072 ( .A(y[2668]), .B(x[2668]), .Z(n37960) );
  XNOR U47073 ( .A(y[2669]), .B(x[2669]), .Z(n37959) );
  XOR U47074 ( .A(n37933), .B(n37934), .Z(n37952) );
  XNOR U47075 ( .A(n37949), .B(n37950), .Z(n37934) );
  XNOR U47076 ( .A(n37944), .B(n37945), .Z(n37950) );
  XNOR U47077 ( .A(n37946), .B(n37947), .Z(n37945) );
  XNOR U47078 ( .A(y[2665]), .B(x[2665]), .Z(n37947) );
  XNOR U47079 ( .A(y[2666]), .B(x[2666]), .Z(n37946) );
  XNOR U47080 ( .A(y[2664]), .B(x[2664]), .Z(n37944) );
  XNOR U47081 ( .A(n37938), .B(n37939), .Z(n37949) );
  XNOR U47082 ( .A(y[2661]), .B(x[2661]), .Z(n37939) );
  XNOR U47083 ( .A(n37940), .B(n37941), .Z(n37938) );
  XNOR U47084 ( .A(y[2662]), .B(x[2662]), .Z(n37941) );
  XNOR U47085 ( .A(y[2663]), .B(x[2663]), .Z(n37940) );
  XOR U47086 ( .A(n37932), .B(n37931), .Z(n37933) );
  XNOR U47087 ( .A(n37927), .B(n37928), .Z(n37931) );
  XNOR U47088 ( .A(y[2658]), .B(x[2658]), .Z(n37928) );
  XNOR U47089 ( .A(n37929), .B(n37930), .Z(n37927) );
  XNOR U47090 ( .A(y[2659]), .B(x[2659]), .Z(n37930) );
  XNOR U47091 ( .A(y[2660]), .B(x[2660]), .Z(n37929) );
  XNOR U47092 ( .A(n37921), .B(n37922), .Z(n37932) );
  XNOR U47093 ( .A(y[2655]), .B(x[2655]), .Z(n37922) );
  XNOR U47094 ( .A(n37923), .B(n37924), .Z(n37921) );
  XNOR U47095 ( .A(y[2656]), .B(x[2656]), .Z(n37924) );
  XNOR U47096 ( .A(y[2657]), .B(x[2657]), .Z(n37923) );
  NAND U47097 ( .A(n37988), .B(n37989), .Z(N62026) );
  NANDN U47098 ( .A(n37990), .B(n37991), .Z(n37989) );
  OR U47099 ( .A(n37992), .B(n37993), .Z(n37991) );
  NAND U47100 ( .A(n37992), .B(n37993), .Z(n37988) );
  XOR U47101 ( .A(n37992), .B(n37994), .Z(N62025) );
  XNOR U47102 ( .A(n37990), .B(n37993), .Z(n37994) );
  AND U47103 ( .A(n37995), .B(n37996), .Z(n37993) );
  NANDN U47104 ( .A(n37997), .B(n37998), .Z(n37996) );
  NANDN U47105 ( .A(n37999), .B(n38000), .Z(n37998) );
  NANDN U47106 ( .A(n38000), .B(n37999), .Z(n37995) );
  NAND U47107 ( .A(n38001), .B(n38002), .Z(n37990) );
  NANDN U47108 ( .A(n38003), .B(n38004), .Z(n38002) );
  OR U47109 ( .A(n38005), .B(n38006), .Z(n38004) );
  NAND U47110 ( .A(n38006), .B(n38005), .Z(n38001) );
  AND U47111 ( .A(n38007), .B(n38008), .Z(n37992) );
  NANDN U47112 ( .A(n38009), .B(n38010), .Z(n38008) );
  NANDN U47113 ( .A(n38011), .B(n38012), .Z(n38010) );
  NANDN U47114 ( .A(n38012), .B(n38011), .Z(n38007) );
  XOR U47115 ( .A(n38006), .B(n38013), .Z(N62024) );
  XOR U47116 ( .A(n38003), .B(n38005), .Z(n38013) );
  XNOR U47117 ( .A(n37999), .B(n38014), .Z(n38005) );
  XNOR U47118 ( .A(n37997), .B(n38000), .Z(n38014) );
  NAND U47119 ( .A(n38015), .B(n38016), .Z(n38000) );
  NAND U47120 ( .A(n38017), .B(n38018), .Z(n38016) );
  OR U47121 ( .A(n38019), .B(n38020), .Z(n38017) );
  NANDN U47122 ( .A(n38021), .B(n38019), .Z(n38015) );
  IV U47123 ( .A(n38020), .Z(n38021) );
  NAND U47124 ( .A(n38022), .B(n38023), .Z(n37997) );
  NAND U47125 ( .A(n38024), .B(n38025), .Z(n38023) );
  NANDN U47126 ( .A(n38026), .B(n38027), .Z(n38024) );
  NANDN U47127 ( .A(n38027), .B(n38026), .Z(n38022) );
  AND U47128 ( .A(n38028), .B(n38029), .Z(n37999) );
  NAND U47129 ( .A(n38030), .B(n38031), .Z(n38029) );
  OR U47130 ( .A(n38032), .B(n38033), .Z(n38030) );
  NANDN U47131 ( .A(n38034), .B(n38032), .Z(n38028) );
  NAND U47132 ( .A(n38035), .B(n38036), .Z(n38003) );
  NANDN U47133 ( .A(n38037), .B(n38038), .Z(n38036) );
  OR U47134 ( .A(n38039), .B(n38040), .Z(n38038) );
  NANDN U47135 ( .A(n38041), .B(n38039), .Z(n38035) );
  IV U47136 ( .A(n38040), .Z(n38041) );
  XNOR U47137 ( .A(n38011), .B(n38042), .Z(n38006) );
  XNOR U47138 ( .A(n38009), .B(n38012), .Z(n38042) );
  NAND U47139 ( .A(n38043), .B(n38044), .Z(n38012) );
  NAND U47140 ( .A(n38045), .B(n38046), .Z(n38044) );
  OR U47141 ( .A(n38047), .B(n38048), .Z(n38045) );
  NANDN U47142 ( .A(n38049), .B(n38047), .Z(n38043) );
  IV U47143 ( .A(n38048), .Z(n38049) );
  NAND U47144 ( .A(n38050), .B(n38051), .Z(n38009) );
  NAND U47145 ( .A(n38052), .B(n38053), .Z(n38051) );
  NANDN U47146 ( .A(n38054), .B(n38055), .Z(n38052) );
  NANDN U47147 ( .A(n38055), .B(n38054), .Z(n38050) );
  AND U47148 ( .A(n38056), .B(n38057), .Z(n38011) );
  NAND U47149 ( .A(n38058), .B(n38059), .Z(n38057) );
  OR U47150 ( .A(n38060), .B(n38061), .Z(n38058) );
  NANDN U47151 ( .A(n38062), .B(n38060), .Z(n38056) );
  XNOR U47152 ( .A(n38037), .B(n38063), .Z(N62023) );
  XOR U47153 ( .A(n38039), .B(n38040), .Z(n38063) );
  XNOR U47154 ( .A(n38053), .B(n38064), .Z(n38040) );
  XOR U47155 ( .A(n38054), .B(n38055), .Z(n38064) );
  XOR U47156 ( .A(n38060), .B(n38065), .Z(n38055) );
  XOR U47157 ( .A(n38059), .B(n38062), .Z(n38065) );
  IV U47158 ( .A(n38061), .Z(n38062) );
  NAND U47159 ( .A(n38066), .B(n38067), .Z(n38061) );
  OR U47160 ( .A(n38068), .B(n38069), .Z(n38067) );
  OR U47161 ( .A(n38070), .B(n38071), .Z(n38066) );
  NAND U47162 ( .A(n38072), .B(n38073), .Z(n38059) );
  OR U47163 ( .A(n38074), .B(n38075), .Z(n38073) );
  OR U47164 ( .A(n38076), .B(n38077), .Z(n38072) );
  NOR U47165 ( .A(n38078), .B(n38079), .Z(n38060) );
  ANDN U47166 ( .B(n38080), .A(n38081), .Z(n38054) );
  XNOR U47167 ( .A(n38047), .B(n38082), .Z(n38053) );
  XNOR U47168 ( .A(n38046), .B(n38048), .Z(n38082) );
  NAND U47169 ( .A(n38083), .B(n38084), .Z(n38048) );
  OR U47170 ( .A(n38085), .B(n38086), .Z(n38084) );
  OR U47171 ( .A(n38087), .B(n38088), .Z(n38083) );
  NAND U47172 ( .A(n38089), .B(n38090), .Z(n38046) );
  OR U47173 ( .A(n38091), .B(n38092), .Z(n38090) );
  OR U47174 ( .A(n38093), .B(n38094), .Z(n38089) );
  ANDN U47175 ( .B(n38095), .A(n38096), .Z(n38047) );
  IV U47176 ( .A(n38097), .Z(n38095) );
  ANDN U47177 ( .B(n38098), .A(n38099), .Z(n38039) );
  XOR U47178 ( .A(n38025), .B(n38100), .Z(n38037) );
  XOR U47179 ( .A(n38026), .B(n38027), .Z(n38100) );
  XOR U47180 ( .A(n38032), .B(n38101), .Z(n38027) );
  XOR U47181 ( .A(n38031), .B(n38034), .Z(n38101) );
  IV U47182 ( .A(n38033), .Z(n38034) );
  NAND U47183 ( .A(n38102), .B(n38103), .Z(n38033) );
  OR U47184 ( .A(n38104), .B(n38105), .Z(n38103) );
  OR U47185 ( .A(n38106), .B(n38107), .Z(n38102) );
  NAND U47186 ( .A(n38108), .B(n38109), .Z(n38031) );
  OR U47187 ( .A(n38110), .B(n38111), .Z(n38109) );
  OR U47188 ( .A(n38112), .B(n38113), .Z(n38108) );
  NOR U47189 ( .A(n38114), .B(n38115), .Z(n38032) );
  ANDN U47190 ( .B(n38116), .A(n38117), .Z(n38026) );
  IV U47191 ( .A(n38118), .Z(n38116) );
  XNOR U47192 ( .A(n38019), .B(n38119), .Z(n38025) );
  XNOR U47193 ( .A(n38018), .B(n38020), .Z(n38119) );
  NAND U47194 ( .A(n38120), .B(n38121), .Z(n38020) );
  OR U47195 ( .A(n38122), .B(n38123), .Z(n38121) );
  OR U47196 ( .A(n38124), .B(n38125), .Z(n38120) );
  NAND U47197 ( .A(n38126), .B(n38127), .Z(n38018) );
  OR U47198 ( .A(n38128), .B(n38129), .Z(n38127) );
  OR U47199 ( .A(n38130), .B(n38131), .Z(n38126) );
  ANDN U47200 ( .B(n38132), .A(n38133), .Z(n38019) );
  IV U47201 ( .A(n38134), .Z(n38132) );
  XNOR U47202 ( .A(n38099), .B(n38098), .Z(N62022) );
  XOR U47203 ( .A(n38118), .B(n38117), .Z(n38098) );
  XNOR U47204 ( .A(n38133), .B(n38134), .Z(n38117) );
  XNOR U47205 ( .A(n38128), .B(n38129), .Z(n38134) );
  XNOR U47206 ( .A(n38130), .B(n38131), .Z(n38129) );
  XNOR U47207 ( .A(y[2653]), .B(x[2653]), .Z(n38131) );
  XNOR U47208 ( .A(y[2654]), .B(x[2654]), .Z(n38130) );
  XNOR U47209 ( .A(y[2652]), .B(x[2652]), .Z(n38128) );
  XNOR U47210 ( .A(n38122), .B(n38123), .Z(n38133) );
  XNOR U47211 ( .A(y[2649]), .B(x[2649]), .Z(n38123) );
  XNOR U47212 ( .A(n38124), .B(n38125), .Z(n38122) );
  XNOR U47213 ( .A(y[2650]), .B(x[2650]), .Z(n38125) );
  XNOR U47214 ( .A(y[2651]), .B(x[2651]), .Z(n38124) );
  XNOR U47215 ( .A(n38115), .B(n38114), .Z(n38118) );
  XNOR U47216 ( .A(n38110), .B(n38111), .Z(n38114) );
  XNOR U47217 ( .A(y[2646]), .B(x[2646]), .Z(n38111) );
  XNOR U47218 ( .A(n38112), .B(n38113), .Z(n38110) );
  XNOR U47219 ( .A(y[2647]), .B(x[2647]), .Z(n38113) );
  XNOR U47220 ( .A(y[2648]), .B(x[2648]), .Z(n38112) );
  XNOR U47221 ( .A(n38104), .B(n38105), .Z(n38115) );
  XNOR U47222 ( .A(y[2643]), .B(x[2643]), .Z(n38105) );
  XNOR U47223 ( .A(n38106), .B(n38107), .Z(n38104) );
  XNOR U47224 ( .A(y[2644]), .B(x[2644]), .Z(n38107) );
  XNOR U47225 ( .A(y[2645]), .B(x[2645]), .Z(n38106) );
  XOR U47226 ( .A(n38080), .B(n38081), .Z(n38099) );
  XNOR U47227 ( .A(n38096), .B(n38097), .Z(n38081) );
  XNOR U47228 ( .A(n38091), .B(n38092), .Z(n38097) );
  XNOR U47229 ( .A(n38093), .B(n38094), .Z(n38092) );
  XNOR U47230 ( .A(y[2641]), .B(x[2641]), .Z(n38094) );
  XNOR U47231 ( .A(y[2642]), .B(x[2642]), .Z(n38093) );
  XNOR U47232 ( .A(y[2640]), .B(x[2640]), .Z(n38091) );
  XNOR U47233 ( .A(n38085), .B(n38086), .Z(n38096) );
  XNOR U47234 ( .A(y[2637]), .B(x[2637]), .Z(n38086) );
  XNOR U47235 ( .A(n38087), .B(n38088), .Z(n38085) );
  XNOR U47236 ( .A(y[2638]), .B(x[2638]), .Z(n38088) );
  XNOR U47237 ( .A(y[2639]), .B(x[2639]), .Z(n38087) );
  XOR U47238 ( .A(n38079), .B(n38078), .Z(n38080) );
  XNOR U47239 ( .A(n38074), .B(n38075), .Z(n38078) );
  XNOR U47240 ( .A(y[2634]), .B(x[2634]), .Z(n38075) );
  XNOR U47241 ( .A(n38076), .B(n38077), .Z(n38074) );
  XNOR U47242 ( .A(y[2635]), .B(x[2635]), .Z(n38077) );
  XNOR U47243 ( .A(y[2636]), .B(x[2636]), .Z(n38076) );
  XNOR U47244 ( .A(n38068), .B(n38069), .Z(n38079) );
  XNOR U47245 ( .A(y[2631]), .B(x[2631]), .Z(n38069) );
  XNOR U47246 ( .A(n38070), .B(n38071), .Z(n38068) );
  XNOR U47247 ( .A(y[2632]), .B(x[2632]), .Z(n38071) );
  XNOR U47248 ( .A(y[2633]), .B(x[2633]), .Z(n38070) );
  NAND U47249 ( .A(n38135), .B(n38136), .Z(N62013) );
  NANDN U47250 ( .A(n38137), .B(n38138), .Z(n38136) );
  OR U47251 ( .A(n38139), .B(n38140), .Z(n38138) );
  NAND U47252 ( .A(n38139), .B(n38140), .Z(n38135) );
  XOR U47253 ( .A(n38139), .B(n38141), .Z(N62012) );
  XNOR U47254 ( .A(n38137), .B(n38140), .Z(n38141) );
  AND U47255 ( .A(n38142), .B(n38143), .Z(n38140) );
  NANDN U47256 ( .A(n38144), .B(n38145), .Z(n38143) );
  NANDN U47257 ( .A(n38146), .B(n38147), .Z(n38145) );
  NANDN U47258 ( .A(n38147), .B(n38146), .Z(n38142) );
  NAND U47259 ( .A(n38148), .B(n38149), .Z(n38137) );
  NANDN U47260 ( .A(n38150), .B(n38151), .Z(n38149) );
  OR U47261 ( .A(n38152), .B(n38153), .Z(n38151) );
  NAND U47262 ( .A(n38153), .B(n38152), .Z(n38148) );
  AND U47263 ( .A(n38154), .B(n38155), .Z(n38139) );
  NANDN U47264 ( .A(n38156), .B(n38157), .Z(n38155) );
  NANDN U47265 ( .A(n38158), .B(n38159), .Z(n38157) );
  NANDN U47266 ( .A(n38159), .B(n38158), .Z(n38154) );
  XOR U47267 ( .A(n38153), .B(n38160), .Z(N62011) );
  XOR U47268 ( .A(n38150), .B(n38152), .Z(n38160) );
  XNOR U47269 ( .A(n38146), .B(n38161), .Z(n38152) );
  XNOR U47270 ( .A(n38144), .B(n38147), .Z(n38161) );
  NAND U47271 ( .A(n38162), .B(n38163), .Z(n38147) );
  NAND U47272 ( .A(n38164), .B(n38165), .Z(n38163) );
  OR U47273 ( .A(n38166), .B(n38167), .Z(n38164) );
  NANDN U47274 ( .A(n38168), .B(n38166), .Z(n38162) );
  IV U47275 ( .A(n38167), .Z(n38168) );
  NAND U47276 ( .A(n38169), .B(n38170), .Z(n38144) );
  NAND U47277 ( .A(n38171), .B(n38172), .Z(n38170) );
  NANDN U47278 ( .A(n38173), .B(n38174), .Z(n38171) );
  NANDN U47279 ( .A(n38174), .B(n38173), .Z(n38169) );
  AND U47280 ( .A(n38175), .B(n38176), .Z(n38146) );
  NAND U47281 ( .A(n38177), .B(n38178), .Z(n38176) );
  OR U47282 ( .A(n38179), .B(n38180), .Z(n38177) );
  NANDN U47283 ( .A(n38181), .B(n38179), .Z(n38175) );
  NAND U47284 ( .A(n38182), .B(n38183), .Z(n38150) );
  NANDN U47285 ( .A(n38184), .B(n38185), .Z(n38183) );
  OR U47286 ( .A(n38186), .B(n38187), .Z(n38185) );
  NANDN U47287 ( .A(n38188), .B(n38186), .Z(n38182) );
  IV U47288 ( .A(n38187), .Z(n38188) );
  XNOR U47289 ( .A(n38158), .B(n38189), .Z(n38153) );
  XNOR U47290 ( .A(n38156), .B(n38159), .Z(n38189) );
  NAND U47291 ( .A(n38190), .B(n38191), .Z(n38159) );
  NAND U47292 ( .A(n38192), .B(n38193), .Z(n38191) );
  OR U47293 ( .A(n38194), .B(n38195), .Z(n38192) );
  NANDN U47294 ( .A(n38196), .B(n38194), .Z(n38190) );
  IV U47295 ( .A(n38195), .Z(n38196) );
  NAND U47296 ( .A(n38197), .B(n38198), .Z(n38156) );
  NAND U47297 ( .A(n38199), .B(n38200), .Z(n38198) );
  NANDN U47298 ( .A(n38201), .B(n38202), .Z(n38199) );
  NANDN U47299 ( .A(n38202), .B(n38201), .Z(n38197) );
  AND U47300 ( .A(n38203), .B(n38204), .Z(n38158) );
  NAND U47301 ( .A(n38205), .B(n38206), .Z(n38204) );
  OR U47302 ( .A(n38207), .B(n38208), .Z(n38205) );
  NANDN U47303 ( .A(n38209), .B(n38207), .Z(n38203) );
  XNOR U47304 ( .A(n38184), .B(n38210), .Z(N62010) );
  XOR U47305 ( .A(n38186), .B(n38187), .Z(n38210) );
  XNOR U47306 ( .A(n38200), .B(n38211), .Z(n38187) );
  XOR U47307 ( .A(n38201), .B(n38202), .Z(n38211) );
  XOR U47308 ( .A(n38207), .B(n38212), .Z(n38202) );
  XOR U47309 ( .A(n38206), .B(n38209), .Z(n38212) );
  IV U47310 ( .A(n38208), .Z(n38209) );
  NAND U47311 ( .A(n38213), .B(n38214), .Z(n38208) );
  OR U47312 ( .A(n38215), .B(n38216), .Z(n38214) );
  OR U47313 ( .A(n38217), .B(n38218), .Z(n38213) );
  NAND U47314 ( .A(n38219), .B(n38220), .Z(n38206) );
  OR U47315 ( .A(n38221), .B(n38222), .Z(n38220) );
  OR U47316 ( .A(n38223), .B(n38224), .Z(n38219) );
  NOR U47317 ( .A(n38225), .B(n38226), .Z(n38207) );
  ANDN U47318 ( .B(n38227), .A(n38228), .Z(n38201) );
  XNOR U47319 ( .A(n38194), .B(n38229), .Z(n38200) );
  XNOR U47320 ( .A(n38193), .B(n38195), .Z(n38229) );
  NAND U47321 ( .A(n38230), .B(n38231), .Z(n38195) );
  OR U47322 ( .A(n38232), .B(n38233), .Z(n38231) );
  OR U47323 ( .A(n38234), .B(n38235), .Z(n38230) );
  NAND U47324 ( .A(n38236), .B(n38237), .Z(n38193) );
  OR U47325 ( .A(n38238), .B(n38239), .Z(n38237) );
  OR U47326 ( .A(n38240), .B(n38241), .Z(n38236) );
  ANDN U47327 ( .B(n38242), .A(n38243), .Z(n38194) );
  IV U47328 ( .A(n38244), .Z(n38242) );
  ANDN U47329 ( .B(n38245), .A(n38246), .Z(n38186) );
  XOR U47330 ( .A(n38172), .B(n38247), .Z(n38184) );
  XOR U47331 ( .A(n38173), .B(n38174), .Z(n38247) );
  XOR U47332 ( .A(n38179), .B(n38248), .Z(n38174) );
  XOR U47333 ( .A(n38178), .B(n38181), .Z(n38248) );
  IV U47334 ( .A(n38180), .Z(n38181) );
  NAND U47335 ( .A(n38249), .B(n38250), .Z(n38180) );
  OR U47336 ( .A(n38251), .B(n38252), .Z(n38250) );
  OR U47337 ( .A(n38253), .B(n38254), .Z(n38249) );
  NAND U47338 ( .A(n38255), .B(n38256), .Z(n38178) );
  OR U47339 ( .A(n38257), .B(n38258), .Z(n38256) );
  OR U47340 ( .A(n38259), .B(n38260), .Z(n38255) );
  NOR U47341 ( .A(n38261), .B(n38262), .Z(n38179) );
  ANDN U47342 ( .B(n38263), .A(n38264), .Z(n38173) );
  IV U47343 ( .A(n38265), .Z(n38263) );
  XNOR U47344 ( .A(n38166), .B(n38266), .Z(n38172) );
  XNOR U47345 ( .A(n38165), .B(n38167), .Z(n38266) );
  NAND U47346 ( .A(n38267), .B(n38268), .Z(n38167) );
  OR U47347 ( .A(n38269), .B(n38270), .Z(n38268) );
  OR U47348 ( .A(n38271), .B(n38272), .Z(n38267) );
  NAND U47349 ( .A(n38273), .B(n38274), .Z(n38165) );
  OR U47350 ( .A(n38275), .B(n38276), .Z(n38274) );
  OR U47351 ( .A(n38277), .B(n38278), .Z(n38273) );
  ANDN U47352 ( .B(n38279), .A(n38280), .Z(n38166) );
  IV U47353 ( .A(n38281), .Z(n38279) );
  XNOR U47354 ( .A(n38246), .B(n38245), .Z(N62009) );
  XOR U47355 ( .A(n38265), .B(n38264), .Z(n38245) );
  XNOR U47356 ( .A(n38280), .B(n38281), .Z(n38264) );
  XNOR U47357 ( .A(n38275), .B(n38276), .Z(n38281) );
  XNOR U47358 ( .A(n38277), .B(n38278), .Z(n38276) );
  XNOR U47359 ( .A(y[2629]), .B(x[2629]), .Z(n38278) );
  XNOR U47360 ( .A(y[2630]), .B(x[2630]), .Z(n38277) );
  XNOR U47361 ( .A(y[2628]), .B(x[2628]), .Z(n38275) );
  XNOR U47362 ( .A(n38269), .B(n38270), .Z(n38280) );
  XNOR U47363 ( .A(y[2625]), .B(x[2625]), .Z(n38270) );
  XNOR U47364 ( .A(n38271), .B(n38272), .Z(n38269) );
  XNOR U47365 ( .A(y[2626]), .B(x[2626]), .Z(n38272) );
  XNOR U47366 ( .A(y[2627]), .B(x[2627]), .Z(n38271) );
  XNOR U47367 ( .A(n38262), .B(n38261), .Z(n38265) );
  XNOR U47368 ( .A(n38257), .B(n38258), .Z(n38261) );
  XNOR U47369 ( .A(y[2622]), .B(x[2622]), .Z(n38258) );
  XNOR U47370 ( .A(n38259), .B(n38260), .Z(n38257) );
  XNOR U47371 ( .A(y[2623]), .B(x[2623]), .Z(n38260) );
  XNOR U47372 ( .A(y[2624]), .B(x[2624]), .Z(n38259) );
  XNOR U47373 ( .A(n38251), .B(n38252), .Z(n38262) );
  XNOR U47374 ( .A(y[2619]), .B(x[2619]), .Z(n38252) );
  XNOR U47375 ( .A(n38253), .B(n38254), .Z(n38251) );
  XNOR U47376 ( .A(y[2620]), .B(x[2620]), .Z(n38254) );
  XNOR U47377 ( .A(y[2621]), .B(x[2621]), .Z(n38253) );
  XOR U47378 ( .A(n38227), .B(n38228), .Z(n38246) );
  XNOR U47379 ( .A(n38243), .B(n38244), .Z(n38228) );
  XNOR U47380 ( .A(n38238), .B(n38239), .Z(n38244) );
  XNOR U47381 ( .A(n38240), .B(n38241), .Z(n38239) );
  XNOR U47382 ( .A(y[2617]), .B(x[2617]), .Z(n38241) );
  XNOR U47383 ( .A(y[2618]), .B(x[2618]), .Z(n38240) );
  XNOR U47384 ( .A(y[2616]), .B(x[2616]), .Z(n38238) );
  XNOR U47385 ( .A(n38232), .B(n38233), .Z(n38243) );
  XNOR U47386 ( .A(y[2613]), .B(x[2613]), .Z(n38233) );
  XNOR U47387 ( .A(n38234), .B(n38235), .Z(n38232) );
  XNOR U47388 ( .A(y[2614]), .B(x[2614]), .Z(n38235) );
  XNOR U47389 ( .A(y[2615]), .B(x[2615]), .Z(n38234) );
  XOR U47390 ( .A(n38226), .B(n38225), .Z(n38227) );
  XNOR U47391 ( .A(n38221), .B(n38222), .Z(n38225) );
  XNOR U47392 ( .A(y[2610]), .B(x[2610]), .Z(n38222) );
  XNOR U47393 ( .A(n38223), .B(n38224), .Z(n38221) );
  XNOR U47394 ( .A(y[2611]), .B(x[2611]), .Z(n38224) );
  XNOR U47395 ( .A(y[2612]), .B(x[2612]), .Z(n38223) );
  XNOR U47396 ( .A(n38215), .B(n38216), .Z(n38226) );
  XNOR U47397 ( .A(y[2607]), .B(x[2607]), .Z(n38216) );
  XNOR U47398 ( .A(n38217), .B(n38218), .Z(n38215) );
  XNOR U47399 ( .A(y[2608]), .B(x[2608]), .Z(n38218) );
  XNOR U47400 ( .A(y[2609]), .B(x[2609]), .Z(n38217) );
  NAND U47401 ( .A(n38282), .B(n38283), .Z(N62000) );
  NANDN U47402 ( .A(n38284), .B(n38285), .Z(n38283) );
  OR U47403 ( .A(n38286), .B(n38287), .Z(n38285) );
  NAND U47404 ( .A(n38286), .B(n38287), .Z(n38282) );
  XOR U47405 ( .A(n38286), .B(n38288), .Z(N61999) );
  XNOR U47406 ( .A(n38284), .B(n38287), .Z(n38288) );
  AND U47407 ( .A(n38289), .B(n38290), .Z(n38287) );
  NANDN U47408 ( .A(n38291), .B(n38292), .Z(n38290) );
  NANDN U47409 ( .A(n38293), .B(n38294), .Z(n38292) );
  NANDN U47410 ( .A(n38294), .B(n38293), .Z(n38289) );
  NAND U47411 ( .A(n38295), .B(n38296), .Z(n38284) );
  NANDN U47412 ( .A(n38297), .B(n38298), .Z(n38296) );
  OR U47413 ( .A(n38299), .B(n38300), .Z(n38298) );
  NAND U47414 ( .A(n38300), .B(n38299), .Z(n38295) );
  AND U47415 ( .A(n38301), .B(n38302), .Z(n38286) );
  NANDN U47416 ( .A(n38303), .B(n38304), .Z(n38302) );
  NANDN U47417 ( .A(n38305), .B(n38306), .Z(n38304) );
  NANDN U47418 ( .A(n38306), .B(n38305), .Z(n38301) );
  XOR U47419 ( .A(n38300), .B(n38307), .Z(N61998) );
  XOR U47420 ( .A(n38297), .B(n38299), .Z(n38307) );
  XNOR U47421 ( .A(n38293), .B(n38308), .Z(n38299) );
  XNOR U47422 ( .A(n38291), .B(n38294), .Z(n38308) );
  NAND U47423 ( .A(n38309), .B(n38310), .Z(n38294) );
  NAND U47424 ( .A(n38311), .B(n38312), .Z(n38310) );
  OR U47425 ( .A(n38313), .B(n38314), .Z(n38311) );
  NANDN U47426 ( .A(n38315), .B(n38313), .Z(n38309) );
  IV U47427 ( .A(n38314), .Z(n38315) );
  NAND U47428 ( .A(n38316), .B(n38317), .Z(n38291) );
  NAND U47429 ( .A(n38318), .B(n38319), .Z(n38317) );
  NANDN U47430 ( .A(n38320), .B(n38321), .Z(n38318) );
  NANDN U47431 ( .A(n38321), .B(n38320), .Z(n38316) );
  AND U47432 ( .A(n38322), .B(n38323), .Z(n38293) );
  NAND U47433 ( .A(n38324), .B(n38325), .Z(n38323) );
  OR U47434 ( .A(n38326), .B(n38327), .Z(n38324) );
  NANDN U47435 ( .A(n38328), .B(n38326), .Z(n38322) );
  NAND U47436 ( .A(n38329), .B(n38330), .Z(n38297) );
  NANDN U47437 ( .A(n38331), .B(n38332), .Z(n38330) );
  OR U47438 ( .A(n38333), .B(n38334), .Z(n38332) );
  NANDN U47439 ( .A(n38335), .B(n38333), .Z(n38329) );
  IV U47440 ( .A(n38334), .Z(n38335) );
  XNOR U47441 ( .A(n38305), .B(n38336), .Z(n38300) );
  XNOR U47442 ( .A(n38303), .B(n38306), .Z(n38336) );
  NAND U47443 ( .A(n38337), .B(n38338), .Z(n38306) );
  NAND U47444 ( .A(n38339), .B(n38340), .Z(n38338) );
  OR U47445 ( .A(n38341), .B(n38342), .Z(n38339) );
  NANDN U47446 ( .A(n38343), .B(n38341), .Z(n38337) );
  IV U47447 ( .A(n38342), .Z(n38343) );
  NAND U47448 ( .A(n38344), .B(n38345), .Z(n38303) );
  NAND U47449 ( .A(n38346), .B(n38347), .Z(n38345) );
  NANDN U47450 ( .A(n38348), .B(n38349), .Z(n38346) );
  NANDN U47451 ( .A(n38349), .B(n38348), .Z(n38344) );
  AND U47452 ( .A(n38350), .B(n38351), .Z(n38305) );
  NAND U47453 ( .A(n38352), .B(n38353), .Z(n38351) );
  OR U47454 ( .A(n38354), .B(n38355), .Z(n38352) );
  NANDN U47455 ( .A(n38356), .B(n38354), .Z(n38350) );
  XNOR U47456 ( .A(n38331), .B(n38357), .Z(N61997) );
  XOR U47457 ( .A(n38333), .B(n38334), .Z(n38357) );
  XNOR U47458 ( .A(n38347), .B(n38358), .Z(n38334) );
  XOR U47459 ( .A(n38348), .B(n38349), .Z(n38358) );
  XOR U47460 ( .A(n38354), .B(n38359), .Z(n38349) );
  XOR U47461 ( .A(n38353), .B(n38356), .Z(n38359) );
  IV U47462 ( .A(n38355), .Z(n38356) );
  NAND U47463 ( .A(n38360), .B(n38361), .Z(n38355) );
  OR U47464 ( .A(n38362), .B(n38363), .Z(n38361) );
  OR U47465 ( .A(n38364), .B(n38365), .Z(n38360) );
  NAND U47466 ( .A(n38366), .B(n38367), .Z(n38353) );
  OR U47467 ( .A(n38368), .B(n38369), .Z(n38367) );
  OR U47468 ( .A(n38370), .B(n38371), .Z(n38366) );
  NOR U47469 ( .A(n38372), .B(n38373), .Z(n38354) );
  ANDN U47470 ( .B(n38374), .A(n38375), .Z(n38348) );
  XNOR U47471 ( .A(n38341), .B(n38376), .Z(n38347) );
  XNOR U47472 ( .A(n38340), .B(n38342), .Z(n38376) );
  NAND U47473 ( .A(n38377), .B(n38378), .Z(n38342) );
  OR U47474 ( .A(n38379), .B(n38380), .Z(n38378) );
  OR U47475 ( .A(n38381), .B(n38382), .Z(n38377) );
  NAND U47476 ( .A(n38383), .B(n38384), .Z(n38340) );
  OR U47477 ( .A(n38385), .B(n38386), .Z(n38384) );
  OR U47478 ( .A(n38387), .B(n38388), .Z(n38383) );
  ANDN U47479 ( .B(n38389), .A(n38390), .Z(n38341) );
  IV U47480 ( .A(n38391), .Z(n38389) );
  ANDN U47481 ( .B(n38392), .A(n38393), .Z(n38333) );
  XOR U47482 ( .A(n38319), .B(n38394), .Z(n38331) );
  XOR U47483 ( .A(n38320), .B(n38321), .Z(n38394) );
  XOR U47484 ( .A(n38326), .B(n38395), .Z(n38321) );
  XOR U47485 ( .A(n38325), .B(n38328), .Z(n38395) );
  IV U47486 ( .A(n38327), .Z(n38328) );
  NAND U47487 ( .A(n38396), .B(n38397), .Z(n38327) );
  OR U47488 ( .A(n38398), .B(n38399), .Z(n38397) );
  OR U47489 ( .A(n38400), .B(n38401), .Z(n38396) );
  NAND U47490 ( .A(n38402), .B(n38403), .Z(n38325) );
  OR U47491 ( .A(n38404), .B(n38405), .Z(n38403) );
  OR U47492 ( .A(n38406), .B(n38407), .Z(n38402) );
  NOR U47493 ( .A(n38408), .B(n38409), .Z(n38326) );
  ANDN U47494 ( .B(n38410), .A(n38411), .Z(n38320) );
  IV U47495 ( .A(n38412), .Z(n38410) );
  XNOR U47496 ( .A(n38313), .B(n38413), .Z(n38319) );
  XNOR U47497 ( .A(n38312), .B(n38314), .Z(n38413) );
  NAND U47498 ( .A(n38414), .B(n38415), .Z(n38314) );
  OR U47499 ( .A(n38416), .B(n38417), .Z(n38415) );
  OR U47500 ( .A(n38418), .B(n38419), .Z(n38414) );
  NAND U47501 ( .A(n38420), .B(n38421), .Z(n38312) );
  OR U47502 ( .A(n38422), .B(n38423), .Z(n38421) );
  OR U47503 ( .A(n38424), .B(n38425), .Z(n38420) );
  ANDN U47504 ( .B(n38426), .A(n38427), .Z(n38313) );
  IV U47505 ( .A(n38428), .Z(n38426) );
  XNOR U47506 ( .A(n38393), .B(n38392), .Z(N61996) );
  XOR U47507 ( .A(n38412), .B(n38411), .Z(n38392) );
  XNOR U47508 ( .A(n38427), .B(n38428), .Z(n38411) );
  XNOR U47509 ( .A(n38422), .B(n38423), .Z(n38428) );
  XNOR U47510 ( .A(n38424), .B(n38425), .Z(n38423) );
  XNOR U47511 ( .A(y[2605]), .B(x[2605]), .Z(n38425) );
  XNOR U47512 ( .A(y[2606]), .B(x[2606]), .Z(n38424) );
  XNOR U47513 ( .A(y[2604]), .B(x[2604]), .Z(n38422) );
  XNOR U47514 ( .A(n38416), .B(n38417), .Z(n38427) );
  XNOR U47515 ( .A(y[2601]), .B(x[2601]), .Z(n38417) );
  XNOR U47516 ( .A(n38418), .B(n38419), .Z(n38416) );
  XNOR U47517 ( .A(y[2602]), .B(x[2602]), .Z(n38419) );
  XNOR U47518 ( .A(y[2603]), .B(x[2603]), .Z(n38418) );
  XNOR U47519 ( .A(n38409), .B(n38408), .Z(n38412) );
  XNOR U47520 ( .A(n38404), .B(n38405), .Z(n38408) );
  XNOR U47521 ( .A(y[2598]), .B(x[2598]), .Z(n38405) );
  XNOR U47522 ( .A(n38406), .B(n38407), .Z(n38404) );
  XNOR U47523 ( .A(y[2599]), .B(x[2599]), .Z(n38407) );
  XNOR U47524 ( .A(y[2600]), .B(x[2600]), .Z(n38406) );
  XNOR U47525 ( .A(n38398), .B(n38399), .Z(n38409) );
  XNOR U47526 ( .A(y[2595]), .B(x[2595]), .Z(n38399) );
  XNOR U47527 ( .A(n38400), .B(n38401), .Z(n38398) );
  XNOR U47528 ( .A(y[2596]), .B(x[2596]), .Z(n38401) );
  XNOR U47529 ( .A(y[2597]), .B(x[2597]), .Z(n38400) );
  XOR U47530 ( .A(n38374), .B(n38375), .Z(n38393) );
  XNOR U47531 ( .A(n38390), .B(n38391), .Z(n38375) );
  XNOR U47532 ( .A(n38385), .B(n38386), .Z(n38391) );
  XNOR U47533 ( .A(n38387), .B(n38388), .Z(n38386) );
  XNOR U47534 ( .A(y[2593]), .B(x[2593]), .Z(n38388) );
  XNOR U47535 ( .A(y[2594]), .B(x[2594]), .Z(n38387) );
  XNOR U47536 ( .A(y[2592]), .B(x[2592]), .Z(n38385) );
  XNOR U47537 ( .A(n38379), .B(n38380), .Z(n38390) );
  XNOR U47538 ( .A(y[2589]), .B(x[2589]), .Z(n38380) );
  XNOR U47539 ( .A(n38381), .B(n38382), .Z(n38379) );
  XNOR U47540 ( .A(y[2590]), .B(x[2590]), .Z(n38382) );
  XNOR U47541 ( .A(y[2591]), .B(x[2591]), .Z(n38381) );
  XOR U47542 ( .A(n38373), .B(n38372), .Z(n38374) );
  XNOR U47543 ( .A(n38368), .B(n38369), .Z(n38372) );
  XNOR U47544 ( .A(y[2586]), .B(x[2586]), .Z(n38369) );
  XNOR U47545 ( .A(n38370), .B(n38371), .Z(n38368) );
  XNOR U47546 ( .A(y[2587]), .B(x[2587]), .Z(n38371) );
  XNOR U47547 ( .A(y[2588]), .B(x[2588]), .Z(n38370) );
  XNOR U47548 ( .A(n38362), .B(n38363), .Z(n38373) );
  XNOR U47549 ( .A(y[2583]), .B(x[2583]), .Z(n38363) );
  XNOR U47550 ( .A(n38364), .B(n38365), .Z(n38362) );
  XNOR U47551 ( .A(y[2584]), .B(x[2584]), .Z(n38365) );
  XNOR U47552 ( .A(y[2585]), .B(x[2585]), .Z(n38364) );
  NAND U47553 ( .A(n38429), .B(n38430), .Z(N61987) );
  NANDN U47554 ( .A(n38431), .B(n38432), .Z(n38430) );
  OR U47555 ( .A(n38433), .B(n38434), .Z(n38432) );
  NAND U47556 ( .A(n38433), .B(n38434), .Z(n38429) );
  XOR U47557 ( .A(n38433), .B(n38435), .Z(N61986) );
  XNOR U47558 ( .A(n38431), .B(n38434), .Z(n38435) );
  AND U47559 ( .A(n38436), .B(n38437), .Z(n38434) );
  NANDN U47560 ( .A(n38438), .B(n38439), .Z(n38437) );
  NANDN U47561 ( .A(n38440), .B(n38441), .Z(n38439) );
  NANDN U47562 ( .A(n38441), .B(n38440), .Z(n38436) );
  NAND U47563 ( .A(n38442), .B(n38443), .Z(n38431) );
  NANDN U47564 ( .A(n38444), .B(n38445), .Z(n38443) );
  OR U47565 ( .A(n38446), .B(n38447), .Z(n38445) );
  NAND U47566 ( .A(n38447), .B(n38446), .Z(n38442) );
  AND U47567 ( .A(n38448), .B(n38449), .Z(n38433) );
  NANDN U47568 ( .A(n38450), .B(n38451), .Z(n38449) );
  NANDN U47569 ( .A(n38452), .B(n38453), .Z(n38451) );
  NANDN U47570 ( .A(n38453), .B(n38452), .Z(n38448) );
  XOR U47571 ( .A(n38447), .B(n38454), .Z(N61985) );
  XOR U47572 ( .A(n38444), .B(n38446), .Z(n38454) );
  XNOR U47573 ( .A(n38440), .B(n38455), .Z(n38446) );
  XNOR U47574 ( .A(n38438), .B(n38441), .Z(n38455) );
  NAND U47575 ( .A(n38456), .B(n38457), .Z(n38441) );
  NAND U47576 ( .A(n38458), .B(n38459), .Z(n38457) );
  OR U47577 ( .A(n38460), .B(n38461), .Z(n38458) );
  NANDN U47578 ( .A(n38462), .B(n38460), .Z(n38456) );
  IV U47579 ( .A(n38461), .Z(n38462) );
  NAND U47580 ( .A(n38463), .B(n38464), .Z(n38438) );
  NAND U47581 ( .A(n38465), .B(n38466), .Z(n38464) );
  NANDN U47582 ( .A(n38467), .B(n38468), .Z(n38465) );
  NANDN U47583 ( .A(n38468), .B(n38467), .Z(n38463) );
  AND U47584 ( .A(n38469), .B(n38470), .Z(n38440) );
  NAND U47585 ( .A(n38471), .B(n38472), .Z(n38470) );
  OR U47586 ( .A(n38473), .B(n38474), .Z(n38471) );
  NANDN U47587 ( .A(n38475), .B(n38473), .Z(n38469) );
  NAND U47588 ( .A(n38476), .B(n38477), .Z(n38444) );
  NANDN U47589 ( .A(n38478), .B(n38479), .Z(n38477) );
  OR U47590 ( .A(n38480), .B(n38481), .Z(n38479) );
  NANDN U47591 ( .A(n38482), .B(n38480), .Z(n38476) );
  IV U47592 ( .A(n38481), .Z(n38482) );
  XNOR U47593 ( .A(n38452), .B(n38483), .Z(n38447) );
  XNOR U47594 ( .A(n38450), .B(n38453), .Z(n38483) );
  NAND U47595 ( .A(n38484), .B(n38485), .Z(n38453) );
  NAND U47596 ( .A(n38486), .B(n38487), .Z(n38485) );
  OR U47597 ( .A(n38488), .B(n38489), .Z(n38486) );
  NANDN U47598 ( .A(n38490), .B(n38488), .Z(n38484) );
  IV U47599 ( .A(n38489), .Z(n38490) );
  NAND U47600 ( .A(n38491), .B(n38492), .Z(n38450) );
  NAND U47601 ( .A(n38493), .B(n38494), .Z(n38492) );
  NANDN U47602 ( .A(n38495), .B(n38496), .Z(n38493) );
  NANDN U47603 ( .A(n38496), .B(n38495), .Z(n38491) );
  AND U47604 ( .A(n38497), .B(n38498), .Z(n38452) );
  NAND U47605 ( .A(n38499), .B(n38500), .Z(n38498) );
  OR U47606 ( .A(n38501), .B(n38502), .Z(n38499) );
  NANDN U47607 ( .A(n38503), .B(n38501), .Z(n38497) );
  XNOR U47608 ( .A(n38478), .B(n38504), .Z(N61984) );
  XOR U47609 ( .A(n38480), .B(n38481), .Z(n38504) );
  XNOR U47610 ( .A(n38494), .B(n38505), .Z(n38481) );
  XOR U47611 ( .A(n38495), .B(n38496), .Z(n38505) );
  XOR U47612 ( .A(n38501), .B(n38506), .Z(n38496) );
  XOR U47613 ( .A(n38500), .B(n38503), .Z(n38506) );
  IV U47614 ( .A(n38502), .Z(n38503) );
  NAND U47615 ( .A(n38507), .B(n38508), .Z(n38502) );
  OR U47616 ( .A(n38509), .B(n38510), .Z(n38508) );
  OR U47617 ( .A(n38511), .B(n38512), .Z(n38507) );
  NAND U47618 ( .A(n38513), .B(n38514), .Z(n38500) );
  OR U47619 ( .A(n38515), .B(n38516), .Z(n38514) );
  OR U47620 ( .A(n38517), .B(n38518), .Z(n38513) );
  NOR U47621 ( .A(n38519), .B(n38520), .Z(n38501) );
  ANDN U47622 ( .B(n38521), .A(n38522), .Z(n38495) );
  XNOR U47623 ( .A(n38488), .B(n38523), .Z(n38494) );
  XNOR U47624 ( .A(n38487), .B(n38489), .Z(n38523) );
  NAND U47625 ( .A(n38524), .B(n38525), .Z(n38489) );
  OR U47626 ( .A(n38526), .B(n38527), .Z(n38525) );
  OR U47627 ( .A(n38528), .B(n38529), .Z(n38524) );
  NAND U47628 ( .A(n38530), .B(n38531), .Z(n38487) );
  OR U47629 ( .A(n38532), .B(n38533), .Z(n38531) );
  OR U47630 ( .A(n38534), .B(n38535), .Z(n38530) );
  ANDN U47631 ( .B(n38536), .A(n38537), .Z(n38488) );
  IV U47632 ( .A(n38538), .Z(n38536) );
  ANDN U47633 ( .B(n38539), .A(n38540), .Z(n38480) );
  XOR U47634 ( .A(n38466), .B(n38541), .Z(n38478) );
  XOR U47635 ( .A(n38467), .B(n38468), .Z(n38541) );
  XOR U47636 ( .A(n38473), .B(n38542), .Z(n38468) );
  XOR U47637 ( .A(n38472), .B(n38475), .Z(n38542) );
  IV U47638 ( .A(n38474), .Z(n38475) );
  NAND U47639 ( .A(n38543), .B(n38544), .Z(n38474) );
  OR U47640 ( .A(n38545), .B(n38546), .Z(n38544) );
  OR U47641 ( .A(n38547), .B(n38548), .Z(n38543) );
  NAND U47642 ( .A(n38549), .B(n38550), .Z(n38472) );
  OR U47643 ( .A(n38551), .B(n38552), .Z(n38550) );
  OR U47644 ( .A(n38553), .B(n38554), .Z(n38549) );
  NOR U47645 ( .A(n38555), .B(n38556), .Z(n38473) );
  ANDN U47646 ( .B(n38557), .A(n38558), .Z(n38467) );
  IV U47647 ( .A(n38559), .Z(n38557) );
  XNOR U47648 ( .A(n38460), .B(n38560), .Z(n38466) );
  XNOR U47649 ( .A(n38459), .B(n38461), .Z(n38560) );
  NAND U47650 ( .A(n38561), .B(n38562), .Z(n38461) );
  OR U47651 ( .A(n38563), .B(n38564), .Z(n38562) );
  OR U47652 ( .A(n38565), .B(n38566), .Z(n38561) );
  NAND U47653 ( .A(n38567), .B(n38568), .Z(n38459) );
  OR U47654 ( .A(n38569), .B(n38570), .Z(n38568) );
  OR U47655 ( .A(n38571), .B(n38572), .Z(n38567) );
  ANDN U47656 ( .B(n38573), .A(n38574), .Z(n38460) );
  IV U47657 ( .A(n38575), .Z(n38573) );
  XNOR U47658 ( .A(n38540), .B(n38539), .Z(N61983) );
  XOR U47659 ( .A(n38559), .B(n38558), .Z(n38539) );
  XNOR U47660 ( .A(n38574), .B(n38575), .Z(n38558) );
  XNOR U47661 ( .A(n38569), .B(n38570), .Z(n38575) );
  XNOR U47662 ( .A(n38571), .B(n38572), .Z(n38570) );
  XNOR U47663 ( .A(y[2581]), .B(x[2581]), .Z(n38572) );
  XNOR U47664 ( .A(y[2582]), .B(x[2582]), .Z(n38571) );
  XNOR U47665 ( .A(y[2580]), .B(x[2580]), .Z(n38569) );
  XNOR U47666 ( .A(n38563), .B(n38564), .Z(n38574) );
  XNOR U47667 ( .A(y[2577]), .B(x[2577]), .Z(n38564) );
  XNOR U47668 ( .A(n38565), .B(n38566), .Z(n38563) );
  XNOR U47669 ( .A(y[2578]), .B(x[2578]), .Z(n38566) );
  XNOR U47670 ( .A(y[2579]), .B(x[2579]), .Z(n38565) );
  XNOR U47671 ( .A(n38556), .B(n38555), .Z(n38559) );
  XNOR U47672 ( .A(n38551), .B(n38552), .Z(n38555) );
  XNOR U47673 ( .A(y[2574]), .B(x[2574]), .Z(n38552) );
  XNOR U47674 ( .A(n38553), .B(n38554), .Z(n38551) );
  XNOR U47675 ( .A(y[2575]), .B(x[2575]), .Z(n38554) );
  XNOR U47676 ( .A(y[2576]), .B(x[2576]), .Z(n38553) );
  XNOR U47677 ( .A(n38545), .B(n38546), .Z(n38556) );
  XNOR U47678 ( .A(y[2571]), .B(x[2571]), .Z(n38546) );
  XNOR U47679 ( .A(n38547), .B(n38548), .Z(n38545) );
  XNOR U47680 ( .A(y[2572]), .B(x[2572]), .Z(n38548) );
  XNOR U47681 ( .A(y[2573]), .B(x[2573]), .Z(n38547) );
  XOR U47682 ( .A(n38521), .B(n38522), .Z(n38540) );
  XNOR U47683 ( .A(n38537), .B(n38538), .Z(n38522) );
  XNOR U47684 ( .A(n38532), .B(n38533), .Z(n38538) );
  XNOR U47685 ( .A(n38534), .B(n38535), .Z(n38533) );
  XNOR U47686 ( .A(y[2569]), .B(x[2569]), .Z(n38535) );
  XNOR U47687 ( .A(y[2570]), .B(x[2570]), .Z(n38534) );
  XNOR U47688 ( .A(y[2568]), .B(x[2568]), .Z(n38532) );
  XNOR U47689 ( .A(n38526), .B(n38527), .Z(n38537) );
  XNOR U47690 ( .A(y[2565]), .B(x[2565]), .Z(n38527) );
  XNOR U47691 ( .A(n38528), .B(n38529), .Z(n38526) );
  XNOR U47692 ( .A(y[2566]), .B(x[2566]), .Z(n38529) );
  XNOR U47693 ( .A(y[2567]), .B(x[2567]), .Z(n38528) );
  XOR U47694 ( .A(n38520), .B(n38519), .Z(n38521) );
  XNOR U47695 ( .A(n38515), .B(n38516), .Z(n38519) );
  XNOR U47696 ( .A(y[2562]), .B(x[2562]), .Z(n38516) );
  XNOR U47697 ( .A(n38517), .B(n38518), .Z(n38515) );
  XNOR U47698 ( .A(y[2563]), .B(x[2563]), .Z(n38518) );
  XNOR U47699 ( .A(y[2564]), .B(x[2564]), .Z(n38517) );
  XNOR U47700 ( .A(n38509), .B(n38510), .Z(n38520) );
  XNOR U47701 ( .A(y[2559]), .B(x[2559]), .Z(n38510) );
  XNOR U47702 ( .A(n38511), .B(n38512), .Z(n38509) );
  XNOR U47703 ( .A(y[2560]), .B(x[2560]), .Z(n38512) );
  XNOR U47704 ( .A(y[2561]), .B(x[2561]), .Z(n38511) );
  NAND U47705 ( .A(n38576), .B(n38577), .Z(N61974) );
  NANDN U47706 ( .A(n38578), .B(n38579), .Z(n38577) );
  OR U47707 ( .A(n38580), .B(n38581), .Z(n38579) );
  NAND U47708 ( .A(n38580), .B(n38581), .Z(n38576) );
  XOR U47709 ( .A(n38580), .B(n38582), .Z(N61973) );
  XNOR U47710 ( .A(n38578), .B(n38581), .Z(n38582) );
  AND U47711 ( .A(n38583), .B(n38584), .Z(n38581) );
  NANDN U47712 ( .A(n38585), .B(n38586), .Z(n38584) );
  NANDN U47713 ( .A(n38587), .B(n38588), .Z(n38586) );
  NANDN U47714 ( .A(n38588), .B(n38587), .Z(n38583) );
  NAND U47715 ( .A(n38589), .B(n38590), .Z(n38578) );
  NANDN U47716 ( .A(n38591), .B(n38592), .Z(n38590) );
  OR U47717 ( .A(n38593), .B(n38594), .Z(n38592) );
  NAND U47718 ( .A(n38594), .B(n38593), .Z(n38589) );
  AND U47719 ( .A(n38595), .B(n38596), .Z(n38580) );
  NANDN U47720 ( .A(n38597), .B(n38598), .Z(n38596) );
  NANDN U47721 ( .A(n38599), .B(n38600), .Z(n38598) );
  NANDN U47722 ( .A(n38600), .B(n38599), .Z(n38595) );
  XOR U47723 ( .A(n38594), .B(n38601), .Z(N61972) );
  XOR U47724 ( .A(n38591), .B(n38593), .Z(n38601) );
  XNOR U47725 ( .A(n38587), .B(n38602), .Z(n38593) );
  XNOR U47726 ( .A(n38585), .B(n38588), .Z(n38602) );
  NAND U47727 ( .A(n38603), .B(n38604), .Z(n38588) );
  NAND U47728 ( .A(n38605), .B(n38606), .Z(n38604) );
  OR U47729 ( .A(n38607), .B(n38608), .Z(n38605) );
  NANDN U47730 ( .A(n38609), .B(n38607), .Z(n38603) );
  IV U47731 ( .A(n38608), .Z(n38609) );
  NAND U47732 ( .A(n38610), .B(n38611), .Z(n38585) );
  NAND U47733 ( .A(n38612), .B(n38613), .Z(n38611) );
  NANDN U47734 ( .A(n38614), .B(n38615), .Z(n38612) );
  NANDN U47735 ( .A(n38615), .B(n38614), .Z(n38610) );
  AND U47736 ( .A(n38616), .B(n38617), .Z(n38587) );
  NAND U47737 ( .A(n38618), .B(n38619), .Z(n38617) );
  OR U47738 ( .A(n38620), .B(n38621), .Z(n38618) );
  NANDN U47739 ( .A(n38622), .B(n38620), .Z(n38616) );
  NAND U47740 ( .A(n38623), .B(n38624), .Z(n38591) );
  NANDN U47741 ( .A(n38625), .B(n38626), .Z(n38624) );
  OR U47742 ( .A(n38627), .B(n38628), .Z(n38626) );
  NANDN U47743 ( .A(n38629), .B(n38627), .Z(n38623) );
  IV U47744 ( .A(n38628), .Z(n38629) );
  XNOR U47745 ( .A(n38599), .B(n38630), .Z(n38594) );
  XNOR U47746 ( .A(n38597), .B(n38600), .Z(n38630) );
  NAND U47747 ( .A(n38631), .B(n38632), .Z(n38600) );
  NAND U47748 ( .A(n38633), .B(n38634), .Z(n38632) );
  OR U47749 ( .A(n38635), .B(n38636), .Z(n38633) );
  NANDN U47750 ( .A(n38637), .B(n38635), .Z(n38631) );
  IV U47751 ( .A(n38636), .Z(n38637) );
  NAND U47752 ( .A(n38638), .B(n38639), .Z(n38597) );
  NAND U47753 ( .A(n38640), .B(n38641), .Z(n38639) );
  NANDN U47754 ( .A(n38642), .B(n38643), .Z(n38640) );
  NANDN U47755 ( .A(n38643), .B(n38642), .Z(n38638) );
  AND U47756 ( .A(n38644), .B(n38645), .Z(n38599) );
  NAND U47757 ( .A(n38646), .B(n38647), .Z(n38645) );
  OR U47758 ( .A(n38648), .B(n38649), .Z(n38646) );
  NANDN U47759 ( .A(n38650), .B(n38648), .Z(n38644) );
  XNOR U47760 ( .A(n38625), .B(n38651), .Z(N61971) );
  XOR U47761 ( .A(n38627), .B(n38628), .Z(n38651) );
  XNOR U47762 ( .A(n38641), .B(n38652), .Z(n38628) );
  XOR U47763 ( .A(n38642), .B(n38643), .Z(n38652) );
  XOR U47764 ( .A(n38648), .B(n38653), .Z(n38643) );
  XOR U47765 ( .A(n38647), .B(n38650), .Z(n38653) );
  IV U47766 ( .A(n38649), .Z(n38650) );
  NAND U47767 ( .A(n38654), .B(n38655), .Z(n38649) );
  OR U47768 ( .A(n38656), .B(n38657), .Z(n38655) );
  OR U47769 ( .A(n38658), .B(n38659), .Z(n38654) );
  NAND U47770 ( .A(n38660), .B(n38661), .Z(n38647) );
  OR U47771 ( .A(n38662), .B(n38663), .Z(n38661) );
  OR U47772 ( .A(n38664), .B(n38665), .Z(n38660) );
  NOR U47773 ( .A(n38666), .B(n38667), .Z(n38648) );
  ANDN U47774 ( .B(n38668), .A(n38669), .Z(n38642) );
  XNOR U47775 ( .A(n38635), .B(n38670), .Z(n38641) );
  XNOR U47776 ( .A(n38634), .B(n38636), .Z(n38670) );
  NAND U47777 ( .A(n38671), .B(n38672), .Z(n38636) );
  OR U47778 ( .A(n38673), .B(n38674), .Z(n38672) );
  OR U47779 ( .A(n38675), .B(n38676), .Z(n38671) );
  NAND U47780 ( .A(n38677), .B(n38678), .Z(n38634) );
  OR U47781 ( .A(n38679), .B(n38680), .Z(n38678) );
  OR U47782 ( .A(n38681), .B(n38682), .Z(n38677) );
  ANDN U47783 ( .B(n38683), .A(n38684), .Z(n38635) );
  IV U47784 ( .A(n38685), .Z(n38683) );
  ANDN U47785 ( .B(n38686), .A(n38687), .Z(n38627) );
  XOR U47786 ( .A(n38613), .B(n38688), .Z(n38625) );
  XOR U47787 ( .A(n38614), .B(n38615), .Z(n38688) );
  XOR U47788 ( .A(n38620), .B(n38689), .Z(n38615) );
  XOR U47789 ( .A(n38619), .B(n38622), .Z(n38689) );
  IV U47790 ( .A(n38621), .Z(n38622) );
  NAND U47791 ( .A(n38690), .B(n38691), .Z(n38621) );
  OR U47792 ( .A(n38692), .B(n38693), .Z(n38691) );
  OR U47793 ( .A(n38694), .B(n38695), .Z(n38690) );
  NAND U47794 ( .A(n38696), .B(n38697), .Z(n38619) );
  OR U47795 ( .A(n38698), .B(n38699), .Z(n38697) );
  OR U47796 ( .A(n38700), .B(n38701), .Z(n38696) );
  NOR U47797 ( .A(n38702), .B(n38703), .Z(n38620) );
  ANDN U47798 ( .B(n38704), .A(n38705), .Z(n38614) );
  IV U47799 ( .A(n38706), .Z(n38704) );
  XNOR U47800 ( .A(n38607), .B(n38707), .Z(n38613) );
  XNOR U47801 ( .A(n38606), .B(n38608), .Z(n38707) );
  NAND U47802 ( .A(n38708), .B(n38709), .Z(n38608) );
  OR U47803 ( .A(n38710), .B(n38711), .Z(n38709) );
  OR U47804 ( .A(n38712), .B(n38713), .Z(n38708) );
  NAND U47805 ( .A(n38714), .B(n38715), .Z(n38606) );
  OR U47806 ( .A(n38716), .B(n38717), .Z(n38715) );
  OR U47807 ( .A(n38718), .B(n38719), .Z(n38714) );
  ANDN U47808 ( .B(n38720), .A(n38721), .Z(n38607) );
  IV U47809 ( .A(n38722), .Z(n38720) );
  XNOR U47810 ( .A(n38687), .B(n38686), .Z(N61970) );
  XOR U47811 ( .A(n38706), .B(n38705), .Z(n38686) );
  XNOR U47812 ( .A(n38721), .B(n38722), .Z(n38705) );
  XNOR U47813 ( .A(n38716), .B(n38717), .Z(n38722) );
  XNOR U47814 ( .A(n38718), .B(n38719), .Z(n38717) );
  XNOR U47815 ( .A(y[2557]), .B(x[2557]), .Z(n38719) );
  XNOR U47816 ( .A(y[2558]), .B(x[2558]), .Z(n38718) );
  XNOR U47817 ( .A(y[2556]), .B(x[2556]), .Z(n38716) );
  XNOR U47818 ( .A(n38710), .B(n38711), .Z(n38721) );
  XNOR U47819 ( .A(y[2553]), .B(x[2553]), .Z(n38711) );
  XNOR U47820 ( .A(n38712), .B(n38713), .Z(n38710) );
  XNOR U47821 ( .A(y[2554]), .B(x[2554]), .Z(n38713) );
  XNOR U47822 ( .A(y[2555]), .B(x[2555]), .Z(n38712) );
  XNOR U47823 ( .A(n38703), .B(n38702), .Z(n38706) );
  XNOR U47824 ( .A(n38698), .B(n38699), .Z(n38702) );
  XNOR U47825 ( .A(y[2550]), .B(x[2550]), .Z(n38699) );
  XNOR U47826 ( .A(n38700), .B(n38701), .Z(n38698) );
  XNOR U47827 ( .A(y[2551]), .B(x[2551]), .Z(n38701) );
  XNOR U47828 ( .A(y[2552]), .B(x[2552]), .Z(n38700) );
  XNOR U47829 ( .A(n38692), .B(n38693), .Z(n38703) );
  XNOR U47830 ( .A(y[2547]), .B(x[2547]), .Z(n38693) );
  XNOR U47831 ( .A(n38694), .B(n38695), .Z(n38692) );
  XNOR U47832 ( .A(y[2548]), .B(x[2548]), .Z(n38695) );
  XNOR U47833 ( .A(y[2549]), .B(x[2549]), .Z(n38694) );
  XOR U47834 ( .A(n38668), .B(n38669), .Z(n38687) );
  XNOR U47835 ( .A(n38684), .B(n38685), .Z(n38669) );
  XNOR U47836 ( .A(n38679), .B(n38680), .Z(n38685) );
  XNOR U47837 ( .A(n38681), .B(n38682), .Z(n38680) );
  XNOR U47838 ( .A(y[2545]), .B(x[2545]), .Z(n38682) );
  XNOR U47839 ( .A(y[2546]), .B(x[2546]), .Z(n38681) );
  XNOR U47840 ( .A(y[2544]), .B(x[2544]), .Z(n38679) );
  XNOR U47841 ( .A(n38673), .B(n38674), .Z(n38684) );
  XNOR U47842 ( .A(y[2541]), .B(x[2541]), .Z(n38674) );
  XNOR U47843 ( .A(n38675), .B(n38676), .Z(n38673) );
  XNOR U47844 ( .A(y[2542]), .B(x[2542]), .Z(n38676) );
  XNOR U47845 ( .A(y[2543]), .B(x[2543]), .Z(n38675) );
  XOR U47846 ( .A(n38667), .B(n38666), .Z(n38668) );
  XNOR U47847 ( .A(n38662), .B(n38663), .Z(n38666) );
  XNOR U47848 ( .A(y[2538]), .B(x[2538]), .Z(n38663) );
  XNOR U47849 ( .A(n38664), .B(n38665), .Z(n38662) );
  XNOR U47850 ( .A(y[2539]), .B(x[2539]), .Z(n38665) );
  XNOR U47851 ( .A(y[2540]), .B(x[2540]), .Z(n38664) );
  XNOR U47852 ( .A(n38656), .B(n38657), .Z(n38667) );
  XNOR U47853 ( .A(y[2535]), .B(x[2535]), .Z(n38657) );
  XNOR U47854 ( .A(n38658), .B(n38659), .Z(n38656) );
  XNOR U47855 ( .A(y[2536]), .B(x[2536]), .Z(n38659) );
  XNOR U47856 ( .A(y[2537]), .B(x[2537]), .Z(n38658) );
  NAND U47857 ( .A(n38723), .B(n38724), .Z(N61961) );
  NANDN U47858 ( .A(n38725), .B(n38726), .Z(n38724) );
  OR U47859 ( .A(n38727), .B(n38728), .Z(n38726) );
  NAND U47860 ( .A(n38727), .B(n38728), .Z(n38723) );
  XOR U47861 ( .A(n38727), .B(n38729), .Z(N61960) );
  XNOR U47862 ( .A(n38725), .B(n38728), .Z(n38729) );
  AND U47863 ( .A(n38730), .B(n38731), .Z(n38728) );
  NANDN U47864 ( .A(n38732), .B(n38733), .Z(n38731) );
  NANDN U47865 ( .A(n38734), .B(n38735), .Z(n38733) );
  NANDN U47866 ( .A(n38735), .B(n38734), .Z(n38730) );
  NAND U47867 ( .A(n38736), .B(n38737), .Z(n38725) );
  NANDN U47868 ( .A(n38738), .B(n38739), .Z(n38737) );
  OR U47869 ( .A(n38740), .B(n38741), .Z(n38739) );
  NAND U47870 ( .A(n38741), .B(n38740), .Z(n38736) );
  AND U47871 ( .A(n38742), .B(n38743), .Z(n38727) );
  NANDN U47872 ( .A(n38744), .B(n38745), .Z(n38743) );
  NANDN U47873 ( .A(n38746), .B(n38747), .Z(n38745) );
  NANDN U47874 ( .A(n38747), .B(n38746), .Z(n38742) );
  XOR U47875 ( .A(n38741), .B(n38748), .Z(N61959) );
  XOR U47876 ( .A(n38738), .B(n38740), .Z(n38748) );
  XNOR U47877 ( .A(n38734), .B(n38749), .Z(n38740) );
  XNOR U47878 ( .A(n38732), .B(n38735), .Z(n38749) );
  NAND U47879 ( .A(n38750), .B(n38751), .Z(n38735) );
  NAND U47880 ( .A(n38752), .B(n38753), .Z(n38751) );
  OR U47881 ( .A(n38754), .B(n38755), .Z(n38752) );
  NANDN U47882 ( .A(n38756), .B(n38754), .Z(n38750) );
  IV U47883 ( .A(n38755), .Z(n38756) );
  NAND U47884 ( .A(n38757), .B(n38758), .Z(n38732) );
  NAND U47885 ( .A(n38759), .B(n38760), .Z(n38758) );
  NANDN U47886 ( .A(n38761), .B(n38762), .Z(n38759) );
  NANDN U47887 ( .A(n38762), .B(n38761), .Z(n38757) );
  AND U47888 ( .A(n38763), .B(n38764), .Z(n38734) );
  NAND U47889 ( .A(n38765), .B(n38766), .Z(n38764) );
  OR U47890 ( .A(n38767), .B(n38768), .Z(n38765) );
  NANDN U47891 ( .A(n38769), .B(n38767), .Z(n38763) );
  NAND U47892 ( .A(n38770), .B(n38771), .Z(n38738) );
  NANDN U47893 ( .A(n38772), .B(n38773), .Z(n38771) );
  OR U47894 ( .A(n38774), .B(n38775), .Z(n38773) );
  NANDN U47895 ( .A(n38776), .B(n38774), .Z(n38770) );
  IV U47896 ( .A(n38775), .Z(n38776) );
  XNOR U47897 ( .A(n38746), .B(n38777), .Z(n38741) );
  XNOR U47898 ( .A(n38744), .B(n38747), .Z(n38777) );
  NAND U47899 ( .A(n38778), .B(n38779), .Z(n38747) );
  NAND U47900 ( .A(n38780), .B(n38781), .Z(n38779) );
  OR U47901 ( .A(n38782), .B(n38783), .Z(n38780) );
  NANDN U47902 ( .A(n38784), .B(n38782), .Z(n38778) );
  IV U47903 ( .A(n38783), .Z(n38784) );
  NAND U47904 ( .A(n38785), .B(n38786), .Z(n38744) );
  NAND U47905 ( .A(n38787), .B(n38788), .Z(n38786) );
  NANDN U47906 ( .A(n38789), .B(n38790), .Z(n38787) );
  NANDN U47907 ( .A(n38790), .B(n38789), .Z(n38785) );
  AND U47908 ( .A(n38791), .B(n38792), .Z(n38746) );
  NAND U47909 ( .A(n38793), .B(n38794), .Z(n38792) );
  OR U47910 ( .A(n38795), .B(n38796), .Z(n38793) );
  NANDN U47911 ( .A(n38797), .B(n38795), .Z(n38791) );
  XNOR U47912 ( .A(n38772), .B(n38798), .Z(N61958) );
  XOR U47913 ( .A(n38774), .B(n38775), .Z(n38798) );
  XNOR U47914 ( .A(n38788), .B(n38799), .Z(n38775) );
  XOR U47915 ( .A(n38789), .B(n38790), .Z(n38799) );
  XOR U47916 ( .A(n38795), .B(n38800), .Z(n38790) );
  XOR U47917 ( .A(n38794), .B(n38797), .Z(n38800) );
  IV U47918 ( .A(n38796), .Z(n38797) );
  NAND U47919 ( .A(n38801), .B(n38802), .Z(n38796) );
  OR U47920 ( .A(n38803), .B(n38804), .Z(n38802) );
  OR U47921 ( .A(n38805), .B(n38806), .Z(n38801) );
  NAND U47922 ( .A(n38807), .B(n38808), .Z(n38794) );
  OR U47923 ( .A(n38809), .B(n38810), .Z(n38808) );
  OR U47924 ( .A(n38811), .B(n38812), .Z(n38807) );
  NOR U47925 ( .A(n38813), .B(n38814), .Z(n38795) );
  ANDN U47926 ( .B(n38815), .A(n38816), .Z(n38789) );
  XNOR U47927 ( .A(n38782), .B(n38817), .Z(n38788) );
  XNOR U47928 ( .A(n38781), .B(n38783), .Z(n38817) );
  NAND U47929 ( .A(n38818), .B(n38819), .Z(n38783) );
  OR U47930 ( .A(n38820), .B(n38821), .Z(n38819) );
  OR U47931 ( .A(n38822), .B(n38823), .Z(n38818) );
  NAND U47932 ( .A(n38824), .B(n38825), .Z(n38781) );
  OR U47933 ( .A(n38826), .B(n38827), .Z(n38825) );
  OR U47934 ( .A(n38828), .B(n38829), .Z(n38824) );
  ANDN U47935 ( .B(n38830), .A(n38831), .Z(n38782) );
  IV U47936 ( .A(n38832), .Z(n38830) );
  ANDN U47937 ( .B(n38833), .A(n38834), .Z(n38774) );
  XOR U47938 ( .A(n38760), .B(n38835), .Z(n38772) );
  XOR U47939 ( .A(n38761), .B(n38762), .Z(n38835) );
  XOR U47940 ( .A(n38767), .B(n38836), .Z(n38762) );
  XOR U47941 ( .A(n38766), .B(n38769), .Z(n38836) );
  IV U47942 ( .A(n38768), .Z(n38769) );
  NAND U47943 ( .A(n38837), .B(n38838), .Z(n38768) );
  OR U47944 ( .A(n38839), .B(n38840), .Z(n38838) );
  OR U47945 ( .A(n38841), .B(n38842), .Z(n38837) );
  NAND U47946 ( .A(n38843), .B(n38844), .Z(n38766) );
  OR U47947 ( .A(n38845), .B(n38846), .Z(n38844) );
  OR U47948 ( .A(n38847), .B(n38848), .Z(n38843) );
  NOR U47949 ( .A(n38849), .B(n38850), .Z(n38767) );
  ANDN U47950 ( .B(n38851), .A(n38852), .Z(n38761) );
  IV U47951 ( .A(n38853), .Z(n38851) );
  XNOR U47952 ( .A(n38754), .B(n38854), .Z(n38760) );
  XNOR U47953 ( .A(n38753), .B(n38755), .Z(n38854) );
  NAND U47954 ( .A(n38855), .B(n38856), .Z(n38755) );
  OR U47955 ( .A(n38857), .B(n38858), .Z(n38856) );
  OR U47956 ( .A(n38859), .B(n38860), .Z(n38855) );
  NAND U47957 ( .A(n38861), .B(n38862), .Z(n38753) );
  OR U47958 ( .A(n38863), .B(n38864), .Z(n38862) );
  OR U47959 ( .A(n38865), .B(n38866), .Z(n38861) );
  ANDN U47960 ( .B(n38867), .A(n38868), .Z(n38754) );
  IV U47961 ( .A(n38869), .Z(n38867) );
  XNOR U47962 ( .A(n38834), .B(n38833), .Z(N61957) );
  XOR U47963 ( .A(n38853), .B(n38852), .Z(n38833) );
  XNOR U47964 ( .A(n38868), .B(n38869), .Z(n38852) );
  XNOR U47965 ( .A(n38863), .B(n38864), .Z(n38869) );
  XNOR U47966 ( .A(n38865), .B(n38866), .Z(n38864) );
  XNOR U47967 ( .A(y[2533]), .B(x[2533]), .Z(n38866) );
  XNOR U47968 ( .A(y[2534]), .B(x[2534]), .Z(n38865) );
  XNOR U47969 ( .A(y[2532]), .B(x[2532]), .Z(n38863) );
  XNOR U47970 ( .A(n38857), .B(n38858), .Z(n38868) );
  XNOR U47971 ( .A(y[2529]), .B(x[2529]), .Z(n38858) );
  XNOR U47972 ( .A(n38859), .B(n38860), .Z(n38857) );
  XNOR U47973 ( .A(y[2530]), .B(x[2530]), .Z(n38860) );
  XNOR U47974 ( .A(y[2531]), .B(x[2531]), .Z(n38859) );
  XNOR U47975 ( .A(n38850), .B(n38849), .Z(n38853) );
  XNOR U47976 ( .A(n38845), .B(n38846), .Z(n38849) );
  XNOR U47977 ( .A(y[2526]), .B(x[2526]), .Z(n38846) );
  XNOR U47978 ( .A(n38847), .B(n38848), .Z(n38845) );
  XNOR U47979 ( .A(y[2527]), .B(x[2527]), .Z(n38848) );
  XNOR U47980 ( .A(y[2528]), .B(x[2528]), .Z(n38847) );
  XNOR U47981 ( .A(n38839), .B(n38840), .Z(n38850) );
  XNOR U47982 ( .A(y[2523]), .B(x[2523]), .Z(n38840) );
  XNOR U47983 ( .A(n38841), .B(n38842), .Z(n38839) );
  XNOR U47984 ( .A(y[2524]), .B(x[2524]), .Z(n38842) );
  XNOR U47985 ( .A(y[2525]), .B(x[2525]), .Z(n38841) );
  XOR U47986 ( .A(n38815), .B(n38816), .Z(n38834) );
  XNOR U47987 ( .A(n38831), .B(n38832), .Z(n38816) );
  XNOR U47988 ( .A(n38826), .B(n38827), .Z(n38832) );
  XNOR U47989 ( .A(n38828), .B(n38829), .Z(n38827) );
  XNOR U47990 ( .A(y[2521]), .B(x[2521]), .Z(n38829) );
  XNOR U47991 ( .A(y[2522]), .B(x[2522]), .Z(n38828) );
  XNOR U47992 ( .A(y[2520]), .B(x[2520]), .Z(n38826) );
  XNOR U47993 ( .A(n38820), .B(n38821), .Z(n38831) );
  XNOR U47994 ( .A(y[2517]), .B(x[2517]), .Z(n38821) );
  XNOR U47995 ( .A(n38822), .B(n38823), .Z(n38820) );
  XNOR U47996 ( .A(y[2518]), .B(x[2518]), .Z(n38823) );
  XNOR U47997 ( .A(y[2519]), .B(x[2519]), .Z(n38822) );
  XOR U47998 ( .A(n38814), .B(n38813), .Z(n38815) );
  XNOR U47999 ( .A(n38809), .B(n38810), .Z(n38813) );
  XNOR U48000 ( .A(y[2514]), .B(x[2514]), .Z(n38810) );
  XNOR U48001 ( .A(n38811), .B(n38812), .Z(n38809) );
  XNOR U48002 ( .A(y[2515]), .B(x[2515]), .Z(n38812) );
  XNOR U48003 ( .A(y[2516]), .B(x[2516]), .Z(n38811) );
  XNOR U48004 ( .A(n38803), .B(n38804), .Z(n38814) );
  XNOR U48005 ( .A(y[2511]), .B(x[2511]), .Z(n38804) );
  XNOR U48006 ( .A(n38805), .B(n38806), .Z(n38803) );
  XNOR U48007 ( .A(y[2512]), .B(x[2512]), .Z(n38806) );
  XNOR U48008 ( .A(y[2513]), .B(x[2513]), .Z(n38805) );
  NAND U48009 ( .A(n38870), .B(n38871), .Z(N61948) );
  NANDN U48010 ( .A(n38872), .B(n38873), .Z(n38871) );
  OR U48011 ( .A(n38874), .B(n38875), .Z(n38873) );
  NAND U48012 ( .A(n38874), .B(n38875), .Z(n38870) );
  XOR U48013 ( .A(n38874), .B(n38876), .Z(N61947) );
  XNOR U48014 ( .A(n38872), .B(n38875), .Z(n38876) );
  AND U48015 ( .A(n38877), .B(n38878), .Z(n38875) );
  NANDN U48016 ( .A(n38879), .B(n38880), .Z(n38878) );
  NANDN U48017 ( .A(n38881), .B(n38882), .Z(n38880) );
  NANDN U48018 ( .A(n38882), .B(n38881), .Z(n38877) );
  NAND U48019 ( .A(n38883), .B(n38884), .Z(n38872) );
  NANDN U48020 ( .A(n38885), .B(n38886), .Z(n38884) );
  OR U48021 ( .A(n38887), .B(n38888), .Z(n38886) );
  NAND U48022 ( .A(n38888), .B(n38887), .Z(n38883) );
  AND U48023 ( .A(n38889), .B(n38890), .Z(n38874) );
  NANDN U48024 ( .A(n38891), .B(n38892), .Z(n38890) );
  NANDN U48025 ( .A(n38893), .B(n38894), .Z(n38892) );
  NANDN U48026 ( .A(n38894), .B(n38893), .Z(n38889) );
  XOR U48027 ( .A(n38888), .B(n38895), .Z(N61946) );
  XOR U48028 ( .A(n38885), .B(n38887), .Z(n38895) );
  XNOR U48029 ( .A(n38881), .B(n38896), .Z(n38887) );
  XNOR U48030 ( .A(n38879), .B(n38882), .Z(n38896) );
  NAND U48031 ( .A(n38897), .B(n38898), .Z(n38882) );
  NAND U48032 ( .A(n38899), .B(n38900), .Z(n38898) );
  OR U48033 ( .A(n38901), .B(n38902), .Z(n38899) );
  NANDN U48034 ( .A(n38903), .B(n38901), .Z(n38897) );
  IV U48035 ( .A(n38902), .Z(n38903) );
  NAND U48036 ( .A(n38904), .B(n38905), .Z(n38879) );
  NAND U48037 ( .A(n38906), .B(n38907), .Z(n38905) );
  NANDN U48038 ( .A(n38908), .B(n38909), .Z(n38906) );
  NANDN U48039 ( .A(n38909), .B(n38908), .Z(n38904) );
  AND U48040 ( .A(n38910), .B(n38911), .Z(n38881) );
  NAND U48041 ( .A(n38912), .B(n38913), .Z(n38911) );
  OR U48042 ( .A(n38914), .B(n38915), .Z(n38912) );
  NANDN U48043 ( .A(n38916), .B(n38914), .Z(n38910) );
  NAND U48044 ( .A(n38917), .B(n38918), .Z(n38885) );
  NANDN U48045 ( .A(n38919), .B(n38920), .Z(n38918) );
  OR U48046 ( .A(n38921), .B(n38922), .Z(n38920) );
  NANDN U48047 ( .A(n38923), .B(n38921), .Z(n38917) );
  IV U48048 ( .A(n38922), .Z(n38923) );
  XNOR U48049 ( .A(n38893), .B(n38924), .Z(n38888) );
  XNOR U48050 ( .A(n38891), .B(n38894), .Z(n38924) );
  NAND U48051 ( .A(n38925), .B(n38926), .Z(n38894) );
  NAND U48052 ( .A(n38927), .B(n38928), .Z(n38926) );
  OR U48053 ( .A(n38929), .B(n38930), .Z(n38927) );
  NANDN U48054 ( .A(n38931), .B(n38929), .Z(n38925) );
  IV U48055 ( .A(n38930), .Z(n38931) );
  NAND U48056 ( .A(n38932), .B(n38933), .Z(n38891) );
  NAND U48057 ( .A(n38934), .B(n38935), .Z(n38933) );
  NANDN U48058 ( .A(n38936), .B(n38937), .Z(n38934) );
  NANDN U48059 ( .A(n38937), .B(n38936), .Z(n38932) );
  AND U48060 ( .A(n38938), .B(n38939), .Z(n38893) );
  NAND U48061 ( .A(n38940), .B(n38941), .Z(n38939) );
  OR U48062 ( .A(n38942), .B(n38943), .Z(n38940) );
  NANDN U48063 ( .A(n38944), .B(n38942), .Z(n38938) );
  XNOR U48064 ( .A(n38919), .B(n38945), .Z(N61945) );
  XOR U48065 ( .A(n38921), .B(n38922), .Z(n38945) );
  XNOR U48066 ( .A(n38935), .B(n38946), .Z(n38922) );
  XOR U48067 ( .A(n38936), .B(n38937), .Z(n38946) );
  XOR U48068 ( .A(n38942), .B(n38947), .Z(n38937) );
  XOR U48069 ( .A(n38941), .B(n38944), .Z(n38947) );
  IV U48070 ( .A(n38943), .Z(n38944) );
  NAND U48071 ( .A(n38948), .B(n38949), .Z(n38943) );
  OR U48072 ( .A(n38950), .B(n38951), .Z(n38949) );
  OR U48073 ( .A(n38952), .B(n38953), .Z(n38948) );
  NAND U48074 ( .A(n38954), .B(n38955), .Z(n38941) );
  OR U48075 ( .A(n38956), .B(n38957), .Z(n38955) );
  OR U48076 ( .A(n38958), .B(n38959), .Z(n38954) );
  NOR U48077 ( .A(n38960), .B(n38961), .Z(n38942) );
  ANDN U48078 ( .B(n38962), .A(n38963), .Z(n38936) );
  XNOR U48079 ( .A(n38929), .B(n38964), .Z(n38935) );
  XNOR U48080 ( .A(n38928), .B(n38930), .Z(n38964) );
  NAND U48081 ( .A(n38965), .B(n38966), .Z(n38930) );
  OR U48082 ( .A(n38967), .B(n38968), .Z(n38966) );
  OR U48083 ( .A(n38969), .B(n38970), .Z(n38965) );
  NAND U48084 ( .A(n38971), .B(n38972), .Z(n38928) );
  OR U48085 ( .A(n38973), .B(n38974), .Z(n38972) );
  OR U48086 ( .A(n38975), .B(n38976), .Z(n38971) );
  ANDN U48087 ( .B(n38977), .A(n38978), .Z(n38929) );
  IV U48088 ( .A(n38979), .Z(n38977) );
  ANDN U48089 ( .B(n38980), .A(n38981), .Z(n38921) );
  XOR U48090 ( .A(n38907), .B(n38982), .Z(n38919) );
  XOR U48091 ( .A(n38908), .B(n38909), .Z(n38982) );
  XOR U48092 ( .A(n38914), .B(n38983), .Z(n38909) );
  XOR U48093 ( .A(n38913), .B(n38916), .Z(n38983) );
  IV U48094 ( .A(n38915), .Z(n38916) );
  NAND U48095 ( .A(n38984), .B(n38985), .Z(n38915) );
  OR U48096 ( .A(n38986), .B(n38987), .Z(n38985) );
  OR U48097 ( .A(n38988), .B(n38989), .Z(n38984) );
  NAND U48098 ( .A(n38990), .B(n38991), .Z(n38913) );
  OR U48099 ( .A(n38992), .B(n38993), .Z(n38991) );
  OR U48100 ( .A(n38994), .B(n38995), .Z(n38990) );
  NOR U48101 ( .A(n38996), .B(n38997), .Z(n38914) );
  ANDN U48102 ( .B(n38998), .A(n38999), .Z(n38908) );
  IV U48103 ( .A(n39000), .Z(n38998) );
  XNOR U48104 ( .A(n38901), .B(n39001), .Z(n38907) );
  XNOR U48105 ( .A(n38900), .B(n38902), .Z(n39001) );
  NAND U48106 ( .A(n39002), .B(n39003), .Z(n38902) );
  OR U48107 ( .A(n39004), .B(n39005), .Z(n39003) );
  OR U48108 ( .A(n39006), .B(n39007), .Z(n39002) );
  NAND U48109 ( .A(n39008), .B(n39009), .Z(n38900) );
  OR U48110 ( .A(n39010), .B(n39011), .Z(n39009) );
  OR U48111 ( .A(n39012), .B(n39013), .Z(n39008) );
  ANDN U48112 ( .B(n39014), .A(n39015), .Z(n38901) );
  IV U48113 ( .A(n39016), .Z(n39014) );
  XNOR U48114 ( .A(n38981), .B(n38980), .Z(N61944) );
  XOR U48115 ( .A(n39000), .B(n38999), .Z(n38980) );
  XNOR U48116 ( .A(n39015), .B(n39016), .Z(n38999) );
  XNOR U48117 ( .A(n39010), .B(n39011), .Z(n39016) );
  XNOR U48118 ( .A(n39012), .B(n39013), .Z(n39011) );
  XNOR U48119 ( .A(y[2509]), .B(x[2509]), .Z(n39013) );
  XNOR U48120 ( .A(y[2510]), .B(x[2510]), .Z(n39012) );
  XNOR U48121 ( .A(y[2508]), .B(x[2508]), .Z(n39010) );
  XNOR U48122 ( .A(n39004), .B(n39005), .Z(n39015) );
  XNOR U48123 ( .A(y[2505]), .B(x[2505]), .Z(n39005) );
  XNOR U48124 ( .A(n39006), .B(n39007), .Z(n39004) );
  XNOR U48125 ( .A(y[2506]), .B(x[2506]), .Z(n39007) );
  XNOR U48126 ( .A(y[2507]), .B(x[2507]), .Z(n39006) );
  XNOR U48127 ( .A(n38997), .B(n38996), .Z(n39000) );
  XNOR U48128 ( .A(n38992), .B(n38993), .Z(n38996) );
  XNOR U48129 ( .A(y[2502]), .B(x[2502]), .Z(n38993) );
  XNOR U48130 ( .A(n38994), .B(n38995), .Z(n38992) );
  XNOR U48131 ( .A(y[2503]), .B(x[2503]), .Z(n38995) );
  XNOR U48132 ( .A(y[2504]), .B(x[2504]), .Z(n38994) );
  XNOR U48133 ( .A(n38986), .B(n38987), .Z(n38997) );
  XNOR U48134 ( .A(y[2499]), .B(x[2499]), .Z(n38987) );
  XNOR U48135 ( .A(n38988), .B(n38989), .Z(n38986) );
  XNOR U48136 ( .A(y[2500]), .B(x[2500]), .Z(n38989) );
  XNOR U48137 ( .A(y[2501]), .B(x[2501]), .Z(n38988) );
  XOR U48138 ( .A(n38962), .B(n38963), .Z(n38981) );
  XNOR U48139 ( .A(n38978), .B(n38979), .Z(n38963) );
  XNOR U48140 ( .A(n38973), .B(n38974), .Z(n38979) );
  XNOR U48141 ( .A(n38975), .B(n38976), .Z(n38974) );
  XNOR U48142 ( .A(y[2497]), .B(x[2497]), .Z(n38976) );
  XNOR U48143 ( .A(y[2498]), .B(x[2498]), .Z(n38975) );
  XNOR U48144 ( .A(y[2496]), .B(x[2496]), .Z(n38973) );
  XNOR U48145 ( .A(n38967), .B(n38968), .Z(n38978) );
  XNOR U48146 ( .A(y[2493]), .B(x[2493]), .Z(n38968) );
  XNOR U48147 ( .A(n38969), .B(n38970), .Z(n38967) );
  XNOR U48148 ( .A(y[2494]), .B(x[2494]), .Z(n38970) );
  XNOR U48149 ( .A(y[2495]), .B(x[2495]), .Z(n38969) );
  XOR U48150 ( .A(n38961), .B(n38960), .Z(n38962) );
  XNOR U48151 ( .A(n38956), .B(n38957), .Z(n38960) );
  XNOR U48152 ( .A(y[2490]), .B(x[2490]), .Z(n38957) );
  XNOR U48153 ( .A(n38958), .B(n38959), .Z(n38956) );
  XNOR U48154 ( .A(y[2491]), .B(x[2491]), .Z(n38959) );
  XNOR U48155 ( .A(y[2492]), .B(x[2492]), .Z(n38958) );
  XNOR U48156 ( .A(n38950), .B(n38951), .Z(n38961) );
  XNOR U48157 ( .A(y[2487]), .B(x[2487]), .Z(n38951) );
  XNOR U48158 ( .A(n38952), .B(n38953), .Z(n38950) );
  XNOR U48159 ( .A(y[2488]), .B(x[2488]), .Z(n38953) );
  XNOR U48160 ( .A(y[2489]), .B(x[2489]), .Z(n38952) );
  NAND U48161 ( .A(n39017), .B(n39018), .Z(N61935) );
  NANDN U48162 ( .A(n39019), .B(n39020), .Z(n39018) );
  OR U48163 ( .A(n39021), .B(n39022), .Z(n39020) );
  NAND U48164 ( .A(n39021), .B(n39022), .Z(n39017) );
  XOR U48165 ( .A(n39021), .B(n39023), .Z(N61934) );
  XNOR U48166 ( .A(n39019), .B(n39022), .Z(n39023) );
  AND U48167 ( .A(n39024), .B(n39025), .Z(n39022) );
  NANDN U48168 ( .A(n39026), .B(n39027), .Z(n39025) );
  NANDN U48169 ( .A(n39028), .B(n39029), .Z(n39027) );
  NANDN U48170 ( .A(n39029), .B(n39028), .Z(n39024) );
  NAND U48171 ( .A(n39030), .B(n39031), .Z(n39019) );
  NANDN U48172 ( .A(n39032), .B(n39033), .Z(n39031) );
  OR U48173 ( .A(n39034), .B(n39035), .Z(n39033) );
  NAND U48174 ( .A(n39035), .B(n39034), .Z(n39030) );
  AND U48175 ( .A(n39036), .B(n39037), .Z(n39021) );
  NANDN U48176 ( .A(n39038), .B(n39039), .Z(n39037) );
  NANDN U48177 ( .A(n39040), .B(n39041), .Z(n39039) );
  NANDN U48178 ( .A(n39041), .B(n39040), .Z(n39036) );
  XOR U48179 ( .A(n39035), .B(n39042), .Z(N61933) );
  XOR U48180 ( .A(n39032), .B(n39034), .Z(n39042) );
  XNOR U48181 ( .A(n39028), .B(n39043), .Z(n39034) );
  XNOR U48182 ( .A(n39026), .B(n39029), .Z(n39043) );
  NAND U48183 ( .A(n39044), .B(n39045), .Z(n39029) );
  NAND U48184 ( .A(n39046), .B(n39047), .Z(n39045) );
  OR U48185 ( .A(n39048), .B(n39049), .Z(n39046) );
  NANDN U48186 ( .A(n39050), .B(n39048), .Z(n39044) );
  IV U48187 ( .A(n39049), .Z(n39050) );
  NAND U48188 ( .A(n39051), .B(n39052), .Z(n39026) );
  NAND U48189 ( .A(n39053), .B(n39054), .Z(n39052) );
  NANDN U48190 ( .A(n39055), .B(n39056), .Z(n39053) );
  NANDN U48191 ( .A(n39056), .B(n39055), .Z(n39051) );
  AND U48192 ( .A(n39057), .B(n39058), .Z(n39028) );
  NAND U48193 ( .A(n39059), .B(n39060), .Z(n39058) );
  OR U48194 ( .A(n39061), .B(n39062), .Z(n39059) );
  NANDN U48195 ( .A(n39063), .B(n39061), .Z(n39057) );
  NAND U48196 ( .A(n39064), .B(n39065), .Z(n39032) );
  NANDN U48197 ( .A(n39066), .B(n39067), .Z(n39065) );
  OR U48198 ( .A(n39068), .B(n39069), .Z(n39067) );
  NANDN U48199 ( .A(n39070), .B(n39068), .Z(n39064) );
  IV U48200 ( .A(n39069), .Z(n39070) );
  XNOR U48201 ( .A(n39040), .B(n39071), .Z(n39035) );
  XNOR U48202 ( .A(n39038), .B(n39041), .Z(n39071) );
  NAND U48203 ( .A(n39072), .B(n39073), .Z(n39041) );
  NAND U48204 ( .A(n39074), .B(n39075), .Z(n39073) );
  OR U48205 ( .A(n39076), .B(n39077), .Z(n39074) );
  NANDN U48206 ( .A(n39078), .B(n39076), .Z(n39072) );
  IV U48207 ( .A(n39077), .Z(n39078) );
  NAND U48208 ( .A(n39079), .B(n39080), .Z(n39038) );
  NAND U48209 ( .A(n39081), .B(n39082), .Z(n39080) );
  NANDN U48210 ( .A(n39083), .B(n39084), .Z(n39081) );
  NANDN U48211 ( .A(n39084), .B(n39083), .Z(n39079) );
  AND U48212 ( .A(n39085), .B(n39086), .Z(n39040) );
  NAND U48213 ( .A(n39087), .B(n39088), .Z(n39086) );
  OR U48214 ( .A(n39089), .B(n39090), .Z(n39087) );
  NANDN U48215 ( .A(n39091), .B(n39089), .Z(n39085) );
  XNOR U48216 ( .A(n39066), .B(n39092), .Z(N61932) );
  XOR U48217 ( .A(n39068), .B(n39069), .Z(n39092) );
  XNOR U48218 ( .A(n39082), .B(n39093), .Z(n39069) );
  XOR U48219 ( .A(n39083), .B(n39084), .Z(n39093) );
  XOR U48220 ( .A(n39089), .B(n39094), .Z(n39084) );
  XOR U48221 ( .A(n39088), .B(n39091), .Z(n39094) );
  IV U48222 ( .A(n39090), .Z(n39091) );
  NAND U48223 ( .A(n39095), .B(n39096), .Z(n39090) );
  OR U48224 ( .A(n39097), .B(n39098), .Z(n39096) );
  OR U48225 ( .A(n39099), .B(n39100), .Z(n39095) );
  NAND U48226 ( .A(n39101), .B(n39102), .Z(n39088) );
  OR U48227 ( .A(n39103), .B(n39104), .Z(n39102) );
  OR U48228 ( .A(n39105), .B(n39106), .Z(n39101) );
  NOR U48229 ( .A(n39107), .B(n39108), .Z(n39089) );
  ANDN U48230 ( .B(n39109), .A(n39110), .Z(n39083) );
  XNOR U48231 ( .A(n39076), .B(n39111), .Z(n39082) );
  XNOR U48232 ( .A(n39075), .B(n39077), .Z(n39111) );
  NAND U48233 ( .A(n39112), .B(n39113), .Z(n39077) );
  OR U48234 ( .A(n39114), .B(n39115), .Z(n39113) );
  OR U48235 ( .A(n39116), .B(n39117), .Z(n39112) );
  NAND U48236 ( .A(n39118), .B(n39119), .Z(n39075) );
  OR U48237 ( .A(n39120), .B(n39121), .Z(n39119) );
  OR U48238 ( .A(n39122), .B(n39123), .Z(n39118) );
  ANDN U48239 ( .B(n39124), .A(n39125), .Z(n39076) );
  IV U48240 ( .A(n39126), .Z(n39124) );
  ANDN U48241 ( .B(n39127), .A(n39128), .Z(n39068) );
  XOR U48242 ( .A(n39054), .B(n39129), .Z(n39066) );
  XOR U48243 ( .A(n39055), .B(n39056), .Z(n39129) );
  XOR U48244 ( .A(n39061), .B(n39130), .Z(n39056) );
  XOR U48245 ( .A(n39060), .B(n39063), .Z(n39130) );
  IV U48246 ( .A(n39062), .Z(n39063) );
  NAND U48247 ( .A(n39131), .B(n39132), .Z(n39062) );
  OR U48248 ( .A(n39133), .B(n39134), .Z(n39132) );
  OR U48249 ( .A(n39135), .B(n39136), .Z(n39131) );
  NAND U48250 ( .A(n39137), .B(n39138), .Z(n39060) );
  OR U48251 ( .A(n39139), .B(n39140), .Z(n39138) );
  OR U48252 ( .A(n39141), .B(n39142), .Z(n39137) );
  NOR U48253 ( .A(n39143), .B(n39144), .Z(n39061) );
  ANDN U48254 ( .B(n39145), .A(n39146), .Z(n39055) );
  IV U48255 ( .A(n39147), .Z(n39145) );
  XNOR U48256 ( .A(n39048), .B(n39148), .Z(n39054) );
  XNOR U48257 ( .A(n39047), .B(n39049), .Z(n39148) );
  NAND U48258 ( .A(n39149), .B(n39150), .Z(n39049) );
  OR U48259 ( .A(n39151), .B(n39152), .Z(n39150) );
  OR U48260 ( .A(n39153), .B(n39154), .Z(n39149) );
  NAND U48261 ( .A(n39155), .B(n39156), .Z(n39047) );
  OR U48262 ( .A(n39157), .B(n39158), .Z(n39156) );
  OR U48263 ( .A(n39159), .B(n39160), .Z(n39155) );
  ANDN U48264 ( .B(n39161), .A(n39162), .Z(n39048) );
  IV U48265 ( .A(n39163), .Z(n39161) );
  XNOR U48266 ( .A(n39128), .B(n39127), .Z(N61931) );
  XOR U48267 ( .A(n39147), .B(n39146), .Z(n39127) );
  XNOR U48268 ( .A(n39162), .B(n39163), .Z(n39146) );
  XNOR U48269 ( .A(n39157), .B(n39158), .Z(n39163) );
  XNOR U48270 ( .A(n39159), .B(n39160), .Z(n39158) );
  XNOR U48271 ( .A(y[2485]), .B(x[2485]), .Z(n39160) );
  XNOR U48272 ( .A(y[2486]), .B(x[2486]), .Z(n39159) );
  XNOR U48273 ( .A(y[2484]), .B(x[2484]), .Z(n39157) );
  XNOR U48274 ( .A(n39151), .B(n39152), .Z(n39162) );
  XNOR U48275 ( .A(y[2481]), .B(x[2481]), .Z(n39152) );
  XNOR U48276 ( .A(n39153), .B(n39154), .Z(n39151) );
  XNOR U48277 ( .A(y[2482]), .B(x[2482]), .Z(n39154) );
  XNOR U48278 ( .A(y[2483]), .B(x[2483]), .Z(n39153) );
  XNOR U48279 ( .A(n39144), .B(n39143), .Z(n39147) );
  XNOR U48280 ( .A(n39139), .B(n39140), .Z(n39143) );
  XNOR U48281 ( .A(y[2478]), .B(x[2478]), .Z(n39140) );
  XNOR U48282 ( .A(n39141), .B(n39142), .Z(n39139) );
  XNOR U48283 ( .A(y[2479]), .B(x[2479]), .Z(n39142) );
  XNOR U48284 ( .A(y[2480]), .B(x[2480]), .Z(n39141) );
  XNOR U48285 ( .A(n39133), .B(n39134), .Z(n39144) );
  XNOR U48286 ( .A(y[2475]), .B(x[2475]), .Z(n39134) );
  XNOR U48287 ( .A(n39135), .B(n39136), .Z(n39133) );
  XNOR U48288 ( .A(y[2476]), .B(x[2476]), .Z(n39136) );
  XNOR U48289 ( .A(y[2477]), .B(x[2477]), .Z(n39135) );
  XOR U48290 ( .A(n39109), .B(n39110), .Z(n39128) );
  XNOR U48291 ( .A(n39125), .B(n39126), .Z(n39110) );
  XNOR U48292 ( .A(n39120), .B(n39121), .Z(n39126) );
  XNOR U48293 ( .A(n39122), .B(n39123), .Z(n39121) );
  XNOR U48294 ( .A(y[2473]), .B(x[2473]), .Z(n39123) );
  XNOR U48295 ( .A(y[2474]), .B(x[2474]), .Z(n39122) );
  XNOR U48296 ( .A(y[2472]), .B(x[2472]), .Z(n39120) );
  XNOR U48297 ( .A(n39114), .B(n39115), .Z(n39125) );
  XNOR U48298 ( .A(y[2469]), .B(x[2469]), .Z(n39115) );
  XNOR U48299 ( .A(n39116), .B(n39117), .Z(n39114) );
  XNOR U48300 ( .A(y[2470]), .B(x[2470]), .Z(n39117) );
  XNOR U48301 ( .A(y[2471]), .B(x[2471]), .Z(n39116) );
  XOR U48302 ( .A(n39108), .B(n39107), .Z(n39109) );
  XNOR U48303 ( .A(n39103), .B(n39104), .Z(n39107) );
  XNOR U48304 ( .A(y[2466]), .B(x[2466]), .Z(n39104) );
  XNOR U48305 ( .A(n39105), .B(n39106), .Z(n39103) );
  XNOR U48306 ( .A(y[2467]), .B(x[2467]), .Z(n39106) );
  XNOR U48307 ( .A(y[2468]), .B(x[2468]), .Z(n39105) );
  XNOR U48308 ( .A(n39097), .B(n39098), .Z(n39108) );
  XNOR U48309 ( .A(y[2463]), .B(x[2463]), .Z(n39098) );
  XNOR U48310 ( .A(n39099), .B(n39100), .Z(n39097) );
  XNOR U48311 ( .A(y[2464]), .B(x[2464]), .Z(n39100) );
  XNOR U48312 ( .A(y[2465]), .B(x[2465]), .Z(n39099) );
  NAND U48313 ( .A(n39164), .B(n39165), .Z(N61922) );
  NANDN U48314 ( .A(n39166), .B(n39167), .Z(n39165) );
  OR U48315 ( .A(n39168), .B(n39169), .Z(n39167) );
  NAND U48316 ( .A(n39168), .B(n39169), .Z(n39164) );
  XOR U48317 ( .A(n39168), .B(n39170), .Z(N61921) );
  XNOR U48318 ( .A(n39166), .B(n39169), .Z(n39170) );
  AND U48319 ( .A(n39171), .B(n39172), .Z(n39169) );
  NANDN U48320 ( .A(n39173), .B(n39174), .Z(n39172) );
  NANDN U48321 ( .A(n39175), .B(n39176), .Z(n39174) );
  NANDN U48322 ( .A(n39176), .B(n39175), .Z(n39171) );
  NAND U48323 ( .A(n39177), .B(n39178), .Z(n39166) );
  NANDN U48324 ( .A(n39179), .B(n39180), .Z(n39178) );
  OR U48325 ( .A(n39181), .B(n39182), .Z(n39180) );
  NAND U48326 ( .A(n39182), .B(n39181), .Z(n39177) );
  AND U48327 ( .A(n39183), .B(n39184), .Z(n39168) );
  NANDN U48328 ( .A(n39185), .B(n39186), .Z(n39184) );
  NANDN U48329 ( .A(n39187), .B(n39188), .Z(n39186) );
  NANDN U48330 ( .A(n39188), .B(n39187), .Z(n39183) );
  XOR U48331 ( .A(n39182), .B(n39189), .Z(N61920) );
  XOR U48332 ( .A(n39179), .B(n39181), .Z(n39189) );
  XNOR U48333 ( .A(n39175), .B(n39190), .Z(n39181) );
  XNOR U48334 ( .A(n39173), .B(n39176), .Z(n39190) );
  NAND U48335 ( .A(n39191), .B(n39192), .Z(n39176) );
  NAND U48336 ( .A(n39193), .B(n39194), .Z(n39192) );
  OR U48337 ( .A(n39195), .B(n39196), .Z(n39193) );
  NANDN U48338 ( .A(n39197), .B(n39195), .Z(n39191) );
  IV U48339 ( .A(n39196), .Z(n39197) );
  NAND U48340 ( .A(n39198), .B(n39199), .Z(n39173) );
  NAND U48341 ( .A(n39200), .B(n39201), .Z(n39199) );
  NANDN U48342 ( .A(n39202), .B(n39203), .Z(n39200) );
  NANDN U48343 ( .A(n39203), .B(n39202), .Z(n39198) );
  AND U48344 ( .A(n39204), .B(n39205), .Z(n39175) );
  NAND U48345 ( .A(n39206), .B(n39207), .Z(n39205) );
  OR U48346 ( .A(n39208), .B(n39209), .Z(n39206) );
  NANDN U48347 ( .A(n39210), .B(n39208), .Z(n39204) );
  NAND U48348 ( .A(n39211), .B(n39212), .Z(n39179) );
  NANDN U48349 ( .A(n39213), .B(n39214), .Z(n39212) );
  OR U48350 ( .A(n39215), .B(n39216), .Z(n39214) );
  NANDN U48351 ( .A(n39217), .B(n39215), .Z(n39211) );
  IV U48352 ( .A(n39216), .Z(n39217) );
  XNOR U48353 ( .A(n39187), .B(n39218), .Z(n39182) );
  XNOR U48354 ( .A(n39185), .B(n39188), .Z(n39218) );
  NAND U48355 ( .A(n39219), .B(n39220), .Z(n39188) );
  NAND U48356 ( .A(n39221), .B(n39222), .Z(n39220) );
  OR U48357 ( .A(n39223), .B(n39224), .Z(n39221) );
  NANDN U48358 ( .A(n39225), .B(n39223), .Z(n39219) );
  IV U48359 ( .A(n39224), .Z(n39225) );
  NAND U48360 ( .A(n39226), .B(n39227), .Z(n39185) );
  NAND U48361 ( .A(n39228), .B(n39229), .Z(n39227) );
  NANDN U48362 ( .A(n39230), .B(n39231), .Z(n39228) );
  NANDN U48363 ( .A(n39231), .B(n39230), .Z(n39226) );
  AND U48364 ( .A(n39232), .B(n39233), .Z(n39187) );
  NAND U48365 ( .A(n39234), .B(n39235), .Z(n39233) );
  OR U48366 ( .A(n39236), .B(n39237), .Z(n39234) );
  NANDN U48367 ( .A(n39238), .B(n39236), .Z(n39232) );
  XNOR U48368 ( .A(n39213), .B(n39239), .Z(N61919) );
  XOR U48369 ( .A(n39215), .B(n39216), .Z(n39239) );
  XNOR U48370 ( .A(n39229), .B(n39240), .Z(n39216) );
  XOR U48371 ( .A(n39230), .B(n39231), .Z(n39240) );
  XOR U48372 ( .A(n39236), .B(n39241), .Z(n39231) );
  XOR U48373 ( .A(n39235), .B(n39238), .Z(n39241) );
  IV U48374 ( .A(n39237), .Z(n39238) );
  NAND U48375 ( .A(n39242), .B(n39243), .Z(n39237) );
  OR U48376 ( .A(n39244), .B(n39245), .Z(n39243) );
  OR U48377 ( .A(n39246), .B(n39247), .Z(n39242) );
  NAND U48378 ( .A(n39248), .B(n39249), .Z(n39235) );
  OR U48379 ( .A(n39250), .B(n39251), .Z(n39249) );
  OR U48380 ( .A(n39252), .B(n39253), .Z(n39248) );
  NOR U48381 ( .A(n39254), .B(n39255), .Z(n39236) );
  ANDN U48382 ( .B(n39256), .A(n39257), .Z(n39230) );
  XNOR U48383 ( .A(n39223), .B(n39258), .Z(n39229) );
  XNOR U48384 ( .A(n39222), .B(n39224), .Z(n39258) );
  NAND U48385 ( .A(n39259), .B(n39260), .Z(n39224) );
  OR U48386 ( .A(n39261), .B(n39262), .Z(n39260) );
  OR U48387 ( .A(n39263), .B(n39264), .Z(n39259) );
  NAND U48388 ( .A(n39265), .B(n39266), .Z(n39222) );
  OR U48389 ( .A(n39267), .B(n39268), .Z(n39266) );
  OR U48390 ( .A(n39269), .B(n39270), .Z(n39265) );
  ANDN U48391 ( .B(n39271), .A(n39272), .Z(n39223) );
  IV U48392 ( .A(n39273), .Z(n39271) );
  ANDN U48393 ( .B(n39274), .A(n39275), .Z(n39215) );
  XOR U48394 ( .A(n39201), .B(n39276), .Z(n39213) );
  XOR U48395 ( .A(n39202), .B(n39203), .Z(n39276) );
  XOR U48396 ( .A(n39208), .B(n39277), .Z(n39203) );
  XOR U48397 ( .A(n39207), .B(n39210), .Z(n39277) );
  IV U48398 ( .A(n39209), .Z(n39210) );
  NAND U48399 ( .A(n39278), .B(n39279), .Z(n39209) );
  OR U48400 ( .A(n39280), .B(n39281), .Z(n39279) );
  OR U48401 ( .A(n39282), .B(n39283), .Z(n39278) );
  NAND U48402 ( .A(n39284), .B(n39285), .Z(n39207) );
  OR U48403 ( .A(n39286), .B(n39287), .Z(n39285) );
  OR U48404 ( .A(n39288), .B(n39289), .Z(n39284) );
  NOR U48405 ( .A(n39290), .B(n39291), .Z(n39208) );
  ANDN U48406 ( .B(n39292), .A(n39293), .Z(n39202) );
  IV U48407 ( .A(n39294), .Z(n39292) );
  XNOR U48408 ( .A(n39195), .B(n39295), .Z(n39201) );
  XNOR U48409 ( .A(n39194), .B(n39196), .Z(n39295) );
  NAND U48410 ( .A(n39296), .B(n39297), .Z(n39196) );
  OR U48411 ( .A(n39298), .B(n39299), .Z(n39297) );
  OR U48412 ( .A(n39300), .B(n39301), .Z(n39296) );
  NAND U48413 ( .A(n39302), .B(n39303), .Z(n39194) );
  OR U48414 ( .A(n39304), .B(n39305), .Z(n39303) );
  OR U48415 ( .A(n39306), .B(n39307), .Z(n39302) );
  ANDN U48416 ( .B(n39308), .A(n39309), .Z(n39195) );
  IV U48417 ( .A(n39310), .Z(n39308) );
  XNOR U48418 ( .A(n39275), .B(n39274), .Z(N61918) );
  XOR U48419 ( .A(n39294), .B(n39293), .Z(n39274) );
  XNOR U48420 ( .A(n39309), .B(n39310), .Z(n39293) );
  XNOR U48421 ( .A(n39304), .B(n39305), .Z(n39310) );
  XNOR U48422 ( .A(n39306), .B(n39307), .Z(n39305) );
  XNOR U48423 ( .A(y[2461]), .B(x[2461]), .Z(n39307) );
  XNOR U48424 ( .A(y[2462]), .B(x[2462]), .Z(n39306) );
  XNOR U48425 ( .A(y[2460]), .B(x[2460]), .Z(n39304) );
  XNOR U48426 ( .A(n39298), .B(n39299), .Z(n39309) );
  XNOR U48427 ( .A(y[2457]), .B(x[2457]), .Z(n39299) );
  XNOR U48428 ( .A(n39300), .B(n39301), .Z(n39298) );
  XNOR U48429 ( .A(y[2458]), .B(x[2458]), .Z(n39301) );
  XNOR U48430 ( .A(y[2459]), .B(x[2459]), .Z(n39300) );
  XNOR U48431 ( .A(n39291), .B(n39290), .Z(n39294) );
  XNOR U48432 ( .A(n39286), .B(n39287), .Z(n39290) );
  XNOR U48433 ( .A(y[2454]), .B(x[2454]), .Z(n39287) );
  XNOR U48434 ( .A(n39288), .B(n39289), .Z(n39286) );
  XNOR U48435 ( .A(y[2455]), .B(x[2455]), .Z(n39289) );
  XNOR U48436 ( .A(y[2456]), .B(x[2456]), .Z(n39288) );
  XNOR U48437 ( .A(n39280), .B(n39281), .Z(n39291) );
  XNOR U48438 ( .A(y[2451]), .B(x[2451]), .Z(n39281) );
  XNOR U48439 ( .A(n39282), .B(n39283), .Z(n39280) );
  XNOR U48440 ( .A(y[2452]), .B(x[2452]), .Z(n39283) );
  XNOR U48441 ( .A(y[2453]), .B(x[2453]), .Z(n39282) );
  XOR U48442 ( .A(n39256), .B(n39257), .Z(n39275) );
  XNOR U48443 ( .A(n39272), .B(n39273), .Z(n39257) );
  XNOR U48444 ( .A(n39267), .B(n39268), .Z(n39273) );
  XNOR U48445 ( .A(n39269), .B(n39270), .Z(n39268) );
  XNOR U48446 ( .A(y[2449]), .B(x[2449]), .Z(n39270) );
  XNOR U48447 ( .A(y[2450]), .B(x[2450]), .Z(n39269) );
  XNOR U48448 ( .A(y[2448]), .B(x[2448]), .Z(n39267) );
  XNOR U48449 ( .A(n39261), .B(n39262), .Z(n39272) );
  XNOR U48450 ( .A(y[2445]), .B(x[2445]), .Z(n39262) );
  XNOR U48451 ( .A(n39263), .B(n39264), .Z(n39261) );
  XNOR U48452 ( .A(y[2446]), .B(x[2446]), .Z(n39264) );
  XNOR U48453 ( .A(y[2447]), .B(x[2447]), .Z(n39263) );
  XOR U48454 ( .A(n39255), .B(n39254), .Z(n39256) );
  XNOR U48455 ( .A(n39250), .B(n39251), .Z(n39254) );
  XNOR U48456 ( .A(y[2442]), .B(x[2442]), .Z(n39251) );
  XNOR U48457 ( .A(n39252), .B(n39253), .Z(n39250) );
  XNOR U48458 ( .A(y[2443]), .B(x[2443]), .Z(n39253) );
  XNOR U48459 ( .A(y[2444]), .B(x[2444]), .Z(n39252) );
  XNOR U48460 ( .A(n39244), .B(n39245), .Z(n39255) );
  XNOR U48461 ( .A(y[2439]), .B(x[2439]), .Z(n39245) );
  XNOR U48462 ( .A(n39246), .B(n39247), .Z(n39244) );
  XNOR U48463 ( .A(y[2440]), .B(x[2440]), .Z(n39247) );
  XNOR U48464 ( .A(y[2441]), .B(x[2441]), .Z(n39246) );
  NAND U48465 ( .A(n39311), .B(n39312), .Z(N61909) );
  NANDN U48466 ( .A(n39313), .B(n39314), .Z(n39312) );
  OR U48467 ( .A(n39315), .B(n39316), .Z(n39314) );
  NAND U48468 ( .A(n39315), .B(n39316), .Z(n39311) );
  XOR U48469 ( .A(n39315), .B(n39317), .Z(N61908) );
  XNOR U48470 ( .A(n39313), .B(n39316), .Z(n39317) );
  AND U48471 ( .A(n39318), .B(n39319), .Z(n39316) );
  NANDN U48472 ( .A(n39320), .B(n39321), .Z(n39319) );
  NANDN U48473 ( .A(n39322), .B(n39323), .Z(n39321) );
  NANDN U48474 ( .A(n39323), .B(n39322), .Z(n39318) );
  NAND U48475 ( .A(n39324), .B(n39325), .Z(n39313) );
  NANDN U48476 ( .A(n39326), .B(n39327), .Z(n39325) );
  OR U48477 ( .A(n39328), .B(n39329), .Z(n39327) );
  NAND U48478 ( .A(n39329), .B(n39328), .Z(n39324) );
  AND U48479 ( .A(n39330), .B(n39331), .Z(n39315) );
  NANDN U48480 ( .A(n39332), .B(n39333), .Z(n39331) );
  NANDN U48481 ( .A(n39334), .B(n39335), .Z(n39333) );
  NANDN U48482 ( .A(n39335), .B(n39334), .Z(n39330) );
  XOR U48483 ( .A(n39329), .B(n39336), .Z(N61907) );
  XOR U48484 ( .A(n39326), .B(n39328), .Z(n39336) );
  XNOR U48485 ( .A(n39322), .B(n39337), .Z(n39328) );
  XNOR U48486 ( .A(n39320), .B(n39323), .Z(n39337) );
  NAND U48487 ( .A(n39338), .B(n39339), .Z(n39323) );
  NAND U48488 ( .A(n39340), .B(n39341), .Z(n39339) );
  OR U48489 ( .A(n39342), .B(n39343), .Z(n39340) );
  NANDN U48490 ( .A(n39344), .B(n39342), .Z(n39338) );
  IV U48491 ( .A(n39343), .Z(n39344) );
  NAND U48492 ( .A(n39345), .B(n39346), .Z(n39320) );
  NAND U48493 ( .A(n39347), .B(n39348), .Z(n39346) );
  NANDN U48494 ( .A(n39349), .B(n39350), .Z(n39347) );
  NANDN U48495 ( .A(n39350), .B(n39349), .Z(n39345) );
  AND U48496 ( .A(n39351), .B(n39352), .Z(n39322) );
  NAND U48497 ( .A(n39353), .B(n39354), .Z(n39352) );
  OR U48498 ( .A(n39355), .B(n39356), .Z(n39353) );
  NANDN U48499 ( .A(n39357), .B(n39355), .Z(n39351) );
  NAND U48500 ( .A(n39358), .B(n39359), .Z(n39326) );
  NANDN U48501 ( .A(n39360), .B(n39361), .Z(n39359) );
  OR U48502 ( .A(n39362), .B(n39363), .Z(n39361) );
  NANDN U48503 ( .A(n39364), .B(n39362), .Z(n39358) );
  IV U48504 ( .A(n39363), .Z(n39364) );
  XNOR U48505 ( .A(n39334), .B(n39365), .Z(n39329) );
  XNOR U48506 ( .A(n39332), .B(n39335), .Z(n39365) );
  NAND U48507 ( .A(n39366), .B(n39367), .Z(n39335) );
  NAND U48508 ( .A(n39368), .B(n39369), .Z(n39367) );
  OR U48509 ( .A(n39370), .B(n39371), .Z(n39368) );
  NANDN U48510 ( .A(n39372), .B(n39370), .Z(n39366) );
  IV U48511 ( .A(n39371), .Z(n39372) );
  NAND U48512 ( .A(n39373), .B(n39374), .Z(n39332) );
  NAND U48513 ( .A(n39375), .B(n39376), .Z(n39374) );
  NANDN U48514 ( .A(n39377), .B(n39378), .Z(n39375) );
  NANDN U48515 ( .A(n39378), .B(n39377), .Z(n39373) );
  AND U48516 ( .A(n39379), .B(n39380), .Z(n39334) );
  NAND U48517 ( .A(n39381), .B(n39382), .Z(n39380) );
  OR U48518 ( .A(n39383), .B(n39384), .Z(n39381) );
  NANDN U48519 ( .A(n39385), .B(n39383), .Z(n39379) );
  XNOR U48520 ( .A(n39360), .B(n39386), .Z(N61906) );
  XOR U48521 ( .A(n39362), .B(n39363), .Z(n39386) );
  XNOR U48522 ( .A(n39376), .B(n39387), .Z(n39363) );
  XOR U48523 ( .A(n39377), .B(n39378), .Z(n39387) );
  XOR U48524 ( .A(n39383), .B(n39388), .Z(n39378) );
  XOR U48525 ( .A(n39382), .B(n39385), .Z(n39388) );
  IV U48526 ( .A(n39384), .Z(n39385) );
  NAND U48527 ( .A(n39389), .B(n39390), .Z(n39384) );
  OR U48528 ( .A(n39391), .B(n39392), .Z(n39390) );
  OR U48529 ( .A(n39393), .B(n39394), .Z(n39389) );
  NAND U48530 ( .A(n39395), .B(n39396), .Z(n39382) );
  OR U48531 ( .A(n39397), .B(n39398), .Z(n39396) );
  OR U48532 ( .A(n39399), .B(n39400), .Z(n39395) );
  NOR U48533 ( .A(n39401), .B(n39402), .Z(n39383) );
  ANDN U48534 ( .B(n39403), .A(n39404), .Z(n39377) );
  XNOR U48535 ( .A(n39370), .B(n39405), .Z(n39376) );
  XNOR U48536 ( .A(n39369), .B(n39371), .Z(n39405) );
  NAND U48537 ( .A(n39406), .B(n39407), .Z(n39371) );
  OR U48538 ( .A(n39408), .B(n39409), .Z(n39407) );
  OR U48539 ( .A(n39410), .B(n39411), .Z(n39406) );
  NAND U48540 ( .A(n39412), .B(n39413), .Z(n39369) );
  OR U48541 ( .A(n39414), .B(n39415), .Z(n39413) );
  OR U48542 ( .A(n39416), .B(n39417), .Z(n39412) );
  ANDN U48543 ( .B(n39418), .A(n39419), .Z(n39370) );
  IV U48544 ( .A(n39420), .Z(n39418) );
  ANDN U48545 ( .B(n39421), .A(n39422), .Z(n39362) );
  XOR U48546 ( .A(n39348), .B(n39423), .Z(n39360) );
  XOR U48547 ( .A(n39349), .B(n39350), .Z(n39423) );
  XOR U48548 ( .A(n39355), .B(n39424), .Z(n39350) );
  XOR U48549 ( .A(n39354), .B(n39357), .Z(n39424) );
  IV U48550 ( .A(n39356), .Z(n39357) );
  NAND U48551 ( .A(n39425), .B(n39426), .Z(n39356) );
  OR U48552 ( .A(n39427), .B(n39428), .Z(n39426) );
  OR U48553 ( .A(n39429), .B(n39430), .Z(n39425) );
  NAND U48554 ( .A(n39431), .B(n39432), .Z(n39354) );
  OR U48555 ( .A(n39433), .B(n39434), .Z(n39432) );
  OR U48556 ( .A(n39435), .B(n39436), .Z(n39431) );
  NOR U48557 ( .A(n39437), .B(n39438), .Z(n39355) );
  ANDN U48558 ( .B(n39439), .A(n39440), .Z(n39349) );
  IV U48559 ( .A(n39441), .Z(n39439) );
  XNOR U48560 ( .A(n39342), .B(n39442), .Z(n39348) );
  XNOR U48561 ( .A(n39341), .B(n39343), .Z(n39442) );
  NAND U48562 ( .A(n39443), .B(n39444), .Z(n39343) );
  OR U48563 ( .A(n39445), .B(n39446), .Z(n39444) );
  OR U48564 ( .A(n39447), .B(n39448), .Z(n39443) );
  NAND U48565 ( .A(n39449), .B(n39450), .Z(n39341) );
  OR U48566 ( .A(n39451), .B(n39452), .Z(n39450) );
  OR U48567 ( .A(n39453), .B(n39454), .Z(n39449) );
  ANDN U48568 ( .B(n39455), .A(n39456), .Z(n39342) );
  IV U48569 ( .A(n39457), .Z(n39455) );
  XNOR U48570 ( .A(n39422), .B(n39421), .Z(N61905) );
  XOR U48571 ( .A(n39441), .B(n39440), .Z(n39421) );
  XNOR U48572 ( .A(n39456), .B(n39457), .Z(n39440) );
  XNOR U48573 ( .A(n39451), .B(n39452), .Z(n39457) );
  XNOR U48574 ( .A(n39453), .B(n39454), .Z(n39452) );
  XNOR U48575 ( .A(y[2437]), .B(x[2437]), .Z(n39454) );
  XNOR U48576 ( .A(y[2438]), .B(x[2438]), .Z(n39453) );
  XNOR U48577 ( .A(y[2436]), .B(x[2436]), .Z(n39451) );
  XNOR U48578 ( .A(n39445), .B(n39446), .Z(n39456) );
  XNOR U48579 ( .A(y[2433]), .B(x[2433]), .Z(n39446) );
  XNOR U48580 ( .A(n39447), .B(n39448), .Z(n39445) );
  XNOR U48581 ( .A(y[2434]), .B(x[2434]), .Z(n39448) );
  XNOR U48582 ( .A(y[2435]), .B(x[2435]), .Z(n39447) );
  XNOR U48583 ( .A(n39438), .B(n39437), .Z(n39441) );
  XNOR U48584 ( .A(n39433), .B(n39434), .Z(n39437) );
  XNOR U48585 ( .A(y[2430]), .B(x[2430]), .Z(n39434) );
  XNOR U48586 ( .A(n39435), .B(n39436), .Z(n39433) );
  XNOR U48587 ( .A(y[2431]), .B(x[2431]), .Z(n39436) );
  XNOR U48588 ( .A(y[2432]), .B(x[2432]), .Z(n39435) );
  XNOR U48589 ( .A(n39427), .B(n39428), .Z(n39438) );
  XNOR U48590 ( .A(y[2427]), .B(x[2427]), .Z(n39428) );
  XNOR U48591 ( .A(n39429), .B(n39430), .Z(n39427) );
  XNOR U48592 ( .A(y[2428]), .B(x[2428]), .Z(n39430) );
  XNOR U48593 ( .A(y[2429]), .B(x[2429]), .Z(n39429) );
  XOR U48594 ( .A(n39403), .B(n39404), .Z(n39422) );
  XNOR U48595 ( .A(n39419), .B(n39420), .Z(n39404) );
  XNOR U48596 ( .A(n39414), .B(n39415), .Z(n39420) );
  XNOR U48597 ( .A(n39416), .B(n39417), .Z(n39415) );
  XNOR U48598 ( .A(y[2425]), .B(x[2425]), .Z(n39417) );
  XNOR U48599 ( .A(y[2426]), .B(x[2426]), .Z(n39416) );
  XNOR U48600 ( .A(y[2424]), .B(x[2424]), .Z(n39414) );
  XNOR U48601 ( .A(n39408), .B(n39409), .Z(n39419) );
  XNOR U48602 ( .A(y[2421]), .B(x[2421]), .Z(n39409) );
  XNOR U48603 ( .A(n39410), .B(n39411), .Z(n39408) );
  XNOR U48604 ( .A(y[2422]), .B(x[2422]), .Z(n39411) );
  XNOR U48605 ( .A(y[2423]), .B(x[2423]), .Z(n39410) );
  XOR U48606 ( .A(n39402), .B(n39401), .Z(n39403) );
  XNOR U48607 ( .A(n39397), .B(n39398), .Z(n39401) );
  XNOR U48608 ( .A(y[2418]), .B(x[2418]), .Z(n39398) );
  XNOR U48609 ( .A(n39399), .B(n39400), .Z(n39397) );
  XNOR U48610 ( .A(y[2419]), .B(x[2419]), .Z(n39400) );
  XNOR U48611 ( .A(y[2420]), .B(x[2420]), .Z(n39399) );
  XNOR U48612 ( .A(n39391), .B(n39392), .Z(n39402) );
  XNOR U48613 ( .A(y[2415]), .B(x[2415]), .Z(n39392) );
  XNOR U48614 ( .A(n39393), .B(n39394), .Z(n39391) );
  XNOR U48615 ( .A(y[2416]), .B(x[2416]), .Z(n39394) );
  XNOR U48616 ( .A(y[2417]), .B(x[2417]), .Z(n39393) );
  NAND U48617 ( .A(n39458), .B(n39459), .Z(N61896) );
  NANDN U48618 ( .A(n39460), .B(n39461), .Z(n39459) );
  OR U48619 ( .A(n39462), .B(n39463), .Z(n39461) );
  NAND U48620 ( .A(n39462), .B(n39463), .Z(n39458) );
  XOR U48621 ( .A(n39462), .B(n39464), .Z(N61895) );
  XNOR U48622 ( .A(n39460), .B(n39463), .Z(n39464) );
  AND U48623 ( .A(n39465), .B(n39466), .Z(n39463) );
  NANDN U48624 ( .A(n39467), .B(n39468), .Z(n39466) );
  NANDN U48625 ( .A(n39469), .B(n39470), .Z(n39468) );
  NANDN U48626 ( .A(n39470), .B(n39469), .Z(n39465) );
  NAND U48627 ( .A(n39471), .B(n39472), .Z(n39460) );
  NANDN U48628 ( .A(n39473), .B(n39474), .Z(n39472) );
  OR U48629 ( .A(n39475), .B(n39476), .Z(n39474) );
  NAND U48630 ( .A(n39476), .B(n39475), .Z(n39471) );
  AND U48631 ( .A(n39477), .B(n39478), .Z(n39462) );
  NANDN U48632 ( .A(n39479), .B(n39480), .Z(n39478) );
  NANDN U48633 ( .A(n39481), .B(n39482), .Z(n39480) );
  NANDN U48634 ( .A(n39482), .B(n39481), .Z(n39477) );
  XOR U48635 ( .A(n39476), .B(n39483), .Z(N61894) );
  XOR U48636 ( .A(n39473), .B(n39475), .Z(n39483) );
  XNOR U48637 ( .A(n39469), .B(n39484), .Z(n39475) );
  XNOR U48638 ( .A(n39467), .B(n39470), .Z(n39484) );
  NAND U48639 ( .A(n39485), .B(n39486), .Z(n39470) );
  NAND U48640 ( .A(n39487), .B(n39488), .Z(n39486) );
  OR U48641 ( .A(n39489), .B(n39490), .Z(n39487) );
  NANDN U48642 ( .A(n39491), .B(n39489), .Z(n39485) );
  IV U48643 ( .A(n39490), .Z(n39491) );
  NAND U48644 ( .A(n39492), .B(n39493), .Z(n39467) );
  NAND U48645 ( .A(n39494), .B(n39495), .Z(n39493) );
  NANDN U48646 ( .A(n39496), .B(n39497), .Z(n39494) );
  NANDN U48647 ( .A(n39497), .B(n39496), .Z(n39492) );
  AND U48648 ( .A(n39498), .B(n39499), .Z(n39469) );
  NAND U48649 ( .A(n39500), .B(n39501), .Z(n39499) );
  OR U48650 ( .A(n39502), .B(n39503), .Z(n39500) );
  NANDN U48651 ( .A(n39504), .B(n39502), .Z(n39498) );
  NAND U48652 ( .A(n39505), .B(n39506), .Z(n39473) );
  NANDN U48653 ( .A(n39507), .B(n39508), .Z(n39506) );
  OR U48654 ( .A(n39509), .B(n39510), .Z(n39508) );
  NANDN U48655 ( .A(n39511), .B(n39509), .Z(n39505) );
  IV U48656 ( .A(n39510), .Z(n39511) );
  XNOR U48657 ( .A(n39481), .B(n39512), .Z(n39476) );
  XNOR U48658 ( .A(n39479), .B(n39482), .Z(n39512) );
  NAND U48659 ( .A(n39513), .B(n39514), .Z(n39482) );
  NAND U48660 ( .A(n39515), .B(n39516), .Z(n39514) );
  OR U48661 ( .A(n39517), .B(n39518), .Z(n39515) );
  NANDN U48662 ( .A(n39519), .B(n39517), .Z(n39513) );
  IV U48663 ( .A(n39518), .Z(n39519) );
  NAND U48664 ( .A(n39520), .B(n39521), .Z(n39479) );
  NAND U48665 ( .A(n39522), .B(n39523), .Z(n39521) );
  NANDN U48666 ( .A(n39524), .B(n39525), .Z(n39522) );
  NANDN U48667 ( .A(n39525), .B(n39524), .Z(n39520) );
  AND U48668 ( .A(n39526), .B(n39527), .Z(n39481) );
  NAND U48669 ( .A(n39528), .B(n39529), .Z(n39527) );
  OR U48670 ( .A(n39530), .B(n39531), .Z(n39528) );
  NANDN U48671 ( .A(n39532), .B(n39530), .Z(n39526) );
  XNOR U48672 ( .A(n39507), .B(n39533), .Z(N61893) );
  XOR U48673 ( .A(n39509), .B(n39510), .Z(n39533) );
  XNOR U48674 ( .A(n39523), .B(n39534), .Z(n39510) );
  XOR U48675 ( .A(n39524), .B(n39525), .Z(n39534) );
  XOR U48676 ( .A(n39530), .B(n39535), .Z(n39525) );
  XOR U48677 ( .A(n39529), .B(n39532), .Z(n39535) );
  IV U48678 ( .A(n39531), .Z(n39532) );
  NAND U48679 ( .A(n39536), .B(n39537), .Z(n39531) );
  OR U48680 ( .A(n39538), .B(n39539), .Z(n39537) );
  OR U48681 ( .A(n39540), .B(n39541), .Z(n39536) );
  NAND U48682 ( .A(n39542), .B(n39543), .Z(n39529) );
  OR U48683 ( .A(n39544), .B(n39545), .Z(n39543) );
  OR U48684 ( .A(n39546), .B(n39547), .Z(n39542) );
  NOR U48685 ( .A(n39548), .B(n39549), .Z(n39530) );
  ANDN U48686 ( .B(n39550), .A(n39551), .Z(n39524) );
  XNOR U48687 ( .A(n39517), .B(n39552), .Z(n39523) );
  XNOR U48688 ( .A(n39516), .B(n39518), .Z(n39552) );
  NAND U48689 ( .A(n39553), .B(n39554), .Z(n39518) );
  OR U48690 ( .A(n39555), .B(n39556), .Z(n39554) );
  OR U48691 ( .A(n39557), .B(n39558), .Z(n39553) );
  NAND U48692 ( .A(n39559), .B(n39560), .Z(n39516) );
  OR U48693 ( .A(n39561), .B(n39562), .Z(n39560) );
  OR U48694 ( .A(n39563), .B(n39564), .Z(n39559) );
  ANDN U48695 ( .B(n39565), .A(n39566), .Z(n39517) );
  IV U48696 ( .A(n39567), .Z(n39565) );
  ANDN U48697 ( .B(n39568), .A(n39569), .Z(n39509) );
  XOR U48698 ( .A(n39495), .B(n39570), .Z(n39507) );
  XOR U48699 ( .A(n39496), .B(n39497), .Z(n39570) );
  XOR U48700 ( .A(n39502), .B(n39571), .Z(n39497) );
  XOR U48701 ( .A(n39501), .B(n39504), .Z(n39571) );
  IV U48702 ( .A(n39503), .Z(n39504) );
  NAND U48703 ( .A(n39572), .B(n39573), .Z(n39503) );
  OR U48704 ( .A(n39574), .B(n39575), .Z(n39573) );
  OR U48705 ( .A(n39576), .B(n39577), .Z(n39572) );
  NAND U48706 ( .A(n39578), .B(n39579), .Z(n39501) );
  OR U48707 ( .A(n39580), .B(n39581), .Z(n39579) );
  OR U48708 ( .A(n39582), .B(n39583), .Z(n39578) );
  NOR U48709 ( .A(n39584), .B(n39585), .Z(n39502) );
  ANDN U48710 ( .B(n39586), .A(n39587), .Z(n39496) );
  IV U48711 ( .A(n39588), .Z(n39586) );
  XNOR U48712 ( .A(n39489), .B(n39589), .Z(n39495) );
  XNOR U48713 ( .A(n39488), .B(n39490), .Z(n39589) );
  NAND U48714 ( .A(n39590), .B(n39591), .Z(n39490) );
  OR U48715 ( .A(n39592), .B(n39593), .Z(n39591) );
  OR U48716 ( .A(n39594), .B(n39595), .Z(n39590) );
  NAND U48717 ( .A(n39596), .B(n39597), .Z(n39488) );
  OR U48718 ( .A(n39598), .B(n39599), .Z(n39597) );
  OR U48719 ( .A(n39600), .B(n39601), .Z(n39596) );
  ANDN U48720 ( .B(n39602), .A(n39603), .Z(n39489) );
  IV U48721 ( .A(n39604), .Z(n39602) );
  XNOR U48722 ( .A(n39569), .B(n39568), .Z(N61892) );
  XOR U48723 ( .A(n39588), .B(n39587), .Z(n39568) );
  XNOR U48724 ( .A(n39603), .B(n39604), .Z(n39587) );
  XNOR U48725 ( .A(n39598), .B(n39599), .Z(n39604) );
  XNOR U48726 ( .A(n39600), .B(n39601), .Z(n39599) );
  XNOR U48727 ( .A(y[2413]), .B(x[2413]), .Z(n39601) );
  XNOR U48728 ( .A(y[2414]), .B(x[2414]), .Z(n39600) );
  XNOR U48729 ( .A(y[2412]), .B(x[2412]), .Z(n39598) );
  XNOR U48730 ( .A(n39592), .B(n39593), .Z(n39603) );
  XNOR U48731 ( .A(y[2409]), .B(x[2409]), .Z(n39593) );
  XNOR U48732 ( .A(n39594), .B(n39595), .Z(n39592) );
  XNOR U48733 ( .A(y[2410]), .B(x[2410]), .Z(n39595) );
  XNOR U48734 ( .A(y[2411]), .B(x[2411]), .Z(n39594) );
  XNOR U48735 ( .A(n39585), .B(n39584), .Z(n39588) );
  XNOR U48736 ( .A(n39580), .B(n39581), .Z(n39584) );
  XNOR U48737 ( .A(y[2406]), .B(x[2406]), .Z(n39581) );
  XNOR U48738 ( .A(n39582), .B(n39583), .Z(n39580) );
  XNOR U48739 ( .A(y[2407]), .B(x[2407]), .Z(n39583) );
  XNOR U48740 ( .A(y[2408]), .B(x[2408]), .Z(n39582) );
  XNOR U48741 ( .A(n39574), .B(n39575), .Z(n39585) );
  XNOR U48742 ( .A(y[2403]), .B(x[2403]), .Z(n39575) );
  XNOR U48743 ( .A(n39576), .B(n39577), .Z(n39574) );
  XNOR U48744 ( .A(y[2404]), .B(x[2404]), .Z(n39577) );
  XNOR U48745 ( .A(y[2405]), .B(x[2405]), .Z(n39576) );
  XOR U48746 ( .A(n39550), .B(n39551), .Z(n39569) );
  XNOR U48747 ( .A(n39566), .B(n39567), .Z(n39551) );
  XNOR U48748 ( .A(n39561), .B(n39562), .Z(n39567) );
  XNOR U48749 ( .A(n39563), .B(n39564), .Z(n39562) );
  XNOR U48750 ( .A(y[2401]), .B(x[2401]), .Z(n39564) );
  XNOR U48751 ( .A(y[2402]), .B(x[2402]), .Z(n39563) );
  XNOR U48752 ( .A(y[2400]), .B(x[2400]), .Z(n39561) );
  XNOR U48753 ( .A(n39555), .B(n39556), .Z(n39566) );
  XNOR U48754 ( .A(y[2397]), .B(x[2397]), .Z(n39556) );
  XNOR U48755 ( .A(n39557), .B(n39558), .Z(n39555) );
  XNOR U48756 ( .A(y[2398]), .B(x[2398]), .Z(n39558) );
  XNOR U48757 ( .A(y[2399]), .B(x[2399]), .Z(n39557) );
  XOR U48758 ( .A(n39549), .B(n39548), .Z(n39550) );
  XNOR U48759 ( .A(n39544), .B(n39545), .Z(n39548) );
  XNOR U48760 ( .A(y[2394]), .B(x[2394]), .Z(n39545) );
  XNOR U48761 ( .A(n39546), .B(n39547), .Z(n39544) );
  XNOR U48762 ( .A(y[2395]), .B(x[2395]), .Z(n39547) );
  XNOR U48763 ( .A(y[2396]), .B(x[2396]), .Z(n39546) );
  XNOR U48764 ( .A(n39538), .B(n39539), .Z(n39549) );
  XNOR U48765 ( .A(y[2391]), .B(x[2391]), .Z(n39539) );
  XNOR U48766 ( .A(n39540), .B(n39541), .Z(n39538) );
  XNOR U48767 ( .A(y[2392]), .B(x[2392]), .Z(n39541) );
  XNOR U48768 ( .A(y[2393]), .B(x[2393]), .Z(n39540) );
  NAND U48769 ( .A(n39605), .B(n39606), .Z(N61883) );
  NANDN U48770 ( .A(n39607), .B(n39608), .Z(n39606) );
  OR U48771 ( .A(n39609), .B(n39610), .Z(n39608) );
  NAND U48772 ( .A(n39609), .B(n39610), .Z(n39605) );
  XOR U48773 ( .A(n39609), .B(n39611), .Z(N61882) );
  XNOR U48774 ( .A(n39607), .B(n39610), .Z(n39611) );
  AND U48775 ( .A(n39612), .B(n39613), .Z(n39610) );
  NANDN U48776 ( .A(n39614), .B(n39615), .Z(n39613) );
  NANDN U48777 ( .A(n39616), .B(n39617), .Z(n39615) );
  NANDN U48778 ( .A(n39617), .B(n39616), .Z(n39612) );
  NAND U48779 ( .A(n39618), .B(n39619), .Z(n39607) );
  NANDN U48780 ( .A(n39620), .B(n39621), .Z(n39619) );
  OR U48781 ( .A(n39622), .B(n39623), .Z(n39621) );
  NAND U48782 ( .A(n39623), .B(n39622), .Z(n39618) );
  AND U48783 ( .A(n39624), .B(n39625), .Z(n39609) );
  NANDN U48784 ( .A(n39626), .B(n39627), .Z(n39625) );
  NANDN U48785 ( .A(n39628), .B(n39629), .Z(n39627) );
  NANDN U48786 ( .A(n39629), .B(n39628), .Z(n39624) );
  XOR U48787 ( .A(n39623), .B(n39630), .Z(N61881) );
  XOR U48788 ( .A(n39620), .B(n39622), .Z(n39630) );
  XNOR U48789 ( .A(n39616), .B(n39631), .Z(n39622) );
  XNOR U48790 ( .A(n39614), .B(n39617), .Z(n39631) );
  NAND U48791 ( .A(n39632), .B(n39633), .Z(n39617) );
  NAND U48792 ( .A(n39634), .B(n39635), .Z(n39633) );
  OR U48793 ( .A(n39636), .B(n39637), .Z(n39634) );
  NANDN U48794 ( .A(n39638), .B(n39636), .Z(n39632) );
  IV U48795 ( .A(n39637), .Z(n39638) );
  NAND U48796 ( .A(n39639), .B(n39640), .Z(n39614) );
  NAND U48797 ( .A(n39641), .B(n39642), .Z(n39640) );
  NANDN U48798 ( .A(n39643), .B(n39644), .Z(n39641) );
  NANDN U48799 ( .A(n39644), .B(n39643), .Z(n39639) );
  AND U48800 ( .A(n39645), .B(n39646), .Z(n39616) );
  NAND U48801 ( .A(n39647), .B(n39648), .Z(n39646) );
  OR U48802 ( .A(n39649), .B(n39650), .Z(n39647) );
  NANDN U48803 ( .A(n39651), .B(n39649), .Z(n39645) );
  NAND U48804 ( .A(n39652), .B(n39653), .Z(n39620) );
  NANDN U48805 ( .A(n39654), .B(n39655), .Z(n39653) );
  OR U48806 ( .A(n39656), .B(n39657), .Z(n39655) );
  NANDN U48807 ( .A(n39658), .B(n39656), .Z(n39652) );
  IV U48808 ( .A(n39657), .Z(n39658) );
  XNOR U48809 ( .A(n39628), .B(n39659), .Z(n39623) );
  XNOR U48810 ( .A(n39626), .B(n39629), .Z(n39659) );
  NAND U48811 ( .A(n39660), .B(n39661), .Z(n39629) );
  NAND U48812 ( .A(n39662), .B(n39663), .Z(n39661) );
  OR U48813 ( .A(n39664), .B(n39665), .Z(n39662) );
  NANDN U48814 ( .A(n39666), .B(n39664), .Z(n39660) );
  IV U48815 ( .A(n39665), .Z(n39666) );
  NAND U48816 ( .A(n39667), .B(n39668), .Z(n39626) );
  NAND U48817 ( .A(n39669), .B(n39670), .Z(n39668) );
  NANDN U48818 ( .A(n39671), .B(n39672), .Z(n39669) );
  NANDN U48819 ( .A(n39672), .B(n39671), .Z(n39667) );
  AND U48820 ( .A(n39673), .B(n39674), .Z(n39628) );
  NAND U48821 ( .A(n39675), .B(n39676), .Z(n39674) );
  OR U48822 ( .A(n39677), .B(n39678), .Z(n39675) );
  NANDN U48823 ( .A(n39679), .B(n39677), .Z(n39673) );
  XNOR U48824 ( .A(n39654), .B(n39680), .Z(N61880) );
  XOR U48825 ( .A(n39656), .B(n39657), .Z(n39680) );
  XNOR U48826 ( .A(n39670), .B(n39681), .Z(n39657) );
  XOR U48827 ( .A(n39671), .B(n39672), .Z(n39681) );
  XOR U48828 ( .A(n39677), .B(n39682), .Z(n39672) );
  XOR U48829 ( .A(n39676), .B(n39679), .Z(n39682) );
  IV U48830 ( .A(n39678), .Z(n39679) );
  NAND U48831 ( .A(n39683), .B(n39684), .Z(n39678) );
  OR U48832 ( .A(n39685), .B(n39686), .Z(n39684) );
  OR U48833 ( .A(n39687), .B(n39688), .Z(n39683) );
  NAND U48834 ( .A(n39689), .B(n39690), .Z(n39676) );
  OR U48835 ( .A(n39691), .B(n39692), .Z(n39690) );
  OR U48836 ( .A(n39693), .B(n39694), .Z(n39689) );
  NOR U48837 ( .A(n39695), .B(n39696), .Z(n39677) );
  ANDN U48838 ( .B(n39697), .A(n39698), .Z(n39671) );
  XNOR U48839 ( .A(n39664), .B(n39699), .Z(n39670) );
  XNOR U48840 ( .A(n39663), .B(n39665), .Z(n39699) );
  NAND U48841 ( .A(n39700), .B(n39701), .Z(n39665) );
  OR U48842 ( .A(n39702), .B(n39703), .Z(n39701) );
  OR U48843 ( .A(n39704), .B(n39705), .Z(n39700) );
  NAND U48844 ( .A(n39706), .B(n39707), .Z(n39663) );
  OR U48845 ( .A(n39708), .B(n39709), .Z(n39707) );
  OR U48846 ( .A(n39710), .B(n39711), .Z(n39706) );
  ANDN U48847 ( .B(n39712), .A(n39713), .Z(n39664) );
  IV U48848 ( .A(n39714), .Z(n39712) );
  ANDN U48849 ( .B(n39715), .A(n39716), .Z(n39656) );
  XOR U48850 ( .A(n39642), .B(n39717), .Z(n39654) );
  XOR U48851 ( .A(n39643), .B(n39644), .Z(n39717) );
  XOR U48852 ( .A(n39649), .B(n39718), .Z(n39644) );
  XOR U48853 ( .A(n39648), .B(n39651), .Z(n39718) );
  IV U48854 ( .A(n39650), .Z(n39651) );
  NAND U48855 ( .A(n39719), .B(n39720), .Z(n39650) );
  OR U48856 ( .A(n39721), .B(n39722), .Z(n39720) );
  OR U48857 ( .A(n39723), .B(n39724), .Z(n39719) );
  NAND U48858 ( .A(n39725), .B(n39726), .Z(n39648) );
  OR U48859 ( .A(n39727), .B(n39728), .Z(n39726) );
  OR U48860 ( .A(n39729), .B(n39730), .Z(n39725) );
  NOR U48861 ( .A(n39731), .B(n39732), .Z(n39649) );
  ANDN U48862 ( .B(n39733), .A(n39734), .Z(n39643) );
  IV U48863 ( .A(n39735), .Z(n39733) );
  XNOR U48864 ( .A(n39636), .B(n39736), .Z(n39642) );
  XNOR U48865 ( .A(n39635), .B(n39637), .Z(n39736) );
  NAND U48866 ( .A(n39737), .B(n39738), .Z(n39637) );
  OR U48867 ( .A(n39739), .B(n39740), .Z(n39738) );
  OR U48868 ( .A(n39741), .B(n39742), .Z(n39737) );
  NAND U48869 ( .A(n39743), .B(n39744), .Z(n39635) );
  OR U48870 ( .A(n39745), .B(n39746), .Z(n39744) );
  OR U48871 ( .A(n39747), .B(n39748), .Z(n39743) );
  ANDN U48872 ( .B(n39749), .A(n39750), .Z(n39636) );
  IV U48873 ( .A(n39751), .Z(n39749) );
  XNOR U48874 ( .A(n39716), .B(n39715), .Z(N61879) );
  XOR U48875 ( .A(n39735), .B(n39734), .Z(n39715) );
  XNOR U48876 ( .A(n39750), .B(n39751), .Z(n39734) );
  XNOR U48877 ( .A(n39745), .B(n39746), .Z(n39751) );
  XNOR U48878 ( .A(n39747), .B(n39748), .Z(n39746) );
  XNOR U48879 ( .A(y[2389]), .B(x[2389]), .Z(n39748) );
  XNOR U48880 ( .A(y[2390]), .B(x[2390]), .Z(n39747) );
  XNOR U48881 ( .A(y[2388]), .B(x[2388]), .Z(n39745) );
  XNOR U48882 ( .A(n39739), .B(n39740), .Z(n39750) );
  XNOR U48883 ( .A(y[2385]), .B(x[2385]), .Z(n39740) );
  XNOR U48884 ( .A(n39741), .B(n39742), .Z(n39739) );
  XNOR U48885 ( .A(y[2386]), .B(x[2386]), .Z(n39742) );
  XNOR U48886 ( .A(y[2387]), .B(x[2387]), .Z(n39741) );
  XNOR U48887 ( .A(n39732), .B(n39731), .Z(n39735) );
  XNOR U48888 ( .A(n39727), .B(n39728), .Z(n39731) );
  XNOR U48889 ( .A(y[2382]), .B(x[2382]), .Z(n39728) );
  XNOR U48890 ( .A(n39729), .B(n39730), .Z(n39727) );
  XNOR U48891 ( .A(y[2383]), .B(x[2383]), .Z(n39730) );
  XNOR U48892 ( .A(y[2384]), .B(x[2384]), .Z(n39729) );
  XNOR U48893 ( .A(n39721), .B(n39722), .Z(n39732) );
  XNOR U48894 ( .A(y[2379]), .B(x[2379]), .Z(n39722) );
  XNOR U48895 ( .A(n39723), .B(n39724), .Z(n39721) );
  XNOR U48896 ( .A(y[2380]), .B(x[2380]), .Z(n39724) );
  XNOR U48897 ( .A(y[2381]), .B(x[2381]), .Z(n39723) );
  XOR U48898 ( .A(n39697), .B(n39698), .Z(n39716) );
  XNOR U48899 ( .A(n39713), .B(n39714), .Z(n39698) );
  XNOR U48900 ( .A(n39708), .B(n39709), .Z(n39714) );
  XNOR U48901 ( .A(n39710), .B(n39711), .Z(n39709) );
  XNOR U48902 ( .A(y[2377]), .B(x[2377]), .Z(n39711) );
  XNOR U48903 ( .A(y[2378]), .B(x[2378]), .Z(n39710) );
  XNOR U48904 ( .A(y[2376]), .B(x[2376]), .Z(n39708) );
  XNOR U48905 ( .A(n39702), .B(n39703), .Z(n39713) );
  XNOR U48906 ( .A(y[2373]), .B(x[2373]), .Z(n39703) );
  XNOR U48907 ( .A(n39704), .B(n39705), .Z(n39702) );
  XNOR U48908 ( .A(y[2374]), .B(x[2374]), .Z(n39705) );
  XNOR U48909 ( .A(y[2375]), .B(x[2375]), .Z(n39704) );
  XOR U48910 ( .A(n39696), .B(n39695), .Z(n39697) );
  XNOR U48911 ( .A(n39691), .B(n39692), .Z(n39695) );
  XNOR U48912 ( .A(y[2370]), .B(x[2370]), .Z(n39692) );
  XNOR U48913 ( .A(n39693), .B(n39694), .Z(n39691) );
  XNOR U48914 ( .A(y[2371]), .B(x[2371]), .Z(n39694) );
  XNOR U48915 ( .A(y[2372]), .B(x[2372]), .Z(n39693) );
  XNOR U48916 ( .A(n39685), .B(n39686), .Z(n39696) );
  XNOR U48917 ( .A(y[2367]), .B(x[2367]), .Z(n39686) );
  XNOR U48918 ( .A(n39687), .B(n39688), .Z(n39685) );
  XNOR U48919 ( .A(y[2368]), .B(x[2368]), .Z(n39688) );
  XNOR U48920 ( .A(y[2369]), .B(x[2369]), .Z(n39687) );
  NAND U48921 ( .A(n39752), .B(n39753), .Z(N61870) );
  NANDN U48922 ( .A(n39754), .B(n39755), .Z(n39753) );
  OR U48923 ( .A(n39756), .B(n39757), .Z(n39755) );
  NAND U48924 ( .A(n39756), .B(n39757), .Z(n39752) );
  XOR U48925 ( .A(n39756), .B(n39758), .Z(N61869) );
  XNOR U48926 ( .A(n39754), .B(n39757), .Z(n39758) );
  AND U48927 ( .A(n39759), .B(n39760), .Z(n39757) );
  NANDN U48928 ( .A(n39761), .B(n39762), .Z(n39760) );
  NANDN U48929 ( .A(n39763), .B(n39764), .Z(n39762) );
  NANDN U48930 ( .A(n39764), .B(n39763), .Z(n39759) );
  NAND U48931 ( .A(n39765), .B(n39766), .Z(n39754) );
  NANDN U48932 ( .A(n39767), .B(n39768), .Z(n39766) );
  OR U48933 ( .A(n39769), .B(n39770), .Z(n39768) );
  NAND U48934 ( .A(n39770), .B(n39769), .Z(n39765) );
  AND U48935 ( .A(n39771), .B(n39772), .Z(n39756) );
  NANDN U48936 ( .A(n39773), .B(n39774), .Z(n39772) );
  NANDN U48937 ( .A(n39775), .B(n39776), .Z(n39774) );
  NANDN U48938 ( .A(n39776), .B(n39775), .Z(n39771) );
  XOR U48939 ( .A(n39770), .B(n39777), .Z(N61868) );
  XOR U48940 ( .A(n39767), .B(n39769), .Z(n39777) );
  XNOR U48941 ( .A(n39763), .B(n39778), .Z(n39769) );
  XNOR U48942 ( .A(n39761), .B(n39764), .Z(n39778) );
  NAND U48943 ( .A(n39779), .B(n39780), .Z(n39764) );
  NAND U48944 ( .A(n39781), .B(n39782), .Z(n39780) );
  OR U48945 ( .A(n39783), .B(n39784), .Z(n39781) );
  NANDN U48946 ( .A(n39785), .B(n39783), .Z(n39779) );
  IV U48947 ( .A(n39784), .Z(n39785) );
  NAND U48948 ( .A(n39786), .B(n39787), .Z(n39761) );
  NAND U48949 ( .A(n39788), .B(n39789), .Z(n39787) );
  NANDN U48950 ( .A(n39790), .B(n39791), .Z(n39788) );
  NANDN U48951 ( .A(n39791), .B(n39790), .Z(n39786) );
  AND U48952 ( .A(n39792), .B(n39793), .Z(n39763) );
  NAND U48953 ( .A(n39794), .B(n39795), .Z(n39793) );
  OR U48954 ( .A(n39796), .B(n39797), .Z(n39794) );
  NANDN U48955 ( .A(n39798), .B(n39796), .Z(n39792) );
  NAND U48956 ( .A(n39799), .B(n39800), .Z(n39767) );
  NANDN U48957 ( .A(n39801), .B(n39802), .Z(n39800) );
  OR U48958 ( .A(n39803), .B(n39804), .Z(n39802) );
  NANDN U48959 ( .A(n39805), .B(n39803), .Z(n39799) );
  IV U48960 ( .A(n39804), .Z(n39805) );
  XNOR U48961 ( .A(n39775), .B(n39806), .Z(n39770) );
  XNOR U48962 ( .A(n39773), .B(n39776), .Z(n39806) );
  NAND U48963 ( .A(n39807), .B(n39808), .Z(n39776) );
  NAND U48964 ( .A(n39809), .B(n39810), .Z(n39808) );
  OR U48965 ( .A(n39811), .B(n39812), .Z(n39809) );
  NANDN U48966 ( .A(n39813), .B(n39811), .Z(n39807) );
  IV U48967 ( .A(n39812), .Z(n39813) );
  NAND U48968 ( .A(n39814), .B(n39815), .Z(n39773) );
  NAND U48969 ( .A(n39816), .B(n39817), .Z(n39815) );
  NANDN U48970 ( .A(n39818), .B(n39819), .Z(n39816) );
  NANDN U48971 ( .A(n39819), .B(n39818), .Z(n39814) );
  AND U48972 ( .A(n39820), .B(n39821), .Z(n39775) );
  NAND U48973 ( .A(n39822), .B(n39823), .Z(n39821) );
  OR U48974 ( .A(n39824), .B(n39825), .Z(n39822) );
  NANDN U48975 ( .A(n39826), .B(n39824), .Z(n39820) );
  XNOR U48976 ( .A(n39801), .B(n39827), .Z(N61867) );
  XOR U48977 ( .A(n39803), .B(n39804), .Z(n39827) );
  XNOR U48978 ( .A(n39817), .B(n39828), .Z(n39804) );
  XOR U48979 ( .A(n39818), .B(n39819), .Z(n39828) );
  XOR U48980 ( .A(n39824), .B(n39829), .Z(n39819) );
  XOR U48981 ( .A(n39823), .B(n39826), .Z(n39829) );
  IV U48982 ( .A(n39825), .Z(n39826) );
  NAND U48983 ( .A(n39830), .B(n39831), .Z(n39825) );
  OR U48984 ( .A(n39832), .B(n39833), .Z(n39831) );
  OR U48985 ( .A(n39834), .B(n39835), .Z(n39830) );
  NAND U48986 ( .A(n39836), .B(n39837), .Z(n39823) );
  OR U48987 ( .A(n39838), .B(n39839), .Z(n39837) );
  OR U48988 ( .A(n39840), .B(n39841), .Z(n39836) );
  NOR U48989 ( .A(n39842), .B(n39843), .Z(n39824) );
  ANDN U48990 ( .B(n39844), .A(n39845), .Z(n39818) );
  XNOR U48991 ( .A(n39811), .B(n39846), .Z(n39817) );
  XNOR U48992 ( .A(n39810), .B(n39812), .Z(n39846) );
  NAND U48993 ( .A(n39847), .B(n39848), .Z(n39812) );
  OR U48994 ( .A(n39849), .B(n39850), .Z(n39848) );
  OR U48995 ( .A(n39851), .B(n39852), .Z(n39847) );
  NAND U48996 ( .A(n39853), .B(n39854), .Z(n39810) );
  OR U48997 ( .A(n39855), .B(n39856), .Z(n39854) );
  OR U48998 ( .A(n39857), .B(n39858), .Z(n39853) );
  ANDN U48999 ( .B(n39859), .A(n39860), .Z(n39811) );
  IV U49000 ( .A(n39861), .Z(n39859) );
  ANDN U49001 ( .B(n39862), .A(n39863), .Z(n39803) );
  XOR U49002 ( .A(n39789), .B(n39864), .Z(n39801) );
  XOR U49003 ( .A(n39790), .B(n39791), .Z(n39864) );
  XOR U49004 ( .A(n39796), .B(n39865), .Z(n39791) );
  XOR U49005 ( .A(n39795), .B(n39798), .Z(n39865) );
  IV U49006 ( .A(n39797), .Z(n39798) );
  NAND U49007 ( .A(n39866), .B(n39867), .Z(n39797) );
  OR U49008 ( .A(n39868), .B(n39869), .Z(n39867) );
  OR U49009 ( .A(n39870), .B(n39871), .Z(n39866) );
  NAND U49010 ( .A(n39872), .B(n39873), .Z(n39795) );
  OR U49011 ( .A(n39874), .B(n39875), .Z(n39873) );
  OR U49012 ( .A(n39876), .B(n39877), .Z(n39872) );
  NOR U49013 ( .A(n39878), .B(n39879), .Z(n39796) );
  ANDN U49014 ( .B(n39880), .A(n39881), .Z(n39790) );
  IV U49015 ( .A(n39882), .Z(n39880) );
  XNOR U49016 ( .A(n39783), .B(n39883), .Z(n39789) );
  XNOR U49017 ( .A(n39782), .B(n39784), .Z(n39883) );
  NAND U49018 ( .A(n39884), .B(n39885), .Z(n39784) );
  OR U49019 ( .A(n39886), .B(n39887), .Z(n39885) );
  OR U49020 ( .A(n39888), .B(n39889), .Z(n39884) );
  NAND U49021 ( .A(n39890), .B(n39891), .Z(n39782) );
  OR U49022 ( .A(n39892), .B(n39893), .Z(n39891) );
  OR U49023 ( .A(n39894), .B(n39895), .Z(n39890) );
  ANDN U49024 ( .B(n39896), .A(n39897), .Z(n39783) );
  IV U49025 ( .A(n39898), .Z(n39896) );
  XNOR U49026 ( .A(n39863), .B(n39862), .Z(N61866) );
  XOR U49027 ( .A(n39882), .B(n39881), .Z(n39862) );
  XNOR U49028 ( .A(n39897), .B(n39898), .Z(n39881) );
  XNOR U49029 ( .A(n39892), .B(n39893), .Z(n39898) );
  XNOR U49030 ( .A(n39894), .B(n39895), .Z(n39893) );
  XNOR U49031 ( .A(y[2365]), .B(x[2365]), .Z(n39895) );
  XNOR U49032 ( .A(y[2366]), .B(x[2366]), .Z(n39894) );
  XNOR U49033 ( .A(y[2364]), .B(x[2364]), .Z(n39892) );
  XNOR U49034 ( .A(n39886), .B(n39887), .Z(n39897) );
  XNOR U49035 ( .A(y[2361]), .B(x[2361]), .Z(n39887) );
  XNOR U49036 ( .A(n39888), .B(n39889), .Z(n39886) );
  XNOR U49037 ( .A(y[2362]), .B(x[2362]), .Z(n39889) );
  XNOR U49038 ( .A(y[2363]), .B(x[2363]), .Z(n39888) );
  XNOR U49039 ( .A(n39879), .B(n39878), .Z(n39882) );
  XNOR U49040 ( .A(n39874), .B(n39875), .Z(n39878) );
  XNOR U49041 ( .A(y[2358]), .B(x[2358]), .Z(n39875) );
  XNOR U49042 ( .A(n39876), .B(n39877), .Z(n39874) );
  XNOR U49043 ( .A(y[2359]), .B(x[2359]), .Z(n39877) );
  XNOR U49044 ( .A(y[2360]), .B(x[2360]), .Z(n39876) );
  XNOR U49045 ( .A(n39868), .B(n39869), .Z(n39879) );
  XNOR U49046 ( .A(y[2355]), .B(x[2355]), .Z(n39869) );
  XNOR U49047 ( .A(n39870), .B(n39871), .Z(n39868) );
  XNOR U49048 ( .A(y[2356]), .B(x[2356]), .Z(n39871) );
  XNOR U49049 ( .A(y[2357]), .B(x[2357]), .Z(n39870) );
  XOR U49050 ( .A(n39844), .B(n39845), .Z(n39863) );
  XNOR U49051 ( .A(n39860), .B(n39861), .Z(n39845) );
  XNOR U49052 ( .A(n39855), .B(n39856), .Z(n39861) );
  XNOR U49053 ( .A(n39857), .B(n39858), .Z(n39856) );
  XNOR U49054 ( .A(y[2353]), .B(x[2353]), .Z(n39858) );
  XNOR U49055 ( .A(y[2354]), .B(x[2354]), .Z(n39857) );
  XNOR U49056 ( .A(y[2352]), .B(x[2352]), .Z(n39855) );
  XNOR U49057 ( .A(n39849), .B(n39850), .Z(n39860) );
  XNOR U49058 ( .A(y[2349]), .B(x[2349]), .Z(n39850) );
  XNOR U49059 ( .A(n39851), .B(n39852), .Z(n39849) );
  XNOR U49060 ( .A(y[2350]), .B(x[2350]), .Z(n39852) );
  XNOR U49061 ( .A(y[2351]), .B(x[2351]), .Z(n39851) );
  XOR U49062 ( .A(n39843), .B(n39842), .Z(n39844) );
  XNOR U49063 ( .A(n39838), .B(n39839), .Z(n39842) );
  XNOR U49064 ( .A(y[2346]), .B(x[2346]), .Z(n39839) );
  XNOR U49065 ( .A(n39840), .B(n39841), .Z(n39838) );
  XNOR U49066 ( .A(y[2347]), .B(x[2347]), .Z(n39841) );
  XNOR U49067 ( .A(y[2348]), .B(x[2348]), .Z(n39840) );
  XNOR U49068 ( .A(n39832), .B(n39833), .Z(n39843) );
  XNOR U49069 ( .A(y[2343]), .B(x[2343]), .Z(n39833) );
  XNOR U49070 ( .A(n39834), .B(n39835), .Z(n39832) );
  XNOR U49071 ( .A(y[2344]), .B(x[2344]), .Z(n39835) );
  XNOR U49072 ( .A(y[2345]), .B(x[2345]), .Z(n39834) );
  NAND U49073 ( .A(n39899), .B(n39900), .Z(N61857) );
  NANDN U49074 ( .A(n39901), .B(n39902), .Z(n39900) );
  OR U49075 ( .A(n39903), .B(n39904), .Z(n39902) );
  NAND U49076 ( .A(n39903), .B(n39904), .Z(n39899) );
  XOR U49077 ( .A(n39903), .B(n39905), .Z(N61856) );
  XNOR U49078 ( .A(n39901), .B(n39904), .Z(n39905) );
  AND U49079 ( .A(n39906), .B(n39907), .Z(n39904) );
  NANDN U49080 ( .A(n39908), .B(n39909), .Z(n39907) );
  NANDN U49081 ( .A(n39910), .B(n39911), .Z(n39909) );
  NANDN U49082 ( .A(n39911), .B(n39910), .Z(n39906) );
  NAND U49083 ( .A(n39912), .B(n39913), .Z(n39901) );
  NANDN U49084 ( .A(n39914), .B(n39915), .Z(n39913) );
  OR U49085 ( .A(n39916), .B(n39917), .Z(n39915) );
  NAND U49086 ( .A(n39917), .B(n39916), .Z(n39912) );
  AND U49087 ( .A(n39918), .B(n39919), .Z(n39903) );
  NANDN U49088 ( .A(n39920), .B(n39921), .Z(n39919) );
  NANDN U49089 ( .A(n39922), .B(n39923), .Z(n39921) );
  NANDN U49090 ( .A(n39923), .B(n39922), .Z(n39918) );
  XOR U49091 ( .A(n39917), .B(n39924), .Z(N61855) );
  XOR U49092 ( .A(n39914), .B(n39916), .Z(n39924) );
  XNOR U49093 ( .A(n39910), .B(n39925), .Z(n39916) );
  XNOR U49094 ( .A(n39908), .B(n39911), .Z(n39925) );
  NAND U49095 ( .A(n39926), .B(n39927), .Z(n39911) );
  NAND U49096 ( .A(n39928), .B(n39929), .Z(n39927) );
  OR U49097 ( .A(n39930), .B(n39931), .Z(n39928) );
  NANDN U49098 ( .A(n39932), .B(n39930), .Z(n39926) );
  IV U49099 ( .A(n39931), .Z(n39932) );
  NAND U49100 ( .A(n39933), .B(n39934), .Z(n39908) );
  NAND U49101 ( .A(n39935), .B(n39936), .Z(n39934) );
  NANDN U49102 ( .A(n39937), .B(n39938), .Z(n39935) );
  NANDN U49103 ( .A(n39938), .B(n39937), .Z(n39933) );
  AND U49104 ( .A(n39939), .B(n39940), .Z(n39910) );
  NAND U49105 ( .A(n39941), .B(n39942), .Z(n39940) );
  OR U49106 ( .A(n39943), .B(n39944), .Z(n39941) );
  NANDN U49107 ( .A(n39945), .B(n39943), .Z(n39939) );
  NAND U49108 ( .A(n39946), .B(n39947), .Z(n39914) );
  NANDN U49109 ( .A(n39948), .B(n39949), .Z(n39947) );
  OR U49110 ( .A(n39950), .B(n39951), .Z(n39949) );
  NANDN U49111 ( .A(n39952), .B(n39950), .Z(n39946) );
  IV U49112 ( .A(n39951), .Z(n39952) );
  XNOR U49113 ( .A(n39922), .B(n39953), .Z(n39917) );
  XNOR U49114 ( .A(n39920), .B(n39923), .Z(n39953) );
  NAND U49115 ( .A(n39954), .B(n39955), .Z(n39923) );
  NAND U49116 ( .A(n39956), .B(n39957), .Z(n39955) );
  OR U49117 ( .A(n39958), .B(n39959), .Z(n39956) );
  NANDN U49118 ( .A(n39960), .B(n39958), .Z(n39954) );
  IV U49119 ( .A(n39959), .Z(n39960) );
  NAND U49120 ( .A(n39961), .B(n39962), .Z(n39920) );
  NAND U49121 ( .A(n39963), .B(n39964), .Z(n39962) );
  NANDN U49122 ( .A(n39965), .B(n39966), .Z(n39963) );
  NANDN U49123 ( .A(n39966), .B(n39965), .Z(n39961) );
  AND U49124 ( .A(n39967), .B(n39968), .Z(n39922) );
  NAND U49125 ( .A(n39969), .B(n39970), .Z(n39968) );
  OR U49126 ( .A(n39971), .B(n39972), .Z(n39969) );
  NANDN U49127 ( .A(n39973), .B(n39971), .Z(n39967) );
  XNOR U49128 ( .A(n39948), .B(n39974), .Z(N61854) );
  XOR U49129 ( .A(n39950), .B(n39951), .Z(n39974) );
  XNOR U49130 ( .A(n39964), .B(n39975), .Z(n39951) );
  XOR U49131 ( .A(n39965), .B(n39966), .Z(n39975) );
  XOR U49132 ( .A(n39971), .B(n39976), .Z(n39966) );
  XOR U49133 ( .A(n39970), .B(n39973), .Z(n39976) );
  IV U49134 ( .A(n39972), .Z(n39973) );
  NAND U49135 ( .A(n39977), .B(n39978), .Z(n39972) );
  OR U49136 ( .A(n39979), .B(n39980), .Z(n39978) );
  OR U49137 ( .A(n39981), .B(n39982), .Z(n39977) );
  NAND U49138 ( .A(n39983), .B(n39984), .Z(n39970) );
  OR U49139 ( .A(n39985), .B(n39986), .Z(n39984) );
  OR U49140 ( .A(n39987), .B(n39988), .Z(n39983) );
  NOR U49141 ( .A(n39989), .B(n39990), .Z(n39971) );
  ANDN U49142 ( .B(n39991), .A(n39992), .Z(n39965) );
  XNOR U49143 ( .A(n39958), .B(n39993), .Z(n39964) );
  XNOR U49144 ( .A(n39957), .B(n39959), .Z(n39993) );
  NAND U49145 ( .A(n39994), .B(n39995), .Z(n39959) );
  OR U49146 ( .A(n39996), .B(n39997), .Z(n39995) );
  OR U49147 ( .A(n39998), .B(n39999), .Z(n39994) );
  NAND U49148 ( .A(n40000), .B(n40001), .Z(n39957) );
  OR U49149 ( .A(n40002), .B(n40003), .Z(n40001) );
  OR U49150 ( .A(n40004), .B(n40005), .Z(n40000) );
  ANDN U49151 ( .B(n40006), .A(n40007), .Z(n39958) );
  IV U49152 ( .A(n40008), .Z(n40006) );
  ANDN U49153 ( .B(n40009), .A(n40010), .Z(n39950) );
  XOR U49154 ( .A(n39936), .B(n40011), .Z(n39948) );
  XOR U49155 ( .A(n39937), .B(n39938), .Z(n40011) );
  XOR U49156 ( .A(n39943), .B(n40012), .Z(n39938) );
  XOR U49157 ( .A(n39942), .B(n39945), .Z(n40012) );
  IV U49158 ( .A(n39944), .Z(n39945) );
  NAND U49159 ( .A(n40013), .B(n40014), .Z(n39944) );
  OR U49160 ( .A(n40015), .B(n40016), .Z(n40014) );
  OR U49161 ( .A(n40017), .B(n40018), .Z(n40013) );
  NAND U49162 ( .A(n40019), .B(n40020), .Z(n39942) );
  OR U49163 ( .A(n40021), .B(n40022), .Z(n40020) );
  OR U49164 ( .A(n40023), .B(n40024), .Z(n40019) );
  NOR U49165 ( .A(n40025), .B(n40026), .Z(n39943) );
  ANDN U49166 ( .B(n40027), .A(n40028), .Z(n39937) );
  IV U49167 ( .A(n40029), .Z(n40027) );
  XNOR U49168 ( .A(n39930), .B(n40030), .Z(n39936) );
  XNOR U49169 ( .A(n39929), .B(n39931), .Z(n40030) );
  NAND U49170 ( .A(n40031), .B(n40032), .Z(n39931) );
  OR U49171 ( .A(n40033), .B(n40034), .Z(n40032) );
  OR U49172 ( .A(n40035), .B(n40036), .Z(n40031) );
  NAND U49173 ( .A(n40037), .B(n40038), .Z(n39929) );
  OR U49174 ( .A(n40039), .B(n40040), .Z(n40038) );
  OR U49175 ( .A(n40041), .B(n40042), .Z(n40037) );
  ANDN U49176 ( .B(n40043), .A(n40044), .Z(n39930) );
  IV U49177 ( .A(n40045), .Z(n40043) );
  XNOR U49178 ( .A(n40010), .B(n40009), .Z(N61853) );
  XOR U49179 ( .A(n40029), .B(n40028), .Z(n40009) );
  XNOR U49180 ( .A(n40044), .B(n40045), .Z(n40028) );
  XNOR U49181 ( .A(n40039), .B(n40040), .Z(n40045) );
  XNOR U49182 ( .A(n40041), .B(n40042), .Z(n40040) );
  XNOR U49183 ( .A(y[2341]), .B(x[2341]), .Z(n40042) );
  XNOR U49184 ( .A(y[2342]), .B(x[2342]), .Z(n40041) );
  XNOR U49185 ( .A(y[2340]), .B(x[2340]), .Z(n40039) );
  XNOR U49186 ( .A(n40033), .B(n40034), .Z(n40044) );
  XNOR U49187 ( .A(y[2337]), .B(x[2337]), .Z(n40034) );
  XNOR U49188 ( .A(n40035), .B(n40036), .Z(n40033) );
  XNOR U49189 ( .A(y[2338]), .B(x[2338]), .Z(n40036) );
  XNOR U49190 ( .A(y[2339]), .B(x[2339]), .Z(n40035) );
  XNOR U49191 ( .A(n40026), .B(n40025), .Z(n40029) );
  XNOR U49192 ( .A(n40021), .B(n40022), .Z(n40025) );
  XNOR U49193 ( .A(y[2334]), .B(x[2334]), .Z(n40022) );
  XNOR U49194 ( .A(n40023), .B(n40024), .Z(n40021) );
  XNOR U49195 ( .A(y[2335]), .B(x[2335]), .Z(n40024) );
  XNOR U49196 ( .A(y[2336]), .B(x[2336]), .Z(n40023) );
  XNOR U49197 ( .A(n40015), .B(n40016), .Z(n40026) );
  XNOR U49198 ( .A(y[2331]), .B(x[2331]), .Z(n40016) );
  XNOR U49199 ( .A(n40017), .B(n40018), .Z(n40015) );
  XNOR U49200 ( .A(y[2332]), .B(x[2332]), .Z(n40018) );
  XNOR U49201 ( .A(y[2333]), .B(x[2333]), .Z(n40017) );
  XOR U49202 ( .A(n39991), .B(n39992), .Z(n40010) );
  XNOR U49203 ( .A(n40007), .B(n40008), .Z(n39992) );
  XNOR U49204 ( .A(n40002), .B(n40003), .Z(n40008) );
  XNOR U49205 ( .A(n40004), .B(n40005), .Z(n40003) );
  XNOR U49206 ( .A(y[2329]), .B(x[2329]), .Z(n40005) );
  XNOR U49207 ( .A(y[2330]), .B(x[2330]), .Z(n40004) );
  XNOR U49208 ( .A(y[2328]), .B(x[2328]), .Z(n40002) );
  XNOR U49209 ( .A(n39996), .B(n39997), .Z(n40007) );
  XNOR U49210 ( .A(y[2325]), .B(x[2325]), .Z(n39997) );
  XNOR U49211 ( .A(n39998), .B(n39999), .Z(n39996) );
  XNOR U49212 ( .A(y[2326]), .B(x[2326]), .Z(n39999) );
  XNOR U49213 ( .A(y[2327]), .B(x[2327]), .Z(n39998) );
  XOR U49214 ( .A(n39990), .B(n39989), .Z(n39991) );
  XNOR U49215 ( .A(n39985), .B(n39986), .Z(n39989) );
  XNOR U49216 ( .A(y[2322]), .B(x[2322]), .Z(n39986) );
  XNOR U49217 ( .A(n39987), .B(n39988), .Z(n39985) );
  XNOR U49218 ( .A(y[2323]), .B(x[2323]), .Z(n39988) );
  XNOR U49219 ( .A(y[2324]), .B(x[2324]), .Z(n39987) );
  XNOR U49220 ( .A(n39979), .B(n39980), .Z(n39990) );
  XNOR U49221 ( .A(y[2319]), .B(x[2319]), .Z(n39980) );
  XNOR U49222 ( .A(n39981), .B(n39982), .Z(n39979) );
  XNOR U49223 ( .A(y[2320]), .B(x[2320]), .Z(n39982) );
  XNOR U49224 ( .A(y[2321]), .B(x[2321]), .Z(n39981) );
  NAND U49225 ( .A(n40046), .B(n40047), .Z(N61844) );
  NANDN U49226 ( .A(n40048), .B(n40049), .Z(n40047) );
  OR U49227 ( .A(n40050), .B(n40051), .Z(n40049) );
  NAND U49228 ( .A(n40050), .B(n40051), .Z(n40046) );
  XOR U49229 ( .A(n40050), .B(n40052), .Z(N61843) );
  XNOR U49230 ( .A(n40048), .B(n40051), .Z(n40052) );
  AND U49231 ( .A(n40053), .B(n40054), .Z(n40051) );
  NANDN U49232 ( .A(n40055), .B(n40056), .Z(n40054) );
  NANDN U49233 ( .A(n40057), .B(n40058), .Z(n40056) );
  NANDN U49234 ( .A(n40058), .B(n40057), .Z(n40053) );
  NAND U49235 ( .A(n40059), .B(n40060), .Z(n40048) );
  NANDN U49236 ( .A(n40061), .B(n40062), .Z(n40060) );
  OR U49237 ( .A(n40063), .B(n40064), .Z(n40062) );
  NAND U49238 ( .A(n40064), .B(n40063), .Z(n40059) );
  AND U49239 ( .A(n40065), .B(n40066), .Z(n40050) );
  NANDN U49240 ( .A(n40067), .B(n40068), .Z(n40066) );
  NANDN U49241 ( .A(n40069), .B(n40070), .Z(n40068) );
  NANDN U49242 ( .A(n40070), .B(n40069), .Z(n40065) );
  XOR U49243 ( .A(n40064), .B(n40071), .Z(N61842) );
  XOR U49244 ( .A(n40061), .B(n40063), .Z(n40071) );
  XNOR U49245 ( .A(n40057), .B(n40072), .Z(n40063) );
  XNOR U49246 ( .A(n40055), .B(n40058), .Z(n40072) );
  NAND U49247 ( .A(n40073), .B(n40074), .Z(n40058) );
  NAND U49248 ( .A(n40075), .B(n40076), .Z(n40074) );
  OR U49249 ( .A(n40077), .B(n40078), .Z(n40075) );
  NANDN U49250 ( .A(n40079), .B(n40077), .Z(n40073) );
  IV U49251 ( .A(n40078), .Z(n40079) );
  NAND U49252 ( .A(n40080), .B(n40081), .Z(n40055) );
  NAND U49253 ( .A(n40082), .B(n40083), .Z(n40081) );
  NANDN U49254 ( .A(n40084), .B(n40085), .Z(n40082) );
  NANDN U49255 ( .A(n40085), .B(n40084), .Z(n40080) );
  AND U49256 ( .A(n40086), .B(n40087), .Z(n40057) );
  NAND U49257 ( .A(n40088), .B(n40089), .Z(n40087) );
  OR U49258 ( .A(n40090), .B(n40091), .Z(n40088) );
  NANDN U49259 ( .A(n40092), .B(n40090), .Z(n40086) );
  NAND U49260 ( .A(n40093), .B(n40094), .Z(n40061) );
  NANDN U49261 ( .A(n40095), .B(n40096), .Z(n40094) );
  OR U49262 ( .A(n40097), .B(n40098), .Z(n40096) );
  NANDN U49263 ( .A(n40099), .B(n40097), .Z(n40093) );
  IV U49264 ( .A(n40098), .Z(n40099) );
  XNOR U49265 ( .A(n40069), .B(n40100), .Z(n40064) );
  XNOR U49266 ( .A(n40067), .B(n40070), .Z(n40100) );
  NAND U49267 ( .A(n40101), .B(n40102), .Z(n40070) );
  NAND U49268 ( .A(n40103), .B(n40104), .Z(n40102) );
  OR U49269 ( .A(n40105), .B(n40106), .Z(n40103) );
  NANDN U49270 ( .A(n40107), .B(n40105), .Z(n40101) );
  IV U49271 ( .A(n40106), .Z(n40107) );
  NAND U49272 ( .A(n40108), .B(n40109), .Z(n40067) );
  NAND U49273 ( .A(n40110), .B(n40111), .Z(n40109) );
  NANDN U49274 ( .A(n40112), .B(n40113), .Z(n40110) );
  NANDN U49275 ( .A(n40113), .B(n40112), .Z(n40108) );
  AND U49276 ( .A(n40114), .B(n40115), .Z(n40069) );
  NAND U49277 ( .A(n40116), .B(n40117), .Z(n40115) );
  OR U49278 ( .A(n40118), .B(n40119), .Z(n40116) );
  NANDN U49279 ( .A(n40120), .B(n40118), .Z(n40114) );
  XNOR U49280 ( .A(n40095), .B(n40121), .Z(N61841) );
  XOR U49281 ( .A(n40097), .B(n40098), .Z(n40121) );
  XNOR U49282 ( .A(n40111), .B(n40122), .Z(n40098) );
  XOR U49283 ( .A(n40112), .B(n40113), .Z(n40122) );
  XOR U49284 ( .A(n40118), .B(n40123), .Z(n40113) );
  XOR U49285 ( .A(n40117), .B(n40120), .Z(n40123) );
  IV U49286 ( .A(n40119), .Z(n40120) );
  NAND U49287 ( .A(n40124), .B(n40125), .Z(n40119) );
  OR U49288 ( .A(n40126), .B(n40127), .Z(n40125) );
  OR U49289 ( .A(n40128), .B(n40129), .Z(n40124) );
  NAND U49290 ( .A(n40130), .B(n40131), .Z(n40117) );
  OR U49291 ( .A(n40132), .B(n40133), .Z(n40131) );
  OR U49292 ( .A(n40134), .B(n40135), .Z(n40130) );
  NOR U49293 ( .A(n40136), .B(n40137), .Z(n40118) );
  ANDN U49294 ( .B(n40138), .A(n40139), .Z(n40112) );
  XNOR U49295 ( .A(n40105), .B(n40140), .Z(n40111) );
  XNOR U49296 ( .A(n40104), .B(n40106), .Z(n40140) );
  NAND U49297 ( .A(n40141), .B(n40142), .Z(n40106) );
  OR U49298 ( .A(n40143), .B(n40144), .Z(n40142) );
  OR U49299 ( .A(n40145), .B(n40146), .Z(n40141) );
  NAND U49300 ( .A(n40147), .B(n40148), .Z(n40104) );
  OR U49301 ( .A(n40149), .B(n40150), .Z(n40148) );
  OR U49302 ( .A(n40151), .B(n40152), .Z(n40147) );
  ANDN U49303 ( .B(n40153), .A(n40154), .Z(n40105) );
  IV U49304 ( .A(n40155), .Z(n40153) );
  ANDN U49305 ( .B(n40156), .A(n40157), .Z(n40097) );
  XOR U49306 ( .A(n40083), .B(n40158), .Z(n40095) );
  XOR U49307 ( .A(n40084), .B(n40085), .Z(n40158) );
  XOR U49308 ( .A(n40090), .B(n40159), .Z(n40085) );
  XOR U49309 ( .A(n40089), .B(n40092), .Z(n40159) );
  IV U49310 ( .A(n40091), .Z(n40092) );
  NAND U49311 ( .A(n40160), .B(n40161), .Z(n40091) );
  OR U49312 ( .A(n40162), .B(n40163), .Z(n40161) );
  OR U49313 ( .A(n40164), .B(n40165), .Z(n40160) );
  NAND U49314 ( .A(n40166), .B(n40167), .Z(n40089) );
  OR U49315 ( .A(n40168), .B(n40169), .Z(n40167) );
  OR U49316 ( .A(n40170), .B(n40171), .Z(n40166) );
  NOR U49317 ( .A(n40172), .B(n40173), .Z(n40090) );
  ANDN U49318 ( .B(n40174), .A(n40175), .Z(n40084) );
  IV U49319 ( .A(n40176), .Z(n40174) );
  XNOR U49320 ( .A(n40077), .B(n40177), .Z(n40083) );
  XNOR U49321 ( .A(n40076), .B(n40078), .Z(n40177) );
  NAND U49322 ( .A(n40178), .B(n40179), .Z(n40078) );
  OR U49323 ( .A(n40180), .B(n40181), .Z(n40179) );
  OR U49324 ( .A(n40182), .B(n40183), .Z(n40178) );
  NAND U49325 ( .A(n40184), .B(n40185), .Z(n40076) );
  OR U49326 ( .A(n40186), .B(n40187), .Z(n40185) );
  OR U49327 ( .A(n40188), .B(n40189), .Z(n40184) );
  ANDN U49328 ( .B(n40190), .A(n40191), .Z(n40077) );
  IV U49329 ( .A(n40192), .Z(n40190) );
  XNOR U49330 ( .A(n40157), .B(n40156), .Z(N61840) );
  XOR U49331 ( .A(n40176), .B(n40175), .Z(n40156) );
  XNOR U49332 ( .A(n40191), .B(n40192), .Z(n40175) );
  XNOR U49333 ( .A(n40186), .B(n40187), .Z(n40192) );
  XNOR U49334 ( .A(n40188), .B(n40189), .Z(n40187) );
  XNOR U49335 ( .A(y[2317]), .B(x[2317]), .Z(n40189) );
  XNOR U49336 ( .A(y[2318]), .B(x[2318]), .Z(n40188) );
  XNOR U49337 ( .A(y[2316]), .B(x[2316]), .Z(n40186) );
  XNOR U49338 ( .A(n40180), .B(n40181), .Z(n40191) );
  XNOR U49339 ( .A(y[2313]), .B(x[2313]), .Z(n40181) );
  XNOR U49340 ( .A(n40182), .B(n40183), .Z(n40180) );
  XNOR U49341 ( .A(y[2314]), .B(x[2314]), .Z(n40183) );
  XNOR U49342 ( .A(y[2315]), .B(x[2315]), .Z(n40182) );
  XNOR U49343 ( .A(n40173), .B(n40172), .Z(n40176) );
  XNOR U49344 ( .A(n40168), .B(n40169), .Z(n40172) );
  XNOR U49345 ( .A(y[2310]), .B(x[2310]), .Z(n40169) );
  XNOR U49346 ( .A(n40170), .B(n40171), .Z(n40168) );
  XNOR U49347 ( .A(y[2311]), .B(x[2311]), .Z(n40171) );
  XNOR U49348 ( .A(y[2312]), .B(x[2312]), .Z(n40170) );
  XNOR U49349 ( .A(n40162), .B(n40163), .Z(n40173) );
  XNOR U49350 ( .A(y[2307]), .B(x[2307]), .Z(n40163) );
  XNOR U49351 ( .A(n40164), .B(n40165), .Z(n40162) );
  XNOR U49352 ( .A(y[2308]), .B(x[2308]), .Z(n40165) );
  XNOR U49353 ( .A(y[2309]), .B(x[2309]), .Z(n40164) );
  XOR U49354 ( .A(n40138), .B(n40139), .Z(n40157) );
  XNOR U49355 ( .A(n40154), .B(n40155), .Z(n40139) );
  XNOR U49356 ( .A(n40149), .B(n40150), .Z(n40155) );
  XNOR U49357 ( .A(n40151), .B(n40152), .Z(n40150) );
  XNOR U49358 ( .A(y[2305]), .B(x[2305]), .Z(n40152) );
  XNOR U49359 ( .A(y[2306]), .B(x[2306]), .Z(n40151) );
  XNOR U49360 ( .A(y[2304]), .B(x[2304]), .Z(n40149) );
  XNOR U49361 ( .A(n40143), .B(n40144), .Z(n40154) );
  XNOR U49362 ( .A(y[2301]), .B(x[2301]), .Z(n40144) );
  XNOR U49363 ( .A(n40145), .B(n40146), .Z(n40143) );
  XNOR U49364 ( .A(y[2302]), .B(x[2302]), .Z(n40146) );
  XNOR U49365 ( .A(y[2303]), .B(x[2303]), .Z(n40145) );
  XOR U49366 ( .A(n40137), .B(n40136), .Z(n40138) );
  XNOR U49367 ( .A(n40132), .B(n40133), .Z(n40136) );
  XNOR U49368 ( .A(y[2298]), .B(x[2298]), .Z(n40133) );
  XNOR U49369 ( .A(n40134), .B(n40135), .Z(n40132) );
  XNOR U49370 ( .A(y[2299]), .B(x[2299]), .Z(n40135) );
  XNOR U49371 ( .A(y[2300]), .B(x[2300]), .Z(n40134) );
  XNOR U49372 ( .A(n40126), .B(n40127), .Z(n40137) );
  XNOR U49373 ( .A(y[2295]), .B(x[2295]), .Z(n40127) );
  XNOR U49374 ( .A(n40128), .B(n40129), .Z(n40126) );
  XNOR U49375 ( .A(y[2296]), .B(x[2296]), .Z(n40129) );
  XNOR U49376 ( .A(y[2297]), .B(x[2297]), .Z(n40128) );
  NAND U49377 ( .A(n40193), .B(n40194), .Z(N61831) );
  NANDN U49378 ( .A(n40195), .B(n40196), .Z(n40194) );
  OR U49379 ( .A(n40197), .B(n40198), .Z(n40196) );
  NAND U49380 ( .A(n40197), .B(n40198), .Z(n40193) );
  XOR U49381 ( .A(n40197), .B(n40199), .Z(N61830) );
  XNOR U49382 ( .A(n40195), .B(n40198), .Z(n40199) );
  AND U49383 ( .A(n40200), .B(n40201), .Z(n40198) );
  NANDN U49384 ( .A(n40202), .B(n40203), .Z(n40201) );
  NANDN U49385 ( .A(n40204), .B(n40205), .Z(n40203) );
  NANDN U49386 ( .A(n40205), .B(n40204), .Z(n40200) );
  NAND U49387 ( .A(n40206), .B(n40207), .Z(n40195) );
  NANDN U49388 ( .A(n40208), .B(n40209), .Z(n40207) );
  OR U49389 ( .A(n40210), .B(n40211), .Z(n40209) );
  NAND U49390 ( .A(n40211), .B(n40210), .Z(n40206) );
  AND U49391 ( .A(n40212), .B(n40213), .Z(n40197) );
  NANDN U49392 ( .A(n40214), .B(n40215), .Z(n40213) );
  NANDN U49393 ( .A(n40216), .B(n40217), .Z(n40215) );
  NANDN U49394 ( .A(n40217), .B(n40216), .Z(n40212) );
  XOR U49395 ( .A(n40211), .B(n40218), .Z(N61829) );
  XOR U49396 ( .A(n40208), .B(n40210), .Z(n40218) );
  XNOR U49397 ( .A(n40204), .B(n40219), .Z(n40210) );
  XNOR U49398 ( .A(n40202), .B(n40205), .Z(n40219) );
  NAND U49399 ( .A(n40220), .B(n40221), .Z(n40205) );
  NAND U49400 ( .A(n40222), .B(n40223), .Z(n40221) );
  OR U49401 ( .A(n40224), .B(n40225), .Z(n40222) );
  NANDN U49402 ( .A(n40226), .B(n40224), .Z(n40220) );
  IV U49403 ( .A(n40225), .Z(n40226) );
  NAND U49404 ( .A(n40227), .B(n40228), .Z(n40202) );
  NAND U49405 ( .A(n40229), .B(n40230), .Z(n40228) );
  NANDN U49406 ( .A(n40231), .B(n40232), .Z(n40229) );
  NANDN U49407 ( .A(n40232), .B(n40231), .Z(n40227) );
  AND U49408 ( .A(n40233), .B(n40234), .Z(n40204) );
  NAND U49409 ( .A(n40235), .B(n40236), .Z(n40234) );
  OR U49410 ( .A(n40237), .B(n40238), .Z(n40235) );
  NANDN U49411 ( .A(n40239), .B(n40237), .Z(n40233) );
  NAND U49412 ( .A(n40240), .B(n40241), .Z(n40208) );
  NANDN U49413 ( .A(n40242), .B(n40243), .Z(n40241) );
  OR U49414 ( .A(n40244), .B(n40245), .Z(n40243) );
  NANDN U49415 ( .A(n40246), .B(n40244), .Z(n40240) );
  IV U49416 ( .A(n40245), .Z(n40246) );
  XNOR U49417 ( .A(n40216), .B(n40247), .Z(n40211) );
  XNOR U49418 ( .A(n40214), .B(n40217), .Z(n40247) );
  NAND U49419 ( .A(n40248), .B(n40249), .Z(n40217) );
  NAND U49420 ( .A(n40250), .B(n40251), .Z(n40249) );
  OR U49421 ( .A(n40252), .B(n40253), .Z(n40250) );
  NANDN U49422 ( .A(n40254), .B(n40252), .Z(n40248) );
  IV U49423 ( .A(n40253), .Z(n40254) );
  NAND U49424 ( .A(n40255), .B(n40256), .Z(n40214) );
  NAND U49425 ( .A(n40257), .B(n40258), .Z(n40256) );
  NANDN U49426 ( .A(n40259), .B(n40260), .Z(n40257) );
  NANDN U49427 ( .A(n40260), .B(n40259), .Z(n40255) );
  AND U49428 ( .A(n40261), .B(n40262), .Z(n40216) );
  NAND U49429 ( .A(n40263), .B(n40264), .Z(n40262) );
  OR U49430 ( .A(n40265), .B(n40266), .Z(n40263) );
  NANDN U49431 ( .A(n40267), .B(n40265), .Z(n40261) );
  XNOR U49432 ( .A(n40242), .B(n40268), .Z(N61828) );
  XOR U49433 ( .A(n40244), .B(n40245), .Z(n40268) );
  XNOR U49434 ( .A(n40258), .B(n40269), .Z(n40245) );
  XOR U49435 ( .A(n40259), .B(n40260), .Z(n40269) );
  XOR U49436 ( .A(n40265), .B(n40270), .Z(n40260) );
  XOR U49437 ( .A(n40264), .B(n40267), .Z(n40270) );
  IV U49438 ( .A(n40266), .Z(n40267) );
  NAND U49439 ( .A(n40271), .B(n40272), .Z(n40266) );
  OR U49440 ( .A(n40273), .B(n40274), .Z(n40272) );
  OR U49441 ( .A(n40275), .B(n40276), .Z(n40271) );
  NAND U49442 ( .A(n40277), .B(n40278), .Z(n40264) );
  OR U49443 ( .A(n40279), .B(n40280), .Z(n40278) );
  OR U49444 ( .A(n40281), .B(n40282), .Z(n40277) );
  NOR U49445 ( .A(n40283), .B(n40284), .Z(n40265) );
  ANDN U49446 ( .B(n40285), .A(n40286), .Z(n40259) );
  XNOR U49447 ( .A(n40252), .B(n40287), .Z(n40258) );
  XNOR U49448 ( .A(n40251), .B(n40253), .Z(n40287) );
  NAND U49449 ( .A(n40288), .B(n40289), .Z(n40253) );
  OR U49450 ( .A(n40290), .B(n40291), .Z(n40289) );
  OR U49451 ( .A(n40292), .B(n40293), .Z(n40288) );
  NAND U49452 ( .A(n40294), .B(n40295), .Z(n40251) );
  OR U49453 ( .A(n40296), .B(n40297), .Z(n40295) );
  OR U49454 ( .A(n40298), .B(n40299), .Z(n40294) );
  ANDN U49455 ( .B(n40300), .A(n40301), .Z(n40252) );
  IV U49456 ( .A(n40302), .Z(n40300) );
  ANDN U49457 ( .B(n40303), .A(n40304), .Z(n40244) );
  XOR U49458 ( .A(n40230), .B(n40305), .Z(n40242) );
  XOR U49459 ( .A(n40231), .B(n40232), .Z(n40305) );
  XOR U49460 ( .A(n40237), .B(n40306), .Z(n40232) );
  XOR U49461 ( .A(n40236), .B(n40239), .Z(n40306) );
  IV U49462 ( .A(n40238), .Z(n40239) );
  NAND U49463 ( .A(n40307), .B(n40308), .Z(n40238) );
  OR U49464 ( .A(n40309), .B(n40310), .Z(n40308) );
  OR U49465 ( .A(n40311), .B(n40312), .Z(n40307) );
  NAND U49466 ( .A(n40313), .B(n40314), .Z(n40236) );
  OR U49467 ( .A(n40315), .B(n40316), .Z(n40314) );
  OR U49468 ( .A(n40317), .B(n40318), .Z(n40313) );
  NOR U49469 ( .A(n40319), .B(n40320), .Z(n40237) );
  ANDN U49470 ( .B(n40321), .A(n40322), .Z(n40231) );
  IV U49471 ( .A(n40323), .Z(n40321) );
  XNOR U49472 ( .A(n40224), .B(n40324), .Z(n40230) );
  XNOR U49473 ( .A(n40223), .B(n40225), .Z(n40324) );
  NAND U49474 ( .A(n40325), .B(n40326), .Z(n40225) );
  OR U49475 ( .A(n40327), .B(n40328), .Z(n40326) );
  OR U49476 ( .A(n40329), .B(n40330), .Z(n40325) );
  NAND U49477 ( .A(n40331), .B(n40332), .Z(n40223) );
  OR U49478 ( .A(n40333), .B(n40334), .Z(n40332) );
  OR U49479 ( .A(n40335), .B(n40336), .Z(n40331) );
  ANDN U49480 ( .B(n40337), .A(n40338), .Z(n40224) );
  IV U49481 ( .A(n40339), .Z(n40337) );
  XNOR U49482 ( .A(n40304), .B(n40303), .Z(N61827) );
  XOR U49483 ( .A(n40323), .B(n40322), .Z(n40303) );
  XNOR U49484 ( .A(n40338), .B(n40339), .Z(n40322) );
  XNOR U49485 ( .A(n40333), .B(n40334), .Z(n40339) );
  XNOR U49486 ( .A(n40335), .B(n40336), .Z(n40334) );
  XNOR U49487 ( .A(y[2293]), .B(x[2293]), .Z(n40336) );
  XNOR U49488 ( .A(y[2294]), .B(x[2294]), .Z(n40335) );
  XNOR U49489 ( .A(y[2292]), .B(x[2292]), .Z(n40333) );
  XNOR U49490 ( .A(n40327), .B(n40328), .Z(n40338) );
  XNOR U49491 ( .A(y[2289]), .B(x[2289]), .Z(n40328) );
  XNOR U49492 ( .A(n40329), .B(n40330), .Z(n40327) );
  XNOR U49493 ( .A(y[2290]), .B(x[2290]), .Z(n40330) );
  XNOR U49494 ( .A(y[2291]), .B(x[2291]), .Z(n40329) );
  XNOR U49495 ( .A(n40320), .B(n40319), .Z(n40323) );
  XNOR U49496 ( .A(n40315), .B(n40316), .Z(n40319) );
  XNOR U49497 ( .A(y[2286]), .B(x[2286]), .Z(n40316) );
  XNOR U49498 ( .A(n40317), .B(n40318), .Z(n40315) );
  XNOR U49499 ( .A(y[2287]), .B(x[2287]), .Z(n40318) );
  XNOR U49500 ( .A(y[2288]), .B(x[2288]), .Z(n40317) );
  XNOR U49501 ( .A(n40309), .B(n40310), .Z(n40320) );
  XNOR U49502 ( .A(y[2283]), .B(x[2283]), .Z(n40310) );
  XNOR U49503 ( .A(n40311), .B(n40312), .Z(n40309) );
  XNOR U49504 ( .A(y[2284]), .B(x[2284]), .Z(n40312) );
  XNOR U49505 ( .A(y[2285]), .B(x[2285]), .Z(n40311) );
  XOR U49506 ( .A(n40285), .B(n40286), .Z(n40304) );
  XNOR U49507 ( .A(n40301), .B(n40302), .Z(n40286) );
  XNOR U49508 ( .A(n40296), .B(n40297), .Z(n40302) );
  XNOR U49509 ( .A(n40298), .B(n40299), .Z(n40297) );
  XNOR U49510 ( .A(y[2281]), .B(x[2281]), .Z(n40299) );
  XNOR U49511 ( .A(y[2282]), .B(x[2282]), .Z(n40298) );
  XNOR U49512 ( .A(y[2280]), .B(x[2280]), .Z(n40296) );
  XNOR U49513 ( .A(n40290), .B(n40291), .Z(n40301) );
  XNOR U49514 ( .A(y[2277]), .B(x[2277]), .Z(n40291) );
  XNOR U49515 ( .A(n40292), .B(n40293), .Z(n40290) );
  XNOR U49516 ( .A(y[2278]), .B(x[2278]), .Z(n40293) );
  XNOR U49517 ( .A(y[2279]), .B(x[2279]), .Z(n40292) );
  XOR U49518 ( .A(n40284), .B(n40283), .Z(n40285) );
  XNOR U49519 ( .A(n40279), .B(n40280), .Z(n40283) );
  XNOR U49520 ( .A(y[2274]), .B(x[2274]), .Z(n40280) );
  XNOR U49521 ( .A(n40281), .B(n40282), .Z(n40279) );
  XNOR U49522 ( .A(y[2275]), .B(x[2275]), .Z(n40282) );
  XNOR U49523 ( .A(y[2276]), .B(x[2276]), .Z(n40281) );
  XNOR U49524 ( .A(n40273), .B(n40274), .Z(n40284) );
  XNOR U49525 ( .A(y[2271]), .B(x[2271]), .Z(n40274) );
  XNOR U49526 ( .A(n40275), .B(n40276), .Z(n40273) );
  XNOR U49527 ( .A(y[2272]), .B(x[2272]), .Z(n40276) );
  XNOR U49528 ( .A(y[2273]), .B(x[2273]), .Z(n40275) );
  NAND U49529 ( .A(n40340), .B(n40341), .Z(N61818) );
  NANDN U49530 ( .A(n40342), .B(n40343), .Z(n40341) );
  OR U49531 ( .A(n40344), .B(n40345), .Z(n40343) );
  NAND U49532 ( .A(n40344), .B(n40345), .Z(n40340) );
  XOR U49533 ( .A(n40344), .B(n40346), .Z(N61817) );
  XNOR U49534 ( .A(n40342), .B(n40345), .Z(n40346) );
  AND U49535 ( .A(n40347), .B(n40348), .Z(n40345) );
  NANDN U49536 ( .A(n40349), .B(n40350), .Z(n40348) );
  NANDN U49537 ( .A(n40351), .B(n40352), .Z(n40350) );
  NANDN U49538 ( .A(n40352), .B(n40351), .Z(n40347) );
  NAND U49539 ( .A(n40353), .B(n40354), .Z(n40342) );
  NANDN U49540 ( .A(n40355), .B(n40356), .Z(n40354) );
  OR U49541 ( .A(n40357), .B(n40358), .Z(n40356) );
  NAND U49542 ( .A(n40358), .B(n40357), .Z(n40353) );
  AND U49543 ( .A(n40359), .B(n40360), .Z(n40344) );
  NANDN U49544 ( .A(n40361), .B(n40362), .Z(n40360) );
  NANDN U49545 ( .A(n40363), .B(n40364), .Z(n40362) );
  NANDN U49546 ( .A(n40364), .B(n40363), .Z(n40359) );
  XOR U49547 ( .A(n40358), .B(n40365), .Z(N61816) );
  XOR U49548 ( .A(n40355), .B(n40357), .Z(n40365) );
  XNOR U49549 ( .A(n40351), .B(n40366), .Z(n40357) );
  XNOR U49550 ( .A(n40349), .B(n40352), .Z(n40366) );
  NAND U49551 ( .A(n40367), .B(n40368), .Z(n40352) );
  NAND U49552 ( .A(n40369), .B(n40370), .Z(n40368) );
  OR U49553 ( .A(n40371), .B(n40372), .Z(n40369) );
  NANDN U49554 ( .A(n40373), .B(n40371), .Z(n40367) );
  IV U49555 ( .A(n40372), .Z(n40373) );
  NAND U49556 ( .A(n40374), .B(n40375), .Z(n40349) );
  NAND U49557 ( .A(n40376), .B(n40377), .Z(n40375) );
  NANDN U49558 ( .A(n40378), .B(n40379), .Z(n40376) );
  NANDN U49559 ( .A(n40379), .B(n40378), .Z(n40374) );
  AND U49560 ( .A(n40380), .B(n40381), .Z(n40351) );
  NAND U49561 ( .A(n40382), .B(n40383), .Z(n40381) );
  OR U49562 ( .A(n40384), .B(n40385), .Z(n40382) );
  NANDN U49563 ( .A(n40386), .B(n40384), .Z(n40380) );
  NAND U49564 ( .A(n40387), .B(n40388), .Z(n40355) );
  NANDN U49565 ( .A(n40389), .B(n40390), .Z(n40388) );
  OR U49566 ( .A(n40391), .B(n40392), .Z(n40390) );
  NANDN U49567 ( .A(n40393), .B(n40391), .Z(n40387) );
  IV U49568 ( .A(n40392), .Z(n40393) );
  XNOR U49569 ( .A(n40363), .B(n40394), .Z(n40358) );
  XNOR U49570 ( .A(n40361), .B(n40364), .Z(n40394) );
  NAND U49571 ( .A(n40395), .B(n40396), .Z(n40364) );
  NAND U49572 ( .A(n40397), .B(n40398), .Z(n40396) );
  OR U49573 ( .A(n40399), .B(n40400), .Z(n40397) );
  NANDN U49574 ( .A(n40401), .B(n40399), .Z(n40395) );
  IV U49575 ( .A(n40400), .Z(n40401) );
  NAND U49576 ( .A(n40402), .B(n40403), .Z(n40361) );
  NAND U49577 ( .A(n40404), .B(n40405), .Z(n40403) );
  NANDN U49578 ( .A(n40406), .B(n40407), .Z(n40404) );
  NANDN U49579 ( .A(n40407), .B(n40406), .Z(n40402) );
  AND U49580 ( .A(n40408), .B(n40409), .Z(n40363) );
  NAND U49581 ( .A(n40410), .B(n40411), .Z(n40409) );
  OR U49582 ( .A(n40412), .B(n40413), .Z(n40410) );
  NANDN U49583 ( .A(n40414), .B(n40412), .Z(n40408) );
  XNOR U49584 ( .A(n40389), .B(n40415), .Z(N61815) );
  XOR U49585 ( .A(n40391), .B(n40392), .Z(n40415) );
  XNOR U49586 ( .A(n40405), .B(n40416), .Z(n40392) );
  XOR U49587 ( .A(n40406), .B(n40407), .Z(n40416) );
  XOR U49588 ( .A(n40412), .B(n40417), .Z(n40407) );
  XOR U49589 ( .A(n40411), .B(n40414), .Z(n40417) );
  IV U49590 ( .A(n40413), .Z(n40414) );
  NAND U49591 ( .A(n40418), .B(n40419), .Z(n40413) );
  OR U49592 ( .A(n40420), .B(n40421), .Z(n40419) );
  OR U49593 ( .A(n40422), .B(n40423), .Z(n40418) );
  NAND U49594 ( .A(n40424), .B(n40425), .Z(n40411) );
  OR U49595 ( .A(n40426), .B(n40427), .Z(n40425) );
  OR U49596 ( .A(n40428), .B(n40429), .Z(n40424) );
  NOR U49597 ( .A(n40430), .B(n40431), .Z(n40412) );
  ANDN U49598 ( .B(n40432), .A(n40433), .Z(n40406) );
  XNOR U49599 ( .A(n40399), .B(n40434), .Z(n40405) );
  XNOR U49600 ( .A(n40398), .B(n40400), .Z(n40434) );
  NAND U49601 ( .A(n40435), .B(n40436), .Z(n40400) );
  OR U49602 ( .A(n40437), .B(n40438), .Z(n40436) );
  OR U49603 ( .A(n40439), .B(n40440), .Z(n40435) );
  NAND U49604 ( .A(n40441), .B(n40442), .Z(n40398) );
  OR U49605 ( .A(n40443), .B(n40444), .Z(n40442) );
  OR U49606 ( .A(n40445), .B(n40446), .Z(n40441) );
  ANDN U49607 ( .B(n40447), .A(n40448), .Z(n40399) );
  IV U49608 ( .A(n40449), .Z(n40447) );
  ANDN U49609 ( .B(n40450), .A(n40451), .Z(n40391) );
  XOR U49610 ( .A(n40377), .B(n40452), .Z(n40389) );
  XOR U49611 ( .A(n40378), .B(n40379), .Z(n40452) );
  XOR U49612 ( .A(n40384), .B(n40453), .Z(n40379) );
  XOR U49613 ( .A(n40383), .B(n40386), .Z(n40453) );
  IV U49614 ( .A(n40385), .Z(n40386) );
  NAND U49615 ( .A(n40454), .B(n40455), .Z(n40385) );
  OR U49616 ( .A(n40456), .B(n40457), .Z(n40455) );
  OR U49617 ( .A(n40458), .B(n40459), .Z(n40454) );
  NAND U49618 ( .A(n40460), .B(n40461), .Z(n40383) );
  OR U49619 ( .A(n40462), .B(n40463), .Z(n40461) );
  OR U49620 ( .A(n40464), .B(n40465), .Z(n40460) );
  NOR U49621 ( .A(n40466), .B(n40467), .Z(n40384) );
  ANDN U49622 ( .B(n40468), .A(n40469), .Z(n40378) );
  IV U49623 ( .A(n40470), .Z(n40468) );
  XNOR U49624 ( .A(n40371), .B(n40471), .Z(n40377) );
  XNOR U49625 ( .A(n40370), .B(n40372), .Z(n40471) );
  NAND U49626 ( .A(n40472), .B(n40473), .Z(n40372) );
  OR U49627 ( .A(n40474), .B(n40475), .Z(n40473) );
  OR U49628 ( .A(n40476), .B(n40477), .Z(n40472) );
  NAND U49629 ( .A(n40478), .B(n40479), .Z(n40370) );
  OR U49630 ( .A(n40480), .B(n40481), .Z(n40479) );
  OR U49631 ( .A(n40482), .B(n40483), .Z(n40478) );
  ANDN U49632 ( .B(n40484), .A(n40485), .Z(n40371) );
  IV U49633 ( .A(n40486), .Z(n40484) );
  XNOR U49634 ( .A(n40451), .B(n40450), .Z(N61814) );
  XOR U49635 ( .A(n40470), .B(n40469), .Z(n40450) );
  XNOR U49636 ( .A(n40485), .B(n40486), .Z(n40469) );
  XNOR U49637 ( .A(n40480), .B(n40481), .Z(n40486) );
  XNOR U49638 ( .A(n40482), .B(n40483), .Z(n40481) );
  XNOR U49639 ( .A(y[2269]), .B(x[2269]), .Z(n40483) );
  XNOR U49640 ( .A(y[2270]), .B(x[2270]), .Z(n40482) );
  XNOR U49641 ( .A(y[2268]), .B(x[2268]), .Z(n40480) );
  XNOR U49642 ( .A(n40474), .B(n40475), .Z(n40485) );
  XNOR U49643 ( .A(y[2265]), .B(x[2265]), .Z(n40475) );
  XNOR U49644 ( .A(n40476), .B(n40477), .Z(n40474) );
  XNOR U49645 ( .A(y[2266]), .B(x[2266]), .Z(n40477) );
  XNOR U49646 ( .A(y[2267]), .B(x[2267]), .Z(n40476) );
  XNOR U49647 ( .A(n40467), .B(n40466), .Z(n40470) );
  XNOR U49648 ( .A(n40462), .B(n40463), .Z(n40466) );
  XNOR U49649 ( .A(y[2262]), .B(x[2262]), .Z(n40463) );
  XNOR U49650 ( .A(n40464), .B(n40465), .Z(n40462) );
  XNOR U49651 ( .A(y[2263]), .B(x[2263]), .Z(n40465) );
  XNOR U49652 ( .A(y[2264]), .B(x[2264]), .Z(n40464) );
  XNOR U49653 ( .A(n40456), .B(n40457), .Z(n40467) );
  XNOR U49654 ( .A(y[2259]), .B(x[2259]), .Z(n40457) );
  XNOR U49655 ( .A(n40458), .B(n40459), .Z(n40456) );
  XNOR U49656 ( .A(y[2260]), .B(x[2260]), .Z(n40459) );
  XNOR U49657 ( .A(y[2261]), .B(x[2261]), .Z(n40458) );
  XOR U49658 ( .A(n40432), .B(n40433), .Z(n40451) );
  XNOR U49659 ( .A(n40448), .B(n40449), .Z(n40433) );
  XNOR U49660 ( .A(n40443), .B(n40444), .Z(n40449) );
  XNOR U49661 ( .A(n40445), .B(n40446), .Z(n40444) );
  XNOR U49662 ( .A(y[2257]), .B(x[2257]), .Z(n40446) );
  XNOR U49663 ( .A(y[2258]), .B(x[2258]), .Z(n40445) );
  XNOR U49664 ( .A(y[2256]), .B(x[2256]), .Z(n40443) );
  XNOR U49665 ( .A(n40437), .B(n40438), .Z(n40448) );
  XNOR U49666 ( .A(y[2253]), .B(x[2253]), .Z(n40438) );
  XNOR U49667 ( .A(n40439), .B(n40440), .Z(n40437) );
  XNOR U49668 ( .A(y[2254]), .B(x[2254]), .Z(n40440) );
  XNOR U49669 ( .A(y[2255]), .B(x[2255]), .Z(n40439) );
  XOR U49670 ( .A(n40431), .B(n40430), .Z(n40432) );
  XNOR U49671 ( .A(n40426), .B(n40427), .Z(n40430) );
  XNOR U49672 ( .A(y[2250]), .B(x[2250]), .Z(n40427) );
  XNOR U49673 ( .A(n40428), .B(n40429), .Z(n40426) );
  XNOR U49674 ( .A(y[2251]), .B(x[2251]), .Z(n40429) );
  XNOR U49675 ( .A(y[2252]), .B(x[2252]), .Z(n40428) );
  XNOR U49676 ( .A(n40420), .B(n40421), .Z(n40431) );
  XNOR U49677 ( .A(y[2247]), .B(x[2247]), .Z(n40421) );
  XNOR U49678 ( .A(n40422), .B(n40423), .Z(n40420) );
  XNOR U49679 ( .A(y[2248]), .B(x[2248]), .Z(n40423) );
  XNOR U49680 ( .A(y[2249]), .B(x[2249]), .Z(n40422) );
  NAND U49681 ( .A(n40487), .B(n40488), .Z(N61805) );
  NANDN U49682 ( .A(n40489), .B(n40490), .Z(n40488) );
  OR U49683 ( .A(n40491), .B(n40492), .Z(n40490) );
  NAND U49684 ( .A(n40491), .B(n40492), .Z(n40487) );
  XOR U49685 ( .A(n40491), .B(n40493), .Z(N61804) );
  XNOR U49686 ( .A(n40489), .B(n40492), .Z(n40493) );
  AND U49687 ( .A(n40494), .B(n40495), .Z(n40492) );
  NANDN U49688 ( .A(n40496), .B(n40497), .Z(n40495) );
  NANDN U49689 ( .A(n40498), .B(n40499), .Z(n40497) );
  NANDN U49690 ( .A(n40499), .B(n40498), .Z(n40494) );
  NAND U49691 ( .A(n40500), .B(n40501), .Z(n40489) );
  NANDN U49692 ( .A(n40502), .B(n40503), .Z(n40501) );
  OR U49693 ( .A(n40504), .B(n40505), .Z(n40503) );
  NAND U49694 ( .A(n40505), .B(n40504), .Z(n40500) );
  AND U49695 ( .A(n40506), .B(n40507), .Z(n40491) );
  NANDN U49696 ( .A(n40508), .B(n40509), .Z(n40507) );
  NANDN U49697 ( .A(n40510), .B(n40511), .Z(n40509) );
  NANDN U49698 ( .A(n40511), .B(n40510), .Z(n40506) );
  XOR U49699 ( .A(n40505), .B(n40512), .Z(N61803) );
  XOR U49700 ( .A(n40502), .B(n40504), .Z(n40512) );
  XNOR U49701 ( .A(n40498), .B(n40513), .Z(n40504) );
  XNOR U49702 ( .A(n40496), .B(n40499), .Z(n40513) );
  NAND U49703 ( .A(n40514), .B(n40515), .Z(n40499) );
  NAND U49704 ( .A(n40516), .B(n40517), .Z(n40515) );
  OR U49705 ( .A(n40518), .B(n40519), .Z(n40516) );
  NANDN U49706 ( .A(n40520), .B(n40518), .Z(n40514) );
  IV U49707 ( .A(n40519), .Z(n40520) );
  NAND U49708 ( .A(n40521), .B(n40522), .Z(n40496) );
  NAND U49709 ( .A(n40523), .B(n40524), .Z(n40522) );
  NANDN U49710 ( .A(n40525), .B(n40526), .Z(n40523) );
  NANDN U49711 ( .A(n40526), .B(n40525), .Z(n40521) );
  AND U49712 ( .A(n40527), .B(n40528), .Z(n40498) );
  NAND U49713 ( .A(n40529), .B(n40530), .Z(n40528) );
  OR U49714 ( .A(n40531), .B(n40532), .Z(n40529) );
  NANDN U49715 ( .A(n40533), .B(n40531), .Z(n40527) );
  NAND U49716 ( .A(n40534), .B(n40535), .Z(n40502) );
  NANDN U49717 ( .A(n40536), .B(n40537), .Z(n40535) );
  OR U49718 ( .A(n40538), .B(n40539), .Z(n40537) );
  NANDN U49719 ( .A(n40540), .B(n40538), .Z(n40534) );
  IV U49720 ( .A(n40539), .Z(n40540) );
  XNOR U49721 ( .A(n40510), .B(n40541), .Z(n40505) );
  XNOR U49722 ( .A(n40508), .B(n40511), .Z(n40541) );
  NAND U49723 ( .A(n40542), .B(n40543), .Z(n40511) );
  NAND U49724 ( .A(n40544), .B(n40545), .Z(n40543) );
  OR U49725 ( .A(n40546), .B(n40547), .Z(n40544) );
  NANDN U49726 ( .A(n40548), .B(n40546), .Z(n40542) );
  IV U49727 ( .A(n40547), .Z(n40548) );
  NAND U49728 ( .A(n40549), .B(n40550), .Z(n40508) );
  NAND U49729 ( .A(n40551), .B(n40552), .Z(n40550) );
  NANDN U49730 ( .A(n40553), .B(n40554), .Z(n40551) );
  NANDN U49731 ( .A(n40554), .B(n40553), .Z(n40549) );
  AND U49732 ( .A(n40555), .B(n40556), .Z(n40510) );
  NAND U49733 ( .A(n40557), .B(n40558), .Z(n40556) );
  OR U49734 ( .A(n40559), .B(n40560), .Z(n40557) );
  NANDN U49735 ( .A(n40561), .B(n40559), .Z(n40555) );
  XNOR U49736 ( .A(n40536), .B(n40562), .Z(N61802) );
  XOR U49737 ( .A(n40538), .B(n40539), .Z(n40562) );
  XNOR U49738 ( .A(n40552), .B(n40563), .Z(n40539) );
  XOR U49739 ( .A(n40553), .B(n40554), .Z(n40563) );
  XOR U49740 ( .A(n40559), .B(n40564), .Z(n40554) );
  XOR U49741 ( .A(n40558), .B(n40561), .Z(n40564) );
  IV U49742 ( .A(n40560), .Z(n40561) );
  NAND U49743 ( .A(n40565), .B(n40566), .Z(n40560) );
  OR U49744 ( .A(n40567), .B(n40568), .Z(n40566) );
  OR U49745 ( .A(n40569), .B(n40570), .Z(n40565) );
  NAND U49746 ( .A(n40571), .B(n40572), .Z(n40558) );
  OR U49747 ( .A(n40573), .B(n40574), .Z(n40572) );
  OR U49748 ( .A(n40575), .B(n40576), .Z(n40571) );
  NOR U49749 ( .A(n40577), .B(n40578), .Z(n40559) );
  ANDN U49750 ( .B(n40579), .A(n40580), .Z(n40553) );
  XNOR U49751 ( .A(n40546), .B(n40581), .Z(n40552) );
  XNOR U49752 ( .A(n40545), .B(n40547), .Z(n40581) );
  NAND U49753 ( .A(n40582), .B(n40583), .Z(n40547) );
  OR U49754 ( .A(n40584), .B(n40585), .Z(n40583) );
  OR U49755 ( .A(n40586), .B(n40587), .Z(n40582) );
  NAND U49756 ( .A(n40588), .B(n40589), .Z(n40545) );
  OR U49757 ( .A(n40590), .B(n40591), .Z(n40589) );
  OR U49758 ( .A(n40592), .B(n40593), .Z(n40588) );
  ANDN U49759 ( .B(n40594), .A(n40595), .Z(n40546) );
  IV U49760 ( .A(n40596), .Z(n40594) );
  ANDN U49761 ( .B(n40597), .A(n40598), .Z(n40538) );
  XOR U49762 ( .A(n40524), .B(n40599), .Z(n40536) );
  XOR U49763 ( .A(n40525), .B(n40526), .Z(n40599) );
  XOR U49764 ( .A(n40531), .B(n40600), .Z(n40526) );
  XOR U49765 ( .A(n40530), .B(n40533), .Z(n40600) );
  IV U49766 ( .A(n40532), .Z(n40533) );
  NAND U49767 ( .A(n40601), .B(n40602), .Z(n40532) );
  OR U49768 ( .A(n40603), .B(n40604), .Z(n40602) );
  OR U49769 ( .A(n40605), .B(n40606), .Z(n40601) );
  NAND U49770 ( .A(n40607), .B(n40608), .Z(n40530) );
  OR U49771 ( .A(n40609), .B(n40610), .Z(n40608) );
  OR U49772 ( .A(n40611), .B(n40612), .Z(n40607) );
  NOR U49773 ( .A(n40613), .B(n40614), .Z(n40531) );
  ANDN U49774 ( .B(n40615), .A(n40616), .Z(n40525) );
  IV U49775 ( .A(n40617), .Z(n40615) );
  XNOR U49776 ( .A(n40518), .B(n40618), .Z(n40524) );
  XNOR U49777 ( .A(n40517), .B(n40519), .Z(n40618) );
  NAND U49778 ( .A(n40619), .B(n40620), .Z(n40519) );
  OR U49779 ( .A(n40621), .B(n40622), .Z(n40620) );
  OR U49780 ( .A(n40623), .B(n40624), .Z(n40619) );
  NAND U49781 ( .A(n40625), .B(n40626), .Z(n40517) );
  OR U49782 ( .A(n40627), .B(n40628), .Z(n40626) );
  OR U49783 ( .A(n40629), .B(n40630), .Z(n40625) );
  ANDN U49784 ( .B(n40631), .A(n40632), .Z(n40518) );
  IV U49785 ( .A(n40633), .Z(n40631) );
  XNOR U49786 ( .A(n40598), .B(n40597), .Z(N61801) );
  XOR U49787 ( .A(n40617), .B(n40616), .Z(n40597) );
  XNOR U49788 ( .A(n40632), .B(n40633), .Z(n40616) );
  XNOR U49789 ( .A(n40627), .B(n40628), .Z(n40633) );
  XNOR U49790 ( .A(n40629), .B(n40630), .Z(n40628) );
  XNOR U49791 ( .A(y[2245]), .B(x[2245]), .Z(n40630) );
  XNOR U49792 ( .A(y[2246]), .B(x[2246]), .Z(n40629) );
  XNOR U49793 ( .A(y[2244]), .B(x[2244]), .Z(n40627) );
  XNOR U49794 ( .A(n40621), .B(n40622), .Z(n40632) );
  XNOR U49795 ( .A(y[2241]), .B(x[2241]), .Z(n40622) );
  XNOR U49796 ( .A(n40623), .B(n40624), .Z(n40621) );
  XNOR U49797 ( .A(y[2242]), .B(x[2242]), .Z(n40624) );
  XNOR U49798 ( .A(y[2243]), .B(x[2243]), .Z(n40623) );
  XNOR U49799 ( .A(n40614), .B(n40613), .Z(n40617) );
  XNOR U49800 ( .A(n40609), .B(n40610), .Z(n40613) );
  XNOR U49801 ( .A(y[2238]), .B(x[2238]), .Z(n40610) );
  XNOR U49802 ( .A(n40611), .B(n40612), .Z(n40609) );
  XNOR U49803 ( .A(y[2239]), .B(x[2239]), .Z(n40612) );
  XNOR U49804 ( .A(y[2240]), .B(x[2240]), .Z(n40611) );
  XNOR U49805 ( .A(n40603), .B(n40604), .Z(n40614) );
  XNOR U49806 ( .A(y[2235]), .B(x[2235]), .Z(n40604) );
  XNOR U49807 ( .A(n40605), .B(n40606), .Z(n40603) );
  XNOR U49808 ( .A(y[2236]), .B(x[2236]), .Z(n40606) );
  XNOR U49809 ( .A(y[2237]), .B(x[2237]), .Z(n40605) );
  XOR U49810 ( .A(n40579), .B(n40580), .Z(n40598) );
  XNOR U49811 ( .A(n40595), .B(n40596), .Z(n40580) );
  XNOR U49812 ( .A(n40590), .B(n40591), .Z(n40596) );
  XNOR U49813 ( .A(n40592), .B(n40593), .Z(n40591) );
  XNOR U49814 ( .A(y[2233]), .B(x[2233]), .Z(n40593) );
  XNOR U49815 ( .A(y[2234]), .B(x[2234]), .Z(n40592) );
  XNOR U49816 ( .A(y[2232]), .B(x[2232]), .Z(n40590) );
  XNOR U49817 ( .A(n40584), .B(n40585), .Z(n40595) );
  XNOR U49818 ( .A(y[2229]), .B(x[2229]), .Z(n40585) );
  XNOR U49819 ( .A(n40586), .B(n40587), .Z(n40584) );
  XNOR U49820 ( .A(y[2230]), .B(x[2230]), .Z(n40587) );
  XNOR U49821 ( .A(y[2231]), .B(x[2231]), .Z(n40586) );
  XOR U49822 ( .A(n40578), .B(n40577), .Z(n40579) );
  XNOR U49823 ( .A(n40573), .B(n40574), .Z(n40577) );
  XNOR U49824 ( .A(y[2226]), .B(x[2226]), .Z(n40574) );
  XNOR U49825 ( .A(n40575), .B(n40576), .Z(n40573) );
  XNOR U49826 ( .A(y[2227]), .B(x[2227]), .Z(n40576) );
  XNOR U49827 ( .A(y[2228]), .B(x[2228]), .Z(n40575) );
  XNOR U49828 ( .A(n40567), .B(n40568), .Z(n40578) );
  XNOR U49829 ( .A(y[2223]), .B(x[2223]), .Z(n40568) );
  XNOR U49830 ( .A(n40569), .B(n40570), .Z(n40567) );
  XNOR U49831 ( .A(y[2224]), .B(x[2224]), .Z(n40570) );
  XNOR U49832 ( .A(y[2225]), .B(x[2225]), .Z(n40569) );
  NAND U49833 ( .A(n40634), .B(n40635), .Z(N61792) );
  NANDN U49834 ( .A(n40636), .B(n40637), .Z(n40635) );
  OR U49835 ( .A(n40638), .B(n40639), .Z(n40637) );
  NAND U49836 ( .A(n40638), .B(n40639), .Z(n40634) );
  XOR U49837 ( .A(n40638), .B(n40640), .Z(N61791) );
  XNOR U49838 ( .A(n40636), .B(n40639), .Z(n40640) );
  AND U49839 ( .A(n40641), .B(n40642), .Z(n40639) );
  NANDN U49840 ( .A(n40643), .B(n40644), .Z(n40642) );
  NANDN U49841 ( .A(n40645), .B(n40646), .Z(n40644) );
  NANDN U49842 ( .A(n40646), .B(n40645), .Z(n40641) );
  NAND U49843 ( .A(n40647), .B(n40648), .Z(n40636) );
  NANDN U49844 ( .A(n40649), .B(n40650), .Z(n40648) );
  OR U49845 ( .A(n40651), .B(n40652), .Z(n40650) );
  NAND U49846 ( .A(n40652), .B(n40651), .Z(n40647) );
  AND U49847 ( .A(n40653), .B(n40654), .Z(n40638) );
  NANDN U49848 ( .A(n40655), .B(n40656), .Z(n40654) );
  NANDN U49849 ( .A(n40657), .B(n40658), .Z(n40656) );
  NANDN U49850 ( .A(n40658), .B(n40657), .Z(n40653) );
  XOR U49851 ( .A(n40652), .B(n40659), .Z(N61790) );
  XOR U49852 ( .A(n40649), .B(n40651), .Z(n40659) );
  XNOR U49853 ( .A(n40645), .B(n40660), .Z(n40651) );
  XNOR U49854 ( .A(n40643), .B(n40646), .Z(n40660) );
  NAND U49855 ( .A(n40661), .B(n40662), .Z(n40646) );
  NAND U49856 ( .A(n40663), .B(n40664), .Z(n40662) );
  OR U49857 ( .A(n40665), .B(n40666), .Z(n40663) );
  NANDN U49858 ( .A(n40667), .B(n40665), .Z(n40661) );
  IV U49859 ( .A(n40666), .Z(n40667) );
  NAND U49860 ( .A(n40668), .B(n40669), .Z(n40643) );
  NAND U49861 ( .A(n40670), .B(n40671), .Z(n40669) );
  NANDN U49862 ( .A(n40672), .B(n40673), .Z(n40670) );
  NANDN U49863 ( .A(n40673), .B(n40672), .Z(n40668) );
  AND U49864 ( .A(n40674), .B(n40675), .Z(n40645) );
  NAND U49865 ( .A(n40676), .B(n40677), .Z(n40675) );
  OR U49866 ( .A(n40678), .B(n40679), .Z(n40676) );
  NANDN U49867 ( .A(n40680), .B(n40678), .Z(n40674) );
  NAND U49868 ( .A(n40681), .B(n40682), .Z(n40649) );
  NANDN U49869 ( .A(n40683), .B(n40684), .Z(n40682) );
  OR U49870 ( .A(n40685), .B(n40686), .Z(n40684) );
  NANDN U49871 ( .A(n40687), .B(n40685), .Z(n40681) );
  IV U49872 ( .A(n40686), .Z(n40687) );
  XNOR U49873 ( .A(n40657), .B(n40688), .Z(n40652) );
  XNOR U49874 ( .A(n40655), .B(n40658), .Z(n40688) );
  NAND U49875 ( .A(n40689), .B(n40690), .Z(n40658) );
  NAND U49876 ( .A(n40691), .B(n40692), .Z(n40690) );
  OR U49877 ( .A(n40693), .B(n40694), .Z(n40691) );
  NANDN U49878 ( .A(n40695), .B(n40693), .Z(n40689) );
  IV U49879 ( .A(n40694), .Z(n40695) );
  NAND U49880 ( .A(n40696), .B(n40697), .Z(n40655) );
  NAND U49881 ( .A(n40698), .B(n40699), .Z(n40697) );
  NANDN U49882 ( .A(n40700), .B(n40701), .Z(n40698) );
  NANDN U49883 ( .A(n40701), .B(n40700), .Z(n40696) );
  AND U49884 ( .A(n40702), .B(n40703), .Z(n40657) );
  NAND U49885 ( .A(n40704), .B(n40705), .Z(n40703) );
  OR U49886 ( .A(n40706), .B(n40707), .Z(n40704) );
  NANDN U49887 ( .A(n40708), .B(n40706), .Z(n40702) );
  XNOR U49888 ( .A(n40683), .B(n40709), .Z(N61789) );
  XOR U49889 ( .A(n40685), .B(n40686), .Z(n40709) );
  XNOR U49890 ( .A(n40699), .B(n40710), .Z(n40686) );
  XOR U49891 ( .A(n40700), .B(n40701), .Z(n40710) );
  XOR U49892 ( .A(n40706), .B(n40711), .Z(n40701) );
  XOR U49893 ( .A(n40705), .B(n40708), .Z(n40711) );
  IV U49894 ( .A(n40707), .Z(n40708) );
  NAND U49895 ( .A(n40712), .B(n40713), .Z(n40707) );
  OR U49896 ( .A(n40714), .B(n40715), .Z(n40713) );
  OR U49897 ( .A(n40716), .B(n40717), .Z(n40712) );
  NAND U49898 ( .A(n40718), .B(n40719), .Z(n40705) );
  OR U49899 ( .A(n40720), .B(n40721), .Z(n40719) );
  OR U49900 ( .A(n40722), .B(n40723), .Z(n40718) );
  NOR U49901 ( .A(n40724), .B(n40725), .Z(n40706) );
  ANDN U49902 ( .B(n40726), .A(n40727), .Z(n40700) );
  XNOR U49903 ( .A(n40693), .B(n40728), .Z(n40699) );
  XNOR U49904 ( .A(n40692), .B(n40694), .Z(n40728) );
  NAND U49905 ( .A(n40729), .B(n40730), .Z(n40694) );
  OR U49906 ( .A(n40731), .B(n40732), .Z(n40730) );
  OR U49907 ( .A(n40733), .B(n40734), .Z(n40729) );
  NAND U49908 ( .A(n40735), .B(n40736), .Z(n40692) );
  OR U49909 ( .A(n40737), .B(n40738), .Z(n40736) );
  OR U49910 ( .A(n40739), .B(n40740), .Z(n40735) );
  ANDN U49911 ( .B(n40741), .A(n40742), .Z(n40693) );
  IV U49912 ( .A(n40743), .Z(n40741) );
  ANDN U49913 ( .B(n40744), .A(n40745), .Z(n40685) );
  XOR U49914 ( .A(n40671), .B(n40746), .Z(n40683) );
  XOR U49915 ( .A(n40672), .B(n40673), .Z(n40746) );
  XOR U49916 ( .A(n40678), .B(n40747), .Z(n40673) );
  XOR U49917 ( .A(n40677), .B(n40680), .Z(n40747) );
  IV U49918 ( .A(n40679), .Z(n40680) );
  NAND U49919 ( .A(n40748), .B(n40749), .Z(n40679) );
  OR U49920 ( .A(n40750), .B(n40751), .Z(n40749) );
  OR U49921 ( .A(n40752), .B(n40753), .Z(n40748) );
  NAND U49922 ( .A(n40754), .B(n40755), .Z(n40677) );
  OR U49923 ( .A(n40756), .B(n40757), .Z(n40755) );
  OR U49924 ( .A(n40758), .B(n40759), .Z(n40754) );
  NOR U49925 ( .A(n40760), .B(n40761), .Z(n40678) );
  ANDN U49926 ( .B(n40762), .A(n40763), .Z(n40672) );
  IV U49927 ( .A(n40764), .Z(n40762) );
  XNOR U49928 ( .A(n40665), .B(n40765), .Z(n40671) );
  XNOR U49929 ( .A(n40664), .B(n40666), .Z(n40765) );
  NAND U49930 ( .A(n40766), .B(n40767), .Z(n40666) );
  OR U49931 ( .A(n40768), .B(n40769), .Z(n40767) );
  OR U49932 ( .A(n40770), .B(n40771), .Z(n40766) );
  NAND U49933 ( .A(n40772), .B(n40773), .Z(n40664) );
  OR U49934 ( .A(n40774), .B(n40775), .Z(n40773) );
  OR U49935 ( .A(n40776), .B(n40777), .Z(n40772) );
  ANDN U49936 ( .B(n40778), .A(n40779), .Z(n40665) );
  IV U49937 ( .A(n40780), .Z(n40778) );
  XNOR U49938 ( .A(n40745), .B(n40744), .Z(N61788) );
  XOR U49939 ( .A(n40764), .B(n40763), .Z(n40744) );
  XNOR U49940 ( .A(n40779), .B(n40780), .Z(n40763) );
  XNOR U49941 ( .A(n40774), .B(n40775), .Z(n40780) );
  XNOR U49942 ( .A(n40776), .B(n40777), .Z(n40775) );
  XNOR U49943 ( .A(y[2221]), .B(x[2221]), .Z(n40777) );
  XNOR U49944 ( .A(y[2222]), .B(x[2222]), .Z(n40776) );
  XNOR U49945 ( .A(y[2220]), .B(x[2220]), .Z(n40774) );
  XNOR U49946 ( .A(n40768), .B(n40769), .Z(n40779) );
  XNOR U49947 ( .A(y[2217]), .B(x[2217]), .Z(n40769) );
  XNOR U49948 ( .A(n40770), .B(n40771), .Z(n40768) );
  XNOR U49949 ( .A(y[2218]), .B(x[2218]), .Z(n40771) );
  XNOR U49950 ( .A(y[2219]), .B(x[2219]), .Z(n40770) );
  XNOR U49951 ( .A(n40761), .B(n40760), .Z(n40764) );
  XNOR U49952 ( .A(n40756), .B(n40757), .Z(n40760) );
  XNOR U49953 ( .A(y[2214]), .B(x[2214]), .Z(n40757) );
  XNOR U49954 ( .A(n40758), .B(n40759), .Z(n40756) );
  XNOR U49955 ( .A(y[2215]), .B(x[2215]), .Z(n40759) );
  XNOR U49956 ( .A(y[2216]), .B(x[2216]), .Z(n40758) );
  XNOR U49957 ( .A(n40750), .B(n40751), .Z(n40761) );
  XNOR U49958 ( .A(y[2211]), .B(x[2211]), .Z(n40751) );
  XNOR U49959 ( .A(n40752), .B(n40753), .Z(n40750) );
  XNOR U49960 ( .A(y[2212]), .B(x[2212]), .Z(n40753) );
  XNOR U49961 ( .A(y[2213]), .B(x[2213]), .Z(n40752) );
  XOR U49962 ( .A(n40726), .B(n40727), .Z(n40745) );
  XNOR U49963 ( .A(n40742), .B(n40743), .Z(n40727) );
  XNOR U49964 ( .A(n40737), .B(n40738), .Z(n40743) );
  XNOR U49965 ( .A(n40739), .B(n40740), .Z(n40738) );
  XNOR U49966 ( .A(y[2209]), .B(x[2209]), .Z(n40740) );
  XNOR U49967 ( .A(y[2210]), .B(x[2210]), .Z(n40739) );
  XNOR U49968 ( .A(y[2208]), .B(x[2208]), .Z(n40737) );
  XNOR U49969 ( .A(n40731), .B(n40732), .Z(n40742) );
  XNOR U49970 ( .A(y[2205]), .B(x[2205]), .Z(n40732) );
  XNOR U49971 ( .A(n40733), .B(n40734), .Z(n40731) );
  XNOR U49972 ( .A(y[2206]), .B(x[2206]), .Z(n40734) );
  XNOR U49973 ( .A(y[2207]), .B(x[2207]), .Z(n40733) );
  XOR U49974 ( .A(n40725), .B(n40724), .Z(n40726) );
  XNOR U49975 ( .A(n40720), .B(n40721), .Z(n40724) );
  XNOR U49976 ( .A(y[2202]), .B(x[2202]), .Z(n40721) );
  XNOR U49977 ( .A(n40722), .B(n40723), .Z(n40720) );
  XNOR U49978 ( .A(y[2203]), .B(x[2203]), .Z(n40723) );
  XNOR U49979 ( .A(y[2204]), .B(x[2204]), .Z(n40722) );
  XNOR U49980 ( .A(n40714), .B(n40715), .Z(n40725) );
  XNOR U49981 ( .A(y[2199]), .B(x[2199]), .Z(n40715) );
  XNOR U49982 ( .A(n40716), .B(n40717), .Z(n40714) );
  XNOR U49983 ( .A(y[2200]), .B(x[2200]), .Z(n40717) );
  XNOR U49984 ( .A(y[2201]), .B(x[2201]), .Z(n40716) );
  NAND U49985 ( .A(n40781), .B(n40782), .Z(N61779) );
  NANDN U49986 ( .A(n40783), .B(n40784), .Z(n40782) );
  OR U49987 ( .A(n40785), .B(n40786), .Z(n40784) );
  NAND U49988 ( .A(n40785), .B(n40786), .Z(n40781) );
  XOR U49989 ( .A(n40785), .B(n40787), .Z(N61778) );
  XNOR U49990 ( .A(n40783), .B(n40786), .Z(n40787) );
  AND U49991 ( .A(n40788), .B(n40789), .Z(n40786) );
  NANDN U49992 ( .A(n40790), .B(n40791), .Z(n40789) );
  NANDN U49993 ( .A(n40792), .B(n40793), .Z(n40791) );
  NANDN U49994 ( .A(n40793), .B(n40792), .Z(n40788) );
  NAND U49995 ( .A(n40794), .B(n40795), .Z(n40783) );
  NANDN U49996 ( .A(n40796), .B(n40797), .Z(n40795) );
  OR U49997 ( .A(n40798), .B(n40799), .Z(n40797) );
  NAND U49998 ( .A(n40799), .B(n40798), .Z(n40794) );
  AND U49999 ( .A(n40800), .B(n40801), .Z(n40785) );
  NANDN U50000 ( .A(n40802), .B(n40803), .Z(n40801) );
  NANDN U50001 ( .A(n40804), .B(n40805), .Z(n40803) );
  NANDN U50002 ( .A(n40805), .B(n40804), .Z(n40800) );
  XOR U50003 ( .A(n40799), .B(n40806), .Z(N61777) );
  XOR U50004 ( .A(n40796), .B(n40798), .Z(n40806) );
  XNOR U50005 ( .A(n40792), .B(n40807), .Z(n40798) );
  XNOR U50006 ( .A(n40790), .B(n40793), .Z(n40807) );
  NAND U50007 ( .A(n40808), .B(n40809), .Z(n40793) );
  NAND U50008 ( .A(n40810), .B(n40811), .Z(n40809) );
  OR U50009 ( .A(n40812), .B(n40813), .Z(n40810) );
  NANDN U50010 ( .A(n40814), .B(n40812), .Z(n40808) );
  IV U50011 ( .A(n40813), .Z(n40814) );
  NAND U50012 ( .A(n40815), .B(n40816), .Z(n40790) );
  NAND U50013 ( .A(n40817), .B(n40818), .Z(n40816) );
  NANDN U50014 ( .A(n40819), .B(n40820), .Z(n40817) );
  NANDN U50015 ( .A(n40820), .B(n40819), .Z(n40815) );
  AND U50016 ( .A(n40821), .B(n40822), .Z(n40792) );
  NAND U50017 ( .A(n40823), .B(n40824), .Z(n40822) );
  OR U50018 ( .A(n40825), .B(n40826), .Z(n40823) );
  NANDN U50019 ( .A(n40827), .B(n40825), .Z(n40821) );
  NAND U50020 ( .A(n40828), .B(n40829), .Z(n40796) );
  NANDN U50021 ( .A(n40830), .B(n40831), .Z(n40829) );
  OR U50022 ( .A(n40832), .B(n40833), .Z(n40831) );
  NANDN U50023 ( .A(n40834), .B(n40832), .Z(n40828) );
  IV U50024 ( .A(n40833), .Z(n40834) );
  XNOR U50025 ( .A(n40804), .B(n40835), .Z(n40799) );
  XNOR U50026 ( .A(n40802), .B(n40805), .Z(n40835) );
  NAND U50027 ( .A(n40836), .B(n40837), .Z(n40805) );
  NAND U50028 ( .A(n40838), .B(n40839), .Z(n40837) );
  OR U50029 ( .A(n40840), .B(n40841), .Z(n40838) );
  NANDN U50030 ( .A(n40842), .B(n40840), .Z(n40836) );
  IV U50031 ( .A(n40841), .Z(n40842) );
  NAND U50032 ( .A(n40843), .B(n40844), .Z(n40802) );
  NAND U50033 ( .A(n40845), .B(n40846), .Z(n40844) );
  NANDN U50034 ( .A(n40847), .B(n40848), .Z(n40845) );
  NANDN U50035 ( .A(n40848), .B(n40847), .Z(n40843) );
  AND U50036 ( .A(n40849), .B(n40850), .Z(n40804) );
  NAND U50037 ( .A(n40851), .B(n40852), .Z(n40850) );
  OR U50038 ( .A(n40853), .B(n40854), .Z(n40851) );
  NANDN U50039 ( .A(n40855), .B(n40853), .Z(n40849) );
  XNOR U50040 ( .A(n40830), .B(n40856), .Z(N61776) );
  XOR U50041 ( .A(n40832), .B(n40833), .Z(n40856) );
  XNOR U50042 ( .A(n40846), .B(n40857), .Z(n40833) );
  XOR U50043 ( .A(n40847), .B(n40848), .Z(n40857) );
  XOR U50044 ( .A(n40853), .B(n40858), .Z(n40848) );
  XOR U50045 ( .A(n40852), .B(n40855), .Z(n40858) );
  IV U50046 ( .A(n40854), .Z(n40855) );
  NAND U50047 ( .A(n40859), .B(n40860), .Z(n40854) );
  OR U50048 ( .A(n40861), .B(n40862), .Z(n40860) );
  OR U50049 ( .A(n40863), .B(n40864), .Z(n40859) );
  NAND U50050 ( .A(n40865), .B(n40866), .Z(n40852) );
  OR U50051 ( .A(n40867), .B(n40868), .Z(n40866) );
  OR U50052 ( .A(n40869), .B(n40870), .Z(n40865) );
  NOR U50053 ( .A(n40871), .B(n40872), .Z(n40853) );
  ANDN U50054 ( .B(n40873), .A(n40874), .Z(n40847) );
  XNOR U50055 ( .A(n40840), .B(n40875), .Z(n40846) );
  XNOR U50056 ( .A(n40839), .B(n40841), .Z(n40875) );
  NAND U50057 ( .A(n40876), .B(n40877), .Z(n40841) );
  OR U50058 ( .A(n40878), .B(n40879), .Z(n40877) );
  OR U50059 ( .A(n40880), .B(n40881), .Z(n40876) );
  NAND U50060 ( .A(n40882), .B(n40883), .Z(n40839) );
  OR U50061 ( .A(n40884), .B(n40885), .Z(n40883) );
  OR U50062 ( .A(n40886), .B(n40887), .Z(n40882) );
  ANDN U50063 ( .B(n40888), .A(n40889), .Z(n40840) );
  IV U50064 ( .A(n40890), .Z(n40888) );
  ANDN U50065 ( .B(n40891), .A(n40892), .Z(n40832) );
  XOR U50066 ( .A(n40818), .B(n40893), .Z(n40830) );
  XOR U50067 ( .A(n40819), .B(n40820), .Z(n40893) );
  XOR U50068 ( .A(n40825), .B(n40894), .Z(n40820) );
  XOR U50069 ( .A(n40824), .B(n40827), .Z(n40894) );
  IV U50070 ( .A(n40826), .Z(n40827) );
  NAND U50071 ( .A(n40895), .B(n40896), .Z(n40826) );
  OR U50072 ( .A(n40897), .B(n40898), .Z(n40896) );
  OR U50073 ( .A(n40899), .B(n40900), .Z(n40895) );
  NAND U50074 ( .A(n40901), .B(n40902), .Z(n40824) );
  OR U50075 ( .A(n40903), .B(n40904), .Z(n40902) );
  OR U50076 ( .A(n40905), .B(n40906), .Z(n40901) );
  NOR U50077 ( .A(n40907), .B(n40908), .Z(n40825) );
  ANDN U50078 ( .B(n40909), .A(n40910), .Z(n40819) );
  IV U50079 ( .A(n40911), .Z(n40909) );
  XNOR U50080 ( .A(n40812), .B(n40912), .Z(n40818) );
  XNOR U50081 ( .A(n40811), .B(n40813), .Z(n40912) );
  NAND U50082 ( .A(n40913), .B(n40914), .Z(n40813) );
  OR U50083 ( .A(n40915), .B(n40916), .Z(n40914) );
  OR U50084 ( .A(n40917), .B(n40918), .Z(n40913) );
  NAND U50085 ( .A(n40919), .B(n40920), .Z(n40811) );
  OR U50086 ( .A(n40921), .B(n40922), .Z(n40920) );
  OR U50087 ( .A(n40923), .B(n40924), .Z(n40919) );
  ANDN U50088 ( .B(n40925), .A(n40926), .Z(n40812) );
  IV U50089 ( .A(n40927), .Z(n40925) );
  XNOR U50090 ( .A(n40892), .B(n40891), .Z(N61775) );
  XOR U50091 ( .A(n40911), .B(n40910), .Z(n40891) );
  XNOR U50092 ( .A(n40926), .B(n40927), .Z(n40910) );
  XNOR U50093 ( .A(n40921), .B(n40922), .Z(n40927) );
  XNOR U50094 ( .A(n40923), .B(n40924), .Z(n40922) );
  XNOR U50095 ( .A(y[2197]), .B(x[2197]), .Z(n40924) );
  XNOR U50096 ( .A(y[2198]), .B(x[2198]), .Z(n40923) );
  XNOR U50097 ( .A(y[2196]), .B(x[2196]), .Z(n40921) );
  XNOR U50098 ( .A(n40915), .B(n40916), .Z(n40926) );
  XNOR U50099 ( .A(y[2193]), .B(x[2193]), .Z(n40916) );
  XNOR U50100 ( .A(n40917), .B(n40918), .Z(n40915) );
  XNOR U50101 ( .A(y[2194]), .B(x[2194]), .Z(n40918) );
  XNOR U50102 ( .A(y[2195]), .B(x[2195]), .Z(n40917) );
  XNOR U50103 ( .A(n40908), .B(n40907), .Z(n40911) );
  XNOR U50104 ( .A(n40903), .B(n40904), .Z(n40907) );
  XNOR U50105 ( .A(y[2190]), .B(x[2190]), .Z(n40904) );
  XNOR U50106 ( .A(n40905), .B(n40906), .Z(n40903) );
  XNOR U50107 ( .A(y[2191]), .B(x[2191]), .Z(n40906) );
  XNOR U50108 ( .A(y[2192]), .B(x[2192]), .Z(n40905) );
  XNOR U50109 ( .A(n40897), .B(n40898), .Z(n40908) );
  XNOR U50110 ( .A(y[2187]), .B(x[2187]), .Z(n40898) );
  XNOR U50111 ( .A(n40899), .B(n40900), .Z(n40897) );
  XNOR U50112 ( .A(y[2188]), .B(x[2188]), .Z(n40900) );
  XNOR U50113 ( .A(y[2189]), .B(x[2189]), .Z(n40899) );
  XOR U50114 ( .A(n40873), .B(n40874), .Z(n40892) );
  XNOR U50115 ( .A(n40889), .B(n40890), .Z(n40874) );
  XNOR U50116 ( .A(n40884), .B(n40885), .Z(n40890) );
  XNOR U50117 ( .A(n40886), .B(n40887), .Z(n40885) );
  XNOR U50118 ( .A(y[2185]), .B(x[2185]), .Z(n40887) );
  XNOR U50119 ( .A(y[2186]), .B(x[2186]), .Z(n40886) );
  XNOR U50120 ( .A(y[2184]), .B(x[2184]), .Z(n40884) );
  XNOR U50121 ( .A(n40878), .B(n40879), .Z(n40889) );
  XNOR U50122 ( .A(y[2181]), .B(x[2181]), .Z(n40879) );
  XNOR U50123 ( .A(n40880), .B(n40881), .Z(n40878) );
  XNOR U50124 ( .A(y[2182]), .B(x[2182]), .Z(n40881) );
  XNOR U50125 ( .A(y[2183]), .B(x[2183]), .Z(n40880) );
  XOR U50126 ( .A(n40872), .B(n40871), .Z(n40873) );
  XNOR U50127 ( .A(n40867), .B(n40868), .Z(n40871) );
  XNOR U50128 ( .A(y[2178]), .B(x[2178]), .Z(n40868) );
  XNOR U50129 ( .A(n40869), .B(n40870), .Z(n40867) );
  XNOR U50130 ( .A(y[2179]), .B(x[2179]), .Z(n40870) );
  XNOR U50131 ( .A(y[2180]), .B(x[2180]), .Z(n40869) );
  XNOR U50132 ( .A(n40861), .B(n40862), .Z(n40872) );
  XNOR U50133 ( .A(y[2175]), .B(x[2175]), .Z(n40862) );
  XNOR U50134 ( .A(n40863), .B(n40864), .Z(n40861) );
  XNOR U50135 ( .A(y[2176]), .B(x[2176]), .Z(n40864) );
  XNOR U50136 ( .A(y[2177]), .B(x[2177]), .Z(n40863) );
  NAND U50137 ( .A(n40928), .B(n40929), .Z(N61766) );
  NANDN U50138 ( .A(n40930), .B(n40931), .Z(n40929) );
  OR U50139 ( .A(n40932), .B(n40933), .Z(n40931) );
  NAND U50140 ( .A(n40932), .B(n40933), .Z(n40928) );
  XOR U50141 ( .A(n40932), .B(n40934), .Z(N61765) );
  XNOR U50142 ( .A(n40930), .B(n40933), .Z(n40934) );
  AND U50143 ( .A(n40935), .B(n40936), .Z(n40933) );
  NANDN U50144 ( .A(n40937), .B(n40938), .Z(n40936) );
  NANDN U50145 ( .A(n40939), .B(n40940), .Z(n40938) );
  NANDN U50146 ( .A(n40940), .B(n40939), .Z(n40935) );
  NAND U50147 ( .A(n40941), .B(n40942), .Z(n40930) );
  NANDN U50148 ( .A(n40943), .B(n40944), .Z(n40942) );
  OR U50149 ( .A(n40945), .B(n40946), .Z(n40944) );
  NAND U50150 ( .A(n40946), .B(n40945), .Z(n40941) );
  AND U50151 ( .A(n40947), .B(n40948), .Z(n40932) );
  NANDN U50152 ( .A(n40949), .B(n40950), .Z(n40948) );
  NANDN U50153 ( .A(n40951), .B(n40952), .Z(n40950) );
  NANDN U50154 ( .A(n40952), .B(n40951), .Z(n40947) );
  XOR U50155 ( .A(n40946), .B(n40953), .Z(N61764) );
  XOR U50156 ( .A(n40943), .B(n40945), .Z(n40953) );
  XNOR U50157 ( .A(n40939), .B(n40954), .Z(n40945) );
  XNOR U50158 ( .A(n40937), .B(n40940), .Z(n40954) );
  NAND U50159 ( .A(n40955), .B(n40956), .Z(n40940) );
  NAND U50160 ( .A(n40957), .B(n40958), .Z(n40956) );
  OR U50161 ( .A(n40959), .B(n40960), .Z(n40957) );
  NANDN U50162 ( .A(n40961), .B(n40959), .Z(n40955) );
  IV U50163 ( .A(n40960), .Z(n40961) );
  NAND U50164 ( .A(n40962), .B(n40963), .Z(n40937) );
  NAND U50165 ( .A(n40964), .B(n40965), .Z(n40963) );
  NANDN U50166 ( .A(n40966), .B(n40967), .Z(n40964) );
  NANDN U50167 ( .A(n40967), .B(n40966), .Z(n40962) );
  AND U50168 ( .A(n40968), .B(n40969), .Z(n40939) );
  NAND U50169 ( .A(n40970), .B(n40971), .Z(n40969) );
  OR U50170 ( .A(n40972), .B(n40973), .Z(n40970) );
  NANDN U50171 ( .A(n40974), .B(n40972), .Z(n40968) );
  NAND U50172 ( .A(n40975), .B(n40976), .Z(n40943) );
  NANDN U50173 ( .A(n40977), .B(n40978), .Z(n40976) );
  OR U50174 ( .A(n40979), .B(n40980), .Z(n40978) );
  NANDN U50175 ( .A(n40981), .B(n40979), .Z(n40975) );
  IV U50176 ( .A(n40980), .Z(n40981) );
  XNOR U50177 ( .A(n40951), .B(n40982), .Z(n40946) );
  XNOR U50178 ( .A(n40949), .B(n40952), .Z(n40982) );
  NAND U50179 ( .A(n40983), .B(n40984), .Z(n40952) );
  NAND U50180 ( .A(n40985), .B(n40986), .Z(n40984) );
  OR U50181 ( .A(n40987), .B(n40988), .Z(n40985) );
  NANDN U50182 ( .A(n40989), .B(n40987), .Z(n40983) );
  IV U50183 ( .A(n40988), .Z(n40989) );
  NAND U50184 ( .A(n40990), .B(n40991), .Z(n40949) );
  NAND U50185 ( .A(n40992), .B(n40993), .Z(n40991) );
  NANDN U50186 ( .A(n40994), .B(n40995), .Z(n40992) );
  NANDN U50187 ( .A(n40995), .B(n40994), .Z(n40990) );
  AND U50188 ( .A(n40996), .B(n40997), .Z(n40951) );
  NAND U50189 ( .A(n40998), .B(n40999), .Z(n40997) );
  OR U50190 ( .A(n41000), .B(n41001), .Z(n40998) );
  NANDN U50191 ( .A(n41002), .B(n41000), .Z(n40996) );
  XNOR U50192 ( .A(n40977), .B(n41003), .Z(N61763) );
  XOR U50193 ( .A(n40979), .B(n40980), .Z(n41003) );
  XNOR U50194 ( .A(n40993), .B(n41004), .Z(n40980) );
  XOR U50195 ( .A(n40994), .B(n40995), .Z(n41004) );
  XOR U50196 ( .A(n41000), .B(n41005), .Z(n40995) );
  XOR U50197 ( .A(n40999), .B(n41002), .Z(n41005) );
  IV U50198 ( .A(n41001), .Z(n41002) );
  NAND U50199 ( .A(n41006), .B(n41007), .Z(n41001) );
  OR U50200 ( .A(n41008), .B(n41009), .Z(n41007) );
  OR U50201 ( .A(n41010), .B(n41011), .Z(n41006) );
  NAND U50202 ( .A(n41012), .B(n41013), .Z(n40999) );
  OR U50203 ( .A(n41014), .B(n41015), .Z(n41013) );
  OR U50204 ( .A(n41016), .B(n41017), .Z(n41012) );
  NOR U50205 ( .A(n41018), .B(n41019), .Z(n41000) );
  ANDN U50206 ( .B(n41020), .A(n41021), .Z(n40994) );
  XNOR U50207 ( .A(n40987), .B(n41022), .Z(n40993) );
  XNOR U50208 ( .A(n40986), .B(n40988), .Z(n41022) );
  NAND U50209 ( .A(n41023), .B(n41024), .Z(n40988) );
  OR U50210 ( .A(n41025), .B(n41026), .Z(n41024) );
  OR U50211 ( .A(n41027), .B(n41028), .Z(n41023) );
  NAND U50212 ( .A(n41029), .B(n41030), .Z(n40986) );
  OR U50213 ( .A(n41031), .B(n41032), .Z(n41030) );
  OR U50214 ( .A(n41033), .B(n41034), .Z(n41029) );
  ANDN U50215 ( .B(n41035), .A(n41036), .Z(n40987) );
  IV U50216 ( .A(n41037), .Z(n41035) );
  ANDN U50217 ( .B(n41038), .A(n41039), .Z(n40979) );
  XOR U50218 ( .A(n40965), .B(n41040), .Z(n40977) );
  XOR U50219 ( .A(n40966), .B(n40967), .Z(n41040) );
  XOR U50220 ( .A(n40972), .B(n41041), .Z(n40967) );
  XOR U50221 ( .A(n40971), .B(n40974), .Z(n41041) );
  IV U50222 ( .A(n40973), .Z(n40974) );
  NAND U50223 ( .A(n41042), .B(n41043), .Z(n40973) );
  OR U50224 ( .A(n41044), .B(n41045), .Z(n41043) );
  OR U50225 ( .A(n41046), .B(n41047), .Z(n41042) );
  NAND U50226 ( .A(n41048), .B(n41049), .Z(n40971) );
  OR U50227 ( .A(n41050), .B(n41051), .Z(n41049) );
  OR U50228 ( .A(n41052), .B(n41053), .Z(n41048) );
  NOR U50229 ( .A(n41054), .B(n41055), .Z(n40972) );
  ANDN U50230 ( .B(n41056), .A(n41057), .Z(n40966) );
  IV U50231 ( .A(n41058), .Z(n41056) );
  XNOR U50232 ( .A(n40959), .B(n41059), .Z(n40965) );
  XNOR U50233 ( .A(n40958), .B(n40960), .Z(n41059) );
  NAND U50234 ( .A(n41060), .B(n41061), .Z(n40960) );
  OR U50235 ( .A(n41062), .B(n41063), .Z(n41061) );
  OR U50236 ( .A(n41064), .B(n41065), .Z(n41060) );
  NAND U50237 ( .A(n41066), .B(n41067), .Z(n40958) );
  OR U50238 ( .A(n41068), .B(n41069), .Z(n41067) );
  OR U50239 ( .A(n41070), .B(n41071), .Z(n41066) );
  ANDN U50240 ( .B(n41072), .A(n41073), .Z(n40959) );
  IV U50241 ( .A(n41074), .Z(n41072) );
  XNOR U50242 ( .A(n41039), .B(n41038), .Z(N61762) );
  XOR U50243 ( .A(n41058), .B(n41057), .Z(n41038) );
  XNOR U50244 ( .A(n41073), .B(n41074), .Z(n41057) );
  XNOR U50245 ( .A(n41068), .B(n41069), .Z(n41074) );
  XNOR U50246 ( .A(n41070), .B(n41071), .Z(n41069) );
  XNOR U50247 ( .A(y[2173]), .B(x[2173]), .Z(n41071) );
  XNOR U50248 ( .A(y[2174]), .B(x[2174]), .Z(n41070) );
  XNOR U50249 ( .A(y[2172]), .B(x[2172]), .Z(n41068) );
  XNOR U50250 ( .A(n41062), .B(n41063), .Z(n41073) );
  XNOR U50251 ( .A(y[2169]), .B(x[2169]), .Z(n41063) );
  XNOR U50252 ( .A(n41064), .B(n41065), .Z(n41062) );
  XNOR U50253 ( .A(y[2170]), .B(x[2170]), .Z(n41065) );
  XNOR U50254 ( .A(y[2171]), .B(x[2171]), .Z(n41064) );
  XNOR U50255 ( .A(n41055), .B(n41054), .Z(n41058) );
  XNOR U50256 ( .A(n41050), .B(n41051), .Z(n41054) );
  XNOR U50257 ( .A(y[2166]), .B(x[2166]), .Z(n41051) );
  XNOR U50258 ( .A(n41052), .B(n41053), .Z(n41050) );
  XNOR U50259 ( .A(y[2167]), .B(x[2167]), .Z(n41053) );
  XNOR U50260 ( .A(y[2168]), .B(x[2168]), .Z(n41052) );
  XNOR U50261 ( .A(n41044), .B(n41045), .Z(n41055) );
  XNOR U50262 ( .A(y[2163]), .B(x[2163]), .Z(n41045) );
  XNOR U50263 ( .A(n41046), .B(n41047), .Z(n41044) );
  XNOR U50264 ( .A(y[2164]), .B(x[2164]), .Z(n41047) );
  XNOR U50265 ( .A(y[2165]), .B(x[2165]), .Z(n41046) );
  XOR U50266 ( .A(n41020), .B(n41021), .Z(n41039) );
  XNOR U50267 ( .A(n41036), .B(n41037), .Z(n41021) );
  XNOR U50268 ( .A(n41031), .B(n41032), .Z(n41037) );
  XNOR U50269 ( .A(n41033), .B(n41034), .Z(n41032) );
  XNOR U50270 ( .A(y[2161]), .B(x[2161]), .Z(n41034) );
  XNOR U50271 ( .A(y[2162]), .B(x[2162]), .Z(n41033) );
  XNOR U50272 ( .A(y[2160]), .B(x[2160]), .Z(n41031) );
  XNOR U50273 ( .A(n41025), .B(n41026), .Z(n41036) );
  XNOR U50274 ( .A(y[2157]), .B(x[2157]), .Z(n41026) );
  XNOR U50275 ( .A(n41027), .B(n41028), .Z(n41025) );
  XNOR U50276 ( .A(y[2158]), .B(x[2158]), .Z(n41028) );
  XNOR U50277 ( .A(y[2159]), .B(x[2159]), .Z(n41027) );
  XOR U50278 ( .A(n41019), .B(n41018), .Z(n41020) );
  XNOR U50279 ( .A(n41014), .B(n41015), .Z(n41018) );
  XNOR U50280 ( .A(y[2154]), .B(x[2154]), .Z(n41015) );
  XNOR U50281 ( .A(n41016), .B(n41017), .Z(n41014) );
  XNOR U50282 ( .A(y[2155]), .B(x[2155]), .Z(n41017) );
  XNOR U50283 ( .A(y[2156]), .B(x[2156]), .Z(n41016) );
  XNOR U50284 ( .A(n41008), .B(n41009), .Z(n41019) );
  XNOR U50285 ( .A(y[2151]), .B(x[2151]), .Z(n41009) );
  XNOR U50286 ( .A(n41010), .B(n41011), .Z(n41008) );
  XNOR U50287 ( .A(y[2152]), .B(x[2152]), .Z(n41011) );
  XNOR U50288 ( .A(y[2153]), .B(x[2153]), .Z(n41010) );
  NAND U50289 ( .A(n41075), .B(n41076), .Z(N61753) );
  NANDN U50290 ( .A(n41077), .B(n41078), .Z(n41076) );
  OR U50291 ( .A(n41079), .B(n41080), .Z(n41078) );
  NAND U50292 ( .A(n41079), .B(n41080), .Z(n41075) );
  XOR U50293 ( .A(n41079), .B(n41081), .Z(N61752) );
  XNOR U50294 ( .A(n41077), .B(n41080), .Z(n41081) );
  AND U50295 ( .A(n41082), .B(n41083), .Z(n41080) );
  NANDN U50296 ( .A(n41084), .B(n41085), .Z(n41083) );
  NANDN U50297 ( .A(n41086), .B(n41087), .Z(n41085) );
  NANDN U50298 ( .A(n41087), .B(n41086), .Z(n41082) );
  NAND U50299 ( .A(n41088), .B(n41089), .Z(n41077) );
  NANDN U50300 ( .A(n41090), .B(n41091), .Z(n41089) );
  OR U50301 ( .A(n41092), .B(n41093), .Z(n41091) );
  NAND U50302 ( .A(n41093), .B(n41092), .Z(n41088) );
  AND U50303 ( .A(n41094), .B(n41095), .Z(n41079) );
  NANDN U50304 ( .A(n41096), .B(n41097), .Z(n41095) );
  NANDN U50305 ( .A(n41098), .B(n41099), .Z(n41097) );
  NANDN U50306 ( .A(n41099), .B(n41098), .Z(n41094) );
  XOR U50307 ( .A(n41093), .B(n41100), .Z(N61751) );
  XOR U50308 ( .A(n41090), .B(n41092), .Z(n41100) );
  XNOR U50309 ( .A(n41086), .B(n41101), .Z(n41092) );
  XNOR U50310 ( .A(n41084), .B(n41087), .Z(n41101) );
  NAND U50311 ( .A(n41102), .B(n41103), .Z(n41087) );
  NAND U50312 ( .A(n41104), .B(n41105), .Z(n41103) );
  OR U50313 ( .A(n41106), .B(n41107), .Z(n41104) );
  NANDN U50314 ( .A(n41108), .B(n41106), .Z(n41102) );
  IV U50315 ( .A(n41107), .Z(n41108) );
  NAND U50316 ( .A(n41109), .B(n41110), .Z(n41084) );
  NAND U50317 ( .A(n41111), .B(n41112), .Z(n41110) );
  NANDN U50318 ( .A(n41113), .B(n41114), .Z(n41111) );
  NANDN U50319 ( .A(n41114), .B(n41113), .Z(n41109) );
  AND U50320 ( .A(n41115), .B(n41116), .Z(n41086) );
  NAND U50321 ( .A(n41117), .B(n41118), .Z(n41116) );
  OR U50322 ( .A(n41119), .B(n41120), .Z(n41117) );
  NANDN U50323 ( .A(n41121), .B(n41119), .Z(n41115) );
  NAND U50324 ( .A(n41122), .B(n41123), .Z(n41090) );
  NANDN U50325 ( .A(n41124), .B(n41125), .Z(n41123) );
  OR U50326 ( .A(n41126), .B(n41127), .Z(n41125) );
  NANDN U50327 ( .A(n41128), .B(n41126), .Z(n41122) );
  IV U50328 ( .A(n41127), .Z(n41128) );
  XNOR U50329 ( .A(n41098), .B(n41129), .Z(n41093) );
  XNOR U50330 ( .A(n41096), .B(n41099), .Z(n41129) );
  NAND U50331 ( .A(n41130), .B(n41131), .Z(n41099) );
  NAND U50332 ( .A(n41132), .B(n41133), .Z(n41131) );
  OR U50333 ( .A(n41134), .B(n41135), .Z(n41132) );
  NANDN U50334 ( .A(n41136), .B(n41134), .Z(n41130) );
  IV U50335 ( .A(n41135), .Z(n41136) );
  NAND U50336 ( .A(n41137), .B(n41138), .Z(n41096) );
  NAND U50337 ( .A(n41139), .B(n41140), .Z(n41138) );
  NANDN U50338 ( .A(n41141), .B(n41142), .Z(n41139) );
  NANDN U50339 ( .A(n41142), .B(n41141), .Z(n41137) );
  AND U50340 ( .A(n41143), .B(n41144), .Z(n41098) );
  NAND U50341 ( .A(n41145), .B(n41146), .Z(n41144) );
  OR U50342 ( .A(n41147), .B(n41148), .Z(n41145) );
  NANDN U50343 ( .A(n41149), .B(n41147), .Z(n41143) );
  XNOR U50344 ( .A(n41124), .B(n41150), .Z(N61750) );
  XOR U50345 ( .A(n41126), .B(n41127), .Z(n41150) );
  XNOR U50346 ( .A(n41140), .B(n41151), .Z(n41127) );
  XOR U50347 ( .A(n41141), .B(n41142), .Z(n41151) );
  XOR U50348 ( .A(n41147), .B(n41152), .Z(n41142) );
  XOR U50349 ( .A(n41146), .B(n41149), .Z(n41152) );
  IV U50350 ( .A(n41148), .Z(n41149) );
  NAND U50351 ( .A(n41153), .B(n41154), .Z(n41148) );
  OR U50352 ( .A(n41155), .B(n41156), .Z(n41154) );
  OR U50353 ( .A(n41157), .B(n41158), .Z(n41153) );
  NAND U50354 ( .A(n41159), .B(n41160), .Z(n41146) );
  OR U50355 ( .A(n41161), .B(n41162), .Z(n41160) );
  OR U50356 ( .A(n41163), .B(n41164), .Z(n41159) );
  NOR U50357 ( .A(n41165), .B(n41166), .Z(n41147) );
  ANDN U50358 ( .B(n41167), .A(n41168), .Z(n41141) );
  XNOR U50359 ( .A(n41134), .B(n41169), .Z(n41140) );
  XNOR U50360 ( .A(n41133), .B(n41135), .Z(n41169) );
  NAND U50361 ( .A(n41170), .B(n41171), .Z(n41135) );
  OR U50362 ( .A(n41172), .B(n41173), .Z(n41171) );
  OR U50363 ( .A(n41174), .B(n41175), .Z(n41170) );
  NAND U50364 ( .A(n41176), .B(n41177), .Z(n41133) );
  OR U50365 ( .A(n41178), .B(n41179), .Z(n41177) );
  OR U50366 ( .A(n41180), .B(n41181), .Z(n41176) );
  ANDN U50367 ( .B(n41182), .A(n41183), .Z(n41134) );
  IV U50368 ( .A(n41184), .Z(n41182) );
  ANDN U50369 ( .B(n41185), .A(n41186), .Z(n41126) );
  XOR U50370 ( .A(n41112), .B(n41187), .Z(n41124) );
  XOR U50371 ( .A(n41113), .B(n41114), .Z(n41187) );
  XOR U50372 ( .A(n41119), .B(n41188), .Z(n41114) );
  XOR U50373 ( .A(n41118), .B(n41121), .Z(n41188) );
  IV U50374 ( .A(n41120), .Z(n41121) );
  NAND U50375 ( .A(n41189), .B(n41190), .Z(n41120) );
  OR U50376 ( .A(n41191), .B(n41192), .Z(n41190) );
  OR U50377 ( .A(n41193), .B(n41194), .Z(n41189) );
  NAND U50378 ( .A(n41195), .B(n41196), .Z(n41118) );
  OR U50379 ( .A(n41197), .B(n41198), .Z(n41196) );
  OR U50380 ( .A(n41199), .B(n41200), .Z(n41195) );
  NOR U50381 ( .A(n41201), .B(n41202), .Z(n41119) );
  ANDN U50382 ( .B(n41203), .A(n41204), .Z(n41113) );
  IV U50383 ( .A(n41205), .Z(n41203) );
  XNOR U50384 ( .A(n41106), .B(n41206), .Z(n41112) );
  XNOR U50385 ( .A(n41105), .B(n41107), .Z(n41206) );
  NAND U50386 ( .A(n41207), .B(n41208), .Z(n41107) );
  OR U50387 ( .A(n41209), .B(n41210), .Z(n41208) );
  OR U50388 ( .A(n41211), .B(n41212), .Z(n41207) );
  NAND U50389 ( .A(n41213), .B(n41214), .Z(n41105) );
  OR U50390 ( .A(n41215), .B(n41216), .Z(n41214) );
  OR U50391 ( .A(n41217), .B(n41218), .Z(n41213) );
  ANDN U50392 ( .B(n41219), .A(n41220), .Z(n41106) );
  IV U50393 ( .A(n41221), .Z(n41219) );
  XNOR U50394 ( .A(n41186), .B(n41185), .Z(N61749) );
  XOR U50395 ( .A(n41205), .B(n41204), .Z(n41185) );
  XNOR U50396 ( .A(n41220), .B(n41221), .Z(n41204) );
  XNOR U50397 ( .A(n41215), .B(n41216), .Z(n41221) );
  XNOR U50398 ( .A(n41217), .B(n41218), .Z(n41216) );
  XNOR U50399 ( .A(y[2149]), .B(x[2149]), .Z(n41218) );
  XNOR U50400 ( .A(y[2150]), .B(x[2150]), .Z(n41217) );
  XNOR U50401 ( .A(y[2148]), .B(x[2148]), .Z(n41215) );
  XNOR U50402 ( .A(n41209), .B(n41210), .Z(n41220) );
  XNOR U50403 ( .A(y[2145]), .B(x[2145]), .Z(n41210) );
  XNOR U50404 ( .A(n41211), .B(n41212), .Z(n41209) );
  XNOR U50405 ( .A(y[2146]), .B(x[2146]), .Z(n41212) );
  XNOR U50406 ( .A(y[2147]), .B(x[2147]), .Z(n41211) );
  XNOR U50407 ( .A(n41202), .B(n41201), .Z(n41205) );
  XNOR U50408 ( .A(n41197), .B(n41198), .Z(n41201) );
  XNOR U50409 ( .A(y[2142]), .B(x[2142]), .Z(n41198) );
  XNOR U50410 ( .A(n41199), .B(n41200), .Z(n41197) );
  XNOR U50411 ( .A(y[2143]), .B(x[2143]), .Z(n41200) );
  XNOR U50412 ( .A(y[2144]), .B(x[2144]), .Z(n41199) );
  XNOR U50413 ( .A(n41191), .B(n41192), .Z(n41202) );
  XNOR U50414 ( .A(y[2139]), .B(x[2139]), .Z(n41192) );
  XNOR U50415 ( .A(n41193), .B(n41194), .Z(n41191) );
  XNOR U50416 ( .A(y[2140]), .B(x[2140]), .Z(n41194) );
  XNOR U50417 ( .A(y[2141]), .B(x[2141]), .Z(n41193) );
  XOR U50418 ( .A(n41167), .B(n41168), .Z(n41186) );
  XNOR U50419 ( .A(n41183), .B(n41184), .Z(n41168) );
  XNOR U50420 ( .A(n41178), .B(n41179), .Z(n41184) );
  XNOR U50421 ( .A(n41180), .B(n41181), .Z(n41179) );
  XNOR U50422 ( .A(y[2137]), .B(x[2137]), .Z(n41181) );
  XNOR U50423 ( .A(y[2138]), .B(x[2138]), .Z(n41180) );
  XNOR U50424 ( .A(y[2136]), .B(x[2136]), .Z(n41178) );
  XNOR U50425 ( .A(n41172), .B(n41173), .Z(n41183) );
  XNOR U50426 ( .A(y[2133]), .B(x[2133]), .Z(n41173) );
  XNOR U50427 ( .A(n41174), .B(n41175), .Z(n41172) );
  XNOR U50428 ( .A(y[2134]), .B(x[2134]), .Z(n41175) );
  XNOR U50429 ( .A(y[2135]), .B(x[2135]), .Z(n41174) );
  XOR U50430 ( .A(n41166), .B(n41165), .Z(n41167) );
  XNOR U50431 ( .A(n41161), .B(n41162), .Z(n41165) );
  XNOR U50432 ( .A(y[2130]), .B(x[2130]), .Z(n41162) );
  XNOR U50433 ( .A(n41163), .B(n41164), .Z(n41161) );
  XNOR U50434 ( .A(y[2131]), .B(x[2131]), .Z(n41164) );
  XNOR U50435 ( .A(y[2132]), .B(x[2132]), .Z(n41163) );
  XNOR U50436 ( .A(n41155), .B(n41156), .Z(n41166) );
  XNOR U50437 ( .A(y[2127]), .B(x[2127]), .Z(n41156) );
  XNOR U50438 ( .A(n41157), .B(n41158), .Z(n41155) );
  XNOR U50439 ( .A(y[2128]), .B(x[2128]), .Z(n41158) );
  XNOR U50440 ( .A(y[2129]), .B(x[2129]), .Z(n41157) );
  NAND U50441 ( .A(n41222), .B(n41223), .Z(N61740) );
  NANDN U50442 ( .A(n41224), .B(n41225), .Z(n41223) );
  OR U50443 ( .A(n41226), .B(n41227), .Z(n41225) );
  NAND U50444 ( .A(n41226), .B(n41227), .Z(n41222) );
  XOR U50445 ( .A(n41226), .B(n41228), .Z(N61739) );
  XNOR U50446 ( .A(n41224), .B(n41227), .Z(n41228) );
  AND U50447 ( .A(n41229), .B(n41230), .Z(n41227) );
  NANDN U50448 ( .A(n41231), .B(n41232), .Z(n41230) );
  NANDN U50449 ( .A(n41233), .B(n41234), .Z(n41232) );
  NANDN U50450 ( .A(n41234), .B(n41233), .Z(n41229) );
  NAND U50451 ( .A(n41235), .B(n41236), .Z(n41224) );
  NANDN U50452 ( .A(n41237), .B(n41238), .Z(n41236) );
  OR U50453 ( .A(n41239), .B(n41240), .Z(n41238) );
  NAND U50454 ( .A(n41240), .B(n41239), .Z(n41235) );
  AND U50455 ( .A(n41241), .B(n41242), .Z(n41226) );
  NANDN U50456 ( .A(n41243), .B(n41244), .Z(n41242) );
  NANDN U50457 ( .A(n41245), .B(n41246), .Z(n41244) );
  NANDN U50458 ( .A(n41246), .B(n41245), .Z(n41241) );
  XOR U50459 ( .A(n41240), .B(n41247), .Z(N61738) );
  XOR U50460 ( .A(n41237), .B(n41239), .Z(n41247) );
  XNOR U50461 ( .A(n41233), .B(n41248), .Z(n41239) );
  XNOR U50462 ( .A(n41231), .B(n41234), .Z(n41248) );
  NAND U50463 ( .A(n41249), .B(n41250), .Z(n41234) );
  NAND U50464 ( .A(n41251), .B(n41252), .Z(n41250) );
  OR U50465 ( .A(n41253), .B(n41254), .Z(n41251) );
  NANDN U50466 ( .A(n41255), .B(n41253), .Z(n41249) );
  IV U50467 ( .A(n41254), .Z(n41255) );
  NAND U50468 ( .A(n41256), .B(n41257), .Z(n41231) );
  NAND U50469 ( .A(n41258), .B(n41259), .Z(n41257) );
  NANDN U50470 ( .A(n41260), .B(n41261), .Z(n41258) );
  NANDN U50471 ( .A(n41261), .B(n41260), .Z(n41256) );
  AND U50472 ( .A(n41262), .B(n41263), .Z(n41233) );
  NAND U50473 ( .A(n41264), .B(n41265), .Z(n41263) );
  OR U50474 ( .A(n41266), .B(n41267), .Z(n41264) );
  NANDN U50475 ( .A(n41268), .B(n41266), .Z(n41262) );
  NAND U50476 ( .A(n41269), .B(n41270), .Z(n41237) );
  NANDN U50477 ( .A(n41271), .B(n41272), .Z(n41270) );
  OR U50478 ( .A(n41273), .B(n41274), .Z(n41272) );
  NANDN U50479 ( .A(n41275), .B(n41273), .Z(n41269) );
  IV U50480 ( .A(n41274), .Z(n41275) );
  XNOR U50481 ( .A(n41245), .B(n41276), .Z(n41240) );
  XNOR U50482 ( .A(n41243), .B(n41246), .Z(n41276) );
  NAND U50483 ( .A(n41277), .B(n41278), .Z(n41246) );
  NAND U50484 ( .A(n41279), .B(n41280), .Z(n41278) );
  OR U50485 ( .A(n41281), .B(n41282), .Z(n41279) );
  NANDN U50486 ( .A(n41283), .B(n41281), .Z(n41277) );
  IV U50487 ( .A(n41282), .Z(n41283) );
  NAND U50488 ( .A(n41284), .B(n41285), .Z(n41243) );
  NAND U50489 ( .A(n41286), .B(n41287), .Z(n41285) );
  NANDN U50490 ( .A(n41288), .B(n41289), .Z(n41286) );
  NANDN U50491 ( .A(n41289), .B(n41288), .Z(n41284) );
  AND U50492 ( .A(n41290), .B(n41291), .Z(n41245) );
  NAND U50493 ( .A(n41292), .B(n41293), .Z(n41291) );
  OR U50494 ( .A(n41294), .B(n41295), .Z(n41292) );
  NANDN U50495 ( .A(n41296), .B(n41294), .Z(n41290) );
  XNOR U50496 ( .A(n41271), .B(n41297), .Z(N61737) );
  XOR U50497 ( .A(n41273), .B(n41274), .Z(n41297) );
  XNOR U50498 ( .A(n41287), .B(n41298), .Z(n41274) );
  XOR U50499 ( .A(n41288), .B(n41289), .Z(n41298) );
  XOR U50500 ( .A(n41294), .B(n41299), .Z(n41289) );
  XOR U50501 ( .A(n41293), .B(n41296), .Z(n41299) );
  IV U50502 ( .A(n41295), .Z(n41296) );
  NAND U50503 ( .A(n41300), .B(n41301), .Z(n41295) );
  OR U50504 ( .A(n41302), .B(n41303), .Z(n41301) );
  OR U50505 ( .A(n41304), .B(n41305), .Z(n41300) );
  NAND U50506 ( .A(n41306), .B(n41307), .Z(n41293) );
  OR U50507 ( .A(n41308), .B(n41309), .Z(n41307) );
  OR U50508 ( .A(n41310), .B(n41311), .Z(n41306) );
  NOR U50509 ( .A(n41312), .B(n41313), .Z(n41294) );
  ANDN U50510 ( .B(n41314), .A(n41315), .Z(n41288) );
  XNOR U50511 ( .A(n41281), .B(n41316), .Z(n41287) );
  XNOR U50512 ( .A(n41280), .B(n41282), .Z(n41316) );
  NAND U50513 ( .A(n41317), .B(n41318), .Z(n41282) );
  OR U50514 ( .A(n41319), .B(n41320), .Z(n41318) );
  OR U50515 ( .A(n41321), .B(n41322), .Z(n41317) );
  NAND U50516 ( .A(n41323), .B(n41324), .Z(n41280) );
  OR U50517 ( .A(n41325), .B(n41326), .Z(n41324) );
  OR U50518 ( .A(n41327), .B(n41328), .Z(n41323) );
  ANDN U50519 ( .B(n41329), .A(n41330), .Z(n41281) );
  IV U50520 ( .A(n41331), .Z(n41329) );
  ANDN U50521 ( .B(n41332), .A(n41333), .Z(n41273) );
  XOR U50522 ( .A(n41259), .B(n41334), .Z(n41271) );
  XOR U50523 ( .A(n41260), .B(n41261), .Z(n41334) );
  XOR U50524 ( .A(n41266), .B(n41335), .Z(n41261) );
  XOR U50525 ( .A(n41265), .B(n41268), .Z(n41335) );
  IV U50526 ( .A(n41267), .Z(n41268) );
  NAND U50527 ( .A(n41336), .B(n41337), .Z(n41267) );
  OR U50528 ( .A(n41338), .B(n41339), .Z(n41337) );
  OR U50529 ( .A(n41340), .B(n41341), .Z(n41336) );
  NAND U50530 ( .A(n41342), .B(n41343), .Z(n41265) );
  OR U50531 ( .A(n41344), .B(n41345), .Z(n41343) );
  OR U50532 ( .A(n41346), .B(n41347), .Z(n41342) );
  NOR U50533 ( .A(n41348), .B(n41349), .Z(n41266) );
  ANDN U50534 ( .B(n41350), .A(n41351), .Z(n41260) );
  IV U50535 ( .A(n41352), .Z(n41350) );
  XNOR U50536 ( .A(n41253), .B(n41353), .Z(n41259) );
  XNOR U50537 ( .A(n41252), .B(n41254), .Z(n41353) );
  NAND U50538 ( .A(n41354), .B(n41355), .Z(n41254) );
  OR U50539 ( .A(n41356), .B(n41357), .Z(n41355) );
  OR U50540 ( .A(n41358), .B(n41359), .Z(n41354) );
  NAND U50541 ( .A(n41360), .B(n41361), .Z(n41252) );
  OR U50542 ( .A(n41362), .B(n41363), .Z(n41361) );
  OR U50543 ( .A(n41364), .B(n41365), .Z(n41360) );
  ANDN U50544 ( .B(n41366), .A(n41367), .Z(n41253) );
  IV U50545 ( .A(n41368), .Z(n41366) );
  XNOR U50546 ( .A(n41333), .B(n41332), .Z(N61736) );
  XOR U50547 ( .A(n41352), .B(n41351), .Z(n41332) );
  XNOR U50548 ( .A(n41367), .B(n41368), .Z(n41351) );
  XNOR U50549 ( .A(n41362), .B(n41363), .Z(n41368) );
  XNOR U50550 ( .A(n41364), .B(n41365), .Z(n41363) );
  XNOR U50551 ( .A(y[2125]), .B(x[2125]), .Z(n41365) );
  XNOR U50552 ( .A(y[2126]), .B(x[2126]), .Z(n41364) );
  XNOR U50553 ( .A(y[2124]), .B(x[2124]), .Z(n41362) );
  XNOR U50554 ( .A(n41356), .B(n41357), .Z(n41367) );
  XNOR U50555 ( .A(y[2121]), .B(x[2121]), .Z(n41357) );
  XNOR U50556 ( .A(n41358), .B(n41359), .Z(n41356) );
  XNOR U50557 ( .A(y[2122]), .B(x[2122]), .Z(n41359) );
  XNOR U50558 ( .A(y[2123]), .B(x[2123]), .Z(n41358) );
  XNOR U50559 ( .A(n41349), .B(n41348), .Z(n41352) );
  XNOR U50560 ( .A(n41344), .B(n41345), .Z(n41348) );
  XNOR U50561 ( .A(y[2118]), .B(x[2118]), .Z(n41345) );
  XNOR U50562 ( .A(n41346), .B(n41347), .Z(n41344) );
  XNOR U50563 ( .A(y[2119]), .B(x[2119]), .Z(n41347) );
  XNOR U50564 ( .A(y[2120]), .B(x[2120]), .Z(n41346) );
  XNOR U50565 ( .A(n41338), .B(n41339), .Z(n41349) );
  XNOR U50566 ( .A(y[2115]), .B(x[2115]), .Z(n41339) );
  XNOR U50567 ( .A(n41340), .B(n41341), .Z(n41338) );
  XNOR U50568 ( .A(y[2116]), .B(x[2116]), .Z(n41341) );
  XNOR U50569 ( .A(y[2117]), .B(x[2117]), .Z(n41340) );
  XOR U50570 ( .A(n41314), .B(n41315), .Z(n41333) );
  XNOR U50571 ( .A(n41330), .B(n41331), .Z(n41315) );
  XNOR U50572 ( .A(n41325), .B(n41326), .Z(n41331) );
  XNOR U50573 ( .A(n41327), .B(n41328), .Z(n41326) );
  XNOR U50574 ( .A(y[2113]), .B(x[2113]), .Z(n41328) );
  XNOR U50575 ( .A(y[2114]), .B(x[2114]), .Z(n41327) );
  XNOR U50576 ( .A(y[2112]), .B(x[2112]), .Z(n41325) );
  XNOR U50577 ( .A(n41319), .B(n41320), .Z(n41330) );
  XNOR U50578 ( .A(y[2109]), .B(x[2109]), .Z(n41320) );
  XNOR U50579 ( .A(n41321), .B(n41322), .Z(n41319) );
  XNOR U50580 ( .A(y[2110]), .B(x[2110]), .Z(n41322) );
  XNOR U50581 ( .A(y[2111]), .B(x[2111]), .Z(n41321) );
  XOR U50582 ( .A(n41313), .B(n41312), .Z(n41314) );
  XNOR U50583 ( .A(n41308), .B(n41309), .Z(n41312) );
  XNOR U50584 ( .A(y[2106]), .B(x[2106]), .Z(n41309) );
  XNOR U50585 ( .A(n41310), .B(n41311), .Z(n41308) );
  XNOR U50586 ( .A(y[2107]), .B(x[2107]), .Z(n41311) );
  XNOR U50587 ( .A(y[2108]), .B(x[2108]), .Z(n41310) );
  XNOR U50588 ( .A(n41302), .B(n41303), .Z(n41313) );
  XNOR U50589 ( .A(y[2103]), .B(x[2103]), .Z(n41303) );
  XNOR U50590 ( .A(n41304), .B(n41305), .Z(n41302) );
  XNOR U50591 ( .A(y[2104]), .B(x[2104]), .Z(n41305) );
  XNOR U50592 ( .A(y[2105]), .B(x[2105]), .Z(n41304) );
  NAND U50593 ( .A(n41369), .B(n41370), .Z(N61727) );
  NANDN U50594 ( .A(n41371), .B(n41372), .Z(n41370) );
  OR U50595 ( .A(n41373), .B(n41374), .Z(n41372) );
  NAND U50596 ( .A(n41373), .B(n41374), .Z(n41369) );
  XOR U50597 ( .A(n41373), .B(n41375), .Z(N61726) );
  XNOR U50598 ( .A(n41371), .B(n41374), .Z(n41375) );
  AND U50599 ( .A(n41376), .B(n41377), .Z(n41374) );
  NANDN U50600 ( .A(n41378), .B(n41379), .Z(n41377) );
  NANDN U50601 ( .A(n41380), .B(n41381), .Z(n41379) );
  NANDN U50602 ( .A(n41381), .B(n41380), .Z(n41376) );
  NAND U50603 ( .A(n41382), .B(n41383), .Z(n41371) );
  NANDN U50604 ( .A(n41384), .B(n41385), .Z(n41383) );
  OR U50605 ( .A(n41386), .B(n41387), .Z(n41385) );
  NAND U50606 ( .A(n41387), .B(n41386), .Z(n41382) );
  AND U50607 ( .A(n41388), .B(n41389), .Z(n41373) );
  NANDN U50608 ( .A(n41390), .B(n41391), .Z(n41389) );
  NANDN U50609 ( .A(n41392), .B(n41393), .Z(n41391) );
  NANDN U50610 ( .A(n41393), .B(n41392), .Z(n41388) );
  XOR U50611 ( .A(n41387), .B(n41394), .Z(N61725) );
  XOR U50612 ( .A(n41384), .B(n41386), .Z(n41394) );
  XNOR U50613 ( .A(n41380), .B(n41395), .Z(n41386) );
  XNOR U50614 ( .A(n41378), .B(n41381), .Z(n41395) );
  NAND U50615 ( .A(n41396), .B(n41397), .Z(n41381) );
  NAND U50616 ( .A(n41398), .B(n41399), .Z(n41397) );
  OR U50617 ( .A(n41400), .B(n41401), .Z(n41398) );
  NANDN U50618 ( .A(n41402), .B(n41400), .Z(n41396) );
  IV U50619 ( .A(n41401), .Z(n41402) );
  NAND U50620 ( .A(n41403), .B(n41404), .Z(n41378) );
  NAND U50621 ( .A(n41405), .B(n41406), .Z(n41404) );
  NANDN U50622 ( .A(n41407), .B(n41408), .Z(n41405) );
  NANDN U50623 ( .A(n41408), .B(n41407), .Z(n41403) );
  AND U50624 ( .A(n41409), .B(n41410), .Z(n41380) );
  NAND U50625 ( .A(n41411), .B(n41412), .Z(n41410) );
  OR U50626 ( .A(n41413), .B(n41414), .Z(n41411) );
  NANDN U50627 ( .A(n41415), .B(n41413), .Z(n41409) );
  NAND U50628 ( .A(n41416), .B(n41417), .Z(n41384) );
  NANDN U50629 ( .A(n41418), .B(n41419), .Z(n41417) );
  OR U50630 ( .A(n41420), .B(n41421), .Z(n41419) );
  NANDN U50631 ( .A(n41422), .B(n41420), .Z(n41416) );
  IV U50632 ( .A(n41421), .Z(n41422) );
  XNOR U50633 ( .A(n41392), .B(n41423), .Z(n41387) );
  XNOR U50634 ( .A(n41390), .B(n41393), .Z(n41423) );
  NAND U50635 ( .A(n41424), .B(n41425), .Z(n41393) );
  NAND U50636 ( .A(n41426), .B(n41427), .Z(n41425) );
  OR U50637 ( .A(n41428), .B(n41429), .Z(n41426) );
  NANDN U50638 ( .A(n41430), .B(n41428), .Z(n41424) );
  IV U50639 ( .A(n41429), .Z(n41430) );
  NAND U50640 ( .A(n41431), .B(n41432), .Z(n41390) );
  NAND U50641 ( .A(n41433), .B(n41434), .Z(n41432) );
  NANDN U50642 ( .A(n41435), .B(n41436), .Z(n41433) );
  NANDN U50643 ( .A(n41436), .B(n41435), .Z(n41431) );
  AND U50644 ( .A(n41437), .B(n41438), .Z(n41392) );
  NAND U50645 ( .A(n41439), .B(n41440), .Z(n41438) );
  OR U50646 ( .A(n41441), .B(n41442), .Z(n41439) );
  NANDN U50647 ( .A(n41443), .B(n41441), .Z(n41437) );
  XNOR U50648 ( .A(n41418), .B(n41444), .Z(N61724) );
  XOR U50649 ( .A(n41420), .B(n41421), .Z(n41444) );
  XNOR U50650 ( .A(n41434), .B(n41445), .Z(n41421) );
  XOR U50651 ( .A(n41435), .B(n41436), .Z(n41445) );
  XOR U50652 ( .A(n41441), .B(n41446), .Z(n41436) );
  XOR U50653 ( .A(n41440), .B(n41443), .Z(n41446) );
  IV U50654 ( .A(n41442), .Z(n41443) );
  NAND U50655 ( .A(n41447), .B(n41448), .Z(n41442) );
  OR U50656 ( .A(n41449), .B(n41450), .Z(n41448) );
  OR U50657 ( .A(n41451), .B(n41452), .Z(n41447) );
  NAND U50658 ( .A(n41453), .B(n41454), .Z(n41440) );
  OR U50659 ( .A(n41455), .B(n41456), .Z(n41454) );
  OR U50660 ( .A(n41457), .B(n41458), .Z(n41453) );
  NOR U50661 ( .A(n41459), .B(n41460), .Z(n41441) );
  ANDN U50662 ( .B(n41461), .A(n41462), .Z(n41435) );
  XNOR U50663 ( .A(n41428), .B(n41463), .Z(n41434) );
  XNOR U50664 ( .A(n41427), .B(n41429), .Z(n41463) );
  NAND U50665 ( .A(n41464), .B(n41465), .Z(n41429) );
  OR U50666 ( .A(n41466), .B(n41467), .Z(n41465) );
  OR U50667 ( .A(n41468), .B(n41469), .Z(n41464) );
  NAND U50668 ( .A(n41470), .B(n41471), .Z(n41427) );
  OR U50669 ( .A(n41472), .B(n41473), .Z(n41471) );
  OR U50670 ( .A(n41474), .B(n41475), .Z(n41470) );
  ANDN U50671 ( .B(n41476), .A(n41477), .Z(n41428) );
  IV U50672 ( .A(n41478), .Z(n41476) );
  ANDN U50673 ( .B(n41479), .A(n41480), .Z(n41420) );
  XOR U50674 ( .A(n41406), .B(n41481), .Z(n41418) );
  XOR U50675 ( .A(n41407), .B(n41408), .Z(n41481) );
  XOR U50676 ( .A(n41413), .B(n41482), .Z(n41408) );
  XOR U50677 ( .A(n41412), .B(n41415), .Z(n41482) );
  IV U50678 ( .A(n41414), .Z(n41415) );
  NAND U50679 ( .A(n41483), .B(n41484), .Z(n41414) );
  OR U50680 ( .A(n41485), .B(n41486), .Z(n41484) );
  OR U50681 ( .A(n41487), .B(n41488), .Z(n41483) );
  NAND U50682 ( .A(n41489), .B(n41490), .Z(n41412) );
  OR U50683 ( .A(n41491), .B(n41492), .Z(n41490) );
  OR U50684 ( .A(n41493), .B(n41494), .Z(n41489) );
  NOR U50685 ( .A(n41495), .B(n41496), .Z(n41413) );
  ANDN U50686 ( .B(n41497), .A(n41498), .Z(n41407) );
  IV U50687 ( .A(n41499), .Z(n41497) );
  XNOR U50688 ( .A(n41400), .B(n41500), .Z(n41406) );
  XNOR U50689 ( .A(n41399), .B(n41401), .Z(n41500) );
  NAND U50690 ( .A(n41501), .B(n41502), .Z(n41401) );
  OR U50691 ( .A(n41503), .B(n41504), .Z(n41502) );
  OR U50692 ( .A(n41505), .B(n41506), .Z(n41501) );
  NAND U50693 ( .A(n41507), .B(n41508), .Z(n41399) );
  OR U50694 ( .A(n41509), .B(n41510), .Z(n41508) );
  OR U50695 ( .A(n41511), .B(n41512), .Z(n41507) );
  ANDN U50696 ( .B(n41513), .A(n41514), .Z(n41400) );
  IV U50697 ( .A(n41515), .Z(n41513) );
  XNOR U50698 ( .A(n41480), .B(n41479), .Z(N61723) );
  XOR U50699 ( .A(n41499), .B(n41498), .Z(n41479) );
  XNOR U50700 ( .A(n41514), .B(n41515), .Z(n41498) );
  XNOR U50701 ( .A(n41509), .B(n41510), .Z(n41515) );
  XNOR U50702 ( .A(n41511), .B(n41512), .Z(n41510) );
  XNOR U50703 ( .A(y[2101]), .B(x[2101]), .Z(n41512) );
  XNOR U50704 ( .A(y[2102]), .B(x[2102]), .Z(n41511) );
  XNOR U50705 ( .A(y[2100]), .B(x[2100]), .Z(n41509) );
  XNOR U50706 ( .A(n41503), .B(n41504), .Z(n41514) );
  XNOR U50707 ( .A(y[2097]), .B(x[2097]), .Z(n41504) );
  XNOR U50708 ( .A(n41505), .B(n41506), .Z(n41503) );
  XNOR U50709 ( .A(y[2098]), .B(x[2098]), .Z(n41506) );
  XNOR U50710 ( .A(y[2099]), .B(x[2099]), .Z(n41505) );
  XNOR U50711 ( .A(n41496), .B(n41495), .Z(n41499) );
  XNOR U50712 ( .A(n41491), .B(n41492), .Z(n41495) );
  XNOR U50713 ( .A(y[2094]), .B(x[2094]), .Z(n41492) );
  XNOR U50714 ( .A(n41493), .B(n41494), .Z(n41491) );
  XNOR U50715 ( .A(y[2095]), .B(x[2095]), .Z(n41494) );
  XNOR U50716 ( .A(y[2096]), .B(x[2096]), .Z(n41493) );
  XNOR U50717 ( .A(n41485), .B(n41486), .Z(n41496) );
  XNOR U50718 ( .A(y[2091]), .B(x[2091]), .Z(n41486) );
  XNOR U50719 ( .A(n41487), .B(n41488), .Z(n41485) );
  XNOR U50720 ( .A(y[2092]), .B(x[2092]), .Z(n41488) );
  XNOR U50721 ( .A(y[2093]), .B(x[2093]), .Z(n41487) );
  XOR U50722 ( .A(n41461), .B(n41462), .Z(n41480) );
  XNOR U50723 ( .A(n41477), .B(n41478), .Z(n41462) );
  XNOR U50724 ( .A(n41472), .B(n41473), .Z(n41478) );
  XNOR U50725 ( .A(n41474), .B(n41475), .Z(n41473) );
  XNOR U50726 ( .A(y[2089]), .B(x[2089]), .Z(n41475) );
  XNOR U50727 ( .A(y[2090]), .B(x[2090]), .Z(n41474) );
  XNOR U50728 ( .A(y[2088]), .B(x[2088]), .Z(n41472) );
  XNOR U50729 ( .A(n41466), .B(n41467), .Z(n41477) );
  XNOR U50730 ( .A(y[2085]), .B(x[2085]), .Z(n41467) );
  XNOR U50731 ( .A(n41468), .B(n41469), .Z(n41466) );
  XNOR U50732 ( .A(y[2086]), .B(x[2086]), .Z(n41469) );
  XNOR U50733 ( .A(y[2087]), .B(x[2087]), .Z(n41468) );
  XOR U50734 ( .A(n41460), .B(n41459), .Z(n41461) );
  XNOR U50735 ( .A(n41455), .B(n41456), .Z(n41459) );
  XNOR U50736 ( .A(y[2082]), .B(x[2082]), .Z(n41456) );
  XNOR U50737 ( .A(n41457), .B(n41458), .Z(n41455) );
  XNOR U50738 ( .A(y[2083]), .B(x[2083]), .Z(n41458) );
  XNOR U50739 ( .A(y[2084]), .B(x[2084]), .Z(n41457) );
  XNOR U50740 ( .A(n41449), .B(n41450), .Z(n41460) );
  XNOR U50741 ( .A(y[2079]), .B(x[2079]), .Z(n41450) );
  XNOR U50742 ( .A(n41451), .B(n41452), .Z(n41449) );
  XNOR U50743 ( .A(y[2080]), .B(x[2080]), .Z(n41452) );
  XNOR U50744 ( .A(y[2081]), .B(x[2081]), .Z(n41451) );
  NAND U50745 ( .A(n41516), .B(n41517), .Z(N61714) );
  NANDN U50746 ( .A(n41518), .B(n41519), .Z(n41517) );
  OR U50747 ( .A(n41520), .B(n41521), .Z(n41519) );
  NAND U50748 ( .A(n41520), .B(n41521), .Z(n41516) );
  XOR U50749 ( .A(n41520), .B(n41522), .Z(N61713) );
  XNOR U50750 ( .A(n41518), .B(n41521), .Z(n41522) );
  AND U50751 ( .A(n41523), .B(n41524), .Z(n41521) );
  NANDN U50752 ( .A(n41525), .B(n41526), .Z(n41524) );
  NANDN U50753 ( .A(n41527), .B(n41528), .Z(n41526) );
  NANDN U50754 ( .A(n41528), .B(n41527), .Z(n41523) );
  NAND U50755 ( .A(n41529), .B(n41530), .Z(n41518) );
  NANDN U50756 ( .A(n41531), .B(n41532), .Z(n41530) );
  OR U50757 ( .A(n41533), .B(n41534), .Z(n41532) );
  NAND U50758 ( .A(n41534), .B(n41533), .Z(n41529) );
  AND U50759 ( .A(n41535), .B(n41536), .Z(n41520) );
  NANDN U50760 ( .A(n41537), .B(n41538), .Z(n41536) );
  NANDN U50761 ( .A(n41539), .B(n41540), .Z(n41538) );
  NANDN U50762 ( .A(n41540), .B(n41539), .Z(n41535) );
  XOR U50763 ( .A(n41534), .B(n41541), .Z(N61712) );
  XOR U50764 ( .A(n41531), .B(n41533), .Z(n41541) );
  XNOR U50765 ( .A(n41527), .B(n41542), .Z(n41533) );
  XNOR U50766 ( .A(n41525), .B(n41528), .Z(n41542) );
  NAND U50767 ( .A(n41543), .B(n41544), .Z(n41528) );
  NAND U50768 ( .A(n41545), .B(n41546), .Z(n41544) );
  OR U50769 ( .A(n41547), .B(n41548), .Z(n41545) );
  NANDN U50770 ( .A(n41549), .B(n41547), .Z(n41543) );
  IV U50771 ( .A(n41548), .Z(n41549) );
  NAND U50772 ( .A(n41550), .B(n41551), .Z(n41525) );
  NAND U50773 ( .A(n41552), .B(n41553), .Z(n41551) );
  NANDN U50774 ( .A(n41554), .B(n41555), .Z(n41552) );
  NANDN U50775 ( .A(n41555), .B(n41554), .Z(n41550) );
  AND U50776 ( .A(n41556), .B(n41557), .Z(n41527) );
  NAND U50777 ( .A(n41558), .B(n41559), .Z(n41557) );
  OR U50778 ( .A(n41560), .B(n41561), .Z(n41558) );
  NANDN U50779 ( .A(n41562), .B(n41560), .Z(n41556) );
  NAND U50780 ( .A(n41563), .B(n41564), .Z(n41531) );
  NANDN U50781 ( .A(n41565), .B(n41566), .Z(n41564) );
  OR U50782 ( .A(n41567), .B(n41568), .Z(n41566) );
  NANDN U50783 ( .A(n41569), .B(n41567), .Z(n41563) );
  IV U50784 ( .A(n41568), .Z(n41569) );
  XNOR U50785 ( .A(n41539), .B(n41570), .Z(n41534) );
  XNOR U50786 ( .A(n41537), .B(n41540), .Z(n41570) );
  NAND U50787 ( .A(n41571), .B(n41572), .Z(n41540) );
  NAND U50788 ( .A(n41573), .B(n41574), .Z(n41572) );
  OR U50789 ( .A(n41575), .B(n41576), .Z(n41573) );
  NANDN U50790 ( .A(n41577), .B(n41575), .Z(n41571) );
  IV U50791 ( .A(n41576), .Z(n41577) );
  NAND U50792 ( .A(n41578), .B(n41579), .Z(n41537) );
  NAND U50793 ( .A(n41580), .B(n41581), .Z(n41579) );
  NANDN U50794 ( .A(n41582), .B(n41583), .Z(n41580) );
  NANDN U50795 ( .A(n41583), .B(n41582), .Z(n41578) );
  AND U50796 ( .A(n41584), .B(n41585), .Z(n41539) );
  NAND U50797 ( .A(n41586), .B(n41587), .Z(n41585) );
  OR U50798 ( .A(n41588), .B(n41589), .Z(n41586) );
  NANDN U50799 ( .A(n41590), .B(n41588), .Z(n41584) );
  XNOR U50800 ( .A(n41565), .B(n41591), .Z(N61711) );
  XOR U50801 ( .A(n41567), .B(n41568), .Z(n41591) );
  XNOR U50802 ( .A(n41581), .B(n41592), .Z(n41568) );
  XOR U50803 ( .A(n41582), .B(n41583), .Z(n41592) );
  XOR U50804 ( .A(n41588), .B(n41593), .Z(n41583) );
  XOR U50805 ( .A(n41587), .B(n41590), .Z(n41593) );
  IV U50806 ( .A(n41589), .Z(n41590) );
  NAND U50807 ( .A(n41594), .B(n41595), .Z(n41589) );
  OR U50808 ( .A(n41596), .B(n41597), .Z(n41595) );
  OR U50809 ( .A(n41598), .B(n41599), .Z(n41594) );
  NAND U50810 ( .A(n41600), .B(n41601), .Z(n41587) );
  OR U50811 ( .A(n41602), .B(n41603), .Z(n41601) );
  OR U50812 ( .A(n41604), .B(n41605), .Z(n41600) );
  NOR U50813 ( .A(n41606), .B(n41607), .Z(n41588) );
  ANDN U50814 ( .B(n41608), .A(n41609), .Z(n41582) );
  XNOR U50815 ( .A(n41575), .B(n41610), .Z(n41581) );
  XNOR U50816 ( .A(n41574), .B(n41576), .Z(n41610) );
  NAND U50817 ( .A(n41611), .B(n41612), .Z(n41576) );
  OR U50818 ( .A(n41613), .B(n41614), .Z(n41612) );
  OR U50819 ( .A(n41615), .B(n41616), .Z(n41611) );
  NAND U50820 ( .A(n41617), .B(n41618), .Z(n41574) );
  OR U50821 ( .A(n41619), .B(n41620), .Z(n41618) );
  OR U50822 ( .A(n41621), .B(n41622), .Z(n41617) );
  ANDN U50823 ( .B(n41623), .A(n41624), .Z(n41575) );
  IV U50824 ( .A(n41625), .Z(n41623) );
  ANDN U50825 ( .B(n41626), .A(n41627), .Z(n41567) );
  XOR U50826 ( .A(n41553), .B(n41628), .Z(n41565) );
  XOR U50827 ( .A(n41554), .B(n41555), .Z(n41628) );
  XOR U50828 ( .A(n41560), .B(n41629), .Z(n41555) );
  XOR U50829 ( .A(n41559), .B(n41562), .Z(n41629) );
  IV U50830 ( .A(n41561), .Z(n41562) );
  NAND U50831 ( .A(n41630), .B(n41631), .Z(n41561) );
  OR U50832 ( .A(n41632), .B(n41633), .Z(n41631) );
  OR U50833 ( .A(n41634), .B(n41635), .Z(n41630) );
  NAND U50834 ( .A(n41636), .B(n41637), .Z(n41559) );
  OR U50835 ( .A(n41638), .B(n41639), .Z(n41637) );
  OR U50836 ( .A(n41640), .B(n41641), .Z(n41636) );
  NOR U50837 ( .A(n41642), .B(n41643), .Z(n41560) );
  ANDN U50838 ( .B(n41644), .A(n41645), .Z(n41554) );
  IV U50839 ( .A(n41646), .Z(n41644) );
  XNOR U50840 ( .A(n41547), .B(n41647), .Z(n41553) );
  XNOR U50841 ( .A(n41546), .B(n41548), .Z(n41647) );
  NAND U50842 ( .A(n41648), .B(n41649), .Z(n41548) );
  OR U50843 ( .A(n41650), .B(n41651), .Z(n41649) );
  OR U50844 ( .A(n41652), .B(n41653), .Z(n41648) );
  NAND U50845 ( .A(n41654), .B(n41655), .Z(n41546) );
  OR U50846 ( .A(n41656), .B(n41657), .Z(n41655) );
  OR U50847 ( .A(n41658), .B(n41659), .Z(n41654) );
  ANDN U50848 ( .B(n41660), .A(n41661), .Z(n41547) );
  IV U50849 ( .A(n41662), .Z(n41660) );
  XNOR U50850 ( .A(n41627), .B(n41626), .Z(N61710) );
  XOR U50851 ( .A(n41646), .B(n41645), .Z(n41626) );
  XNOR U50852 ( .A(n41661), .B(n41662), .Z(n41645) );
  XNOR U50853 ( .A(n41656), .B(n41657), .Z(n41662) );
  XNOR U50854 ( .A(n41658), .B(n41659), .Z(n41657) );
  XNOR U50855 ( .A(y[2077]), .B(x[2077]), .Z(n41659) );
  XNOR U50856 ( .A(y[2078]), .B(x[2078]), .Z(n41658) );
  XNOR U50857 ( .A(y[2076]), .B(x[2076]), .Z(n41656) );
  XNOR U50858 ( .A(n41650), .B(n41651), .Z(n41661) );
  XNOR U50859 ( .A(y[2073]), .B(x[2073]), .Z(n41651) );
  XNOR U50860 ( .A(n41652), .B(n41653), .Z(n41650) );
  XNOR U50861 ( .A(y[2074]), .B(x[2074]), .Z(n41653) );
  XNOR U50862 ( .A(y[2075]), .B(x[2075]), .Z(n41652) );
  XNOR U50863 ( .A(n41643), .B(n41642), .Z(n41646) );
  XNOR U50864 ( .A(n41638), .B(n41639), .Z(n41642) );
  XNOR U50865 ( .A(y[2070]), .B(x[2070]), .Z(n41639) );
  XNOR U50866 ( .A(n41640), .B(n41641), .Z(n41638) );
  XNOR U50867 ( .A(y[2071]), .B(x[2071]), .Z(n41641) );
  XNOR U50868 ( .A(y[2072]), .B(x[2072]), .Z(n41640) );
  XNOR U50869 ( .A(n41632), .B(n41633), .Z(n41643) );
  XNOR U50870 ( .A(y[2067]), .B(x[2067]), .Z(n41633) );
  XNOR U50871 ( .A(n41634), .B(n41635), .Z(n41632) );
  XNOR U50872 ( .A(y[2068]), .B(x[2068]), .Z(n41635) );
  XNOR U50873 ( .A(y[2069]), .B(x[2069]), .Z(n41634) );
  XOR U50874 ( .A(n41608), .B(n41609), .Z(n41627) );
  XNOR U50875 ( .A(n41624), .B(n41625), .Z(n41609) );
  XNOR U50876 ( .A(n41619), .B(n41620), .Z(n41625) );
  XNOR U50877 ( .A(n41621), .B(n41622), .Z(n41620) );
  XNOR U50878 ( .A(y[2065]), .B(x[2065]), .Z(n41622) );
  XNOR U50879 ( .A(y[2066]), .B(x[2066]), .Z(n41621) );
  XNOR U50880 ( .A(y[2064]), .B(x[2064]), .Z(n41619) );
  XNOR U50881 ( .A(n41613), .B(n41614), .Z(n41624) );
  XNOR U50882 ( .A(y[2061]), .B(x[2061]), .Z(n41614) );
  XNOR U50883 ( .A(n41615), .B(n41616), .Z(n41613) );
  XNOR U50884 ( .A(y[2062]), .B(x[2062]), .Z(n41616) );
  XNOR U50885 ( .A(y[2063]), .B(x[2063]), .Z(n41615) );
  XOR U50886 ( .A(n41607), .B(n41606), .Z(n41608) );
  XNOR U50887 ( .A(n41602), .B(n41603), .Z(n41606) );
  XNOR U50888 ( .A(y[2058]), .B(x[2058]), .Z(n41603) );
  XNOR U50889 ( .A(n41604), .B(n41605), .Z(n41602) );
  XNOR U50890 ( .A(y[2059]), .B(x[2059]), .Z(n41605) );
  XNOR U50891 ( .A(y[2060]), .B(x[2060]), .Z(n41604) );
  XNOR U50892 ( .A(n41596), .B(n41597), .Z(n41607) );
  XNOR U50893 ( .A(y[2055]), .B(x[2055]), .Z(n41597) );
  XNOR U50894 ( .A(n41598), .B(n41599), .Z(n41596) );
  XNOR U50895 ( .A(y[2056]), .B(x[2056]), .Z(n41599) );
  XNOR U50896 ( .A(y[2057]), .B(x[2057]), .Z(n41598) );
  NAND U50897 ( .A(n41663), .B(n41664), .Z(N61701) );
  NANDN U50898 ( .A(n41665), .B(n41666), .Z(n41664) );
  OR U50899 ( .A(n41667), .B(n41668), .Z(n41666) );
  NAND U50900 ( .A(n41667), .B(n41668), .Z(n41663) );
  XOR U50901 ( .A(n41667), .B(n41669), .Z(N61700) );
  XNOR U50902 ( .A(n41665), .B(n41668), .Z(n41669) );
  AND U50903 ( .A(n41670), .B(n41671), .Z(n41668) );
  NANDN U50904 ( .A(n41672), .B(n41673), .Z(n41671) );
  NANDN U50905 ( .A(n41674), .B(n41675), .Z(n41673) );
  NANDN U50906 ( .A(n41675), .B(n41674), .Z(n41670) );
  NAND U50907 ( .A(n41676), .B(n41677), .Z(n41665) );
  NANDN U50908 ( .A(n41678), .B(n41679), .Z(n41677) );
  OR U50909 ( .A(n41680), .B(n41681), .Z(n41679) );
  NAND U50910 ( .A(n41681), .B(n41680), .Z(n41676) );
  AND U50911 ( .A(n41682), .B(n41683), .Z(n41667) );
  NANDN U50912 ( .A(n41684), .B(n41685), .Z(n41683) );
  NANDN U50913 ( .A(n41686), .B(n41687), .Z(n41685) );
  NANDN U50914 ( .A(n41687), .B(n41686), .Z(n41682) );
  XOR U50915 ( .A(n41681), .B(n41688), .Z(N61699) );
  XOR U50916 ( .A(n41678), .B(n41680), .Z(n41688) );
  XNOR U50917 ( .A(n41674), .B(n41689), .Z(n41680) );
  XNOR U50918 ( .A(n41672), .B(n41675), .Z(n41689) );
  NAND U50919 ( .A(n41690), .B(n41691), .Z(n41675) );
  NAND U50920 ( .A(n41692), .B(n41693), .Z(n41691) );
  OR U50921 ( .A(n41694), .B(n41695), .Z(n41692) );
  NANDN U50922 ( .A(n41696), .B(n41694), .Z(n41690) );
  IV U50923 ( .A(n41695), .Z(n41696) );
  NAND U50924 ( .A(n41697), .B(n41698), .Z(n41672) );
  NAND U50925 ( .A(n41699), .B(n41700), .Z(n41698) );
  NANDN U50926 ( .A(n41701), .B(n41702), .Z(n41699) );
  NANDN U50927 ( .A(n41702), .B(n41701), .Z(n41697) );
  AND U50928 ( .A(n41703), .B(n41704), .Z(n41674) );
  NAND U50929 ( .A(n41705), .B(n41706), .Z(n41704) );
  OR U50930 ( .A(n41707), .B(n41708), .Z(n41705) );
  NANDN U50931 ( .A(n41709), .B(n41707), .Z(n41703) );
  NAND U50932 ( .A(n41710), .B(n41711), .Z(n41678) );
  NANDN U50933 ( .A(n41712), .B(n41713), .Z(n41711) );
  OR U50934 ( .A(n41714), .B(n41715), .Z(n41713) );
  NANDN U50935 ( .A(n41716), .B(n41714), .Z(n41710) );
  IV U50936 ( .A(n41715), .Z(n41716) );
  XNOR U50937 ( .A(n41686), .B(n41717), .Z(n41681) );
  XNOR U50938 ( .A(n41684), .B(n41687), .Z(n41717) );
  NAND U50939 ( .A(n41718), .B(n41719), .Z(n41687) );
  NAND U50940 ( .A(n41720), .B(n41721), .Z(n41719) );
  OR U50941 ( .A(n41722), .B(n41723), .Z(n41720) );
  NANDN U50942 ( .A(n41724), .B(n41722), .Z(n41718) );
  IV U50943 ( .A(n41723), .Z(n41724) );
  NAND U50944 ( .A(n41725), .B(n41726), .Z(n41684) );
  NAND U50945 ( .A(n41727), .B(n41728), .Z(n41726) );
  NANDN U50946 ( .A(n41729), .B(n41730), .Z(n41727) );
  NANDN U50947 ( .A(n41730), .B(n41729), .Z(n41725) );
  AND U50948 ( .A(n41731), .B(n41732), .Z(n41686) );
  NAND U50949 ( .A(n41733), .B(n41734), .Z(n41732) );
  OR U50950 ( .A(n41735), .B(n41736), .Z(n41733) );
  NANDN U50951 ( .A(n41737), .B(n41735), .Z(n41731) );
  XNOR U50952 ( .A(n41712), .B(n41738), .Z(N61698) );
  XOR U50953 ( .A(n41714), .B(n41715), .Z(n41738) );
  XNOR U50954 ( .A(n41728), .B(n41739), .Z(n41715) );
  XOR U50955 ( .A(n41729), .B(n41730), .Z(n41739) );
  XOR U50956 ( .A(n41735), .B(n41740), .Z(n41730) );
  XOR U50957 ( .A(n41734), .B(n41737), .Z(n41740) );
  IV U50958 ( .A(n41736), .Z(n41737) );
  NAND U50959 ( .A(n41741), .B(n41742), .Z(n41736) );
  OR U50960 ( .A(n41743), .B(n41744), .Z(n41742) );
  OR U50961 ( .A(n41745), .B(n41746), .Z(n41741) );
  NAND U50962 ( .A(n41747), .B(n41748), .Z(n41734) );
  OR U50963 ( .A(n41749), .B(n41750), .Z(n41748) );
  OR U50964 ( .A(n41751), .B(n41752), .Z(n41747) );
  NOR U50965 ( .A(n41753), .B(n41754), .Z(n41735) );
  ANDN U50966 ( .B(n41755), .A(n41756), .Z(n41729) );
  XNOR U50967 ( .A(n41722), .B(n41757), .Z(n41728) );
  XNOR U50968 ( .A(n41721), .B(n41723), .Z(n41757) );
  NAND U50969 ( .A(n41758), .B(n41759), .Z(n41723) );
  OR U50970 ( .A(n41760), .B(n41761), .Z(n41759) );
  OR U50971 ( .A(n41762), .B(n41763), .Z(n41758) );
  NAND U50972 ( .A(n41764), .B(n41765), .Z(n41721) );
  OR U50973 ( .A(n41766), .B(n41767), .Z(n41765) );
  OR U50974 ( .A(n41768), .B(n41769), .Z(n41764) );
  ANDN U50975 ( .B(n41770), .A(n41771), .Z(n41722) );
  IV U50976 ( .A(n41772), .Z(n41770) );
  ANDN U50977 ( .B(n41773), .A(n41774), .Z(n41714) );
  XOR U50978 ( .A(n41700), .B(n41775), .Z(n41712) );
  XOR U50979 ( .A(n41701), .B(n41702), .Z(n41775) );
  XOR U50980 ( .A(n41707), .B(n41776), .Z(n41702) );
  XOR U50981 ( .A(n41706), .B(n41709), .Z(n41776) );
  IV U50982 ( .A(n41708), .Z(n41709) );
  NAND U50983 ( .A(n41777), .B(n41778), .Z(n41708) );
  OR U50984 ( .A(n41779), .B(n41780), .Z(n41778) );
  OR U50985 ( .A(n41781), .B(n41782), .Z(n41777) );
  NAND U50986 ( .A(n41783), .B(n41784), .Z(n41706) );
  OR U50987 ( .A(n41785), .B(n41786), .Z(n41784) );
  OR U50988 ( .A(n41787), .B(n41788), .Z(n41783) );
  NOR U50989 ( .A(n41789), .B(n41790), .Z(n41707) );
  ANDN U50990 ( .B(n41791), .A(n41792), .Z(n41701) );
  IV U50991 ( .A(n41793), .Z(n41791) );
  XNOR U50992 ( .A(n41694), .B(n41794), .Z(n41700) );
  XNOR U50993 ( .A(n41693), .B(n41695), .Z(n41794) );
  NAND U50994 ( .A(n41795), .B(n41796), .Z(n41695) );
  OR U50995 ( .A(n41797), .B(n41798), .Z(n41796) );
  OR U50996 ( .A(n41799), .B(n41800), .Z(n41795) );
  NAND U50997 ( .A(n41801), .B(n41802), .Z(n41693) );
  OR U50998 ( .A(n41803), .B(n41804), .Z(n41802) );
  OR U50999 ( .A(n41805), .B(n41806), .Z(n41801) );
  ANDN U51000 ( .B(n41807), .A(n41808), .Z(n41694) );
  IV U51001 ( .A(n41809), .Z(n41807) );
  XNOR U51002 ( .A(n41774), .B(n41773), .Z(N61697) );
  XOR U51003 ( .A(n41793), .B(n41792), .Z(n41773) );
  XNOR U51004 ( .A(n41808), .B(n41809), .Z(n41792) );
  XNOR U51005 ( .A(n41803), .B(n41804), .Z(n41809) );
  XNOR U51006 ( .A(n41805), .B(n41806), .Z(n41804) );
  XNOR U51007 ( .A(y[2053]), .B(x[2053]), .Z(n41806) );
  XNOR U51008 ( .A(y[2054]), .B(x[2054]), .Z(n41805) );
  XNOR U51009 ( .A(y[2052]), .B(x[2052]), .Z(n41803) );
  XNOR U51010 ( .A(n41797), .B(n41798), .Z(n41808) );
  XNOR U51011 ( .A(y[2049]), .B(x[2049]), .Z(n41798) );
  XNOR U51012 ( .A(n41799), .B(n41800), .Z(n41797) );
  XNOR U51013 ( .A(y[2050]), .B(x[2050]), .Z(n41800) );
  XNOR U51014 ( .A(y[2051]), .B(x[2051]), .Z(n41799) );
  XNOR U51015 ( .A(n41790), .B(n41789), .Z(n41793) );
  XNOR U51016 ( .A(n41785), .B(n41786), .Z(n41789) );
  XNOR U51017 ( .A(y[2046]), .B(x[2046]), .Z(n41786) );
  XNOR U51018 ( .A(n41787), .B(n41788), .Z(n41785) );
  XNOR U51019 ( .A(y[2047]), .B(x[2047]), .Z(n41788) );
  XNOR U51020 ( .A(y[2048]), .B(x[2048]), .Z(n41787) );
  XNOR U51021 ( .A(n41779), .B(n41780), .Z(n41790) );
  XNOR U51022 ( .A(y[2043]), .B(x[2043]), .Z(n41780) );
  XNOR U51023 ( .A(n41781), .B(n41782), .Z(n41779) );
  XNOR U51024 ( .A(y[2044]), .B(x[2044]), .Z(n41782) );
  XNOR U51025 ( .A(y[2045]), .B(x[2045]), .Z(n41781) );
  XOR U51026 ( .A(n41755), .B(n41756), .Z(n41774) );
  XNOR U51027 ( .A(n41771), .B(n41772), .Z(n41756) );
  XNOR U51028 ( .A(n41766), .B(n41767), .Z(n41772) );
  XNOR U51029 ( .A(n41768), .B(n41769), .Z(n41767) );
  XNOR U51030 ( .A(y[2041]), .B(x[2041]), .Z(n41769) );
  XNOR U51031 ( .A(y[2042]), .B(x[2042]), .Z(n41768) );
  XNOR U51032 ( .A(y[2040]), .B(x[2040]), .Z(n41766) );
  XNOR U51033 ( .A(n41760), .B(n41761), .Z(n41771) );
  XNOR U51034 ( .A(y[2037]), .B(x[2037]), .Z(n41761) );
  XNOR U51035 ( .A(n41762), .B(n41763), .Z(n41760) );
  XNOR U51036 ( .A(y[2038]), .B(x[2038]), .Z(n41763) );
  XNOR U51037 ( .A(y[2039]), .B(x[2039]), .Z(n41762) );
  XOR U51038 ( .A(n41754), .B(n41753), .Z(n41755) );
  XNOR U51039 ( .A(n41749), .B(n41750), .Z(n41753) );
  XNOR U51040 ( .A(y[2034]), .B(x[2034]), .Z(n41750) );
  XNOR U51041 ( .A(n41751), .B(n41752), .Z(n41749) );
  XNOR U51042 ( .A(y[2035]), .B(x[2035]), .Z(n41752) );
  XNOR U51043 ( .A(y[2036]), .B(x[2036]), .Z(n41751) );
  XNOR U51044 ( .A(n41743), .B(n41744), .Z(n41754) );
  XNOR U51045 ( .A(y[2031]), .B(x[2031]), .Z(n41744) );
  XNOR U51046 ( .A(n41745), .B(n41746), .Z(n41743) );
  XNOR U51047 ( .A(y[2032]), .B(x[2032]), .Z(n41746) );
  XNOR U51048 ( .A(y[2033]), .B(x[2033]), .Z(n41745) );
  NAND U51049 ( .A(n41810), .B(n41811), .Z(N61688) );
  NANDN U51050 ( .A(n41812), .B(n41813), .Z(n41811) );
  OR U51051 ( .A(n41814), .B(n41815), .Z(n41813) );
  NAND U51052 ( .A(n41814), .B(n41815), .Z(n41810) );
  XOR U51053 ( .A(n41814), .B(n41816), .Z(N61687) );
  XNOR U51054 ( .A(n41812), .B(n41815), .Z(n41816) );
  AND U51055 ( .A(n41817), .B(n41818), .Z(n41815) );
  NANDN U51056 ( .A(n41819), .B(n41820), .Z(n41818) );
  NANDN U51057 ( .A(n41821), .B(n41822), .Z(n41820) );
  NANDN U51058 ( .A(n41822), .B(n41821), .Z(n41817) );
  NAND U51059 ( .A(n41823), .B(n41824), .Z(n41812) );
  NANDN U51060 ( .A(n41825), .B(n41826), .Z(n41824) );
  OR U51061 ( .A(n41827), .B(n41828), .Z(n41826) );
  NAND U51062 ( .A(n41828), .B(n41827), .Z(n41823) );
  AND U51063 ( .A(n41829), .B(n41830), .Z(n41814) );
  NANDN U51064 ( .A(n41831), .B(n41832), .Z(n41830) );
  NANDN U51065 ( .A(n41833), .B(n41834), .Z(n41832) );
  NANDN U51066 ( .A(n41834), .B(n41833), .Z(n41829) );
  XOR U51067 ( .A(n41828), .B(n41835), .Z(N61686) );
  XOR U51068 ( .A(n41825), .B(n41827), .Z(n41835) );
  XNOR U51069 ( .A(n41821), .B(n41836), .Z(n41827) );
  XNOR U51070 ( .A(n41819), .B(n41822), .Z(n41836) );
  NAND U51071 ( .A(n41837), .B(n41838), .Z(n41822) );
  NAND U51072 ( .A(n41839), .B(n41840), .Z(n41838) );
  OR U51073 ( .A(n41841), .B(n41842), .Z(n41839) );
  NANDN U51074 ( .A(n41843), .B(n41841), .Z(n41837) );
  IV U51075 ( .A(n41842), .Z(n41843) );
  NAND U51076 ( .A(n41844), .B(n41845), .Z(n41819) );
  NAND U51077 ( .A(n41846), .B(n41847), .Z(n41845) );
  NANDN U51078 ( .A(n41848), .B(n41849), .Z(n41846) );
  NANDN U51079 ( .A(n41849), .B(n41848), .Z(n41844) );
  AND U51080 ( .A(n41850), .B(n41851), .Z(n41821) );
  NAND U51081 ( .A(n41852), .B(n41853), .Z(n41851) );
  OR U51082 ( .A(n41854), .B(n41855), .Z(n41852) );
  NANDN U51083 ( .A(n41856), .B(n41854), .Z(n41850) );
  NAND U51084 ( .A(n41857), .B(n41858), .Z(n41825) );
  NANDN U51085 ( .A(n41859), .B(n41860), .Z(n41858) );
  OR U51086 ( .A(n41861), .B(n41862), .Z(n41860) );
  NANDN U51087 ( .A(n41863), .B(n41861), .Z(n41857) );
  IV U51088 ( .A(n41862), .Z(n41863) );
  XNOR U51089 ( .A(n41833), .B(n41864), .Z(n41828) );
  XNOR U51090 ( .A(n41831), .B(n41834), .Z(n41864) );
  NAND U51091 ( .A(n41865), .B(n41866), .Z(n41834) );
  NAND U51092 ( .A(n41867), .B(n41868), .Z(n41866) );
  OR U51093 ( .A(n41869), .B(n41870), .Z(n41867) );
  NANDN U51094 ( .A(n41871), .B(n41869), .Z(n41865) );
  IV U51095 ( .A(n41870), .Z(n41871) );
  NAND U51096 ( .A(n41872), .B(n41873), .Z(n41831) );
  NAND U51097 ( .A(n41874), .B(n41875), .Z(n41873) );
  NANDN U51098 ( .A(n41876), .B(n41877), .Z(n41874) );
  NANDN U51099 ( .A(n41877), .B(n41876), .Z(n41872) );
  AND U51100 ( .A(n41878), .B(n41879), .Z(n41833) );
  NAND U51101 ( .A(n41880), .B(n41881), .Z(n41879) );
  OR U51102 ( .A(n41882), .B(n41883), .Z(n41880) );
  NANDN U51103 ( .A(n41884), .B(n41882), .Z(n41878) );
  XNOR U51104 ( .A(n41859), .B(n41885), .Z(N61685) );
  XOR U51105 ( .A(n41861), .B(n41862), .Z(n41885) );
  XNOR U51106 ( .A(n41875), .B(n41886), .Z(n41862) );
  XOR U51107 ( .A(n41876), .B(n41877), .Z(n41886) );
  XOR U51108 ( .A(n41882), .B(n41887), .Z(n41877) );
  XOR U51109 ( .A(n41881), .B(n41884), .Z(n41887) );
  IV U51110 ( .A(n41883), .Z(n41884) );
  NAND U51111 ( .A(n41888), .B(n41889), .Z(n41883) );
  OR U51112 ( .A(n41890), .B(n41891), .Z(n41889) );
  OR U51113 ( .A(n41892), .B(n41893), .Z(n41888) );
  NAND U51114 ( .A(n41894), .B(n41895), .Z(n41881) );
  OR U51115 ( .A(n41896), .B(n41897), .Z(n41895) );
  OR U51116 ( .A(n41898), .B(n41899), .Z(n41894) );
  NOR U51117 ( .A(n41900), .B(n41901), .Z(n41882) );
  ANDN U51118 ( .B(n41902), .A(n41903), .Z(n41876) );
  XNOR U51119 ( .A(n41869), .B(n41904), .Z(n41875) );
  XNOR U51120 ( .A(n41868), .B(n41870), .Z(n41904) );
  NAND U51121 ( .A(n41905), .B(n41906), .Z(n41870) );
  OR U51122 ( .A(n41907), .B(n41908), .Z(n41906) );
  OR U51123 ( .A(n41909), .B(n41910), .Z(n41905) );
  NAND U51124 ( .A(n41911), .B(n41912), .Z(n41868) );
  OR U51125 ( .A(n41913), .B(n41914), .Z(n41912) );
  OR U51126 ( .A(n41915), .B(n41916), .Z(n41911) );
  ANDN U51127 ( .B(n41917), .A(n41918), .Z(n41869) );
  IV U51128 ( .A(n41919), .Z(n41917) );
  ANDN U51129 ( .B(n41920), .A(n41921), .Z(n41861) );
  XOR U51130 ( .A(n41847), .B(n41922), .Z(n41859) );
  XOR U51131 ( .A(n41848), .B(n41849), .Z(n41922) );
  XOR U51132 ( .A(n41854), .B(n41923), .Z(n41849) );
  XOR U51133 ( .A(n41853), .B(n41856), .Z(n41923) );
  IV U51134 ( .A(n41855), .Z(n41856) );
  NAND U51135 ( .A(n41924), .B(n41925), .Z(n41855) );
  OR U51136 ( .A(n41926), .B(n41927), .Z(n41925) );
  OR U51137 ( .A(n41928), .B(n41929), .Z(n41924) );
  NAND U51138 ( .A(n41930), .B(n41931), .Z(n41853) );
  OR U51139 ( .A(n41932), .B(n41933), .Z(n41931) );
  OR U51140 ( .A(n41934), .B(n41935), .Z(n41930) );
  NOR U51141 ( .A(n41936), .B(n41937), .Z(n41854) );
  ANDN U51142 ( .B(n41938), .A(n41939), .Z(n41848) );
  IV U51143 ( .A(n41940), .Z(n41938) );
  XNOR U51144 ( .A(n41841), .B(n41941), .Z(n41847) );
  XNOR U51145 ( .A(n41840), .B(n41842), .Z(n41941) );
  NAND U51146 ( .A(n41942), .B(n41943), .Z(n41842) );
  OR U51147 ( .A(n41944), .B(n41945), .Z(n41943) );
  OR U51148 ( .A(n41946), .B(n41947), .Z(n41942) );
  NAND U51149 ( .A(n41948), .B(n41949), .Z(n41840) );
  OR U51150 ( .A(n41950), .B(n41951), .Z(n41949) );
  OR U51151 ( .A(n41952), .B(n41953), .Z(n41948) );
  ANDN U51152 ( .B(n41954), .A(n41955), .Z(n41841) );
  IV U51153 ( .A(n41956), .Z(n41954) );
  XNOR U51154 ( .A(n41921), .B(n41920), .Z(N61684) );
  XOR U51155 ( .A(n41940), .B(n41939), .Z(n41920) );
  XNOR U51156 ( .A(n41955), .B(n41956), .Z(n41939) );
  XNOR U51157 ( .A(n41950), .B(n41951), .Z(n41956) );
  XNOR U51158 ( .A(n41952), .B(n41953), .Z(n41951) );
  XNOR U51159 ( .A(y[2029]), .B(x[2029]), .Z(n41953) );
  XNOR U51160 ( .A(y[2030]), .B(x[2030]), .Z(n41952) );
  XNOR U51161 ( .A(y[2028]), .B(x[2028]), .Z(n41950) );
  XNOR U51162 ( .A(n41944), .B(n41945), .Z(n41955) );
  XNOR U51163 ( .A(y[2025]), .B(x[2025]), .Z(n41945) );
  XNOR U51164 ( .A(n41946), .B(n41947), .Z(n41944) );
  XNOR U51165 ( .A(y[2026]), .B(x[2026]), .Z(n41947) );
  XNOR U51166 ( .A(y[2027]), .B(x[2027]), .Z(n41946) );
  XNOR U51167 ( .A(n41937), .B(n41936), .Z(n41940) );
  XNOR U51168 ( .A(n41932), .B(n41933), .Z(n41936) );
  XNOR U51169 ( .A(y[2022]), .B(x[2022]), .Z(n41933) );
  XNOR U51170 ( .A(n41934), .B(n41935), .Z(n41932) );
  XNOR U51171 ( .A(y[2023]), .B(x[2023]), .Z(n41935) );
  XNOR U51172 ( .A(y[2024]), .B(x[2024]), .Z(n41934) );
  XNOR U51173 ( .A(n41926), .B(n41927), .Z(n41937) );
  XNOR U51174 ( .A(y[2019]), .B(x[2019]), .Z(n41927) );
  XNOR U51175 ( .A(n41928), .B(n41929), .Z(n41926) );
  XNOR U51176 ( .A(y[2020]), .B(x[2020]), .Z(n41929) );
  XNOR U51177 ( .A(y[2021]), .B(x[2021]), .Z(n41928) );
  XOR U51178 ( .A(n41902), .B(n41903), .Z(n41921) );
  XNOR U51179 ( .A(n41918), .B(n41919), .Z(n41903) );
  XNOR U51180 ( .A(n41913), .B(n41914), .Z(n41919) );
  XNOR U51181 ( .A(n41915), .B(n41916), .Z(n41914) );
  XNOR U51182 ( .A(y[2017]), .B(x[2017]), .Z(n41916) );
  XNOR U51183 ( .A(y[2018]), .B(x[2018]), .Z(n41915) );
  XNOR U51184 ( .A(y[2016]), .B(x[2016]), .Z(n41913) );
  XNOR U51185 ( .A(n41907), .B(n41908), .Z(n41918) );
  XNOR U51186 ( .A(y[2013]), .B(x[2013]), .Z(n41908) );
  XNOR U51187 ( .A(n41909), .B(n41910), .Z(n41907) );
  XNOR U51188 ( .A(y[2014]), .B(x[2014]), .Z(n41910) );
  XNOR U51189 ( .A(y[2015]), .B(x[2015]), .Z(n41909) );
  XOR U51190 ( .A(n41901), .B(n41900), .Z(n41902) );
  XNOR U51191 ( .A(n41896), .B(n41897), .Z(n41900) );
  XNOR U51192 ( .A(y[2010]), .B(x[2010]), .Z(n41897) );
  XNOR U51193 ( .A(n41898), .B(n41899), .Z(n41896) );
  XNOR U51194 ( .A(y[2011]), .B(x[2011]), .Z(n41899) );
  XNOR U51195 ( .A(y[2012]), .B(x[2012]), .Z(n41898) );
  XNOR U51196 ( .A(n41890), .B(n41891), .Z(n41901) );
  XNOR U51197 ( .A(y[2007]), .B(x[2007]), .Z(n41891) );
  XNOR U51198 ( .A(n41892), .B(n41893), .Z(n41890) );
  XNOR U51199 ( .A(y[2008]), .B(x[2008]), .Z(n41893) );
  XNOR U51200 ( .A(y[2009]), .B(x[2009]), .Z(n41892) );
  NAND U51201 ( .A(n41957), .B(n41958), .Z(N61675) );
  NANDN U51202 ( .A(n41959), .B(n41960), .Z(n41958) );
  OR U51203 ( .A(n41961), .B(n41962), .Z(n41960) );
  NAND U51204 ( .A(n41961), .B(n41962), .Z(n41957) );
  XOR U51205 ( .A(n41961), .B(n41963), .Z(N61674) );
  XNOR U51206 ( .A(n41959), .B(n41962), .Z(n41963) );
  AND U51207 ( .A(n41964), .B(n41965), .Z(n41962) );
  NANDN U51208 ( .A(n41966), .B(n41967), .Z(n41965) );
  NANDN U51209 ( .A(n41968), .B(n41969), .Z(n41967) );
  NANDN U51210 ( .A(n41969), .B(n41968), .Z(n41964) );
  NAND U51211 ( .A(n41970), .B(n41971), .Z(n41959) );
  NANDN U51212 ( .A(n41972), .B(n41973), .Z(n41971) );
  OR U51213 ( .A(n41974), .B(n41975), .Z(n41973) );
  NAND U51214 ( .A(n41975), .B(n41974), .Z(n41970) );
  AND U51215 ( .A(n41976), .B(n41977), .Z(n41961) );
  NANDN U51216 ( .A(n41978), .B(n41979), .Z(n41977) );
  NANDN U51217 ( .A(n41980), .B(n41981), .Z(n41979) );
  NANDN U51218 ( .A(n41981), .B(n41980), .Z(n41976) );
  XOR U51219 ( .A(n41975), .B(n41982), .Z(N61673) );
  XOR U51220 ( .A(n41972), .B(n41974), .Z(n41982) );
  XNOR U51221 ( .A(n41968), .B(n41983), .Z(n41974) );
  XNOR U51222 ( .A(n41966), .B(n41969), .Z(n41983) );
  NAND U51223 ( .A(n41984), .B(n41985), .Z(n41969) );
  NAND U51224 ( .A(n41986), .B(n41987), .Z(n41985) );
  OR U51225 ( .A(n41988), .B(n41989), .Z(n41986) );
  NANDN U51226 ( .A(n41990), .B(n41988), .Z(n41984) );
  IV U51227 ( .A(n41989), .Z(n41990) );
  NAND U51228 ( .A(n41991), .B(n41992), .Z(n41966) );
  NAND U51229 ( .A(n41993), .B(n41994), .Z(n41992) );
  NANDN U51230 ( .A(n41995), .B(n41996), .Z(n41993) );
  NANDN U51231 ( .A(n41996), .B(n41995), .Z(n41991) );
  AND U51232 ( .A(n41997), .B(n41998), .Z(n41968) );
  NAND U51233 ( .A(n41999), .B(n42000), .Z(n41998) );
  OR U51234 ( .A(n42001), .B(n42002), .Z(n41999) );
  NANDN U51235 ( .A(n42003), .B(n42001), .Z(n41997) );
  NAND U51236 ( .A(n42004), .B(n42005), .Z(n41972) );
  NANDN U51237 ( .A(n42006), .B(n42007), .Z(n42005) );
  OR U51238 ( .A(n42008), .B(n42009), .Z(n42007) );
  NANDN U51239 ( .A(n42010), .B(n42008), .Z(n42004) );
  IV U51240 ( .A(n42009), .Z(n42010) );
  XNOR U51241 ( .A(n41980), .B(n42011), .Z(n41975) );
  XNOR U51242 ( .A(n41978), .B(n41981), .Z(n42011) );
  NAND U51243 ( .A(n42012), .B(n42013), .Z(n41981) );
  NAND U51244 ( .A(n42014), .B(n42015), .Z(n42013) );
  OR U51245 ( .A(n42016), .B(n42017), .Z(n42014) );
  NANDN U51246 ( .A(n42018), .B(n42016), .Z(n42012) );
  IV U51247 ( .A(n42017), .Z(n42018) );
  NAND U51248 ( .A(n42019), .B(n42020), .Z(n41978) );
  NAND U51249 ( .A(n42021), .B(n42022), .Z(n42020) );
  NANDN U51250 ( .A(n42023), .B(n42024), .Z(n42021) );
  NANDN U51251 ( .A(n42024), .B(n42023), .Z(n42019) );
  AND U51252 ( .A(n42025), .B(n42026), .Z(n41980) );
  NAND U51253 ( .A(n42027), .B(n42028), .Z(n42026) );
  OR U51254 ( .A(n42029), .B(n42030), .Z(n42027) );
  NANDN U51255 ( .A(n42031), .B(n42029), .Z(n42025) );
  XNOR U51256 ( .A(n42006), .B(n42032), .Z(N61672) );
  XOR U51257 ( .A(n42008), .B(n42009), .Z(n42032) );
  XNOR U51258 ( .A(n42022), .B(n42033), .Z(n42009) );
  XOR U51259 ( .A(n42023), .B(n42024), .Z(n42033) );
  XOR U51260 ( .A(n42029), .B(n42034), .Z(n42024) );
  XOR U51261 ( .A(n42028), .B(n42031), .Z(n42034) );
  IV U51262 ( .A(n42030), .Z(n42031) );
  NAND U51263 ( .A(n42035), .B(n42036), .Z(n42030) );
  OR U51264 ( .A(n42037), .B(n42038), .Z(n42036) );
  OR U51265 ( .A(n42039), .B(n42040), .Z(n42035) );
  NAND U51266 ( .A(n42041), .B(n42042), .Z(n42028) );
  OR U51267 ( .A(n42043), .B(n42044), .Z(n42042) );
  OR U51268 ( .A(n42045), .B(n42046), .Z(n42041) );
  NOR U51269 ( .A(n42047), .B(n42048), .Z(n42029) );
  ANDN U51270 ( .B(n42049), .A(n42050), .Z(n42023) );
  XNOR U51271 ( .A(n42016), .B(n42051), .Z(n42022) );
  XNOR U51272 ( .A(n42015), .B(n42017), .Z(n42051) );
  NAND U51273 ( .A(n42052), .B(n42053), .Z(n42017) );
  OR U51274 ( .A(n42054), .B(n42055), .Z(n42053) );
  OR U51275 ( .A(n42056), .B(n42057), .Z(n42052) );
  NAND U51276 ( .A(n42058), .B(n42059), .Z(n42015) );
  OR U51277 ( .A(n42060), .B(n42061), .Z(n42059) );
  OR U51278 ( .A(n42062), .B(n42063), .Z(n42058) );
  ANDN U51279 ( .B(n42064), .A(n42065), .Z(n42016) );
  IV U51280 ( .A(n42066), .Z(n42064) );
  ANDN U51281 ( .B(n42067), .A(n42068), .Z(n42008) );
  XOR U51282 ( .A(n41994), .B(n42069), .Z(n42006) );
  XOR U51283 ( .A(n41995), .B(n41996), .Z(n42069) );
  XOR U51284 ( .A(n42001), .B(n42070), .Z(n41996) );
  XOR U51285 ( .A(n42000), .B(n42003), .Z(n42070) );
  IV U51286 ( .A(n42002), .Z(n42003) );
  NAND U51287 ( .A(n42071), .B(n42072), .Z(n42002) );
  OR U51288 ( .A(n42073), .B(n42074), .Z(n42072) );
  OR U51289 ( .A(n42075), .B(n42076), .Z(n42071) );
  NAND U51290 ( .A(n42077), .B(n42078), .Z(n42000) );
  OR U51291 ( .A(n42079), .B(n42080), .Z(n42078) );
  OR U51292 ( .A(n42081), .B(n42082), .Z(n42077) );
  NOR U51293 ( .A(n42083), .B(n42084), .Z(n42001) );
  ANDN U51294 ( .B(n42085), .A(n42086), .Z(n41995) );
  IV U51295 ( .A(n42087), .Z(n42085) );
  XNOR U51296 ( .A(n41988), .B(n42088), .Z(n41994) );
  XNOR U51297 ( .A(n41987), .B(n41989), .Z(n42088) );
  NAND U51298 ( .A(n42089), .B(n42090), .Z(n41989) );
  OR U51299 ( .A(n42091), .B(n42092), .Z(n42090) );
  OR U51300 ( .A(n42093), .B(n42094), .Z(n42089) );
  NAND U51301 ( .A(n42095), .B(n42096), .Z(n41987) );
  OR U51302 ( .A(n42097), .B(n42098), .Z(n42096) );
  OR U51303 ( .A(n42099), .B(n42100), .Z(n42095) );
  ANDN U51304 ( .B(n42101), .A(n42102), .Z(n41988) );
  IV U51305 ( .A(n42103), .Z(n42101) );
  XNOR U51306 ( .A(n42068), .B(n42067), .Z(N61671) );
  XOR U51307 ( .A(n42087), .B(n42086), .Z(n42067) );
  XNOR U51308 ( .A(n42102), .B(n42103), .Z(n42086) );
  XNOR U51309 ( .A(n42097), .B(n42098), .Z(n42103) );
  XNOR U51310 ( .A(n42099), .B(n42100), .Z(n42098) );
  XNOR U51311 ( .A(y[2005]), .B(x[2005]), .Z(n42100) );
  XNOR U51312 ( .A(y[2006]), .B(x[2006]), .Z(n42099) );
  XNOR U51313 ( .A(y[2004]), .B(x[2004]), .Z(n42097) );
  XNOR U51314 ( .A(n42091), .B(n42092), .Z(n42102) );
  XNOR U51315 ( .A(y[2001]), .B(x[2001]), .Z(n42092) );
  XNOR U51316 ( .A(n42093), .B(n42094), .Z(n42091) );
  XNOR U51317 ( .A(y[2002]), .B(x[2002]), .Z(n42094) );
  XNOR U51318 ( .A(y[2003]), .B(x[2003]), .Z(n42093) );
  XNOR U51319 ( .A(n42084), .B(n42083), .Z(n42087) );
  XNOR U51320 ( .A(n42079), .B(n42080), .Z(n42083) );
  XNOR U51321 ( .A(y[1998]), .B(x[1998]), .Z(n42080) );
  XNOR U51322 ( .A(n42081), .B(n42082), .Z(n42079) );
  XNOR U51323 ( .A(y[1999]), .B(x[1999]), .Z(n42082) );
  XNOR U51324 ( .A(y[2000]), .B(x[2000]), .Z(n42081) );
  XNOR U51325 ( .A(n42073), .B(n42074), .Z(n42084) );
  XNOR U51326 ( .A(y[1995]), .B(x[1995]), .Z(n42074) );
  XNOR U51327 ( .A(n42075), .B(n42076), .Z(n42073) );
  XNOR U51328 ( .A(y[1996]), .B(x[1996]), .Z(n42076) );
  XNOR U51329 ( .A(y[1997]), .B(x[1997]), .Z(n42075) );
  XOR U51330 ( .A(n42049), .B(n42050), .Z(n42068) );
  XNOR U51331 ( .A(n42065), .B(n42066), .Z(n42050) );
  XNOR U51332 ( .A(n42060), .B(n42061), .Z(n42066) );
  XNOR U51333 ( .A(n42062), .B(n42063), .Z(n42061) );
  XNOR U51334 ( .A(y[1993]), .B(x[1993]), .Z(n42063) );
  XNOR U51335 ( .A(y[1994]), .B(x[1994]), .Z(n42062) );
  XNOR U51336 ( .A(y[1992]), .B(x[1992]), .Z(n42060) );
  XNOR U51337 ( .A(n42054), .B(n42055), .Z(n42065) );
  XNOR U51338 ( .A(y[1989]), .B(x[1989]), .Z(n42055) );
  XNOR U51339 ( .A(n42056), .B(n42057), .Z(n42054) );
  XNOR U51340 ( .A(y[1990]), .B(x[1990]), .Z(n42057) );
  XNOR U51341 ( .A(y[1991]), .B(x[1991]), .Z(n42056) );
  XOR U51342 ( .A(n42048), .B(n42047), .Z(n42049) );
  XNOR U51343 ( .A(n42043), .B(n42044), .Z(n42047) );
  XNOR U51344 ( .A(y[1986]), .B(x[1986]), .Z(n42044) );
  XNOR U51345 ( .A(n42045), .B(n42046), .Z(n42043) );
  XNOR U51346 ( .A(y[1987]), .B(x[1987]), .Z(n42046) );
  XNOR U51347 ( .A(y[1988]), .B(x[1988]), .Z(n42045) );
  XNOR U51348 ( .A(n42037), .B(n42038), .Z(n42048) );
  XNOR U51349 ( .A(y[1983]), .B(x[1983]), .Z(n42038) );
  XNOR U51350 ( .A(n42039), .B(n42040), .Z(n42037) );
  XNOR U51351 ( .A(y[1984]), .B(x[1984]), .Z(n42040) );
  XNOR U51352 ( .A(y[1985]), .B(x[1985]), .Z(n42039) );
  NAND U51353 ( .A(n42104), .B(n42105), .Z(N61662) );
  NANDN U51354 ( .A(n42106), .B(n42107), .Z(n42105) );
  OR U51355 ( .A(n42108), .B(n42109), .Z(n42107) );
  NAND U51356 ( .A(n42108), .B(n42109), .Z(n42104) );
  XOR U51357 ( .A(n42108), .B(n42110), .Z(N61661) );
  XNOR U51358 ( .A(n42106), .B(n42109), .Z(n42110) );
  AND U51359 ( .A(n42111), .B(n42112), .Z(n42109) );
  NANDN U51360 ( .A(n42113), .B(n42114), .Z(n42112) );
  NANDN U51361 ( .A(n42115), .B(n42116), .Z(n42114) );
  NANDN U51362 ( .A(n42116), .B(n42115), .Z(n42111) );
  NAND U51363 ( .A(n42117), .B(n42118), .Z(n42106) );
  NANDN U51364 ( .A(n42119), .B(n42120), .Z(n42118) );
  OR U51365 ( .A(n42121), .B(n42122), .Z(n42120) );
  NAND U51366 ( .A(n42122), .B(n42121), .Z(n42117) );
  AND U51367 ( .A(n42123), .B(n42124), .Z(n42108) );
  NANDN U51368 ( .A(n42125), .B(n42126), .Z(n42124) );
  NANDN U51369 ( .A(n42127), .B(n42128), .Z(n42126) );
  NANDN U51370 ( .A(n42128), .B(n42127), .Z(n42123) );
  XOR U51371 ( .A(n42122), .B(n42129), .Z(N61660) );
  XOR U51372 ( .A(n42119), .B(n42121), .Z(n42129) );
  XNOR U51373 ( .A(n42115), .B(n42130), .Z(n42121) );
  XNOR U51374 ( .A(n42113), .B(n42116), .Z(n42130) );
  NAND U51375 ( .A(n42131), .B(n42132), .Z(n42116) );
  NAND U51376 ( .A(n42133), .B(n42134), .Z(n42132) );
  OR U51377 ( .A(n42135), .B(n42136), .Z(n42133) );
  NANDN U51378 ( .A(n42137), .B(n42135), .Z(n42131) );
  IV U51379 ( .A(n42136), .Z(n42137) );
  NAND U51380 ( .A(n42138), .B(n42139), .Z(n42113) );
  NAND U51381 ( .A(n42140), .B(n42141), .Z(n42139) );
  NANDN U51382 ( .A(n42142), .B(n42143), .Z(n42140) );
  NANDN U51383 ( .A(n42143), .B(n42142), .Z(n42138) );
  AND U51384 ( .A(n42144), .B(n42145), .Z(n42115) );
  NAND U51385 ( .A(n42146), .B(n42147), .Z(n42145) );
  OR U51386 ( .A(n42148), .B(n42149), .Z(n42146) );
  NANDN U51387 ( .A(n42150), .B(n42148), .Z(n42144) );
  NAND U51388 ( .A(n42151), .B(n42152), .Z(n42119) );
  NANDN U51389 ( .A(n42153), .B(n42154), .Z(n42152) );
  OR U51390 ( .A(n42155), .B(n42156), .Z(n42154) );
  NANDN U51391 ( .A(n42157), .B(n42155), .Z(n42151) );
  IV U51392 ( .A(n42156), .Z(n42157) );
  XNOR U51393 ( .A(n42127), .B(n42158), .Z(n42122) );
  XNOR U51394 ( .A(n42125), .B(n42128), .Z(n42158) );
  NAND U51395 ( .A(n42159), .B(n42160), .Z(n42128) );
  NAND U51396 ( .A(n42161), .B(n42162), .Z(n42160) );
  OR U51397 ( .A(n42163), .B(n42164), .Z(n42161) );
  NANDN U51398 ( .A(n42165), .B(n42163), .Z(n42159) );
  IV U51399 ( .A(n42164), .Z(n42165) );
  NAND U51400 ( .A(n42166), .B(n42167), .Z(n42125) );
  NAND U51401 ( .A(n42168), .B(n42169), .Z(n42167) );
  NANDN U51402 ( .A(n42170), .B(n42171), .Z(n42168) );
  NANDN U51403 ( .A(n42171), .B(n42170), .Z(n42166) );
  AND U51404 ( .A(n42172), .B(n42173), .Z(n42127) );
  NAND U51405 ( .A(n42174), .B(n42175), .Z(n42173) );
  OR U51406 ( .A(n42176), .B(n42177), .Z(n42174) );
  NANDN U51407 ( .A(n42178), .B(n42176), .Z(n42172) );
  XNOR U51408 ( .A(n42153), .B(n42179), .Z(N61659) );
  XOR U51409 ( .A(n42155), .B(n42156), .Z(n42179) );
  XNOR U51410 ( .A(n42169), .B(n42180), .Z(n42156) );
  XOR U51411 ( .A(n42170), .B(n42171), .Z(n42180) );
  XOR U51412 ( .A(n42176), .B(n42181), .Z(n42171) );
  XOR U51413 ( .A(n42175), .B(n42178), .Z(n42181) );
  IV U51414 ( .A(n42177), .Z(n42178) );
  NAND U51415 ( .A(n42182), .B(n42183), .Z(n42177) );
  OR U51416 ( .A(n42184), .B(n42185), .Z(n42183) );
  OR U51417 ( .A(n42186), .B(n42187), .Z(n42182) );
  NAND U51418 ( .A(n42188), .B(n42189), .Z(n42175) );
  OR U51419 ( .A(n42190), .B(n42191), .Z(n42189) );
  OR U51420 ( .A(n42192), .B(n42193), .Z(n42188) );
  NOR U51421 ( .A(n42194), .B(n42195), .Z(n42176) );
  ANDN U51422 ( .B(n42196), .A(n42197), .Z(n42170) );
  XNOR U51423 ( .A(n42163), .B(n42198), .Z(n42169) );
  XNOR U51424 ( .A(n42162), .B(n42164), .Z(n42198) );
  NAND U51425 ( .A(n42199), .B(n42200), .Z(n42164) );
  OR U51426 ( .A(n42201), .B(n42202), .Z(n42200) );
  OR U51427 ( .A(n42203), .B(n42204), .Z(n42199) );
  NAND U51428 ( .A(n42205), .B(n42206), .Z(n42162) );
  OR U51429 ( .A(n42207), .B(n42208), .Z(n42206) );
  OR U51430 ( .A(n42209), .B(n42210), .Z(n42205) );
  ANDN U51431 ( .B(n42211), .A(n42212), .Z(n42163) );
  IV U51432 ( .A(n42213), .Z(n42211) );
  ANDN U51433 ( .B(n42214), .A(n42215), .Z(n42155) );
  XOR U51434 ( .A(n42141), .B(n42216), .Z(n42153) );
  XOR U51435 ( .A(n42142), .B(n42143), .Z(n42216) );
  XOR U51436 ( .A(n42148), .B(n42217), .Z(n42143) );
  XOR U51437 ( .A(n42147), .B(n42150), .Z(n42217) );
  IV U51438 ( .A(n42149), .Z(n42150) );
  NAND U51439 ( .A(n42218), .B(n42219), .Z(n42149) );
  OR U51440 ( .A(n42220), .B(n42221), .Z(n42219) );
  OR U51441 ( .A(n42222), .B(n42223), .Z(n42218) );
  NAND U51442 ( .A(n42224), .B(n42225), .Z(n42147) );
  OR U51443 ( .A(n42226), .B(n42227), .Z(n42225) );
  OR U51444 ( .A(n42228), .B(n42229), .Z(n42224) );
  NOR U51445 ( .A(n42230), .B(n42231), .Z(n42148) );
  ANDN U51446 ( .B(n42232), .A(n42233), .Z(n42142) );
  IV U51447 ( .A(n42234), .Z(n42232) );
  XNOR U51448 ( .A(n42135), .B(n42235), .Z(n42141) );
  XNOR U51449 ( .A(n42134), .B(n42136), .Z(n42235) );
  NAND U51450 ( .A(n42236), .B(n42237), .Z(n42136) );
  OR U51451 ( .A(n42238), .B(n42239), .Z(n42237) );
  OR U51452 ( .A(n42240), .B(n42241), .Z(n42236) );
  NAND U51453 ( .A(n42242), .B(n42243), .Z(n42134) );
  OR U51454 ( .A(n42244), .B(n42245), .Z(n42243) );
  OR U51455 ( .A(n42246), .B(n42247), .Z(n42242) );
  ANDN U51456 ( .B(n42248), .A(n42249), .Z(n42135) );
  IV U51457 ( .A(n42250), .Z(n42248) );
  XNOR U51458 ( .A(n42215), .B(n42214), .Z(N61658) );
  XOR U51459 ( .A(n42234), .B(n42233), .Z(n42214) );
  XNOR U51460 ( .A(n42249), .B(n42250), .Z(n42233) );
  XNOR U51461 ( .A(n42244), .B(n42245), .Z(n42250) );
  XNOR U51462 ( .A(n42246), .B(n42247), .Z(n42245) );
  XNOR U51463 ( .A(y[1981]), .B(x[1981]), .Z(n42247) );
  XNOR U51464 ( .A(y[1982]), .B(x[1982]), .Z(n42246) );
  XNOR U51465 ( .A(y[1980]), .B(x[1980]), .Z(n42244) );
  XNOR U51466 ( .A(n42238), .B(n42239), .Z(n42249) );
  XNOR U51467 ( .A(y[1977]), .B(x[1977]), .Z(n42239) );
  XNOR U51468 ( .A(n42240), .B(n42241), .Z(n42238) );
  XNOR U51469 ( .A(y[1978]), .B(x[1978]), .Z(n42241) );
  XNOR U51470 ( .A(y[1979]), .B(x[1979]), .Z(n42240) );
  XNOR U51471 ( .A(n42231), .B(n42230), .Z(n42234) );
  XNOR U51472 ( .A(n42226), .B(n42227), .Z(n42230) );
  XNOR U51473 ( .A(y[1974]), .B(x[1974]), .Z(n42227) );
  XNOR U51474 ( .A(n42228), .B(n42229), .Z(n42226) );
  XNOR U51475 ( .A(y[1975]), .B(x[1975]), .Z(n42229) );
  XNOR U51476 ( .A(y[1976]), .B(x[1976]), .Z(n42228) );
  XNOR U51477 ( .A(n42220), .B(n42221), .Z(n42231) );
  XNOR U51478 ( .A(y[1971]), .B(x[1971]), .Z(n42221) );
  XNOR U51479 ( .A(n42222), .B(n42223), .Z(n42220) );
  XNOR U51480 ( .A(y[1972]), .B(x[1972]), .Z(n42223) );
  XNOR U51481 ( .A(y[1973]), .B(x[1973]), .Z(n42222) );
  XOR U51482 ( .A(n42196), .B(n42197), .Z(n42215) );
  XNOR U51483 ( .A(n42212), .B(n42213), .Z(n42197) );
  XNOR U51484 ( .A(n42207), .B(n42208), .Z(n42213) );
  XNOR U51485 ( .A(n42209), .B(n42210), .Z(n42208) );
  XNOR U51486 ( .A(y[1969]), .B(x[1969]), .Z(n42210) );
  XNOR U51487 ( .A(y[1970]), .B(x[1970]), .Z(n42209) );
  XNOR U51488 ( .A(y[1968]), .B(x[1968]), .Z(n42207) );
  XNOR U51489 ( .A(n42201), .B(n42202), .Z(n42212) );
  XNOR U51490 ( .A(y[1965]), .B(x[1965]), .Z(n42202) );
  XNOR U51491 ( .A(n42203), .B(n42204), .Z(n42201) );
  XNOR U51492 ( .A(y[1966]), .B(x[1966]), .Z(n42204) );
  XNOR U51493 ( .A(y[1967]), .B(x[1967]), .Z(n42203) );
  XOR U51494 ( .A(n42195), .B(n42194), .Z(n42196) );
  XNOR U51495 ( .A(n42190), .B(n42191), .Z(n42194) );
  XNOR U51496 ( .A(y[1962]), .B(x[1962]), .Z(n42191) );
  XNOR U51497 ( .A(n42192), .B(n42193), .Z(n42190) );
  XNOR U51498 ( .A(y[1963]), .B(x[1963]), .Z(n42193) );
  XNOR U51499 ( .A(y[1964]), .B(x[1964]), .Z(n42192) );
  XNOR U51500 ( .A(n42184), .B(n42185), .Z(n42195) );
  XNOR U51501 ( .A(y[1959]), .B(x[1959]), .Z(n42185) );
  XNOR U51502 ( .A(n42186), .B(n42187), .Z(n42184) );
  XNOR U51503 ( .A(y[1960]), .B(x[1960]), .Z(n42187) );
  XNOR U51504 ( .A(y[1961]), .B(x[1961]), .Z(n42186) );
  NAND U51505 ( .A(n42251), .B(n42252), .Z(N61649) );
  NANDN U51506 ( .A(n42253), .B(n42254), .Z(n42252) );
  OR U51507 ( .A(n42255), .B(n42256), .Z(n42254) );
  NAND U51508 ( .A(n42255), .B(n42256), .Z(n42251) );
  XOR U51509 ( .A(n42255), .B(n42257), .Z(N61648) );
  XNOR U51510 ( .A(n42253), .B(n42256), .Z(n42257) );
  AND U51511 ( .A(n42258), .B(n42259), .Z(n42256) );
  NANDN U51512 ( .A(n42260), .B(n42261), .Z(n42259) );
  NANDN U51513 ( .A(n42262), .B(n42263), .Z(n42261) );
  NANDN U51514 ( .A(n42263), .B(n42262), .Z(n42258) );
  NAND U51515 ( .A(n42264), .B(n42265), .Z(n42253) );
  NANDN U51516 ( .A(n42266), .B(n42267), .Z(n42265) );
  OR U51517 ( .A(n42268), .B(n42269), .Z(n42267) );
  NAND U51518 ( .A(n42269), .B(n42268), .Z(n42264) );
  AND U51519 ( .A(n42270), .B(n42271), .Z(n42255) );
  NANDN U51520 ( .A(n42272), .B(n42273), .Z(n42271) );
  NANDN U51521 ( .A(n42274), .B(n42275), .Z(n42273) );
  NANDN U51522 ( .A(n42275), .B(n42274), .Z(n42270) );
  XOR U51523 ( .A(n42269), .B(n42276), .Z(N61647) );
  XOR U51524 ( .A(n42266), .B(n42268), .Z(n42276) );
  XNOR U51525 ( .A(n42262), .B(n42277), .Z(n42268) );
  XNOR U51526 ( .A(n42260), .B(n42263), .Z(n42277) );
  NAND U51527 ( .A(n42278), .B(n42279), .Z(n42263) );
  NAND U51528 ( .A(n42280), .B(n42281), .Z(n42279) );
  OR U51529 ( .A(n42282), .B(n42283), .Z(n42280) );
  NANDN U51530 ( .A(n42284), .B(n42282), .Z(n42278) );
  IV U51531 ( .A(n42283), .Z(n42284) );
  NAND U51532 ( .A(n42285), .B(n42286), .Z(n42260) );
  NAND U51533 ( .A(n42287), .B(n42288), .Z(n42286) );
  NANDN U51534 ( .A(n42289), .B(n42290), .Z(n42287) );
  NANDN U51535 ( .A(n42290), .B(n42289), .Z(n42285) );
  AND U51536 ( .A(n42291), .B(n42292), .Z(n42262) );
  NAND U51537 ( .A(n42293), .B(n42294), .Z(n42292) );
  OR U51538 ( .A(n42295), .B(n42296), .Z(n42293) );
  NANDN U51539 ( .A(n42297), .B(n42295), .Z(n42291) );
  NAND U51540 ( .A(n42298), .B(n42299), .Z(n42266) );
  NANDN U51541 ( .A(n42300), .B(n42301), .Z(n42299) );
  OR U51542 ( .A(n42302), .B(n42303), .Z(n42301) );
  NANDN U51543 ( .A(n42304), .B(n42302), .Z(n42298) );
  IV U51544 ( .A(n42303), .Z(n42304) );
  XNOR U51545 ( .A(n42274), .B(n42305), .Z(n42269) );
  XNOR U51546 ( .A(n42272), .B(n42275), .Z(n42305) );
  NAND U51547 ( .A(n42306), .B(n42307), .Z(n42275) );
  NAND U51548 ( .A(n42308), .B(n42309), .Z(n42307) );
  OR U51549 ( .A(n42310), .B(n42311), .Z(n42308) );
  NANDN U51550 ( .A(n42312), .B(n42310), .Z(n42306) );
  IV U51551 ( .A(n42311), .Z(n42312) );
  NAND U51552 ( .A(n42313), .B(n42314), .Z(n42272) );
  NAND U51553 ( .A(n42315), .B(n42316), .Z(n42314) );
  NANDN U51554 ( .A(n42317), .B(n42318), .Z(n42315) );
  NANDN U51555 ( .A(n42318), .B(n42317), .Z(n42313) );
  AND U51556 ( .A(n42319), .B(n42320), .Z(n42274) );
  NAND U51557 ( .A(n42321), .B(n42322), .Z(n42320) );
  OR U51558 ( .A(n42323), .B(n42324), .Z(n42321) );
  NANDN U51559 ( .A(n42325), .B(n42323), .Z(n42319) );
  XNOR U51560 ( .A(n42300), .B(n42326), .Z(N61646) );
  XOR U51561 ( .A(n42302), .B(n42303), .Z(n42326) );
  XNOR U51562 ( .A(n42316), .B(n42327), .Z(n42303) );
  XOR U51563 ( .A(n42317), .B(n42318), .Z(n42327) );
  XOR U51564 ( .A(n42323), .B(n42328), .Z(n42318) );
  XOR U51565 ( .A(n42322), .B(n42325), .Z(n42328) );
  IV U51566 ( .A(n42324), .Z(n42325) );
  NAND U51567 ( .A(n42329), .B(n42330), .Z(n42324) );
  OR U51568 ( .A(n42331), .B(n42332), .Z(n42330) );
  OR U51569 ( .A(n42333), .B(n42334), .Z(n42329) );
  NAND U51570 ( .A(n42335), .B(n42336), .Z(n42322) );
  OR U51571 ( .A(n42337), .B(n42338), .Z(n42336) );
  OR U51572 ( .A(n42339), .B(n42340), .Z(n42335) );
  NOR U51573 ( .A(n42341), .B(n42342), .Z(n42323) );
  ANDN U51574 ( .B(n42343), .A(n42344), .Z(n42317) );
  XNOR U51575 ( .A(n42310), .B(n42345), .Z(n42316) );
  XNOR U51576 ( .A(n42309), .B(n42311), .Z(n42345) );
  NAND U51577 ( .A(n42346), .B(n42347), .Z(n42311) );
  OR U51578 ( .A(n42348), .B(n42349), .Z(n42347) );
  OR U51579 ( .A(n42350), .B(n42351), .Z(n42346) );
  NAND U51580 ( .A(n42352), .B(n42353), .Z(n42309) );
  OR U51581 ( .A(n42354), .B(n42355), .Z(n42353) );
  OR U51582 ( .A(n42356), .B(n42357), .Z(n42352) );
  ANDN U51583 ( .B(n42358), .A(n42359), .Z(n42310) );
  IV U51584 ( .A(n42360), .Z(n42358) );
  ANDN U51585 ( .B(n42361), .A(n42362), .Z(n42302) );
  XOR U51586 ( .A(n42288), .B(n42363), .Z(n42300) );
  XOR U51587 ( .A(n42289), .B(n42290), .Z(n42363) );
  XOR U51588 ( .A(n42295), .B(n42364), .Z(n42290) );
  XOR U51589 ( .A(n42294), .B(n42297), .Z(n42364) );
  IV U51590 ( .A(n42296), .Z(n42297) );
  NAND U51591 ( .A(n42365), .B(n42366), .Z(n42296) );
  OR U51592 ( .A(n42367), .B(n42368), .Z(n42366) );
  OR U51593 ( .A(n42369), .B(n42370), .Z(n42365) );
  NAND U51594 ( .A(n42371), .B(n42372), .Z(n42294) );
  OR U51595 ( .A(n42373), .B(n42374), .Z(n42372) );
  OR U51596 ( .A(n42375), .B(n42376), .Z(n42371) );
  NOR U51597 ( .A(n42377), .B(n42378), .Z(n42295) );
  ANDN U51598 ( .B(n42379), .A(n42380), .Z(n42289) );
  IV U51599 ( .A(n42381), .Z(n42379) );
  XNOR U51600 ( .A(n42282), .B(n42382), .Z(n42288) );
  XNOR U51601 ( .A(n42281), .B(n42283), .Z(n42382) );
  NAND U51602 ( .A(n42383), .B(n42384), .Z(n42283) );
  OR U51603 ( .A(n42385), .B(n42386), .Z(n42384) );
  OR U51604 ( .A(n42387), .B(n42388), .Z(n42383) );
  NAND U51605 ( .A(n42389), .B(n42390), .Z(n42281) );
  OR U51606 ( .A(n42391), .B(n42392), .Z(n42390) );
  OR U51607 ( .A(n42393), .B(n42394), .Z(n42389) );
  ANDN U51608 ( .B(n42395), .A(n42396), .Z(n42282) );
  IV U51609 ( .A(n42397), .Z(n42395) );
  XNOR U51610 ( .A(n42362), .B(n42361), .Z(N61645) );
  XOR U51611 ( .A(n42381), .B(n42380), .Z(n42361) );
  XNOR U51612 ( .A(n42396), .B(n42397), .Z(n42380) );
  XNOR U51613 ( .A(n42391), .B(n42392), .Z(n42397) );
  XNOR U51614 ( .A(n42393), .B(n42394), .Z(n42392) );
  XNOR U51615 ( .A(y[1957]), .B(x[1957]), .Z(n42394) );
  XNOR U51616 ( .A(y[1958]), .B(x[1958]), .Z(n42393) );
  XNOR U51617 ( .A(y[1956]), .B(x[1956]), .Z(n42391) );
  XNOR U51618 ( .A(n42385), .B(n42386), .Z(n42396) );
  XNOR U51619 ( .A(y[1953]), .B(x[1953]), .Z(n42386) );
  XNOR U51620 ( .A(n42387), .B(n42388), .Z(n42385) );
  XNOR U51621 ( .A(y[1954]), .B(x[1954]), .Z(n42388) );
  XNOR U51622 ( .A(y[1955]), .B(x[1955]), .Z(n42387) );
  XNOR U51623 ( .A(n42378), .B(n42377), .Z(n42381) );
  XNOR U51624 ( .A(n42373), .B(n42374), .Z(n42377) );
  XNOR U51625 ( .A(y[1950]), .B(x[1950]), .Z(n42374) );
  XNOR U51626 ( .A(n42375), .B(n42376), .Z(n42373) );
  XNOR U51627 ( .A(y[1951]), .B(x[1951]), .Z(n42376) );
  XNOR U51628 ( .A(y[1952]), .B(x[1952]), .Z(n42375) );
  XNOR U51629 ( .A(n42367), .B(n42368), .Z(n42378) );
  XNOR U51630 ( .A(y[1947]), .B(x[1947]), .Z(n42368) );
  XNOR U51631 ( .A(n42369), .B(n42370), .Z(n42367) );
  XNOR U51632 ( .A(y[1948]), .B(x[1948]), .Z(n42370) );
  XNOR U51633 ( .A(y[1949]), .B(x[1949]), .Z(n42369) );
  XOR U51634 ( .A(n42343), .B(n42344), .Z(n42362) );
  XNOR U51635 ( .A(n42359), .B(n42360), .Z(n42344) );
  XNOR U51636 ( .A(n42354), .B(n42355), .Z(n42360) );
  XNOR U51637 ( .A(n42356), .B(n42357), .Z(n42355) );
  XNOR U51638 ( .A(y[1945]), .B(x[1945]), .Z(n42357) );
  XNOR U51639 ( .A(y[1946]), .B(x[1946]), .Z(n42356) );
  XNOR U51640 ( .A(y[1944]), .B(x[1944]), .Z(n42354) );
  XNOR U51641 ( .A(n42348), .B(n42349), .Z(n42359) );
  XNOR U51642 ( .A(y[1941]), .B(x[1941]), .Z(n42349) );
  XNOR U51643 ( .A(n42350), .B(n42351), .Z(n42348) );
  XNOR U51644 ( .A(y[1942]), .B(x[1942]), .Z(n42351) );
  XNOR U51645 ( .A(y[1943]), .B(x[1943]), .Z(n42350) );
  XOR U51646 ( .A(n42342), .B(n42341), .Z(n42343) );
  XNOR U51647 ( .A(n42337), .B(n42338), .Z(n42341) );
  XNOR U51648 ( .A(y[1938]), .B(x[1938]), .Z(n42338) );
  XNOR U51649 ( .A(n42339), .B(n42340), .Z(n42337) );
  XNOR U51650 ( .A(y[1939]), .B(x[1939]), .Z(n42340) );
  XNOR U51651 ( .A(y[1940]), .B(x[1940]), .Z(n42339) );
  XNOR U51652 ( .A(n42331), .B(n42332), .Z(n42342) );
  XNOR U51653 ( .A(y[1935]), .B(x[1935]), .Z(n42332) );
  XNOR U51654 ( .A(n42333), .B(n42334), .Z(n42331) );
  XNOR U51655 ( .A(y[1936]), .B(x[1936]), .Z(n42334) );
  XNOR U51656 ( .A(y[1937]), .B(x[1937]), .Z(n42333) );
  NAND U51657 ( .A(n42398), .B(n42399), .Z(N61636) );
  NANDN U51658 ( .A(n42400), .B(n42401), .Z(n42399) );
  OR U51659 ( .A(n42402), .B(n42403), .Z(n42401) );
  NAND U51660 ( .A(n42402), .B(n42403), .Z(n42398) );
  XOR U51661 ( .A(n42402), .B(n42404), .Z(N61635) );
  XNOR U51662 ( .A(n42400), .B(n42403), .Z(n42404) );
  AND U51663 ( .A(n42405), .B(n42406), .Z(n42403) );
  NANDN U51664 ( .A(n42407), .B(n42408), .Z(n42406) );
  NANDN U51665 ( .A(n42409), .B(n42410), .Z(n42408) );
  NANDN U51666 ( .A(n42410), .B(n42409), .Z(n42405) );
  NAND U51667 ( .A(n42411), .B(n42412), .Z(n42400) );
  NANDN U51668 ( .A(n42413), .B(n42414), .Z(n42412) );
  OR U51669 ( .A(n42415), .B(n42416), .Z(n42414) );
  NAND U51670 ( .A(n42416), .B(n42415), .Z(n42411) );
  AND U51671 ( .A(n42417), .B(n42418), .Z(n42402) );
  NANDN U51672 ( .A(n42419), .B(n42420), .Z(n42418) );
  NANDN U51673 ( .A(n42421), .B(n42422), .Z(n42420) );
  NANDN U51674 ( .A(n42422), .B(n42421), .Z(n42417) );
  XOR U51675 ( .A(n42416), .B(n42423), .Z(N61634) );
  XOR U51676 ( .A(n42413), .B(n42415), .Z(n42423) );
  XNOR U51677 ( .A(n42409), .B(n42424), .Z(n42415) );
  XNOR U51678 ( .A(n42407), .B(n42410), .Z(n42424) );
  NAND U51679 ( .A(n42425), .B(n42426), .Z(n42410) );
  NAND U51680 ( .A(n42427), .B(n42428), .Z(n42426) );
  OR U51681 ( .A(n42429), .B(n42430), .Z(n42427) );
  NANDN U51682 ( .A(n42431), .B(n42429), .Z(n42425) );
  IV U51683 ( .A(n42430), .Z(n42431) );
  NAND U51684 ( .A(n42432), .B(n42433), .Z(n42407) );
  NAND U51685 ( .A(n42434), .B(n42435), .Z(n42433) );
  NANDN U51686 ( .A(n42436), .B(n42437), .Z(n42434) );
  NANDN U51687 ( .A(n42437), .B(n42436), .Z(n42432) );
  AND U51688 ( .A(n42438), .B(n42439), .Z(n42409) );
  NAND U51689 ( .A(n42440), .B(n42441), .Z(n42439) );
  OR U51690 ( .A(n42442), .B(n42443), .Z(n42440) );
  NANDN U51691 ( .A(n42444), .B(n42442), .Z(n42438) );
  NAND U51692 ( .A(n42445), .B(n42446), .Z(n42413) );
  NANDN U51693 ( .A(n42447), .B(n42448), .Z(n42446) );
  OR U51694 ( .A(n42449), .B(n42450), .Z(n42448) );
  NANDN U51695 ( .A(n42451), .B(n42449), .Z(n42445) );
  IV U51696 ( .A(n42450), .Z(n42451) );
  XNOR U51697 ( .A(n42421), .B(n42452), .Z(n42416) );
  XNOR U51698 ( .A(n42419), .B(n42422), .Z(n42452) );
  NAND U51699 ( .A(n42453), .B(n42454), .Z(n42422) );
  NAND U51700 ( .A(n42455), .B(n42456), .Z(n42454) );
  OR U51701 ( .A(n42457), .B(n42458), .Z(n42455) );
  NANDN U51702 ( .A(n42459), .B(n42457), .Z(n42453) );
  IV U51703 ( .A(n42458), .Z(n42459) );
  NAND U51704 ( .A(n42460), .B(n42461), .Z(n42419) );
  NAND U51705 ( .A(n42462), .B(n42463), .Z(n42461) );
  NANDN U51706 ( .A(n42464), .B(n42465), .Z(n42462) );
  NANDN U51707 ( .A(n42465), .B(n42464), .Z(n42460) );
  AND U51708 ( .A(n42466), .B(n42467), .Z(n42421) );
  NAND U51709 ( .A(n42468), .B(n42469), .Z(n42467) );
  OR U51710 ( .A(n42470), .B(n42471), .Z(n42468) );
  NANDN U51711 ( .A(n42472), .B(n42470), .Z(n42466) );
  XNOR U51712 ( .A(n42447), .B(n42473), .Z(N61633) );
  XOR U51713 ( .A(n42449), .B(n42450), .Z(n42473) );
  XNOR U51714 ( .A(n42463), .B(n42474), .Z(n42450) );
  XOR U51715 ( .A(n42464), .B(n42465), .Z(n42474) );
  XOR U51716 ( .A(n42470), .B(n42475), .Z(n42465) );
  XOR U51717 ( .A(n42469), .B(n42472), .Z(n42475) );
  IV U51718 ( .A(n42471), .Z(n42472) );
  NAND U51719 ( .A(n42476), .B(n42477), .Z(n42471) );
  OR U51720 ( .A(n42478), .B(n42479), .Z(n42477) );
  OR U51721 ( .A(n42480), .B(n42481), .Z(n42476) );
  NAND U51722 ( .A(n42482), .B(n42483), .Z(n42469) );
  OR U51723 ( .A(n42484), .B(n42485), .Z(n42483) );
  OR U51724 ( .A(n42486), .B(n42487), .Z(n42482) );
  NOR U51725 ( .A(n42488), .B(n42489), .Z(n42470) );
  ANDN U51726 ( .B(n42490), .A(n42491), .Z(n42464) );
  XNOR U51727 ( .A(n42457), .B(n42492), .Z(n42463) );
  XNOR U51728 ( .A(n42456), .B(n42458), .Z(n42492) );
  NAND U51729 ( .A(n42493), .B(n42494), .Z(n42458) );
  OR U51730 ( .A(n42495), .B(n42496), .Z(n42494) );
  OR U51731 ( .A(n42497), .B(n42498), .Z(n42493) );
  NAND U51732 ( .A(n42499), .B(n42500), .Z(n42456) );
  OR U51733 ( .A(n42501), .B(n42502), .Z(n42500) );
  OR U51734 ( .A(n42503), .B(n42504), .Z(n42499) );
  ANDN U51735 ( .B(n42505), .A(n42506), .Z(n42457) );
  IV U51736 ( .A(n42507), .Z(n42505) );
  ANDN U51737 ( .B(n42508), .A(n42509), .Z(n42449) );
  XOR U51738 ( .A(n42435), .B(n42510), .Z(n42447) );
  XOR U51739 ( .A(n42436), .B(n42437), .Z(n42510) );
  XOR U51740 ( .A(n42442), .B(n42511), .Z(n42437) );
  XOR U51741 ( .A(n42441), .B(n42444), .Z(n42511) );
  IV U51742 ( .A(n42443), .Z(n42444) );
  NAND U51743 ( .A(n42512), .B(n42513), .Z(n42443) );
  OR U51744 ( .A(n42514), .B(n42515), .Z(n42513) );
  OR U51745 ( .A(n42516), .B(n42517), .Z(n42512) );
  NAND U51746 ( .A(n42518), .B(n42519), .Z(n42441) );
  OR U51747 ( .A(n42520), .B(n42521), .Z(n42519) );
  OR U51748 ( .A(n42522), .B(n42523), .Z(n42518) );
  NOR U51749 ( .A(n42524), .B(n42525), .Z(n42442) );
  ANDN U51750 ( .B(n42526), .A(n42527), .Z(n42436) );
  IV U51751 ( .A(n42528), .Z(n42526) );
  XNOR U51752 ( .A(n42429), .B(n42529), .Z(n42435) );
  XNOR U51753 ( .A(n42428), .B(n42430), .Z(n42529) );
  NAND U51754 ( .A(n42530), .B(n42531), .Z(n42430) );
  OR U51755 ( .A(n42532), .B(n42533), .Z(n42531) );
  OR U51756 ( .A(n42534), .B(n42535), .Z(n42530) );
  NAND U51757 ( .A(n42536), .B(n42537), .Z(n42428) );
  OR U51758 ( .A(n42538), .B(n42539), .Z(n42537) );
  OR U51759 ( .A(n42540), .B(n42541), .Z(n42536) );
  ANDN U51760 ( .B(n42542), .A(n42543), .Z(n42429) );
  IV U51761 ( .A(n42544), .Z(n42542) );
  XNOR U51762 ( .A(n42509), .B(n42508), .Z(N61632) );
  XOR U51763 ( .A(n42528), .B(n42527), .Z(n42508) );
  XNOR U51764 ( .A(n42543), .B(n42544), .Z(n42527) );
  XNOR U51765 ( .A(n42538), .B(n42539), .Z(n42544) );
  XNOR U51766 ( .A(n42540), .B(n42541), .Z(n42539) );
  XNOR U51767 ( .A(y[1933]), .B(x[1933]), .Z(n42541) );
  XNOR U51768 ( .A(y[1934]), .B(x[1934]), .Z(n42540) );
  XNOR U51769 ( .A(y[1932]), .B(x[1932]), .Z(n42538) );
  XNOR U51770 ( .A(n42532), .B(n42533), .Z(n42543) );
  XNOR U51771 ( .A(y[1929]), .B(x[1929]), .Z(n42533) );
  XNOR U51772 ( .A(n42534), .B(n42535), .Z(n42532) );
  XNOR U51773 ( .A(y[1930]), .B(x[1930]), .Z(n42535) );
  XNOR U51774 ( .A(y[1931]), .B(x[1931]), .Z(n42534) );
  XNOR U51775 ( .A(n42525), .B(n42524), .Z(n42528) );
  XNOR U51776 ( .A(n42520), .B(n42521), .Z(n42524) );
  XNOR U51777 ( .A(y[1926]), .B(x[1926]), .Z(n42521) );
  XNOR U51778 ( .A(n42522), .B(n42523), .Z(n42520) );
  XNOR U51779 ( .A(y[1927]), .B(x[1927]), .Z(n42523) );
  XNOR U51780 ( .A(y[1928]), .B(x[1928]), .Z(n42522) );
  XNOR U51781 ( .A(n42514), .B(n42515), .Z(n42525) );
  XNOR U51782 ( .A(y[1923]), .B(x[1923]), .Z(n42515) );
  XNOR U51783 ( .A(n42516), .B(n42517), .Z(n42514) );
  XNOR U51784 ( .A(y[1924]), .B(x[1924]), .Z(n42517) );
  XNOR U51785 ( .A(y[1925]), .B(x[1925]), .Z(n42516) );
  XOR U51786 ( .A(n42490), .B(n42491), .Z(n42509) );
  XNOR U51787 ( .A(n42506), .B(n42507), .Z(n42491) );
  XNOR U51788 ( .A(n42501), .B(n42502), .Z(n42507) );
  XNOR U51789 ( .A(n42503), .B(n42504), .Z(n42502) );
  XNOR U51790 ( .A(y[1921]), .B(x[1921]), .Z(n42504) );
  XNOR U51791 ( .A(y[1922]), .B(x[1922]), .Z(n42503) );
  XNOR U51792 ( .A(y[1920]), .B(x[1920]), .Z(n42501) );
  XNOR U51793 ( .A(n42495), .B(n42496), .Z(n42506) );
  XNOR U51794 ( .A(y[1917]), .B(x[1917]), .Z(n42496) );
  XNOR U51795 ( .A(n42497), .B(n42498), .Z(n42495) );
  XNOR U51796 ( .A(y[1918]), .B(x[1918]), .Z(n42498) );
  XNOR U51797 ( .A(y[1919]), .B(x[1919]), .Z(n42497) );
  XOR U51798 ( .A(n42489), .B(n42488), .Z(n42490) );
  XNOR U51799 ( .A(n42484), .B(n42485), .Z(n42488) );
  XNOR U51800 ( .A(y[1914]), .B(x[1914]), .Z(n42485) );
  XNOR U51801 ( .A(n42486), .B(n42487), .Z(n42484) );
  XNOR U51802 ( .A(y[1915]), .B(x[1915]), .Z(n42487) );
  XNOR U51803 ( .A(y[1916]), .B(x[1916]), .Z(n42486) );
  XNOR U51804 ( .A(n42478), .B(n42479), .Z(n42489) );
  XNOR U51805 ( .A(y[1911]), .B(x[1911]), .Z(n42479) );
  XNOR U51806 ( .A(n42480), .B(n42481), .Z(n42478) );
  XNOR U51807 ( .A(y[1912]), .B(x[1912]), .Z(n42481) );
  XNOR U51808 ( .A(y[1913]), .B(x[1913]), .Z(n42480) );
  NAND U51809 ( .A(n42545), .B(n42546), .Z(N61623) );
  NANDN U51810 ( .A(n42547), .B(n42548), .Z(n42546) );
  OR U51811 ( .A(n42549), .B(n42550), .Z(n42548) );
  NAND U51812 ( .A(n42549), .B(n42550), .Z(n42545) );
  XOR U51813 ( .A(n42549), .B(n42551), .Z(N61622) );
  XNOR U51814 ( .A(n42547), .B(n42550), .Z(n42551) );
  AND U51815 ( .A(n42552), .B(n42553), .Z(n42550) );
  NANDN U51816 ( .A(n42554), .B(n42555), .Z(n42553) );
  NANDN U51817 ( .A(n42556), .B(n42557), .Z(n42555) );
  NANDN U51818 ( .A(n42557), .B(n42556), .Z(n42552) );
  NAND U51819 ( .A(n42558), .B(n42559), .Z(n42547) );
  NANDN U51820 ( .A(n42560), .B(n42561), .Z(n42559) );
  OR U51821 ( .A(n42562), .B(n42563), .Z(n42561) );
  NAND U51822 ( .A(n42563), .B(n42562), .Z(n42558) );
  AND U51823 ( .A(n42564), .B(n42565), .Z(n42549) );
  NANDN U51824 ( .A(n42566), .B(n42567), .Z(n42565) );
  NANDN U51825 ( .A(n42568), .B(n42569), .Z(n42567) );
  NANDN U51826 ( .A(n42569), .B(n42568), .Z(n42564) );
  XOR U51827 ( .A(n42563), .B(n42570), .Z(N61621) );
  XOR U51828 ( .A(n42560), .B(n42562), .Z(n42570) );
  XNOR U51829 ( .A(n42556), .B(n42571), .Z(n42562) );
  XNOR U51830 ( .A(n42554), .B(n42557), .Z(n42571) );
  NAND U51831 ( .A(n42572), .B(n42573), .Z(n42557) );
  NAND U51832 ( .A(n42574), .B(n42575), .Z(n42573) );
  OR U51833 ( .A(n42576), .B(n42577), .Z(n42574) );
  NANDN U51834 ( .A(n42578), .B(n42576), .Z(n42572) );
  IV U51835 ( .A(n42577), .Z(n42578) );
  NAND U51836 ( .A(n42579), .B(n42580), .Z(n42554) );
  NAND U51837 ( .A(n42581), .B(n42582), .Z(n42580) );
  NANDN U51838 ( .A(n42583), .B(n42584), .Z(n42581) );
  NANDN U51839 ( .A(n42584), .B(n42583), .Z(n42579) );
  AND U51840 ( .A(n42585), .B(n42586), .Z(n42556) );
  NAND U51841 ( .A(n42587), .B(n42588), .Z(n42586) );
  OR U51842 ( .A(n42589), .B(n42590), .Z(n42587) );
  NANDN U51843 ( .A(n42591), .B(n42589), .Z(n42585) );
  NAND U51844 ( .A(n42592), .B(n42593), .Z(n42560) );
  NANDN U51845 ( .A(n42594), .B(n42595), .Z(n42593) );
  OR U51846 ( .A(n42596), .B(n42597), .Z(n42595) );
  NANDN U51847 ( .A(n42598), .B(n42596), .Z(n42592) );
  IV U51848 ( .A(n42597), .Z(n42598) );
  XNOR U51849 ( .A(n42568), .B(n42599), .Z(n42563) );
  XNOR U51850 ( .A(n42566), .B(n42569), .Z(n42599) );
  NAND U51851 ( .A(n42600), .B(n42601), .Z(n42569) );
  NAND U51852 ( .A(n42602), .B(n42603), .Z(n42601) );
  OR U51853 ( .A(n42604), .B(n42605), .Z(n42602) );
  NANDN U51854 ( .A(n42606), .B(n42604), .Z(n42600) );
  IV U51855 ( .A(n42605), .Z(n42606) );
  NAND U51856 ( .A(n42607), .B(n42608), .Z(n42566) );
  NAND U51857 ( .A(n42609), .B(n42610), .Z(n42608) );
  NANDN U51858 ( .A(n42611), .B(n42612), .Z(n42609) );
  NANDN U51859 ( .A(n42612), .B(n42611), .Z(n42607) );
  AND U51860 ( .A(n42613), .B(n42614), .Z(n42568) );
  NAND U51861 ( .A(n42615), .B(n42616), .Z(n42614) );
  OR U51862 ( .A(n42617), .B(n42618), .Z(n42615) );
  NANDN U51863 ( .A(n42619), .B(n42617), .Z(n42613) );
  XNOR U51864 ( .A(n42594), .B(n42620), .Z(N61620) );
  XOR U51865 ( .A(n42596), .B(n42597), .Z(n42620) );
  XNOR U51866 ( .A(n42610), .B(n42621), .Z(n42597) );
  XOR U51867 ( .A(n42611), .B(n42612), .Z(n42621) );
  XOR U51868 ( .A(n42617), .B(n42622), .Z(n42612) );
  XOR U51869 ( .A(n42616), .B(n42619), .Z(n42622) );
  IV U51870 ( .A(n42618), .Z(n42619) );
  NAND U51871 ( .A(n42623), .B(n42624), .Z(n42618) );
  OR U51872 ( .A(n42625), .B(n42626), .Z(n42624) );
  OR U51873 ( .A(n42627), .B(n42628), .Z(n42623) );
  NAND U51874 ( .A(n42629), .B(n42630), .Z(n42616) );
  OR U51875 ( .A(n42631), .B(n42632), .Z(n42630) );
  OR U51876 ( .A(n42633), .B(n42634), .Z(n42629) );
  NOR U51877 ( .A(n42635), .B(n42636), .Z(n42617) );
  ANDN U51878 ( .B(n42637), .A(n42638), .Z(n42611) );
  XNOR U51879 ( .A(n42604), .B(n42639), .Z(n42610) );
  XNOR U51880 ( .A(n42603), .B(n42605), .Z(n42639) );
  NAND U51881 ( .A(n42640), .B(n42641), .Z(n42605) );
  OR U51882 ( .A(n42642), .B(n42643), .Z(n42641) );
  OR U51883 ( .A(n42644), .B(n42645), .Z(n42640) );
  NAND U51884 ( .A(n42646), .B(n42647), .Z(n42603) );
  OR U51885 ( .A(n42648), .B(n42649), .Z(n42647) );
  OR U51886 ( .A(n42650), .B(n42651), .Z(n42646) );
  ANDN U51887 ( .B(n42652), .A(n42653), .Z(n42604) );
  IV U51888 ( .A(n42654), .Z(n42652) );
  ANDN U51889 ( .B(n42655), .A(n42656), .Z(n42596) );
  XOR U51890 ( .A(n42582), .B(n42657), .Z(n42594) );
  XOR U51891 ( .A(n42583), .B(n42584), .Z(n42657) );
  XOR U51892 ( .A(n42589), .B(n42658), .Z(n42584) );
  XOR U51893 ( .A(n42588), .B(n42591), .Z(n42658) );
  IV U51894 ( .A(n42590), .Z(n42591) );
  NAND U51895 ( .A(n42659), .B(n42660), .Z(n42590) );
  OR U51896 ( .A(n42661), .B(n42662), .Z(n42660) );
  OR U51897 ( .A(n42663), .B(n42664), .Z(n42659) );
  NAND U51898 ( .A(n42665), .B(n42666), .Z(n42588) );
  OR U51899 ( .A(n42667), .B(n42668), .Z(n42666) );
  OR U51900 ( .A(n42669), .B(n42670), .Z(n42665) );
  NOR U51901 ( .A(n42671), .B(n42672), .Z(n42589) );
  ANDN U51902 ( .B(n42673), .A(n42674), .Z(n42583) );
  IV U51903 ( .A(n42675), .Z(n42673) );
  XNOR U51904 ( .A(n42576), .B(n42676), .Z(n42582) );
  XNOR U51905 ( .A(n42575), .B(n42577), .Z(n42676) );
  NAND U51906 ( .A(n42677), .B(n42678), .Z(n42577) );
  OR U51907 ( .A(n42679), .B(n42680), .Z(n42678) );
  OR U51908 ( .A(n42681), .B(n42682), .Z(n42677) );
  NAND U51909 ( .A(n42683), .B(n42684), .Z(n42575) );
  OR U51910 ( .A(n42685), .B(n42686), .Z(n42684) );
  OR U51911 ( .A(n42687), .B(n42688), .Z(n42683) );
  ANDN U51912 ( .B(n42689), .A(n42690), .Z(n42576) );
  IV U51913 ( .A(n42691), .Z(n42689) );
  XNOR U51914 ( .A(n42656), .B(n42655), .Z(N61619) );
  XOR U51915 ( .A(n42675), .B(n42674), .Z(n42655) );
  XNOR U51916 ( .A(n42690), .B(n42691), .Z(n42674) );
  XNOR U51917 ( .A(n42685), .B(n42686), .Z(n42691) );
  XNOR U51918 ( .A(n42687), .B(n42688), .Z(n42686) );
  XNOR U51919 ( .A(y[1909]), .B(x[1909]), .Z(n42688) );
  XNOR U51920 ( .A(y[1910]), .B(x[1910]), .Z(n42687) );
  XNOR U51921 ( .A(y[1908]), .B(x[1908]), .Z(n42685) );
  XNOR U51922 ( .A(n42679), .B(n42680), .Z(n42690) );
  XNOR U51923 ( .A(y[1905]), .B(x[1905]), .Z(n42680) );
  XNOR U51924 ( .A(n42681), .B(n42682), .Z(n42679) );
  XNOR U51925 ( .A(y[1906]), .B(x[1906]), .Z(n42682) );
  XNOR U51926 ( .A(y[1907]), .B(x[1907]), .Z(n42681) );
  XNOR U51927 ( .A(n42672), .B(n42671), .Z(n42675) );
  XNOR U51928 ( .A(n42667), .B(n42668), .Z(n42671) );
  XNOR U51929 ( .A(y[1902]), .B(x[1902]), .Z(n42668) );
  XNOR U51930 ( .A(n42669), .B(n42670), .Z(n42667) );
  XNOR U51931 ( .A(y[1903]), .B(x[1903]), .Z(n42670) );
  XNOR U51932 ( .A(y[1904]), .B(x[1904]), .Z(n42669) );
  XNOR U51933 ( .A(n42661), .B(n42662), .Z(n42672) );
  XNOR U51934 ( .A(y[1899]), .B(x[1899]), .Z(n42662) );
  XNOR U51935 ( .A(n42663), .B(n42664), .Z(n42661) );
  XNOR U51936 ( .A(y[1900]), .B(x[1900]), .Z(n42664) );
  XNOR U51937 ( .A(y[1901]), .B(x[1901]), .Z(n42663) );
  XOR U51938 ( .A(n42637), .B(n42638), .Z(n42656) );
  XNOR U51939 ( .A(n42653), .B(n42654), .Z(n42638) );
  XNOR U51940 ( .A(n42648), .B(n42649), .Z(n42654) );
  XNOR U51941 ( .A(n42650), .B(n42651), .Z(n42649) );
  XNOR U51942 ( .A(y[1897]), .B(x[1897]), .Z(n42651) );
  XNOR U51943 ( .A(y[1898]), .B(x[1898]), .Z(n42650) );
  XNOR U51944 ( .A(y[1896]), .B(x[1896]), .Z(n42648) );
  XNOR U51945 ( .A(n42642), .B(n42643), .Z(n42653) );
  XNOR U51946 ( .A(y[1893]), .B(x[1893]), .Z(n42643) );
  XNOR U51947 ( .A(n42644), .B(n42645), .Z(n42642) );
  XNOR U51948 ( .A(y[1894]), .B(x[1894]), .Z(n42645) );
  XNOR U51949 ( .A(y[1895]), .B(x[1895]), .Z(n42644) );
  XOR U51950 ( .A(n42636), .B(n42635), .Z(n42637) );
  XNOR U51951 ( .A(n42631), .B(n42632), .Z(n42635) );
  XNOR U51952 ( .A(y[1890]), .B(x[1890]), .Z(n42632) );
  XNOR U51953 ( .A(n42633), .B(n42634), .Z(n42631) );
  XNOR U51954 ( .A(y[1891]), .B(x[1891]), .Z(n42634) );
  XNOR U51955 ( .A(y[1892]), .B(x[1892]), .Z(n42633) );
  XNOR U51956 ( .A(n42625), .B(n42626), .Z(n42636) );
  XNOR U51957 ( .A(y[1887]), .B(x[1887]), .Z(n42626) );
  XNOR U51958 ( .A(n42627), .B(n42628), .Z(n42625) );
  XNOR U51959 ( .A(y[1888]), .B(x[1888]), .Z(n42628) );
  XNOR U51960 ( .A(y[1889]), .B(x[1889]), .Z(n42627) );
  NAND U51961 ( .A(n42692), .B(n42693), .Z(N61610) );
  NANDN U51962 ( .A(n42694), .B(n42695), .Z(n42693) );
  OR U51963 ( .A(n42696), .B(n42697), .Z(n42695) );
  NAND U51964 ( .A(n42696), .B(n42697), .Z(n42692) );
  XOR U51965 ( .A(n42696), .B(n42698), .Z(N61609) );
  XNOR U51966 ( .A(n42694), .B(n42697), .Z(n42698) );
  AND U51967 ( .A(n42699), .B(n42700), .Z(n42697) );
  NANDN U51968 ( .A(n42701), .B(n42702), .Z(n42700) );
  NANDN U51969 ( .A(n42703), .B(n42704), .Z(n42702) );
  NANDN U51970 ( .A(n42704), .B(n42703), .Z(n42699) );
  NAND U51971 ( .A(n42705), .B(n42706), .Z(n42694) );
  NANDN U51972 ( .A(n42707), .B(n42708), .Z(n42706) );
  OR U51973 ( .A(n42709), .B(n42710), .Z(n42708) );
  NAND U51974 ( .A(n42710), .B(n42709), .Z(n42705) );
  AND U51975 ( .A(n42711), .B(n42712), .Z(n42696) );
  NANDN U51976 ( .A(n42713), .B(n42714), .Z(n42712) );
  NANDN U51977 ( .A(n42715), .B(n42716), .Z(n42714) );
  NANDN U51978 ( .A(n42716), .B(n42715), .Z(n42711) );
  XOR U51979 ( .A(n42710), .B(n42717), .Z(N61608) );
  XOR U51980 ( .A(n42707), .B(n42709), .Z(n42717) );
  XNOR U51981 ( .A(n42703), .B(n42718), .Z(n42709) );
  XNOR U51982 ( .A(n42701), .B(n42704), .Z(n42718) );
  NAND U51983 ( .A(n42719), .B(n42720), .Z(n42704) );
  NAND U51984 ( .A(n42721), .B(n42722), .Z(n42720) );
  OR U51985 ( .A(n42723), .B(n42724), .Z(n42721) );
  NANDN U51986 ( .A(n42725), .B(n42723), .Z(n42719) );
  IV U51987 ( .A(n42724), .Z(n42725) );
  NAND U51988 ( .A(n42726), .B(n42727), .Z(n42701) );
  NAND U51989 ( .A(n42728), .B(n42729), .Z(n42727) );
  NANDN U51990 ( .A(n42730), .B(n42731), .Z(n42728) );
  NANDN U51991 ( .A(n42731), .B(n42730), .Z(n42726) );
  AND U51992 ( .A(n42732), .B(n42733), .Z(n42703) );
  NAND U51993 ( .A(n42734), .B(n42735), .Z(n42733) );
  OR U51994 ( .A(n42736), .B(n42737), .Z(n42734) );
  NANDN U51995 ( .A(n42738), .B(n42736), .Z(n42732) );
  NAND U51996 ( .A(n42739), .B(n42740), .Z(n42707) );
  NANDN U51997 ( .A(n42741), .B(n42742), .Z(n42740) );
  OR U51998 ( .A(n42743), .B(n42744), .Z(n42742) );
  NANDN U51999 ( .A(n42745), .B(n42743), .Z(n42739) );
  IV U52000 ( .A(n42744), .Z(n42745) );
  XNOR U52001 ( .A(n42715), .B(n42746), .Z(n42710) );
  XNOR U52002 ( .A(n42713), .B(n42716), .Z(n42746) );
  NAND U52003 ( .A(n42747), .B(n42748), .Z(n42716) );
  NAND U52004 ( .A(n42749), .B(n42750), .Z(n42748) );
  OR U52005 ( .A(n42751), .B(n42752), .Z(n42749) );
  NANDN U52006 ( .A(n42753), .B(n42751), .Z(n42747) );
  IV U52007 ( .A(n42752), .Z(n42753) );
  NAND U52008 ( .A(n42754), .B(n42755), .Z(n42713) );
  NAND U52009 ( .A(n42756), .B(n42757), .Z(n42755) );
  NANDN U52010 ( .A(n42758), .B(n42759), .Z(n42756) );
  NANDN U52011 ( .A(n42759), .B(n42758), .Z(n42754) );
  AND U52012 ( .A(n42760), .B(n42761), .Z(n42715) );
  NAND U52013 ( .A(n42762), .B(n42763), .Z(n42761) );
  OR U52014 ( .A(n42764), .B(n42765), .Z(n42762) );
  NANDN U52015 ( .A(n42766), .B(n42764), .Z(n42760) );
  XNOR U52016 ( .A(n42741), .B(n42767), .Z(N61607) );
  XOR U52017 ( .A(n42743), .B(n42744), .Z(n42767) );
  XNOR U52018 ( .A(n42757), .B(n42768), .Z(n42744) );
  XOR U52019 ( .A(n42758), .B(n42759), .Z(n42768) );
  XOR U52020 ( .A(n42764), .B(n42769), .Z(n42759) );
  XOR U52021 ( .A(n42763), .B(n42766), .Z(n42769) );
  IV U52022 ( .A(n42765), .Z(n42766) );
  NAND U52023 ( .A(n42770), .B(n42771), .Z(n42765) );
  OR U52024 ( .A(n42772), .B(n42773), .Z(n42771) );
  OR U52025 ( .A(n42774), .B(n42775), .Z(n42770) );
  NAND U52026 ( .A(n42776), .B(n42777), .Z(n42763) );
  OR U52027 ( .A(n42778), .B(n42779), .Z(n42777) );
  OR U52028 ( .A(n42780), .B(n42781), .Z(n42776) );
  NOR U52029 ( .A(n42782), .B(n42783), .Z(n42764) );
  ANDN U52030 ( .B(n42784), .A(n42785), .Z(n42758) );
  XNOR U52031 ( .A(n42751), .B(n42786), .Z(n42757) );
  XNOR U52032 ( .A(n42750), .B(n42752), .Z(n42786) );
  NAND U52033 ( .A(n42787), .B(n42788), .Z(n42752) );
  OR U52034 ( .A(n42789), .B(n42790), .Z(n42788) );
  OR U52035 ( .A(n42791), .B(n42792), .Z(n42787) );
  NAND U52036 ( .A(n42793), .B(n42794), .Z(n42750) );
  OR U52037 ( .A(n42795), .B(n42796), .Z(n42794) );
  OR U52038 ( .A(n42797), .B(n42798), .Z(n42793) );
  ANDN U52039 ( .B(n42799), .A(n42800), .Z(n42751) );
  IV U52040 ( .A(n42801), .Z(n42799) );
  ANDN U52041 ( .B(n42802), .A(n42803), .Z(n42743) );
  XOR U52042 ( .A(n42729), .B(n42804), .Z(n42741) );
  XOR U52043 ( .A(n42730), .B(n42731), .Z(n42804) );
  XOR U52044 ( .A(n42736), .B(n42805), .Z(n42731) );
  XOR U52045 ( .A(n42735), .B(n42738), .Z(n42805) );
  IV U52046 ( .A(n42737), .Z(n42738) );
  NAND U52047 ( .A(n42806), .B(n42807), .Z(n42737) );
  OR U52048 ( .A(n42808), .B(n42809), .Z(n42807) );
  OR U52049 ( .A(n42810), .B(n42811), .Z(n42806) );
  NAND U52050 ( .A(n42812), .B(n42813), .Z(n42735) );
  OR U52051 ( .A(n42814), .B(n42815), .Z(n42813) );
  OR U52052 ( .A(n42816), .B(n42817), .Z(n42812) );
  NOR U52053 ( .A(n42818), .B(n42819), .Z(n42736) );
  ANDN U52054 ( .B(n42820), .A(n42821), .Z(n42730) );
  IV U52055 ( .A(n42822), .Z(n42820) );
  XNOR U52056 ( .A(n42723), .B(n42823), .Z(n42729) );
  XNOR U52057 ( .A(n42722), .B(n42724), .Z(n42823) );
  NAND U52058 ( .A(n42824), .B(n42825), .Z(n42724) );
  OR U52059 ( .A(n42826), .B(n42827), .Z(n42825) );
  OR U52060 ( .A(n42828), .B(n42829), .Z(n42824) );
  NAND U52061 ( .A(n42830), .B(n42831), .Z(n42722) );
  OR U52062 ( .A(n42832), .B(n42833), .Z(n42831) );
  OR U52063 ( .A(n42834), .B(n42835), .Z(n42830) );
  ANDN U52064 ( .B(n42836), .A(n42837), .Z(n42723) );
  IV U52065 ( .A(n42838), .Z(n42836) );
  XNOR U52066 ( .A(n42803), .B(n42802), .Z(N61606) );
  XOR U52067 ( .A(n42822), .B(n42821), .Z(n42802) );
  XNOR U52068 ( .A(n42837), .B(n42838), .Z(n42821) );
  XNOR U52069 ( .A(n42832), .B(n42833), .Z(n42838) );
  XNOR U52070 ( .A(n42834), .B(n42835), .Z(n42833) );
  XNOR U52071 ( .A(y[1885]), .B(x[1885]), .Z(n42835) );
  XNOR U52072 ( .A(y[1886]), .B(x[1886]), .Z(n42834) );
  XNOR U52073 ( .A(y[1884]), .B(x[1884]), .Z(n42832) );
  XNOR U52074 ( .A(n42826), .B(n42827), .Z(n42837) );
  XNOR U52075 ( .A(y[1881]), .B(x[1881]), .Z(n42827) );
  XNOR U52076 ( .A(n42828), .B(n42829), .Z(n42826) );
  XNOR U52077 ( .A(y[1882]), .B(x[1882]), .Z(n42829) );
  XNOR U52078 ( .A(y[1883]), .B(x[1883]), .Z(n42828) );
  XNOR U52079 ( .A(n42819), .B(n42818), .Z(n42822) );
  XNOR U52080 ( .A(n42814), .B(n42815), .Z(n42818) );
  XNOR U52081 ( .A(y[1878]), .B(x[1878]), .Z(n42815) );
  XNOR U52082 ( .A(n42816), .B(n42817), .Z(n42814) );
  XNOR U52083 ( .A(y[1879]), .B(x[1879]), .Z(n42817) );
  XNOR U52084 ( .A(y[1880]), .B(x[1880]), .Z(n42816) );
  XNOR U52085 ( .A(n42808), .B(n42809), .Z(n42819) );
  XNOR U52086 ( .A(y[1875]), .B(x[1875]), .Z(n42809) );
  XNOR U52087 ( .A(n42810), .B(n42811), .Z(n42808) );
  XNOR U52088 ( .A(y[1876]), .B(x[1876]), .Z(n42811) );
  XNOR U52089 ( .A(y[1877]), .B(x[1877]), .Z(n42810) );
  XOR U52090 ( .A(n42784), .B(n42785), .Z(n42803) );
  XNOR U52091 ( .A(n42800), .B(n42801), .Z(n42785) );
  XNOR U52092 ( .A(n42795), .B(n42796), .Z(n42801) );
  XNOR U52093 ( .A(n42797), .B(n42798), .Z(n42796) );
  XNOR U52094 ( .A(y[1873]), .B(x[1873]), .Z(n42798) );
  XNOR U52095 ( .A(y[1874]), .B(x[1874]), .Z(n42797) );
  XNOR U52096 ( .A(y[1872]), .B(x[1872]), .Z(n42795) );
  XNOR U52097 ( .A(n42789), .B(n42790), .Z(n42800) );
  XNOR U52098 ( .A(y[1869]), .B(x[1869]), .Z(n42790) );
  XNOR U52099 ( .A(n42791), .B(n42792), .Z(n42789) );
  XNOR U52100 ( .A(y[1870]), .B(x[1870]), .Z(n42792) );
  XNOR U52101 ( .A(y[1871]), .B(x[1871]), .Z(n42791) );
  XOR U52102 ( .A(n42783), .B(n42782), .Z(n42784) );
  XNOR U52103 ( .A(n42778), .B(n42779), .Z(n42782) );
  XNOR U52104 ( .A(y[1866]), .B(x[1866]), .Z(n42779) );
  XNOR U52105 ( .A(n42780), .B(n42781), .Z(n42778) );
  XNOR U52106 ( .A(y[1867]), .B(x[1867]), .Z(n42781) );
  XNOR U52107 ( .A(y[1868]), .B(x[1868]), .Z(n42780) );
  XNOR U52108 ( .A(n42772), .B(n42773), .Z(n42783) );
  XNOR U52109 ( .A(y[1863]), .B(x[1863]), .Z(n42773) );
  XNOR U52110 ( .A(n42774), .B(n42775), .Z(n42772) );
  XNOR U52111 ( .A(y[1864]), .B(x[1864]), .Z(n42775) );
  XNOR U52112 ( .A(y[1865]), .B(x[1865]), .Z(n42774) );
  NAND U52113 ( .A(n42839), .B(n42840), .Z(N61597) );
  NANDN U52114 ( .A(n42841), .B(n42842), .Z(n42840) );
  OR U52115 ( .A(n42843), .B(n42844), .Z(n42842) );
  NAND U52116 ( .A(n42843), .B(n42844), .Z(n42839) );
  XOR U52117 ( .A(n42843), .B(n42845), .Z(N61596) );
  XNOR U52118 ( .A(n42841), .B(n42844), .Z(n42845) );
  AND U52119 ( .A(n42846), .B(n42847), .Z(n42844) );
  NANDN U52120 ( .A(n42848), .B(n42849), .Z(n42847) );
  NANDN U52121 ( .A(n42850), .B(n42851), .Z(n42849) );
  NANDN U52122 ( .A(n42851), .B(n42850), .Z(n42846) );
  NAND U52123 ( .A(n42852), .B(n42853), .Z(n42841) );
  NANDN U52124 ( .A(n42854), .B(n42855), .Z(n42853) );
  OR U52125 ( .A(n42856), .B(n42857), .Z(n42855) );
  NAND U52126 ( .A(n42857), .B(n42856), .Z(n42852) );
  AND U52127 ( .A(n42858), .B(n42859), .Z(n42843) );
  NANDN U52128 ( .A(n42860), .B(n42861), .Z(n42859) );
  NANDN U52129 ( .A(n42862), .B(n42863), .Z(n42861) );
  NANDN U52130 ( .A(n42863), .B(n42862), .Z(n42858) );
  XOR U52131 ( .A(n42857), .B(n42864), .Z(N61595) );
  XOR U52132 ( .A(n42854), .B(n42856), .Z(n42864) );
  XNOR U52133 ( .A(n42850), .B(n42865), .Z(n42856) );
  XNOR U52134 ( .A(n42848), .B(n42851), .Z(n42865) );
  NAND U52135 ( .A(n42866), .B(n42867), .Z(n42851) );
  NAND U52136 ( .A(n42868), .B(n42869), .Z(n42867) );
  OR U52137 ( .A(n42870), .B(n42871), .Z(n42868) );
  NANDN U52138 ( .A(n42872), .B(n42870), .Z(n42866) );
  IV U52139 ( .A(n42871), .Z(n42872) );
  NAND U52140 ( .A(n42873), .B(n42874), .Z(n42848) );
  NAND U52141 ( .A(n42875), .B(n42876), .Z(n42874) );
  NANDN U52142 ( .A(n42877), .B(n42878), .Z(n42875) );
  NANDN U52143 ( .A(n42878), .B(n42877), .Z(n42873) );
  AND U52144 ( .A(n42879), .B(n42880), .Z(n42850) );
  NAND U52145 ( .A(n42881), .B(n42882), .Z(n42880) );
  OR U52146 ( .A(n42883), .B(n42884), .Z(n42881) );
  NANDN U52147 ( .A(n42885), .B(n42883), .Z(n42879) );
  NAND U52148 ( .A(n42886), .B(n42887), .Z(n42854) );
  NANDN U52149 ( .A(n42888), .B(n42889), .Z(n42887) );
  OR U52150 ( .A(n42890), .B(n42891), .Z(n42889) );
  NANDN U52151 ( .A(n42892), .B(n42890), .Z(n42886) );
  IV U52152 ( .A(n42891), .Z(n42892) );
  XNOR U52153 ( .A(n42862), .B(n42893), .Z(n42857) );
  XNOR U52154 ( .A(n42860), .B(n42863), .Z(n42893) );
  NAND U52155 ( .A(n42894), .B(n42895), .Z(n42863) );
  NAND U52156 ( .A(n42896), .B(n42897), .Z(n42895) );
  OR U52157 ( .A(n42898), .B(n42899), .Z(n42896) );
  NANDN U52158 ( .A(n42900), .B(n42898), .Z(n42894) );
  IV U52159 ( .A(n42899), .Z(n42900) );
  NAND U52160 ( .A(n42901), .B(n42902), .Z(n42860) );
  NAND U52161 ( .A(n42903), .B(n42904), .Z(n42902) );
  NANDN U52162 ( .A(n42905), .B(n42906), .Z(n42903) );
  NANDN U52163 ( .A(n42906), .B(n42905), .Z(n42901) );
  AND U52164 ( .A(n42907), .B(n42908), .Z(n42862) );
  NAND U52165 ( .A(n42909), .B(n42910), .Z(n42908) );
  OR U52166 ( .A(n42911), .B(n42912), .Z(n42909) );
  NANDN U52167 ( .A(n42913), .B(n42911), .Z(n42907) );
  XNOR U52168 ( .A(n42888), .B(n42914), .Z(N61594) );
  XOR U52169 ( .A(n42890), .B(n42891), .Z(n42914) );
  XNOR U52170 ( .A(n42904), .B(n42915), .Z(n42891) );
  XOR U52171 ( .A(n42905), .B(n42906), .Z(n42915) );
  XOR U52172 ( .A(n42911), .B(n42916), .Z(n42906) );
  XOR U52173 ( .A(n42910), .B(n42913), .Z(n42916) );
  IV U52174 ( .A(n42912), .Z(n42913) );
  NAND U52175 ( .A(n42917), .B(n42918), .Z(n42912) );
  OR U52176 ( .A(n42919), .B(n42920), .Z(n42918) );
  OR U52177 ( .A(n42921), .B(n42922), .Z(n42917) );
  NAND U52178 ( .A(n42923), .B(n42924), .Z(n42910) );
  OR U52179 ( .A(n42925), .B(n42926), .Z(n42924) );
  OR U52180 ( .A(n42927), .B(n42928), .Z(n42923) );
  NOR U52181 ( .A(n42929), .B(n42930), .Z(n42911) );
  ANDN U52182 ( .B(n42931), .A(n42932), .Z(n42905) );
  XNOR U52183 ( .A(n42898), .B(n42933), .Z(n42904) );
  XNOR U52184 ( .A(n42897), .B(n42899), .Z(n42933) );
  NAND U52185 ( .A(n42934), .B(n42935), .Z(n42899) );
  OR U52186 ( .A(n42936), .B(n42937), .Z(n42935) );
  OR U52187 ( .A(n42938), .B(n42939), .Z(n42934) );
  NAND U52188 ( .A(n42940), .B(n42941), .Z(n42897) );
  OR U52189 ( .A(n42942), .B(n42943), .Z(n42941) );
  OR U52190 ( .A(n42944), .B(n42945), .Z(n42940) );
  ANDN U52191 ( .B(n42946), .A(n42947), .Z(n42898) );
  IV U52192 ( .A(n42948), .Z(n42946) );
  ANDN U52193 ( .B(n42949), .A(n42950), .Z(n42890) );
  XOR U52194 ( .A(n42876), .B(n42951), .Z(n42888) );
  XOR U52195 ( .A(n42877), .B(n42878), .Z(n42951) );
  XOR U52196 ( .A(n42883), .B(n42952), .Z(n42878) );
  XOR U52197 ( .A(n42882), .B(n42885), .Z(n42952) );
  IV U52198 ( .A(n42884), .Z(n42885) );
  NAND U52199 ( .A(n42953), .B(n42954), .Z(n42884) );
  OR U52200 ( .A(n42955), .B(n42956), .Z(n42954) );
  OR U52201 ( .A(n42957), .B(n42958), .Z(n42953) );
  NAND U52202 ( .A(n42959), .B(n42960), .Z(n42882) );
  OR U52203 ( .A(n42961), .B(n42962), .Z(n42960) );
  OR U52204 ( .A(n42963), .B(n42964), .Z(n42959) );
  NOR U52205 ( .A(n42965), .B(n42966), .Z(n42883) );
  ANDN U52206 ( .B(n42967), .A(n42968), .Z(n42877) );
  IV U52207 ( .A(n42969), .Z(n42967) );
  XNOR U52208 ( .A(n42870), .B(n42970), .Z(n42876) );
  XNOR U52209 ( .A(n42869), .B(n42871), .Z(n42970) );
  NAND U52210 ( .A(n42971), .B(n42972), .Z(n42871) );
  OR U52211 ( .A(n42973), .B(n42974), .Z(n42972) );
  OR U52212 ( .A(n42975), .B(n42976), .Z(n42971) );
  NAND U52213 ( .A(n42977), .B(n42978), .Z(n42869) );
  OR U52214 ( .A(n42979), .B(n42980), .Z(n42978) );
  OR U52215 ( .A(n42981), .B(n42982), .Z(n42977) );
  ANDN U52216 ( .B(n42983), .A(n42984), .Z(n42870) );
  IV U52217 ( .A(n42985), .Z(n42983) );
  XNOR U52218 ( .A(n42950), .B(n42949), .Z(N61593) );
  XOR U52219 ( .A(n42969), .B(n42968), .Z(n42949) );
  XNOR U52220 ( .A(n42984), .B(n42985), .Z(n42968) );
  XNOR U52221 ( .A(n42979), .B(n42980), .Z(n42985) );
  XNOR U52222 ( .A(n42981), .B(n42982), .Z(n42980) );
  XNOR U52223 ( .A(y[1861]), .B(x[1861]), .Z(n42982) );
  XNOR U52224 ( .A(y[1862]), .B(x[1862]), .Z(n42981) );
  XNOR U52225 ( .A(y[1860]), .B(x[1860]), .Z(n42979) );
  XNOR U52226 ( .A(n42973), .B(n42974), .Z(n42984) );
  XNOR U52227 ( .A(y[1857]), .B(x[1857]), .Z(n42974) );
  XNOR U52228 ( .A(n42975), .B(n42976), .Z(n42973) );
  XNOR U52229 ( .A(y[1858]), .B(x[1858]), .Z(n42976) );
  XNOR U52230 ( .A(y[1859]), .B(x[1859]), .Z(n42975) );
  XNOR U52231 ( .A(n42966), .B(n42965), .Z(n42969) );
  XNOR U52232 ( .A(n42961), .B(n42962), .Z(n42965) );
  XNOR U52233 ( .A(y[1854]), .B(x[1854]), .Z(n42962) );
  XNOR U52234 ( .A(n42963), .B(n42964), .Z(n42961) );
  XNOR U52235 ( .A(y[1855]), .B(x[1855]), .Z(n42964) );
  XNOR U52236 ( .A(y[1856]), .B(x[1856]), .Z(n42963) );
  XNOR U52237 ( .A(n42955), .B(n42956), .Z(n42966) );
  XNOR U52238 ( .A(y[1851]), .B(x[1851]), .Z(n42956) );
  XNOR U52239 ( .A(n42957), .B(n42958), .Z(n42955) );
  XNOR U52240 ( .A(y[1852]), .B(x[1852]), .Z(n42958) );
  XNOR U52241 ( .A(y[1853]), .B(x[1853]), .Z(n42957) );
  XOR U52242 ( .A(n42931), .B(n42932), .Z(n42950) );
  XNOR U52243 ( .A(n42947), .B(n42948), .Z(n42932) );
  XNOR U52244 ( .A(n42942), .B(n42943), .Z(n42948) );
  XNOR U52245 ( .A(n42944), .B(n42945), .Z(n42943) );
  XNOR U52246 ( .A(y[1849]), .B(x[1849]), .Z(n42945) );
  XNOR U52247 ( .A(y[1850]), .B(x[1850]), .Z(n42944) );
  XNOR U52248 ( .A(y[1848]), .B(x[1848]), .Z(n42942) );
  XNOR U52249 ( .A(n42936), .B(n42937), .Z(n42947) );
  XNOR U52250 ( .A(y[1845]), .B(x[1845]), .Z(n42937) );
  XNOR U52251 ( .A(n42938), .B(n42939), .Z(n42936) );
  XNOR U52252 ( .A(y[1846]), .B(x[1846]), .Z(n42939) );
  XNOR U52253 ( .A(y[1847]), .B(x[1847]), .Z(n42938) );
  XOR U52254 ( .A(n42930), .B(n42929), .Z(n42931) );
  XNOR U52255 ( .A(n42925), .B(n42926), .Z(n42929) );
  XNOR U52256 ( .A(y[1842]), .B(x[1842]), .Z(n42926) );
  XNOR U52257 ( .A(n42927), .B(n42928), .Z(n42925) );
  XNOR U52258 ( .A(y[1843]), .B(x[1843]), .Z(n42928) );
  XNOR U52259 ( .A(y[1844]), .B(x[1844]), .Z(n42927) );
  XNOR U52260 ( .A(n42919), .B(n42920), .Z(n42930) );
  XNOR U52261 ( .A(y[1839]), .B(x[1839]), .Z(n42920) );
  XNOR U52262 ( .A(n42921), .B(n42922), .Z(n42919) );
  XNOR U52263 ( .A(y[1840]), .B(x[1840]), .Z(n42922) );
  XNOR U52264 ( .A(y[1841]), .B(x[1841]), .Z(n42921) );
  NAND U52265 ( .A(n42986), .B(n42987), .Z(N61584) );
  NANDN U52266 ( .A(n42988), .B(n42989), .Z(n42987) );
  OR U52267 ( .A(n42990), .B(n42991), .Z(n42989) );
  NAND U52268 ( .A(n42990), .B(n42991), .Z(n42986) );
  XOR U52269 ( .A(n42990), .B(n42992), .Z(N61583) );
  XNOR U52270 ( .A(n42988), .B(n42991), .Z(n42992) );
  AND U52271 ( .A(n42993), .B(n42994), .Z(n42991) );
  NANDN U52272 ( .A(n42995), .B(n42996), .Z(n42994) );
  NANDN U52273 ( .A(n42997), .B(n42998), .Z(n42996) );
  NANDN U52274 ( .A(n42998), .B(n42997), .Z(n42993) );
  NAND U52275 ( .A(n42999), .B(n43000), .Z(n42988) );
  NANDN U52276 ( .A(n43001), .B(n43002), .Z(n43000) );
  OR U52277 ( .A(n43003), .B(n43004), .Z(n43002) );
  NAND U52278 ( .A(n43004), .B(n43003), .Z(n42999) );
  AND U52279 ( .A(n43005), .B(n43006), .Z(n42990) );
  NANDN U52280 ( .A(n43007), .B(n43008), .Z(n43006) );
  NANDN U52281 ( .A(n43009), .B(n43010), .Z(n43008) );
  NANDN U52282 ( .A(n43010), .B(n43009), .Z(n43005) );
  XOR U52283 ( .A(n43004), .B(n43011), .Z(N61582) );
  XOR U52284 ( .A(n43001), .B(n43003), .Z(n43011) );
  XNOR U52285 ( .A(n42997), .B(n43012), .Z(n43003) );
  XNOR U52286 ( .A(n42995), .B(n42998), .Z(n43012) );
  NAND U52287 ( .A(n43013), .B(n43014), .Z(n42998) );
  NAND U52288 ( .A(n43015), .B(n43016), .Z(n43014) );
  OR U52289 ( .A(n43017), .B(n43018), .Z(n43015) );
  NANDN U52290 ( .A(n43019), .B(n43017), .Z(n43013) );
  IV U52291 ( .A(n43018), .Z(n43019) );
  NAND U52292 ( .A(n43020), .B(n43021), .Z(n42995) );
  NAND U52293 ( .A(n43022), .B(n43023), .Z(n43021) );
  NANDN U52294 ( .A(n43024), .B(n43025), .Z(n43022) );
  NANDN U52295 ( .A(n43025), .B(n43024), .Z(n43020) );
  AND U52296 ( .A(n43026), .B(n43027), .Z(n42997) );
  NAND U52297 ( .A(n43028), .B(n43029), .Z(n43027) );
  OR U52298 ( .A(n43030), .B(n43031), .Z(n43028) );
  NANDN U52299 ( .A(n43032), .B(n43030), .Z(n43026) );
  NAND U52300 ( .A(n43033), .B(n43034), .Z(n43001) );
  NANDN U52301 ( .A(n43035), .B(n43036), .Z(n43034) );
  OR U52302 ( .A(n43037), .B(n43038), .Z(n43036) );
  NANDN U52303 ( .A(n43039), .B(n43037), .Z(n43033) );
  IV U52304 ( .A(n43038), .Z(n43039) );
  XNOR U52305 ( .A(n43009), .B(n43040), .Z(n43004) );
  XNOR U52306 ( .A(n43007), .B(n43010), .Z(n43040) );
  NAND U52307 ( .A(n43041), .B(n43042), .Z(n43010) );
  NAND U52308 ( .A(n43043), .B(n43044), .Z(n43042) );
  OR U52309 ( .A(n43045), .B(n43046), .Z(n43043) );
  NANDN U52310 ( .A(n43047), .B(n43045), .Z(n43041) );
  IV U52311 ( .A(n43046), .Z(n43047) );
  NAND U52312 ( .A(n43048), .B(n43049), .Z(n43007) );
  NAND U52313 ( .A(n43050), .B(n43051), .Z(n43049) );
  NANDN U52314 ( .A(n43052), .B(n43053), .Z(n43050) );
  NANDN U52315 ( .A(n43053), .B(n43052), .Z(n43048) );
  AND U52316 ( .A(n43054), .B(n43055), .Z(n43009) );
  NAND U52317 ( .A(n43056), .B(n43057), .Z(n43055) );
  OR U52318 ( .A(n43058), .B(n43059), .Z(n43056) );
  NANDN U52319 ( .A(n43060), .B(n43058), .Z(n43054) );
  XNOR U52320 ( .A(n43035), .B(n43061), .Z(N61581) );
  XOR U52321 ( .A(n43037), .B(n43038), .Z(n43061) );
  XNOR U52322 ( .A(n43051), .B(n43062), .Z(n43038) );
  XOR U52323 ( .A(n43052), .B(n43053), .Z(n43062) );
  XOR U52324 ( .A(n43058), .B(n43063), .Z(n43053) );
  XOR U52325 ( .A(n43057), .B(n43060), .Z(n43063) );
  IV U52326 ( .A(n43059), .Z(n43060) );
  NAND U52327 ( .A(n43064), .B(n43065), .Z(n43059) );
  OR U52328 ( .A(n43066), .B(n43067), .Z(n43065) );
  OR U52329 ( .A(n43068), .B(n43069), .Z(n43064) );
  NAND U52330 ( .A(n43070), .B(n43071), .Z(n43057) );
  OR U52331 ( .A(n43072), .B(n43073), .Z(n43071) );
  OR U52332 ( .A(n43074), .B(n43075), .Z(n43070) );
  NOR U52333 ( .A(n43076), .B(n43077), .Z(n43058) );
  ANDN U52334 ( .B(n43078), .A(n43079), .Z(n43052) );
  XNOR U52335 ( .A(n43045), .B(n43080), .Z(n43051) );
  XNOR U52336 ( .A(n43044), .B(n43046), .Z(n43080) );
  NAND U52337 ( .A(n43081), .B(n43082), .Z(n43046) );
  OR U52338 ( .A(n43083), .B(n43084), .Z(n43082) );
  OR U52339 ( .A(n43085), .B(n43086), .Z(n43081) );
  NAND U52340 ( .A(n43087), .B(n43088), .Z(n43044) );
  OR U52341 ( .A(n43089), .B(n43090), .Z(n43088) );
  OR U52342 ( .A(n43091), .B(n43092), .Z(n43087) );
  ANDN U52343 ( .B(n43093), .A(n43094), .Z(n43045) );
  IV U52344 ( .A(n43095), .Z(n43093) );
  ANDN U52345 ( .B(n43096), .A(n43097), .Z(n43037) );
  XOR U52346 ( .A(n43023), .B(n43098), .Z(n43035) );
  XOR U52347 ( .A(n43024), .B(n43025), .Z(n43098) );
  XOR U52348 ( .A(n43030), .B(n43099), .Z(n43025) );
  XOR U52349 ( .A(n43029), .B(n43032), .Z(n43099) );
  IV U52350 ( .A(n43031), .Z(n43032) );
  NAND U52351 ( .A(n43100), .B(n43101), .Z(n43031) );
  OR U52352 ( .A(n43102), .B(n43103), .Z(n43101) );
  OR U52353 ( .A(n43104), .B(n43105), .Z(n43100) );
  NAND U52354 ( .A(n43106), .B(n43107), .Z(n43029) );
  OR U52355 ( .A(n43108), .B(n43109), .Z(n43107) );
  OR U52356 ( .A(n43110), .B(n43111), .Z(n43106) );
  NOR U52357 ( .A(n43112), .B(n43113), .Z(n43030) );
  ANDN U52358 ( .B(n43114), .A(n43115), .Z(n43024) );
  IV U52359 ( .A(n43116), .Z(n43114) );
  XNOR U52360 ( .A(n43017), .B(n43117), .Z(n43023) );
  XNOR U52361 ( .A(n43016), .B(n43018), .Z(n43117) );
  NAND U52362 ( .A(n43118), .B(n43119), .Z(n43018) );
  OR U52363 ( .A(n43120), .B(n43121), .Z(n43119) );
  OR U52364 ( .A(n43122), .B(n43123), .Z(n43118) );
  NAND U52365 ( .A(n43124), .B(n43125), .Z(n43016) );
  OR U52366 ( .A(n43126), .B(n43127), .Z(n43125) );
  OR U52367 ( .A(n43128), .B(n43129), .Z(n43124) );
  ANDN U52368 ( .B(n43130), .A(n43131), .Z(n43017) );
  IV U52369 ( .A(n43132), .Z(n43130) );
  XNOR U52370 ( .A(n43097), .B(n43096), .Z(N61580) );
  XOR U52371 ( .A(n43116), .B(n43115), .Z(n43096) );
  XNOR U52372 ( .A(n43131), .B(n43132), .Z(n43115) );
  XNOR U52373 ( .A(n43126), .B(n43127), .Z(n43132) );
  XNOR U52374 ( .A(n43128), .B(n43129), .Z(n43127) );
  XNOR U52375 ( .A(y[1837]), .B(x[1837]), .Z(n43129) );
  XNOR U52376 ( .A(y[1838]), .B(x[1838]), .Z(n43128) );
  XNOR U52377 ( .A(y[1836]), .B(x[1836]), .Z(n43126) );
  XNOR U52378 ( .A(n43120), .B(n43121), .Z(n43131) );
  XNOR U52379 ( .A(y[1833]), .B(x[1833]), .Z(n43121) );
  XNOR U52380 ( .A(n43122), .B(n43123), .Z(n43120) );
  XNOR U52381 ( .A(y[1834]), .B(x[1834]), .Z(n43123) );
  XNOR U52382 ( .A(y[1835]), .B(x[1835]), .Z(n43122) );
  XNOR U52383 ( .A(n43113), .B(n43112), .Z(n43116) );
  XNOR U52384 ( .A(n43108), .B(n43109), .Z(n43112) );
  XNOR U52385 ( .A(y[1830]), .B(x[1830]), .Z(n43109) );
  XNOR U52386 ( .A(n43110), .B(n43111), .Z(n43108) );
  XNOR U52387 ( .A(y[1831]), .B(x[1831]), .Z(n43111) );
  XNOR U52388 ( .A(y[1832]), .B(x[1832]), .Z(n43110) );
  XNOR U52389 ( .A(n43102), .B(n43103), .Z(n43113) );
  XNOR U52390 ( .A(y[1827]), .B(x[1827]), .Z(n43103) );
  XNOR U52391 ( .A(n43104), .B(n43105), .Z(n43102) );
  XNOR U52392 ( .A(y[1828]), .B(x[1828]), .Z(n43105) );
  XNOR U52393 ( .A(y[1829]), .B(x[1829]), .Z(n43104) );
  XOR U52394 ( .A(n43078), .B(n43079), .Z(n43097) );
  XNOR U52395 ( .A(n43094), .B(n43095), .Z(n43079) );
  XNOR U52396 ( .A(n43089), .B(n43090), .Z(n43095) );
  XNOR U52397 ( .A(n43091), .B(n43092), .Z(n43090) );
  XNOR U52398 ( .A(y[1825]), .B(x[1825]), .Z(n43092) );
  XNOR U52399 ( .A(y[1826]), .B(x[1826]), .Z(n43091) );
  XNOR U52400 ( .A(y[1824]), .B(x[1824]), .Z(n43089) );
  XNOR U52401 ( .A(n43083), .B(n43084), .Z(n43094) );
  XNOR U52402 ( .A(y[1821]), .B(x[1821]), .Z(n43084) );
  XNOR U52403 ( .A(n43085), .B(n43086), .Z(n43083) );
  XNOR U52404 ( .A(y[1822]), .B(x[1822]), .Z(n43086) );
  XNOR U52405 ( .A(y[1823]), .B(x[1823]), .Z(n43085) );
  XOR U52406 ( .A(n43077), .B(n43076), .Z(n43078) );
  XNOR U52407 ( .A(n43072), .B(n43073), .Z(n43076) );
  XNOR U52408 ( .A(y[1818]), .B(x[1818]), .Z(n43073) );
  XNOR U52409 ( .A(n43074), .B(n43075), .Z(n43072) );
  XNOR U52410 ( .A(y[1819]), .B(x[1819]), .Z(n43075) );
  XNOR U52411 ( .A(y[1820]), .B(x[1820]), .Z(n43074) );
  XNOR U52412 ( .A(n43066), .B(n43067), .Z(n43077) );
  XNOR U52413 ( .A(y[1815]), .B(x[1815]), .Z(n43067) );
  XNOR U52414 ( .A(n43068), .B(n43069), .Z(n43066) );
  XNOR U52415 ( .A(y[1816]), .B(x[1816]), .Z(n43069) );
  XNOR U52416 ( .A(y[1817]), .B(x[1817]), .Z(n43068) );
  NAND U52417 ( .A(n43133), .B(n43134), .Z(N61571) );
  NANDN U52418 ( .A(n43135), .B(n43136), .Z(n43134) );
  OR U52419 ( .A(n43137), .B(n43138), .Z(n43136) );
  NAND U52420 ( .A(n43137), .B(n43138), .Z(n43133) );
  XOR U52421 ( .A(n43137), .B(n43139), .Z(N61570) );
  XNOR U52422 ( .A(n43135), .B(n43138), .Z(n43139) );
  AND U52423 ( .A(n43140), .B(n43141), .Z(n43138) );
  NANDN U52424 ( .A(n43142), .B(n43143), .Z(n43141) );
  NANDN U52425 ( .A(n43144), .B(n43145), .Z(n43143) );
  NANDN U52426 ( .A(n43145), .B(n43144), .Z(n43140) );
  NAND U52427 ( .A(n43146), .B(n43147), .Z(n43135) );
  NANDN U52428 ( .A(n43148), .B(n43149), .Z(n43147) );
  OR U52429 ( .A(n43150), .B(n43151), .Z(n43149) );
  NAND U52430 ( .A(n43151), .B(n43150), .Z(n43146) );
  AND U52431 ( .A(n43152), .B(n43153), .Z(n43137) );
  NANDN U52432 ( .A(n43154), .B(n43155), .Z(n43153) );
  NANDN U52433 ( .A(n43156), .B(n43157), .Z(n43155) );
  NANDN U52434 ( .A(n43157), .B(n43156), .Z(n43152) );
  XOR U52435 ( .A(n43151), .B(n43158), .Z(N61569) );
  XOR U52436 ( .A(n43148), .B(n43150), .Z(n43158) );
  XNOR U52437 ( .A(n43144), .B(n43159), .Z(n43150) );
  XNOR U52438 ( .A(n43142), .B(n43145), .Z(n43159) );
  NAND U52439 ( .A(n43160), .B(n43161), .Z(n43145) );
  NAND U52440 ( .A(n43162), .B(n43163), .Z(n43161) );
  OR U52441 ( .A(n43164), .B(n43165), .Z(n43162) );
  NANDN U52442 ( .A(n43166), .B(n43164), .Z(n43160) );
  IV U52443 ( .A(n43165), .Z(n43166) );
  NAND U52444 ( .A(n43167), .B(n43168), .Z(n43142) );
  NAND U52445 ( .A(n43169), .B(n43170), .Z(n43168) );
  NANDN U52446 ( .A(n43171), .B(n43172), .Z(n43169) );
  NANDN U52447 ( .A(n43172), .B(n43171), .Z(n43167) );
  AND U52448 ( .A(n43173), .B(n43174), .Z(n43144) );
  NAND U52449 ( .A(n43175), .B(n43176), .Z(n43174) );
  OR U52450 ( .A(n43177), .B(n43178), .Z(n43175) );
  NANDN U52451 ( .A(n43179), .B(n43177), .Z(n43173) );
  NAND U52452 ( .A(n43180), .B(n43181), .Z(n43148) );
  NANDN U52453 ( .A(n43182), .B(n43183), .Z(n43181) );
  OR U52454 ( .A(n43184), .B(n43185), .Z(n43183) );
  NANDN U52455 ( .A(n43186), .B(n43184), .Z(n43180) );
  IV U52456 ( .A(n43185), .Z(n43186) );
  XNOR U52457 ( .A(n43156), .B(n43187), .Z(n43151) );
  XNOR U52458 ( .A(n43154), .B(n43157), .Z(n43187) );
  NAND U52459 ( .A(n43188), .B(n43189), .Z(n43157) );
  NAND U52460 ( .A(n43190), .B(n43191), .Z(n43189) );
  OR U52461 ( .A(n43192), .B(n43193), .Z(n43190) );
  NANDN U52462 ( .A(n43194), .B(n43192), .Z(n43188) );
  IV U52463 ( .A(n43193), .Z(n43194) );
  NAND U52464 ( .A(n43195), .B(n43196), .Z(n43154) );
  NAND U52465 ( .A(n43197), .B(n43198), .Z(n43196) );
  NANDN U52466 ( .A(n43199), .B(n43200), .Z(n43197) );
  NANDN U52467 ( .A(n43200), .B(n43199), .Z(n43195) );
  AND U52468 ( .A(n43201), .B(n43202), .Z(n43156) );
  NAND U52469 ( .A(n43203), .B(n43204), .Z(n43202) );
  OR U52470 ( .A(n43205), .B(n43206), .Z(n43203) );
  NANDN U52471 ( .A(n43207), .B(n43205), .Z(n43201) );
  XNOR U52472 ( .A(n43182), .B(n43208), .Z(N61568) );
  XOR U52473 ( .A(n43184), .B(n43185), .Z(n43208) );
  XNOR U52474 ( .A(n43198), .B(n43209), .Z(n43185) );
  XOR U52475 ( .A(n43199), .B(n43200), .Z(n43209) );
  XOR U52476 ( .A(n43205), .B(n43210), .Z(n43200) );
  XOR U52477 ( .A(n43204), .B(n43207), .Z(n43210) );
  IV U52478 ( .A(n43206), .Z(n43207) );
  NAND U52479 ( .A(n43211), .B(n43212), .Z(n43206) );
  OR U52480 ( .A(n43213), .B(n43214), .Z(n43212) );
  OR U52481 ( .A(n43215), .B(n43216), .Z(n43211) );
  NAND U52482 ( .A(n43217), .B(n43218), .Z(n43204) );
  OR U52483 ( .A(n43219), .B(n43220), .Z(n43218) );
  OR U52484 ( .A(n43221), .B(n43222), .Z(n43217) );
  NOR U52485 ( .A(n43223), .B(n43224), .Z(n43205) );
  ANDN U52486 ( .B(n43225), .A(n43226), .Z(n43199) );
  XNOR U52487 ( .A(n43192), .B(n43227), .Z(n43198) );
  XNOR U52488 ( .A(n43191), .B(n43193), .Z(n43227) );
  NAND U52489 ( .A(n43228), .B(n43229), .Z(n43193) );
  OR U52490 ( .A(n43230), .B(n43231), .Z(n43229) );
  OR U52491 ( .A(n43232), .B(n43233), .Z(n43228) );
  NAND U52492 ( .A(n43234), .B(n43235), .Z(n43191) );
  OR U52493 ( .A(n43236), .B(n43237), .Z(n43235) );
  OR U52494 ( .A(n43238), .B(n43239), .Z(n43234) );
  ANDN U52495 ( .B(n43240), .A(n43241), .Z(n43192) );
  IV U52496 ( .A(n43242), .Z(n43240) );
  ANDN U52497 ( .B(n43243), .A(n43244), .Z(n43184) );
  XOR U52498 ( .A(n43170), .B(n43245), .Z(n43182) );
  XOR U52499 ( .A(n43171), .B(n43172), .Z(n43245) );
  XOR U52500 ( .A(n43177), .B(n43246), .Z(n43172) );
  XOR U52501 ( .A(n43176), .B(n43179), .Z(n43246) );
  IV U52502 ( .A(n43178), .Z(n43179) );
  NAND U52503 ( .A(n43247), .B(n43248), .Z(n43178) );
  OR U52504 ( .A(n43249), .B(n43250), .Z(n43248) );
  OR U52505 ( .A(n43251), .B(n43252), .Z(n43247) );
  NAND U52506 ( .A(n43253), .B(n43254), .Z(n43176) );
  OR U52507 ( .A(n43255), .B(n43256), .Z(n43254) );
  OR U52508 ( .A(n43257), .B(n43258), .Z(n43253) );
  NOR U52509 ( .A(n43259), .B(n43260), .Z(n43177) );
  ANDN U52510 ( .B(n43261), .A(n43262), .Z(n43171) );
  IV U52511 ( .A(n43263), .Z(n43261) );
  XNOR U52512 ( .A(n43164), .B(n43264), .Z(n43170) );
  XNOR U52513 ( .A(n43163), .B(n43165), .Z(n43264) );
  NAND U52514 ( .A(n43265), .B(n43266), .Z(n43165) );
  OR U52515 ( .A(n43267), .B(n43268), .Z(n43266) );
  OR U52516 ( .A(n43269), .B(n43270), .Z(n43265) );
  NAND U52517 ( .A(n43271), .B(n43272), .Z(n43163) );
  OR U52518 ( .A(n43273), .B(n43274), .Z(n43272) );
  OR U52519 ( .A(n43275), .B(n43276), .Z(n43271) );
  ANDN U52520 ( .B(n43277), .A(n43278), .Z(n43164) );
  IV U52521 ( .A(n43279), .Z(n43277) );
  XNOR U52522 ( .A(n43244), .B(n43243), .Z(N61567) );
  XOR U52523 ( .A(n43263), .B(n43262), .Z(n43243) );
  XNOR U52524 ( .A(n43278), .B(n43279), .Z(n43262) );
  XNOR U52525 ( .A(n43273), .B(n43274), .Z(n43279) );
  XNOR U52526 ( .A(n43275), .B(n43276), .Z(n43274) );
  XNOR U52527 ( .A(y[1813]), .B(x[1813]), .Z(n43276) );
  XNOR U52528 ( .A(y[1814]), .B(x[1814]), .Z(n43275) );
  XNOR U52529 ( .A(y[1812]), .B(x[1812]), .Z(n43273) );
  XNOR U52530 ( .A(n43267), .B(n43268), .Z(n43278) );
  XNOR U52531 ( .A(y[1809]), .B(x[1809]), .Z(n43268) );
  XNOR U52532 ( .A(n43269), .B(n43270), .Z(n43267) );
  XNOR U52533 ( .A(y[1810]), .B(x[1810]), .Z(n43270) );
  XNOR U52534 ( .A(y[1811]), .B(x[1811]), .Z(n43269) );
  XNOR U52535 ( .A(n43260), .B(n43259), .Z(n43263) );
  XNOR U52536 ( .A(n43255), .B(n43256), .Z(n43259) );
  XNOR U52537 ( .A(y[1806]), .B(x[1806]), .Z(n43256) );
  XNOR U52538 ( .A(n43257), .B(n43258), .Z(n43255) );
  XNOR U52539 ( .A(y[1807]), .B(x[1807]), .Z(n43258) );
  XNOR U52540 ( .A(y[1808]), .B(x[1808]), .Z(n43257) );
  XNOR U52541 ( .A(n43249), .B(n43250), .Z(n43260) );
  XNOR U52542 ( .A(y[1803]), .B(x[1803]), .Z(n43250) );
  XNOR U52543 ( .A(n43251), .B(n43252), .Z(n43249) );
  XNOR U52544 ( .A(y[1804]), .B(x[1804]), .Z(n43252) );
  XNOR U52545 ( .A(y[1805]), .B(x[1805]), .Z(n43251) );
  XOR U52546 ( .A(n43225), .B(n43226), .Z(n43244) );
  XNOR U52547 ( .A(n43241), .B(n43242), .Z(n43226) );
  XNOR U52548 ( .A(n43236), .B(n43237), .Z(n43242) );
  XNOR U52549 ( .A(n43238), .B(n43239), .Z(n43237) );
  XNOR U52550 ( .A(y[1801]), .B(x[1801]), .Z(n43239) );
  XNOR U52551 ( .A(y[1802]), .B(x[1802]), .Z(n43238) );
  XNOR U52552 ( .A(y[1800]), .B(x[1800]), .Z(n43236) );
  XNOR U52553 ( .A(n43230), .B(n43231), .Z(n43241) );
  XNOR U52554 ( .A(y[1797]), .B(x[1797]), .Z(n43231) );
  XNOR U52555 ( .A(n43232), .B(n43233), .Z(n43230) );
  XNOR U52556 ( .A(y[1798]), .B(x[1798]), .Z(n43233) );
  XNOR U52557 ( .A(y[1799]), .B(x[1799]), .Z(n43232) );
  XOR U52558 ( .A(n43224), .B(n43223), .Z(n43225) );
  XNOR U52559 ( .A(n43219), .B(n43220), .Z(n43223) );
  XNOR U52560 ( .A(y[1794]), .B(x[1794]), .Z(n43220) );
  XNOR U52561 ( .A(n43221), .B(n43222), .Z(n43219) );
  XNOR U52562 ( .A(y[1795]), .B(x[1795]), .Z(n43222) );
  XNOR U52563 ( .A(y[1796]), .B(x[1796]), .Z(n43221) );
  XNOR U52564 ( .A(n43213), .B(n43214), .Z(n43224) );
  XNOR U52565 ( .A(y[1791]), .B(x[1791]), .Z(n43214) );
  XNOR U52566 ( .A(n43215), .B(n43216), .Z(n43213) );
  XNOR U52567 ( .A(y[1792]), .B(x[1792]), .Z(n43216) );
  XNOR U52568 ( .A(y[1793]), .B(x[1793]), .Z(n43215) );
  NAND U52569 ( .A(n43280), .B(n43281), .Z(N61558) );
  NANDN U52570 ( .A(n43282), .B(n43283), .Z(n43281) );
  OR U52571 ( .A(n43284), .B(n43285), .Z(n43283) );
  NAND U52572 ( .A(n43284), .B(n43285), .Z(n43280) );
  XOR U52573 ( .A(n43284), .B(n43286), .Z(N61557) );
  XNOR U52574 ( .A(n43282), .B(n43285), .Z(n43286) );
  AND U52575 ( .A(n43287), .B(n43288), .Z(n43285) );
  NANDN U52576 ( .A(n43289), .B(n43290), .Z(n43288) );
  NANDN U52577 ( .A(n43291), .B(n43292), .Z(n43290) );
  NANDN U52578 ( .A(n43292), .B(n43291), .Z(n43287) );
  NAND U52579 ( .A(n43293), .B(n43294), .Z(n43282) );
  NANDN U52580 ( .A(n43295), .B(n43296), .Z(n43294) );
  OR U52581 ( .A(n43297), .B(n43298), .Z(n43296) );
  NAND U52582 ( .A(n43298), .B(n43297), .Z(n43293) );
  AND U52583 ( .A(n43299), .B(n43300), .Z(n43284) );
  NANDN U52584 ( .A(n43301), .B(n43302), .Z(n43300) );
  NANDN U52585 ( .A(n43303), .B(n43304), .Z(n43302) );
  NANDN U52586 ( .A(n43304), .B(n43303), .Z(n43299) );
  XOR U52587 ( .A(n43298), .B(n43305), .Z(N61556) );
  XOR U52588 ( .A(n43295), .B(n43297), .Z(n43305) );
  XNOR U52589 ( .A(n43291), .B(n43306), .Z(n43297) );
  XNOR U52590 ( .A(n43289), .B(n43292), .Z(n43306) );
  NAND U52591 ( .A(n43307), .B(n43308), .Z(n43292) );
  NAND U52592 ( .A(n43309), .B(n43310), .Z(n43308) );
  OR U52593 ( .A(n43311), .B(n43312), .Z(n43309) );
  NANDN U52594 ( .A(n43313), .B(n43311), .Z(n43307) );
  IV U52595 ( .A(n43312), .Z(n43313) );
  NAND U52596 ( .A(n43314), .B(n43315), .Z(n43289) );
  NAND U52597 ( .A(n43316), .B(n43317), .Z(n43315) );
  NANDN U52598 ( .A(n43318), .B(n43319), .Z(n43316) );
  NANDN U52599 ( .A(n43319), .B(n43318), .Z(n43314) );
  AND U52600 ( .A(n43320), .B(n43321), .Z(n43291) );
  NAND U52601 ( .A(n43322), .B(n43323), .Z(n43321) );
  OR U52602 ( .A(n43324), .B(n43325), .Z(n43322) );
  NANDN U52603 ( .A(n43326), .B(n43324), .Z(n43320) );
  NAND U52604 ( .A(n43327), .B(n43328), .Z(n43295) );
  NANDN U52605 ( .A(n43329), .B(n43330), .Z(n43328) );
  OR U52606 ( .A(n43331), .B(n43332), .Z(n43330) );
  NANDN U52607 ( .A(n43333), .B(n43331), .Z(n43327) );
  IV U52608 ( .A(n43332), .Z(n43333) );
  XNOR U52609 ( .A(n43303), .B(n43334), .Z(n43298) );
  XNOR U52610 ( .A(n43301), .B(n43304), .Z(n43334) );
  NAND U52611 ( .A(n43335), .B(n43336), .Z(n43304) );
  NAND U52612 ( .A(n43337), .B(n43338), .Z(n43336) );
  OR U52613 ( .A(n43339), .B(n43340), .Z(n43337) );
  NANDN U52614 ( .A(n43341), .B(n43339), .Z(n43335) );
  IV U52615 ( .A(n43340), .Z(n43341) );
  NAND U52616 ( .A(n43342), .B(n43343), .Z(n43301) );
  NAND U52617 ( .A(n43344), .B(n43345), .Z(n43343) );
  NANDN U52618 ( .A(n43346), .B(n43347), .Z(n43344) );
  NANDN U52619 ( .A(n43347), .B(n43346), .Z(n43342) );
  AND U52620 ( .A(n43348), .B(n43349), .Z(n43303) );
  NAND U52621 ( .A(n43350), .B(n43351), .Z(n43349) );
  OR U52622 ( .A(n43352), .B(n43353), .Z(n43350) );
  NANDN U52623 ( .A(n43354), .B(n43352), .Z(n43348) );
  XNOR U52624 ( .A(n43329), .B(n43355), .Z(N61555) );
  XOR U52625 ( .A(n43331), .B(n43332), .Z(n43355) );
  XNOR U52626 ( .A(n43345), .B(n43356), .Z(n43332) );
  XOR U52627 ( .A(n43346), .B(n43347), .Z(n43356) );
  XOR U52628 ( .A(n43352), .B(n43357), .Z(n43347) );
  XOR U52629 ( .A(n43351), .B(n43354), .Z(n43357) );
  IV U52630 ( .A(n43353), .Z(n43354) );
  NAND U52631 ( .A(n43358), .B(n43359), .Z(n43353) );
  OR U52632 ( .A(n43360), .B(n43361), .Z(n43359) );
  OR U52633 ( .A(n43362), .B(n43363), .Z(n43358) );
  NAND U52634 ( .A(n43364), .B(n43365), .Z(n43351) );
  OR U52635 ( .A(n43366), .B(n43367), .Z(n43365) );
  OR U52636 ( .A(n43368), .B(n43369), .Z(n43364) );
  NOR U52637 ( .A(n43370), .B(n43371), .Z(n43352) );
  ANDN U52638 ( .B(n43372), .A(n43373), .Z(n43346) );
  XNOR U52639 ( .A(n43339), .B(n43374), .Z(n43345) );
  XNOR U52640 ( .A(n43338), .B(n43340), .Z(n43374) );
  NAND U52641 ( .A(n43375), .B(n43376), .Z(n43340) );
  OR U52642 ( .A(n43377), .B(n43378), .Z(n43376) );
  OR U52643 ( .A(n43379), .B(n43380), .Z(n43375) );
  NAND U52644 ( .A(n43381), .B(n43382), .Z(n43338) );
  OR U52645 ( .A(n43383), .B(n43384), .Z(n43382) );
  OR U52646 ( .A(n43385), .B(n43386), .Z(n43381) );
  ANDN U52647 ( .B(n43387), .A(n43388), .Z(n43339) );
  IV U52648 ( .A(n43389), .Z(n43387) );
  ANDN U52649 ( .B(n43390), .A(n43391), .Z(n43331) );
  XOR U52650 ( .A(n43317), .B(n43392), .Z(n43329) );
  XOR U52651 ( .A(n43318), .B(n43319), .Z(n43392) );
  XOR U52652 ( .A(n43324), .B(n43393), .Z(n43319) );
  XOR U52653 ( .A(n43323), .B(n43326), .Z(n43393) );
  IV U52654 ( .A(n43325), .Z(n43326) );
  NAND U52655 ( .A(n43394), .B(n43395), .Z(n43325) );
  OR U52656 ( .A(n43396), .B(n43397), .Z(n43395) );
  OR U52657 ( .A(n43398), .B(n43399), .Z(n43394) );
  NAND U52658 ( .A(n43400), .B(n43401), .Z(n43323) );
  OR U52659 ( .A(n43402), .B(n43403), .Z(n43401) );
  OR U52660 ( .A(n43404), .B(n43405), .Z(n43400) );
  NOR U52661 ( .A(n43406), .B(n43407), .Z(n43324) );
  ANDN U52662 ( .B(n43408), .A(n43409), .Z(n43318) );
  IV U52663 ( .A(n43410), .Z(n43408) );
  XNOR U52664 ( .A(n43311), .B(n43411), .Z(n43317) );
  XNOR U52665 ( .A(n43310), .B(n43312), .Z(n43411) );
  NAND U52666 ( .A(n43412), .B(n43413), .Z(n43312) );
  OR U52667 ( .A(n43414), .B(n43415), .Z(n43413) );
  OR U52668 ( .A(n43416), .B(n43417), .Z(n43412) );
  NAND U52669 ( .A(n43418), .B(n43419), .Z(n43310) );
  OR U52670 ( .A(n43420), .B(n43421), .Z(n43419) );
  OR U52671 ( .A(n43422), .B(n43423), .Z(n43418) );
  ANDN U52672 ( .B(n43424), .A(n43425), .Z(n43311) );
  IV U52673 ( .A(n43426), .Z(n43424) );
  XNOR U52674 ( .A(n43391), .B(n43390), .Z(N61554) );
  XOR U52675 ( .A(n43410), .B(n43409), .Z(n43390) );
  XNOR U52676 ( .A(n43425), .B(n43426), .Z(n43409) );
  XNOR U52677 ( .A(n43420), .B(n43421), .Z(n43426) );
  XNOR U52678 ( .A(n43422), .B(n43423), .Z(n43421) );
  XNOR U52679 ( .A(y[1789]), .B(x[1789]), .Z(n43423) );
  XNOR U52680 ( .A(y[1790]), .B(x[1790]), .Z(n43422) );
  XNOR U52681 ( .A(y[1788]), .B(x[1788]), .Z(n43420) );
  XNOR U52682 ( .A(n43414), .B(n43415), .Z(n43425) );
  XNOR U52683 ( .A(y[1785]), .B(x[1785]), .Z(n43415) );
  XNOR U52684 ( .A(n43416), .B(n43417), .Z(n43414) );
  XNOR U52685 ( .A(y[1786]), .B(x[1786]), .Z(n43417) );
  XNOR U52686 ( .A(y[1787]), .B(x[1787]), .Z(n43416) );
  XNOR U52687 ( .A(n43407), .B(n43406), .Z(n43410) );
  XNOR U52688 ( .A(n43402), .B(n43403), .Z(n43406) );
  XNOR U52689 ( .A(y[1782]), .B(x[1782]), .Z(n43403) );
  XNOR U52690 ( .A(n43404), .B(n43405), .Z(n43402) );
  XNOR U52691 ( .A(y[1783]), .B(x[1783]), .Z(n43405) );
  XNOR U52692 ( .A(y[1784]), .B(x[1784]), .Z(n43404) );
  XNOR U52693 ( .A(n43396), .B(n43397), .Z(n43407) );
  XNOR U52694 ( .A(y[1779]), .B(x[1779]), .Z(n43397) );
  XNOR U52695 ( .A(n43398), .B(n43399), .Z(n43396) );
  XNOR U52696 ( .A(y[1780]), .B(x[1780]), .Z(n43399) );
  XNOR U52697 ( .A(y[1781]), .B(x[1781]), .Z(n43398) );
  XOR U52698 ( .A(n43372), .B(n43373), .Z(n43391) );
  XNOR U52699 ( .A(n43388), .B(n43389), .Z(n43373) );
  XNOR U52700 ( .A(n43383), .B(n43384), .Z(n43389) );
  XNOR U52701 ( .A(n43385), .B(n43386), .Z(n43384) );
  XNOR U52702 ( .A(y[1777]), .B(x[1777]), .Z(n43386) );
  XNOR U52703 ( .A(y[1778]), .B(x[1778]), .Z(n43385) );
  XNOR U52704 ( .A(y[1776]), .B(x[1776]), .Z(n43383) );
  XNOR U52705 ( .A(n43377), .B(n43378), .Z(n43388) );
  XNOR U52706 ( .A(y[1773]), .B(x[1773]), .Z(n43378) );
  XNOR U52707 ( .A(n43379), .B(n43380), .Z(n43377) );
  XNOR U52708 ( .A(y[1774]), .B(x[1774]), .Z(n43380) );
  XNOR U52709 ( .A(y[1775]), .B(x[1775]), .Z(n43379) );
  XOR U52710 ( .A(n43371), .B(n43370), .Z(n43372) );
  XNOR U52711 ( .A(n43366), .B(n43367), .Z(n43370) );
  XNOR U52712 ( .A(y[1770]), .B(x[1770]), .Z(n43367) );
  XNOR U52713 ( .A(n43368), .B(n43369), .Z(n43366) );
  XNOR U52714 ( .A(y[1771]), .B(x[1771]), .Z(n43369) );
  XNOR U52715 ( .A(y[1772]), .B(x[1772]), .Z(n43368) );
  XNOR U52716 ( .A(n43360), .B(n43361), .Z(n43371) );
  XNOR U52717 ( .A(y[1767]), .B(x[1767]), .Z(n43361) );
  XNOR U52718 ( .A(n43362), .B(n43363), .Z(n43360) );
  XNOR U52719 ( .A(y[1768]), .B(x[1768]), .Z(n43363) );
  XNOR U52720 ( .A(y[1769]), .B(x[1769]), .Z(n43362) );
  NAND U52721 ( .A(n43427), .B(n43428), .Z(N61545) );
  NANDN U52722 ( .A(n43429), .B(n43430), .Z(n43428) );
  OR U52723 ( .A(n43431), .B(n43432), .Z(n43430) );
  NAND U52724 ( .A(n43431), .B(n43432), .Z(n43427) );
  XOR U52725 ( .A(n43431), .B(n43433), .Z(N61544) );
  XNOR U52726 ( .A(n43429), .B(n43432), .Z(n43433) );
  AND U52727 ( .A(n43434), .B(n43435), .Z(n43432) );
  NANDN U52728 ( .A(n43436), .B(n43437), .Z(n43435) );
  NANDN U52729 ( .A(n43438), .B(n43439), .Z(n43437) );
  NANDN U52730 ( .A(n43439), .B(n43438), .Z(n43434) );
  NAND U52731 ( .A(n43440), .B(n43441), .Z(n43429) );
  NANDN U52732 ( .A(n43442), .B(n43443), .Z(n43441) );
  OR U52733 ( .A(n43444), .B(n43445), .Z(n43443) );
  NAND U52734 ( .A(n43445), .B(n43444), .Z(n43440) );
  AND U52735 ( .A(n43446), .B(n43447), .Z(n43431) );
  NANDN U52736 ( .A(n43448), .B(n43449), .Z(n43447) );
  NANDN U52737 ( .A(n43450), .B(n43451), .Z(n43449) );
  NANDN U52738 ( .A(n43451), .B(n43450), .Z(n43446) );
  XOR U52739 ( .A(n43445), .B(n43452), .Z(N61543) );
  XOR U52740 ( .A(n43442), .B(n43444), .Z(n43452) );
  XNOR U52741 ( .A(n43438), .B(n43453), .Z(n43444) );
  XNOR U52742 ( .A(n43436), .B(n43439), .Z(n43453) );
  NAND U52743 ( .A(n43454), .B(n43455), .Z(n43439) );
  NAND U52744 ( .A(n43456), .B(n43457), .Z(n43455) );
  OR U52745 ( .A(n43458), .B(n43459), .Z(n43456) );
  NANDN U52746 ( .A(n43460), .B(n43458), .Z(n43454) );
  IV U52747 ( .A(n43459), .Z(n43460) );
  NAND U52748 ( .A(n43461), .B(n43462), .Z(n43436) );
  NAND U52749 ( .A(n43463), .B(n43464), .Z(n43462) );
  NANDN U52750 ( .A(n43465), .B(n43466), .Z(n43463) );
  NANDN U52751 ( .A(n43466), .B(n43465), .Z(n43461) );
  AND U52752 ( .A(n43467), .B(n43468), .Z(n43438) );
  NAND U52753 ( .A(n43469), .B(n43470), .Z(n43468) );
  OR U52754 ( .A(n43471), .B(n43472), .Z(n43469) );
  NANDN U52755 ( .A(n43473), .B(n43471), .Z(n43467) );
  NAND U52756 ( .A(n43474), .B(n43475), .Z(n43442) );
  NANDN U52757 ( .A(n43476), .B(n43477), .Z(n43475) );
  OR U52758 ( .A(n43478), .B(n43479), .Z(n43477) );
  NANDN U52759 ( .A(n43480), .B(n43478), .Z(n43474) );
  IV U52760 ( .A(n43479), .Z(n43480) );
  XNOR U52761 ( .A(n43450), .B(n43481), .Z(n43445) );
  XNOR U52762 ( .A(n43448), .B(n43451), .Z(n43481) );
  NAND U52763 ( .A(n43482), .B(n43483), .Z(n43451) );
  NAND U52764 ( .A(n43484), .B(n43485), .Z(n43483) );
  OR U52765 ( .A(n43486), .B(n43487), .Z(n43484) );
  NANDN U52766 ( .A(n43488), .B(n43486), .Z(n43482) );
  IV U52767 ( .A(n43487), .Z(n43488) );
  NAND U52768 ( .A(n43489), .B(n43490), .Z(n43448) );
  NAND U52769 ( .A(n43491), .B(n43492), .Z(n43490) );
  NANDN U52770 ( .A(n43493), .B(n43494), .Z(n43491) );
  NANDN U52771 ( .A(n43494), .B(n43493), .Z(n43489) );
  AND U52772 ( .A(n43495), .B(n43496), .Z(n43450) );
  NAND U52773 ( .A(n43497), .B(n43498), .Z(n43496) );
  OR U52774 ( .A(n43499), .B(n43500), .Z(n43497) );
  NANDN U52775 ( .A(n43501), .B(n43499), .Z(n43495) );
  XNOR U52776 ( .A(n43476), .B(n43502), .Z(N61542) );
  XOR U52777 ( .A(n43478), .B(n43479), .Z(n43502) );
  XNOR U52778 ( .A(n43492), .B(n43503), .Z(n43479) );
  XOR U52779 ( .A(n43493), .B(n43494), .Z(n43503) );
  XOR U52780 ( .A(n43499), .B(n43504), .Z(n43494) );
  XOR U52781 ( .A(n43498), .B(n43501), .Z(n43504) );
  IV U52782 ( .A(n43500), .Z(n43501) );
  NAND U52783 ( .A(n43505), .B(n43506), .Z(n43500) );
  OR U52784 ( .A(n43507), .B(n43508), .Z(n43506) );
  OR U52785 ( .A(n43509), .B(n43510), .Z(n43505) );
  NAND U52786 ( .A(n43511), .B(n43512), .Z(n43498) );
  OR U52787 ( .A(n43513), .B(n43514), .Z(n43512) );
  OR U52788 ( .A(n43515), .B(n43516), .Z(n43511) );
  NOR U52789 ( .A(n43517), .B(n43518), .Z(n43499) );
  ANDN U52790 ( .B(n43519), .A(n43520), .Z(n43493) );
  XNOR U52791 ( .A(n43486), .B(n43521), .Z(n43492) );
  XNOR U52792 ( .A(n43485), .B(n43487), .Z(n43521) );
  NAND U52793 ( .A(n43522), .B(n43523), .Z(n43487) );
  OR U52794 ( .A(n43524), .B(n43525), .Z(n43523) );
  OR U52795 ( .A(n43526), .B(n43527), .Z(n43522) );
  NAND U52796 ( .A(n43528), .B(n43529), .Z(n43485) );
  OR U52797 ( .A(n43530), .B(n43531), .Z(n43529) );
  OR U52798 ( .A(n43532), .B(n43533), .Z(n43528) );
  ANDN U52799 ( .B(n43534), .A(n43535), .Z(n43486) );
  IV U52800 ( .A(n43536), .Z(n43534) );
  ANDN U52801 ( .B(n43537), .A(n43538), .Z(n43478) );
  XOR U52802 ( .A(n43464), .B(n43539), .Z(n43476) );
  XOR U52803 ( .A(n43465), .B(n43466), .Z(n43539) );
  XOR U52804 ( .A(n43471), .B(n43540), .Z(n43466) );
  XOR U52805 ( .A(n43470), .B(n43473), .Z(n43540) );
  IV U52806 ( .A(n43472), .Z(n43473) );
  NAND U52807 ( .A(n43541), .B(n43542), .Z(n43472) );
  OR U52808 ( .A(n43543), .B(n43544), .Z(n43542) );
  OR U52809 ( .A(n43545), .B(n43546), .Z(n43541) );
  NAND U52810 ( .A(n43547), .B(n43548), .Z(n43470) );
  OR U52811 ( .A(n43549), .B(n43550), .Z(n43548) );
  OR U52812 ( .A(n43551), .B(n43552), .Z(n43547) );
  NOR U52813 ( .A(n43553), .B(n43554), .Z(n43471) );
  ANDN U52814 ( .B(n43555), .A(n43556), .Z(n43465) );
  IV U52815 ( .A(n43557), .Z(n43555) );
  XNOR U52816 ( .A(n43458), .B(n43558), .Z(n43464) );
  XNOR U52817 ( .A(n43457), .B(n43459), .Z(n43558) );
  NAND U52818 ( .A(n43559), .B(n43560), .Z(n43459) );
  OR U52819 ( .A(n43561), .B(n43562), .Z(n43560) );
  OR U52820 ( .A(n43563), .B(n43564), .Z(n43559) );
  NAND U52821 ( .A(n43565), .B(n43566), .Z(n43457) );
  OR U52822 ( .A(n43567), .B(n43568), .Z(n43566) );
  OR U52823 ( .A(n43569), .B(n43570), .Z(n43565) );
  ANDN U52824 ( .B(n43571), .A(n43572), .Z(n43458) );
  IV U52825 ( .A(n43573), .Z(n43571) );
  XNOR U52826 ( .A(n43538), .B(n43537), .Z(N61541) );
  XOR U52827 ( .A(n43557), .B(n43556), .Z(n43537) );
  XNOR U52828 ( .A(n43572), .B(n43573), .Z(n43556) );
  XNOR U52829 ( .A(n43567), .B(n43568), .Z(n43573) );
  XNOR U52830 ( .A(n43569), .B(n43570), .Z(n43568) );
  XNOR U52831 ( .A(y[1765]), .B(x[1765]), .Z(n43570) );
  XNOR U52832 ( .A(y[1766]), .B(x[1766]), .Z(n43569) );
  XNOR U52833 ( .A(y[1764]), .B(x[1764]), .Z(n43567) );
  XNOR U52834 ( .A(n43561), .B(n43562), .Z(n43572) );
  XNOR U52835 ( .A(y[1761]), .B(x[1761]), .Z(n43562) );
  XNOR U52836 ( .A(n43563), .B(n43564), .Z(n43561) );
  XNOR U52837 ( .A(y[1762]), .B(x[1762]), .Z(n43564) );
  XNOR U52838 ( .A(y[1763]), .B(x[1763]), .Z(n43563) );
  XNOR U52839 ( .A(n43554), .B(n43553), .Z(n43557) );
  XNOR U52840 ( .A(n43549), .B(n43550), .Z(n43553) );
  XNOR U52841 ( .A(y[1758]), .B(x[1758]), .Z(n43550) );
  XNOR U52842 ( .A(n43551), .B(n43552), .Z(n43549) );
  XNOR U52843 ( .A(y[1759]), .B(x[1759]), .Z(n43552) );
  XNOR U52844 ( .A(y[1760]), .B(x[1760]), .Z(n43551) );
  XNOR U52845 ( .A(n43543), .B(n43544), .Z(n43554) );
  XNOR U52846 ( .A(y[1755]), .B(x[1755]), .Z(n43544) );
  XNOR U52847 ( .A(n43545), .B(n43546), .Z(n43543) );
  XNOR U52848 ( .A(y[1756]), .B(x[1756]), .Z(n43546) );
  XNOR U52849 ( .A(y[1757]), .B(x[1757]), .Z(n43545) );
  XOR U52850 ( .A(n43519), .B(n43520), .Z(n43538) );
  XNOR U52851 ( .A(n43535), .B(n43536), .Z(n43520) );
  XNOR U52852 ( .A(n43530), .B(n43531), .Z(n43536) );
  XNOR U52853 ( .A(n43532), .B(n43533), .Z(n43531) );
  XNOR U52854 ( .A(y[1753]), .B(x[1753]), .Z(n43533) );
  XNOR U52855 ( .A(y[1754]), .B(x[1754]), .Z(n43532) );
  XNOR U52856 ( .A(y[1752]), .B(x[1752]), .Z(n43530) );
  XNOR U52857 ( .A(n43524), .B(n43525), .Z(n43535) );
  XNOR U52858 ( .A(y[1749]), .B(x[1749]), .Z(n43525) );
  XNOR U52859 ( .A(n43526), .B(n43527), .Z(n43524) );
  XNOR U52860 ( .A(y[1750]), .B(x[1750]), .Z(n43527) );
  XNOR U52861 ( .A(y[1751]), .B(x[1751]), .Z(n43526) );
  XOR U52862 ( .A(n43518), .B(n43517), .Z(n43519) );
  XNOR U52863 ( .A(n43513), .B(n43514), .Z(n43517) );
  XNOR U52864 ( .A(y[1746]), .B(x[1746]), .Z(n43514) );
  XNOR U52865 ( .A(n43515), .B(n43516), .Z(n43513) );
  XNOR U52866 ( .A(y[1747]), .B(x[1747]), .Z(n43516) );
  XNOR U52867 ( .A(y[1748]), .B(x[1748]), .Z(n43515) );
  XNOR U52868 ( .A(n43507), .B(n43508), .Z(n43518) );
  XNOR U52869 ( .A(y[1743]), .B(x[1743]), .Z(n43508) );
  XNOR U52870 ( .A(n43509), .B(n43510), .Z(n43507) );
  XNOR U52871 ( .A(y[1744]), .B(x[1744]), .Z(n43510) );
  XNOR U52872 ( .A(y[1745]), .B(x[1745]), .Z(n43509) );
  NAND U52873 ( .A(n43574), .B(n43575), .Z(N61532) );
  NANDN U52874 ( .A(n43576), .B(n43577), .Z(n43575) );
  OR U52875 ( .A(n43578), .B(n43579), .Z(n43577) );
  NAND U52876 ( .A(n43578), .B(n43579), .Z(n43574) );
  XOR U52877 ( .A(n43578), .B(n43580), .Z(N61531) );
  XNOR U52878 ( .A(n43576), .B(n43579), .Z(n43580) );
  AND U52879 ( .A(n43581), .B(n43582), .Z(n43579) );
  NANDN U52880 ( .A(n43583), .B(n43584), .Z(n43582) );
  NANDN U52881 ( .A(n43585), .B(n43586), .Z(n43584) );
  NANDN U52882 ( .A(n43586), .B(n43585), .Z(n43581) );
  NAND U52883 ( .A(n43587), .B(n43588), .Z(n43576) );
  NANDN U52884 ( .A(n43589), .B(n43590), .Z(n43588) );
  OR U52885 ( .A(n43591), .B(n43592), .Z(n43590) );
  NAND U52886 ( .A(n43592), .B(n43591), .Z(n43587) );
  AND U52887 ( .A(n43593), .B(n43594), .Z(n43578) );
  NANDN U52888 ( .A(n43595), .B(n43596), .Z(n43594) );
  NANDN U52889 ( .A(n43597), .B(n43598), .Z(n43596) );
  NANDN U52890 ( .A(n43598), .B(n43597), .Z(n43593) );
  XOR U52891 ( .A(n43592), .B(n43599), .Z(N61530) );
  XOR U52892 ( .A(n43589), .B(n43591), .Z(n43599) );
  XNOR U52893 ( .A(n43585), .B(n43600), .Z(n43591) );
  XNOR U52894 ( .A(n43583), .B(n43586), .Z(n43600) );
  NAND U52895 ( .A(n43601), .B(n43602), .Z(n43586) );
  NAND U52896 ( .A(n43603), .B(n43604), .Z(n43602) );
  OR U52897 ( .A(n43605), .B(n43606), .Z(n43603) );
  NANDN U52898 ( .A(n43607), .B(n43605), .Z(n43601) );
  IV U52899 ( .A(n43606), .Z(n43607) );
  NAND U52900 ( .A(n43608), .B(n43609), .Z(n43583) );
  NAND U52901 ( .A(n43610), .B(n43611), .Z(n43609) );
  NANDN U52902 ( .A(n43612), .B(n43613), .Z(n43610) );
  NANDN U52903 ( .A(n43613), .B(n43612), .Z(n43608) );
  AND U52904 ( .A(n43614), .B(n43615), .Z(n43585) );
  NAND U52905 ( .A(n43616), .B(n43617), .Z(n43615) );
  OR U52906 ( .A(n43618), .B(n43619), .Z(n43616) );
  NANDN U52907 ( .A(n43620), .B(n43618), .Z(n43614) );
  NAND U52908 ( .A(n43621), .B(n43622), .Z(n43589) );
  NANDN U52909 ( .A(n43623), .B(n43624), .Z(n43622) );
  OR U52910 ( .A(n43625), .B(n43626), .Z(n43624) );
  NANDN U52911 ( .A(n43627), .B(n43625), .Z(n43621) );
  IV U52912 ( .A(n43626), .Z(n43627) );
  XNOR U52913 ( .A(n43597), .B(n43628), .Z(n43592) );
  XNOR U52914 ( .A(n43595), .B(n43598), .Z(n43628) );
  NAND U52915 ( .A(n43629), .B(n43630), .Z(n43598) );
  NAND U52916 ( .A(n43631), .B(n43632), .Z(n43630) );
  OR U52917 ( .A(n43633), .B(n43634), .Z(n43631) );
  NANDN U52918 ( .A(n43635), .B(n43633), .Z(n43629) );
  IV U52919 ( .A(n43634), .Z(n43635) );
  NAND U52920 ( .A(n43636), .B(n43637), .Z(n43595) );
  NAND U52921 ( .A(n43638), .B(n43639), .Z(n43637) );
  NANDN U52922 ( .A(n43640), .B(n43641), .Z(n43638) );
  NANDN U52923 ( .A(n43641), .B(n43640), .Z(n43636) );
  AND U52924 ( .A(n43642), .B(n43643), .Z(n43597) );
  NAND U52925 ( .A(n43644), .B(n43645), .Z(n43643) );
  OR U52926 ( .A(n43646), .B(n43647), .Z(n43644) );
  NANDN U52927 ( .A(n43648), .B(n43646), .Z(n43642) );
  XNOR U52928 ( .A(n43623), .B(n43649), .Z(N61529) );
  XOR U52929 ( .A(n43625), .B(n43626), .Z(n43649) );
  XNOR U52930 ( .A(n43639), .B(n43650), .Z(n43626) );
  XOR U52931 ( .A(n43640), .B(n43641), .Z(n43650) );
  XOR U52932 ( .A(n43646), .B(n43651), .Z(n43641) );
  XOR U52933 ( .A(n43645), .B(n43648), .Z(n43651) );
  IV U52934 ( .A(n43647), .Z(n43648) );
  NAND U52935 ( .A(n43652), .B(n43653), .Z(n43647) );
  OR U52936 ( .A(n43654), .B(n43655), .Z(n43653) );
  OR U52937 ( .A(n43656), .B(n43657), .Z(n43652) );
  NAND U52938 ( .A(n43658), .B(n43659), .Z(n43645) );
  OR U52939 ( .A(n43660), .B(n43661), .Z(n43659) );
  OR U52940 ( .A(n43662), .B(n43663), .Z(n43658) );
  NOR U52941 ( .A(n43664), .B(n43665), .Z(n43646) );
  ANDN U52942 ( .B(n43666), .A(n43667), .Z(n43640) );
  XNOR U52943 ( .A(n43633), .B(n43668), .Z(n43639) );
  XNOR U52944 ( .A(n43632), .B(n43634), .Z(n43668) );
  NAND U52945 ( .A(n43669), .B(n43670), .Z(n43634) );
  OR U52946 ( .A(n43671), .B(n43672), .Z(n43670) );
  OR U52947 ( .A(n43673), .B(n43674), .Z(n43669) );
  NAND U52948 ( .A(n43675), .B(n43676), .Z(n43632) );
  OR U52949 ( .A(n43677), .B(n43678), .Z(n43676) );
  OR U52950 ( .A(n43679), .B(n43680), .Z(n43675) );
  ANDN U52951 ( .B(n43681), .A(n43682), .Z(n43633) );
  IV U52952 ( .A(n43683), .Z(n43681) );
  ANDN U52953 ( .B(n43684), .A(n43685), .Z(n43625) );
  XOR U52954 ( .A(n43611), .B(n43686), .Z(n43623) );
  XOR U52955 ( .A(n43612), .B(n43613), .Z(n43686) );
  XOR U52956 ( .A(n43618), .B(n43687), .Z(n43613) );
  XOR U52957 ( .A(n43617), .B(n43620), .Z(n43687) );
  IV U52958 ( .A(n43619), .Z(n43620) );
  NAND U52959 ( .A(n43688), .B(n43689), .Z(n43619) );
  OR U52960 ( .A(n43690), .B(n43691), .Z(n43689) );
  OR U52961 ( .A(n43692), .B(n43693), .Z(n43688) );
  NAND U52962 ( .A(n43694), .B(n43695), .Z(n43617) );
  OR U52963 ( .A(n43696), .B(n43697), .Z(n43695) );
  OR U52964 ( .A(n43698), .B(n43699), .Z(n43694) );
  NOR U52965 ( .A(n43700), .B(n43701), .Z(n43618) );
  ANDN U52966 ( .B(n43702), .A(n43703), .Z(n43612) );
  IV U52967 ( .A(n43704), .Z(n43702) );
  XNOR U52968 ( .A(n43605), .B(n43705), .Z(n43611) );
  XNOR U52969 ( .A(n43604), .B(n43606), .Z(n43705) );
  NAND U52970 ( .A(n43706), .B(n43707), .Z(n43606) );
  OR U52971 ( .A(n43708), .B(n43709), .Z(n43707) );
  OR U52972 ( .A(n43710), .B(n43711), .Z(n43706) );
  NAND U52973 ( .A(n43712), .B(n43713), .Z(n43604) );
  OR U52974 ( .A(n43714), .B(n43715), .Z(n43713) );
  OR U52975 ( .A(n43716), .B(n43717), .Z(n43712) );
  ANDN U52976 ( .B(n43718), .A(n43719), .Z(n43605) );
  IV U52977 ( .A(n43720), .Z(n43718) );
  XNOR U52978 ( .A(n43685), .B(n43684), .Z(N61528) );
  XOR U52979 ( .A(n43704), .B(n43703), .Z(n43684) );
  XNOR U52980 ( .A(n43719), .B(n43720), .Z(n43703) );
  XNOR U52981 ( .A(n43714), .B(n43715), .Z(n43720) );
  XNOR U52982 ( .A(n43716), .B(n43717), .Z(n43715) );
  XNOR U52983 ( .A(y[1741]), .B(x[1741]), .Z(n43717) );
  XNOR U52984 ( .A(y[1742]), .B(x[1742]), .Z(n43716) );
  XNOR U52985 ( .A(y[1740]), .B(x[1740]), .Z(n43714) );
  XNOR U52986 ( .A(n43708), .B(n43709), .Z(n43719) );
  XNOR U52987 ( .A(y[1737]), .B(x[1737]), .Z(n43709) );
  XNOR U52988 ( .A(n43710), .B(n43711), .Z(n43708) );
  XNOR U52989 ( .A(y[1738]), .B(x[1738]), .Z(n43711) );
  XNOR U52990 ( .A(y[1739]), .B(x[1739]), .Z(n43710) );
  XNOR U52991 ( .A(n43701), .B(n43700), .Z(n43704) );
  XNOR U52992 ( .A(n43696), .B(n43697), .Z(n43700) );
  XNOR U52993 ( .A(y[1734]), .B(x[1734]), .Z(n43697) );
  XNOR U52994 ( .A(n43698), .B(n43699), .Z(n43696) );
  XNOR U52995 ( .A(y[1735]), .B(x[1735]), .Z(n43699) );
  XNOR U52996 ( .A(y[1736]), .B(x[1736]), .Z(n43698) );
  XNOR U52997 ( .A(n43690), .B(n43691), .Z(n43701) );
  XNOR U52998 ( .A(y[1731]), .B(x[1731]), .Z(n43691) );
  XNOR U52999 ( .A(n43692), .B(n43693), .Z(n43690) );
  XNOR U53000 ( .A(y[1732]), .B(x[1732]), .Z(n43693) );
  XNOR U53001 ( .A(y[1733]), .B(x[1733]), .Z(n43692) );
  XOR U53002 ( .A(n43666), .B(n43667), .Z(n43685) );
  XNOR U53003 ( .A(n43682), .B(n43683), .Z(n43667) );
  XNOR U53004 ( .A(n43677), .B(n43678), .Z(n43683) );
  XNOR U53005 ( .A(n43679), .B(n43680), .Z(n43678) );
  XNOR U53006 ( .A(y[1729]), .B(x[1729]), .Z(n43680) );
  XNOR U53007 ( .A(y[1730]), .B(x[1730]), .Z(n43679) );
  XNOR U53008 ( .A(y[1728]), .B(x[1728]), .Z(n43677) );
  XNOR U53009 ( .A(n43671), .B(n43672), .Z(n43682) );
  XNOR U53010 ( .A(y[1725]), .B(x[1725]), .Z(n43672) );
  XNOR U53011 ( .A(n43673), .B(n43674), .Z(n43671) );
  XNOR U53012 ( .A(y[1726]), .B(x[1726]), .Z(n43674) );
  XNOR U53013 ( .A(y[1727]), .B(x[1727]), .Z(n43673) );
  XOR U53014 ( .A(n43665), .B(n43664), .Z(n43666) );
  XNOR U53015 ( .A(n43660), .B(n43661), .Z(n43664) );
  XNOR U53016 ( .A(y[1722]), .B(x[1722]), .Z(n43661) );
  XNOR U53017 ( .A(n43662), .B(n43663), .Z(n43660) );
  XNOR U53018 ( .A(y[1723]), .B(x[1723]), .Z(n43663) );
  XNOR U53019 ( .A(y[1724]), .B(x[1724]), .Z(n43662) );
  XNOR U53020 ( .A(n43654), .B(n43655), .Z(n43665) );
  XNOR U53021 ( .A(y[1719]), .B(x[1719]), .Z(n43655) );
  XNOR U53022 ( .A(n43656), .B(n43657), .Z(n43654) );
  XNOR U53023 ( .A(y[1720]), .B(x[1720]), .Z(n43657) );
  XNOR U53024 ( .A(y[1721]), .B(x[1721]), .Z(n43656) );
  NAND U53025 ( .A(n43721), .B(n43722), .Z(N61519) );
  NANDN U53026 ( .A(n43723), .B(n43724), .Z(n43722) );
  OR U53027 ( .A(n43725), .B(n43726), .Z(n43724) );
  NAND U53028 ( .A(n43725), .B(n43726), .Z(n43721) );
  XOR U53029 ( .A(n43725), .B(n43727), .Z(N61518) );
  XNOR U53030 ( .A(n43723), .B(n43726), .Z(n43727) );
  AND U53031 ( .A(n43728), .B(n43729), .Z(n43726) );
  NANDN U53032 ( .A(n43730), .B(n43731), .Z(n43729) );
  NANDN U53033 ( .A(n43732), .B(n43733), .Z(n43731) );
  NANDN U53034 ( .A(n43733), .B(n43732), .Z(n43728) );
  NAND U53035 ( .A(n43734), .B(n43735), .Z(n43723) );
  NANDN U53036 ( .A(n43736), .B(n43737), .Z(n43735) );
  OR U53037 ( .A(n43738), .B(n43739), .Z(n43737) );
  NAND U53038 ( .A(n43739), .B(n43738), .Z(n43734) );
  AND U53039 ( .A(n43740), .B(n43741), .Z(n43725) );
  NANDN U53040 ( .A(n43742), .B(n43743), .Z(n43741) );
  NANDN U53041 ( .A(n43744), .B(n43745), .Z(n43743) );
  NANDN U53042 ( .A(n43745), .B(n43744), .Z(n43740) );
  XOR U53043 ( .A(n43739), .B(n43746), .Z(N61517) );
  XOR U53044 ( .A(n43736), .B(n43738), .Z(n43746) );
  XNOR U53045 ( .A(n43732), .B(n43747), .Z(n43738) );
  XNOR U53046 ( .A(n43730), .B(n43733), .Z(n43747) );
  NAND U53047 ( .A(n43748), .B(n43749), .Z(n43733) );
  NAND U53048 ( .A(n43750), .B(n43751), .Z(n43749) );
  OR U53049 ( .A(n43752), .B(n43753), .Z(n43750) );
  NANDN U53050 ( .A(n43754), .B(n43752), .Z(n43748) );
  IV U53051 ( .A(n43753), .Z(n43754) );
  NAND U53052 ( .A(n43755), .B(n43756), .Z(n43730) );
  NAND U53053 ( .A(n43757), .B(n43758), .Z(n43756) );
  NANDN U53054 ( .A(n43759), .B(n43760), .Z(n43757) );
  NANDN U53055 ( .A(n43760), .B(n43759), .Z(n43755) );
  AND U53056 ( .A(n43761), .B(n43762), .Z(n43732) );
  NAND U53057 ( .A(n43763), .B(n43764), .Z(n43762) );
  OR U53058 ( .A(n43765), .B(n43766), .Z(n43763) );
  NANDN U53059 ( .A(n43767), .B(n43765), .Z(n43761) );
  NAND U53060 ( .A(n43768), .B(n43769), .Z(n43736) );
  NANDN U53061 ( .A(n43770), .B(n43771), .Z(n43769) );
  OR U53062 ( .A(n43772), .B(n43773), .Z(n43771) );
  NANDN U53063 ( .A(n43774), .B(n43772), .Z(n43768) );
  IV U53064 ( .A(n43773), .Z(n43774) );
  XNOR U53065 ( .A(n43744), .B(n43775), .Z(n43739) );
  XNOR U53066 ( .A(n43742), .B(n43745), .Z(n43775) );
  NAND U53067 ( .A(n43776), .B(n43777), .Z(n43745) );
  NAND U53068 ( .A(n43778), .B(n43779), .Z(n43777) );
  OR U53069 ( .A(n43780), .B(n43781), .Z(n43778) );
  NANDN U53070 ( .A(n43782), .B(n43780), .Z(n43776) );
  IV U53071 ( .A(n43781), .Z(n43782) );
  NAND U53072 ( .A(n43783), .B(n43784), .Z(n43742) );
  NAND U53073 ( .A(n43785), .B(n43786), .Z(n43784) );
  NANDN U53074 ( .A(n43787), .B(n43788), .Z(n43785) );
  NANDN U53075 ( .A(n43788), .B(n43787), .Z(n43783) );
  AND U53076 ( .A(n43789), .B(n43790), .Z(n43744) );
  NAND U53077 ( .A(n43791), .B(n43792), .Z(n43790) );
  OR U53078 ( .A(n43793), .B(n43794), .Z(n43791) );
  NANDN U53079 ( .A(n43795), .B(n43793), .Z(n43789) );
  XNOR U53080 ( .A(n43770), .B(n43796), .Z(N61516) );
  XOR U53081 ( .A(n43772), .B(n43773), .Z(n43796) );
  XNOR U53082 ( .A(n43786), .B(n43797), .Z(n43773) );
  XOR U53083 ( .A(n43787), .B(n43788), .Z(n43797) );
  XOR U53084 ( .A(n43793), .B(n43798), .Z(n43788) );
  XOR U53085 ( .A(n43792), .B(n43795), .Z(n43798) );
  IV U53086 ( .A(n43794), .Z(n43795) );
  NAND U53087 ( .A(n43799), .B(n43800), .Z(n43794) );
  OR U53088 ( .A(n43801), .B(n43802), .Z(n43800) );
  OR U53089 ( .A(n43803), .B(n43804), .Z(n43799) );
  NAND U53090 ( .A(n43805), .B(n43806), .Z(n43792) );
  OR U53091 ( .A(n43807), .B(n43808), .Z(n43806) );
  OR U53092 ( .A(n43809), .B(n43810), .Z(n43805) );
  NOR U53093 ( .A(n43811), .B(n43812), .Z(n43793) );
  ANDN U53094 ( .B(n43813), .A(n43814), .Z(n43787) );
  XNOR U53095 ( .A(n43780), .B(n43815), .Z(n43786) );
  XNOR U53096 ( .A(n43779), .B(n43781), .Z(n43815) );
  NAND U53097 ( .A(n43816), .B(n43817), .Z(n43781) );
  OR U53098 ( .A(n43818), .B(n43819), .Z(n43817) );
  OR U53099 ( .A(n43820), .B(n43821), .Z(n43816) );
  NAND U53100 ( .A(n43822), .B(n43823), .Z(n43779) );
  OR U53101 ( .A(n43824), .B(n43825), .Z(n43823) );
  OR U53102 ( .A(n43826), .B(n43827), .Z(n43822) );
  ANDN U53103 ( .B(n43828), .A(n43829), .Z(n43780) );
  IV U53104 ( .A(n43830), .Z(n43828) );
  ANDN U53105 ( .B(n43831), .A(n43832), .Z(n43772) );
  XOR U53106 ( .A(n43758), .B(n43833), .Z(n43770) );
  XOR U53107 ( .A(n43759), .B(n43760), .Z(n43833) );
  XOR U53108 ( .A(n43765), .B(n43834), .Z(n43760) );
  XOR U53109 ( .A(n43764), .B(n43767), .Z(n43834) );
  IV U53110 ( .A(n43766), .Z(n43767) );
  NAND U53111 ( .A(n43835), .B(n43836), .Z(n43766) );
  OR U53112 ( .A(n43837), .B(n43838), .Z(n43836) );
  OR U53113 ( .A(n43839), .B(n43840), .Z(n43835) );
  NAND U53114 ( .A(n43841), .B(n43842), .Z(n43764) );
  OR U53115 ( .A(n43843), .B(n43844), .Z(n43842) );
  OR U53116 ( .A(n43845), .B(n43846), .Z(n43841) );
  NOR U53117 ( .A(n43847), .B(n43848), .Z(n43765) );
  ANDN U53118 ( .B(n43849), .A(n43850), .Z(n43759) );
  IV U53119 ( .A(n43851), .Z(n43849) );
  XNOR U53120 ( .A(n43752), .B(n43852), .Z(n43758) );
  XNOR U53121 ( .A(n43751), .B(n43753), .Z(n43852) );
  NAND U53122 ( .A(n43853), .B(n43854), .Z(n43753) );
  OR U53123 ( .A(n43855), .B(n43856), .Z(n43854) );
  OR U53124 ( .A(n43857), .B(n43858), .Z(n43853) );
  NAND U53125 ( .A(n43859), .B(n43860), .Z(n43751) );
  OR U53126 ( .A(n43861), .B(n43862), .Z(n43860) );
  OR U53127 ( .A(n43863), .B(n43864), .Z(n43859) );
  ANDN U53128 ( .B(n43865), .A(n43866), .Z(n43752) );
  IV U53129 ( .A(n43867), .Z(n43865) );
  XNOR U53130 ( .A(n43832), .B(n43831), .Z(N61515) );
  XOR U53131 ( .A(n43851), .B(n43850), .Z(n43831) );
  XNOR U53132 ( .A(n43866), .B(n43867), .Z(n43850) );
  XNOR U53133 ( .A(n43861), .B(n43862), .Z(n43867) );
  XNOR U53134 ( .A(n43863), .B(n43864), .Z(n43862) );
  XNOR U53135 ( .A(y[1717]), .B(x[1717]), .Z(n43864) );
  XNOR U53136 ( .A(y[1718]), .B(x[1718]), .Z(n43863) );
  XNOR U53137 ( .A(y[1716]), .B(x[1716]), .Z(n43861) );
  XNOR U53138 ( .A(n43855), .B(n43856), .Z(n43866) );
  XNOR U53139 ( .A(y[1713]), .B(x[1713]), .Z(n43856) );
  XNOR U53140 ( .A(n43857), .B(n43858), .Z(n43855) );
  XNOR U53141 ( .A(y[1714]), .B(x[1714]), .Z(n43858) );
  XNOR U53142 ( .A(y[1715]), .B(x[1715]), .Z(n43857) );
  XNOR U53143 ( .A(n43848), .B(n43847), .Z(n43851) );
  XNOR U53144 ( .A(n43843), .B(n43844), .Z(n43847) );
  XNOR U53145 ( .A(y[1710]), .B(x[1710]), .Z(n43844) );
  XNOR U53146 ( .A(n43845), .B(n43846), .Z(n43843) );
  XNOR U53147 ( .A(y[1711]), .B(x[1711]), .Z(n43846) );
  XNOR U53148 ( .A(y[1712]), .B(x[1712]), .Z(n43845) );
  XNOR U53149 ( .A(n43837), .B(n43838), .Z(n43848) );
  XNOR U53150 ( .A(y[1707]), .B(x[1707]), .Z(n43838) );
  XNOR U53151 ( .A(n43839), .B(n43840), .Z(n43837) );
  XNOR U53152 ( .A(y[1708]), .B(x[1708]), .Z(n43840) );
  XNOR U53153 ( .A(y[1709]), .B(x[1709]), .Z(n43839) );
  XOR U53154 ( .A(n43813), .B(n43814), .Z(n43832) );
  XNOR U53155 ( .A(n43829), .B(n43830), .Z(n43814) );
  XNOR U53156 ( .A(n43824), .B(n43825), .Z(n43830) );
  XNOR U53157 ( .A(n43826), .B(n43827), .Z(n43825) );
  XNOR U53158 ( .A(y[1705]), .B(x[1705]), .Z(n43827) );
  XNOR U53159 ( .A(y[1706]), .B(x[1706]), .Z(n43826) );
  XNOR U53160 ( .A(y[1704]), .B(x[1704]), .Z(n43824) );
  XNOR U53161 ( .A(n43818), .B(n43819), .Z(n43829) );
  XNOR U53162 ( .A(y[1701]), .B(x[1701]), .Z(n43819) );
  XNOR U53163 ( .A(n43820), .B(n43821), .Z(n43818) );
  XNOR U53164 ( .A(y[1702]), .B(x[1702]), .Z(n43821) );
  XNOR U53165 ( .A(y[1703]), .B(x[1703]), .Z(n43820) );
  XOR U53166 ( .A(n43812), .B(n43811), .Z(n43813) );
  XNOR U53167 ( .A(n43807), .B(n43808), .Z(n43811) );
  XNOR U53168 ( .A(y[1698]), .B(x[1698]), .Z(n43808) );
  XNOR U53169 ( .A(n43809), .B(n43810), .Z(n43807) );
  XNOR U53170 ( .A(y[1699]), .B(x[1699]), .Z(n43810) );
  XNOR U53171 ( .A(y[1700]), .B(x[1700]), .Z(n43809) );
  XNOR U53172 ( .A(n43801), .B(n43802), .Z(n43812) );
  XNOR U53173 ( .A(y[1695]), .B(x[1695]), .Z(n43802) );
  XNOR U53174 ( .A(n43803), .B(n43804), .Z(n43801) );
  XNOR U53175 ( .A(y[1696]), .B(x[1696]), .Z(n43804) );
  XNOR U53176 ( .A(y[1697]), .B(x[1697]), .Z(n43803) );
  NAND U53177 ( .A(n43868), .B(n43869), .Z(N61506) );
  NANDN U53178 ( .A(n43870), .B(n43871), .Z(n43869) );
  OR U53179 ( .A(n43872), .B(n43873), .Z(n43871) );
  NAND U53180 ( .A(n43872), .B(n43873), .Z(n43868) );
  XOR U53181 ( .A(n43872), .B(n43874), .Z(N61505) );
  XNOR U53182 ( .A(n43870), .B(n43873), .Z(n43874) );
  AND U53183 ( .A(n43875), .B(n43876), .Z(n43873) );
  NANDN U53184 ( .A(n43877), .B(n43878), .Z(n43876) );
  NANDN U53185 ( .A(n43879), .B(n43880), .Z(n43878) );
  NANDN U53186 ( .A(n43880), .B(n43879), .Z(n43875) );
  NAND U53187 ( .A(n43881), .B(n43882), .Z(n43870) );
  NANDN U53188 ( .A(n43883), .B(n43884), .Z(n43882) );
  OR U53189 ( .A(n43885), .B(n43886), .Z(n43884) );
  NAND U53190 ( .A(n43886), .B(n43885), .Z(n43881) );
  AND U53191 ( .A(n43887), .B(n43888), .Z(n43872) );
  NANDN U53192 ( .A(n43889), .B(n43890), .Z(n43888) );
  NANDN U53193 ( .A(n43891), .B(n43892), .Z(n43890) );
  NANDN U53194 ( .A(n43892), .B(n43891), .Z(n43887) );
  XOR U53195 ( .A(n43886), .B(n43893), .Z(N61504) );
  XOR U53196 ( .A(n43883), .B(n43885), .Z(n43893) );
  XNOR U53197 ( .A(n43879), .B(n43894), .Z(n43885) );
  XNOR U53198 ( .A(n43877), .B(n43880), .Z(n43894) );
  NAND U53199 ( .A(n43895), .B(n43896), .Z(n43880) );
  NAND U53200 ( .A(n43897), .B(n43898), .Z(n43896) );
  OR U53201 ( .A(n43899), .B(n43900), .Z(n43897) );
  NANDN U53202 ( .A(n43901), .B(n43899), .Z(n43895) );
  IV U53203 ( .A(n43900), .Z(n43901) );
  NAND U53204 ( .A(n43902), .B(n43903), .Z(n43877) );
  NAND U53205 ( .A(n43904), .B(n43905), .Z(n43903) );
  NANDN U53206 ( .A(n43906), .B(n43907), .Z(n43904) );
  NANDN U53207 ( .A(n43907), .B(n43906), .Z(n43902) );
  AND U53208 ( .A(n43908), .B(n43909), .Z(n43879) );
  NAND U53209 ( .A(n43910), .B(n43911), .Z(n43909) );
  OR U53210 ( .A(n43912), .B(n43913), .Z(n43910) );
  NANDN U53211 ( .A(n43914), .B(n43912), .Z(n43908) );
  NAND U53212 ( .A(n43915), .B(n43916), .Z(n43883) );
  NANDN U53213 ( .A(n43917), .B(n43918), .Z(n43916) );
  OR U53214 ( .A(n43919), .B(n43920), .Z(n43918) );
  NANDN U53215 ( .A(n43921), .B(n43919), .Z(n43915) );
  IV U53216 ( .A(n43920), .Z(n43921) );
  XNOR U53217 ( .A(n43891), .B(n43922), .Z(n43886) );
  XNOR U53218 ( .A(n43889), .B(n43892), .Z(n43922) );
  NAND U53219 ( .A(n43923), .B(n43924), .Z(n43892) );
  NAND U53220 ( .A(n43925), .B(n43926), .Z(n43924) );
  OR U53221 ( .A(n43927), .B(n43928), .Z(n43925) );
  NANDN U53222 ( .A(n43929), .B(n43927), .Z(n43923) );
  IV U53223 ( .A(n43928), .Z(n43929) );
  NAND U53224 ( .A(n43930), .B(n43931), .Z(n43889) );
  NAND U53225 ( .A(n43932), .B(n43933), .Z(n43931) );
  NANDN U53226 ( .A(n43934), .B(n43935), .Z(n43932) );
  NANDN U53227 ( .A(n43935), .B(n43934), .Z(n43930) );
  AND U53228 ( .A(n43936), .B(n43937), .Z(n43891) );
  NAND U53229 ( .A(n43938), .B(n43939), .Z(n43937) );
  OR U53230 ( .A(n43940), .B(n43941), .Z(n43938) );
  NANDN U53231 ( .A(n43942), .B(n43940), .Z(n43936) );
  XNOR U53232 ( .A(n43917), .B(n43943), .Z(N61503) );
  XOR U53233 ( .A(n43919), .B(n43920), .Z(n43943) );
  XNOR U53234 ( .A(n43933), .B(n43944), .Z(n43920) );
  XOR U53235 ( .A(n43934), .B(n43935), .Z(n43944) );
  XOR U53236 ( .A(n43940), .B(n43945), .Z(n43935) );
  XOR U53237 ( .A(n43939), .B(n43942), .Z(n43945) );
  IV U53238 ( .A(n43941), .Z(n43942) );
  NAND U53239 ( .A(n43946), .B(n43947), .Z(n43941) );
  OR U53240 ( .A(n43948), .B(n43949), .Z(n43947) );
  OR U53241 ( .A(n43950), .B(n43951), .Z(n43946) );
  NAND U53242 ( .A(n43952), .B(n43953), .Z(n43939) );
  OR U53243 ( .A(n43954), .B(n43955), .Z(n43953) );
  OR U53244 ( .A(n43956), .B(n43957), .Z(n43952) );
  NOR U53245 ( .A(n43958), .B(n43959), .Z(n43940) );
  ANDN U53246 ( .B(n43960), .A(n43961), .Z(n43934) );
  XNOR U53247 ( .A(n43927), .B(n43962), .Z(n43933) );
  XNOR U53248 ( .A(n43926), .B(n43928), .Z(n43962) );
  NAND U53249 ( .A(n43963), .B(n43964), .Z(n43928) );
  OR U53250 ( .A(n43965), .B(n43966), .Z(n43964) );
  OR U53251 ( .A(n43967), .B(n43968), .Z(n43963) );
  NAND U53252 ( .A(n43969), .B(n43970), .Z(n43926) );
  OR U53253 ( .A(n43971), .B(n43972), .Z(n43970) );
  OR U53254 ( .A(n43973), .B(n43974), .Z(n43969) );
  ANDN U53255 ( .B(n43975), .A(n43976), .Z(n43927) );
  IV U53256 ( .A(n43977), .Z(n43975) );
  ANDN U53257 ( .B(n43978), .A(n43979), .Z(n43919) );
  XOR U53258 ( .A(n43905), .B(n43980), .Z(n43917) );
  XOR U53259 ( .A(n43906), .B(n43907), .Z(n43980) );
  XOR U53260 ( .A(n43912), .B(n43981), .Z(n43907) );
  XOR U53261 ( .A(n43911), .B(n43914), .Z(n43981) );
  IV U53262 ( .A(n43913), .Z(n43914) );
  NAND U53263 ( .A(n43982), .B(n43983), .Z(n43913) );
  OR U53264 ( .A(n43984), .B(n43985), .Z(n43983) );
  OR U53265 ( .A(n43986), .B(n43987), .Z(n43982) );
  NAND U53266 ( .A(n43988), .B(n43989), .Z(n43911) );
  OR U53267 ( .A(n43990), .B(n43991), .Z(n43989) );
  OR U53268 ( .A(n43992), .B(n43993), .Z(n43988) );
  NOR U53269 ( .A(n43994), .B(n43995), .Z(n43912) );
  ANDN U53270 ( .B(n43996), .A(n43997), .Z(n43906) );
  IV U53271 ( .A(n43998), .Z(n43996) );
  XNOR U53272 ( .A(n43899), .B(n43999), .Z(n43905) );
  XNOR U53273 ( .A(n43898), .B(n43900), .Z(n43999) );
  NAND U53274 ( .A(n44000), .B(n44001), .Z(n43900) );
  OR U53275 ( .A(n44002), .B(n44003), .Z(n44001) );
  OR U53276 ( .A(n44004), .B(n44005), .Z(n44000) );
  NAND U53277 ( .A(n44006), .B(n44007), .Z(n43898) );
  OR U53278 ( .A(n44008), .B(n44009), .Z(n44007) );
  OR U53279 ( .A(n44010), .B(n44011), .Z(n44006) );
  ANDN U53280 ( .B(n44012), .A(n44013), .Z(n43899) );
  IV U53281 ( .A(n44014), .Z(n44012) );
  XNOR U53282 ( .A(n43979), .B(n43978), .Z(N61502) );
  XOR U53283 ( .A(n43998), .B(n43997), .Z(n43978) );
  XNOR U53284 ( .A(n44013), .B(n44014), .Z(n43997) );
  XNOR U53285 ( .A(n44008), .B(n44009), .Z(n44014) );
  XNOR U53286 ( .A(n44010), .B(n44011), .Z(n44009) );
  XNOR U53287 ( .A(y[1693]), .B(x[1693]), .Z(n44011) );
  XNOR U53288 ( .A(y[1694]), .B(x[1694]), .Z(n44010) );
  XNOR U53289 ( .A(y[1692]), .B(x[1692]), .Z(n44008) );
  XNOR U53290 ( .A(n44002), .B(n44003), .Z(n44013) );
  XNOR U53291 ( .A(y[1689]), .B(x[1689]), .Z(n44003) );
  XNOR U53292 ( .A(n44004), .B(n44005), .Z(n44002) );
  XNOR U53293 ( .A(y[1690]), .B(x[1690]), .Z(n44005) );
  XNOR U53294 ( .A(y[1691]), .B(x[1691]), .Z(n44004) );
  XNOR U53295 ( .A(n43995), .B(n43994), .Z(n43998) );
  XNOR U53296 ( .A(n43990), .B(n43991), .Z(n43994) );
  XNOR U53297 ( .A(y[1686]), .B(x[1686]), .Z(n43991) );
  XNOR U53298 ( .A(n43992), .B(n43993), .Z(n43990) );
  XNOR U53299 ( .A(y[1687]), .B(x[1687]), .Z(n43993) );
  XNOR U53300 ( .A(y[1688]), .B(x[1688]), .Z(n43992) );
  XNOR U53301 ( .A(n43984), .B(n43985), .Z(n43995) );
  XNOR U53302 ( .A(y[1683]), .B(x[1683]), .Z(n43985) );
  XNOR U53303 ( .A(n43986), .B(n43987), .Z(n43984) );
  XNOR U53304 ( .A(y[1684]), .B(x[1684]), .Z(n43987) );
  XNOR U53305 ( .A(y[1685]), .B(x[1685]), .Z(n43986) );
  XOR U53306 ( .A(n43960), .B(n43961), .Z(n43979) );
  XNOR U53307 ( .A(n43976), .B(n43977), .Z(n43961) );
  XNOR U53308 ( .A(n43971), .B(n43972), .Z(n43977) );
  XNOR U53309 ( .A(n43973), .B(n43974), .Z(n43972) );
  XNOR U53310 ( .A(y[1681]), .B(x[1681]), .Z(n43974) );
  XNOR U53311 ( .A(y[1682]), .B(x[1682]), .Z(n43973) );
  XNOR U53312 ( .A(y[1680]), .B(x[1680]), .Z(n43971) );
  XNOR U53313 ( .A(n43965), .B(n43966), .Z(n43976) );
  XNOR U53314 ( .A(y[1677]), .B(x[1677]), .Z(n43966) );
  XNOR U53315 ( .A(n43967), .B(n43968), .Z(n43965) );
  XNOR U53316 ( .A(y[1678]), .B(x[1678]), .Z(n43968) );
  XNOR U53317 ( .A(y[1679]), .B(x[1679]), .Z(n43967) );
  XOR U53318 ( .A(n43959), .B(n43958), .Z(n43960) );
  XNOR U53319 ( .A(n43954), .B(n43955), .Z(n43958) );
  XNOR U53320 ( .A(y[1674]), .B(x[1674]), .Z(n43955) );
  XNOR U53321 ( .A(n43956), .B(n43957), .Z(n43954) );
  XNOR U53322 ( .A(y[1675]), .B(x[1675]), .Z(n43957) );
  XNOR U53323 ( .A(y[1676]), .B(x[1676]), .Z(n43956) );
  XNOR U53324 ( .A(n43948), .B(n43949), .Z(n43959) );
  XNOR U53325 ( .A(y[1671]), .B(x[1671]), .Z(n43949) );
  XNOR U53326 ( .A(n43950), .B(n43951), .Z(n43948) );
  XNOR U53327 ( .A(y[1672]), .B(x[1672]), .Z(n43951) );
  XNOR U53328 ( .A(y[1673]), .B(x[1673]), .Z(n43950) );
  NAND U53329 ( .A(n44015), .B(n44016), .Z(N61493) );
  NANDN U53330 ( .A(n44017), .B(n44018), .Z(n44016) );
  OR U53331 ( .A(n44019), .B(n44020), .Z(n44018) );
  NAND U53332 ( .A(n44019), .B(n44020), .Z(n44015) );
  XOR U53333 ( .A(n44019), .B(n44021), .Z(N61492) );
  XNOR U53334 ( .A(n44017), .B(n44020), .Z(n44021) );
  AND U53335 ( .A(n44022), .B(n44023), .Z(n44020) );
  NANDN U53336 ( .A(n44024), .B(n44025), .Z(n44023) );
  NANDN U53337 ( .A(n44026), .B(n44027), .Z(n44025) );
  NANDN U53338 ( .A(n44027), .B(n44026), .Z(n44022) );
  NAND U53339 ( .A(n44028), .B(n44029), .Z(n44017) );
  NANDN U53340 ( .A(n44030), .B(n44031), .Z(n44029) );
  OR U53341 ( .A(n44032), .B(n44033), .Z(n44031) );
  NAND U53342 ( .A(n44033), .B(n44032), .Z(n44028) );
  AND U53343 ( .A(n44034), .B(n44035), .Z(n44019) );
  NANDN U53344 ( .A(n44036), .B(n44037), .Z(n44035) );
  NANDN U53345 ( .A(n44038), .B(n44039), .Z(n44037) );
  NANDN U53346 ( .A(n44039), .B(n44038), .Z(n44034) );
  XOR U53347 ( .A(n44033), .B(n44040), .Z(N61491) );
  XOR U53348 ( .A(n44030), .B(n44032), .Z(n44040) );
  XNOR U53349 ( .A(n44026), .B(n44041), .Z(n44032) );
  XNOR U53350 ( .A(n44024), .B(n44027), .Z(n44041) );
  NAND U53351 ( .A(n44042), .B(n44043), .Z(n44027) );
  NAND U53352 ( .A(n44044), .B(n44045), .Z(n44043) );
  OR U53353 ( .A(n44046), .B(n44047), .Z(n44044) );
  NANDN U53354 ( .A(n44048), .B(n44046), .Z(n44042) );
  IV U53355 ( .A(n44047), .Z(n44048) );
  NAND U53356 ( .A(n44049), .B(n44050), .Z(n44024) );
  NAND U53357 ( .A(n44051), .B(n44052), .Z(n44050) );
  NANDN U53358 ( .A(n44053), .B(n44054), .Z(n44051) );
  NANDN U53359 ( .A(n44054), .B(n44053), .Z(n44049) );
  AND U53360 ( .A(n44055), .B(n44056), .Z(n44026) );
  NAND U53361 ( .A(n44057), .B(n44058), .Z(n44056) );
  OR U53362 ( .A(n44059), .B(n44060), .Z(n44057) );
  NANDN U53363 ( .A(n44061), .B(n44059), .Z(n44055) );
  NAND U53364 ( .A(n44062), .B(n44063), .Z(n44030) );
  NANDN U53365 ( .A(n44064), .B(n44065), .Z(n44063) );
  OR U53366 ( .A(n44066), .B(n44067), .Z(n44065) );
  NANDN U53367 ( .A(n44068), .B(n44066), .Z(n44062) );
  IV U53368 ( .A(n44067), .Z(n44068) );
  XNOR U53369 ( .A(n44038), .B(n44069), .Z(n44033) );
  XNOR U53370 ( .A(n44036), .B(n44039), .Z(n44069) );
  NAND U53371 ( .A(n44070), .B(n44071), .Z(n44039) );
  NAND U53372 ( .A(n44072), .B(n44073), .Z(n44071) );
  OR U53373 ( .A(n44074), .B(n44075), .Z(n44072) );
  NANDN U53374 ( .A(n44076), .B(n44074), .Z(n44070) );
  IV U53375 ( .A(n44075), .Z(n44076) );
  NAND U53376 ( .A(n44077), .B(n44078), .Z(n44036) );
  NAND U53377 ( .A(n44079), .B(n44080), .Z(n44078) );
  NANDN U53378 ( .A(n44081), .B(n44082), .Z(n44079) );
  NANDN U53379 ( .A(n44082), .B(n44081), .Z(n44077) );
  AND U53380 ( .A(n44083), .B(n44084), .Z(n44038) );
  NAND U53381 ( .A(n44085), .B(n44086), .Z(n44084) );
  OR U53382 ( .A(n44087), .B(n44088), .Z(n44085) );
  NANDN U53383 ( .A(n44089), .B(n44087), .Z(n44083) );
  XNOR U53384 ( .A(n44064), .B(n44090), .Z(N61490) );
  XOR U53385 ( .A(n44066), .B(n44067), .Z(n44090) );
  XNOR U53386 ( .A(n44080), .B(n44091), .Z(n44067) );
  XOR U53387 ( .A(n44081), .B(n44082), .Z(n44091) );
  XOR U53388 ( .A(n44087), .B(n44092), .Z(n44082) );
  XOR U53389 ( .A(n44086), .B(n44089), .Z(n44092) );
  IV U53390 ( .A(n44088), .Z(n44089) );
  NAND U53391 ( .A(n44093), .B(n44094), .Z(n44088) );
  OR U53392 ( .A(n44095), .B(n44096), .Z(n44094) );
  OR U53393 ( .A(n44097), .B(n44098), .Z(n44093) );
  NAND U53394 ( .A(n44099), .B(n44100), .Z(n44086) );
  OR U53395 ( .A(n44101), .B(n44102), .Z(n44100) );
  OR U53396 ( .A(n44103), .B(n44104), .Z(n44099) );
  NOR U53397 ( .A(n44105), .B(n44106), .Z(n44087) );
  ANDN U53398 ( .B(n44107), .A(n44108), .Z(n44081) );
  XNOR U53399 ( .A(n44074), .B(n44109), .Z(n44080) );
  XNOR U53400 ( .A(n44073), .B(n44075), .Z(n44109) );
  NAND U53401 ( .A(n44110), .B(n44111), .Z(n44075) );
  OR U53402 ( .A(n44112), .B(n44113), .Z(n44111) );
  OR U53403 ( .A(n44114), .B(n44115), .Z(n44110) );
  NAND U53404 ( .A(n44116), .B(n44117), .Z(n44073) );
  OR U53405 ( .A(n44118), .B(n44119), .Z(n44117) );
  OR U53406 ( .A(n44120), .B(n44121), .Z(n44116) );
  ANDN U53407 ( .B(n44122), .A(n44123), .Z(n44074) );
  IV U53408 ( .A(n44124), .Z(n44122) );
  ANDN U53409 ( .B(n44125), .A(n44126), .Z(n44066) );
  XOR U53410 ( .A(n44052), .B(n44127), .Z(n44064) );
  XOR U53411 ( .A(n44053), .B(n44054), .Z(n44127) );
  XOR U53412 ( .A(n44059), .B(n44128), .Z(n44054) );
  XOR U53413 ( .A(n44058), .B(n44061), .Z(n44128) );
  IV U53414 ( .A(n44060), .Z(n44061) );
  NAND U53415 ( .A(n44129), .B(n44130), .Z(n44060) );
  OR U53416 ( .A(n44131), .B(n44132), .Z(n44130) );
  OR U53417 ( .A(n44133), .B(n44134), .Z(n44129) );
  NAND U53418 ( .A(n44135), .B(n44136), .Z(n44058) );
  OR U53419 ( .A(n44137), .B(n44138), .Z(n44136) );
  OR U53420 ( .A(n44139), .B(n44140), .Z(n44135) );
  NOR U53421 ( .A(n44141), .B(n44142), .Z(n44059) );
  ANDN U53422 ( .B(n44143), .A(n44144), .Z(n44053) );
  IV U53423 ( .A(n44145), .Z(n44143) );
  XNOR U53424 ( .A(n44046), .B(n44146), .Z(n44052) );
  XNOR U53425 ( .A(n44045), .B(n44047), .Z(n44146) );
  NAND U53426 ( .A(n44147), .B(n44148), .Z(n44047) );
  OR U53427 ( .A(n44149), .B(n44150), .Z(n44148) );
  OR U53428 ( .A(n44151), .B(n44152), .Z(n44147) );
  NAND U53429 ( .A(n44153), .B(n44154), .Z(n44045) );
  OR U53430 ( .A(n44155), .B(n44156), .Z(n44154) );
  OR U53431 ( .A(n44157), .B(n44158), .Z(n44153) );
  ANDN U53432 ( .B(n44159), .A(n44160), .Z(n44046) );
  IV U53433 ( .A(n44161), .Z(n44159) );
  XNOR U53434 ( .A(n44126), .B(n44125), .Z(N61489) );
  XOR U53435 ( .A(n44145), .B(n44144), .Z(n44125) );
  XNOR U53436 ( .A(n44160), .B(n44161), .Z(n44144) );
  XNOR U53437 ( .A(n44155), .B(n44156), .Z(n44161) );
  XNOR U53438 ( .A(n44157), .B(n44158), .Z(n44156) );
  XNOR U53439 ( .A(y[1669]), .B(x[1669]), .Z(n44158) );
  XNOR U53440 ( .A(y[1670]), .B(x[1670]), .Z(n44157) );
  XNOR U53441 ( .A(y[1668]), .B(x[1668]), .Z(n44155) );
  XNOR U53442 ( .A(n44149), .B(n44150), .Z(n44160) );
  XNOR U53443 ( .A(y[1665]), .B(x[1665]), .Z(n44150) );
  XNOR U53444 ( .A(n44151), .B(n44152), .Z(n44149) );
  XNOR U53445 ( .A(y[1666]), .B(x[1666]), .Z(n44152) );
  XNOR U53446 ( .A(y[1667]), .B(x[1667]), .Z(n44151) );
  XNOR U53447 ( .A(n44142), .B(n44141), .Z(n44145) );
  XNOR U53448 ( .A(n44137), .B(n44138), .Z(n44141) );
  XNOR U53449 ( .A(y[1662]), .B(x[1662]), .Z(n44138) );
  XNOR U53450 ( .A(n44139), .B(n44140), .Z(n44137) );
  XNOR U53451 ( .A(y[1663]), .B(x[1663]), .Z(n44140) );
  XNOR U53452 ( .A(y[1664]), .B(x[1664]), .Z(n44139) );
  XNOR U53453 ( .A(n44131), .B(n44132), .Z(n44142) );
  XNOR U53454 ( .A(y[1659]), .B(x[1659]), .Z(n44132) );
  XNOR U53455 ( .A(n44133), .B(n44134), .Z(n44131) );
  XNOR U53456 ( .A(y[1660]), .B(x[1660]), .Z(n44134) );
  XNOR U53457 ( .A(y[1661]), .B(x[1661]), .Z(n44133) );
  XOR U53458 ( .A(n44107), .B(n44108), .Z(n44126) );
  XNOR U53459 ( .A(n44123), .B(n44124), .Z(n44108) );
  XNOR U53460 ( .A(n44118), .B(n44119), .Z(n44124) );
  XNOR U53461 ( .A(n44120), .B(n44121), .Z(n44119) );
  XNOR U53462 ( .A(y[1657]), .B(x[1657]), .Z(n44121) );
  XNOR U53463 ( .A(y[1658]), .B(x[1658]), .Z(n44120) );
  XNOR U53464 ( .A(y[1656]), .B(x[1656]), .Z(n44118) );
  XNOR U53465 ( .A(n44112), .B(n44113), .Z(n44123) );
  XNOR U53466 ( .A(y[1653]), .B(x[1653]), .Z(n44113) );
  XNOR U53467 ( .A(n44114), .B(n44115), .Z(n44112) );
  XNOR U53468 ( .A(y[1654]), .B(x[1654]), .Z(n44115) );
  XNOR U53469 ( .A(y[1655]), .B(x[1655]), .Z(n44114) );
  XOR U53470 ( .A(n44106), .B(n44105), .Z(n44107) );
  XNOR U53471 ( .A(n44101), .B(n44102), .Z(n44105) );
  XNOR U53472 ( .A(y[1650]), .B(x[1650]), .Z(n44102) );
  XNOR U53473 ( .A(n44103), .B(n44104), .Z(n44101) );
  XNOR U53474 ( .A(y[1651]), .B(x[1651]), .Z(n44104) );
  XNOR U53475 ( .A(y[1652]), .B(x[1652]), .Z(n44103) );
  XNOR U53476 ( .A(n44095), .B(n44096), .Z(n44106) );
  XNOR U53477 ( .A(y[1647]), .B(x[1647]), .Z(n44096) );
  XNOR U53478 ( .A(n44097), .B(n44098), .Z(n44095) );
  XNOR U53479 ( .A(y[1648]), .B(x[1648]), .Z(n44098) );
  XNOR U53480 ( .A(y[1649]), .B(x[1649]), .Z(n44097) );
  NAND U53481 ( .A(n44162), .B(n44163), .Z(N61480) );
  NANDN U53482 ( .A(n44164), .B(n44165), .Z(n44163) );
  OR U53483 ( .A(n44166), .B(n44167), .Z(n44165) );
  NAND U53484 ( .A(n44166), .B(n44167), .Z(n44162) );
  XOR U53485 ( .A(n44166), .B(n44168), .Z(N61479) );
  XNOR U53486 ( .A(n44164), .B(n44167), .Z(n44168) );
  AND U53487 ( .A(n44169), .B(n44170), .Z(n44167) );
  NANDN U53488 ( .A(n44171), .B(n44172), .Z(n44170) );
  NANDN U53489 ( .A(n44173), .B(n44174), .Z(n44172) );
  NANDN U53490 ( .A(n44174), .B(n44173), .Z(n44169) );
  NAND U53491 ( .A(n44175), .B(n44176), .Z(n44164) );
  NANDN U53492 ( .A(n44177), .B(n44178), .Z(n44176) );
  OR U53493 ( .A(n44179), .B(n44180), .Z(n44178) );
  NAND U53494 ( .A(n44180), .B(n44179), .Z(n44175) );
  AND U53495 ( .A(n44181), .B(n44182), .Z(n44166) );
  NANDN U53496 ( .A(n44183), .B(n44184), .Z(n44182) );
  NANDN U53497 ( .A(n44185), .B(n44186), .Z(n44184) );
  NANDN U53498 ( .A(n44186), .B(n44185), .Z(n44181) );
  XOR U53499 ( .A(n44180), .B(n44187), .Z(N61478) );
  XOR U53500 ( .A(n44177), .B(n44179), .Z(n44187) );
  XNOR U53501 ( .A(n44173), .B(n44188), .Z(n44179) );
  XNOR U53502 ( .A(n44171), .B(n44174), .Z(n44188) );
  NAND U53503 ( .A(n44189), .B(n44190), .Z(n44174) );
  NAND U53504 ( .A(n44191), .B(n44192), .Z(n44190) );
  OR U53505 ( .A(n44193), .B(n44194), .Z(n44191) );
  NANDN U53506 ( .A(n44195), .B(n44193), .Z(n44189) );
  IV U53507 ( .A(n44194), .Z(n44195) );
  NAND U53508 ( .A(n44196), .B(n44197), .Z(n44171) );
  NAND U53509 ( .A(n44198), .B(n44199), .Z(n44197) );
  NANDN U53510 ( .A(n44200), .B(n44201), .Z(n44198) );
  NANDN U53511 ( .A(n44201), .B(n44200), .Z(n44196) );
  AND U53512 ( .A(n44202), .B(n44203), .Z(n44173) );
  NAND U53513 ( .A(n44204), .B(n44205), .Z(n44203) );
  OR U53514 ( .A(n44206), .B(n44207), .Z(n44204) );
  NANDN U53515 ( .A(n44208), .B(n44206), .Z(n44202) );
  NAND U53516 ( .A(n44209), .B(n44210), .Z(n44177) );
  NANDN U53517 ( .A(n44211), .B(n44212), .Z(n44210) );
  OR U53518 ( .A(n44213), .B(n44214), .Z(n44212) );
  NANDN U53519 ( .A(n44215), .B(n44213), .Z(n44209) );
  IV U53520 ( .A(n44214), .Z(n44215) );
  XNOR U53521 ( .A(n44185), .B(n44216), .Z(n44180) );
  XNOR U53522 ( .A(n44183), .B(n44186), .Z(n44216) );
  NAND U53523 ( .A(n44217), .B(n44218), .Z(n44186) );
  NAND U53524 ( .A(n44219), .B(n44220), .Z(n44218) );
  OR U53525 ( .A(n44221), .B(n44222), .Z(n44219) );
  NANDN U53526 ( .A(n44223), .B(n44221), .Z(n44217) );
  IV U53527 ( .A(n44222), .Z(n44223) );
  NAND U53528 ( .A(n44224), .B(n44225), .Z(n44183) );
  NAND U53529 ( .A(n44226), .B(n44227), .Z(n44225) );
  NANDN U53530 ( .A(n44228), .B(n44229), .Z(n44226) );
  NANDN U53531 ( .A(n44229), .B(n44228), .Z(n44224) );
  AND U53532 ( .A(n44230), .B(n44231), .Z(n44185) );
  NAND U53533 ( .A(n44232), .B(n44233), .Z(n44231) );
  OR U53534 ( .A(n44234), .B(n44235), .Z(n44232) );
  NANDN U53535 ( .A(n44236), .B(n44234), .Z(n44230) );
  XNOR U53536 ( .A(n44211), .B(n44237), .Z(N61477) );
  XOR U53537 ( .A(n44213), .B(n44214), .Z(n44237) );
  XNOR U53538 ( .A(n44227), .B(n44238), .Z(n44214) );
  XOR U53539 ( .A(n44228), .B(n44229), .Z(n44238) );
  XOR U53540 ( .A(n44234), .B(n44239), .Z(n44229) );
  XOR U53541 ( .A(n44233), .B(n44236), .Z(n44239) );
  IV U53542 ( .A(n44235), .Z(n44236) );
  NAND U53543 ( .A(n44240), .B(n44241), .Z(n44235) );
  OR U53544 ( .A(n44242), .B(n44243), .Z(n44241) );
  OR U53545 ( .A(n44244), .B(n44245), .Z(n44240) );
  NAND U53546 ( .A(n44246), .B(n44247), .Z(n44233) );
  OR U53547 ( .A(n44248), .B(n44249), .Z(n44247) );
  OR U53548 ( .A(n44250), .B(n44251), .Z(n44246) );
  NOR U53549 ( .A(n44252), .B(n44253), .Z(n44234) );
  ANDN U53550 ( .B(n44254), .A(n44255), .Z(n44228) );
  XNOR U53551 ( .A(n44221), .B(n44256), .Z(n44227) );
  XNOR U53552 ( .A(n44220), .B(n44222), .Z(n44256) );
  NAND U53553 ( .A(n44257), .B(n44258), .Z(n44222) );
  OR U53554 ( .A(n44259), .B(n44260), .Z(n44258) );
  OR U53555 ( .A(n44261), .B(n44262), .Z(n44257) );
  NAND U53556 ( .A(n44263), .B(n44264), .Z(n44220) );
  OR U53557 ( .A(n44265), .B(n44266), .Z(n44264) );
  OR U53558 ( .A(n44267), .B(n44268), .Z(n44263) );
  ANDN U53559 ( .B(n44269), .A(n44270), .Z(n44221) );
  IV U53560 ( .A(n44271), .Z(n44269) );
  ANDN U53561 ( .B(n44272), .A(n44273), .Z(n44213) );
  XOR U53562 ( .A(n44199), .B(n44274), .Z(n44211) );
  XOR U53563 ( .A(n44200), .B(n44201), .Z(n44274) );
  XOR U53564 ( .A(n44206), .B(n44275), .Z(n44201) );
  XOR U53565 ( .A(n44205), .B(n44208), .Z(n44275) );
  IV U53566 ( .A(n44207), .Z(n44208) );
  NAND U53567 ( .A(n44276), .B(n44277), .Z(n44207) );
  OR U53568 ( .A(n44278), .B(n44279), .Z(n44277) );
  OR U53569 ( .A(n44280), .B(n44281), .Z(n44276) );
  NAND U53570 ( .A(n44282), .B(n44283), .Z(n44205) );
  OR U53571 ( .A(n44284), .B(n44285), .Z(n44283) );
  OR U53572 ( .A(n44286), .B(n44287), .Z(n44282) );
  NOR U53573 ( .A(n44288), .B(n44289), .Z(n44206) );
  ANDN U53574 ( .B(n44290), .A(n44291), .Z(n44200) );
  IV U53575 ( .A(n44292), .Z(n44290) );
  XNOR U53576 ( .A(n44193), .B(n44293), .Z(n44199) );
  XNOR U53577 ( .A(n44192), .B(n44194), .Z(n44293) );
  NAND U53578 ( .A(n44294), .B(n44295), .Z(n44194) );
  OR U53579 ( .A(n44296), .B(n44297), .Z(n44295) );
  OR U53580 ( .A(n44298), .B(n44299), .Z(n44294) );
  NAND U53581 ( .A(n44300), .B(n44301), .Z(n44192) );
  OR U53582 ( .A(n44302), .B(n44303), .Z(n44301) );
  OR U53583 ( .A(n44304), .B(n44305), .Z(n44300) );
  ANDN U53584 ( .B(n44306), .A(n44307), .Z(n44193) );
  IV U53585 ( .A(n44308), .Z(n44306) );
  XNOR U53586 ( .A(n44273), .B(n44272), .Z(N61476) );
  XOR U53587 ( .A(n44292), .B(n44291), .Z(n44272) );
  XNOR U53588 ( .A(n44307), .B(n44308), .Z(n44291) );
  XNOR U53589 ( .A(n44302), .B(n44303), .Z(n44308) );
  XNOR U53590 ( .A(n44304), .B(n44305), .Z(n44303) );
  XNOR U53591 ( .A(y[1645]), .B(x[1645]), .Z(n44305) );
  XNOR U53592 ( .A(y[1646]), .B(x[1646]), .Z(n44304) );
  XNOR U53593 ( .A(y[1644]), .B(x[1644]), .Z(n44302) );
  XNOR U53594 ( .A(n44296), .B(n44297), .Z(n44307) );
  XNOR U53595 ( .A(y[1641]), .B(x[1641]), .Z(n44297) );
  XNOR U53596 ( .A(n44298), .B(n44299), .Z(n44296) );
  XNOR U53597 ( .A(y[1642]), .B(x[1642]), .Z(n44299) );
  XNOR U53598 ( .A(y[1643]), .B(x[1643]), .Z(n44298) );
  XNOR U53599 ( .A(n44289), .B(n44288), .Z(n44292) );
  XNOR U53600 ( .A(n44284), .B(n44285), .Z(n44288) );
  XNOR U53601 ( .A(y[1638]), .B(x[1638]), .Z(n44285) );
  XNOR U53602 ( .A(n44286), .B(n44287), .Z(n44284) );
  XNOR U53603 ( .A(y[1639]), .B(x[1639]), .Z(n44287) );
  XNOR U53604 ( .A(y[1640]), .B(x[1640]), .Z(n44286) );
  XNOR U53605 ( .A(n44278), .B(n44279), .Z(n44289) );
  XNOR U53606 ( .A(y[1635]), .B(x[1635]), .Z(n44279) );
  XNOR U53607 ( .A(n44280), .B(n44281), .Z(n44278) );
  XNOR U53608 ( .A(y[1636]), .B(x[1636]), .Z(n44281) );
  XNOR U53609 ( .A(y[1637]), .B(x[1637]), .Z(n44280) );
  XOR U53610 ( .A(n44254), .B(n44255), .Z(n44273) );
  XNOR U53611 ( .A(n44270), .B(n44271), .Z(n44255) );
  XNOR U53612 ( .A(n44265), .B(n44266), .Z(n44271) );
  XNOR U53613 ( .A(n44267), .B(n44268), .Z(n44266) );
  XNOR U53614 ( .A(y[1633]), .B(x[1633]), .Z(n44268) );
  XNOR U53615 ( .A(y[1634]), .B(x[1634]), .Z(n44267) );
  XNOR U53616 ( .A(y[1632]), .B(x[1632]), .Z(n44265) );
  XNOR U53617 ( .A(n44259), .B(n44260), .Z(n44270) );
  XNOR U53618 ( .A(y[1629]), .B(x[1629]), .Z(n44260) );
  XNOR U53619 ( .A(n44261), .B(n44262), .Z(n44259) );
  XNOR U53620 ( .A(y[1630]), .B(x[1630]), .Z(n44262) );
  XNOR U53621 ( .A(y[1631]), .B(x[1631]), .Z(n44261) );
  XOR U53622 ( .A(n44253), .B(n44252), .Z(n44254) );
  XNOR U53623 ( .A(n44248), .B(n44249), .Z(n44252) );
  XNOR U53624 ( .A(y[1626]), .B(x[1626]), .Z(n44249) );
  XNOR U53625 ( .A(n44250), .B(n44251), .Z(n44248) );
  XNOR U53626 ( .A(y[1627]), .B(x[1627]), .Z(n44251) );
  XNOR U53627 ( .A(y[1628]), .B(x[1628]), .Z(n44250) );
  XNOR U53628 ( .A(n44242), .B(n44243), .Z(n44253) );
  XNOR U53629 ( .A(y[1623]), .B(x[1623]), .Z(n44243) );
  XNOR U53630 ( .A(n44244), .B(n44245), .Z(n44242) );
  XNOR U53631 ( .A(y[1624]), .B(x[1624]), .Z(n44245) );
  XNOR U53632 ( .A(y[1625]), .B(x[1625]), .Z(n44244) );
  NAND U53633 ( .A(n44309), .B(n44310), .Z(N61467) );
  NANDN U53634 ( .A(n44311), .B(n44312), .Z(n44310) );
  OR U53635 ( .A(n44313), .B(n44314), .Z(n44312) );
  NAND U53636 ( .A(n44313), .B(n44314), .Z(n44309) );
  XOR U53637 ( .A(n44313), .B(n44315), .Z(N61466) );
  XNOR U53638 ( .A(n44311), .B(n44314), .Z(n44315) );
  AND U53639 ( .A(n44316), .B(n44317), .Z(n44314) );
  NANDN U53640 ( .A(n44318), .B(n44319), .Z(n44317) );
  NANDN U53641 ( .A(n44320), .B(n44321), .Z(n44319) );
  NANDN U53642 ( .A(n44321), .B(n44320), .Z(n44316) );
  NAND U53643 ( .A(n44322), .B(n44323), .Z(n44311) );
  NANDN U53644 ( .A(n44324), .B(n44325), .Z(n44323) );
  OR U53645 ( .A(n44326), .B(n44327), .Z(n44325) );
  NAND U53646 ( .A(n44327), .B(n44326), .Z(n44322) );
  AND U53647 ( .A(n44328), .B(n44329), .Z(n44313) );
  NANDN U53648 ( .A(n44330), .B(n44331), .Z(n44329) );
  NANDN U53649 ( .A(n44332), .B(n44333), .Z(n44331) );
  NANDN U53650 ( .A(n44333), .B(n44332), .Z(n44328) );
  XOR U53651 ( .A(n44327), .B(n44334), .Z(N61465) );
  XOR U53652 ( .A(n44324), .B(n44326), .Z(n44334) );
  XNOR U53653 ( .A(n44320), .B(n44335), .Z(n44326) );
  XNOR U53654 ( .A(n44318), .B(n44321), .Z(n44335) );
  NAND U53655 ( .A(n44336), .B(n44337), .Z(n44321) );
  NAND U53656 ( .A(n44338), .B(n44339), .Z(n44337) );
  OR U53657 ( .A(n44340), .B(n44341), .Z(n44338) );
  NANDN U53658 ( .A(n44342), .B(n44340), .Z(n44336) );
  IV U53659 ( .A(n44341), .Z(n44342) );
  NAND U53660 ( .A(n44343), .B(n44344), .Z(n44318) );
  NAND U53661 ( .A(n44345), .B(n44346), .Z(n44344) );
  NANDN U53662 ( .A(n44347), .B(n44348), .Z(n44345) );
  NANDN U53663 ( .A(n44348), .B(n44347), .Z(n44343) );
  AND U53664 ( .A(n44349), .B(n44350), .Z(n44320) );
  NAND U53665 ( .A(n44351), .B(n44352), .Z(n44350) );
  OR U53666 ( .A(n44353), .B(n44354), .Z(n44351) );
  NANDN U53667 ( .A(n44355), .B(n44353), .Z(n44349) );
  NAND U53668 ( .A(n44356), .B(n44357), .Z(n44324) );
  NANDN U53669 ( .A(n44358), .B(n44359), .Z(n44357) );
  OR U53670 ( .A(n44360), .B(n44361), .Z(n44359) );
  NANDN U53671 ( .A(n44362), .B(n44360), .Z(n44356) );
  IV U53672 ( .A(n44361), .Z(n44362) );
  XNOR U53673 ( .A(n44332), .B(n44363), .Z(n44327) );
  XNOR U53674 ( .A(n44330), .B(n44333), .Z(n44363) );
  NAND U53675 ( .A(n44364), .B(n44365), .Z(n44333) );
  NAND U53676 ( .A(n44366), .B(n44367), .Z(n44365) );
  OR U53677 ( .A(n44368), .B(n44369), .Z(n44366) );
  NANDN U53678 ( .A(n44370), .B(n44368), .Z(n44364) );
  IV U53679 ( .A(n44369), .Z(n44370) );
  NAND U53680 ( .A(n44371), .B(n44372), .Z(n44330) );
  NAND U53681 ( .A(n44373), .B(n44374), .Z(n44372) );
  NANDN U53682 ( .A(n44375), .B(n44376), .Z(n44373) );
  NANDN U53683 ( .A(n44376), .B(n44375), .Z(n44371) );
  AND U53684 ( .A(n44377), .B(n44378), .Z(n44332) );
  NAND U53685 ( .A(n44379), .B(n44380), .Z(n44378) );
  OR U53686 ( .A(n44381), .B(n44382), .Z(n44379) );
  NANDN U53687 ( .A(n44383), .B(n44381), .Z(n44377) );
  XNOR U53688 ( .A(n44358), .B(n44384), .Z(N61464) );
  XOR U53689 ( .A(n44360), .B(n44361), .Z(n44384) );
  XNOR U53690 ( .A(n44374), .B(n44385), .Z(n44361) );
  XOR U53691 ( .A(n44375), .B(n44376), .Z(n44385) );
  XOR U53692 ( .A(n44381), .B(n44386), .Z(n44376) );
  XOR U53693 ( .A(n44380), .B(n44383), .Z(n44386) );
  IV U53694 ( .A(n44382), .Z(n44383) );
  NAND U53695 ( .A(n44387), .B(n44388), .Z(n44382) );
  OR U53696 ( .A(n44389), .B(n44390), .Z(n44388) );
  OR U53697 ( .A(n44391), .B(n44392), .Z(n44387) );
  NAND U53698 ( .A(n44393), .B(n44394), .Z(n44380) );
  OR U53699 ( .A(n44395), .B(n44396), .Z(n44394) );
  OR U53700 ( .A(n44397), .B(n44398), .Z(n44393) );
  NOR U53701 ( .A(n44399), .B(n44400), .Z(n44381) );
  ANDN U53702 ( .B(n44401), .A(n44402), .Z(n44375) );
  XNOR U53703 ( .A(n44368), .B(n44403), .Z(n44374) );
  XNOR U53704 ( .A(n44367), .B(n44369), .Z(n44403) );
  NAND U53705 ( .A(n44404), .B(n44405), .Z(n44369) );
  OR U53706 ( .A(n44406), .B(n44407), .Z(n44405) );
  OR U53707 ( .A(n44408), .B(n44409), .Z(n44404) );
  NAND U53708 ( .A(n44410), .B(n44411), .Z(n44367) );
  OR U53709 ( .A(n44412), .B(n44413), .Z(n44411) );
  OR U53710 ( .A(n44414), .B(n44415), .Z(n44410) );
  ANDN U53711 ( .B(n44416), .A(n44417), .Z(n44368) );
  IV U53712 ( .A(n44418), .Z(n44416) );
  ANDN U53713 ( .B(n44419), .A(n44420), .Z(n44360) );
  XOR U53714 ( .A(n44346), .B(n44421), .Z(n44358) );
  XOR U53715 ( .A(n44347), .B(n44348), .Z(n44421) );
  XOR U53716 ( .A(n44353), .B(n44422), .Z(n44348) );
  XOR U53717 ( .A(n44352), .B(n44355), .Z(n44422) );
  IV U53718 ( .A(n44354), .Z(n44355) );
  NAND U53719 ( .A(n44423), .B(n44424), .Z(n44354) );
  OR U53720 ( .A(n44425), .B(n44426), .Z(n44424) );
  OR U53721 ( .A(n44427), .B(n44428), .Z(n44423) );
  NAND U53722 ( .A(n44429), .B(n44430), .Z(n44352) );
  OR U53723 ( .A(n44431), .B(n44432), .Z(n44430) );
  OR U53724 ( .A(n44433), .B(n44434), .Z(n44429) );
  NOR U53725 ( .A(n44435), .B(n44436), .Z(n44353) );
  ANDN U53726 ( .B(n44437), .A(n44438), .Z(n44347) );
  IV U53727 ( .A(n44439), .Z(n44437) );
  XNOR U53728 ( .A(n44340), .B(n44440), .Z(n44346) );
  XNOR U53729 ( .A(n44339), .B(n44341), .Z(n44440) );
  NAND U53730 ( .A(n44441), .B(n44442), .Z(n44341) );
  OR U53731 ( .A(n44443), .B(n44444), .Z(n44442) );
  OR U53732 ( .A(n44445), .B(n44446), .Z(n44441) );
  NAND U53733 ( .A(n44447), .B(n44448), .Z(n44339) );
  OR U53734 ( .A(n44449), .B(n44450), .Z(n44448) );
  OR U53735 ( .A(n44451), .B(n44452), .Z(n44447) );
  ANDN U53736 ( .B(n44453), .A(n44454), .Z(n44340) );
  IV U53737 ( .A(n44455), .Z(n44453) );
  XNOR U53738 ( .A(n44420), .B(n44419), .Z(N61463) );
  XOR U53739 ( .A(n44439), .B(n44438), .Z(n44419) );
  XNOR U53740 ( .A(n44454), .B(n44455), .Z(n44438) );
  XNOR U53741 ( .A(n44449), .B(n44450), .Z(n44455) );
  XNOR U53742 ( .A(n44451), .B(n44452), .Z(n44450) );
  XNOR U53743 ( .A(y[1621]), .B(x[1621]), .Z(n44452) );
  XNOR U53744 ( .A(y[1622]), .B(x[1622]), .Z(n44451) );
  XNOR U53745 ( .A(y[1620]), .B(x[1620]), .Z(n44449) );
  XNOR U53746 ( .A(n44443), .B(n44444), .Z(n44454) );
  XNOR U53747 ( .A(y[1617]), .B(x[1617]), .Z(n44444) );
  XNOR U53748 ( .A(n44445), .B(n44446), .Z(n44443) );
  XNOR U53749 ( .A(y[1618]), .B(x[1618]), .Z(n44446) );
  XNOR U53750 ( .A(y[1619]), .B(x[1619]), .Z(n44445) );
  XNOR U53751 ( .A(n44436), .B(n44435), .Z(n44439) );
  XNOR U53752 ( .A(n44431), .B(n44432), .Z(n44435) );
  XNOR U53753 ( .A(y[1614]), .B(x[1614]), .Z(n44432) );
  XNOR U53754 ( .A(n44433), .B(n44434), .Z(n44431) );
  XNOR U53755 ( .A(y[1615]), .B(x[1615]), .Z(n44434) );
  XNOR U53756 ( .A(y[1616]), .B(x[1616]), .Z(n44433) );
  XNOR U53757 ( .A(n44425), .B(n44426), .Z(n44436) );
  XNOR U53758 ( .A(y[1611]), .B(x[1611]), .Z(n44426) );
  XNOR U53759 ( .A(n44427), .B(n44428), .Z(n44425) );
  XNOR U53760 ( .A(y[1612]), .B(x[1612]), .Z(n44428) );
  XNOR U53761 ( .A(y[1613]), .B(x[1613]), .Z(n44427) );
  XOR U53762 ( .A(n44401), .B(n44402), .Z(n44420) );
  XNOR U53763 ( .A(n44417), .B(n44418), .Z(n44402) );
  XNOR U53764 ( .A(n44412), .B(n44413), .Z(n44418) );
  XNOR U53765 ( .A(n44414), .B(n44415), .Z(n44413) );
  XNOR U53766 ( .A(y[1609]), .B(x[1609]), .Z(n44415) );
  XNOR U53767 ( .A(y[1610]), .B(x[1610]), .Z(n44414) );
  XNOR U53768 ( .A(y[1608]), .B(x[1608]), .Z(n44412) );
  XNOR U53769 ( .A(n44406), .B(n44407), .Z(n44417) );
  XNOR U53770 ( .A(y[1605]), .B(x[1605]), .Z(n44407) );
  XNOR U53771 ( .A(n44408), .B(n44409), .Z(n44406) );
  XNOR U53772 ( .A(y[1606]), .B(x[1606]), .Z(n44409) );
  XNOR U53773 ( .A(y[1607]), .B(x[1607]), .Z(n44408) );
  XOR U53774 ( .A(n44400), .B(n44399), .Z(n44401) );
  XNOR U53775 ( .A(n44395), .B(n44396), .Z(n44399) );
  XNOR U53776 ( .A(y[1602]), .B(x[1602]), .Z(n44396) );
  XNOR U53777 ( .A(n44397), .B(n44398), .Z(n44395) );
  XNOR U53778 ( .A(y[1603]), .B(x[1603]), .Z(n44398) );
  XNOR U53779 ( .A(y[1604]), .B(x[1604]), .Z(n44397) );
  XNOR U53780 ( .A(n44389), .B(n44390), .Z(n44400) );
  XNOR U53781 ( .A(y[1599]), .B(x[1599]), .Z(n44390) );
  XNOR U53782 ( .A(n44391), .B(n44392), .Z(n44389) );
  XNOR U53783 ( .A(y[1600]), .B(x[1600]), .Z(n44392) );
  XNOR U53784 ( .A(y[1601]), .B(x[1601]), .Z(n44391) );
  NAND U53785 ( .A(n44456), .B(n44457), .Z(N61454) );
  NANDN U53786 ( .A(n44458), .B(n44459), .Z(n44457) );
  OR U53787 ( .A(n44460), .B(n44461), .Z(n44459) );
  NAND U53788 ( .A(n44460), .B(n44461), .Z(n44456) );
  XOR U53789 ( .A(n44460), .B(n44462), .Z(N61453) );
  XNOR U53790 ( .A(n44458), .B(n44461), .Z(n44462) );
  AND U53791 ( .A(n44463), .B(n44464), .Z(n44461) );
  NANDN U53792 ( .A(n44465), .B(n44466), .Z(n44464) );
  NANDN U53793 ( .A(n44467), .B(n44468), .Z(n44466) );
  NANDN U53794 ( .A(n44468), .B(n44467), .Z(n44463) );
  NAND U53795 ( .A(n44469), .B(n44470), .Z(n44458) );
  NANDN U53796 ( .A(n44471), .B(n44472), .Z(n44470) );
  OR U53797 ( .A(n44473), .B(n44474), .Z(n44472) );
  NAND U53798 ( .A(n44474), .B(n44473), .Z(n44469) );
  AND U53799 ( .A(n44475), .B(n44476), .Z(n44460) );
  NANDN U53800 ( .A(n44477), .B(n44478), .Z(n44476) );
  NANDN U53801 ( .A(n44479), .B(n44480), .Z(n44478) );
  NANDN U53802 ( .A(n44480), .B(n44479), .Z(n44475) );
  XOR U53803 ( .A(n44474), .B(n44481), .Z(N61452) );
  XOR U53804 ( .A(n44471), .B(n44473), .Z(n44481) );
  XNOR U53805 ( .A(n44467), .B(n44482), .Z(n44473) );
  XNOR U53806 ( .A(n44465), .B(n44468), .Z(n44482) );
  NAND U53807 ( .A(n44483), .B(n44484), .Z(n44468) );
  NAND U53808 ( .A(n44485), .B(n44486), .Z(n44484) );
  OR U53809 ( .A(n44487), .B(n44488), .Z(n44485) );
  NANDN U53810 ( .A(n44489), .B(n44487), .Z(n44483) );
  IV U53811 ( .A(n44488), .Z(n44489) );
  NAND U53812 ( .A(n44490), .B(n44491), .Z(n44465) );
  NAND U53813 ( .A(n44492), .B(n44493), .Z(n44491) );
  NANDN U53814 ( .A(n44494), .B(n44495), .Z(n44492) );
  NANDN U53815 ( .A(n44495), .B(n44494), .Z(n44490) );
  AND U53816 ( .A(n44496), .B(n44497), .Z(n44467) );
  NAND U53817 ( .A(n44498), .B(n44499), .Z(n44497) );
  OR U53818 ( .A(n44500), .B(n44501), .Z(n44498) );
  NANDN U53819 ( .A(n44502), .B(n44500), .Z(n44496) );
  NAND U53820 ( .A(n44503), .B(n44504), .Z(n44471) );
  NANDN U53821 ( .A(n44505), .B(n44506), .Z(n44504) );
  OR U53822 ( .A(n44507), .B(n44508), .Z(n44506) );
  NANDN U53823 ( .A(n44509), .B(n44507), .Z(n44503) );
  IV U53824 ( .A(n44508), .Z(n44509) );
  XNOR U53825 ( .A(n44479), .B(n44510), .Z(n44474) );
  XNOR U53826 ( .A(n44477), .B(n44480), .Z(n44510) );
  NAND U53827 ( .A(n44511), .B(n44512), .Z(n44480) );
  NAND U53828 ( .A(n44513), .B(n44514), .Z(n44512) );
  OR U53829 ( .A(n44515), .B(n44516), .Z(n44513) );
  NANDN U53830 ( .A(n44517), .B(n44515), .Z(n44511) );
  IV U53831 ( .A(n44516), .Z(n44517) );
  NAND U53832 ( .A(n44518), .B(n44519), .Z(n44477) );
  NAND U53833 ( .A(n44520), .B(n44521), .Z(n44519) );
  NANDN U53834 ( .A(n44522), .B(n44523), .Z(n44520) );
  NANDN U53835 ( .A(n44523), .B(n44522), .Z(n44518) );
  AND U53836 ( .A(n44524), .B(n44525), .Z(n44479) );
  NAND U53837 ( .A(n44526), .B(n44527), .Z(n44525) );
  OR U53838 ( .A(n44528), .B(n44529), .Z(n44526) );
  NANDN U53839 ( .A(n44530), .B(n44528), .Z(n44524) );
  XNOR U53840 ( .A(n44505), .B(n44531), .Z(N61451) );
  XOR U53841 ( .A(n44507), .B(n44508), .Z(n44531) );
  XNOR U53842 ( .A(n44521), .B(n44532), .Z(n44508) );
  XOR U53843 ( .A(n44522), .B(n44523), .Z(n44532) );
  XOR U53844 ( .A(n44528), .B(n44533), .Z(n44523) );
  XOR U53845 ( .A(n44527), .B(n44530), .Z(n44533) );
  IV U53846 ( .A(n44529), .Z(n44530) );
  NAND U53847 ( .A(n44534), .B(n44535), .Z(n44529) );
  OR U53848 ( .A(n44536), .B(n44537), .Z(n44535) );
  OR U53849 ( .A(n44538), .B(n44539), .Z(n44534) );
  NAND U53850 ( .A(n44540), .B(n44541), .Z(n44527) );
  OR U53851 ( .A(n44542), .B(n44543), .Z(n44541) );
  OR U53852 ( .A(n44544), .B(n44545), .Z(n44540) );
  NOR U53853 ( .A(n44546), .B(n44547), .Z(n44528) );
  ANDN U53854 ( .B(n44548), .A(n44549), .Z(n44522) );
  XNOR U53855 ( .A(n44515), .B(n44550), .Z(n44521) );
  XNOR U53856 ( .A(n44514), .B(n44516), .Z(n44550) );
  NAND U53857 ( .A(n44551), .B(n44552), .Z(n44516) );
  OR U53858 ( .A(n44553), .B(n44554), .Z(n44552) );
  OR U53859 ( .A(n44555), .B(n44556), .Z(n44551) );
  NAND U53860 ( .A(n44557), .B(n44558), .Z(n44514) );
  OR U53861 ( .A(n44559), .B(n44560), .Z(n44558) );
  OR U53862 ( .A(n44561), .B(n44562), .Z(n44557) );
  ANDN U53863 ( .B(n44563), .A(n44564), .Z(n44515) );
  IV U53864 ( .A(n44565), .Z(n44563) );
  ANDN U53865 ( .B(n44566), .A(n44567), .Z(n44507) );
  XOR U53866 ( .A(n44493), .B(n44568), .Z(n44505) );
  XOR U53867 ( .A(n44494), .B(n44495), .Z(n44568) );
  XOR U53868 ( .A(n44500), .B(n44569), .Z(n44495) );
  XOR U53869 ( .A(n44499), .B(n44502), .Z(n44569) );
  IV U53870 ( .A(n44501), .Z(n44502) );
  NAND U53871 ( .A(n44570), .B(n44571), .Z(n44501) );
  OR U53872 ( .A(n44572), .B(n44573), .Z(n44571) );
  OR U53873 ( .A(n44574), .B(n44575), .Z(n44570) );
  NAND U53874 ( .A(n44576), .B(n44577), .Z(n44499) );
  OR U53875 ( .A(n44578), .B(n44579), .Z(n44577) );
  OR U53876 ( .A(n44580), .B(n44581), .Z(n44576) );
  NOR U53877 ( .A(n44582), .B(n44583), .Z(n44500) );
  ANDN U53878 ( .B(n44584), .A(n44585), .Z(n44494) );
  IV U53879 ( .A(n44586), .Z(n44584) );
  XNOR U53880 ( .A(n44487), .B(n44587), .Z(n44493) );
  XNOR U53881 ( .A(n44486), .B(n44488), .Z(n44587) );
  NAND U53882 ( .A(n44588), .B(n44589), .Z(n44488) );
  OR U53883 ( .A(n44590), .B(n44591), .Z(n44589) );
  OR U53884 ( .A(n44592), .B(n44593), .Z(n44588) );
  NAND U53885 ( .A(n44594), .B(n44595), .Z(n44486) );
  OR U53886 ( .A(n44596), .B(n44597), .Z(n44595) );
  OR U53887 ( .A(n44598), .B(n44599), .Z(n44594) );
  ANDN U53888 ( .B(n44600), .A(n44601), .Z(n44487) );
  IV U53889 ( .A(n44602), .Z(n44600) );
  XNOR U53890 ( .A(n44567), .B(n44566), .Z(N61450) );
  XOR U53891 ( .A(n44586), .B(n44585), .Z(n44566) );
  XNOR U53892 ( .A(n44601), .B(n44602), .Z(n44585) );
  XNOR U53893 ( .A(n44596), .B(n44597), .Z(n44602) );
  XNOR U53894 ( .A(n44598), .B(n44599), .Z(n44597) );
  XNOR U53895 ( .A(y[1597]), .B(x[1597]), .Z(n44599) );
  XNOR U53896 ( .A(y[1598]), .B(x[1598]), .Z(n44598) );
  XNOR U53897 ( .A(y[1596]), .B(x[1596]), .Z(n44596) );
  XNOR U53898 ( .A(n44590), .B(n44591), .Z(n44601) );
  XNOR U53899 ( .A(y[1593]), .B(x[1593]), .Z(n44591) );
  XNOR U53900 ( .A(n44592), .B(n44593), .Z(n44590) );
  XNOR U53901 ( .A(y[1594]), .B(x[1594]), .Z(n44593) );
  XNOR U53902 ( .A(y[1595]), .B(x[1595]), .Z(n44592) );
  XNOR U53903 ( .A(n44583), .B(n44582), .Z(n44586) );
  XNOR U53904 ( .A(n44578), .B(n44579), .Z(n44582) );
  XNOR U53905 ( .A(y[1590]), .B(x[1590]), .Z(n44579) );
  XNOR U53906 ( .A(n44580), .B(n44581), .Z(n44578) );
  XNOR U53907 ( .A(y[1591]), .B(x[1591]), .Z(n44581) );
  XNOR U53908 ( .A(y[1592]), .B(x[1592]), .Z(n44580) );
  XNOR U53909 ( .A(n44572), .B(n44573), .Z(n44583) );
  XNOR U53910 ( .A(y[1587]), .B(x[1587]), .Z(n44573) );
  XNOR U53911 ( .A(n44574), .B(n44575), .Z(n44572) );
  XNOR U53912 ( .A(y[1588]), .B(x[1588]), .Z(n44575) );
  XNOR U53913 ( .A(y[1589]), .B(x[1589]), .Z(n44574) );
  XOR U53914 ( .A(n44548), .B(n44549), .Z(n44567) );
  XNOR U53915 ( .A(n44564), .B(n44565), .Z(n44549) );
  XNOR U53916 ( .A(n44559), .B(n44560), .Z(n44565) );
  XNOR U53917 ( .A(n44561), .B(n44562), .Z(n44560) );
  XNOR U53918 ( .A(y[1585]), .B(x[1585]), .Z(n44562) );
  XNOR U53919 ( .A(y[1586]), .B(x[1586]), .Z(n44561) );
  XNOR U53920 ( .A(y[1584]), .B(x[1584]), .Z(n44559) );
  XNOR U53921 ( .A(n44553), .B(n44554), .Z(n44564) );
  XNOR U53922 ( .A(y[1581]), .B(x[1581]), .Z(n44554) );
  XNOR U53923 ( .A(n44555), .B(n44556), .Z(n44553) );
  XNOR U53924 ( .A(y[1582]), .B(x[1582]), .Z(n44556) );
  XNOR U53925 ( .A(y[1583]), .B(x[1583]), .Z(n44555) );
  XOR U53926 ( .A(n44547), .B(n44546), .Z(n44548) );
  XNOR U53927 ( .A(n44542), .B(n44543), .Z(n44546) );
  XNOR U53928 ( .A(y[1578]), .B(x[1578]), .Z(n44543) );
  XNOR U53929 ( .A(n44544), .B(n44545), .Z(n44542) );
  XNOR U53930 ( .A(y[1579]), .B(x[1579]), .Z(n44545) );
  XNOR U53931 ( .A(y[1580]), .B(x[1580]), .Z(n44544) );
  XNOR U53932 ( .A(n44536), .B(n44537), .Z(n44547) );
  XNOR U53933 ( .A(y[1575]), .B(x[1575]), .Z(n44537) );
  XNOR U53934 ( .A(n44538), .B(n44539), .Z(n44536) );
  XNOR U53935 ( .A(y[1576]), .B(x[1576]), .Z(n44539) );
  XNOR U53936 ( .A(y[1577]), .B(x[1577]), .Z(n44538) );
  NAND U53937 ( .A(n44603), .B(n44604), .Z(N61441) );
  NANDN U53938 ( .A(n44605), .B(n44606), .Z(n44604) );
  OR U53939 ( .A(n44607), .B(n44608), .Z(n44606) );
  NAND U53940 ( .A(n44607), .B(n44608), .Z(n44603) );
  XOR U53941 ( .A(n44607), .B(n44609), .Z(N61440) );
  XNOR U53942 ( .A(n44605), .B(n44608), .Z(n44609) );
  AND U53943 ( .A(n44610), .B(n44611), .Z(n44608) );
  NANDN U53944 ( .A(n44612), .B(n44613), .Z(n44611) );
  NANDN U53945 ( .A(n44614), .B(n44615), .Z(n44613) );
  NANDN U53946 ( .A(n44615), .B(n44614), .Z(n44610) );
  NAND U53947 ( .A(n44616), .B(n44617), .Z(n44605) );
  NANDN U53948 ( .A(n44618), .B(n44619), .Z(n44617) );
  OR U53949 ( .A(n44620), .B(n44621), .Z(n44619) );
  NAND U53950 ( .A(n44621), .B(n44620), .Z(n44616) );
  AND U53951 ( .A(n44622), .B(n44623), .Z(n44607) );
  NANDN U53952 ( .A(n44624), .B(n44625), .Z(n44623) );
  NANDN U53953 ( .A(n44626), .B(n44627), .Z(n44625) );
  NANDN U53954 ( .A(n44627), .B(n44626), .Z(n44622) );
  XOR U53955 ( .A(n44621), .B(n44628), .Z(N61439) );
  XOR U53956 ( .A(n44618), .B(n44620), .Z(n44628) );
  XNOR U53957 ( .A(n44614), .B(n44629), .Z(n44620) );
  XNOR U53958 ( .A(n44612), .B(n44615), .Z(n44629) );
  NAND U53959 ( .A(n44630), .B(n44631), .Z(n44615) );
  NAND U53960 ( .A(n44632), .B(n44633), .Z(n44631) );
  OR U53961 ( .A(n44634), .B(n44635), .Z(n44632) );
  NANDN U53962 ( .A(n44636), .B(n44634), .Z(n44630) );
  IV U53963 ( .A(n44635), .Z(n44636) );
  NAND U53964 ( .A(n44637), .B(n44638), .Z(n44612) );
  NAND U53965 ( .A(n44639), .B(n44640), .Z(n44638) );
  NANDN U53966 ( .A(n44641), .B(n44642), .Z(n44639) );
  NANDN U53967 ( .A(n44642), .B(n44641), .Z(n44637) );
  AND U53968 ( .A(n44643), .B(n44644), .Z(n44614) );
  NAND U53969 ( .A(n44645), .B(n44646), .Z(n44644) );
  OR U53970 ( .A(n44647), .B(n44648), .Z(n44645) );
  NANDN U53971 ( .A(n44649), .B(n44647), .Z(n44643) );
  NAND U53972 ( .A(n44650), .B(n44651), .Z(n44618) );
  NANDN U53973 ( .A(n44652), .B(n44653), .Z(n44651) );
  OR U53974 ( .A(n44654), .B(n44655), .Z(n44653) );
  NANDN U53975 ( .A(n44656), .B(n44654), .Z(n44650) );
  IV U53976 ( .A(n44655), .Z(n44656) );
  XNOR U53977 ( .A(n44626), .B(n44657), .Z(n44621) );
  XNOR U53978 ( .A(n44624), .B(n44627), .Z(n44657) );
  NAND U53979 ( .A(n44658), .B(n44659), .Z(n44627) );
  NAND U53980 ( .A(n44660), .B(n44661), .Z(n44659) );
  OR U53981 ( .A(n44662), .B(n44663), .Z(n44660) );
  NANDN U53982 ( .A(n44664), .B(n44662), .Z(n44658) );
  IV U53983 ( .A(n44663), .Z(n44664) );
  NAND U53984 ( .A(n44665), .B(n44666), .Z(n44624) );
  NAND U53985 ( .A(n44667), .B(n44668), .Z(n44666) );
  NANDN U53986 ( .A(n44669), .B(n44670), .Z(n44667) );
  NANDN U53987 ( .A(n44670), .B(n44669), .Z(n44665) );
  AND U53988 ( .A(n44671), .B(n44672), .Z(n44626) );
  NAND U53989 ( .A(n44673), .B(n44674), .Z(n44672) );
  OR U53990 ( .A(n44675), .B(n44676), .Z(n44673) );
  NANDN U53991 ( .A(n44677), .B(n44675), .Z(n44671) );
  XNOR U53992 ( .A(n44652), .B(n44678), .Z(N61438) );
  XOR U53993 ( .A(n44654), .B(n44655), .Z(n44678) );
  XNOR U53994 ( .A(n44668), .B(n44679), .Z(n44655) );
  XOR U53995 ( .A(n44669), .B(n44670), .Z(n44679) );
  XOR U53996 ( .A(n44675), .B(n44680), .Z(n44670) );
  XOR U53997 ( .A(n44674), .B(n44677), .Z(n44680) );
  IV U53998 ( .A(n44676), .Z(n44677) );
  NAND U53999 ( .A(n44681), .B(n44682), .Z(n44676) );
  OR U54000 ( .A(n44683), .B(n44684), .Z(n44682) );
  OR U54001 ( .A(n44685), .B(n44686), .Z(n44681) );
  NAND U54002 ( .A(n44687), .B(n44688), .Z(n44674) );
  OR U54003 ( .A(n44689), .B(n44690), .Z(n44688) );
  OR U54004 ( .A(n44691), .B(n44692), .Z(n44687) );
  NOR U54005 ( .A(n44693), .B(n44694), .Z(n44675) );
  ANDN U54006 ( .B(n44695), .A(n44696), .Z(n44669) );
  XNOR U54007 ( .A(n44662), .B(n44697), .Z(n44668) );
  XNOR U54008 ( .A(n44661), .B(n44663), .Z(n44697) );
  NAND U54009 ( .A(n44698), .B(n44699), .Z(n44663) );
  OR U54010 ( .A(n44700), .B(n44701), .Z(n44699) );
  OR U54011 ( .A(n44702), .B(n44703), .Z(n44698) );
  NAND U54012 ( .A(n44704), .B(n44705), .Z(n44661) );
  OR U54013 ( .A(n44706), .B(n44707), .Z(n44705) );
  OR U54014 ( .A(n44708), .B(n44709), .Z(n44704) );
  ANDN U54015 ( .B(n44710), .A(n44711), .Z(n44662) );
  IV U54016 ( .A(n44712), .Z(n44710) );
  ANDN U54017 ( .B(n44713), .A(n44714), .Z(n44654) );
  XOR U54018 ( .A(n44640), .B(n44715), .Z(n44652) );
  XOR U54019 ( .A(n44641), .B(n44642), .Z(n44715) );
  XOR U54020 ( .A(n44647), .B(n44716), .Z(n44642) );
  XOR U54021 ( .A(n44646), .B(n44649), .Z(n44716) );
  IV U54022 ( .A(n44648), .Z(n44649) );
  NAND U54023 ( .A(n44717), .B(n44718), .Z(n44648) );
  OR U54024 ( .A(n44719), .B(n44720), .Z(n44718) );
  OR U54025 ( .A(n44721), .B(n44722), .Z(n44717) );
  NAND U54026 ( .A(n44723), .B(n44724), .Z(n44646) );
  OR U54027 ( .A(n44725), .B(n44726), .Z(n44724) );
  OR U54028 ( .A(n44727), .B(n44728), .Z(n44723) );
  NOR U54029 ( .A(n44729), .B(n44730), .Z(n44647) );
  ANDN U54030 ( .B(n44731), .A(n44732), .Z(n44641) );
  IV U54031 ( .A(n44733), .Z(n44731) );
  XNOR U54032 ( .A(n44634), .B(n44734), .Z(n44640) );
  XNOR U54033 ( .A(n44633), .B(n44635), .Z(n44734) );
  NAND U54034 ( .A(n44735), .B(n44736), .Z(n44635) );
  OR U54035 ( .A(n44737), .B(n44738), .Z(n44736) );
  OR U54036 ( .A(n44739), .B(n44740), .Z(n44735) );
  NAND U54037 ( .A(n44741), .B(n44742), .Z(n44633) );
  OR U54038 ( .A(n44743), .B(n44744), .Z(n44742) );
  OR U54039 ( .A(n44745), .B(n44746), .Z(n44741) );
  ANDN U54040 ( .B(n44747), .A(n44748), .Z(n44634) );
  IV U54041 ( .A(n44749), .Z(n44747) );
  XNOR U54042 ( .A(n44714), .B(n44713), .Z(N61437) );
  XOR U54043 ( .A(n44733), .B(n44732), .Z(n44713) );
  XNOR U54044 ( .A(n44748), .B(n44749), .Z(n44732) );
  XNOR U54045 ( .A(n44743), .B(n44744), .Z(n44749) );
  XNOR U54046 ( .A(n44745), .B(n44746), .Z(n44744) );
  XNOR U54047 ( .A(y[1573]), .B(x[1573]), .Z(n44746) );
  XNOR U54048 ( .A(y[1574]), .B(x[1574]), .Z(n44745) );
  XNOR U54049 ( .A(y[1572]), .B(x[1572]), .Z(n44743) );
  XNOR U54050 ( .A(n44737), .B(n44738), .Z(n44748) );
  XNOR U54051 ( .A(y[1569]), .B(x[1569]), .Z(n44738) );
  XNOR U54052 ( .A(n44739), .B(n44740), .Z(n44737) );
  XNOR U54053 ( .A(y[1570]), .B(x[1570]), .Z(n44740) );
  XNOR U54054 ( .A(y[1571]), .B(x[1571]), .Z(n44739) );
  XNOR U54055 ( .A(n44730), .B(n44729), .Z(n44733) );
  XNOR U54056 ( .A(n44725), .B(n44726), .Z(n44729) );
  XNOR U54057 ( .A(y[1566]), .B(x[1566]), .Z(n44726) );
  XNOR U54058 ( .A(n44727), .B(n44728), .Z(n44725) );
  XNOR U54059 ( .A(y[1567]), .B(x[1567]), .Z(n44728) );
  XNOR U54060 ( .A(y[1568]), .B(x[1568]), .Z(n44727) );
  XNOR U54061 ( .A(n44719), .B(n44720), .Z(n44730) );
  XNOR U54062 ( .A(y[1563]), .B(x[1563]), .Z(n44720) );
  XNOR U54063 ( .A(n44721), .B(n44722), .Z(n44719) );
  XNOR U54064 ( .A(y[1564]), .B(x[1564]), .Z(n44722) );
  XNOR U54065 ( .A(y[1565]), .B(x[1565]), .Z(n44721) );
  XOR U54066 ( .A(n44695), .B(n44696), .Z(n44714) );
  XNOR U54067 ( .A(n44711), .B(n44712), .Z(n44696) );
  XNOR U54068 ( .A(n44706), .B(n44707), .Z(n44712) );
  XNOR U54069 ( .A(n44708), .B(n44709), .Z(n44707) );
  XNOR U54070 ( .A(y[1561]), .B(x[1561]), .Z(n44709) );
  XNOR U54071 ( .A(y[1562]), .B(x[1562]), .Z(n44708) );
  XNOR U54072 ( .A(y[1560]), .B(x[1560]), .Z(n44706) );
  XNOR U54073 ( .A(n44700), .B(n44701), .Z(n44711) );
  XNOR U54074 ( .A(y[1557]), .B(x[1557]), .Z(n44701) );
  XNOR U54075 ( .A(n44702), .B(n44703), .Z(n44700) );
  XNOR U54076 ( .A(y[1558]), .B(x[1558]), .Z(n44703) );
  XNOR U54077 ( .A(y[1559]), .B(x[1559]), .Z(n44702) );
  XOR U54078 ( .A(n44694), .B(n44693), .Z(n44695) );
  XNOR U54079 ( .A(n44689), .B(n44690), .Z(n44693) );
  XNOR U54080 ( .A(y[1554]), .B(x[1554]), .Z(n44690) );
  XNOR U54081 ( .A(n44691), .B(n44692), .Z(n44689) );
  XNOR U54082 ( .A(y[1555]), .B(x[1555]), .Z(n44692) );
  XNOR U54083 ( .A(y[1556]), .B(x[1556]), .Z(n44691) );
  XNOR U54084 ( .A(n44683), .B(n44684), .Z(n44694) );
  XNOR U54085 ( .A(y[1551]), .B(x[1551]), .Z(n44684) );
  XNOR U54086 ( .A(n44685), .B(n44686), .Z(n44683) );
  XNOR U54087 ( .A(y[1552]), .B(x[1552]), .Z(n44686) );
  XNOR U54088 ( .A(y[1553]), .B(x[1553]), .Z(n44685) );
  NAND U54089 ( .A(n44750), .B(n44751), .Z(N61428) );
  NANDN U54090 ( .A(n44752), .B(n44753), .Z(n44751) );
  OR U54091 ( .A(n44754), .B(n44755), .Z(n44753) );
  NAND U54092 ( .A(n44754), .B(n44755), .Z(n44750) );
  XOR U54093 ( .A(n44754), .B(n44756), .Z(N61427) );
  XNOR U54094 ( .A(n44752), .B(n44755), .Z(n44756) );
  AND U54095 ( .A(n44757), .B(n44758), .Z(n44755) );
  NANDN U54096 ( .A(n44759), .B(n44760), .Z(n44758) );
  NANDN U54097 ( .A(n44761), .B(n44762), .Z(n44760) );
  NANDN U54098 ( .A(n44762), .B(n44761), .Z(n44757) );
  NAND U54099 ( .A(n44763), .B(n44764), .Z(n44752) );
  NANDN U54100 ( .A(n44765), .B(n44766), .Z(n44764) );
  OR U54101 ( .A(n44767), .B(n44768), .Z(n44766) );
  NAND U54102 ( .A(n44768), .B(n44767), .Z(n44763) );
  AND U54103 ( .A(n44769), .B(n44770), .Z(n44754) );
  NANDN U54104 ( .A(n44771), .B(n44772), .Z(n44770) );
  NANDN U54105 ( .A(n44773), .B(n44774), .Z(n44772) );
  NANDN U54106 ( .A(n44774), .B(n44773), .Z(n44769) );
  XOR U54107 ( .A(n44768), .B(n44775), .Z(N61426) );
  XOR U54108 ( .A(n44765), .B(n44767), .Z(n44775) );
  XNOR U54109 ( .A(n44761), .B(n44776), .Z(n44767) );
  XNOR U54110 ( .A(n44759), .B(n44762), .Z(n44776) );
  NAND U54111 ( .A(n44777), .B(n44778), .Z(n44762) );
  NAND U54112 ( .A(n44779), .B(n44780), .Z(n44778) );
  OR U54113 ( .A(n44781), .B(n44782), .Z(n44779) );
  NANDN U54114 ( .A(n44783), .B(n44781), .Z(n44777) );
  IV U54115 ( .A(n44782), .Z(n44783) );
  NAND U54116 ( .A(n44784), .B(n44785), .Z(n44759) );
  NAND U54117 ( .A(n44786), .B(n44787), .Z(n44785) );
  NANDN U54118 ( .A(n44788), .B(n44789), .Z(n44786) );
  NANDN U54119 ( .A(n44789), .B(n44788), .Z(n44784) );
  AND U54120 ( .A(n44790), .B(n44791), .Z(n44761) );
  NAND U54121 ( .A(n44792), .B(n44793), .Z(n44791) );
  OR U54122 ( .A(n44794), .B(n44795), .Z(n44792) );
  NANDN U54123 ( .A(n44796), .B(n44794), .Z(n44790) );
  NAND U54124 ( .A(n44797), .B(n44798), .Z(n44765) );
  NANDN U54125 ( .A(n44799), .B(n44800), .Z(n44798) );
  OR U54126 ( .A(n44801), .B(n44802), .Z(n44800) );
  NANDN U54127 ( .A(n44803), .B(n44801), .Z(n44797) );
  IV U54128 ( .A(n44802), .Z(n44803) );
  XNOR U54129 ( .A(n44773), .B(n44804), .Z(n44768) );
  XNOR U54130 ( .A(n44771), .B(n44774), .Z(n44804) );
  NAND U54131 ( .A(n44805), .B(n44806), .Z(n44774) );
  NAND U54132 ( .A(n44807), .B(n44808), .Z(n44806) );
  OR U54133 ( .A(n44809), .B(n44810), .Z(n44807) );
  NANDN U54134 ( .A(n44811), .B(n44809), .Z(n44805) );
  IV U54135 ( .A(n44810), .Z(n44811) );
  NAND U54136 ( .A(n44812), .B(n44813), .Z(n44771) );
  NAND U54137 ( .A(n44814), .B(n44815), .Z(n44813) );
  NANDN U54138 ( .A(n44816), .B(n44817), .Z(n44814) );
  NANDN U54139 ( .A(n44817), .B(n44816), .Z(n44812) );
  AND U54140 ( .A(n44818), .B(n44819), .Z(n44773) );
  NAND U54141 ( .A(n44820), .B(n44821), .Z(n44819) );
  OR U54142 ( .A(n44822), .B(n44823), .Z(n44820) );
  NANDN U54143 ( .A(n44824), .B(n44822), .Z(n44818) );
  XNOR U54144 ( .A(n44799), .B(n44825), .Z(N61425) );
  XOR U54145 ( .A(n44801), .B(n44802), .Z(n44825) );
  XNOR U54146 ( .A(n44815), .B(n44826), .Z(n44802) );
  XOR U54147 ( .A(n44816), .B(n44817), .Z(n44826) );
  XOR U54148 ( .A(n44822), .B(n44827), .Z(n44817) );
  XOR U54149 ( .A(n44821), .B(n44824), .Z(n44827) );
  IV U54150 ( .A(n44823), .Z(n44824) );
  NAND U54151 ( .A(n44828), .B(n44829), .Z(n44823) );
  OR U54152 ( .A(n44830), .B(n44831), .Z(n44829) );
  OR U54153 ( .A(n44832), .B(n44833), .Z(n44828) );
  NAND U54154 ( .A(n44834), .B(n44835), .Z(n44821) );
  OR U54155 ( .A(n44836), .B(n44837), .Z(n44835) );
  OR U54156 ( .A(n44838), .B(n44839), .Z(n44834) );
  NOR U54157 ( .A(n44840), .B(n44841), .Z(n44822) );
  ANDN U54158 ( .B(n44842), .A(n44843), .Z(n44816) );
  XNOR U54159 ( .A(n44809), .B(n44844), .Z(n44815) );
  XNOR U54160 ( .A(n44808), .B(n44810), .Z(n44844) );
  NAND U54161 ( .A(n44845), .B(n44846), .Z(n44810) );
  OR U54162 ( .A(n44847), .B(n44848), .Z(n44846) );
  OR U54163 ( .A(n44849), .B(n44850), .Z(n44845) );
  NAND U54164 ( .A(n44851), .B(n44852), .Z(n44808) );
  OR U54165 ( .A(n44853), .B(n44854), .Z(n44852) );
  OR U54166 ( .A(n44855), .B(n44856), .Z(n44851) );
  ANDN U54167 ( .B(n44857), .A(n44858), .Z(n44809) );
  IV U54168 ( .A(n44859), .Z(n44857) );
  ANDN U54169 ( .B(n44860), .A(n44861), .Z(n44801) );
  XOR U54170 ( .A(n44787), .B(n44862), .Z(n44799) );
  XOR U54171 ( .A(n44788), .B(n44789), .Z(n44862) );
  XOR U54172 ( .A(n44794), .B(n44863), .Z(n44789) );
  XOR U54173 ( .A(n44793), .B(n44796), .Z(n44863) );
  IV U54174 ( .A(n44795), .Z(n44796) );
  NAND U54175 ( .A(n44864), .B(n44865), .Z(n44795) );
  OR U54176 ( .A(n44866), .B(n44867), .Z(n44865) );
  OR U54177 ( .A(n44868), .B(n44869), .Z(n44864) );
  NAND U54178 ( .A(n44870), .B(n44871), .Z(n44793) );
  OR U54179 ( .A(n44872), .B(n44873), .Z(n44871) );
  OR U54180 ( .A(n44874), .B(n44875), .Z(n44870) );
  NOR U54181 ( .A(n44876), .B(n44877), .Z(n44794) );
  ANDN U54182 ( .B(n44878), .A(n44879), .Z(n44788) );
  IV U54183 ( .A(n44880), .Z(n44878) );
  XNOR U54184 ( .A(n44781), .B(n44881), .Z(n44787) );
  XNOR U54185 ( .A(n44780), .B(n44782), .Z(n44881) );
  NAND U54186 ( .A(n44882), .B(n44883), .Z(n44782) );
  OR U54187 ( .A(n44884), .B(n44885), .Z(n44883) );
  OR U54188 ( .A(n44886), .B(n44887), .Z(n44882) );
  NAND U54189 ( .A(n44888), .B(n44889), .Z(n44780) );
  OR U54190 ( .A(n44890), .B(n44891), .Z(n44889) );
  OR U54191 ( .A(n44892), .B(n44893), .Z(n44888) );
  ANDN U54192 ( .B(n44894), .A(n44895), .Z(n44781) );
  IV U54193 ( .A(n44896), .Z(n44894) );
  XNOR U54194 ( .A(n44861), .B(n44860), .Z(N61424) );
  XOR U54195 ( .A(n44880), .B(n44879), .Z(n44860) );
  XNOR U54196 ( .A(n44895), .B(n44896), .Z(n44879) );
  XNOR U54197 ( .A(n44890), .B(n44891), .Z(n44896) );
  XNOR U54198 ( .A(n44892), .B(n44893), .Z(n44891) );
  XNOR U54199 ( .A(y[1549]), .B(x[1549]), .Z(n44893) );
  XNOR U54200 ( .A(y[1550]), .B(x[1550]), .Z(n44892) );
  XNOR U54201 ( .A(y[1548]), .B(x[1548]), .Z(n44890) );
  XNOR U54202 ( .A(n44884), .B(n44885), .Z(n44895) );
  XNOR U54203 ( .A(y[1545]), .B(x[1545]), .Z(n44885) );
  XNOR U54204 ( .A(n44886), .B(n44887), .Z(n44884) );
  XNOR U54205 ( .A(y[1546]), .B(x[1546]), .Z(n44887) );
  XNOR U54206 ( .A(y[1547]), .B(x[1547]), .Z(n44886) );
  XNOR U54207 ( .A(n44877), .B(n44876), .Z(n44880) );
  XNOR U54208 ( .A(n44872), .B(n44873), .Z(n44876) );
  XNOR U54209 ( .A(y[1542]), .B(x[1542]), .Z(n44873) );
  XNOR U54210 ( .A(n44874), .B(n44875), .Z(n44872) );
  XNOR U54211 ( .A(y[1543]), .B(x[1543]), .Z(n44875) );
  XNOR U54212 ( .A(y[1544]), .B(x[1544]), .Z(n44874) );
  XNOR U54213 ( .A(n44866), .B(n44867), .Z(n44877) );
  XNOR U54214 ( .A(y[1539]), .B(x[1539]), .Z(n44867) );
  XNOR U54215 ( .A(n44868), .B(n44869), .Z(n44866) );
  XNOR U54216 ( .A(y[1540]), .B(x[1540]), .Z(n44869) );
  XNOR U54217 ( .A(y[1541]), .B(x[1541]), .Z(n44868) );
  XOR U54218 ( .A(n44842), .B(n44843), .Z(n44861) );
  XNOR U54219 ( .A(n44858), .B(n44859), .Z(n44843) );
  XNOR U54220 ( .A(n44853), .B(n44854), .Z(n44859) );
  XNOR U54221 ( .A(n44855), .B(n44856), .Z(n44854) );
  XNOR U54222 ( .A(y[1537]), .B(x[1537]), .Z(n44856) );
  XNOR U54223 ( .A(y[1538]), .B(x[1538]), .Z(n44855) );
  XNOR U54224 ( .A(y[1536]), .B(x[1536]), .Z(n44853) );
  XNOR U54225 ( .A(n44847), .B(n44848), .Z(n44858) );
  XNOR U54226 ( .A(y[1533]), .B(x[1533]), .Z(n44848) );
  XNOR U54227 ( .A(n44849), .B(n44850), .Z(n44847) );
  XNOR U54228 ( .A(y[1534]), .B(x[1534]), .Z(n44850) );
  XNOR U54229 ( .A(y[1535]), .B(x[1535]), .Z(n44849) );
  XOR U54230 ( .A(n44841), .B(n44840), .Z(n44842) );
  XNOR U54231 ( .A(n44836), .B(n44837), .Z(n44840) );
  XNOR U54232 ( .A(y[1530]), .B(x[1530]), .Z(n44837) );
  XNOR U54233 ( .A(n44838), .B(n44839), .Z(n44836) );
  XNOR U54234 ( .A(y[1531]), .B(x[1531]), .Z(n44839) );
  XNOR U54235 ( .A(y[1532]), .B(x[1532]), .Z(n44838) );
  XNOR U54236 ( .A(n44830), .B(n44831), .Z(n44841) );
  XNOR U54237 ( .A(y[1527]), .B(x[1527]), .Z(n44831) );
  XNOR U54238 ( .A(n44832), .B(n44833), .Z(n44830) );
  XNOR U54239 ( .A(y[1528]), .B(x[1528]), .Z(n44833) );
  XNOR U54240 ( .A(y[1529]), .B(x[1529]), .Z(n44832) );
  NAND U54241 ( .A(n44897), .B(n44898), .Z(N61415) );
  NANDN U54242 ( .A(n44899), .B(n44900), .Z(n44898) );
  OR U54243 ( .A(n44901), .B(n44902), .Z(n44900) );
  NAND U54244 ( .A(n44901), .B(n44902), .Z(n44897) );
  XOR U54245 ( .A(n44901), .B(n44903), .Z(N61414) );
  XNOR U54246 ( .A(n44899), .B(n44902), .Z(n44903) );
  AND U54247 ( .A(n44904), .B(n44905), .Z(n44902) );
  NANDN U54248 ( .A(n44906), .B(n44907), .Z(n44905) );
  NANDN U54249 ( .A(n44908), .B(n44909), .Z(n44907) );
  NANDN U54250 ( .A(n44909), .B(n44908), .Z(n44904) );
  NAND U54251 ( .A(n44910), .B(n44911), .Z(n44899) );
  NANDN U54252 ( .A(n44912), .B(n44913), .Z(n44911) );
  OR U54253 ( .A(n44914), .B(n44915), .Z(n44913) );
  NAND U54254 ( .A(n44915), .B(n44914), .Z(n44910) );
  AND U54255 ( .A(n44916), .B(n44917), .Z(n44901) );
  NANDN U54256 ( .A(n44918), .B(n44919), .Z(n44917) );
  NANDN U54257 ( .A(n44920), .B(n44921), .Z(n44919) );
  NANDN U54258 ( .A(n44921), .B(n44920), .Z(n44916) );
  XOR U54259 ( .A(n44915), .B(n44922), .Z(N61413) );
  XOR U54260 ( .A(n44912), .B(n44914), .Z(n44922) );
  XNOR U54261 ( .A(n44908), .B(n44923), .Z(n44914) );
  XNOR U54262 ( .A(n44906), .B(n44909), .Z(n44923) );
  NAND U54263 ( .A(n44924), .B(n44925), .Z(n44909) );
  NAND U54264 ( .A(n44926), .B(n44927), .Z(n44925) );
  OR U54265 ( .A(n44928), .B(n44929), .Z(n44926) );
  NANDN U54266 ( .A(n44930), .B(n44928), .Z(n44924) );
  IV U54267 ( .A(n44929), .Z(n44930) );
  NAND U54268 ( .A(n44931), .B(n44932), .Z(n44906) );
  NAND U54269 ( .A(n44933), .B(n44934), .Z(n44932) );
  NANDN U54270 ( .A(n44935), .B(n44936), .Z(n44933) );
  NANDN U54271 ( .A(n44936), .B(n44935), .Z(n44931) );
  AND U54272 ( .A(n44937), .B(n44938), .Z(n44908) );
  NAND U54273 ( .A(n44939), .B(n44940), .Z(n44938) );
  OR U54274 ( .A(n44941), .B(n44942), .Z(n44939) );
  NANDN U54275 ( .A(n44943), .B(n44941), .Z(n44937) );
  NAND U54276 ( .A(n44944), .B(n44945), .Z(n44912) );
  NANDN U54277 ( .A(n44946), .B(n44947), .Z(n44945) );
  OR U54278 ( .A(n44948), .B(n44949), .Z(n44947) );
  NANDN U54279 ( .A(n44950), .B(n44948), .Z(n44944) );
  IV U54280 ( .A(n44949), .Z(n44950) );
  XNOR U54281 ( .A(n44920), .B(n44951), .Z(n44915) );
  XNOR U54282 ( .A(n44918), .B(n44921), .Z(n44951) );
  NAND U54283 ( .A(n44952), .B(n44953), .Z(n44921) );
  NAND U54284 ( .A(n44954), .B(n44955), .Z(n44953) );
  OR U54285 ( .A(n44956), .B(n44957), .Z(n44954) );
  NANDN U54286 ( .A(n44958), .B(n44956), .Z(n44952) );
  IV U54287 ( .A(n44957), .Z(n44958) );
  NAND U54288 ( .A(n44959), .B(n44960), .Z(n44918) );
  NAND U54289 ( .A(n44961), .B(n44962), .Z(n44960) );
  NANDN U54290 ( .A(n44963), .B(n44964), .Z(n44961) );
  NANDN U54291 ( .A(n44964), .B(n44963), .Z(n44959) );
  AND U54292 ( .A(n44965), .B(n44966), .Z(n44920) );
  NAND U54293 ( .A(n44967), .B(n44968), .Z(n44966) );
  OR U54294 ( .A(n44969), .B(n44970), .Z(n44967) );
  NANDN U54295 ( .A(n44971), .B(n44969), .Z(n44965) );
  XNOR U54296 ( .A(n44946), .B(n44972), .Z(N61412) );
  XOR U54297 ( .A(n44948), .B(n44949), .Z(n44972) );
  XNOR U54298 ( .A(n44962), .B(n44973), .Z(n44949) );
  XOR U54299 ( .A(n44963), .B(n44964), .Z(n44973) );
  XOR U54300 ( .A(n44969), .B(n44974), .Z(n44964) );
  XOR U54301 ( .A(n44968), .B(n44971), .Z(n44974) );
  IV U54302 ( .A(n44970), .Z(n44971) );
  NAND U54303 ( .A(n44975), .B(n44976), .Z(n44970) );
  OR U54304 ( .A(n44977), .B(n44978), .Z(n44976) );
  OR U54305 ( .A(n44979), .B(n44980), .Z(n44975) );
  NAND U54306 ( .A(n44981), .B(n44982), .Z(n44968) );
  OR U54307 ( .A(n44983), .B(n44984), .Z(n44982) );
  OR U54308 ( .A(n44985), .B(n44986), .Z(n44981) );
  NOR U54309 ( .A(n44987), .B(n44988), .Z(n44969) );
  ANDN U54310 ( .B(n44989), .A(n44990), .Z(n44963) );
  XNOR U54311 ( .A(n44956), .B(n44991), .Z(n44962) );
  XNOR U54312 ( .A(n44955), .B(n44957), .Z(n44991) );
  NAND U54313 ( .A(n44992), .B(n44993), .Z(n44957) );
  OR U54314 ( .A(n44994), .B(n44995), .Z(n44993) );
  OR U54315 ( .A(n44996), .B(n44997), .Z(n44992) );
  NAND U54316 ( .A(n44998), .B(n44999), .Z(n44955) );
  OR U54317 ( .A(n45000), .B(n45001), .Z(n44999) );
  OR U54318 ( .A(n45002), .B(n45003), .Z(n44998) );
  ANDN U54319 ( .B(n45004), .A(n45005), .Z(n44956) );
  IV U54320 ( .A(n45006), .Z(n45004) );
  ANDN U54321 ( .B(n45007), .A(n45008), .Z(n44948) );
  XOR U54322 ( .A(n44934), .B(n45009), .Z(n44946) );
  XOR U54323 ( .A(n44935), .B(n44936), .Z(n45009) );
  XOR U54324 ( .A(n44941), .B(n45010), .Z(n44936) );
  XOR U54325 ( .A(n44940), .B(n44943), .Z(n45010) );
  IV U54326 ( .A(n44942), .Z(n44943) );
  NAND U54327 ( .A(n45011), .B(n45012), .Z(n44942) );
  OR U54328 ( .A(n45013), .B(n45014), .Z(n45012) );
  OR U54329 ( .A(n45015), .B(n45016), .Z(n45011) );
  NAND U54330 ( .A(n45017), .B(n45018), .Z(n44940) );
  OR U54331 ( .A(n45019), .B(n45020), .Z(n45018) );
  OR U54332 ( .A(n45021), .B(n45022), .Z(n45017) );
  NOR U54333 ( .A(n45023), .B(n45024), .Z(n44941) );
  ANDN U54334 ( .B(n45025), .A(n45026), .Z(n44935) );
  IV U54335 ( .A(n45027), .Z(n45025) );
  XNOR U54336 ( .A(n44928), .B(n45028), .Z(n44934) );
  XNOR U54337 ( .A(n44927), .B(n44929), .Z(n45028) );
  NAND U54338 ( .A(n45029), .B(n45030), .Z(n44929) );
  OR U54339 ( .A(n45031), .B(n45032), .Z(n45030) );
  OR U54340 ( .A(n45033), .B(n45034), .Z(n45029) );
  NAND U54341 ( .A(n45035), .B(n45036), .Z(n44927) );
  OR U54342 ( .A(n45037), .B(n45038), .Z(n45036) );
  OR U54343 ( .A(n45039), .B(n45040), .Z(n45035) );
  ANDN U54344 ( .B(n45041), .A(n45042), .Z(n44928) );
  IV U54345 ( .A(n45043), .Z(n45041) );
  XNOR U54346 ( .A(n45008), .B(n45007), .Z(N61411) );
  XOR U54347 ( .A(n45027), .B(n45026), .Z(n45007) );
  XNOR U54348 ( .A(n45042), .B(n45043), .Z(n45026) );
  XNOR U54349 ( .A(n45037), .B(n45038), .Z(n45043) );
  XNOR U54350 ( .A(n45039), .B(n45040), .Z(n45038) );
  XNOR U54351 ( .A(y[1525]), .B(x[1525]), .Z(n45040) );
  XNOR U54352 ( .A(y[1526]), .B(x[1526]), .Z(n45039) );
  XNOR U54353 ( .A(y[1524]), .B(x[1524]), .Z(n45037) );
  XNOR U54354 ( .A(n45031), .B(n45032), .Z(n45042) );
  XNOR U54355 ( .A(y[1521]), .B(x[1521]), .Z(n45032) );
  XNOR U54356 ( .A(n45033), .B(n45034), .Z(n45031) );
  XNOR U54357 ( .A(y[1522]), .B(x[1522]), .Z(n45034) );
  XNOR U54358 ( .A(y[1523]), .B(x[1523]), .Z(n45033) );
  XNOR U54359 ( .A(n45024), .B(n45023), .Z(n45027) );
  XNOR U54360 ( .A(n45019), .B(n45020), .Z(n45023) );
  XNOR U54361 ( .A(y[1518]), .B(x[1518]), .Z(n45020) );
  XNOR U54362 ( .A(n45021), .B(n45022), .Z(n45019) );
  XNOR U54363 ( .A(y[1519]), .B(x[1519]), .Z(n45022) );
  XNOR U54364 ( .A(y[1520]), .B(x[1520]), .Z(n45021) );
  XNOR U54365 ( .A(n45013), .B(n45014), .Z(n45024) );
  XNOR U54366 ( .A(y[1515]), .B(x[1515]), .Z(n45014) );
  XNOR U54367 ( .A(n45015), .B(n45016), .Z(n45013) );
  XNOR U54368 ( .A(y[1516]), .B(x[1516]), .Z(n45016) );
  XNOR U54369 ( .A(y[1517]), .B(x[1517]), .Z(n45015) );
  XOR U54370 ( .A(n44989), .B(n44990), .Z(n45008) );
  XNOR U54371 ( .A(n45005), .B(n45006), .Z(n44990) );
  XNOR U54372 ( .A(n45000), .B(n45001), .Z(n45006) );
  XNOR U54373 ( .A(n45002), .B(n45003), .Z(n45001) );
  XNOR U54374 ( .A(y[1513]), .B(x[1513]), .Z(n45003) );
  XNOR U54375 ( .A(y[1514]), .B(x[1514]), .Z(n45002) );
  XNOR U54376 ( .A(y[1512]), .B(x[1512]), .Z(n45000) );
  XNOR U54377 ( .A(n44994), .B(n44995), .Z(n45005) );
  XNOR U54378 ( .A(y[1509]), .B(x[1509]), .Z(n44995) );
  XNOR U54379 ( .A(n44996), .B(n44997), .Z(n44994) );
  XNOR U54380 ( .A(y[1510]), .B(x[1510]), .Z(n44997) );
  XNOR U54381 ( .A(y[1511]), .B(x[1511]), .Z(n44996) );
  XOR U54382 ( .A(n44988), .B(n44987), .Z(n44989) );
  XNOR U54383 ( .A(n44983), .B(n44984), .Z(n44987) );
  XNOR U54384 ( .A(y[1506]), .B(x[1506]), .Z(n44984) );
  XNOR U54385 ( .A(n44985), .B(n44986), .Z(n44983) );
  XNOR U54386 ( .A(y[1507]), .B(x[1507]), .Z(n44986) );
  XNOR U54387 ( .A(y[1508]), .B(x[1508]), .Z(n44985) );
  XNOR U54388 ( .A(n44977), .B(n44978), .Z(n44988) );
  XNOR U54389 ( .A(y[1503]), .B(x[1503]), .Z(n44978) );
  XNOR U54390 ( .A(n44979), .B(n44980), .Z(n44977) );
  XNOR U54391 ( .A(y[1504]), .B(x[1504]), .Z(n44980) );
  XNOR U54392 ( .A(y[1505]), .B(x[1505]), .Z(n44979) );
  NAND U54393 ( .A(n45044), .B(n45045), .Z(N61402) );
  NANDN U54394 ( .A(n45046), .B(n45047), .Z(n45045) );
  OR U54395 ( .A(n45048), .B(n45049), .Z(n45047) );
  NAND U54396 ( .A(n45048), .B(n45049), .Z(n45044) );
  XOR U54397 ( .A(n45048), .B(n45050), .Z(N61401) );
  XNOR U54398 ( .A(n45046), .B(n45049), .Z(n45050) );
  AND U54399 ( .A(n45051), .B(n45052), .Z(n45049) );
  NANDN U54400 ( .A(n45053), .B(n45054), .Z(n45052) );
  NANDN U54401 ( .A(n45055), .B(n45056), .Z(n45054) );
  NANDN U54402 ( .A(n45056), .B(n45055), .Z(n45051) );
  NAND U54403 ( .A(n45057), .B(n45058), .Z(n45046) );
  NANDN U54404 ( .A(n45059), .B(n45060), .Z(n45058) );
  OR U54405 ( .A(n45061), .B(n45062), .Z(n45060) );
  NAND U54406 ( .A(n45062), .B(n45061), .Z(n45057) );
  AND U54407 ( .A(n45063), .B(n45064), .Z(n45048) );
  NANDN U54408 ( .A(n45065), .B(n45066), .Z(n45064) );
  NANDN U54409 ( .A(n45067), .B(n45068), .Z(n45066) );
  NANDN U54410 ( .A(n45068), .B(n45067), .Z(n45063) );
  XOR U54411 ( .A(n45062), .B(n45069), .Z(N61400) );
  XOR U54412 ( .A(n45059), .B(n45061), .Z(n45069) );
  XNOR U54413 ( .A(n45055), .B(n45070), .Z(n45061) );
  XNOR U54414 ( .A(n45053), .B(n45056), .Z(n45070) );
  NAND U54415 ( .A(n45071), .B(n45072), .Z(n45056) );
  NAND U54416 ( .A(n45073), .B(n45074), .Z(n45072) );
  OR U54417 ( .A(n45075), .B(n45076), .Z(n45073) );
  NANDN U54418 ( .A(n45077), .B(n45075), .Z(n45071) );
  IV U54419 ( .A(n45076), .Z(n45077) );
  NAND U54420 ( .A(n45078), .B(n45079), .Z(n45053) );
  NAND U54421 ( .A(n45080), .B(n45081), .Z(n45079) );
  NANDN U54422 ( .A(n45082), .B(n45083), .Z(n45080) );
  NANDN U54423 ( .A(n45083), .B(n45082), .Z(n45078) );
  AND U54424 ( .A(n45084), .B(n45085), .Z(n45055) );
  NAND U54425 ( .A(n45086), .B(n45087), .Z(n45085) );
  OR U54426 ( .A(n45088), .B(n45089), .Z(n45086) );
  NANDN U54427 ( .A(n45090), .B(n45088), .Z(n45084) );
  NAND U54428 ( .A(n45091), .B(n45092), .Z(n45059) );
  NANDN U54429 ( .A(n45093), .B(n45094), .Z(n45092) );
  OR U54430 ( .A(n45095), .B(n45096), .Z(n45094) );
  NANDN U54431 ( .A(n45097), .B(n45095), .Z(n45091) );
  IV U54432 ( .A(n45096), .Z(n45097) );
  XNOR U54433 ( .A(n45067), .B(n45098), .Z(n45062) );
  XNOR U54434 ( .A(n45065), .B(n45068), .Z(n45098) );
  NAND U54435 ( .A(n45099), .B(n45100), .Z(n45068) );
  NAND U54436 ( .A(n45101), .B(n45102), .Z(n45100) );
  OR U54437 ( .A(n45103), .B(n45104), .Z(n45101) );
  NANDN U54438 ( .A(n45105), .B(n45103), .Z(n45099) );
  IV U54439 ( .A(n45104), .Z(n45105) );
  NAND U54440 ( .A(n45106), .B(n45107), .Z(n45065) );
  NAND U54441 ( .A(n45108), .B(n45109), .Z(n45107) );
  NANDN U54442 ( .A(n45110), .B(n45111), .Z(n45108) );
  NANDN U54443 ( .A(n45111), .B(n45110), .Z(n45106) );
  AND U54444 ( .A(n45112), .B(n45113), .Z(n45067) );
  NAND U54445 ( .A(n45114), .B(n45115), .Z(n45113) );
  OR U54446 ( .A(n45116), .B(n45117), .Z(n45114) );
  NANDN U54447 ( .A(n45118), .B(n45116), .Z(n45112) );
  XNOR U54448 ( .A(n45093), .B(n45119), .Z(N61399) );
  XOR U54449 ( .A(n45095), .B(n45096), .Z(n45119) );
  XNOR U54450 ( .A(n45109), .B(n45120), .Z(n45096) );
  XOR U54451 ( .A(n45110), .B(n45111), .Z(n45120) );
  XOR U54452 ( .A(n45116), .B(n45121), .Z(n45111) );
  XOR U54453 ( .A(n45115), .B(n45118), .Z(n45121) );
  IV U54454 ( .A(n45117), .Z(n45118) );
  NAND U54455 ( .A(n45122), .B(n45123), .Z(n45117) );
  OR U54456 ( .A(n45124), .B(n45125), .Z(n45123) );
  OR U54457 ( .A(n45126), .B(n45127), .Z(n45122) );
  NAND U54458 ( .A(n45128), .B(n45129), .Z(n45115) );
  OR U54459 ( .A(n45130), .B(n45131), .Z(n45129) );
  OR U54460 ( .A(n45132), .B(n45133), .Z(n45128) );
  NOR U54461 ( .A(n45134), .B(n45135), .Z(n45116) );
  ANDN U54462 ( .B(n45136), .A(n45137), .Z(n45110) );
  XNOR U54463 ( .A(n45103), .B(n45138), .Z(n45109) );
  XNOR U54464 ( .A(n45102), .B(n45104), .Z(n45138) );
  NAND U54465 ( .A(n45139), .B(n45140), .Z(n45104) );
  OR U54466 ( .A(n45141), .B(n45142), .Z(n45140) );
  OR U54467 ( .A(n45143), .B(n45144), .Z(n45139) );
  NAND U54468 ( .A(n45145), .B(n45146), .Z(n45102) );
  OR U54469 ( .A(n45147), .B(n45148), .Z(n45146) );
  OR U54470 ( .A(n45149), .B(n45150), .Z(n45145) );
  ANDN U54471 ( .B(n45151), .A(n45152), .Z(n45103) );
  IV U54472 ( .A(n45153), .Z(n45151) );
  ANDN U54473 ( .B(n45154), .A(n45155), .Z(n45095) );
  XOR U54474 ( .A(n45081), .B(n45156), .Z(n45093) );
  XOR U54475 ( .A(n45082), .B(n45083), .Z(n45156) );
  XOR U54476 ( .A(n45088), .B(n45157), .Z(n45083) );
  XOR U54477 ( .A(n45087), .B(n45090), .Z(n45157) );
  IV U54478 ( .A(n45089), .Z(n45090) );
  NAND U54479 ( .A(n45158), .B(n45159), .Z(n45089) );
  OR U54480 ( .A(n45160), .B(n45161), .Z(n45159) );
  OR U54481 ( .A(n45162), .B(n45163), .Z(n45158) );
  NAND U54482 ( .A(n45164), .B(n45165), .Z(n45087) );
  OR U54483 ( .A(n45166), .B(n45167), .Z(n45165) );
  OR U54484 ( .A(n45168), .B(n45169), .Z(n45164) );
  NOR U54485 ( .A(n45170), .B(n45171), .Z(n45088) );
  ANDN U54486 ( .B(n45172), .A(n45173), .Z(n45082) );
  IV U54487 ( .A(n45174), .Z(n45172) );
  XNOR U54488 ( .A(n45075), .B(n45175), .Z(n45081) );
  XNOR U54489 ( .A(n45074), .B(n45076), .Z(n45175) );
  NAND U54490 ( .A(n45176), .B(n45177), .Z(n45076) );
  OR U54491 ( .A(n45178), .B(n45179), .Z(n45177) );
  OR U54492 ( .A(n45180), .B(n45181), .Z(n45176) );
  NAND U54493 ( .A(n45182), .B(n45183), .Z(n45074) );
  OR U54494 ( .A(n45184), .B(n45185), .Z(n45183) );
  OR U54495 ( .A(n45186), .B(n45187), .Z(n45182) );
  ANDN U54496 ( .B(n45188), .A(n45189), .Z(n45075) );
  IV U54497 ( .A(n45190), .Z(n45188) );
  XNOR U54498 ( .A(n45155), .B(n45154), .Z(N61398) );
  XOR U54499 ( .A(n45174), .B(n45173), .Z(n45154) );
  XNOR U54500 ( .A(n45189), .B(n45190), .Z(n45173) );
  XNOR U54501 ( .A(n45184), .B(n45185), .Z(n45190) );
  XNOR U54502 ( .A(n45186), .B(n45187), .Z(n45185) );
  XNOR U54503 ( .A(y[1501]), .B(x[1501]), .Z(n45187) );
  XNOR U54504 ( .A(y[1502]), .B(x[1502]), .Z(n45186) );
  XNOR U54505 ( .A(y[1500]), .B(x[1500]), .Z(n45184) );
  XNOR U54506 ( .A(n45178), .B(n45179), .Z(n45189) );
  XNOR U54507 ( .A(y[1497]), .B(x[1497]), .Z(n45179) );
  XNOR U54508 ( .A(n45180), .B(n45181), .Z(n45178) );
  XNOR U54509 ( .A(y[1498]), .B(x[1498]), .Z(n45181) );
  XNOR U54510 ( .A(y[1499]), .B(x[1499]), .Z(n45180) );
  XNOR U54511 ( .A(n45171), .B(n45170), .Z(n45174) );
  XNOR U54512 ( .A(n45166), .B(n45167), .Z(n45170) );
  XNOR U54513 ( .A(y[1494]), .B(x[1494]), .Z(n45167) );
  XNOR U54514 ( .A(n45168), .B(n45169), .Z(n45166) );
  XNOR U54515 ( .A(y[1495]), .B(x[1495]), .Z(n45169) );
  XNOR U54516 ( .A(y[1496]), .B(x[1496]), .Z(n45168) );
  XNOR U54517 ( .A(n45160), .B(n45161), .Z(n45171) );
  XNOR U54518 ( .A(y[1491]), .B(x[1491]), .Z(n45161) );
  XNOR U54519 ( .A(n45162), .B(n45163), .Z(n45160) );
  XNOR U54520 ( .A(y[1492]), .B(x[1492]), .Z(n45163) );
  XNOR U54521 ( .A(y[1493]), .B(x[1493]), .Z(n45162) );
  XOR U54522 ( .A(n45136), .B(n45137), .Z(n45155) );
  XNOR U54523 ( .A(n45152), .B(n45153), .Z(n45137) );
  XNOR U54524 ( .A(n45147), .B(n45148), .Z(n45153) );
  XNOR U54525 ( .A(n45149), .B(n45150), .Z(n45148) );
  XNOR U54526 ( .A(y[1489]), .B(x[1489]), .Z(n45150) );
  XNOR U54527 ( .A(y[1490]), .B(x[1490]), .Z(n45149) );
  XNOR U54528 ( .A(y[1488]), .B(x[1488]), .Z(n45147) );
  XNOR U54529 ( .A(n45141), .B(n45142), .Z(n45152) );
  XNOR U54530 ( .A(y[1485]), .B(x[1485]), .Z(n45142) );
  XNOR U54531 ( .A(n45143), .B(n45144), .Z(n45141) );
  XNOR U54532 ( .A(y[1486]), .B(x[1486]), .Z(n45144) );
  XNOR U54533 ( .A(y[1487]), .B(x[1487]), .Z(n45143) );
  XOR U54534 ( .A(n45135), .B(n45134), .Z(n45136) );
  XNOR U54535 ( .A(n45130), .B(n45131), .Z(n45134) );
  XNOR U54536 ( .A(y[1482]), .B(x[1482]), .Z(n45131) );
  XNOR U54537 ( .A(n45132), .B(n45133), .Z(n45130) );
  XNOR U54538 ( .A(y[1483]), .B(x[1483]), .Z(n45133) );
  XNOR U54539 ( .A(y[1484]), .B(x[1484]), .Z(n45132) );
  XNOR U54540 ( .A(n45124), .B(n45125), .Z(n45135) );
  XNOR U54541 ( .A(y[1479]), .B(x[1479]), .Z(n45125) );
  XNOR U54542 ( .A(n45126), .B(n45127), .Z(n45124) );
  XNOR U54543 ( .A(y[1480]), .B(x[1480]), .Z(n45127) );
  XNOR U54544 ( .A(y[1481]), .B(x[1481]), .Z(n45126) );
  NAND U54545 ( .A(n45191), .B(n45192), .Z(N61389) );
  NANDN U54546 ( .A(n45193), .B(n45194), .Z(n45192) );
  OR U54547 ( .A(n45195), .B(n45196), .Z(n45194) );
  NAND U54548 ( .A(n45195), .B(n45196), .Z(n45191) );
  XOR U54549 ( .A(n45195), .B(n45197), .Z(N61388) );
  XNOR U54550 ( .A(n45193), .B(n45196), .Z(n45197) );
  AND U54551 ( .A(n45198), .B(n45199), .Z(n45196) );
  NANDN U54552 ( .A(n45200), .B(n45201), .Z(n45199) );
  NANDN U54553 ( .A(n45202), .B(n45203), .Z(n45201) );
  NANDN U54554 ( .A(n45203), .B(n45202), .Z(n45198) );
  NAND U54555 ( .A(n45204), .B(n45205), .Z(n45193) );
  NANDN U54556 ( .A(n45206), .B(n45207), .Z(n45205) );
  OR U54557 ( .A(n45208), .B(n45209), .Z(n45207) );
  NAND U54558 ( .A(n45209), .B(n45208), .Z(n45204) );
  AND U54559 ( .A(n45210), .B(n45211), .Z(n45195) );
  NANDN U54560 ( .A(n45212), .B(n45213), .Z(n45211) );
  NANDN U54561 ( .A(n45214), .B(n45215), .Z(n45213) );
  NANDN U54562 ( .A(n45215), .B(n45214), .Z(n45210) );
  XOR U54563 ( .A(n45209), .B(n45216), .Z(N61387) );
  XOR U54564 ( .A(n45206), .B(n45208), .Z(n45216) );
  XNOR U54565 ( .A(n45202), .B(n45217), .Z(n45208) );
  XNOR U54566 ( .A(n45200), .B(n45203), .Z(n45217) );
  NAND U54567 ( .A(n45218), .B(n45219), .Z(n45203) );
  NAND U54568 ( .A(n45220), .B(n45221), .Z(n45219) );
  OR U54569 ( .A(n45222), .B(n45223), .Z(n45220) );
  NANDN U54570 ( .A(n45224), .B(n45222), .Z(n45218) );
  IV U54571 ( .A(n45223), .Z(n45224) );
  NAND U54572 ( .A(n45225), .B(n45226), .Z(n45200) );
  NAND U54573 ( .A(n45227), .B(n45228), .Z(n45226) );
  NANDN U54574 ( .A(n45229), .B(n45230), .Z(n45227) );
  NANDN U54575 ( .A(n45230), .B(n45229), .Z(n45225) );
  AND U54576 ( .A(n45231), .B(n45232), .Z(n45202) );
  NAND U54577 ( .A(n45233), .B(n45234), .Z(n45232) );
  OR U54578 ( .A(n45235), .B(n45236), .Z(n45233) );
  NANDN U54579 ( .A(n45237), .B(n45235), .Z(n45231) );
  NAND U54580 ( .A(n45238), .B(n45239), .Z(n45206) );
  NANDN U54581 ( .A(n45240), .B(n45241), .Z(n45239) );
  OR U54582 ( .A(n45242), .B(n45243), .Z(n45241) );
  NANDN U54583 ( .A(n45244), .B(n45242), .Z(n45238) );
  IV U54584 ( .A(n45243), .Z(n45244) );
  XNOR U54585 ( .A(n45214), .B(n45245), .Z(n45209) );
  XNOR U54586 ( .A(n45212), .B(n45215), .Z(n45245) );
  NAND U54587 ( .A(n45246), .B(n45247), .Z(n45215) );
  NAND U54588 ( .A(n45248), .B(n45249), .Z(n45247) );
  OR U54589 ( .A(n45250), .B(n45251), .Z(n45248) );
  NANDN U54590 ( .A(n45252), .B(n45250), .Z(n45246) );
  IV U54591 ( .A(n45251), .Z(n45252) );
  NAND U54592 ( .A(n45253), .B(n45254), .Z(n45212) );
  NAND U54593 ( .A(n45255), .B(n45256), .Z(n45254) );
  NANDN U54594 ( .A(n45257), .B(n45258), .Z(n45255) );
  NANDN U54595 ( .A(n45258), .B(n45257), .Z(n45253) );
  AND U54596 ( .A(n45259), .B(n45260), .Z(n45214) );
  NAND U54597 ( .A(n45261), .B(n45262), .Z(n45260) );
  OR U54598 ( .A(n45263), .B(n45264), .Z(n45261) );
  NANDN U54599 ( .A(n45265), .B(n45263), .Z(n45259) );
  XNOR U54600 ( .A(n45240), .B(n45266), .Z(N61386) );
  XOR U54601 ( .A(n45242), .B(n45243), .Z(n45266) );
  XNOR U54602 ( .A(n45256), .B(n45267), .Z(n45243) );
  XOR U54603 ( .A(n45257), .B(n45258), .Z(n45267) );
  XOR U54604 ( .A(n45263), .B(n45268), .Z(n45258) );
  XOR U54605 ( .A(n45262), .B(n45265), .Z(n45268) );
  IV U54606 ( .A(n45264), .Z(n45265) );
  NAND U54607 ( .A(n45269), .B(n45270), .Z(n45264) );
  OR U54608 ( .A(n45271), .B(n45272), .Z(n45270) );
  OR U54609 ( .A(n45273), .B(n45274), .Z(n45269) );
  NAND U54610 ( .A(n45275), .B(n45276), .Z(n45262) );
  OR U54611 ( .A(n45277), .B(n45278), .Z(n45276) );
  OR U54612 ( .A(n45279), .B(n45280), .Z(n45275) );
  NOR U54613 ( .A(n45281), .B(n45282), .Z(n45263) );
  ANDN U54614 ( .B(n45283), .A(n45284), .Z(n45257) );
  XNOR U54615 ( .A(n45250), .B(n45285), .Z(n45256) );
  XNOR U54616 ( .A(n45249), .B(n45251), .Z(n45285) );
  NAND U54617 ( .A(n45286), .B(n45287), .Z(n45251) );
  OR U54618 ( .A(n45288), .B(n45289), .Z(n45287) );
  OR U54619 ( .A(n45290), .B(n45291), .Z(n45286) );
  NAND U54620 ( .A(n45292), .B(n45293), .Z(n45249) );
  OR U54621 ( .A(n45294), .B(n45295), .Z(n45293) );
  OR U54622 ( .A(n45296), .B(n45297), .Z(n45292) );
  ANDN U54623 ( .B(n45298), .A(n45299), .Z(n45250) );
  IV U54624 ( .A(n45300), .Z(n45298) );
  ANDN U54625 ( .B(n45301), .A(n45302), .Z(n45242) );
  XOR U54626 ( .A(n45228), .B(n45303), .Z(n45240) );
  XOR U54627 ( .A(n45229), .B(n45230), .Z(n45303) );
  XOR U54628 ( .A(n45235), .B(n45304), .Z(n45230) );
  XOR U54629 ( .A(n45234), .B(n45237), .Z(n45304) );
  IV U54630 ( .A(n45236), .Z(n45237) );
  NAND U54631 ( .A(n45305), .B(n45306), .Z(n45236) );
  OR U54632 ( .A(n45307), .B(n45308), .Z(n45306) );
  OR U54633 ( .A(n45309), .B(n45310), .Z(n45305) );
  NAND U54634 ( .A(n45311), .B(n45312), .Z(n45234) );
  OR U54635 ( .A(n45313), .B(n45314), .Z(n45312) );
  OR U54636 ( .A(n45315), .B(n45316), .Z(n45311) );
  NOR U54637 ( .A(n45317), .B(n45318), .Z(n45235) );
  ANDN U54638 ( .B(n45319), .A(n45320), .Z(n45229) );
  IV U54639 ( .A(n45321), .Z(n45319) );
  XNOR U54640 ( .A(n45222), .B(n45322), .Z(n45228) );
  XNOR U54641 ( .A(n45221), .B(n45223), .Z(n45322) );
  NAND U54642 ( .A(n45323), .B(n45324), .Z(n45223) );
  OR U54643 ( .A(n45325), .B(n45326), .Z(n45324) );
  OR U54644 ( .A(n45327), .B(n45328), .Z(n45323) );
  NAND U54645 ( .A(n45329), .B(n45330), .Z(n45221) );
  OR U54646 ( .A(n45331), .B(n45332), .Z(n45330) );
  OR U54647 ( .A(n45333), .B(n45334), .Z(n45329) );
  ANDN U54648 ( .B(n45335), .A(n45336), .Z(n45222) );
  IV U54649 ( .A(n45337), .Z(n45335) );
  XNOR U54650 ( .A(n45302), .B(n45301), .Z(N61385) );
  XOR U54651 ( .A(n45321), .B(n45320), .Z(n45301) );
  XNOR U54652 ( .A(n45336), .B(n45337), .Z(n45320) );
  XNOR U54653 ( .A(n45331), .B(n45332), .Z(n45337) );
  XNOR U54654 ( .A(n45333), .B(n45334), .Z(n45332) );
  XNOR U54655 ( .A(y[1477]), .B(x[1477]), .Z(n45334) );
  XNOR U54656 ( .A(y[1478]), .B(x[1478]), .Z(n45333) );
  XNOR U54657 ( .A(y[1476]), .B(x[1476]), .Z(n45331) );
  XNOR U54658 ( .A(n45325), .B(n45326), .Z(n45336) );
  XNOR U54659 ( .A(y[1473]), .B(x[1473]), .Z(n45326) );
  XNOR U54660 ( .A(n45327), .B(n45328), .Z(n45325) );
  XNOR U54661 ( .A(y[1474]), .B(x[1474]), .Z(n45328) );
  XNOR U54662 ( .A(y[1475]), .B(x[1475]), .Z(n45327) );
  XNOR U54663 ( .A(n45318), .B(n45317), .Z(n45321) );
  XNOR U54664 ( .A(n45313), .B(n45314), .Z(n45317) );
  XNOR U54665 ( .A(y[1470]), .B(x[1470]), .Z(n45314) );
  XNOR U54666 ( .A(n45315), .B(n45316), .Z(n45313) );
  XNOR U54667 ( .A(y[1471]), .B(x[1471]), .Z(n45316) );
  XNOR U54668 ( .A(y[1472]), .B(x[1472]), .Z(n45315) );
  XNOR U54669 ( .A(n45307), .B(n45308), .Z(n45318) );
  XNOR U54670 ( .A(y[1467]), .B(x[1467]), .Z(n45308) );
  XNOR U54671 ( .A(n45309), .B(n45310), .Z(n45307) );
  XNOR U54672 ( .A(y[1468]), .B(x[1468]), .Z(n45310) );
  XNOR U54673 ( .A(y[1469]), .B(x[1469]), .Z(n45309) );
  XOR U54674 ( .A(n45283), .B(n45284), .Z(n45302) );
  XNOR U54675 ( .A(n45299), .B(n45300), .Z(n45284) );
  XNOR U54676 ( .A(n45294), .B(n45295), .Z(n45300) );
  XNOR U54677 ( .A(n45296), .B(n45297), .Z(n45295) );
  XNOR U54678 ( .A(y[1465]), .B(x[1465]), .Z(n45297) );
  XNOR U54679 ( .A(y[1466]), .B(x[1466]), .Z(n45296) );
  XNOR U54680 ( .A(y[1464]), .B(x[1464]), .Z(n45294) );
  XNOR U54681 ( .A(n45288), .B(n45289), .Z(n45299) );
  XNOR U54682 ( .A(y[1461]), .B(x[1461]), .Z(n45289) );
  XNOR U54683 ( .A(n45290), .B(n45291), .Z(n45288) );
  XNOR U54684 ( .A(y[1462]), .B(x[1462]), .Z(n45291) );
  XNOR U54685 ( .A(y[1463]), .B(x[1463]), .Z(n45290) );
  XOR U54686 ( .A(n45282), .B(n45281), .Z(n45283) );
  XNOR U54687 ( .A(n45277), .B(n45278), .Z(n45281) );
  XNOR U54688 ( .A(y[1458]), .B(x[1458]), .Z(n45278) );
  XNOR U54689 ( .A(n45279), .B(n45280), .Z(n45277) );
  XNOR U54690 ( .A(y[1459]), .B(x[1459]), .Z(n45280) );
  XNOR U54691 ( .A(y[1460]), .B(x[1460]), .Z(n45279) );
  XNOR U54692 ( .A(n45271), .B(n45272), .Z(n45282) );
  XNOR U54693 ( .A(y[1455]), .B(x[1455]), .Z(n45272) );
  XNOR U54694 ( .A(n45273), .B(n45274), .Z(n45271) );
  XNOR U54695 ( .A(y[1456]), .B(x[1456]), .Z(n45274) );
  XNOR U54696 ( .A(y[1457]), .B(x[1457]), .Z(n45273) );
  NAND U54697 ( .A(n45338), .B(n45339), .Z(N61376) );
  NANDN U54698 ( .A(n45340), .B(n45341), .Z(n45339) );
  OR U54699 ( .A(n45342), .B(n45343), .Z(n45341) );
  NAND U54700 ( .A(n45342), .B(n45343), .Z(n45338) );
  XOR U54701 ( .A(n45342), .B(n45344), .Z(N61375) );
  XNOR U54702 ( .A(n45340), .B(n45343), .Z(n45344) );
  AND U54703 ( .A(n45345), .B(n45346), .Z(n45343) );
  NANDN U54704 ( .A(n45347), .B(n45348), .Z(n45346) );
  NANDN U54705 ( .A(n45349), .B(n45350), .Z(n45348) );
  NANDN U54706 ( .A(n45350), .B(n45349), .Z(n45345) );
  NAND U54707 ( .A(n45351), .B(n45352), .Z(n45340) );
  NANDN U54708 ( .A(n45353), .B(n45354), .Z(n45352) );
  OR U54709 ( .A(n45355), .B(n45356), .Z(n45354) );
  NAND U54710 ( .A(n45356), .B(n45355), .Z(n45351) );
  AND U54711 ( .A(n45357), .B(n45358), .Z(n45342) );
  NANDN U54712 ( .A(n45359), .B(n45360), .Z(n45358) );
  NANDN U54713 ( .A(n45361), .B(n45362), .Z(n45360) );
  NANDN U54714 ( .A(n45362), .B(n45361), .Z(n45357) );
  XOR U54715 ( .A(n45356), .B(n45363), .Z(N61374) );
  XOR U54716 ( .A(n45353), .B(n45355), .Z(n45363) );
  XNOR U54717 ( .A(n45349), .B(n45364), .Z(n45355) );
  XNOR U54718 ( .A(n45347), .B(n45350), .Z(n45364) );
  NAND U54719 ( .A(n45365), .B(n45366), .Z(n45350) );
  NAND U54720 ( .A(n45367), .B(n45368), .Z(n45366) );
  OR U54721 ( .A(n45369), .B(n45370), .Z(n45367) );
  NANDN U54722 ( .A(n45371), .B(n45369), .Z(n45365) );
  IV U54723 ( .A(n45370), .Z(n45371) );
  NAND U54724 ( .A(n45372), .B(n45373), .Z(n45347) );
  NAND U54725 ( .A(n45374), .B(n45375), .Z(n45373) );
  NANDN U54726 ( .A(n45376), .B(n45377), .Z(n45374) );
  NANDN U54727 ( .A(n45377), .B(n45376), .Z(n45372) );
  AND U54728 ( .A(n45378), .B(n45379), .Z(n45349) );
  NAND U54729 ( .A(n45380), .B(n45381), .Z(n45379) );
  OR U54730 ( .A(n45382), .B(n45383), .Z(n45380) );
  NANDN U54731 ( .A(n45384), .B(n45382), .Z(n45378) );
  NAND U54732 ( .A(n45385), .B(n45386), .Z(n45353) );
  NANDN U54733 ( .A(n45387), .B(n45388), .Z(n45386) );
  OR U54734 ( .A(n45389), .B(n45390), .Z(n45388) );
  NANDN U54735 ( .A(n45391), .B(n45389), .Z(n45385) );
  IV U54736 ( .A(n45390), .Z(n45391) );
  XNOR U54737 ( .A(n45361), .B(n45392), .Z(n45356) );
  XNOR U54738 ( .A(n45359), .B(n45362), .Z(n45392) );
  NAND U54739 ( .A(n45393), .B(n45394), .Z(n45362) );
  NAND U54740 ( .A(n45395), .B(n45396), .Z(n45394) );
  OR U54741 ( .A(n45397), .B(n45398), .Z(n45395) );
  NANDN U54742 ( .A(n45399), .B(n45397), .Z(n45393) );
  IV U54743 ( .A(n45398), .Z(n45399) );
  NAND U54744 ( .A(n45400), .B(n45401), .Z(n45359) );
  NAND U54745 ( .A(n45402), .B(n45403), .Z(n45401) );
  NANDN U54746 ( .A(n45404), .B(n45405), .Z(n45402) );
  NANDN U54747 ( .A(n45405), .B(n45404), .Z(n45400) );
  AND U54748 ( .A(n45406), .B(n45407), .Z(n45361) );
  NAND U54749 ( .A(n45408), .B(n45409), .Z(n45407) );
  OR U54750 ( .A(n45410), .B(n45411), .Z(n45408) );
  NANDN U54751 ( .A(n45412), .B(n45410), .Z(n45406) );
  XNOR U54752 ( .A(n45387), .B(n45413), .Z(N61373) );
  XOR U54753 ( .A(n45389), .B(n45390), .Z(n45413) );
  XNOR U54754 ( .A(n45403), .B(n45414), .Z(n45390) );
  XOR U54755 ( .A(n45404), .B(n45405), .Z(n45414) );
  XOR U54756 ( .A(n45410), .B(n45415), .Z(n45405) );
  XOR U54757 ( .A(n45409), .B(n45412), .Z(n45415) );
  IV U54758 ( .A(n45411), .Z(n45412) );
  NAND U54759 ( .A(n45416), .B(n45417), .Z(n45411) );
  OR U54760 ( .A(n45418), .B(n45419), .Z(n45417) );
  OR U54761 ( .A(n45420), .B(n45421), .Z(n45416) );
  NAND U54762 ( .A(n45422), .B(n45423), .Z(n45409) );
  OR U54763 ( .A(n45424), .B(n45425), .Z(n45423) );
  OR U54764 ( .A(n45426), .B(n45427), .Z(n45422) );
  NOR U54765 ( .A(n45428), .B(n45429), .Z(n45410) );
  ANDN U54766 ( .B(n45430), .A(n45431), .Z(n45404) );
  XNOR U54767 ( .A(n45397), .B(n45432), .Z(n45403) );
  XNOR U54768 ( .A(n45396), .B(n45398), .Z(n45432) );
  NAND U54769 ( .A(n45433), .B(n45434), .Z(n45398) );
  OR U54770 ( .A(n45435), .B(n45436), .Z(n45434) );
  OR U54771 ( .A(n45437), .B(n45438), .Z(n45433) );
  NAND U54772 ( .A(n45439), .B(n45440), .Z(n45396) );
  OR U54773 ( .A(n45441), .B(n45442), .Z(n45440) );
  OR U54774 ( .A(n45443), .B(n45444), .Z(n45439) );
  ANDN U54775 ( .B(n45445), .A(n45446), .Z(n45397) );
  IV U54776 ( .A(n45447), .Z(n45445) );
  ANDN U54777 ( .B(n45448), .A(n45449), .Z(n45389) );
  XOR U54778 ( .A(n45375), .B(n45450), .Z(n45387) );
  XOR U54779 ( .A(n45376), .B(n45377), .Z(n45450) );
  XOR U54780 ( .A(n45382), .B(n45451), .Z(n45377) );
  XOR U54781 ( .A(n45381), .B(n45384), .Z(n45451) );
  IV U54782 ( .A(n45383), .Z(n45384) );
  NAND U54783 ( .A(n45452), .B(n45453), .Z(n45383) );
  OR U54784 ( .A(n45454), .B(n45455), .Z(n45453) );
  OR U54785 ( .A(n45456), .B(n45457), .Z(n45452) );
  NAND U54786 ( .A(n45458), .B(n45459), .Z(n45381) );
  OR U54787 ( .A(n45460), .B(n45461), .Z(n45459) );
  OR U54788 ( .A(n45462), .B(n45463), .Z(n45458) );
  NOR U54789 ( .A(n45464), .B(n45465), .Z(n45382) );
  ANDN U54790 ( .B(n45466), .A(n45467), .Z(n45376) );
  IV U54791 ( .A(n45468), .Z(n45466) );
  XNOR U54792 ( .A(n45369), .B(n45469), .Z(n45375) );
  XNOR U54793 ( .A(n45368), .B(n45370), .Z(n45469) );
  NAND U54794 ( .A(n45470), .B(n45471), .Z(n45370) );
  OR U54795 ( .A(n45472), .B(n45473), .Z(n45471) );
  OR U54796 ( .A(n45474), .B(n45475), .Z(n45470) );
  NAND U54797 ( .A(n45476), .B(n45477), .Z(n45368) );
  OR U54798 ( .A(n45478), .B(n45479), .Z(n45477) );
  OR U54799 ( .A(n45480), .B(n45481), .Z(n45476) );
  ANDN U54800 ( .B(n45482), .A(n45483), .Z(n45369) );
  IV U54801 ( .A(n45484), .Z(n45482) );
  XNOR U54802 ( .A(n45449), .B(n45448), .Z(N61372) );
  XOR U54803 ( .A(n45468), .B(n45467), .Z(n45448) );
  XNOR U54804 ( .A(n45483), .B(n45484), .Z(n45467) );
  XNOR U54805 ( .A(n45478), .B(n45479), .Z(n45484) );
  XNOR U54806 ( .A(n45480), .B(n45481), .Z(n45479) );
  XNOR U54807 ( .A(y[1453]), .B(x[1453]), .Z(n45481) );
  XNOR U54808 ( .A(y[1454]), .B(x[1454]), .Z(n45480) );
  XNOR U54809 ( .A(y[1452]), .B(x[1452]), .Z(n45478) );
  XNOR U54810 ( .A(n45472), .B(n45473), .Z(n45483) );
  XNOR U54811 ( .A(y[1449]), .B(x[1449]), .Z(n45473) );
  XNOR U54812 ( .A(n45474), .B(n45475), .Z(n45472) );
  XNOR U54813 ( .A(y[1450]), .B(x[1450]), .Z(n45475) );
  XNOR U54814 ( .A(y[1451]), .B(x[1451]), .Z(n45474) );
  XNOR U54815 ( .A(n45465), .B(n45464), .Z(n45468) );
  XNOR U54816 ( .A(n45460), .B(n45461), .Z(n45464) );
  XNOR U54817 ( .A(y[1446]), .B(x[1446]), .Z(n45461) );
  XNOR U54818 ( .A(n45462), .B(n45463), .Z(n45460) );
  XNOR U54819 ( .A(y[1447]), .B(x[1447]), .Z(n45463) );
  XNOR U54820 ( .A(y[1448]), .B(x[1448]), .Z(n45462) );
  XNOR U54821 ( .A(n45454), .B(n45455), .Z(n45465) );
  XNOR U54822 ( .A(y[1443]), .B(x[1443]), .Z(n45455) );
  XNOR U54823 ( .A(n45456), .B(n45457), .Z(n45454) );
  XNOR U54824 ( .A(y[1444]), .B(x[1444]), .Z(n45457) );
  XNOR U54825 ( .A(y[1445]), .B(x[1445]), .Z(n45456) );
  XOR U54826 ( .A(n45430), .B(n45431), .Z(n45449) );
  XNOR U54827 ( .A(n45446), .B(n45447), .Z(n45431) );
  XNOR U54828 ( .A(n45441), .B(n45442), .Z(n45447) );
  XNOR U54829 ( .A(n45443), .B(n45444), .Z(n45442) );
  XNOR U54830 ( .A(y[1441]), .B(x[1441]), .Z(n45444) );
  XNOR U54831 ( .A(y[1442]), .B(x[1442]), .Z(n45443) );
  XNOR U54832 ( .A(y[1440]), .B(x[1440]), .Z(n45441) );
  XNOR U54833 ( .A(n45435), .B(n45436), .Z(n45446) );
  XNOR U54834 ( .A(y[1437]), .B(x[1437]), .Z(n45436) );
  XNOR U54835 ( .A(n45437), .B(n45438), .Z(n45435) );
  XNOR U54836 ( .A(y[1438]), .B(x[1438]), .Z(n45438) );
  XNOR U54837 ( .A(y[1439]), .B(x[1439]), .Z(n45437) );
  XOR U54838 ( .A(n45429), .B(n45428), .Z(n45430) );
  XNOR U54839 ( .A(n45424), .B(n45425), .Z(n45428) );
  XNOR U54840 ( .A(y[1434]), .B(x[1434]), .Z(n45425) );
  XNOR U54841 ( .A(n45426), .B(n45427), .Z(n45424) );
  XNOR U54842 ( .A(y[1435]), .B(x[1435]), .Z(n45427) );
  XNOR U54843 ( .A(y[1436]), .B(x[1436]), .Z(n45426) );
  XNOR U54844 ( .A(n45418), .B(n45419), .Z(n45429) );
  XNOR U54845 ( .A(y[1431]), .B(x[1431]), .Z(n45419) );
  XNOR U54846 ( .A(n45420), .B(n45421), .Z(n45418) );
  XNOR U54847 ( .A(y[1432]), .B(x[1432]), .Z(n45421) );
  XNOR U54848 ( .A(y[1433]), .B(x[1433]), .Z(n45420) );
  NAND U54849 ( .A(n45485), .B(n45486), .Z(N61363) );
  NANDN U54850 ( .A(n45487), .B(n45488), .Z(n45486) );
  OR U54851 ( .A(n45489), .B(n45490), .Z(n45488) );
  NAND U54852 ( .A(n45489), .B(n45490), .Z(n45485) );
  XOR U54853 ( .A(n45489), .B(n45491), .Z(N61362) );
  XNOR U54854 ( .A(n45487), .B(n45490), .Z(n45491) );
  AND U54855 ( .A(n45492), .B(n45493), .Z(n45490) );
  NANDN U54856 ( .A(n45494), .B(n45495), .Z(n45493) );
  NANDN U54857 ( .A(n45496), .B(n45497), .Z(n45495) );
  NANDN U54858 ( .A(n45497), .B(n45496), .Z(n45492) );
  NAND U54859 ( .A(n45498), .B(n45499), .Z(n45487) );
  NANDN U54860 ( .A(n45500), .B(n45501), .Z(n45499) );
  OR U54861 ( .A(n45502), .B(n45503), .Z(n45501) );
  NAND U54862 ( .A(n45503), .B(n45502), .Z(n45498) );
  AND U54863 ( .A(n45504), .B(n45505), .Z(n45489) );
  NANDN U54864 ( .A(n45506), .B(n45507), .Z(n45505) );
  NANDN U54865 ( .A(n45508), .B(n45509), .Z(n45507) );
  NANDN U54866 ( .A(n45509), .B(n45508), .Z(n45504) );
  XOR U54867 ( .A(n45503), .B(n45510), .Z(N61361) );
  XOR U54868 ( .A(n45500), .B(n45502), .Z(n45510) );
  XNOR U54869 ( .A(n45496), .B(n45511), .Z(n45502) );
  XNOR U54870 ( .A(n45494), .B(n45497), .Z(n45511) );
  NAND U54871 ( .A(n45512), .B(n45513), .Z(n45497) );
  NAND U54872 ( .A(n45514), .B(n45515), .Z(n45513) );
  OR U54873 ( .A(n45516), .B(n45517), .Z(n45514) );
  NANDN U54874 ( .A(n45518), .B(n45516), .Z(n45512) );
  IV U54875 ( .A(n45517), .Z(n45518) );
  NAND U54876 ( .A(n45519), .B(n45520), .Z(n45494) );
  NAND U54877 ( .A(n45521), .B(n45522), .Z(n45520) );
  NANDN U54878 ( .A(n45523), .B(n45524), .Z(n45521) );
  NANDN U54879 ( .A(n45524), .B(n45523), .Z(n45519) );
  AND U54880 ( .A(n45525), .B(n45526), .Z(n45496) );
  NAND U54881 ( .A(n45527), .B(n45528), .Z(n45526) );
  OR U54882 ( .A(n45529), .B(n45530), .Z(n45527) );
  NANDN U54883 ( .A(n45531), .B(n45529), .Z(n45525) );
  NAND U54884 ( .A(n45532), .B(n45533), .Z(n45500) );
  NANDN U54885 ( .A(n45534), .B(n45535), .Z(n45533) );
  OR U54886 ( .A(n45536), .B(n45537), .Z(n45535) );
  NANDN U54887 ( .A(n45538), .B(n45536), .Z(n45532) );
  IV U54888 ( .A(n45537), .Z(n45538) );
  XNOR U54889 ( .A(n45508), .B(n45539), .Z(n45503) );
  XNOR U54890 ( .A(n45506), .B(n45509), .Z(n45539) );
  NAND U54891 ( .A(n45540), .B(n45541), .Z(n45509) );
  NAND U54892 ( .A(n45542), .B(n45543), .Z(n45541) );
  OR U54893 ( .A(n45544), .B(n45545), .Z(n45542) );
  NANDN U54894 ( .A(n45546), .B(n45544), .Z(n45540) );
  IV U54895 ( .A(n45545), .Z(n45546) );
  NAND U54896 ( .A(n45547), .B(n45548), .Z(n45506) );
  NAND U54897 ( .A(n45549), .B(n45550), .Z(n45548) );
  NANDN U54898 ( .A(n45551), .B(n45552), .Z(n45549) );
  NANDN U54899 ( .A(n45552), .B(n45551), .Z(n45547) );
  AND U54900 ( .A(n45553), .B(n45554), .Z(n45508) );
  NAND U54901 ( .A(n45555), .B(n45556), .Z(n45554) );
  OR U54902 ( .A(n45557), .B(n45558), .Z(n45555) );
  NANDN U54903 ( .A(n45559), .B(n45557), .Z(n45553) );
  XNOR U54904 ( .A(n45534), .B(n45560), .Z(N61360) );
  XOR U54905 ( .A(n45536), .B(n45537), .Z(n45560) );
  XNOR U54906 ( .A(n45550), .B(n45561), .Z(n45537) );
  XOR U54907 ( .A(n45551), .B(n45552), .Z(n45561) );
  XOR U54908 ( .A(n45557), .B(n45562), .Z(n45552) );
  XOR U54909 ( .A(n45556), .B(n45559), .Z(n45562) );
  IV U54910 ( .A(n45558), .Z(n45559) );
  NAND U54911 ( .A(n45563), .B(n45564), .Z(n45558) );
  OR U54912 ( .A(n45565), .B(n45566), .Z(n45564) );
  OR U54913 ( .A(n45567), .B(n45568), .Z(n45563) );
  NAND U54914 ( .A(n45569), .B(n45570), .Z(n45556) );
  OR U54915 ( .A(n45571), .B(n45572), .Z(n45570) );
  OR U54916 ( .A(n45573), .B(n45574), .Z(n45569) );
  NOR U54917 ( .A(n45575), .B(n45576), .Z(n45557) );
  ANDN U54918 ( .B(n45577), .A(n45578), .Z(n45551) );
  XNOR U54919 ( .A(n45544), .B(n45579), .Z(n45550) );
  XNOR U54920 ( .A(n45543), .B(n45545), .Z(n45579) );
  NAND U54921 ( .A(n45580), .B(n45581), .Z(n45545) );
  OR U54922 ( .A(n45582), .B(n45583), .Z(n45581) );
  OR U54923 ( .A(n45584), .B(n45585), .Z(n45580) );
  NAND U54924 ( .A(n45586), .B(n45587), .Z(n45543) );
  OR U54925 ( .A(n45588), .B(n45589), .Z(n45587) );
  OR U54926 ( .A(n45590), .B(n45591), .Z(n45586) );
  ANDN U54927 ( .B(n45592), .A(n45593), .Z(n45544) );
  IV U54928 ( .A(n45594), .Z(n45592) );
  ANDN U54929 ( .B(n45595), .A(n45596), .Z(n45536) );
  XOR U54930 ( .A(n45522), .B(n45597), .Z(n45534) );
  XOR U54931 ( .A(n45523), .B(n45524), .Z(n45597) );
  XOR U54932 ( .A(n45529), .B(n45598), .Z(n45524) );
  XOR U54933 ( .A(n45528), .B(n45531), .Z(n45598) );
  IV U54934 ( .A(n45530), .Z(n45531) );
  NAND U54935 ( .A(n45599), .B(n45600), .Z(n45530) );
  OR U54936 ( .A(n45601), .B(n45602), .Z(n45600) );
  OR U54937 ( .A(n45603), .B(n45604), .Z(n45599) );
  NAND U54938 ( .A(n45605), .B(n45606), .Z(n45528) );
  OR U54939 ( .A(n45607), .B(n45608), .Z(n45606) );
  OR U54940 ( .A(n45609), .B(n45610), .Z(n45605) );
  NOR U54941 ( .A(n45611), .B(n45612), .Z(n45529) );
  ANDN U54942 ( .B(n45613), .A(n45614), .Z(n45523) );
  IV U54943 ( .A(n45615), .Z(n45613) );
  XNOR U54944 ( .A(n45516), .B(n45616), .Z(n45522) );
  XNOR U54945 ( .A(n45515), .B(n45517), .Z(n45616) );
  NAND U54946 ( .A(n45617), .B(n45618), .Z(n45517) );
  OR U54947 ( .A(n45619), .B(n45620), .Z(n45618) );
  OR U54948 ( .A(n45621), .B(n45622), .Z(n45617) );
  NAND U54949 ( .A(n45623), .B(n45624), .Z(n45515) );
  OR U54950 ( .A(n45625), .B(n45626), .Z(n45624) );
  OR U54951 ( .A(n45627), .B(n45628), .Z(n45623) );
  ANDN U54952 ( .B(n45629), .A(n45630), .Z(n45516) );
  IV U54953 ( .A(n45631), .Z(n45629) );
  XNOR U54954 ( .A(n45596), .B(n45595), .Z(N61359) );
  XOR U54955 ( .A(n45615), .B(n45614), .Z(n45595) );
  XNOR U54956 ( .A(n45630), .B(n45631), .Z(n45614) );
  XNOR U54957 ( .A(n45625), .B(n45626), .Z(n45631) );
  XNOR U54958 ( .A(n45627), .B(n45628), .Z(n45626) );
  XNOR U54959 ( .A(y[1429]), .B(x[1429]), .Z(n45628) );
  XNOR U54960 ( .A(y[1430]), .B(x[1430]), .Z(n45627) );
  XNOR U54961 ( .A(y[1428]), .B(x[1428]), .Z(n45625) );
  XNOR U54962 ( .A(n45619), .B(n45620), .Z(n45630) );
  XNOR U54963 ( .A(y[1425]), .B(x[1425]), .Z(n45620) );
  XNOR U54964 ( .A(n45621), .B(n45622), .Z(n45619) );
  XNOR U54965 ( .A(y[1426]), .B(x[1426]), .Z(n45622) );
  XNOR U54966 ( .A(y[1427]), .B(x[1427]), .Z(n45621) );
  XNOR U54967 ( .A(n45612), .B(n45611), .Z(n45615) );
  XNOR U54968 ( .A(n45607), .B(n45608), .Z(n45611) );
  XNOR U54969 ( .A(y[1422]), .B(x[1422]), .Z(n45608) );
  XNOR U54970 ( .A(n45609), .B(n45610), .Z(n45607) );
  XNOR U54971 ( .A(y[1423]), .B(x[1423]), .Z(n45610) );
  XNOR U54972 ( .A(y[1424]), .B(x[1424]), .Z(n45609) );
  XNOR U54973 ( .A(n45601), .B(n45602), .Z(n45612) );
  XNOR U54974 ( .A(y[1419]), .B(x[1419]), .Z(n45602) );
  XNOR U54975 ( .A(n45603), .B(n45604), .Z(n45601) );
  XNOR U54976 ( .A(y[1420]), .B(x[1420]), .Z(n45604) );
  XNOR U54977 ( .A(y[1421]), .B(x[1421]), .Z(n45603) );
  XOR U54978 ( .A(n45577), .B(n45578), .Z(n45596) );
  XNOR U54979 ( .A(n45593), .B(n45594), .Z(n45578) );
  XNOR U54980 ( .A(n45588), .B(n45589), .Z(n45594) );
  XNOR U54981 ( .A(n45590), .B(n45591), .Z(n45589) );
  XNOR U54982 ( .A(y[1417]), .B(x[1417]), .Z(n45591) );
  XNOR U54983 ( .A(y[1418]), .B(x[1418]), .Z(n45590) );
  XNOR U54984 ( .A(y[1416]), .B(x[1416]), .Z(n45588) );
  XNOR U54985 ( .A(n45582), .B(n45583), .Z(n45593) );
  XNOR U54986 ( .A(y[1413]), .B(x[1413]), .Z(n45583) );
  XNOR U54987 ( .A(n45584), .B(n45585), .Z(n45582) );
  XNOR U54988 ( .A(y[1414]), .B(x[1414]), .Z(n45585) );
  XNOR U54989 ( .A(y[1415]), .B(x[1415]), .Z(n45584) );
  XOR U54990 ( .A(n45576), .B(n45575), .Z(n45577) );
  XNOR U54991 ( .A(n45571), .B(n45572), .Z(n45575) );
  XNOR U54992 ( .A(y[1410]), .B(x[1410]), .Z(n45572) );
  XNOR U54993 ( .A(n45573), .B(n45574), .Z(n45571) );
  XNOR U54994 ( .A(y[1411]), .B(x[1411]), .Z(n45574) );
  XNOR U54995 ( .A(y[1412]), .B(x[1412]), .Z(n45573) );
  XNOR U54996 ( .A(n45565), .B(n45566), .Z(n45576) );
  XNOR U54997 ( .A(y[1407]), .B(x[1407]), .Z(n45566) );
  XNOR U54998 ( .A(n45567), .B(n45568), .Z(n45565) );
  XNOR U54999 ( .A(y[1408]), .B(x[1408]), .Z(n45568) );
  XNOR U55000 ( .A(y[1409]), .B(x[1409]), .Z(n45567) );
  NAND U55001 ( .A(n45632), .B(n45633), .Z(N61350) );
  NANDN U55002 ( .A(n45634), .B(n45635), .Z(n45633) );
  OR U55003 ( .A(n45636), .B(n45637), .Z(n45635) );
  NAND U55004 ( .A(n45636), .B(n45637), .Z(n45632) );
  XOR U55005 ( .A(n45636), .B(n45638), .Z(N61349) );
  XNOR U55006 ( .A(n45634), .B(n45637), .Z(n45638) );
  AND U55007 ( .A(n45639), .B(n45640), .Z(n45637) );
  NANDN U55008 ( .A(n45641), .B(n45642), .Z(n45640) );
  NANDN U55009 ( .A(n45643), .B(n45644), .Z(n45642) );
  NANDN U55010 ( .A(n45644), .B(n45643), .Z(n45639) );
  NAND U55011 ( .A(n45645), .B(n45646), .Z(n45634) );
  NANDN U55012 ( .A(n45647), .B(n45648), .Z(n45646) );
  OR U55013 ( .A(n45649), .B(n45650), .Z(n45648) );
  NAND U55014 ( .A(n45650), .B(n45649), .Z(n45645) );
  AND U55015 ( .A(n45651), .B(n45652), .Z(n45636) );
  NANDN U55016 ( .A(n45653), .B(n45654), .Z(n45652) );
  NANDN U55017 ( .A(n45655), .B(n45656), .Z(n45654) );
  NANDN U55018 ( .A(n45656), .B(n45655), .Z(n45651) );
  XOR U55019 ( .A(n45650), .B(n45657), .Z(N61348) );
  XOR U55020 ( .A(n45647), .B(n45649), .Z(n45657) );
  XNOR U55021 ( .A(n45643), .B(n45658), .Z(n45649) );
  XNOR U55022 ( .A(n45641), .B(n45644), .Z(n45658) );
  NAND U55023 ( .A(n45659), .B(n45660), .Z(n45644) );
  NAND U55024 ( .A(n45661), .B(n45662), .Z(n45660) );
  OR U55025 ( .A(n45663), .B(n45664), .Z(n45661) );
  NANDN U55026 ( .A(n45665), .B(n45663), .Z(n45659) );
  IV U55027 ( .A(n45664), .Z(n45665) );
  NAND U55028 ( .A(n45666), .B(n45667), .Z(n45641) );
  NAND U55029 ( .A(n45668), .B(n45669), .Z(n45667) );
  NANDN U55030 ( .A(n45670), .B(n45671), .Z(n45668) );
  NANDN U55031 ( .A(n45671), .B(n45670), .Z(n45666) );
  AND U55032 ( .A(n45672), .B(n45673), .Z(n45643) );
  NAND U55033 ( .A(n45674), .B(n45675), .Z(n45673) );
  OR U55034 ( .A(n45676), .B(n45677), .Z(n45674) );
  NANDN U55035 ( .A(n45678), .B(n45676), .Z(n45672) );
  NAND U55036 ( .A(n45679), .B(n45680), .Z(n45647) );
  NANDN U55037 ( .A(n45681), .B(n45682), .Z(n45680) );
  OR U55038 ( .A(n45683), .B(n45684), .Z(n45682) );
  NANDN U55039 ( .A(n45685), .B(n45683), .Z(n45679) );
  IV U55040 ( .A(n45684), .Z(n45685) );
  XNOR U55041 ( .A(n45655), .B(n45686), .Z(n45650) );
  XNOR U55042 ( .A(n45653), .B(n45656), .Z(n45686) );
  NAND U55043 ( .A(n45687), .B(n45688), .Z(n45656) );
  NAND U55044 ( .A(n45689), .B(n45690), .Z(n45688) );
  OR U55045 ( .A(n45691), .B(n45692), .Z(n45689) );
  NANDN U55046 ( .A(n45693), .B(n45691), .Z(n45687) );
  IV U55047 ( .A(n45692), .Z(n45693) );
  NAND U55048 ( .A(n45694), .B(n45695), .Z(n45653) );
  NAND U55049 ( .A(n45696), .B(n45697), .Z(n45695) );
  NANDN U55050 ( .A(n45698), .B(n45699), .Z(n45696) );
  NANDN U55051 ( .A(n45699), .B(n45698), .Z(n45694) );
  AND U55052 ( .A(n45700), .B(n45701), .Z(n45655) );
  NAND U55053 ( .A(n45702), .B(n45703), .Z(n45701) );
  OR U55054 ( .A(n45704), .B(n45705), .Z(n45702) );
  NANDN U55055 ( .A(n45706), .B(n45704), .Z(n45700) );
  XNOR U55056 ( .A(n45681), .B(n45707), .Z(N61347) );
  XOR U55057 ( .A(n45683), .B(n45684), .Z(n45707) );
  XNOR U55058 ( .A(n45697), .B(n45708), .Z(n45684) );
  XOR U55059 ( .A(n45698), .B(n45699), .Z(n45708) );
  XOR U55060 ( .A(n45704), .B(n45709), .Z(n45699) );
  XOR U55061 ( .A(n45703), .B(n45706), .Z(n45709) );
  IV U55062 ( .A(n45705), .Z(n45706) );
  NAND U55063 ( .A(n45710), .B(n45711), .Z(n45705) );
  OR U55064 ( .A(n45712), .B(n45713), .Z(n45711) );
  OR U55065 ( .A(n45714), .B(n45715), .Z(n45710) );
  NAND U55066 ( .A(n45716), .B(n45717), .Z(n45703) );
  OR U55067 ( .A(n45718), .B(n45719), .Z(n45717) );
  OR U55068 ( .A(n45720), .B(n45721), .Z(n45716) );
  NOR U55069 ( .A(n45722), .B(n45723), .Z(n45704) );
  ANDN U55070 ( .B(n45724), .A(n45725), .Z(n45698) );
  XNOR U55071 ( .A(n45691), .B(n45726), .Z(n45697) );
  XNOR U55072 ( .A(n45690), .B(n45692), .Z(n45726) );
  NAND U55073 ( .A(n45727), .B(n45728), .Z(n45692) );
  OR U55074 ( .A(n45729), .B(n45730), .Z(n45728) );
  OR U55075 ( .A(n45731), .B(n45732), .Z(n45727) );
  NAND U55076 ( .A(n45733), .B(n45734), .Z(n45690) );
  OR U55077 ( .A(n45735), .B(n45736), .Z(n45734) );
  OR U55078 ( .A(n45737), .B(n45738), .Z(n45733) );
  ANDN U55079 ( .B(n45739), .A(n45740), .Z(n45691) );
  IV U55080 ( .A(n45741), .Z(n45739) );
  ANDN U55081 ( .B(n45742), .A(n45743), .Z(n45683) );
  XOR U55082 ( .A(n45669), .B(n45744), .Z(n45681) );
  XOR U55083 ( .A(n45670), .B(n45671), .Z(n45744) );
  XOR U55084 ( .A(n45676), .B(n45745), .Z(n45671) );
  XOR U55085 ( .A(n45675), .B(n45678), .Z(n45745) );
  IV U55086 ( .A(n45677), .Z(n45678) );
  NAND U55087 ( .A(n45746), .B(n45747), .Z(n45677) );
  OR U55088 ( .A(n45748), .B(n45749), .Z(n45747) );
  OR U55089 ( .A(n45750), .B(n45751), .Z(n45746) );
  NAND U55090 ( .A(n45752), .B(n45753), .Z(n45675) );
  OR U55091 ( .A(n45754), .B(n45755), .Z(n45753) );
  OR U55092 ( .A(n45756), .B(n45757), .Z(n45752) );
  NOR U55093 ( .A(n45758), .B(n45759), .Z(n45676) );
  ANDN U55094 ( .B(n45760), .A(n45761), .Z(n45670) );
  IV U55095 ( .A(n45762), .Z(n45760) );
  XNOR U55096 ( .A(n45663), .B(n45763), .Z(n45669) );
  XNOR U55097 ( .A(n45662), .B(n45664), .Z(n45763) );
  NAND U55098 ( .A(n45764), .B(n45765), .Z(n45664) );
  OR U55099 ( .A(n45766), .B(n45767), .Z(n45765) );
  OR U55100 ( .A(n45768), .B(n45769), .Z(n45764) );
  NAND U55101 ( .A(n45770), .B(n45771), .Z(n45662) );
  OR U55102 ( .A(n45772), .B(n45773), .Z(n45771) );
  OR U55103 ( .A(n45774), .B(n45775), .Z(n45770) );
  ANDN U55104 ( .B(n45776), .A(n45777), .Z(n45663) );
  IV U55105 ( .A(n45778), .Z(n45776) );
  XNOR U55106 ( .A(n45743), .B(n45742), .Z(N61346) );
  XOR U55107 ( .A(n45762), .B(n45761), .Z(n45742) );
  XNOR U55108 ( .A(n45777), .B(n45778), .Z(n45761) );
  XNOR U55109 ( .A(n45772), .B(n45773), .Z(n45778) );
  XNOR U55110 ( .A(n45774), .B(n45775), .Z(n45773) );
  XNOR U55111 ( .A(y[1405]), .B(x[1405]), .Z(n45775) );
  XNOR U55112 ( .A(y[1406]), .B(x[1406]), .Z(n45774) );
  XNOR U55113 ( .A(y[1404]), .B(x[1404]), .Z(n45772) );
  XNOR U55114 ( .A(n45766), .B(n45767), .Z(n45777) );
  XNOR U55115 ( .A(y[1401]), .B(x[1401]), .Z(n45767) );
  XNOR U55116 ( .A(n45768), .B(n45769), .Z(n45766) );
  XNOR U55117 ( .A(y[1402]), .B(x[1402]), .Z(n45769) );
  XNOR U55118 ( .A(y[1403]), .B(x[1403]), .Z(n45768) );
  XNOR U55119 ( .A(n45759), .B(n45758), .Z(n45762) );
  XNOR U55120 ( .A(n45754), .B(n45755), .Z(n45758) );
  XNOR U55121 ( .A(y[1398]), .B(x[1398]), .Z(n45755) );
  XNOR U55122 ( .A(n45756), .B(n45757), .Z(n45754) );
  XNOR U55123 ( .A(y[1399]), .B(x[1399]), .Z(n45757) );
  XNOR U55124 ( .A(y[1400]), .B(x[1400]), .Z(n45756) );
  XNOR U55125 ( .A(n45748), .B(n45749), .Z(n45759) );
  XNOR U55126 ( .A(y[1395]), .B(x[1395]), .Z(n45749) );
  XNOR U55127 ( .A(n45750), .B(n45751), .Z(n45748) );
  XNOR U55128 ( .A(y[1396]), .B(x[1396]), .Z(n45751) );
  XNOR U55129 ( .A(y[1397]), .B(x[1397]), .Z(n45750) );
  XOR U55130 ( .A(n45724), .B(n45725), .Z(n45743) );
  XNOR U55131 ( .A(n45740), .B(n45741), .Z(n45725) );
  XNOR U55132 ( .A(n45735), .B(n45736), .Z(n45741) );
  XNOR U55133 ( .A(n45737), .B(n45738), .Z(n45736) );
  XNOR U55134 ( .A(y[1393]), .B(x[1393]), .Z(n45738) );
  XNOR U55135 ( .A(y[1394]), .B(x[1394]), .Z(n45737) );
  XNOR U55136 ( .A(y[1392]), .B(x[1392]), .Z(n45735) );
  XNOR U55137 ( .A(n45729), .B(n45730), .Z(n45740) );
  XNOR U55138 ( .A(y[1389]), .B(x[1389]), .Z(n45730) );
  XNOR U55139 ( .A(n45731), .B(n45732), .Z(n45729) );
  XNOR U55140 ( .A(y[1390]), .B(x[1390]), .Z(n45732) );
  XNOR U55141 ( .A(y[1391]), .B(x[1391]), .Z(n45731) );
  XOR U55142 ( .A(n45723), .B(n45722), .Z(n45724) );
  XNOR U55143 ( .A(n45718), .B(n45719), .Z(n45722) );
  XNOR U55144 ( .A(y[1386]), .B(x[1386]), .Z(n45719) );
  XNOR U55145 ( .A(n45720), .B(n45721), .Z(n45718) );
  XNOR U55146 ( .A(y[1387]), .B(x[1387]), .Z(n45721) );
  XNOR U55147 ( .A(y[1388]), .B(x[1388]), .Z(n45720) );
  XNOR U55148 ( .A(n45712), .B(n45713), .Z(n45723) );
  XNOR U55149 ( .A(y[1383]), .B(x[1383]), .Z(n45713) );
  XNOR U55150 ( .A(n45714), .B(n45715), .Z(n45712) );
  XNOR U55151 ( .A(y[1384]), .B(x[1384]), .Z(n45715) );
  XNOR U55152 ( .A(y[1385]), .B(x[1385]), .Z(n45714) );
  NAND U55153 ( .A(n45779), .B(n45780), .Z(N61337) );
  NANDN U55154 ( .A(n45781), .B(n45782), .Z(n45780) );
  OR U55155 ( .A(n45783), .B(n45784), .Z(n45782) );
  NAND U55156 ( .A(n45783), .B(n45784), .Z(n45779) );
  XOR U55157 ( .A(n45783), .B(n45785), .Z(N61336) );
  XNOR U55158 ( .A(n45781), .B(n45784), .Z(n45785) );
  AND U55159 ( .A(n45786), .B(n45787), .Z(n45784) );
  NANDN U55160 ( .A(n45788), .B(n45789), .Z(n45787) );
  NANDN U55161 ( .A(n45790), .B(n45791), .Z(n45789) );
  NANDN U55162 ( .A(n45791), .B(n45790), .Z(n45786) );
  NAND U55163 ( .A(n45792), .B(n45793), .Z(n45781) );
  NANDN U55164 ( .A(n45794), .B(n45795), .Z(n45793) );
  OR U55165 ( .A(n45796), .B(n45797), .Z(n45795) );
  NAND U55166 ( .A(n45797), .B(n45796), .Z(n45792) );
  AND U55167 ( .A(n45798), .B(n45799), .Z(n45783) );
  NANDN U55168 ( .A(n45800), .B(n45801), .Z(n45799) );
  NANDN U55169 ( .A(n45802), .B(n45803), .Z(n45801) );
  NANDN U55170 ( .A(n45803), .B(n45802), .Z(n45798) );
  XOR U55171 ( .A(n45797), .B(n45804), .Z(N61335) );
  XOR U55172 ( .A(n45794), .B(n45796), .Z(n45804) );
  XNOR U55173 ( .A(n45790), .B(n45805), .Z(n45796) );
  XNOR U55174 ( .A(n45788), .B(n45791), .Z(n45805) );
  NAND U55175 ( .A(n45806), .B(n45807), .Z(n45791) );
  NAND U55176 ( .A(n45808), .B(n45809), .Z(n45807) );
  OR U55177 ( .A(n45810), .B(n45811), .Z(n45808) );
  NANDN U55178 ( .A(n45812), .B(n45810), .Z(n45806) );
  IV U55179 ( .A(n45811), .Z(n45812) );
  NAND U55180 ( .A(n45813), .B(n45814), .Z(n45788) );
  NAND U55181 ( .A(n45815), .B(n45816), .Z(n45814) );
  NANDN U55182 ( .A(n45817), .B(n45818), .Z(n45815) );
  NANDN U55183 ( .A(n45818), .B(n45817), .Z(n45813) );
  AND U55184 ( .A(n45819), .B(n45820), .Z(n45790) );
  NAND U55185 ( .A(n45821), .B(n45822), .Z(n45820) );
  OR U55186 ( .A(n45823), .B(n45824), .Z(n45821) );
  NANDN U55187 ( .A(n45825), .B(n45823), .Z(n45819) );
  NAND U55188 ( .A(n45826), .B(n45827), .Z(n45794) );
  NANDN U55189 ( .A(n45828), .B(n45829), .Z(n45827) );
  OR U55190 ( .A(n45830), .B(n45831), .Z(n45829) );
  NANDN U55191 ( .A(n45832), .B(n45830), .Z(n45826) );
  IV U55192 ( .A(n45831), .Z(n45832) );
  XNOR U55193 ( .A(n45802), .B(n45833), .Z(n45797) );
  XNOR U55194 ( .A(n45800), .B(n45803), .Z(n45833) );
  NAND U55195 ( .A(n45834), .B(n45835), .Z(n45803) );
  NAND U55196 ( .A(n45836), .B(n45837), .Z(n45835) );
  OR U55197 ( .A(n45838), .B(n45839), .Z(n45836) );
  NANDN U55198 ( .A(n45840), .B(n45838), .Z(n45834) );
  IV U55199 ( .A(n45839), .Z(n45840) );
  NAND U55200 ( .A(n45841), .B(n45842), .Z(n45800) );
  NAND U55201 ( .A(n45843), .B(n45844), .Z(n45842) );
  NANDN U55202 ( .A(n45845), .B(n45846), .Z(n45843) );
  NANDN U55203 ( .A(n45846), .B(n45845), .Z(n45841) );
  AND U55204 ( .A(n45847), .B(n45848), .Z(n45802) );
  NAND U55205 ( .A(n45849), .B(n45850), .Z(n45848) );
  OR U55206 ( .A(n45851), .B(n45852), .Z(n45849) );
  NANDN U55207 ( .A(n45853), .B(n45851), .Z(n45847) );
  XNOR U55208 ( .A(n45828), .B(n45854), .Z(N61334) );
  XOR U55209 ( .A(n45830), .B(n45831), .Z(n45854) );
  XNOR U55210 ( .A(n45844), .B(n45855), .Z(n45831) );
  XOR U55211 ( .A(n45845), .B(n45846), .Z(n45855) );
  XOR U55212 ( .A(n45851), .B(n45856), .Z(n45846) );
  XOR U55213 ( .A(n45850), .B(n45853), .Z(n45856) );
  IV U55214 ( .A(n45852), .Z(n45853) );
  NAND U55215 ( .A(n45857), .B(n45858), .Z(n45852) );
  OR U55216 ( .A(n45859), .B(n45860), .Z(n45858) );
  OR U55217 ( .A(n45861), .B(n45862), .Z(n45857) );
  NAND U55218 ( .A(n45863), .B(n45864), .Z(n45850) );
  OR U55219 ( .A(n45865), .B(n45866), .Z(n45864) );
  OR U55220 ( .A(n45867), .B(n45868), .Z(n45863) );
  NOR U55221 ( .A(n45869), .B(n45870), .Z(n45851) );
  ANDN U55222 ( .B(n45871), .A(n45872), .Z(n45845) );
  XNOR U55223 ( .A(n45838), .B(n45873), .Z(n45844) );
  XNOR U55224 ( .A(n45837), .B(n45839), .Z(n45873) );
  NAND U55225 ( .A(n45874), .B(n45875), .Z(n45839) );
  OR U55226 ( .A(n45876), .B(n45877), .Z(n45875) );
  OR U55227 ( .A(n45878), .B(n45879), .Z(n45874) );
  NAND U55228 ( .A(n45880), .B(n45881), .Z(n45837) );
  OR U55229 ( .A(n45882), .B(n45883), .Z(n45881) );
  OR U55230 ( .A(n45884), .B(n45885), .Z(n45880) );
  ANDN U55231 ( .B(n45886), .A(n45887), .Z(n45838) );
  IV U55232 ( .A(n45888), .Z(n45886) );
  ANDN U55233 ( .B(n45889), .A(n45890), .Z(n45830) );
  XOR U55234 ( .A(n45816), .B(n45891), .Z(n45828) );
  XOR U55235 ( .A(n45817), .B(n45818), .Z(n45891) );
  XOR U55236 ( .A(n45823), .B(n45892), .Z(n45818) );
  XOR U55237 ( .A(n45822), .B(n45825), .Z(n45892) );
  IV U55238 ( .A(n45824), .Z(n45825) );
  NAND U55239 ( .A(n45893), .B(n45894), .Z(n45824) );
  OR U55240 ( .A(n45895), .B(n45896), .Z(n45894) );
  OR U55241 ( .A(n45897), .B(n45898), .Z(n45893) );
  NAND U55242 ( .A(n45899), .B(n45900), .Z(n45822) );
  OR U55243 ( .A(n45901), .B(n45902), .Z(n45900) );
  OR U55244 ( .A(n45903), .B(n45904), .Z(n45899) );
  NOR U55245 ( .A(n45905), .B(n45906), .Z(n45823) );
  ANDN U55246 ( .B(n45907), .A(n45908), .Z(n45817) );
  IV U55247 ( .A(n45909), .Z(n45907) );
  XNOR U55248 ( .A(n45810), .B(n45910), .Z(n45816) );
  XNOR U55249 ( .A(n45809), .B(n45811), .Z(n45910) );
  NAND U55250 ( .A(n45911), .B(n45912), .Z(n45811) );
  OR U55251 ( .A(n45913), .B(n45914), .Z(n45912) );
  OR U55252 ( .A(n45915), .B(n45916), .Z(n45911) );
  NAND U55253 ( .A(n45917), .B(n45918), .Z(n45809) );
  OR U55254 ( .A(n45919), .B(n45920), .Z(n45918) );
  OR U55255 ( .A(n45921), .B(n45922), .Z(n45917) );
  ANDN U55256 ( .B(n45923), .A(n45924), .Z(n45810) );
  IV U55257 ( .A(n45925), .Z(n45923) );
  XNOR U55258 ( .A(n45890), .B(n45889), .Z(N61333) );
  XOR U55259 ( .A(n45909), .B(n45908), .Z(n45889) );
  XNOR U55260 ( .A(n45924), .B(n45925), .Z(n45908) );
  XNOR U55261 ( .A(n45919), .B(n45920), .Z(n45925) );
  XNOR U55262 ( .A(n45921), .B(n45922), .Z(n45920) );
  XNOR U55263 ( .A(y[1381]), .B(x[1381]), .Z(n45922) );
  XNOR U55264 ( .A(y[1382]), .B(x[1382]), .Z(n45921) );
  XNOR U55265 ( .A(y[1380]), .B(x[1380]), .Z(n45919) );
  XNOR U55266 ( .A(n45913), .B(n45914), .Z(n45924) );
  XNOR U55267 ( .A(y[1377]), .B(x[1377]), .Z(n45914) );
  XNOR U55268 ( .A(n45915), .B(n45916), .Z(n45913) );
  XNOR U55269 ( .A(y[1378]), .B(x[1378]), .Z(n45916) );
  XNOR U55270 ( .A(y[1379]), .B(x[1379]), .Z(n45915) );
  XNOR U55271 ( .A(n45906), .B(n45905), .Z(n45909) );
  XNOR U55272 ( .A(n45901), .B(n45902), .Z(n45905) );
  XNOR U55273 ( .A(y[1374]), .B(x[1374]), .Z(n45902) );
  XNOR U55274 ( .A(n45903), .B(n45904), .Z(n45901) );
  XNOR U55275 ( .A(y[1375]), .B(x[1375]), .Z(n45904) );
  XNOR U55276 ( .A(y[1376]), .B(x[1376]), .Z(n45903) );
  XNOR U55277 ( .A(n45895), .B(n45896), .Z(n45906) );
  XNOR U55278 ( .A(y[1371]), .B(x[1371]), .Z(n45896) );
  XNOR U55279 ( .A(n45897), .B(n45898), .Z(n45895) );
  XNOR U55280 ( .A(y[1372]), .B(x[1372]), .Z(n45898) );
  XNOR U55281 ( .A(y[1373]), .B(x[1373]), .Z(n45897) );
  XOR U55282 ( .A(n45871), .B(n45872), .Z(n45890) );
  XNOR U55283 ( .A(n45887), .B(n45888), .Z(n45872) );
  XNOR U55284 ( .A(n45882), .B(n45883), .Z(n45888) );
  XNOR U55285 ( .A(n45884), .B(n45885), .Z(n45883) );
  XNOR U55286 ( .A(y[1369]), .B(x[1369]), .Z(n45885) );
  XNOR U55287 ( .A(y[1370]), .B(x[1370]), .Z(n45884) );
  XNOR U55288 ( .A(y[1368]), .B(x[1368]), .Z(n45882) );
  XNOR U55289 ( .A(n45876), .B(n45877), .Z(n45887) );
  XNOR U55290 ( .A(y[1365]), .B(x[1365]), .Z(n45877) );
  XNOR U55291 ( .A(n45878), .B(n45879), .Z(n45876) );
  XNOR U55292 ( .A(y[1366]), .B(x[1366]), .Z(n45879) );
  XNOR U55293 ( .A(y[1367]), .B(x[1367]), .Z(n45878) );
  XOR U55294 ( .A(n45870), .B(n45869), .Z(n45871) );
  XNOR U55295 ( .A(n45865), .B(n45866), .Z(n45869) );
  XNOR U55296 ( .A(y[1362]), .B(x[1362]), .Z(n45866) );
  XNOR U55297 ( .A(n45867), .B(n45868), .Z(n45865) );
  XNOR U55298 ( .A(y[1363]), .B(x[1363]), .Z(n45868) );
  XNOR U55299 ( .A(y[1364]), .B(x[1364]), .Z(n45867) );
  XNOR U55300 ( .A(n45859), .B(n45860), .Z(n45870) );
  XNOR U55301 ( .A(y[1359]), .B(x[1359]), .Z(n45860) );
  XNOR U55302 ( .A(n45861), .B(n45862), .Z(n45859) );
  XNOR U55303 ( .A(y[1360]), .B(x[1360]), .Z(n45862) );
  XNOR U55304 ( .A(y[1361]), .B(x[1361]), .Z(n45861) );
  NAND U55305 ( .A(n45926), .B(n45927), .Z(N61324) );
  NANDN U55306 ( .A(n45928), .B(n45929), .Z(n45927) );
  OR U55307 ( .A(n45930), .B(n45931), .Z(n45929) );
  NAND U55308 ( .A(n45930), .B(n45931), .Z(n45926) );
  XOR U55309 ( .A(n45930), .B(n45932), .Z(N61323) );
  XNOR U55310 ( .A(n45928), .B(n45931), .Z(n45932) );
  AND U55311 ( .A(n45933), .B(n45934), .Z(n45931) );
  NANDN U55312 ( .A(n45935), .B(n45936), .Z(n45934) );
  NANDN U55313 ( .A(n45937), .B(n45938), .Z(n45936) );
  NANDN U55314 ( .A(n45938), .B(n45937), .Z(n45933) );
  NAND U55315 ( .A(n45939), .B(n45940), .Z(n45928) );
  NANDN U55316 ( .A(n45941), .B(n45942), .Z(n45940) );
  OR U55317 ( .A(n45943), .B(n45944), .Z(n45942) );
  NAND U55318 ( .A(n45944), .B(n45943), .Z(n45939) );
  AND U55319 ( .A(n45945), .B(n45946), .Z(n45930) );
  NANDN U55320 ( .A(n45947), .B(n45948), .Z(n45946) );
  NANDN U55321 ( .A(n45949), .B(n45950), .Z(n45948) );
  NANDN U55322 ( .A(n45950), .B(n45949), .Z(n45945) );
  XOR U55323 ( .A(n45944), .B(n45951), .Z(N61322) );
  XOR U55324 ( .A(n45941), .B(n45943), .Z(n45951) );
  XNOR U55325 ( .A(n45937), .B(n45952), .Z(n45943) );
  XNOR U55326 ( .A(n45935), .B(n45938), .Z(n45952) );
  NAND U55327 ( .A(n45953), .B(n45954), .Z(n45938) );
  NAND U55328 ( .A(n45955), .B(n45956), .Z(n45954) );
  OR U55329 ( .A(n45957), .B(n45958), .Z(n45955) );
  NANDN U55330 ( .A(n45959), .B(n45957), .Z(n45953) );
  IV U55331 ( .A(n45958), .Z(n45959) );
  NAND U55332 ( .A(n45960), .B(n45961), .Z(n45935) );
  NAND U55333 ( .A(n45962), .B(n45963), .Z(n45961) );
  NANDN U55334 ( .A(n45964), .B(n45965), .Z(n45962) );
  NANDN U55335 ( .A(n45965), .B(n45964), .Z(n45960) );
  AND U55336 ( .A(n45966), .B(n45967), .Z(n45937) );
  NAND U55337 ( .A(n45968), .B(n45969), .Z(n45967) );
  OR U55338 ( .A(n45970), .B(n45971), .Z(n45968) );
  NANDN U55339 ( .A(n45972), .B(n45970), .Z(n45966) );
  NAND U55340 ( .A(n45973), .B(n45974), .Z(n45941) );
  NANDN U55341 ( .A(n45975), .B(n45976), .Z(n45974) );
  OR U55342 ( .A(n45977), .B(n45978), .Z(n45976) );
  NANDN U55343 ( .A(n45979), .B(n45977), .Z(n45973) );
  IV U55344 ( .A(n45978), .Z(n45979) );
  XNOR U55345 ( .A(n45949), .B(n45980), .Z(n45944) );
  XNOR U55346 ( .A(n45947), .B(n45950), .Z(n45980) );
  NAND U55347 ( .A(n45981), .B(n45982), .Z(n45950) );
  NAND U55348 ( .A(n45983), .B(n45984), .Z(n45982) );
  OR U55349 ( .A(n45985), .B(n45986), .Z(n45983) );
  NANDN U55350 ( .A(n45987), .B(n45985), .Z(n45981) );
  IV U55351 ( .A(n45986), .Z(n45987) );
  NAND U55352 ( .A(n45988), .B(n45989), .Z(n45947) );
  NAND U55353 ( .A(n45990), .B(n45991), .Z(n45989) );
  NANDN U55354 ( .A(n45992), .B(n45993), .Z(n45990) );
  NANDN U55355 ( .A(n45993), .B(n45992), .Z(n45988) );
  AND U55356 ( .A(n45994), .B(n45995), .Z(n45949) );
  NAND U55357 ( .A(n45996), .B(n45997), .Z(n45995) );
  OR U55358 ( .A(n45998), .B(n45999), .Z(n45996) );
  NANDN U55359 ( .A(n46000), .B(n45998), .Z(n45994) );
  XNOR U55360 ( .A(n45975), .B(n46001), .Z(N61321) );
  XOR U55361 ( .A(n45977), .B(n45978), .Z(n46001) );
  XNOR U55362 ( .A(n45991), .B(n46002), .Z(n45978) );
  XOR U55363 ( .A(n45992), .B(n45993), .Z(n46002) );
  XOR U55364 ( .A(n45998), .B(n46003), .Z(n45993) );
  XOR U55365 ( .A(n45997), .B(n46000), .Z(n46003) );
  IV U55366 ( .A(n45999), .Z(n46000) );
  NAND U55367 ( .A(n46004), .B(n46005), .Z(n45999) );
  OR U55368 ( .A(n46006), .B(n46007), .Z(n46005) );
  OR U55369 ( .A(n46008), .B(n46009), .Z(n46004) );
  NAND U55370 ( .A(n46010), .B(n46011), .Z(n45997) );
  OR U55371 ( .A(n46012), .B(n46013), .Z(n46011) );
  OR U55372 ( .A(n46014), .B(n46015), .Z(n46010) );
  NOR U55373 ( .A(n46016), .B(n46017), .Z(n45998) );
  ANDN U55374 ( .B(n46018), .A(n46019), .Z(n45992) );
  XNOR U55375 ( .A(n45985), .B(n46020), .Z(n45991) );
  XNOR U55376 ( .A(n45984), .B(n45986), .Z(n46020) );
  NAND U55377 ( .A(n46021), .B(n46022), .Z(n45986) );
  OR U55378 ( .A(n46023), .B(n46024), .Z(n46022) );
  OR U55379 ( .A(n46025), .B(n46026), .Z(n46021) );
  NAND U55380 ( .A(n46027), .B(n46028), .Z(n45984) );
  OR U55381 ( .A(n46029), .B(n46030), .Z(n46028) );
  OR U55382 ( .A(n46031), .B(n46032), .Z(n46027) );
  ANDN U55383 ( .B(n46033), .A(n46034), .Z(n45985) );
  IV U55384 ( .A(n46035), .Z(n46033) );
  ANDN U55385 ( .B(n46036), .A(n46037), .Z(n45977) );
  XOR U55386 ( .A(n45963), .B(n46038), .Z(n45975) );
  XOR U55387 ( .A(n45964), .B(n45965), .Z(n46038) );
  XOR U55388 ( .A(n45970), .B(n46039), .Z(n45965) );
  XOR U55389 ( .A(n45969), .B(n45972), .Z(n46039) );
  IV U55390 ( .A(n45971), .Z(n45972) );
  NAND U55391 ( .A(n46040), .B(n46041), .Z(n45971) );
  OR U55392 ( .A(n46042), .B(n46043), .Z(n46041) );
  OR U55393 ( .A(n46044), .B(n46045), .Z(n46040) );
  NAND U55394 ( .A(n46046), .B(n46047), .Z(n45969) );
  OR U55395 ( .A(n46048), .B(n46049), .Z(n46047) );
  OR U55396 ( .A(n46050), .B(n46051), .Z(n46046) );
  NOR U55397 ( .A(n46052), .B(n46053), .Z(n45970) );
  ANDN U55398 ( .B(n46054), .A(n46055), .Z(n45964) );
  IV U55399 ( .A(n46056), .Z(n46054) );
  XNOR U55400 ( .A(n45957), .B(n46057), .Z(n45963) );
  XNOR U55401 ( .A(n45956), .B(n45958), .Z(n46057) );
  NAND U55402 ( .A(n46058), .B(n46059), .Z(n45958) );
  OR U55403 ( .A(n46060), .B(n46061), .Z(n46059) );
  OR U55404 ( .A(n46062), .B(n46063), .Z(n46058) );
  NAND U55405 ( .A(n46064), .B(n46065), .Z(n45956) );
  OR U55406 ( .A(n46066), .B(n46067), .Z(n46065) );
  OR U55407 ( .A(n46068), .B(n46069), .Z(n46064) );
  ANDN U55408 ( .B(n46070), .A(n46071), .Z(n45957) );
  IV U55409 ( .A(n46072), .Z(n46070) );
  XNOR U55410 ( .A(n46037), .B(n46036), .Z(N61320) );
  XOR U55411 ( .A(n46056), .B(n46055), .Z(n46036) );
  XNOR U55412 ( .A(n46071), .B(n46072), .Z(n46055) );
  XNOR U55413 ( .A(n46066), .B(n46067), .Z(n46072) );
  XNOR U55414 ( .A(n46068), .B(n46069), .Z(n46067) );
  XNOR U55415 ( .A(y[1357]), .B(x[1357]), .Z(n46069) );
  XNOR U55416 ( .A(y[1358]), .B(x[1358]), .Z(n46068) );
  XNOR U55417 ( .A(y[1356]), .B(x[1356]), .Z(n46066) );
  XNOR U55418 ( .A(n46060), .B(n46061), .Z(n46071) );
  XNOR U55419 ( .A(y[1353]), .B(x[1353]), .Z(n46061) );
  XNOR U55420 ( .A(n46062), .B(n46063), .Z(n46060) );
  XNOR U55421 ( .A(y[1354]), .B(x[1354]), .Z(n46063) );
  XNOR U55422 ( .A(y[1355]), .B(x[1355]), .Z(n46062) );
  XNOR U55423 ( .A(n46053), .B(n46052), .Z(n46056) );
  XNOR U55424 ( .A(n46048), .B(n46049), .Z(n46052) );
  XNOR U55425 ( .A(y[1350]), .B(x[1350]), .Z(n46049) );
  XNOR U55426 ( .A(n46050), .B(n46051), .Z(n46048) );
  XNOR U55427 ( .A(y[1351]), .B(x[1351]), .Z(n46051) );
  XNOR U55428 ( .A(y[1352]), .B(x[1352]), .Z(n46050) );
  XNOR U55429 ( .A(n46042), .B(n46043), .Z(n46053) );
  XNOR U55430 ( .A(y[1347]), .B(x[1347]), .Z(n46043) );
  XNOR U55431 ( .A(n46044), .B(n46045), .Z(n46042) );
  XNOR U55432 ( .A(y[1348]), .B(x[1348]), .Z(n46045) );
  XNOR U55433 ( .A(y[1349]), .B(x[1349]), .Z(n46044) );
  XOR U55434 ( .A(n46018), .B(n46019), .Z(n46037) );
  XNOR U55435 ( .A(n46034), .B(n46035), .Z(n46019) );
  XNOR U55436 ( .A(n46029), .B(n46030), .Z(n46035) );
  XNOR U55437 ( .A(n46031), .B(n46032), .Z(n46030) );
  XNOR U55438 ( .A(y[1345]), .B(x[1345]), .Z(n46032) );
  XNOR U55439 ( .A(y[1346]), .B(x[1346]), .Z(n46031) );
  XNOR U55440 ( .A(y[1344]), .B(x[1344]), .Z(n46029) );
  XNOR U55441 ( .A(n46023), .B(n46024), .Z(n46034) );
  XNOR U55442 ( .A(y[1341]), .B(x[1341]), .Z(n46024) );
  XNOR U55443 ( .A(n46025), .B(n46026), .Z(n46023) );
  XNOR U55444 ( .A(y[1342]), .B(x[1342]), .Z(n46026) );
  XNOR U55445 ( .A(y[1343]), .B(x[1343]), .Z(n46025) );
  XOR U55446 ( .A(n46017), .B(n46016), .Z(n46018) );
  XNOR U55447 ( .A(n46012), .B(n46013), .Z(n46016) );
  XNOR U55448 ( .A(y[1338]), .B(x[1338]), .Z(n46013) );
  XNOR U55449 ( .A(n46014), .B(n46015), .Z(n46012) );
  XNOR U55450 ( .A(y[1339]), .B(x[1339]), .Z(n46015) );
  XNOR U55451 ( .A(y[1340]), .B(x[1340]), .Z(n46014) );
  XNOR U55452 ( .A(n46006), .B(n46007), .Z(n46017) );
  XNOR U55453 ( .A(y[1335]), .B(x[1335]), .Z(n46007) );
  XNOR U55454 ( .A(n46008), .B(n46009), .Z(n46006) );
  XNOR U55455 ( .A(y[1336]), .B(x[1336]), .Z(n46009) );
  XNOR U55456 ( .A(y[1337]), .B(x[1337]), .Z(n46008) );
  NAND U55457 ( .A(n46073), .B(n46074), .Z(N61311) );
  NANDN U55458 ( .A(n46075), .B(n46076), .Z(n46074) );
  OR U55459 ( .A(n46077), .B(n46078), .Z(n46076) );
  NAND U55460 ( .A(n46077), .B(n46078), .Z(n46073) );
  XOR U55461 ( .A(n46077), .B(n46079), .Z(N61310) );
  XNOR U55462 ( .A(n46075), .B(n46078), .Z(n46079) );
  AND U55463 ( .A(n46080), .B(n46081), .Z(n46078) );
  NANDN U55464 ( .A(n46082), .B(n46083), .Z(n46081) );
  NANDN U55465 ( .A(n46084), .B(n46085), .Z(n46083) );
  NANDN U55466 ( .A(n46085), .B(n46084), .Z(n46080) );
  NAND U55467 ( .A(n46086), .B(n46087), .Z(n46075) );
  NANDN U55468 ( .A(n46088), .B(n46089), .Z(n46087) );
  OR U55469 ( .A(n46090), .B(n46091), .Z(n46089) );
  NAND U55470 ( .A(n46091), .B(n46090), .Z(n46086) );
  AND U55471 ( .A(n46092), .B(n46093), .Z(n46077) );
  NANDN U55472 ( .A(n46094), .B(n46095), .Z(n46093) );
  NANDN U55473 ( .A(n46096), .B(n46097), .Z(n46095) );
  NANDN U55474 ( .A(n46097), .B(n46096), .Z(n46092) );
  XOR U55475 ( .A(n46091), .B(n46098), .Z(N61309) );
  XOR U55476 ( .A(n46088), .B(n46090), .Z(n46098) );
  XNOR U55477 ( .A(n46084), .B(n46099), .Z(n46090) );
  XNOR U55478 ( .A(n46082), .B(n46085), .Z(n46099) );
  NAND U55479 ( .A(n46100), .B(n46101), .Z(n46085) );
  NAND U55480 ( .A(n46102), .B(n46103), .Z(n46101) );
  OR U55481 ( .A(n46104), .B(n46105), .Z(n46102) );
  NANDN U55482 ( .A(n46106), .B(n46104), .Z(n46100) );
  IV U55483 ( .A(n46105), .Z(n46106) );
  NAND U55484 ( .A(n46107), .B(n46108), .Z(n46082) );
  NAND U55485 ( .A(n46109), .B(n46110), .Z(n46108) );
  NANDN U55486 ( .A(n46111), .B(n46112), .Z(n46109) );
  NANDN U55487 ( .A(n46112), .B(n46111), .Z(n46107) );
  AND U55488 ( .A(n46113), .B(n46114), .Z(n46084) );
  NAND U55489 ( .A(n46115), .B(n46116), .Z(n46114) );
  OR U55490 ( .A(n46117), .B(n46118), .Z(n46115) );
  NANDN U55491 ( .A(n46119), .B(n46117), .Z(n46113) );
  NAND U55492 ( .A(n46120), .B(n46121), .Z(n46088) );
  NANDN U55493 ( .A(n46122), .B(n46123), .Z(n46121) );
  OR U55494 ( .A(n46124), .B(n46125), .Z(n46123) );
  NANDN U55495 ( .A(n46126), .B(n46124), .Z(n46120) );
  IV U55496 ( .A(n46125), .Z(n46126) );
  XNOR U55497 ( .A(n46096), .B(n46127), .Z(n46091) );
  XNOR U55498 ( .A(n46094), .B(n46097), .Z(n46127) );
  NAND U55499 ( .A(n46128), .B(n46129), .Z(n46097) );
  NAND U55500 ( .A(n46130), .B(n46131), .Z(n46129) );
  OR U55501 ( .A(n46132), .B(n46133), .Z(n46130) );
  NANDN U55502 ( .A(n46134), .B(n46132), .Z(n46128) );
  IV U55503 ( .A(n46133), .Z(n46134) );
  NAND U55504 ( .A(n46135), .B(n46136), .Z(n46094) );
  NAND U55505 ( .A(n46137), .B(n46138), .Z(n46136) );
  NANDN U55506 ( .A(n46139), .B(n46140), .Z(n46137) );
  NANDN U55507 ( .A(n46140), .B(n46139), .Z(n46135) );
  AND U55508 ( .A(n46141), .B(n46142), .Z(n46096) );
  NAND U55509 ( .A(n46143), .B(n46144), .Z(n46142) );
  OR U55510 ( .A(n46145), .B(n46146), .Z(n46143) );
  NANDN U55511 ( .A(n46147), .B(n46145), .Z(n46141) );
  XNOR U55512 ( .A(n46122), .B(n46148), .Z(N61308) );
  XOR U55513 ( .A(n46124), .B(n46125), .Z(n46148) );
  XNOR U55514 ( .A(n46138), .B(n46149), .Z(n46125) );
  XOR U55515 ( .A(n46139), .B(n46140), .Z(n46149) );
  XOR U55516 ( .A(n46145), .B(n46150), .Z(n46140) );
  XOR U55517 ( .A(n46144), .B(n46147), .Z(n46150) );
  IV U55518 ( .A(n46146), .Z(n46147) );
  NAND U55519 ( .A(n46151), .B(n46152), .Z(n46146) );
  OR U55520 ( .A(n46153), .B(n46154), .Z(n46152) );
  OR U55521 ( .A(n46155), .B(n46156), .Z(n46151) );
  NAND U55522 ( .A(n46157), .B(n46158), .Z(n46144) );
  OR U55523 ( .A(n46159), .B(n46160), .Z(n46158) );
  OR U55524 ( .A(n46161), .B(n46162), .Z(n46157) );
  NOR U55525 ( .A(n46163), .B(n46164), .Z(n46145) );
  ANDN U55526 ( .B(n46165), .A(n46166), .Z(n46139) );
  XNOR U55527 ( .A(n46132), .B(n46167), .Z(n46138) );
  XNOR U55528 ( .A(n46131), .B(n46133), .Z(n46167) );
  NAND U55529 ( .A(n46168), .B(n46169), .Z(n46133) );
  OR U55530 ( .A(n46170), .B(n46171), .Z(n46169) );
  OR U55531 ( .A(n46172), .B(n46173), .Z(n46168) );
  NAND U55532 ( .A(n46174), .B(n46175), .Z(n46131) );
  OR U55533 ( .A(n46176), .B(n46177), .Z(n46175) );
  OR U55534 ( .A(n46178), .B(n46179), .Z(n46174) );
  ANDN U55535 ( .B(n46180), .A(n46181), .Z(n46132) );
  IV U55536 ( .A(n46182), .Z(n46180) );
  ANDN U55537 ( .B(n46183), .A(n46184), .Z(n46124) );
  XOR U55538 ( .A(n46110), .B(n46185), .Z(n46122) );
  XOR U55539 ( .A(n46111), .B(n46112), .Z(n46185) );
  XOR U55540 ( .A(n46117), .B(n46186), .Z(n46112) );
  XOR U55541 ( .A(n46116), .B(n46119), .Z(n46186) );
  IV U55542 ( .A(n46118), .Z(n46119) );
  NAND U55543 ( .A(n46187), .B(n46188), .Z(n46118) );
  OR U55544 ( .A(n46189), .B(n46190), .Z(n46188) );
  OR U55545 ( .A(n46191), .B(n46192), .Z(n46187) );
  NAND U55546 ( .A(n46193), .B(n46194), .Z(n46116) );
  OR U55547 ( .A(n46195), .B(n46196), .Z(n46194) );
  OR U55548 ( .A(n46197), .B(n46198), .Z(n46193) );
  NOR U55549 ( .A(n46199), .B(n46200), .Z(n46117) );
  ANDN U55550 ( .B(n46201), .A(n46202), .Z(n46111) );
  IV U55551 ( .A(n46203), .Z(n46201) );
  XNOR U55552 ( .A(n46104), .B(n46204), .Z(n46110) );
  XNOR U55553 ( .A(n46103), .B(n46105), .Z(n46204) );
  NAND U55554 ( .A(n46205), .B(n46206), .Z(n46105) );
  OR U55555 ( .A(n46207), .B(n46208), .Z(n46206) );
  OR U55556 ( .A(n46209), .B(n46210), .Z(n46205) );
  NAND U55557 ( .A(n46211), .B(n46212), .Z(n46103) );
  OR U55558 ( .A(n46213), .B(n46214), .Z(n46212) );
  OR U55559 ( .A(n46215), .B(n46216), .Z(n46211) );
  ANDN U55560 ( .B(n46217), .A(n46218), .Z(n46104) );
  IV U55561 ( .A(n46219), .Z(n46217) );
  XNOR U55562 ( .A(n46184), .B(n46183), .Z(N61307) );
  XOR U55563 ( .A(n46203), .B(n46202), .Z(n46183) );
  XNOR U55564 ( .A(n46218), .B(n46219), .Z(n46202) );
  XNOR U55565 ( .A(n46213), .B(n46214), .Z(n46219) );
  XNOR U55566 ( .A(n46215), .B(n46216), .Z(n46214) );
  XNOR U55567 ( .A(y[1333]), .B(x[1333]), .Z(n46216) );
  XNOR U55568 ( .A(y[1334]), .B(x[1334]), .Z(n46215) );
  XNOR U55569 ( .A(y[1332]), .B(x[1332]), .Z(n46213) );
  XNOR U55570 ( .A(n46207), .B(n46208), .Z(n46218) );
  XNOR U55571 ( .A(y[1329]), .B(x[1329]), .Z(n46208) );
  XNOR U55572 ( .A(n46209), .B(n46210), .Z(n46207) );
  XNOR U55573 ( .A(y[1330]), .B(x[1330]), .Z(n46210) );
  XNOR U55574 ( .A(y[1331]), .B(x[1331]), .Z(n46209) );
  XNOR U55575 ( .A(n46200), .B(n46199), .Z(n46203) );
  XNOR U55576 ( .A(n46195), .B(n46196), .Z(n46199) );
  XNOR U55577 ( .A(y[1326]), .B(x[1326]), .Z(n46196) );
  XNOR U55578 ( .A(n46197), .B(n46198), .Z(n46195) );
  XNOR U55579 ( .A(y[1327]), .B(x[1327]), .Z(n46198) );
  XNOR U55580 ( .A(y[1328]), .B(x[1328]), .Z(n46197) );
  XNOR U55581 ( .A(n46189), .B(n46190), .Z(n46200) );
  XNOR U55582 ( .A(y[1323]), .B(x[1323]), .Z(n46190) );
  XNOR U55583 ( .A(n46191), .B(n46192), .Z(n46189) );
  XNOR U55584 ( .A(y[1324]), .B(x[1324]), .Z(n46192) );
  XNOR U55585 ( .A(y[1325]), .B(x[1325]), .Z(n46191) );
  XOR U55586 ( .A(n46165), .B(n46166), .Z(n46184) );
  XNOR U55587 ( .A(n46181), .B(n46182), .Z(n46166) );
  XNOR U55588 ( .A(n46176), .B(n46177), .Z(n46182) );
  XNOR U55589 ( .A(n46178), .B(n46179), .Z(n46177) );
  XNOR U55590 ( .A(y[1321]), .B(x[1321]), .Z(n46179) );
  XNOR U55591 ( .A(y[1322]), .B(x[1322]), .Z(n46178) );
  XNOR U55592 ( .A(y[1320]), .B(x[1320]), .Z(n46176) );
  XNOR U55593 ( .A(n46170), .B(n46171), .Z(n46181) );
  XNOR U55594 ( .A(y[1317]), .B(x[1317]), .Z(n46171) );
  XNOR U55595 ( .A(n46172), .B(n46173), .Z(n46170) );
  XNOR U55596 ( .A(y[1318]), .B(x[1318]), .Z(n46173) );
  XNOR U55597 ( .A(y[1319]), .B(x[1319]), .Z(n46172) );
  XOR U55598 ( .A(n46164), .B(n46163), .Z(n46165) );
  XNOR U55599 ( .A(n46159), .B(n46160), .Z(n46163) );
  XNOR U55600 ( .A(y[1314]), .B(x[1314]), .Z(n46160) );
  XNOR U55601 ( .A(n46161), .B(n46162), .Z(n46159) );
  XNOR U55602 ( .A(y[1315]), .B(x[1315]), .Z(n46162) );
  XNOR U55603 ( .A(y[1316]), .B(x[1316]), .Z(n46161) );
  XNOR U55604 ( .A(n46153), .B(n46154), .Z(n46164) );
  XNOR U55605 ( .A(y[1311]), .B(x[1311]), .Z(n46154) );
  XNOR U55606 ( .A(n46155), .B(n46156), .Z(n46153) );
  XNOR U55607 ( .A(y[1312]), .B(x[1312]), .Z(n46156) );
  XNOR U55608 ( .A(y[1313]), .B(x[1313]), .Z(n46155) );
  NAND U55609 ( .A(n46220), .B(n46221), .Z(N61298) );
  NANDN U55610 ( .A(n46222), .B(n46223), .Z(n46221) );
  OR U55611 ( .A(n46224), .B(n46225), .Z(n46223) );
  NAND U55612 ( .A(n46224), .B(n46225), .Z(n46220) );
  XOR U55613 ( .A(n46224), .B(n46226), .Z(N61297) );
  XNOR U55614 ( .A(n46222), .B(n46225), .Z(n46226) );
  AND U55615 ( .A(n46227), .B(n46228), .Z(n46225) );
  NANDN U55616 ( .A(n46229), .B(n46230), .Z(n46228) );
  NANDN U55617 ( .A(n46231), .B(n46232), .Z(n46230) );
  NANDN U55618 ( .A(n46232), .B(n46231), .Z(n46227) );
  NAND U55619 ( .A(n46233), .B(n46234), .Z(n46222) );
  NANDN U55620 ( .A(n46235), .B(n46236), .Z(n46234) );
  OR U55621 ( .A(n46237), .B(n46238), .Z(n46236) );
  NAND U55622 ( .A(n46238), .B(n46237), .Z(n46233) );
  AND U55623 ( .A(n46239), .B(n46240), .Z(n46224) );
  NANDN U55624 ( .A(n46241), .B(n46242), .Z(n46240) );
  NANDN U55625 ( .A(n46243), .B(n46244), .Z(n46242) );
  NANDN U55626 ( .A(n46244), .B(n46243), .Z(n46239) );
  XOR U55627 ( .A(n46238), .B(n46245), .Z(N61296) );
  XOR U55628 ( .A(n46235), .B(n46237), .Z(n46245) );
  XNOR U55629 ( .A(n46231), .B(n46246), .Z(n46237) );
  XNOR U55630 ( .A(n46229), .B(n46232), .Z(n46246) );
  NAND U55631 ( .A(n46247), .B(n46248), .Z(n46232) );
  NAND U55632 ( .A(n46249), .B(n46250), .Z(n46248) );
  OR U55633 ( .A(n46251), .B(n46252), .Z(n46249) );
  NANDN U55634 ( .A(n46253), .B(n46251), .Z(n46247) );
  IV U55635 ( .A(n46252), .Z(n46253) );
  NAND U55636 ( .A(n46254), .B(n46255), .Z(n46229) );
  NAND U55637 ( .A(n46256), .B(n46257), .Z(n46255) );
  NANDN U55638 ( .A(n46258), .B(n46259), .Z(n46256) );
  NANDN U55639 ( .A(n46259), .B(n46258), .Z(n46254) );
  AND U55640 ( .A(n46260), .B(n46261), .Z(n46231) );
  NAND U55641 ( .A(n46262), .B(n46263), .Z(n46261) );
  OR U55642 ( .A(n46264), .B(n46265), .Z(n46262) );
  NANDN U55643 ( .A(n46266), .B(n46264), .Z(n46260) );
  NAND U55644 ( .A(n46267), .B(n46268), .Z(n46235) );
  NANDN U55645 ( .A(n46269), .B(n46270), .Z(n46268) );
  OR U55646 ( .A(n46271), .B(n46272), .Z(n46270) );
  NANDN U55647 ( .A(n46273), .B(n46271), .Z(n46267) );
  IV U55648 ( .A(n46272), .Z(n46273) );
  XNOR U55649 ( .A(n46243), .B(n46274), .Z(n46238) );
  XNOR U55650 ( .A(n46241), .B(n46244), .Z(n46274) );
  NAND U55651 ( .A(n46275), .B(n46276), .Z(n46244) );
  NAND U55652 ( .A(n46277), .B(n46278), .Z(n46276) );
  OR U55653 ( .A(n46279), .B(n46280), .Z(n46277) );
  NANDN U55654 ( .A(n46281), .B(n46279), .Z(n46275) );
  IV U55655 ( .A(n46280), .Z(n46281) );
  NAND U55656 ( .A(n46282), .B(n46283), .Z(n46241) );
  NAND U55657 ( .A(n46284), .B(n46285), .Z(n46283) );
  NANDN U55658 ( .A(n46286), .B(n46287), .Z(n46284) );
  NANDN U55659 ( .A(n46287), .B(n46286), .Z(n46282) );
  AND U55660 ( .A(n46288), .B(n46289), .Z(n46243) );
  NAND U55661 ( .A(n46290), .B(n46291), .Z(n46289) );
  OR U55662 ( .A(n46292), .B(n46293), .Z(n46290) );
  NANDN U55663 ( .A(n46294), .B(n46292), .Z(n46288) );
  XNOR U55664 ( .A(n46269), .B(n46295), .Z(N61295) );
  XOR U55665 ( .A(n46271), .B(n46272), .Z(n46295) );
  XNOR U55666 ( .A(n46285), .B(n46296), .Z(n46272) );
  XOR U55667 ( .A(n46286), .B(n46287), .Z(n46296) );
  XOR U55668 ( .A(n46292), .B(n46297), .Z(n46287) );
  XOR U55669 ( .A(n46291), .B(n46294), .Z(n46297) );
  IV U55670 ( .A(n46293), .Z(n46294) );
  NAND U55671 ( .A(n46298), .B(n46299), .Z(n46293) );
  OR U55672 ( .A(n46300), .B(n46301), .Z(n46299) );
  OR U55673 ( .A(n46302), .B(n46303), .Z(n46298) );
  NAND U55674 ( .A(n46304), .B(n46305), .Z(n46291) );
  OR U55675 ( .A(n46306), .B(n46307), .Z(n46305) );
  OR U55676 ( .A(n46308), .B(n46309), .Z(n46304) );
  NOR U55677 ( .A(n46310), .B(n46311), .Z(n46292) );
  ANDN U55678 ( .B(n46312), .A(n46313), .Z(n46286) );
  XNOR U55679 ( .A(n46279), .B(n46314), .Z(n46285) );
  XNOR U55680 ( .A(n46278), .B(n46280), .Z(n46314) );
  NAND U55681 ( .A(n46315), .B(n46316), .Z(n46280) );
  OR U55682 ( .A(n46317), .B(n46318), .Z(n46316) );
  OR U55683 ( .A(n46319), .B(n46320), .Z(n46315) );
  NAND U55684 ( .A(n46321), .B(n46322), .Z(n46278) );
  OR U55685 ( .A(n46323), .B(n46324), .Z(n46322) );
  OR U55686 ( .A(n46325), .B(n46326), .Z(n46321) );
  ANDN U55687 ( .B(n46327), .A(n46328), .Z(n46279) );
  IV U55688 ( .A(n46329), .Z(n46327) );
  ANDN U55689 ( .B(n46330), .A(n46331), .Z(n46271) );
  XOR U55690 ( .A(n46257), .B(n46332), .Z(n46269) );
  XOR U55691 ( .A(n46258), .B(n46259), .Z(n46332) );
  XOR U55692 ( .A(n46264), .B(n46333), .Z(n46259) );
  XOR U55693 ( .A(n46263), .B(n46266), .Z(n46333) );
  IV U55694 ( .A(n46265), .Z(n46266) );
  NAND U55695 ( .A(n46334), .B(n46335), .Z(n46265) );
  OR U55696 ( .A(n46336), .B(n46337), .Z(n46335) );
  OR U55697 ( .A(n46338), .B(n46339), .Z(n46334) );
  NAND U55698 ( .A(n46340), .B(n46341), .Z(n46263) );
  OR U55699 ( .A(n46342), .B(n46343), .Z(n46341) );
  OR U55700 ( .A(n46344), .B(n46345), .Z(n46340) );
  NOR U55701 ( .A(n46346), .B(n46347), .Z(n46264) );
  ANDN U55702 ( .B(n46348), .A(n46349), .Z(n46258) );
  IV U55703 ( .A(n46350), .Z(n46348) );
  XNOR U55704 ( .A(n46251), .B(n46351), .Z(n46257) );
  XNOR U55705 ( .A(n46250), .B(n46252), .Z(n46351) );
  NAND U55706 ( .A(n46352), .B(n46353), .Z(n46252) );
  OR U55707 ( .A(n46354), .B(n46355), .Z(n46353) );
  OR U55708 ( .A(n46356), .B(n46357), .Z(n46352) );
  NAND U55709 ( .A(n46358), .B(n46359), .Z(n46250) );
  OR U55710 ( .A(n46360), .B(n46361), .Z(n46359) );
  OR U55711 ( .A(n46362), .B(n46363), .Z(n46358) );
  ANDN U55712 ( .B(n46364), .A(n46365), .Z(n46251) );
  IV U55713 ( .A(n46366), .Z(n46364) );
  XNOR U55714 ( .A(n46331), .B(n46330), .Z(N61294) );
  XOR U55715 ( .A(n46350), .B(n46349), .Z(n46330) );
  XNOR U55716 ( .A(n46365), .B(n46366), .Z(n46349) );
  XNOR U55717 ( .A(n46360), .B(n46361), .Z(n46366) );
  XNOR U55718 ( .A(n46362), .B(n46363), .Z(n46361) );
  XNOR U55719 ( .A(y[1309]), .B(x[1309]), .Z(n46363) );
  XNOR U55720 ( .A(y[1310]), .B(x[1310]), .Z(n46362) );
  XNOR U55721 ( .A(y[1308]), .B(x[1308]), .Z(n46360) );
  XNOR U55722 ( .A(n46354), .B(n46355), .Z(n46365) );
  XNOR U55723 ( .A(y[1305]), .B(x[1305]), .Z(n46355) );
  XNOR U55724 ( .A(n46356), .B(n46357), .Z(n46354) );
  XNOR U55725 ( .A(y[1306]), .B(x[1306]), .Z(n46357) );
  XNOR U55726 ( .A(y[1307]), .B(x[1307]), .Z(n46356) );
  XNOR U55727 ( .A(n46347), .B(n46346), .Z(n46350) );
  XNOR U55728 ( .A(n46342), .B(n46343), .Z(n46346) );
  XNOR U55729 ( .A(y[1302]), .B(x[1302]), .Z(n46343) );
  XNOR U55730 ( .A(n46344), .B(n46345), .Z(n46342) );
  XNOR U55731 ( .A(y[1303]), .B(x[1303]), .Z(n46345) );
  XNOR U55732 ( .A(y[1304]), .B(x[1304]), .Z(n46344) );
  XNOR U55733 ( .A(n46336), .B(n46337), .Z(n46347) );
  XNOR U55734 ( .A(y[1299]), .B(x[1299]), .Z(n46337) );
  XNOR U55735 ( .A(n46338), .B(n46339), .Z(n46336) );
  XNOR U55736 ( .A(y[1300]), .B(x[1300]), .Z(n46339) );
  XNOR U55737 ( .A(y[1301]), .B(x[1301]), .Z(n46338) );
  XOR U55738 ( .A(n46312), .B(n46313), .Z(n46331) );
  XNOR U55739 ( .A(n46328), .B(n46329), .Z(n46313) );
  XNOR U55740 ( .A(n46323), .B(n46324), .Z(n46329) );
  XNOR U55741 ( .A(n46325), .B(n46326), .Z(n46324) );
  XNOR U55742 ( .A(y[1297]), .B(x[1297]), .Z(n46326) );
  XNOR U55743 ( .A(y[1298]), .B(x[1298]), .Z(n46325) );
  XNOR U55744 ( .A(y[1296]), .B(x[1296]), .Z(n46323) );
  XNOR U55745 ( .A(n46317), .B(n46318), .Z(n46328) );
  XNOR U55746 ( .A(y[1293]), .B(x[1293]), .Z(n46318) );
  XNOR U55747 ( .A(n46319), .B(n46320), .Z(n46317) );
  XNOR U55748 ( .A(y[1294]), .B(x[1294]), .Z(n46320) );
  XNOR U55749 ( .A(y[1295]), .B(x[1295]), .Z(n46319) );
  XOR U55750 ( .A(n46311), .B(n46310), .Z(n46312) );
  XNOR U55751 ( .A(n46306), .B(n46307), .Z(n46310) );
  XNOR U55752 ( .A(y[1290]), .B(x[1290]), .Z(n46307) );
  XNOR U55753 ( .A(n46308), .B(n46309), .Z(n46306) );
  XNOR U55754 ( .A(y[1291]), .B(x[1291]), .Z(n46309) );
  XNOR U55755 ( .A(y[1292]), .B(x[1292]), .Z(n46308) );
  XNOR U55756 ( .A(n46300), .B(n46301), .Z(n46311) );
  XNOR U55757 ( .A(y[1287]), .B(x[1287]), .Z(n46301) );
  XNOR U55758 ( .A(n46302), .B(n46303), .Z(n46300) );
  XNOR U55759 ( .A(y[1288]), .B(x[1288]), .Z(n46303) );
  XNOR U55760 ( .A(y[1289]), .B(x[1289]), .Z(n46302) );
  NAND U55761 ( .A(n46367), .B(n46368), .Z(N61285) );
  NANDN U55762 ( .A(n46369), .B(n46370), .Z(n46368) );
  OR U55763 ( .A(n46371), .B(n46372), .Z(n46370) );
  NAND U55764 ( .A(n46371), .B(n46372), .Z(n46367) );
  XOR U55765 ( .A(n46371), .B(n46373), .Z(N61284) );
  XNOR U55766 ( .A(n46369), .B(n46372), .Z(n46373) );
  AND U55767 ( .A(n46374), .B(n46375), .Z(n46372) );
  NANDN U55768 ( .A(n46376), .B(n46377), .Z(n46375) );
  NANDN U55769 ( .A(n46378), .B(n46379), .Z(n46377) );
  NANDN U55770 ( .A(n46379), .B(n46378), .Z(n46374) );
  NAND U55771 ( .A(n46380), .B(n46381), .Z(n46369) );
  NANDN U55772 ( .A(n46382), .B(n46383), .Z(n46381) );
  OR U55773 ( .A(n46384), .B(n46385), .Z(n46383) );
  NAND U55774 ( .A(n46385), .B(n46384), .Z(n46380) );
  AND U55775 ( .A(n46386), .B(n46387), .Z(n46371) );
  NANDN U55776 ( .A(n46388), .B(n46389), .Z(n46387) );
  NANDN U55777 ( .A(n46390), .B(n46391), .Z(n46389) );
  NANDN U55778 ( .A(n46391), .B(n46390), .Z(n46386) );
  XOR U55779 ( .A(n46385), .B(n46392), .Z(N61283) );
  XOR U55780 ( .A(n46382), .B(n46384), .Z(n46392) );
  XNOR U55781 ( .A(n46378), .B(n46393), .Z(n46384) );
  XNOR U55782 ( .A(n46376), .B(n46379), .Z(n46393) );
  NAND U55783 ( .A(n46394), .B(n46395), .Z(n46379) );
  NAND U55784 ( .A(n46396), .B(n46397), .Z(n46395) );
  OR U55785 ( .A(n46398), .B(n46399), .Z(n46396) );
  NANDN U55786 ( .A(n46400), .B(n46398), .Z(n46394) );
  IV U55787 ( .A(n46399), .Z(n46400) );
  NAND U55788 ( .A(n46401), .B(n46402), .Z(n46376) );
  NAND U55789 ( .A(n46403), .B(n46404), .Z(n46402) );
  NANDN U55790 ( .A(n46405), .B(n46406), .Z(n46403) );
  NANDN U55791 ( .A(n46406), .B(n46405), .Z(n46401) );
  AND U55792 ( .A(n46407), .B(n46408), .Z(n46378) );
  NAND U55793 ( .A(n46409), .B(n46410), .Z(n46408) );
  OR U55794 ( .A(n46411), .B(n46412), .Z(n46409) );
  NANDN U55795 ( .A(n46413), .B(n46411), .Z(n46407) );
  NAND U55796 ( .A(n46414), .B(n46415), .Z(n46382) );
  NANDN U55797 ( .A(n46416), .B(n46417), .Z(n46415) );
  OR U55798 ( .A(n46418), .B(n46419), .Z(n46417) );
  NANDN U55799 ( .A(n46420), .B(n46418), .Z(n46414) );
  IV U55800 ( .A(n46419), .Z(n46420) );
  XNOR U55801 ( .A(n46390), .B(n46421), .Z(n46385) );
  XNOR U55802 ( .A(n46388), .B(n46391), .Z(n46421) );
  NAND U55803 ( .A(n46422), .B(n46423), .Z(n46391) );
  NAND U55804 ( .A(n46424), .B(n46425), .Z(n46423) );
  OR U55805 ( .A(n46426), .B(n46427), .Z(n46424) );
  NANDN U55806 ( .A(n46428), .B(n46426), .Z(n46422) );
  IV U55807 ( .A(n46427), .Z(n46428) );
  NAND U55808 ( .A(n46429), .B(n46430), .Z(n46388) );
  NAND U55809 ( .A(n46431), .B(n46432), .Z(n46430) );
  NANDN U55810 ( .A(n46433), .B(n46434), .Z(n46431) );
  NANDN U55811 ( .A(n46434), .B(n46433), .Z(n46429) );
  AND U55812 ( .A(n46435), .B(n46436), .Z(n46390) );
  NAND U55813 ( .A(n46437), .B(n46438), .Z(n46436) );
  OR U55814 ( .A(n46439), .B(n46440), .Z(n46437) );
  NANDN U55815 ( .A(n46441), .B(n46439), .Z(n46435) );
  XNOR U55816 ( .A(n46416), .B(n46442), .Z(N61282) );
  XOR U55817 ( .A(n46418), .B(n46419), .Z(n46442) );
  XNOR U55818 ( .A(n46432), .B(n46443), .Z(n46419) );
  XOR U55819 ( .A(n46433), .B(n46434), .Z(n46443) );
  XOR U55820 ( .A(n46439), .B(n46444), .Z(n46434) );
  XOR U55821 ( .A(n46438), .B(n46441), .Z(n46444) );
  IV U55822 ( .A(n46440), .Z(n46441) );
  NAND U55823 ( .A(n46445), .B(n46446), .Z(n46440) );
  OR U55824 ( .A(n46447), .B(n46448), .Z(n46446) );
  OR U55825 ( .A(n46449), .B(n46450), .Z(n46445) );
  NAND U55826 ( .A(n46451), .B(n46452), .Z(n46438) );
  OR U55827 ( .A(n46453), .B(n46454), .Z(n46452) );
  OR U55828 ( .A(n46455), .B(n46456), .Z(n46451) );
  NOR U55829 ( .A(n46457), .B(n46458), .Z(n46439) );
  ANDN U55830 ( .B(n46459), .A(n46460), .Z(n46433) );
  XNOR U55831 ( .A(n46426), .B(n46461), .Z(n46432) );
  XNOR U55832 ( .A(n46425), .B(n46427), .Z(n46461) );
  NAND U55833 ( .A(n46462), .B(n46463), .Z(n46427) );
  OR U55834 ( .A(n46464), .B(n46465), .Z(n46463) );
  OR U55835 ( .A(n46466), .B(n46467), .Z(n46462) );
  NAND U55836 ( .A(n46468), .B(n46469), .Z(n46425) );
  OR U55837 ( .A(n46470), .B(n46471), .Z(n46469) );
  OR U55838 ( .A(n46472), .B(n46473), .Z(n46468) );
  ANDN U55839 ( .B(n46474), .A(n46475), .Z(n46426) );
  IV U55840 ( .A(n46476), .Z(n46474) );
  ANDN U55841 ( .B(n46477), .A(n46478), .Z(n46418) );
  XOR U55842 ( .A(n46404), .B(n46479), .Z(n46416) );
  XOR U55843 ( .A(n46405), .B(n46406), .Z(n46479) );
  XOR U55844 ( .A(n46411), .B(n46480), .Z(n46406) );
  XOR U55845 ( .A(n46410), .B(n46413), .Z(n46480) );
  IV U55846 ( .A(n46412), .Z(n46413) );
  NAND U55847 ( .A(n46481), .B(n46482), .Z(n46412) );
  OR U55848 ( .A(n46483), .B(n46484), .Z(n46482) );
  OR U55849 ( .A(n46485), .B(n46486), .Z(n46481) );
  NAND U55850 ( .A(n46487), .B(n46488), .Z(n46410) );
  OR U55851 ( .A(n46489), .B(n46490), .Z(n46488) );
  OR U55852 ( .A(n46491), .B(n46492), .Z(n46487) );
  NOR U55853 ( .A(n46493), .B(n46494), .Z(n46411) );
  ANDN U55854 ( .B(n46495), .A(n46496), .Z(n46405) );
  IV U55855 ( .A(n46497), .Z(n46495) );
  XNOR U55856 ( .A(n46398), .B(n46498), .Z(n46404) );
  XNOR U55857 ( .A(n46397), .B(n46399), .Z(n46498) );
  NAND U55858 ( .A(n46499), .B(n46500), .Z(n46399) );
  OR U55859 ( .A(n46501), .B(n46502), .Z(n46500) );
  OR U55860 ( .A(n46503), .B(n46504), .Z(n46499) );
  NAND U55861 ( .A(n46505), .B(n46506), .Z(n46397) );
  OR U55862 ( .A(n46507), .B(n46508), .Z(n46506) );
  OR U55863 ( .A(n46509), .B(n46510), .Z(n46505) );
  ANDN U55864 ( .B(n46511), .A(n46512), .Z(n46398) );
  IV U55865 ( .A(n46513), .Z(n46511) );
  XNOR U55866 ( .A(n46478), .B(n46477), .Z(N61281) );
  XOR U55867 ( .A(n46497), .B(n46496), .Z(n46477) );
  XNOR U55868 ( .A(n46512), .B(n46513), .Z(n46496) );
  XNOR U55869 ( .A(n46507), .B(n46508), .Z(n46513) );
  XNOR U55870 ( .A(n46509), .B(n46510), .Z(n46508) );
  XNOR U55871 ( .A(y[1285]), .B(x[1285]), .Z(n46510) );
  XNOR U55872 ( .A(y[1286]), .B(x[1286]), .Z(n46509) );
  XNOR U55873 ( .A(y[1284]), .B(x[1284]), .Z(n46507) );
  XNOR U55874 ( .A(n46501), .B(n46502), .Z(n46512) );
  XNOR U55875 ( .A(y[1281]), .B(x[1281]), .Z(n46502) );
  XNOR U55876 ( .A(n46503), .B(n46504), .Z(n46501) );
  XNOR U55877 ( .A(y[1282]), .B(x[1282]), .Z(n46504) );
  XNOR U55878 ( .A(y[1283]), .B(x[1283]), .Z(n46503) );
  XNOR U55879 ( .A(n46494), .B(n46493), .Z(n46497) );
  XNOR U55880 ( .A(n46489), .B(n46490), .Z(n46493) );
  XNOR U55881 ( .A(y[1278]), .B(x[1278]), .Z(n46490) );
  XNOR U55882 ( .A(n46491), .B(n46492), .Z(n46489) );
  XNOR U55883 ( .A(y[1279]), .B(x[1279]), .Z(n46492) );
  XNOR U55884 ( .A(y[1280]), .B(x[1280]), .Z(n46491) );
  XNOR U55885 ( .A(n46483), .B(n46484), .Z(n46494) );
  XNOR U55886 ( .A(y[1275]), .B(x[1275]), .Z(n46484) );
  XNOR U55887 ( .A(n46485), .B(n46486), .Z(n46483) );
  XNOR U55888 ( .A(y[1276]), .B(x[1276]), .Z(n46486) );
  XNOR U55889 ( .A(y[1277]), .B(x[1277]), .Z(n46485) );
  XOR U55890 ( .A(n46459), .B(n46460), .Z(n46478) );
  XNOR U55891 ( .A(n46475), .B(n46476), .Z(n46460) );
  XNOR U55892 ( .A(n46470), .B(n46471), .Z(n46476) );
  XNOR U55893 ( .A(n46472), .B(n46473), .Z(n46471) );
  XNOR U55894 ( .A(y[1273]), .B(x[1273]), .Z(n46473) );
  XNOR U55895 ( .A(y[1274]), .B(x[1274]), .Z(n46472) );
  XNOR U55896 ( .A(y[1272]), .B(x[1272]), .Z(n46470) );
  XNOR U55897 ( .A(n46464), .B(n46465), .Z(n46475) );
  XNOR U55898 ( .A(y[1269]), .B(x[1269]), .Z(n46465) );
  XNOR U55899 ( .A(n46466), .B(n46467), .Z(n46464) );
  XNOR U55900 ( .A(y[1270]), .B(x[1270]), .Z(n46467) );
  XNOR U55901 ( .A(y[1271]), .B(x[1271]), .Z(n46466) );
  XOR U55902 ( .A(n46458), .B(n46457), .Z(n46459) );
  XNOR U55903 ( .A(n46453), .B(n46454), .Z(n46457) );
  XNOR U55904 ( .A(y[1266]), .B(x[1266]), .Z(n46454) );
  XNOR U55905 ( .A(n46455), .B(n46456), .Z(n46453) );
  XNOR U55906 ( .A(y[1267]), .B(x[1267]), .Z(n46456) );
  XNOR U55907 ( .A(y[1268]), .B(x[1268]), .Z(n46455) );
  XNOR U55908 ( .A(n46447), .B(n46448), .Z(n46458) );
  XNOR U55909 ( .A(y[1263]), .B(x[1263]), .Z(n46448) );
  XNOR U55910 ( .A(n46449), .B(n46450), .Z(n46447) );
  XNOR U55911 ( .A(y[1264]), .B(x[1264]), .Z(n46450) );
  XNOR U55912 ( .A(y[1265]), .B(x[1265]), .Z(n46449) );
  NAND U55913 ( .A(n46514), .B(n46515), .Z(N61272) );
  NANDN U55914 ( .A(n46516), .B(n46517), .Z(n46515) );
  OR U55915 ( .A(n46518), .B(n46519), .Z(n46517) );
  NAND U55916 ( .A(n46518), .B(n46519), .Z(n46514) );
  XOR U55917 ( .A(n46518), .B(n46520), .Z(N61271) );
  XNOR U55918 ( .A(n46516), .B(n46519), .Z(n46520) );
  AND U55919 ( .A(n46521), .B(n46522), .Z(n46519) );
  NANDN U55920 ( .A(n46523), .B(n46524), .Z(n46522) );
  NANDN U55921 ( .A(n46525), .B(n46526), .Z(n46524) );
  NANDN U55922 ( .A(n46526), .B(n46525), .Z(n46521) );
  NAND U55923 ( .A(n46527), .B(n46528), .Z(n46516) );
  NANDN U55924 ( .A(n46529), .B(n46530), .Z(n46528) );
  OR U55925 ( .A(n46531), .B(n46532), .Z(n46530) );
  NAND U55926 ( .A(n46532), .B(n46531), .Z(n46527) );
  AND U55927 ( .A(n46533), .B(n46534), .Z(n46518) );
  NANDN U55928 ( .A(n46535), .B(n46536), .Z(n46534) );
  NANDN U55929 ( .A(n46537), .B(n46538), .Z(n46536) );
  NANDN U55930 ( .A(n46538), .B(n46537), .Z(n46533) );
  XOR U55931 ( .A(n46532), .B(n46539), .Z(N61270) );
  XOR U55932 ( .A(n46529), .B(n46531), .Z(n46539) );
  XNOR U55933 ( .A(n46525), .B(n46540), .Z(n46531) );
  XNOR U55934 ( .A(n46523), .B(n46526), .Z(n46540) );
  NAND U55935 ( .A(n46541), .B(n46542), .Z(n46526) );
  NAND U55936 ( .A(n46543), .B(n46544), .Z(n46542) );
  OR U55937 ( .A(n46545), .B(n46546), .Z(n46543) );
  NANDN U55938 ( .A(n46547), .B(n46545), .Z(n46541) );
  IV U55939 ( .A(n46546), .Z(n46547) );
  NAND U55940 ( .A(n46548), .B(n46549), .Z(n46523) );
  NAND U55941 ( .A(n46550), .B(n46551), .Z(n46549) );
  NANDN U55942 ( .A(n46552), .B(n46553), .Z(n46550) );
  NANDN U55943 ( .A(n46553), .B(n46552), .Z(n46548) );
  AND U55944 ( .A(n46554), .B(n46555), .Z(n46525) );
  NAND U55945 ( .A(n46556), .B(n46557), .Z(n46555) );
  OR U55946 ( .A(n46558), .B(n46559), .Z(n46556) );
  NANDN U55947 ( .A(n46560), .B(n46558), .Z(n46554) );
  NAND U55948 ( .A(n46561), .B(n46562), .Z(n46529) );
  NANDN U55949 ( .A(n46563), .B(n46564), .Z(n46562) );
  OR U55950 ( .A(n46565), .B(n46566), .Z(n46564) );
  NANDN U55951 ( .A(n46567), .B(n46565), .Z(n46561) );
  IV U55952 ( .A(n46566), .Z(n46567) );
  XNOR U55953 ( .A(n46537), .B(n46568), .Z(n46532) );
  XNOR U55954 ( .A(n46535), .B(n46538), .Z(n46568) );
  NAND U55955 ( .A(n46569), .B(n46570), .Z(n46538) );
  NAND U55956 ( .A(n46571), .B(n46572), .Z(n46570) );
  OR U55957 ( .A(n46573), .B(n46574), .Z(n46571) );
  NANDN U55958 ( .A(n46575), .B(n46573), .Z(n46569) );
  IV U55959 ( .A(n46574), .Z(n46575) );
  NAND U55960 ( .A(n46576), .B(n46577), .Z(n46535) );
  NAND U55961 ( .A(n46578), .B(n46579), .Z(n46577) );
  NANDN U55962 ( .A(n46580), .B(n46581), .Z(n46578) );
  NANDN U55963 ( .A(n46581), .B(n46580), .Z(n46576) );
  AND U55964 ( .A(n46582), .B(n46583), .Z(n46537) );
  NAND U55965 ( .A(n46584), .B(n46585), .Z(n46583) );
  OR U55966 ( .A(n46586), .B(n46587), .Z(n46584) );
  NANDN U55967 ( .A(n46588), .B(n46586), .Z(n46582) );
  XNOR U55968 ( .A(n46563), .B(n46589), .Z(N61269) );
  XOR U55969 ( .A(n46565), .B(n46566), .Z(n46589) );
  XNOR U55970 ( .A(n46579), .B(n46590), .Z(n46566) );
  XOR U55971 ( .A(n46580), .B(n46581), .Z(n46590) );
  XOR U55972 ( .A(n46586), .B(n46591), .Z(n46581) );
  XOR U55973 ( .A(n46585), .B(n46588), .Z(n46591) );
  IV U55974 ( .A(n46587), .Z(n46588) );
  NAND U55975 ( .A(n46592), .B(n46593), .Z(n46587) );
  OR U55976 ( .A(n46594), .B(n46595), .Z(n46593) );
  OR U55977 ( .A(n46596), .B(n46597), .Z(n46592) );
  NAND U55978 ( .A(n46598), .B(n46599), .Z(n46585) );
  OR U55979 ( .A(n46600), .B(n46601), .Z(n46599) );
  OR U55980 ( .A(n46602), .B(n46603), .Z(n46598) );
  NOR U55981 ( .A(n46604), .B(n46605), .Z(n46586) );
  ANDN U55982 ( .B(n46606), .A(n46607), .Z(n46580) );
  XNOR U55983 ( .A(n46573), .B(n46608), .Z(n46579) );
  XNOR U55984 ( .A(n46572), .B(n46574), .Z(n46608) );
  NAND U55985 ( .A(n46609), .B(n46610), .Z(n46574) );
  OR U55986 ( .A(n46611), .B(n46612), .Z(n46610) );
  OR U55987 ( .A(n46613), .B(n46614), .Z(n46609) );
  NAND U55988 ( .A(n46615), .B(n46616), .Z(n46572) );
  OR U55989 ( .A(n46617), .B(n46618), .Z(n46616) );
  OR U55990 ( .A(n46619), .B(n46620), .Z(n46615) );
  ANDN U55991 ( .B(n46621), .A(n46622), .Z(n46573) );
  IV U55992 ( .A(n46623), .Z(n46621) );
  ANDN U55993 ( .B(n46624), .A(n46625), .Z(n46565) );
  XOR U55994 ( .A(n46551), .B(n46626), .Z(n46563) );
  XOR U55995 ( .A(n46552), .B(n46553), .Z(n46626) );
  XOR U55996 ( .A(n46558), .B(n46627), .Z(n46553) );
  XOR U55997 ( .A(n46557), .B(n46560), .Z(n46627) );
  IV U55998 ( .A(n46559), .Z(n46560) );
  NAND U55999 ( .A(n46628), .B(n46629), .Z(n46559) );
  OR U56000 ( .A(n46630), .B(n46631), .Z(n46629) );
  OR U56001 ( .A(n46632), .B(n46633), .Z(n46628) );
  NAND U56002 ( .A(n46634), .B(n46635), .Z(n46557) );
  OR U56003 ( .A(n46636), .B(n46637), .Z(n46635) );
  OR U56004 ( .A(n46638), .B(n46639), .Z(n46634) );
  NOR U56005 ( .A(n46640), .B(n46641), .Z(n46558) );
  ANDN U56006 ( .B(n46642), .A(n46643), .Z(n46552) );
  IV U56007 ( .A(n46644), .Z(n46642) );
  XNOR U56008 ( .A(n46545), .B(n46645), .Z(n46551) );
  XNOR U56009 ( .A(n46544), .B(n46546), .Z(n46645) );
  NAND U56010 ( .A(n46646), .B(n46647), .Z(n46546) );
  OR U56011 ( .A(n46648), .B(n46649), .Z(n46647) );
  OR U56012 ( .A(n46650), .B(n46651), .Z(n46646) );
  NAND U56013 ( .A(n46652), .B(n46653), .Z(n46544) );
  OR U56014 ( .A(n46654), .B(n46655), .Z(n46653) );
  OR U56015 ( .A(n46656), .B(n46657), .Z(n46652) );
  ANDN U56016 ( .B(n46658), .A(n46659), .Z(n46545) );
  IV U56017 ( .A(n46660), .Z(n46658) );
  XNOR U56018 ( .A(n46625), .B(n46624), .Z(N61268) );
  XOR U56019 ( .A(n46644), .B(n46643), .Z(n46624) );
  XNOR U56020 ( .A(n46659), .B(n46660), .Z(n46643) );
  XNOR U56021 ( .A(n46654), .B(n46655), .Z(n46660) );
  XNOR U56022 ( .A(n46656), .B(n46657), .Z(n46655) );
  XNOR U56023 ( .A(y[1261]), .B(x[1261]), .Z(n46657) );
  XNOR U56024 ( .A(y[1262]), .B(x[1262]), .Z(n46656) );
  XNOR U56025 ( .A(y[1260]), .B(x[1260]), .Z(n46654) );
  XNOR U56026 ( .A(n46648), .B(n46649), .Z(n46659) );
  XNOR U56027 ( .A(y[1257]), .B(x[1257]), .Z(n46649) );
  XNOR U56028 ( .A(n46650), .B(n46651), .Z(n46648) );
  XNOR U56029 ( .A(y[1258]), .B(x[1258]), .Z(n46651) );
  XNOR U56030 ( .A(y[1259]), .B(x[1259]), .Z(n46650) );
  XNOR U56031 ( .A(n46641), .B(n46640), .Z(n46644) );
  XNOR U56032 ( .A(n46636), .B(n46637), .Z(n46640) );
  XNOR U56033 ( .A(y[1254]), .B(x[1254]), .Z(n46637) );
  XNOR U56034 ( .A(n46638), .B(n46639), .Z(n46636) );
  XNOR U56035 ( .A(y[1255]), .B(x[1255]), .Z(n46639) );
  XNOR U56036 ( .A(y[1256]), .B(x[1256]), .Z(n46638) );
  XNOR U56037 ( .A(n46630), .B(n46631), .Z(n46641) );
  XNOR U56038 ( .A(y[1251]), .B(x[1251]), .Z(n46631) );
  XNOR U56039 ( .A(n46632), .B(n46633), .Z(n46630) );
  XNOR U56040 ( .A(y[1252]), .B(x[1252]), .Z(n46633) );
  XNOR U56041 ( .A(y[1253]), .B(x[1253]), .Z(n46632) );
  XOR U56042 ( .A(n46606), .B(n46607), .Z(n46625) );
  XNOR U56043 ( .A(n46622), .B(n46623), .Z(n46607) );
  XNOR U56044 ( .A(n46617), .B(n46618), .Z(n46623) );
  XNOR U56045 ( .A(n46619), .B(n46620), .Z(n46618) );
  XNOR U56046 ( .A(y[1249]), .B(x[1249]), .Z(n46620) );
  XNOR U56047 ( .A(y[1250]), .B(x[1250]), .Z(n46619) );
  XNOR U56048 ( .A(y[1248]), .B(x[1248]), .Z(n46617) );
  XNOR U56049 ( .A(n46611), .B(n46612), .Z(n46622) );
  XNOR U56050 ( .A(y[1245]), .B(x[1245]), .Z(n46612) );
  XNOR U56051 ( .A(n46613), .B(n46614), .Z(n46611) );
  XNOR U56052 ( .A(y[1246]), .B(x[1246]), .Z(n46614) );
  XNOR U56053 ( .A(y[1247]), .B(x[1247]), .Z(n46613) );
  XOR U56054 ( .A(n46605), .B(n46604), .Z(n46606) );
  XNOR U56055 ( .A(n46600), .B(n46601), .Z(n46604) );
  XNOR U56056 ( .A(y[1242]), .B(x[1242]), .Z(n46601) );
  XNOR U56057 ( .A(n46602), .B(n46603), .Z(n46600) );
  XNOR U56058 ( .A(y[1243]), .B(x[1243]), .Z(n46603) );
  XNOR U56059 ( .A(y[1244]), .B(x[1244]), .Z(n46602) );
  XNOR U56060 ( .A(n46594), .B(n46595), .Z(n46605) );
  XNOR U56061 ( .A(y[1239]), .B(x[1239]), .Z(n46595) );
  XNOR U56062 ( .A(n46596), .B(n46597), .Z(n46594) );
  XNOR U56063 ( .A(y[1240]), .B(x[1240]), .Z(n46597) );
  XNOR U56064 ( .A(y[1241]), .B(x[1241]), .Z(n46596) );
  NAND U56065 ( .A(n46661), .B(n46662), .Z(N61259) );
  NANDN U56066 ( .A(n46663), .B(n46664), .Z(n46662) );
  OR U56067 ( .A(n46665), .B(n46666), .Z(n46664) );
  NAND U56068 ( .A(n46665), .B(n46666), .Z(n46661) );
  XOR U56069 ( .A(n46665), .B(n46667), .Z(N61258) );
  XNOR U56070 ( .A(n46663), .B(n46666), .Z(n46667) );
  AND U56071 ( .A(n46668), .B(n46669), .Z(n46666) );
  NANDN U56072 ( .A(n46670), .B(n46671), .Z(n46669) );
  NANDN U56073 ( .A(n46672), .B(n46673), .Z(n46671) );
  NANDN U56074 ( .A(n46673), .B(n46672), .Z(n46668) );
  NAND U56075 ( .A(n46674), .B(n46675), .Z(n46663) );
  NANDN U56076 ( .A(n46676), .B(n46677), .Z(n46675) );
  OR U56077 ( .A(n46678), .B(n46679), .Z(n46677) );
  NAND U56078 ( .A(n46679), .B(n46678), .Z(n46674) );
  AND U56079 ( .A(n46680), .B(n46681), .Z(n46665) );
  NANDN U56080 ( .A(n46682), .B(n46683), .Z(n46681) );
  NANDN U56081 ( .A(n46684), .B(n46685), .Z(n46683) );
  NANDN U56082 ( .A(n46685), .B(n46684), .Z(n46680) );
  XOR U56083 ( .A(n46679), .B(n46686), .Z(N61257) );
  XOR U56084 ( .A(n46676), .B(n46678), .Z(n46686) );
  XNOR U56085 ( .A(n46672), .B(n46687), .Z(n46678) );
  XNOR U56086 ( .A(n46670), .B(n46673), .Z(n46687) );
  NAND U56087 ( .A(n46688), .B(n46689), .Z(n46673) );
  NAND U56088 ( .A(n46690), .B(n46691), .Z(n46689) );
  OR U56089 ( .A(n46692), .B(n46693), .Z(n46690) );
  NANDN U56090 ( .A(n46694), .B(n46692), .Z(n46688) );
  IV U56091 ( .A(n46693), .Z(n46694) );
  NAND U56092 ( .A(n46695), .B(n46696), .Z(n46670) );
  NAND U56093 ( .A(n46697), .B(n46698), .Z(n46696) );
  NANDN U56094 ( .A(n46699), .B(n46700), .Z(n46697) );
  NANDN U56095 ( .A(n46700), .B(n46699), .Z(n46695) );
  AND U56096 ( .A(n46701), .B(n46702), .Z(n46672) );
  NAND U56097 ( .A(n46703), .B(n46704), .Z(n46702) );
  OR U56098 ( .A(n46705), .B(n46706), .Z(n46703) );
  NANDN U56099 ( .A(n46707), .B(n46705), .Z(n46701) );
  NAND U56100 ( .A(n46708), .B(n46709), .Z(n46676) );
  NANDN U56101 ( .A(n46710), .B(n46711), .Z(n46709) );
  OR U56102 ( .A(n46712), .B(n46713), .Z(n46711) );
  NANDN U56103 ( .A(n46714), .B(n46712), .Z(n46708) );
  IV U56104 ( .A(n46713), .Z(n46714) );
  XNOR U56105 ( .A(n46684), .B(n46715), .Z(n46679) );
  XNOR U56106 ( .A(n46682), .B(n46685), .Z(n46715) );
  NAND U56107 ( .A(n46716), .B(n46717), .Z(n46685) );
  NAND U56108 ( .A(n46718), .B(n46719), .Z(n46717) );
  OR U56109 ( .A(n46720), .B(n46721), .Z(n46718) );
  NANDN U56110 ( .A(n46722), .B(n46720), .Z(n46716) );
  IV U56111 ( .A(n46721), .Z(n46722) );
  NAND U56112 ( .A(n46723), .B(n46724), .Z(n46682) );
  NAND U56113 ( .A(n46725), .B(n46726), .Z(n46724) );
  NANDN U56114 ( .A(n46727), .B(n46728), .Z(n46725) );
  NANDN U56115 ( .A(n46728), .B(n46727), .Z(n46723) );
  AND U56116 ( .A(n46729), .B(n46730), .Z(n46684) );
  NAND U56117 ( .A(n46731), .B(n46732), .Z(n46730) );
  OR U56118 ( .A(n46733), .B(n46734), .Z(n46731) );
  NANDN U56119 ( .A(n46735), .B(n46733), .Z(n46729) );
  XNOR U56120 ( .A(n46710), .B(n46736), .Z(N61256) );
  XOR U56121 ( .A(n46712), .B(n46713), .Z(n46736) );
  XNOR U56122 ( .A(n46726), .B(n46737), .Z(n46713) );
  XOR U56123 ( .A(n46727), .B(n46728), .Z(n46737) );
  XOR U56124 ( .A(n46733), .B(n46738), .Z(n46728) );
  XOR U56125 ( .A(n46732), .B(n46735), .Z(n46738) );
  IV U56126 ( .A(n46734), .Z(n46735) );
  NAND U56127 ( .A(n46739), .B(n46740), .Z(n46734) );
  OR U56128 ( .A(n46741), .B(n46742), .Z(n46740) );
  OR U56129 ( .A(n46743), .B(n46744), .Z(n46739) );
  NAND U56130 ( .A(n46745), .B(n46746), .Z(n46732) );
  OR U56131 ( .A(n46747), .B(n46748), .Z(n46746) );
  OR U56132 ( .A(n46749), .B(n46750), .Z(n46745) );
  NOR U56133 ( .A(n46751), .B(n46752), .Z(n46733) );
  ANDN U56134 ( .B(n46753), .A(n46754), .Z(n46727) );
  XNOR U56135 ( .A(n46720), .B(n46755), .Z(n46726) );
  XNOR U56136 ( .A(n46719), .B(n46721), .Z(n46755) );
  NAND U56137 ( .A(n46756), .B(n46757), .Z(n46721) );
  OR U56138 ( .A(n46758), .B(n46759), .Z(n46757) );
  OR U56139 ( .A(n46760), .B(n46761), .Z(n46756) );
  NAND U56140 ( .A(n46762), .B(n46763), .Z(n46719) );
  OR U56141 ( .A(n46764), .B(n46765), .Z(n46763) );
  OR U56142 ( .A(n46766), .B(n46767), .Z(n46762) );
  ANDN U56143 ( .B(n46768), .A(n46769), .Z(n46720) );
  IV U56144 ( .A(n46770), .Z(n46768) );
  ANDN U56145 ( .B(n46771), .A(n46772), .Z(n46712) );
  XOR U56146 ( .A(n46698), .B(n46773), .Z(n46710) );
  XOR U56147 ( .A(n46699), .B(n46700), .Z(n46773) );
  XOR U56148 ( .A(n46705), .B(n46774), .Z(n46700) );
  XOR U56149 ( .A(n46704), .B(n46707), .Z(n46774) );
  IV U56150 ( .A(n46706), .Z(n46707) );
  NAND U56151 ( .A(n46775), .B(n46776), .Z(n46706) );
  OR U56152 ( .A(n46777), .B(n46778), .Z(n46776) );
  OR U56153 ( .A(n46779), .B(n46780), .Z(n46775) );
  NAND U56154 ( .A(n46781), .B(n46782), .Z(n46704) );
  OR U56155 ( .A(n46783), .B(n46784), .Z(n46782) );
  OR U56156 ( .A(n46785), .B(n46786), .Z(n46781) );
  NOR U56157 ( .A(n46787), .B(n46788), .Z(n46705) );
  ANDN U56158 ( .B(n46789), .A(n46790), .Z(n46699) );
  IV U56159 ( .A(n46791), .Z(n46789) );
  XNOR U56160 ( .A(n46692), .B(n46792), .Z(n46698) );
  XNOR U56161 ( .A(n46691), .B(n46693), .Z(n46792) );
  NAND U56162 ( .A(n46793), .B(n46794), .Z(n46693) );
  OR U56163 ( .A(n46795), .B(n46796), .Z(n46794) );
  OR U56164 ( .A(n46797), .B(n46798), .Z(n46793) );
  NAND U56165 ( .A(n46799), .B(n46800), .Z(n46691) );
  OR U56166 ( .A(n46801), .B(n46802), .Z(n46800) );
  OR U56167 ( .A(n46803), .B(n46804), .Z(n46799) );
  ANDN U56168 ( .B(n46805), .A(n46806), .Z(n46692) );
  IV U56169 ( .A(n46807), .Z(n46805) );
  XNOR U56170 ( .A(n46772), .B(n46771), .Z(N61255) );
  XOR U56171 ( .A(n46791), .B(n46790), .Z(n46771) );
  XNOR U56172 ( .A(n46806), .B(n46807), .Z(n46790) );
  XNOR U56173 ( .A(n46801), .B(n46802), .Z(n46807) );
  XNOR U56174 ( .A(n46803), .B(n46804), .Z(n46802) );
  XNOR U56175 ( .A(y[1237]), .B(x[1237]), .Z(n46804) );
  XNOR U56176 ( .A(y[1238]), .B(x[1238]), .Z(n46803) );
  XNOR U56177 ( .A(y[1236]), .B(x[1236]), .Z(n46801) );
  XNOR U56178 ( .A(n46795), .B(n46796), .Z(n46806) );
  XNOR U56179 ( .A(y[1233]), .B(x[1233]), .Z(n46796) );
  XNOR U56180 ( .A(n46797), .B(n46798), .Z(n46795) );
  XNOR U56181 ( .A(y[1234]), .B(x[1234]), .Z(n46798) );
  XNOR U56182 ( .A(y[1235]), .B(x[1235]), .Z(n46797) );
  XNOR U56183 ( .A(n46788), .B(n46787), .Z(n46791) );
  XNOR U56184 ( .A(n46783), .B(n46784), .Z(n46787) );
  XNOR U56185 ( .A(y[1230]), .B(x[1230]), .Z(n46784) );
  XNOR U56186 ( .A(n46785), .B(n46786), .Z(n46783) );
  XNOR U56187 ( .A(y[1231]), .B(x[1231]), .Z(n46786) );
  XNOR U56188 ( .A(y[1232]), .B(x[1232]), .Z(n46785) );
  XNOR U56189 ( .A(n46777), .B(n46778), .Z(n46788) );
  XNOR U56190 ( .A(y[1227]), .B(x[1227]), .Z(n46778) );
  XNOR U56191 ( .A(n46779), .B(n46780), .Z(n46777) );
  XNOR U56192 ( .A(y[1228]), .B(x[1228]), .Z(n46780) );
  XNOR U56193 ( .A(y[1229]), .B(x[1229]), .Z(n46779) );
  XOR U56194 ( .A(n46753), .B(n46754), .Z(n46772) );
  XNOR U56195 ( .A(n46769), .B(n46770), .Z(n46754) );
  XNOR U56196 ( .A(n46764), .B(n46765), .Z(n46770) );
  XNOR U56197 ( .A(n46766), .B(n46767), .Z(n46765) );
  XNOR U56198 ( .A(y[1225]), .B(x[1225]), .Z(n46767) );
  XNOR U56199 ( .A(y[1226]), .B(x[1226]), .Z(n46766) );
  XNOR U56200 ( .A(y[1224]), .B(x[1224]), .Z(n46764) );
  XNOR U56201 ( .A(n46758), .B(n46759), .Z(n46769) );
  XNOR U56202 ( .A(y[1221]), .B(x[1221]), .Z(n46759) );
  XNOR U56203 ( .A(n46760), .B(n46761), .Z(n46758) );
  XNOR U56204 ( .A(y[1222]), .B(x[1222]), .Z(n46761) );
  XNOR U56205 ( .A(y[1223]), .B(x[1223]), .Z(n46760) );
  XOR U56206 ( .A(n46752), .B(n46751), .Z(n46753) );
  XNOR U56207 ( .A(n46747), .B(n46748), .Z(n46751) );
  XNOR U56208 ( .A(y[1218]), .B(x[1218]), .Z(n46748) );
  XNOR U56209 ( .A(n46749), .B(n46750), .Z(n46747) );
  XNOR U56210 ( .A(y[1219]), .B(x[1219]), .Z(n46750) );
  XNOR U56211 ( .A(y[1220]), .B(x[1220]), .Z(n46749) );
  XNOR U56212 ( .A(n46741), .B(n46742), .Z(n46752) );
  XNOR U56213 ( .A(y[1215]), .B(x[1215]), .Z(n46742) );
  XNOR U56214 ( .A(n46743), .B(n46744), .Z(n46741) );
  XNOR U56215 ( .A(y[1216]), .B(x[1216]), .Z(n46744) );
  XNOR U56216 ( .A(y[1217]), .B(x[1217]), .Z(n46743) );
  NAND U56217 ( .A(n46808), .B(n46809), .Z(N61246) );
  NANDN U56218 ( .A(n46810), .B(n46811), .Z(n46809) );
  OR U56219 ( .A(n46812), .B(n46813), .Z(n46811) );
  NAND U56220 ( .A(n46812), .B(n46813), .Z(n46808) );
  XOR U56221 ( .A(n46812), .B(n46814), .Z(N61245) );
  XNOR U56222 ( .A(n46810), .B(n46813), .Z(n46814) );
  AND U56223 ( .A(n46815), .B(n46816), .Z(n46813) );
  NANDN U56224 ( .A(n46817), .B(n46818), .Z(n46816) );
  NANDN U56225 ( .A(n46819), .B(n46820), .Z(n46818) );
  NANDN U56226 ( .A(n46820), .B(n46819), .Z(n46815) );
  NAND U56227 ( .A(n46821), .B(n46822), .Z(n46810) );
  NANDN U56228 ( .A(n46823), .B(n46824), .Z(n46822) );
  OR U56229 ( .A(n46825), .B(n46826), .Z(n46824) );
  NAND U56230 ( .A(n46826), .B(n46825), .Z(n46821) );
  AND U56231 ( .A(n46827), .B(n46828), .Z(n46812) );
  NANDN U56232 ( .A(n46829), .B(n46830), .Z(n46828) );
  NANDN U56233 ( .A(n46831), .B(n46832), .Z(n46830) );
  NANDN U56234 ( .A(n46832), .B(n46831), .Z(n46827) );
  XOR U56235 ( .A(n46826), .B(n46833), .Z(N61244) );
  XOR U56236 ( .A(n46823), .B(n46825), .Z(n46833) );
  XNOR U56237 ( .A(n46819), .B(n46834), .Z(n46825) );
  XNOR U56238 ( .A(n46817), .B(n46820), .Z(n46834) );
  NAND U56239 ( .A(n46835), .B(n46836), .Z(n46820) );
  NAND U56240 ( .A(n46837), .B(n46838), .Z(n46836) );
  OR U56241 ( .A(n46839), .B(n46840), .Z(n46837) );
  NANDN U56242 ( .A(n46841), .B(n46839), .Z(n46835) );
  IV U56243 ( .A(n46840), .Z(n46841) );
  NAND U56244 ( .A(n46842), .B(n46843), .Z(n46817) );
  NAND U56245 ( .A(n46844), .B(n46845), .Z(n46843) );
  NANDN U56246 ( .A(n46846), .B(n46847), .Z(n46844) );
  NANDN U56247 ( .A(n46847), .B(n46846), .Z(n46842) );
  AND U56248 ( .A(n46848), .B(n46849), .Z(n46819) );
  NAND U56249 ( .A(n46850), .B(n46851), .Z(n46849) );
  OR U56250 ( .A(n46852), .B(n46853), .Z(n46850) );
  NANDN U56251 ( .A(n46854), .B(n46852), .Z(n46848) );
  NAND U56252 ( .A(n46855), .B(n46856), .Z(n46823) );
  NANDN U56253 ( .A(n46857), .B(n46858), .Z(n46856) );
  OR U56254 ( .A(n46859), .B(n46860), .Z(n46858) );
  NANDN U56255 ( .A(n46861), .B(n46859), .Z(n46855) );
  IV U56256 ( .A(n46860), .Z(n46861) );
  XNOR U56257 ( .A(n46831), .B(n46862), .Z(n46826) );
  XNOR U56258 ( .A(n46829), .B(n46832), .Z(n46862) );
  NAND U56259 ( .A(n46863), .B(n46864), .Z(n46832) );
  NAND U56260 ( .A(n46865), .B(n46866), .Z(n46864) );
  OR U56261 ( .A(n46867), .B(n46868), .Z(n46865) );
  NANDN U56262 ( .A(n46869), .B(n46867), .Z(n46863) );
  IV U56263 ( .A(n46868), .Z(n46869) );
  NAND U56264 ( .A(n46870), .B(n46871), .Z(n46829) );
  NAND U56265 ( .A(n46872), .B(n46873), .Z(n46871) );
  NANDN U56266 ( .A(n46874), .B(n46875), .Z(n46872) );
  NANDN U56267 ( .A(n46875), .B(n46874), .Z(n46870) );
  AND U56268 ( .A(n46876), .B(n46877), .Z(n46831) );
  NAND U56269 ( .A(n46878), .B(n46879), .Z(n46877) );
  OR U56270 ( .A(n46880), .B(n46881), .Z(n46878) );
  NANDN U56271 ( .A(n46882), .B(n46880), .Z(n46876) );
  XNOR U56272 ( .A(n46857), .B(n46883), .Z(N61243) );
  XOR U56273 ( .A(n46859), .B(n46860), .Z(n46883) );
  XNOR U56274 ( .A(n46873), .B(n46884), .Z(n46860) );
  XOR U56275 ( .A(n46874), .B(n46875), .Z(n46884) );
  XOR U56276 ( .A(n46880), .B(n46885), .Z(n46875) );
  XOR U56277 ( .A(n46879), .B(n46882), .Z(n46885) );
  IV U56278 ( .A(n46881), .Z(n46882) );
  NAND U56279 ( .A(n46886), .B(n46887), .Z(n46881) );
  OR U56280 ( .A(n46888), .B(n46889), .Z(n46887) );
  OR U56281 ( .A(n46890), .B(n46891), .Z(n46886) );
  NAND U56282 ( .A(n46892), .B(n46893), .Z(n46879) );
  OR U56283 ( .A(n46894), .B(n46895), .Z(n46893) );
  OR U56284 ( .A(n46896), .B(n46897), .Z(n46892) );
  NOR U56285 ( .A(n46898), .B(n46899), .Z(n46880) );
  ANDN U56286 ( .B(n46900), .A(n46901), .Z(n46874) );
  XNOR U56287 ( .A(n46867), .B(n46902), .Z(n46873) );
  XNOR U56288 ( .A(n46866), .B(n46868), .Z(n46902) );
  NAND U56289 ( .A(n46903), .B(n46904), .Z(n46868) );
  OR U56290 ( .A(n46905), .B(n46906), .Z(n46904) );
  OR U56291 ( .A(n46907), .B(n46908), .Z(n46903) );
  NAND U56292 ( .A(n46909), .B(n46910), .Z(n46866) );
  OR U56293 ( .A(n46911), .B(n46912), .Z(n46910) );
  OR U56294 ( .A(n46913), .B(n46914), .Z(n46909) );
  ANDN U56295 ( .B(n46915), .A(n46916), .Z(n46867) );
  IV U56296 ( .A(n46917), .Z(n46915) );
  ANDN U56297 ( .B(n46918), .A(n46919), .Z(n46859) );
  XOR U56298 ( .A(n46845), .B(n46920), .Z(n46857) );
  XOR U56299 ( .A(n46846), .B(n46847), .Z(n46920) );
  XOR U56300 ( .A(n46852), .B(n46921), .Z(n46847) );
  XOR U56301 ( .A(n46851), .B(n46854), .Z(n46921) );
  IV U56302 ( .A(n46853), .Z(n46854) );
  NAND U56303 ( .A(n46922), .B(n46923), .Z(n46853) );
  OR U56304 ( .A(n46924), .B(n46925), .Z(n46923) );
  OR U56305 ( .A(n46926), .B(n46927), .Z(n46922) );
  NAND U56306 ( .A(n46928), .B(n46929), .Z(n46851) );
  OR U56307 ( .A(n46930), .B(n46931), .Z(n46929) );
  OR U56308 ( .A(n46932), .B(n46933), .Z(n46928) );
  NOR U56309 ( .A(n46934), .B(n46935), .Z(n46852) );
  ANDN U56310 ( .B(n46936), .A(n46937), .Z(n46846) );
  IV U56311 ( .A(n46938), .Z(n46936) );
  XNOR U56312 ( .A(n46839), .B(n46939), .Z(n46845) );
  XNOR U56313 ( .A(n46838), .B(n46840), .Z(n46939) );
  NAND U56314 ( .A(n46940), .B(n46941), .Z(n46840) );
  OR U56315 ( .A(n46942), .B(n46943), .Z(n46941) );
  OR U56316 ( .A(n46944), .B(n46945), .Z(n46940) );
  NAND U56317 ( .A(n46946), .B(n46947), .Z(n46838) );
  OR U56318 ( .A(n46948), .B(n46949), .Z(n46947) );
  OR U56319 ( .A(n46950), .B(n46951), .Z(n46946) );
  ANDN U56320 ( .B(n46952), .A(n46953), .Z(n46839) );
  IV U56321 ( .A(n46954), .Z(n46952) );
  XNOR U56322 ( .A(n46919), .B(n46918), .Z(N61242) );
  XOR U56323 ( .A(n46938), .B(n46937), .Z(n46918) );
  XNOR U56324 ( .A(n46953), .B(n46954), .Z(n46937) );
  XNOR U56325 ( .A(n46948), .B(n46949), .Z(n46954) );
  XNOR U56326 ( .A(n46950), .B(n46951), .Z(n46949) );
  XNOR U56327 ( .A(y[1213]), .B(x[1213]), .Z(n46951) );
  XNOR U56328 ( .A(y[1214]), .B(x[1214]), .Z(n46950) );
  XNOR U56329 ( .A(y[1212]), .B(x[1212]), .Z(n46948) );
  XNOR U56330 ( .A(n46942), .B(n46943), .Z(n46953) );
  XNOR U56331 ( .A(y[1209]), .B(x[1209]), .Z(n46943) );
  XNOR U56332 ( .A(n46944), .B(n46945), .Z(n46942) );
  XNOR U56333 ( .A(y[1210]), .B(x[1210]), .Z(n46945) );
  XNOR U56334 ( .A(y[1211]), .B(x[1211]), .Z(n46944) );
  XNOR U56335 ( .A(n46935), .B(n46934), .Z(n46938) );
  XNOR U56336 ( .A(n46930), .B(n46931), .Z(n46934) );
  XNOR U56337 ( .A(y[1206]), .B(x[1206]), .Z(n46931) );
  XNOR U56338 ( .A(n46932), .B(n46933), .Z(n46930) );
  XNOR U56339 ( .A(y[1207]), .B(x[1207]), .Z(n46933) );
  XNOR U56340 ( .A(y[1208]), .B(x[1208]), .Z(n46932) );
  XNOR U56341 ( .A(n46924), .B(n46925), .Z(n46935) );
  XNOR U56342 ( .A(y[1203]), .B(x[1203]), .Z(n46925) );
  XNOR U56343 ( .A(n46926), .B(n46927), .Z(n46924) );
  XNOR U56344 ( .A(y[1204]), .B(x[1204]), .Z(n46927) );
  XNOR U56345 ( .A(y[1205]), .B(x[1205]), .Z(n46926) );
  XOR U56346 ( .A(n46900), .B(n46901), .Z(n46919) );
  XNOR U56347 ( .A(n46916), .B(n46917), .Z(n46901) );
  XNOR U56348 ( .A(n46911), .B(n46912), .Z(n46917) );
  XNOR U56349 ( .A(n46913), .B(n46914), .Z(n46912) );
  XNOR U56350 ( .A(y[1201]), .B(x[1201]), .Z(n46914) );
  XNOR U56351 ( .A(y[1202]), .B(x[1202]), .Z(n46913) );
  XNOR U56352 ( .A(y[1200]), .B(x[1200]), .Z(n46911) );
  XNOR U56353 ( .A(n46905), .B(n46906), .Z(n46916) );
  XNOR U56354 ( .A(y[1197]), .B(x[1197]), .Z(n46906) );
  XNOR U56355 ( .A(n46907), .B(n46908), .Z(n46905) );
  XNOR U56356 ( .A(y[1198]), .B(x[1198]), .Z(n46908) );
  XNOR U56357 ( .A(y[1199]), .B(x[1199]), .Z(n46907) );
  XOR U56358 ( .A(n46899), .B(n46898), .Z(n46900) );
  XNOR U56359 ( .A(n46894), .B(n46895), .Z(n46898) );
  XNOR U56360 ( .A(y[1194]), .B(x[1194]), .Z(n46895) );
  XNOR U56361 ( .A(n46896), .B(n46897), .Z(n46894) );
  XNOR U56362 ( .A(y[1195]), .B(x[1195]), .Z(n46897) );
  XNOR U56363 ( .A(y[1196]), .B(x[1196]), .Z(n46896) );
  XNOR U56364 ( .A(n46888), .B(n46889), .Z(n46899) );
  XNOR U56365 ( .A(y[1191]), .B(x[1191]), .Z(n46889) );
  XNOR U56366 ( .A(n46890), .B(n46891), .Z(n46888) );
  XNOR U56367 ( .A(y[1192]), .B(x[1192]), .Z(n46891) );
  XNOR U56368 ( .A(y[1193]), .B(x[1193]), .Z(n46890) );
  NAND U56369 ( .A(n46955), .B(n46956), .Z(N61233) );
  NANDN U56370 ( .A(n46957), .B(n46958), .Z(n46956) );
  OR U56371 ( .A(n46959), .B(n46960), .Z(n46958) );
  NAND U56372 ( .A(n46959), .B(n46960), .Z(n46955) );
  XOR U56373 ( .A(n46959), .B(n46961), .Z(N61232) );
  XNOR U56374 ( .A(n46957), .B(n46960), .Z(n46961) );
  AND U56375 ( .A(n46962), .B(n46963), .Z(n46960) );
  NANDN U56376 ( .A(n46964), .B(n46965), .Z(n46963) );
  NANDN U56377 ( .A(n46966), .B(n46967), .Z(n46965) );
  NANDN U56378 ( .A(n46967), .B(n46966), .Z(n46962) );
  NAND U56379 ( .A(n46968), .B(n46969), .Z(n46957) );
  NANDN U56380 ( .A(n46970), .B(n46971), .Z(n46969) );
  OR U56381 ( .A(n46972), .B(n46973), .Z(n46971) );
  NAND U56382 ( .A(n46973), .B(n46972), .Z(n46968) );
  AND U56383 ( .A(n46974), .B(n46975), .Z(n46959) );
  NANDN U56384 ( .A(n46976), .B(n46977), .Z(n46975) );
  NANDN U56385 ( .A(n46978), .B(n46979), .Z(n46977) );
  NANDN U56386 ( .A(n46979), .B(n46978), .Z(n46974) );
  XOR U56387 ( .A(n46973), .B(n46980), .Z(N61231) );
  XOR U56388 ( .A(n46970), .B(n46972), .Z(n46980) );
  XNOR U56389 ( .A(n46966), .B(n46981), .Z(n46972) );
  XNOR U56390 ( .A(n46964), .B(n46967), .Z(n46981) );
  NAND U56391 ( .A(n46982), .B(n46983), .Z(n46967) );
  NAND U56392 ( .A(n46984), .B(n46985), .Z(n46983) );
  OR U56393 ( .A(n46986), .B(n46987), .Z(n46984) );
  NANDN U56394 ( .A(n46988), .B(n46986), .Z(n46982) );
  IV U56395 ( .A(n46987), .Z(n46988) );
  NAND U56396 ( .A(n46989), .B(n46990), .Z(n46964) );
  NAND U56397 ( .A(n46991), .B(n46992), .Z(n46990) );
  NANDN U56398 ( .A(n46993), .B(n46994), .Z(n46991) );
  NANDN U56399 ( .A(n46994), .B(n46993), .Z(n46989) );
  AND U56400 ( .A(n46995), .B(n46996), .Z(n46966) );
  NAND U56401 ( .A(n46997), .B(n46998), .Z(n46996) );
  OR U56402 ( .A(n46999), .B(n47000), .Z(n46997) );
  NANDN U56403 ( .A(n47001), .B(n46999), .Z(n46995) );
  NAND U56404 ( .A(n47002), .B(n47003), .Z(n46970) );
  NANDN U56405 ( .A(n47004), .B(n47005), .Z(n47003) );
  OR U56406 ( .A(n47006), .B(n47007), .Z(n47005) );
  NANDN U56407 ( .A(n47008), .B(n47006), .Z(n47002) );
  IV U56408 ( .A(n47007), .Z(n47008) );
  XNOR U56409 ( .A(n46978), .B(n47009), .Z(n46973) );
  XNOR U56410 ( .A(n46976), .B(n46979), .Z(n47009) );
  NAND U56411 ( .A(n47010), .B(n47011), .Z(n46979) );
  NAND U56412 ( .A(n47012), .B(n47013), .Z(n47011) );
  OR U56413 ( .A(n47014), .B(n47015), .Z(n47012) );
  NANDN U56414 ( .A(n47016), .B(n47014), .Z(n47010) );
  IV U56415 ( .A(n47015), .Z(n47016) );
  NAND U56416 ( .A(n47017), .B(n47018), .Z(n46976) );
  NAND U56417 ( .A(n47019), .B(n47020), .Z(n47018) );
  NANDN U56418 ( .A(n47021), .B(n47022), .Z(n47019) );
  NANDN U56419 ( .A(n47022), .B(n47021), .Z(n47017) );
  AND U56420 ( .A(n47023), .B(n47024), .Z(n46978) );
  NAND U56421 ( .A(n47025), .B(n47026), .Z(n47024) );
  OR U56422 ( .A(n47027), .B(n47028), .Z(n47025) );
  NANDN U56423 ( .A(n47029), .B(n47027), .Z(n47023) );
  XNOR U56424 ( .A(n47004), .B(n47030), .Z(N61230) );
  XOR U56425 ( .A(n47006), .B(n47007), .Z(n47030) );
  XNOR U56426 ( .A(n47020), .B(n47031), .Z(n47007) );
  XOR U56427 ( .A(n47021), .B(n47022), .Z(n47031) );
  XOR U56428 ( .A(n47027), .B(n47032), .Z(n47022) );
  XOR U56429 ( .A(n47026), .B(n47029), .Z(n47032) );
  IV U56430 ( .A(n47028), .Z(n47029) );
  NAND U56431 ( .A(n47033), .B(n47034), .Z(n47028) );
  OR U56432 ( .A(n47035), .B(n47036), .Z(n47034) );
  OR U56433 ( .A(n47037), .B(n47038), .Z(n47033) );
  NAND U56434 ( .A(n47039), .B(n47040), .Z(n47026) );
  OR U56435 ( .A(n47041), .B(n47042), .Z(n47040) );
  OR U56436 ( .A(n47043), .B(n47044), .Z(n47039) );
  NOR U56437 ( .A(n47045), .B(n47046), .Z(n47027) );
  ANDN U56438 ( .B(n47047), .A(n47048), .Z(n47021) );
  XNOR U56439 ( .A(n47014), .B(n47049), .Z(n47020) );
  XNOR U56440 ( .A(n47013), .B(n47015), .Z(n47049) );
  NAND U56441 ( .A(n47050), .B(n47051), .Z(n47015) );
  OR U56442 ( .A(n47052), .B(n47053), .Z(n47051) );
  OR U56443 ( .A(n47054), .B(n47055), .Z(n47050) );
  NAND U56444 ( .A(n47056), .B(n47057), .Z(n47013) );
  OR U56445 ( .A(n47058), .B(n47059), .Z(n47057) );
  OR U56446 ( .A(n47060), .B(n47061), .Z(n47056) );
  ANDN U56447 ( .B(n47062), .A(n47063), .Z(n47014) );
  IV U56448 ( .A(n47064), .Z(n47062) );
  ANDN U56449 ( .B(n47065), .A(n47066), .Z(n47006) );
  XOR U56450 ( .A(n46992), .B(n47067), .Z(n47004) );
  XOR U56451 ( .A(n46993), .B(n46994), .Z(n47067) );
  XOR U56452 ( .A(n46999), .B(n47068), .Z(n46994) );
  XOR U56453 ( .A(n46998), .B(n47001), .Z(n47068) );
  IV U56454 ( .A(n47000), .Z(n47001) );
  NAND U56455 ( .A(n47069), .B(n47070), .Z(n47000) );
  OR U56456 ( .A(n47071), .B(n47072), .Z(n47070) );
  OR U56457 ( .A(n47073), .B(n47074), .Z(n47069) );
  NAND U56458 ( .A(n47075), .B(n47076), .Z(n46998) );
  OR U56459 ( .A(n47077), .B(n47078), .Z(n47076) );
  OR U56460 ( .A(n47079), .B(n47080), .Z(n47075) );
  NOR U56461 ( .A(n47081), .B(n47082), .Z(n46999) );
  ANDN U56462 ( .B(n47083), .A(n47084), .Z(n46993) );
  IV U56463 ( .A(n47085), .Z(n47083) );
  XNOR U56464 ( .A(n46986), .B(n47086), .Z(n46992) );
  XNOR U56465 ( .A(n46985), .B(n46987), .Z(n47086) );
  NAND U56466 ( .A(n47087), .B(n47088), .Z(n46987) );
  OR U56467 ( .A(n47089), .B(n47090), .Z(n47088) );
  OR U56468 ( .A(n47091), .B(n47092), .Z(n47087) );
  NAND U56469 ( .A(n47093), .B(n47094), .Z(n46985) );
  OR U56470 ( .A(n47095), .B(n47096), .Z(n47094) );
  OR U56471 ( .A(n47097), .B(n47098), .Z(n47093) );
  ANDN U56472 ( .B(n47099), .A(n47100), .Z(n46986) );
  IV U56473 ( .A(n47101), .Z(n47099) );
  XNOR U56474 ( .A(n47066), .B(n47065), .Z(N61229) );
  XOR U56475 ( .A(n47085), .B(n47084), .Z(n47065) );
  XNOR U56476 ( .A(n47100), .B(n47101), .Z(n47084) );
  XNOR U56477 ( .A(n47095), .B(n47096), .Z(n47101) );
  XNOR U56478 ( .A(n47097), .B(n47098), .Z(n47096) );
  XNOR U56479 ( .A(y[1189]), .B(x[1189]), .Z(n47098) );
  XNOR U56480 ( .A(y[1190]), .B(x[1190]), .Z(n47097) );
  XNOR U56481 ( .A(y[1188]), .B(x[1188]), .Z(n47095) );
  XNOR U56482 ( .A(n47089), .B(n47090), .Z(n47100) );
  XNOR U56483 ( .A(y[1185]), .B(x[1185]), .Z(n47090) );
  XNOR U56484 ( .A(n47091), .B(n47092), .Z(n47089) );
  XNOR U56485 ( .A(y[1186]), .B(x[1186]), .Z(n47092) );
  XNOR U56486 ( .A(y[1187]), .B(x[1187]), .Z(n47091) );
  XNOR U56487 ( .A(n47082), .B(n47081), .Z(n47085) );
  XNOR U56488 ( .A(n47077), .B(n47078), .Z(n47081) );
  XNOR U56489 ( .A(y[1182]), .B(x[1182]), .Z(n47078) );
  XNOR U56490 ( .A(n47079), .B(n47080), .Z(n47077) );
  XNOR U56491 ( .A(y[1183]), .B(x[1183]), .Z(n47080) );
  XNOR U56492 ( .A(y[1184]), .B(x[1184]), .Z(n47079) );
  XNOR U56493 ( .A(n47071), .B(n47072), .Z(n47082) );
  XNOR U56494 ( .A(y[1179]), .B(x[1179]), .Z(n47072) );
  XNOR U56495 ( .A(n47073), .B(n47074), .Z(n47071) );
  XNOR U56496 ( .A(y[1180]), .B(x[1180]), .Z(n47074) );
  XNOR U56497 ( .A(y[1181]), .B(x[1181]), .Z(n47073) );
  XOR U56498 ( .A(n47047), .B(n47048), .Z(n47066) );
  XNOR U56499 ( .A(n47063), .B(n47064), .Z(n47048) );
  XNOR U56500 ( .A(n47058), .B(n47059), .Z(n47064) );
  XNOR U56501 ( .A(n47060), .B(n47061), .Z(n47059) );
  XNOR U56502 ( .A(y[1177]), .B(x[1177]), .Z(n47061) );
  XNOR U56503 ( .A(y[1178]), .B(x[1178]), .Z(n47060) );
  XNOR U56504 ( .A(y[1176]), .B(x[1176]), .Z(n47058) );
  XNOR U56505 ( .A(n47052), .B(n47053), .Z(n47063) );
  XNOR U56506 ( .A(y[1173]), .B(x[1173]), .Z(n47053) );
  XNOR U56507 ( .A(n47054), .B(n47055), .Z(n47052) );
  XNOR U56508 ( .A(y[1174]), .B(x[1174]), .Z(n47055) );
  XNOR U56509 ( .A(y[1175]), .B(x[1175]), .Z(n47054) );
  XOR U56510 ( .A(n47046), .B(n47045), .Z(n47047) );
  XNOR U56511 ( .A(n47041), .B(n47042), .Z(n47045) );
  XNOR U56512 ( .A(y[1170]), .B(x[1170]), .Z(n47042) );
  XNOR U56513 ( .A(n47043), .B(n47044), .Z(n47041) );
  XNOR U56514 ( .A(y[1171]), .B(x[1171]), .Z(n47044) );
  XNOR U56515 ( .A(y[1172]), .B(x[1172]), .Z(n47043) );
  XNOR U56516 ( .A(n47035), .B(n47036), .Z(n47046) );
  XNOR U56517 ( .A(y[1167]), .B(x[1167]), .Z(n47036) );
  XNOR U56518 ( .A(n47037), .B(n47038), .Z(n47035) );
  XNOR U56519 ( .A(y[1168]), .B(x[1168]), .Z(n47038) );
  XNOR U56520 ( .A(y[1169]), .B(x[1169]), .Z(n47037) );
  NAND U56521 ( .A(n47102), .B(n47103), .Z(N61220) );
  NANDN U56522 ( .A(n47104), .B(n47105), .Z(n47103) );
  OR U56523 ( .A(n47106), .B(n47107), .Z(n47105) );
  NAND U56524 ( .A(n47106), .B(n47107), .Z(n47102) );
  XOR U56525 ( .A(n47106), .B(n47108), .Z(N61219) );
  XNOR U56526 ( .A(n47104), .B(n47107), .Z(n47108) );
  AND U56527 ( .A(n47109), .B(n47110), .Z(n47107) );
  NANDN U56528 ( .A(n47111), .B(n47112), .Z(n47110) );
  NANDN U56529 ( .A(n47113), .B(n47114), .Z(n47112) );
  NANDN U56530 ( .A(n47114), .B(n47113), .Z(n47109) );
  NAND U56531 ( .A(n47115), .B(n47116), .Z(n47104) );
  NANDN U56532 ( .A(n47117), .B(n47118), .Z(n47116) );
  OR U56533 ( .A(n47119), .B(n47120), .Z(n47118) );
  NAND U56534 ( .A(n47120), .B(n47119), .Z(n47115) );
  AND U56535 ( .A(n47121), .B(n47122), .Z(n47106) );
  NANDN U56536 ( .A(n47123), .B(n47124), .Z(n47122) );
  NANDN U56537 ( .A(n47125), .B(n47126), .Z(n47124) );
  NANDN U56538 ( .A(n47126), .B(n47125), .Z(n47121) );
  XOR U56539 ( .A(n47120), .B(n47127), .Z(N61218) );
  XOR U56540 ( .A(n47117), .B(n47119), .Z(n47127) );
  XNOR U56541 ( .A(n47113), .B(n47128), .Z(n47119) );
  XNOR U56542 ( .A(n47111), .B(n47114), .Z(n47128) );
  NAND U56543 ( .A(n47129), .B(n47130), .Z(n47114) );
  NAND U56544 ( .A(n47131), .B(n47132), .Z(n47130) );
  OR U56545 ( .A(n47133), .B(n47134), .Z(n47131) );
  NANDN U56546 ( .A(n47135), .B(n47133), .Z(n47129) );
  IV U56547 ( .A(n47134), .Z(n47135) );
  NAND U56548 ( .A(n47136), .B(n47137), .Z(n47111) );
  NAND U56549 ( .A(n47138), .B(n47139), .Z(n47137) );
  NANDN U56550 ( .A(n47140), .B(n47141), .Z(n47138) );
  NANDN U56551 ( .A(n47141), .B(n47140), .Z(n47136) );
  AND U56552 ( .A(n47142), .B(n47143), .Z(n47113) );
  NAND U56553 ( .A(n47144), .B(n47145), .Z(n47143) );
  OR U56554 ( .A(n47146), .B(n47147), .Z(n47144) );
  NANDN U56555 ( .A(n47148), .B(n47146), .Z(n47142) );
  NAND U56556 ( .A(n47149), .B(n47150), .Z(n47117) );
  NANDN U56557 ( .A(n47151), .B(n47152), .Z(n47150) );
  OR U56558 ( .A(n47153), .B(n47154), .Z(n47152) );
  NANDN U56559 ( .A(n47155), .B(n47153), .Z(n47149) );
  IV U56560 ( .A(n47154), .Z(n47155) );
  XNOR U56561 ( .A(n47125), .B(n47156), .Z(n47120) );
  XNOR U56562 ( .A(n47123), .B(n47126), .Z(n47156) );
  NAND U56563 ( .A(n47157), .B(n47158), .Z(n47126) );
  NAND U56564 ( .A(n47159), .B(n47160), .Z(n47158) );
  OR U56565 ( .A(n47161), .B(n47162), .Z(n47159) );
  NANDN U56566 ( .A(n47163), .B(n47161), .Z(n47157) );
  IV U56567 ( .A(n47162), .Z(n47163) );
  NAND U56568 ( .A(n47164), .B(n47165), .Z(n47123) );
  NAND U56569 ( .A(n47166), .B(n47167), .Z(n47165) );
  NANDN U56570 ( .A(n47168), .B(n47169), .Z(n47166) );
  NANDN U56571 ( .A(n47169), .B(n47168), .Z(n47164) );
  AND U56572 ( .A(n47170), .B(n47171), .Z(n47125) );
  NAND U56573 ( .A(n47172), .B(n47173), .Z(n47171) );
  OR U56574 ( .A(n47174), .B(n47175), .Z(n47172) );
  NANDN U56575 ( .A(n47176), .B(n47174), .Z(n47170) );
  XNOR U56576 ( .A(n47151), .B(n47177), .Z(N61217) );
  XOR U56577 ( .A(n47153), .B(n47154), .Z(n47177) );
  XNOR U56578 ( .A(n47167), .B(n47178), .Z(n47154) );
  XOR U56579 ( .A(n47168), .B(n47169), .Z(n47178) );
  XOR U56580 ( .A(n47174), .B(n47179), .Z(n47169) );
  XOR U56581 ( .A(n47173), .B(n47176), .Z(n47179) );
  IV U56582 ( .A(n47175), .Z(n47176) );
  NAND U56583 ( .A(n47180), .B(n47181), .Z(n47175) );
  OR U56584 ( .A(n47182), .B(n47183), .Z(n47181) );
  OR U56585 ( .A(n47184), .B(n47185), .Z(n47180) );
  NAND U56586 ( .A(n47186), .B(n47187), .Z(n47173) );
  OR U56587 ( .A(n47188), .B(n47189), .Z(n47187) );
  OR U56588 ( .A(n47190), .B(n47191), .Z(n47186) );
  NOR U56589 ( .A(n47192), .B(n47193), .Z(n47174) );
  ANDN U56590 ( .B(n47194), .A(n47195), .Z(n47168) );
  XNOR U56591 ( .A(n47161), .B(n47196), .Z(n47167) );
  XNOR U56592 ( .A(n47160), .B(n47162), .Z(n47196) );
  NAND U56593 ( .A(n47197), .B(n47198), .Z(n47162) );
  OR U56594 ( .A(n47199), .B(n47200), .Z(n47198) );
  OR U56595 ( .A(n47201), .B(n47202), .Z(n47197) );
  NAND U56596 ( .A(n47203), .B(n47204), .Z(n47160) );
  OR U56597 ( .A(n47205), .B(n47206), .Z(n47204) );
  OR U56598 ( .A(n47207), .B(n47208), .Z(n47203) );
  ANDN U56599 ( .B(n47209), .A(n47210), .Z(n47161) );
  IV U56600 ( .A(n47211), .Z(n47209) );
  ANDN U56601 ( .B(n47212), .A(n47213), .Z(n47153) );
  XOR U56602 ( .A(n47139), .B(n47214), .Z(n47151) );
  XOR U56603 ( .A(n47140), .B(n47141), .Z(n47214) );
  XOR U56604 ( .A(n47146), .B(n47215), .Z(n47141) );
  XOR U56605 ( .A(n47145), .B(n47148), .Z(n47215) );
  IV U56606 ( .A(n47147), .Z(n47148) );
  NAND U56607 ( .A(n47216), .B(n47217), .Z(n47147) );
  OR U56608 ( .A(n47218), .B(n47219), .Z(n47217) );
  OR U56609 ( .A(n47220), .B(n47221), .Z(n47216) );
  NAND U56610 ( .A(n47222), .B(n47223), .Z(n47145) );
  OR U56611 ( .A(n47224), .B(n47225), .Z(n47223) );
  OR U56612 ( .A(n47226), .B(n47227), .Z(n47222) );
  NOR U56613 ( .A(n47228), .B(n47229), .Z(n47146) );
  ANDN U56614 ( .B(n47230), .A(n47231), .Z(n47140) );
  IV U56615 ( .A(n47232), .Z(n47230) );
  XNOR U56616 ( .A(n47133), .B(n47233), .Z(n47139) );
  XNOR U56617 ( .A(n47132), .B(n47134), .Z(n47233) );
  NAND U56618 ( .A(n47234), .B(n47235), .Z(n47134) );
  OR U56619 ( .A(n47236), .B(n47237), .Z(n47235) );
  OR U56620 ( .A(n47238), .B(n47239), .Z(n47234) );
  NAND U56621 ( .A(n47240), .B(n47241), .Z(n47132) );
  OR U56622 ( .A(n47242), .B(n47243), .Z(n47241) );
  OR U56623 ( .A(n47244), .B(n47245), .Z(n47240) );
  ANDN U56624 ( .B(n47246), .A(n47247), .Z(n47133) );
  IV U56625 ( .A(n47248), .Z(n47246) );
  XNOR U56626 ( .A(n47213), .B(n47212), .Z(N61216) );
  XOR U56627 ( .A(n47232), .B(n47231), .Z(n47212) );
  XNOR U56628 ( .A(n47247), .B(n47248), .Z(n47231) );
  XNOR U56629 ( .A(n47242), .B(n47243), .Z(n47248) );
  XNOR U56630 ( .A(n47244), .B(n47245), .Z(n47243) );
  XNOR U56631 ( .A(y[1165]), .B(x[1165]), .Z(n47245) );
  XNOR U56632 ( .A(y[1166]), .B(x[1166]), .Z(n47244) );
  XNOR U56633 ( .A(y[1164]), .B(x[1164]), .Z(n47242) );
  XNOR U56634 ( .A(n47236), .B(n47237), .Z(n47247) );
  XNOR U56635 ( .A(y[1161]), .B(x[1161]), .Z(n47237) );
  XNOR U56636 ( .A(n47238), .B(n47239), .Z(n47236) );
  XNOR U56637 ( .A(y[1162]), .B(x[1162]), .Z(n47239) );
  XNOR U56638 ( .A(y[1163]), .B(x[1163]), .Z(n47238) );
  XNOR U56639 ( .A(n47229), .B(n47228), .Z(n47232) );
  XNOR U56640 ( .A(n47224), .B(n47225), .Z(n47228) );
  XNOR U56641 ( .A(y[1158]), .B(x[1158]), .Z(n47225) );
  XNOR U56642 ( .A(n47226), .B(n47227), .Z(n47224) );
  XNOR U56643 ( .A(y[1159]), .B(x[1159]), .Z(n47227) );
  XNOR U56644 ( .A(y[1160]), .B(x[1160]), .Z(n47226) );
  XNOR U56645 ( .A(n47218), .B(n47219), .Z(n47229) );
  XNOR U56646 ( .A(y[1155]), .B(x[1155]), .Z(n47219) );
  XNOR U56647 ( .A(n47220), .B(n47221), .Z(n47218) );
  XNOR U56648 ( .A(y[1156]), .B(x[1156]), .Z(n47221) );
  XNOR U56649 ( .A(y[1157]), .B(x[1157]), .Z(n47220) );
  XOR U56650 ( .A(n47194), .B(n47195), .Z(n47213) );
  XNOR U56651 ( .A(n47210), .B(n47211), .Z(n47195) );
  XNOR U56652 ( .A(n47205), .B(n47206), .Z(n47211) );
  XNOR U56653 ( .A(n47207), .B(n47208), .Z(n47206) );
  XNOR U56654 ( .A(y[1153]), .B(x[1153]), .Z(n47208) );
  XNOR U56655 ( .A(y[1154]), .B(x[1154]), .Z(n47207) );
  XNOR U56656 ( .A(y[1152]), .B(x[1152]), .Z(n47205) );
  XNOR U56657 ( .A(n47199), .B(n47200), .Z(n47210) );
  XNOR U56658 ( .A(y[1149]), .B(x[1149]), .Z(n47200) );
  XNOR U56659 ( .A(n47201), .B(n47202), .Z(n47199) );
  XNOR U56660 ( .A(y[1150]), .B(x[1150]), .Z(n47202) );
  XNOR U56661 ( .A(y[1151]), .B(x[1151]), .Z(n47201) );
  XOR U56662 ( .A(n47193), .B(n47192), .Z(n47194) );
  XNOR U56663 ( .A(n47188), .B(n47189), .Z(n47192) );
  XNOR U56664 ( .A(y[1146]), .B(x[1146]), .Z(n47189) );
  XNOR U56665 ( .A(n47190), .B(n47191), .Z(n47188) );
  XNOR U56666 ( .A(y[1147]), .B(x[1147]), .Z(n47191) );
  XNOR U56667 ( .A(y[1148]), .B(x[1148]), .Z(n47190) );
  XNOR U56668 ( .A(n47182), .B(n47183), .Z(n47193) );
  XNOR U56669 ( .A(y[1143]), .B(x[1143]), .Z(n47183) );
  XNOR U56670 ( .A(n47184), .B(n47185), .Z(n47182) );
  XNOR U56671 ( .A(y[1144]), .B(x[1144]), .Z(n47185) );
  XNOR U56672 ( .A(y[1145]), .B(x[1145]), .Z(n47184) );
  NAND U56673 ( .A(n47249), .B(n47250), .Z(N61207) );
  NANDN U56674 ( .A(n47251), .B(n47252), .Z(n47250) );
  OR U56675 ( .A(n47253), .B(n47254), .Z(n47252) );
  NAND U56676 ( .A(n47253), .B(n47254), .Z(n47249) );
  XOR U56677 ( .A(n47253), .B(n47255), .Z(N61206) );
  XNOR U56678 ( .A(n47251), .B(n47254), .Z(n47255) );
  AND U56679 ( .A(n47256), .B(n47257), .Z(n47254) );
  NANDN U56680 ( .A(n47258), .B(n47259), .Z(n47257) );
  NANDN U56681 ( .A(n47260), .B(n47261), .Z(n47259) );
  NANDN U56682 ( .A(n47261), .B(n47260), .Z(n47256) );
  NAND U56683 ( .A(n47262), .B(n47263), .Z(n47251) );
  NANDN U56684 ( .A(n47264), .B(n47265), .Z(n47263) );
  OR U56685 ( .A(n47266), .B(n47267), .Z(n47265) );
  NAND U56686 ( .A(n47267), .B(n47266), .Z(n47262) );
  AND U56687 ( .A(n47268), .B(n47269), .Z(n47253) );
  NANDN U56688 ( .A(n47270), .B(n47271), .Z(n47269) );
  NANDN U56689 ( .A(n47272), .B(n47273), .Z(n47271) );
  NANDN U56690 ( .A(n47273), .B(n47272), .Z(n47268) );
  XOR U56691 ( .A(n47267), .B(n47274), .Z(N61205) );
  XOR U56692 ( .A(n47264), .B(n47266), .Z(n47274) );
  XNOR U56693 ( .A(n47260), .B(n47275), .Z(n47266) );
  XNOR U56694 ( .A(n47258), .B(n47261), .Z(n47275) );
  NAND U56695 ( .A(n47276), .B(n47277), .Z(n47261) );
  NAND U56696 ( .A(n47278), .B(n47279), .Z(n47277) );
  OR U56697 ( .A(n47280), .B(n47281), .Z(n47278) );
  NANDN U56698 ( .A(n47282), .B(n47280), .Z(n47276) );
  IV U56699 ( .A(n47281), .Z(n47282) );
  NAND U56700 ( .A(n47283), .B(n47284), .Z(n47258) );
  NAND U56701 ( .A(n47285), .B(n47286), .Z(n47284) );
  NANDN U56702 ( .A(n47287), .B(n47288), .Z(n47285) );
  NANDN U56703 ( .A(n47288), .B(n47287), .Z(n47283) );
  AND U56704 ( .A(n47289), .B(n47290), .Z(n47260) );
  NAND U56705 ( .A(n47291), .B(n47292), .Z(n47290) );
  OR U56706 ( .A(n47293), .B(n47294), .Z(n47291) );
  NANDN U56707 ( .A(n47295), .B(n47293), .Z(n47289) );
  NAND U56708 ( .A(n47296), .B(n47297), .Z(n47264) );
  NANDN U56709 ( .A(n47298), .B(n47299), .Z(n47297) );
  OR U56710 ( .A(n47300), .B(n47301), .Z(n47299) );
  NANDN U56711 ( .A(n47302), .B(n47300), .Z(n47296) );
  IV U56712 ( .A(n47301), .Z(n47302) );
  XNOR U56713 ( .A(n47272), .B(n47303), .Z(n47267) );
  XNOR U56714 ( .A(n47270), .B(n47273), .Z(n47303) );
  NAND U56715 ( .A(n47304), .B(n47305), .Z(n47273) );
  NAND U56716 ( .A(n47306), .B(n47307), .Z(n47305) );
  OR U56717 ( .A(n47308), .B(n47309), .Z(n47306) );
  NANDN U56718 ( .A(n47310), .B(n47308), .Z(n47304) );
  IV U56719 ( .A(n47309), .Z(n47310) );
  NAND U56720 ( .A(n47311), .B(n47312), .Z(n47270) );
  NAND U56721 ( .A(n47313), .B(n47314), .Z(n47312) );
  NANDN U56722 ( .A(n47315), .B(n47316), .Z(n47313) );
  NANDN U56723 ( .A(n47316), .B(n47315), .Z(n47311) );
  AND U56724 ( .A(n47317), .B(n47318), .Z(n47272) );
  NAND U56725 ( .A(n47319), .B(n47320), .Z(n47318) );
  OR U56726 ( .A(n47321), .B(n47322), .Z(n47319) );
  NANDN U56727 ( .A(n47323), .B(n47321), .Z(n47317) );
  XNOR U56728 ( .A(n47298), .B(n47324), .Z(N61204) );
  XOR U56729 ( .A(n47300), .B(n47301), .Z(n47324) );
  XNOR U56730 ( .A(n47314), .B(n47325), .Z(n47301) );
  XOR U56731 ( .A(n47315), .B(n47316), .Z(n47325) );
  XOR U56732 ( .A(n47321), .B(n47326), .Z(n47316) );
  XOR U56733 ( .A(n47320), .B(n47323), .Z(n47326) );
  IV U56734 ( .A(n47322), .Z(n47323) );
  NAND U56735 ( .A(n47327), .B(n47328), .Z(n47322) );
  OR U56736 ( .A(n47329), .B(n47330), .Z(n47328) );
  OR U56737 ( .A(n47331), .B(n47332), .Z(n47327) );
  NAND U56738 ( .A(n47333), .B(n47334), .Z(n47320) );
  OR U56739 ( .A(n47335), .B(n47336), .Z(n47334) );
  OR U56740 ( .A(n47337), .B(n47338), .Z(n47333) );
  NOR U56741 ( .A(n47339), .B(n47340), .Z(n47321) );
  ANDN U56742 ( .B(n47341), .A(n47342), .Z(n47315) );
  XNOR U56743 ( .A(n47308), .B(n47343), .Z(n47314) );
  XNOR U56744 ( .A(n47307), .B(n47309), .Z(n47343) );
  NAND U56745 ( .A(n47344), .B(n47345), .Z(n47309) );
  OR U56746 ( .A(n47346), .B(n47347), .Z(n47345) );
  OR U56747 ( .A(n47348), .B(n47349), .Z(n47344) );
  NAND U56748 ( .A(n47350), .B(n47351), .Z(n47307) );
  OR U56749 ( .A(n47352), .B(n47353), .Z(n47351) );
  OR U56750 ( .A(n47354), .B(n47355), .Z(n47350) );
  ANDN U56751 ( .B(n47356), .A(n47357), .Z(n47308) );
  IV U56752 ( .A(n47358), .Z(n47356) );
  ANDN U56753 ( .B(n47359), .A(n47360), .Z(n47300) );
  XOR U56754 ( .A(n47286), .B(n47361), .Z(n47298) );
  XOR U56755 ( .A(n47287), .B(n47288), .Z(n47361) );
  XOR U56756 ( .A(n47293), .B(n47362), .Z(n47288) );
  XOR U56757 ( .A(n47292), .B(n47295), .Z(n47362) );
  IV U56758 ( .A(n47294), .Z(n47295) );
  NAND U56759 ( .A(n47363), .B(n47364), .Z(n47294) );
  OR U56760 ( .A(n47365), .B(n47366), .Z(n47364) );
  OR U56761 ( .A(n47367), .B(n47368), .Z(n47363) );
  NAND U56762 ( .A(n47369), .B(n47370), .Z(n47292) );
  OR U56763 ( .A(n47371), .B(n47372), .Z(n47370) );
  OR U56764 ( .A(n47373), .B(n47374), .Z(n47369) );
  NOR U56765 ( .A(n47375), .B(n47376), .Z(n47293) );
  ANDN U56766 ( .B(n47377), .A(n47378), .Z(n47287) );
  IV U56767 ( .A(n47379), .Z(n47377) );
  XNOR U56768 ( .A(n47280), .B(n47380), .Z(n47286) );
  XNOR U56769 ( .A(n47279), .B(n47281), .Z(n47380) );
  NAND U56770 ( .A(n47381), .B(n47382), .Z(n47281) );
  OR U56771 ( .A(n47383), .B(n47384), .Z(n47382) );
  OR U56772 ( .A(n47385), .B(n47386), .Z(n47381) );
  NAND U56773 ( .A(n47387), .B(n47388), .Z(n47279) );
  OR U56774 ( .A(n47389), .B(n47390), .Z(n47388) );
  OR U56775 ( .A(n47391), .B(n47392), .Z(n47387) );
  ANDN U56776 ( .B(n47393), .A(n47394), .Z(n47280) );
  IV U56777 ( .A(n47395), .Z(n47393) );
  XNOR U56778 ( .A(n47360), .B(n47359), .Z(N61203) );
  XOR U56779 ( .A(n47379), .B(n47378), .Z(n47359) );
  XNOR U56780 ( .A(n47394), .B(n47395), .Z(n47378) );
  XNOR U56781 ( .A(n47389), .B(n47390), .Z(n47395) );
  XNOR U56782 ( .A(n47391), .B(n47392), .Z(n47390) );
  XNOR U56783 ( .A(y[1141]), .B(x[1141]), .Z(n47392) );
  XNOR U56784 ( .A(y[1142]), .B(x[1142]), .Z(n47391) );
  XNOR U56785 ( .A(y[1140]), .B(x[1140]), .Z(n47389) );
  XNOR U56786 ( .A(n47383), .B(n47384), .Z(n47394) );
  XNOR U56787 ( .A(y[1137]), .B(x[1137]), .Z(n47384) );
  XNOR U56788 ( .A(n47385), .B(n47386), .Z(n47383) );
  XNOR U56789 ( .A(y[1138]), .B(x[1138]), .Z(n47386) );
  XNOR U56790 ( .A(y[1139]), .B(x[1139]), .Z(n47385) );
  XNOR U56791 ( .A(n47376), .B(n47375), .Z(n47379) );
  XNOR U56792 ( .A(n47371), .B(n47372), .Z(n47375) );
  XNOR U56793 ( .A(y[1134]), .B(x[1134]), .Z(n47372) );
  XNOR U56794 ( .A(n47373), .B(n47374), .Z(n47371) );
  XNOR U56795 ( .A(y[1135]), .B(x[1135]), .Z(n47374) );
  XNOR U56796 ( .A(y[1136]), .B(x[1136]), .Z(n47373) );
  XNOR U56797 ( .A(n47365), .B(n47366), .Z(n47376) );
  XNOR U56798 ( .A(y[1131]), .B(x[1131]), .Z(n47366) );
  XNOR U56799 ( .A(n47367), .B(n47368), .Z(n47365) );
  XNOR U56800 ( .A(y[1132]), .B(x[1132]), .Z(n47368) );
  XNOR U56801 ( .A(y[1133]), .B(x[1133]), .Z(n47367) );
  XOR U56802 ( .A(n47341), .B(n47342), .Z(n47360) );
  XNOR U56803 ( .A(n47357), .B(n47358), .Z(n47342) );
  XNOR U56804 ( .A(n47352), .B(n47353), .Z(n47358) );
  XNOR U56805 ( .A(n47354), .B(n47355), .Z(n47353) );
  XNOR U56806 ( .A(y[1129]), .B(x[1129]), .Z(n47355) );
  XNOR U56807 ( .A(y[1130]), .B(x[1130]), .Z(n47354) );
  XNOR U56808 ( .A(y[1128]), .B(x[1128]), .Z(n47352) );
  XNOR U56809 ( .A(n47346), .B(n47347), .Z(n47357) );
  XNOR U56810 ( .A(y[1125]), .B(x[1125]), .Z(n47347) );
  XNOR U56811 ( .A(n47348), .B(n47349), .Z(n47346) );
  XNOR U56812 ( .A(y[1126]), .B(x[1126]), .Z(n47349) );
  XNOR U56813 ( .A(y[1127]), .B(x[1127]), .Z(n47348) );
  XOR U56814 ( .A(n47340), .B(n47339), .Z(n47341) );
  XNOR U56815 ( .A(n47335), .B(n47336), .Z(n47339) );
  XNOR U56816 ( .A(y[1122]), .B(x[1122]), .Z(n47336) );
  XNOR U56817 ( .A(n47337), .B(n47338), .Z(n47335) );
  XNOR U56818 ( .A(y[1123]), .B(x[1123]), .Z(n47338) );
  XNOR U56819 ( .A(y[1124]), .B(x[1124]), .Z(n47337) );
  XNOR U56820 ( .A(n47329), .B(n47330), .Z(n47340) );
  XNOR U56821 ( .A(y[1119]), .B(x[1119]), .Z(n47330) );
  XNOR U56822 ( .A(n47331), .B(n47332), .Z(n47329) );
  XNOR U56823 ( .A(y[1120]), .B(x[1120]), .Z(n47332) );
  XNOR U56824 ( .A(y[1121]), .B(x[1121]), .Z(n47331) );
  NAND U56825 ( .A(n47396), .B(n47397), .Z(N61194) );
  NANDN U56826 ( .A(n47398), .B(n47399), .Z(n47397) );
  OR U56827 ( .A(n47400), .B(n47401), .Z(n47399) );
  NAND U56828 ( .A(n47400), .B(n47401), .Z(n47396) );
  XOR U56829 ( .A(n47400), .B(n47402), .Z(N61193) );
  XNOR U56830 ( .A(n47398), .B(n47401), .Z(n47402) );
  AND U56831 ( .A(n47403), .B(n47404), .Z(n47401) );
  NANDN U56832 ( .A(n47405), .B(n47406), .Z(n47404) );
  NANDN U56833 ( .A(n47407), .B(n47408), .Z(n47406) );
  NANDN U56834 ( .A(n47408), .B(n47407), .Z(n47403) );
  NAND U56835 ( .A(n47409), .B(n47410), .Z(n47398) );
  NANDN U56836 ( .A(n47411), .B(n47412), .Z(n47410) );
  OR U56837 ( .A(n47413), .B(n47414), .Z(n47412) );
  NAND U56838 ( .A(n47414), .B(n47413), .Z(n47409) );
  AND U56839 ( .A(n47415), .B(n47416), .Z(n47400) );
  NANDN U56840 ( .A(n47417), .B(n47418), .Z(n47416) );
  NANDN U56841 ( .A(n47419), .B(n47420), .Z(n47418) );
  NANDN U56842 ( .A(n47420), .B(n47419), .Z(n47415) );
  XOR U56843 ( .A(n47414), .B(n47421), .Z(N61192) );
  XOR U56844 ( .A(n47411), .B(n47413), .Z(n47421) );
  XNOR U56845 ( .A(n47407), .B(n47422), .Z(n47413) );
  XNOR U56846 ( .A(n47405), .B(n47408), .Z(n47422) );
  NAND U56847 ( .A(n47423), .B(n47424), .Z(n47408) );
  NAND U56848 ( .A(n47425), .B(n47426), .Z(n47424) );
  OR U56849 ( .A(n47427), .B(n47428), .Z(n47425) );
  NANDN U56850 ( .A(n47429), .B(n47427), .Z(n47423) );
  IV U56851 ( .A(n47428), .Z(n47429) );
  NAND U56852 ( .A(n47430), .B(n47431), .Z(n47405) );
  NAND U56853 ( .A(n47432), .B(n47433), .Z(n47431) );
  NANDN U56854 ( .A(n47434), .B(n47435), .Z(n47432) );
  NANDN U56855 ( .A(n47435), .B(n47434), .Z(n47430) );
  AND U56856 ( .A(n47436), .B(n47437), .Z(n47407) );
  NAND U56857 ( .A(n47438), .B(n47439), .Z(n47437) );
  OR U56858 ( .A(n47440), .B(n47441), .Z(n47438) );
  NANDN U56859 ( .A(n47442), .B(n47440), .Z(n47436) );
  NAND U56860 ( .A(n47443), .B(n47444), .Z(n47411) );
  NANDN U56861 ( .A(n47445), .B(n47446), .Z(n47444) );
  OR U56862 ( .A(n47447), .B(n47448), .Z(n47446) );
  NANDN U56863 ( .A(n47449), .B(n47447), .Z(n47443) );
  IV U56864 ( .A(n47448), .Z(n47449) );
  XNOR U56865 ( .A(n47419), .B(n47450), .Z(n47414) );
  XNOR U56866 ( .A(n47417), .B(n47420), .Z(n47450) );
  NAND U56867 ( .A(n47451), .B(n47452), .Z(n47420) );
  NAND U56868 ( .A(n47453), .B(n47454), .Z(n47452) );
  OR U56869 ( .A(n47455), .B(n47456), .Z(n47453) );
  NANDN U56870 ( .A(n47457), .B(n47455), .Z(n47451) );
  IV U56871 ( .A(n47456), .Z(n47457) );
  NAND U56872 ( .A(n47458), .B(n47459), .Z(n47417) );
  NAND U56873 ( .A(n47460), .B(n47461), .Z(n47459) );
  NANDN U56874 ( .A(n47462), .B(n47463), .Z(n47460) );
  NANDN U56875 ( .A(n47463), .B(n47462), .Z(n47458) );
  AND U56876 ( .A(n47464), .B(n47465), .Z(n47419) );
  NAND U56877 ( .A(n47466), .B(n47467), .Z(n47465) );
  OR U56878 ( .A(n47468), .B(n47469), .Z(n47466) );
  NANDN U56879 ( .A(n47470), .B(n47468), .Z(n47464) );
  XNOR U56880 ( .A(n47445), .B(n47471), .Z(N61191) );
  XOR U56881 ( .A(n47447), .B(n47448), .Z(n47471) );
  XNOR U56882 ( .A(n47461), .B(n47472), .Z(n47448) );
  XOR U56883 ( .A(n47462), .B(n47463), .Z(n47472) );
  XOR U56884 ( .A(n47468), .B(n47473), .Z(n47463) );
  XOR U56885 ( .A(n47467), .B(n47470), .Z(n47473) );
  IV U56886 ( .A(n47469), .Z(n47470) );
  NAND U56887 ( .A(n47474), .B(n47475), .Z(n47469) );
  OR U56888 ( .A(n47476), .B(n47477), .Z(n47475) );
  OR U56889 ( .A(n47478), .B(n47479), .Z(n47474) );
  NAND U56890 ( .A(n47480), .B(n47481), .Z(n47467) );
  OR U56891 ( .A(n47482), .B(n47483), .Z(n47481) );
  OR U56892 ( .A(n47484), .B(n47485), .Z(n47480) );
  NOR U56893 ( .A(n47486), .B(n47487), .Z(n47468) );
  ANDN U56894 ( .B(n47488), .A(n47489), .Z(n47462) );
  XNOR U56895 ( .A(n47455), .B(n47490), .Z(n47461) );
  XNOR U56896 ( .A(n47454), .B(n47456), .Z(n47490) );
  NAND U56897 ( .A(n47491), .B(n47492), .Z(n47456) );
  OR U56898 ( .A(n47493), .B(n47494), .Z(n47492) );
  OR U56899 ( .A(n47495), .B(n47496), .Z(n47491) );
  NAND U56900 ( .A(n47497), .B(n47498), .Z(n47454) );
  OR U56901 ( .A(n47499), .B(n47500), .Z(n47498) );
  OR U56902 ( .A(n47501), .B(n47502), .Z(n47497) );
  ANDN U56903 ( .B(n47503), .A(n47504), .Z(n47455) );
  IV U56904 ( .A(n47505), .Z(n47503) );
  ANDN U56905 ( .B(n47506), .A(n47507), .Z(n47447) );
  XOR U56906 ( .A(n47433), .B(n47508), .Z(n47445) );
  XOR U56907 ( .A(n47434), .B(n47435), .Z(n47508) );
  XOR U56908 ( .A(n47440), .B(n47509), .Z(n47435) );
  XOR U56909 ( .A(n47439), .B(n47442), .Z(n47509) );
  IV U56910 ( .A(n47441), .Z(n47442) );
  NAND U56911 ( .A(n47510), .B(n47511), .Z(n47441) );
  OR U56912 ( .A(n47512), .B(n47513), .Z(n47511) );
  OR U56913 ( .A(n47514), .B(n47515), .Z(n47510) );
  NAND U56914 ( .A(n47516), .B(n47517), .Z(n47439) );
  OR U56915 ( .A(n47518), .B(n47519), .Z(n47517) );
  OR U56916 ( .A(n47520), .B(n47521), .Z(n47516) );
  NOR U56917 ( .A(n47522), .B(n47523), .Z(n47440) );
  ANDN U56918 ( .B(n47524), .A(n47525), .Z(n47434) );
  IV U56919 ( .A(n47526), .Z(n47524) );
  XNOR U56920 ( .A(n47427), .B(n47527), .Z(n47433) );
  XNOR U56921 ( .A(n47426), .B(n47428), .Z(n47527) );
  NAND U56922 ( .A(n47528), .B(n47529), .Z(n47428) );
  OR U56923 ( .A(n47530), .B(n47531), .Z(n47529) );
  OR U56924 ( .A(n47532), .B(n47533), .Z(n47528) );
  NAND U56925 ( .A(n47534), .B(n47535), .Z(n47426) );
  OR U56926 ( .A(n47536), .B(n47537), .Z(n47535) );
  OR U56927 ( .A(n47538), .B(n47539), .Z(n47534) );
  ANDN U56928 ( .B(n47540), .A(n47541), .Z(n47427) );
  IV U56929 ( .A(n47542), .Z(n47540) );
  XNOR U56930 ( .A(n47507), .B(n47506), .Z(N61190) );
  XOR U56931 ( .A(n47526), .B(n47525), .Z(n47506) );
  XNOR U56932 ( .A(n47541), .B(n47542), .Z(n47525) );
  XNOR U56933 ( .A(n47536), .B(n47537), .Z(n47542) );
  XNOR U56934 ( .A(n47538), .B(n47539), .Z(n47537) );
  XNOR U56935 ( .A(y[1117]), .B(x[1117]), .Z(n47539) );
  XNOR U56936 ( .A(y[1118]), .B(x[1118]), .Z(n47538) );
  XNOR U56937 ( .A(y[1116]), .B(x[1116]), .Z(n47536) );
  XNOR U56938 ( .A(n47530), .B(n47531), .Z(n47541) );
  XNOR U56939 ( .A(y[1113]), .B(x[1113]), .Z(n47531) );
  XNOR U56940 ( .A(n47532), .B(n47533), .Z(n47530) );
  XNOR U56941 ( .A(y[1114]), .B(x[1114]), .Z(n47533) );
  XNOR U56942 ( .A(y[1115]), .B(x[1115]), .Z(n47532) );
  XNOR U56943 ( .A(n47523), .B(n47522), .Z(n47526) );
  XNOR U56944 ( .A(n47518), .B(n47519), .Z(n47522) );
  XNOR U56945 ( .A(y[1110]), .B(x[1110]), .Z(n47519) );
  XNOR U56946 ( .A(n47520), .B(n47521), .Z(n47518) );
  XNOR U56947 ( .A(y[1111]), .B(x[1111]), .Z(n47521) );
  XNOR U56948 ( .A(y[1112]), .B(x[1112]), .Z(n47520) );
  XNOR U56949 ( .A(n47512), .B(n47513), .Z(n47523) );
  XNOR U56950 ( .A(y[1107]), .B(x[1107]), .Z(n47513) );
  XNOR U56951 ( .A(n47514), .B(n47515), .Z(n47512) );
  XNOR U56952 ( .A(y[1108]), .B(x[1108]), .Z(n47515) );
  XNOR U56953 ( .A(y[1109]), .B(x[1109]), .Z(n47514) );
  XOR U56954 ( .A(n47488), .B(n47489), .Z(n47507) );
  XNOR U56955 ( .A(n47504), .B(n47505), .Z(n47489) );
  XNOR U56956 ( .A(n47499), .B(n47500), .Z(n47505) );
  XNOR U56957 ( .A(n47501), .B(n47502), .Z(n47500) );
  XNOR U56958 ( .A(y[1105]), .B(x[1105]), .Z(n47502) );
  XNOR U56959 ( .A(y[1106]), .B(x[1106]), .Z(n47501) );
  XNOR U56960 ( .A(y[1104]), .B(x[1104]), .Z(n47499) );
  XNOR U56961 ( .A(n47493), .B(n47494), .Z(n47504) );
  XNOR U56962 ( .A(y[1101]), .B(x[1101]), .Z(n47494) );
  XNOR U56963 ( .A(n47495), .B(n47496), .Z(n47493) );
  XNOR U56964 ( .A(y[1102]), .B(x[1102]), .Z(n47496) );
  XNOR U56965 ( .A(y[1103]), .B(x[1103]), .Z(n47495) );
  XOR U56966 ( .A(n47487), .B(n47486), .Z(n47488) );
  XNOR U56967 ( .A(n47482), .B(n47483), .Z(n47486) );
  XNOR U56968 ( .A(y[1098]), .B(x[1098]), .Z(n47483) );
  XNOR U56969 ( .A(n47484), .B(n47485), .Z(n47482) );
  XNOR U56970 ( .A(y[1099]), .B(x[1099]), .Z(n47485) );
  XNOR U56971 ( .A(y[1100]), .B(x[1100]), .Z(n47484) );
  XNOR U56972 ( .A(n47476), .B(n47477), .Z(n47487) );
  XNOR U56973 ( .A(y[1095]), .B(x[1095]), .Z(n47477) );
  XNOR U56974 ( .A(n47478), .B(n47479), .Z(n47476) );
  XNOR U56975 ( .A(y[1096]), .B(x[1096]), .Z(n47479) );
  XNOR U56976 ( .A(y[1097]), .B(x[1097]), .Z(n47478) );
  NAND U56977 ( .A(n47543), .B(n47544), .Z(N61181) );
  NANDN U56978 ( .A(n47545), .B(n47546), .Z(n47544) );
  OR U56979 ( .A(n47547), .B(n47548), .Z(n47546) );
  NAND U56980 ( .A(n47547), .B(n47548), .Z(n47543) );
  XOR U56981 ( .A(n47547), .B(n47549), .Z(N61180) );
  XNOR U56982 ( .A(n47545), .B(n47548), .Z(n47549) );
  AND U56983 ( .A(n47550), .B(n47551), .Z(n47548) );
  NANDN U56984 ( .A(n47552), .B(n47553), .Z(n47551) );
  NANDN U56985 ( .A(n47554), .B(n47555), .Z(n47553) );
  NANDN U56986 ( .A(n47555), .B(n47554), .Z(n47550) );
  NAND U56987 ( .A(n47556), .B(n47557), .Z(n47545) );
  NANDN U56988 ( .A(n47558), .B(n47559), .Z(n47557) );
  OR U56989 ( .A(n47560), .B(n47561), .Z(n47559) );
  NAND U56990 ( .A(n47561), .B(n47560), .Z(n47556) );
  AND U56991 ( .A(n47562), .B(n47563), .Z(n47547) );
  NANDN U56992 ( .A(n47564), .B(n47565), .Z(n47563) );
  NANDN U56993 ( .A(n47566), .B(n47567), .Z(n47565) );
  NANDN U56994 ( .A(n47567), .B(n47566), .Z(n47562) );
  XOR U56995 ( .A(n47561), .B(n47568), .Z(N61179) );
  XOR U56996 ( .A(n47558), .B(n47560), .Z(n47568) );
  XNOR U56997 ( .A(n47554), .B(n47569), .Z(n47560) );
  XNOR U56998 ( .A(n47552), .B(n47555), .Z(n47569) );
  NAND U56999 ( .A(n47570), .B(n47571), .Z(n47555) );
  NAND U57000 ( .A(n47572), .B(n47573), .Z(n47571) );
  OR U57001 ( .A(n47574), .B(n47575), .Z(n47572) );
  NANDN U57002 ( .A(n47576), .B(n47574), .Z(n47570) );
  IV U57003 ( .A(n47575), .Z(n47576) );
  NAND U57004 ( .A(n47577), .B(n47578), .Z(n47552) );
  NAND U57005 ( .A(n47579), .B(n47580), .Z(n47578) );
  NANDN U57006 ( .A(n47581), .B(n47582), .Z(n47579) );
  NANDN U57007 ( .A(n47582), .B(n47581), .Z(n47577) );
  AND U57008 ( .A(n47583), .B(n47584), .Z(n47554) );
  NAND U57009 ( .A(n47585), .B(n47586), .Z(n47584) );
  OR U57010 ( .A(n47587), .B(n47588), .Z(n47585) );
  NANDN U57011 ( .A(n47589), .B(n47587), .Z(n47583) );
  NAND U57012 ( .A(n47590), .B(n47591), .Z(n47558) );
  NANDN U57013 ( .A(n47592), .B(n47593), .Z(n47591) );
  OR U57014 ( .A(n47594), .B(n47595), .Z(n47593) );
  NANDN U57015 ( .A(n47596), .B(n47594), .Z(n47590) );
  IV U57016 ( .A(n47595), .Z(n47596) );
  XNOR U57017 ( .A(n47566), .B(n47597), .Z(n47561) );
  XNOR U57018 ( .A(n47564), .B(n47567), .Z(n47597) );
  NAND U57019 ( .A(n47598), .B(n47599), .Z(n47567) );
  NAND U57020 ( .A(n47600), .B(n47601), .Z(n47599) );
  OR U57021 ( .A(n47602), .B(n47603), .Z(n47600) );
  NANDN U57022 ( .A(n47604), .B(n47602), .Z(n47598) );
  IV U57023 ( .A(n47603), .Z(n47604) );
  NAND U57024 ( .A(n47605), .B(n47606), .Z(n47564) );
  NAND U57025 ( .A(n47607), .B(n47608), .Z(n47606) );
  NANDN U57026 ( .A(n47609), .B(n47610), .Z(n47607) );
  NANDN U57027 ( .A(n47610), .B(n47609), .Z(n47605) );
  AND U57028 ( .A(n47611), .B(n47612), .Z(n47566) );
  NAND U57029 ( .A(n47613), .B(n47614), .Z(n47612) );
  OR U57030 ( .A(n47615), .B(n47616), .Z(n47613) );
  NANDN U57031 ( .A(n47617), .B(n47615), .Z(n47611) );
  XNOR U57032 ( .A(n47592), .B(n47618), .Z(N61178) );
  XOR U57033 ( .A(n47594), .B(n47595), .Z(n47618) );
  XNOR U57034 ( .A(n47608), .B(n47619), .Z(n47595) );
  XOR U57035 ( .A(n47609), .B(n47610), .Z(n47619) );
  XOR U57036 ( .A(n47615), .B(n47620), .Z(n47610) );
  XOR U57037 ( .A(n47614), .B(n47617), .Z(n47620) );
  IV U57038 ( .A(n47616), .Z(n47617) );
  NAND U57039 ( .A(n47621), .B(n47622), .Z(n47616) );
  OR U57040 ( .A(n47623), .B(n47624), .Z(n47622) );
  OR U57041 ( .A(n47625), .B(n47626), .Z(n47621) );
  NAND U57042 ( .A(n47627), .B(n47628), .Z(n47614) );
  OR U57043 ( .A(n47629), .B(n47630), .Z(n47628) );
  OR U57044 ( .A(n47631), .B(n47632), .Z(n47627) );
  NOR U57045 ( .A(n47633), .B(n47634), .Z(n47615) );
  ANDN U57046 ( .B(n47635), .A(n47636), .Z(n47609) );
  XNOR U57047 ( .A(n47602), .B(n47637), .Z(n47608) );
  XNOR U57048 ( .A(n47601), .B(n47603), .Z(n47637) );
  NAND U57049 ( .A(n47638), .B(n47639), .Z(n47603) );
  OR U57050 ( .A(n47640), .B(n47641), .Z(n47639) );
  OR U57051 ( .A(n47642), .B(n47643), .Z(n47638) );
  NAND U57052 ( .A(n47644), .B(n47645), .Z(n47601) );
  OR U57053 ( .A(n47646), .B(n47647), .Z(n47645) );
  OR U57054 ( .A(n47648), .B(n47649), .Z(n47644) );
  ANDN U57055 ( .B(n47650), .A(n47651), .Z(n47602) );
  IV U57056 ( .A(n47652), .Z(n47650) );
  ANDN U57057 ( .B(n47653), .A(n47654), .Z(n47594) );
  XOR U57058 ( .A(n47580), .B(n47655), .Z(n47592) );
  XOR U57059 ( .A(n47581), .B(n47582), .Z(n47655) );
  XOR U57060 ( .A(n47587), .B(n47656), .Z(n47582) );
  XOR U57061 ( .A(n47586), .B(n47589), .Z(n47656) );
  IV U57062 ( .A(n47588), .Z(n47589) );
  NAND U57063 ( .A(n47657), .B(n47658), .Z(n47588) );
  OR U57064 ( .A(n47659), .B(n47660), .Z(n47658) );
  OR U57065 ( .A(n47661), .B(n47662), .Z(n47657) );
  NAND U57066 ( .A(n47663), .B(n47664), .Z(n47586) );
  OR U57067 ( .A(n47665), .B(n47666), .Z(n47664) );
  OR U57068 ( .A(n47667), .B(n47668), .Z(n47663) );
  NOR U57069 ( .A(n47669), .B(n47670), .Z(n47587) );
  ANDN U57070 ( .B(n47671), .A(n47672), .Z(n47581) );
  IV U57071 ( .A(n47673), .Z(n47671) );
  XNOR U57072 ( .A(n47574), .B(n47674), .Z(n47580) );
  XNOR U57073 ( .A(n47573), .B(n47575), .Z(n47674) );
  NAND U57074 ( .A(n47675), .B(n47676), .Z(n47575) );
  OR U57075 ( .A(n47677), .B(n47678), .Z(n47676) );
  OR U57076 ( .A(n47679), .B(n47680), .Z(n47675) );
  NAND U57077 ( .A(n47681), .B(n47682), .Z(n47573) );
  OR U57078 ( .A(n47683), .B(n47684), .Z(n47682) );
  OR U57079 ( .A(n47685), .B(n47686), .Z(n47681) );
  ANDN U57080 ( .B(n47687), .A(n47688), .Z(n47574) );
  IV U57081 ( .A(n47689), .Z(n47687) );
  XNOR U57082 ( .A(n47654), .B(n47653), .Z(N61177) );
  XOR U57083 ( .A(n47673), .B(n47672), .Z(n47653) );
  XNOR U57084 ( .A(n47688), .B(n47689), .Z(n47672) );
  XNOR U57085 ( .A(n47683), .B(n47684), .Z(n47689) );
  XNOR U57086 ( .A(n47685), .B(n47686), .Z(n47684) );
  XNOR U57087 ( .A(y[1093]), .B(x[1093]), .Z(n47686) );
  XNOR U57088 ( .A(y[1094]), .B(x[1094]), .Z(n47685) );
  XNOR U57089 ( .A(y[1092]), .B(x[1092]), .Z(n47683) );
  XNOR U57090 ( .A(n47677), .B(n47678), .Z(n47688) );
  XNOR U57091 ( .A(y[1089]), .B(x[1089]), .Z(n47678) );
  XNOR U57092 ( .A(n47679), .B(n47680), .Z(n47677) );
  XNOR U57093 ( .A(y[1090]), .B(x[1090]), .Z(n47680) );
  XNOR U57094 ( .A(y[1091]), .B(x[1091]), .Z(n47679) );
  XNOR U57095 ( .A(n47670), .B(n47669), .Z(n47673) );
  XNOR U57096 ( .A(n47665), .B(n47666), .Z(n47669) );
  XNOR U57097 ( .A(y[1086]), .B(x[1086]), .Z(n47666) );
  XNOR U57098 ( .A(n47667), .B(n47668), .Z(n47665) );
  XNOR U57099 ( .A(y[1087]), .B(x[1087]), .Z(n47668) );
  XNOR U57100 ( .A(y[1088]), .B(x[1088]), .Z(n47667) );
  XNOR U57101 ( .A(n47659), .B(n47660), .Z(n47670) );
  XNOR U57102 ( .A(y[1083]), .B(x[1083]), .Z(n47660) );
  XNOR U57103 ( .A(n47661), .B(n47662), .Z(n47659) );
  XNOR U57104 ( .A(y[1084]), .B(x[1084]), .Z(n47662) );
  XNOR U57105 ( .A(y[1085]), .B(x[1085]), .Z(n47661) );
  XOR U57106 ( .A(n47635), .B(n47636), .Z(n47654) );
  XNOR U57107 ( .A(n47651), .B(n47652), .Z(n47636) );
  XNOR U57108 ( .A(n47646), .B(n47647), .Z(n47652) );
  XNOR U57109 ( .A(n47648), .B(n47649), .Z(n47647) );
  XNOR U57110 ( .A(y[1081]), .B(x[1081]), .Z(n47649) );
  XNOR U57111 ( .A(y[1082]), .B(x[1082]), .Z(n47648) );
  XNOR U57112 ( .A(y[1080]), .B(x[1080]), .Z(n47646) );
  XNOR U57113 ( .A(n47640), .B(n47641), .Z(n47651) );
  XNOR U57114 ( .A(y[1077]), .B(x[1077]), .Z(n47641) );
  XNOR U57115 ( .A(n47642), .B(n47643), .Z(n47640) );
  XNOR U57116 ( .A(y[1078]), .B(x[1078]), .Z(n47643) );
  XNOR U57117 ( .A(y[1079]), .B(x[1079]), .Z(n47642) );
  XOR U57118 ( .A(n47634), .B(n47633), .Z(n47635) );
  XNOR U57119 ( .A(n47629), .B(n47630), .Z(n47633) );
  XNOR U57120 ( .A(y[1074]), .B(x[1074]), .Z(n47630) );
  XNOR U57121 ( .A(n47631), .B(n47632), .Z(n47629) );
  XNOR U57122 ( .A(y[1075]), .B(x[1075]), .Z(n47632) );
  XNOR U57123 ( .A(y[1076]), .B(x[1076]), .Z(n47631) );
  XNOR U57124 ( .A(n47623), .B(n47624), .Z(n47634) );
  XNOR U57125 ( .A(y[1071]), .B(x[1071]), .Z(n47624) );
  XNOR U57126 ( .A(n47625), .B(n47626), .Z(n47623) );
  XNOR U57127 ( .A(y[1072]), .B(x[1072]), .Z(n47626) );
  XNOR U57128 ( .A(y[1073]), .B(x[1073]), .Z(n47625) );
  NAND U57129 ( .A(n47690), .B(n47691), .Z(N61168) );
  NANDN U57130 ( .A(n47692), .B(n47693), .Z(n47691) );
  OR U57131 ( .A(n47694), .B(n47695), .Z(n47693) );
  NAND U57132 ( .A(n47694), .B(n47695), .Z(n47690) );
  XOR U57133 ( .A(n47694), .B(n47696), .Z(N61167) );
  XNOR U57134 ( .A(n47692), .B(n47695), .Z(n47696) );
  AND U57135 ( .A(n47697), .B(n47698), .Z(n47695) );
  NANDN U57136 ( .A(n47699), .B(n47700), .Z(n47698) );
  NANDN U57137 ( .A(n47701), .B(n47702), .Z(n47700) );
  NANDN U57138 ( .A(n47702), .B(n47701), .Z(n47697) );
  NAND U57139 ( .A(n47703), .B(n47704), .Z(n47692) );
  NANDN U57140 ( .A(n47705), .B(n47706), .Z(n47704) );
  OR U57141 ( .A(n47707), .B(n47708), .Z(n47706) );
  NAND U57142 ( .A(n47708), .B(n47707), .Z(n47703) );
  AND U57143 ( .A(n47709), .B(n47710), .Z(n47694) );
  NANDN U57144 ( .A(n47711), .B(n47712), .Z(n47710) );
  NANDN U57145 ( .A(n47713), .B(n47714), .Z(n47712) );
  NANDN U57146 ( .A(n47714), .B(n47713), .Z(n47709) );
  XOR U57147 ( .A(n47708), .B(n47715), .Z(N61166) );
  XOR U57148 ( .A(n47705), .B(n47707), .Z(n47715) );
  XNOR U57149 ( .A(n47701), .B(n47716), .Z(n47707) );
  XNOR U57150 ( .A(n47699), .B(n47702), .Z(n47716) );
  NAND U57151 ( .A(n47717), .B(n47718), .Z(n47702) );
  NAND U57152 ( .A(n47719), .B(n47720), .Z(n47718) );
  OR U57153 ( .A(n47721), .B(n47722), .Z(n47719) );
  NANDN U57154 ( .A(n47723), .B(n47721), .Z(n47717) );
  IV U57155 ( .A(n47722), .Z(n47723) );
  NAND U57156 ( .A(n47724), .B(n47725), .Z(n47699) );
  NAND U57157 ( .A(n47726), .B(n47727), .Z(n47725) );
  NANDN U57158 ( .A(n47728), .B(n47729), .Z(n47726) );
  NANDN U57159 ( .A(n47729), .B(n47728), .Z(n47724) );
  AND U57160 ( .A(n47730), .B(n47731), .Z(n47701) );
  NAND U57161 ( .A(n47732), .B(n47733), .Z(n47731) );
  OR U57162 ( .A(n47734), .B(n47735), .Z(n47732) );
  NANDN U57163 ( .A(n47736), .B(n47734), .Z(n47730) );
  NAND U57164 ( .A(n47737), .B(n47738), .Z(n47705) );
  NANDN U57165 ( .A(n47739), .B(n47740), .Z(n47738) );
  OR U57166 ( .A(n47741), .B(n47742), .Z(n47740) );
  NANDN U57167 ( .A(n47743), .B(n47741), .Z(n47737) );
  IV U57168 ( .A(n47742), .Z(n47743) );
  XNOR U57169 ( .A(n47713), .B(n47744), .Z(n47708) );
  XNOR U57170 ( .A(n47711), .B(n47714), .Z(n47744) );
  NAND U57171 ( .A(n47745), .B(n47746), .Z(n47714) );
  NAND U57172 ( .A(n47747), .B(n47748), .Z(n47746) );
  OR U57173 ( .A(n47749), .B(n47750), .Z(n47747) );
  NANDN U57174 ( .A(n47751), .B(n47749), .Z(n47745) );
  IV U57175 ( .A(n47750), .Z(n47751) );
  NAND U57176 ( .A(n47752), .B(n47753), .Z(n47711) );
  NAND U57177 ( .A(n47754), .B(n47755), .Z(n47753) );
  NANDN U57178 ( .A(n47756), .B(n47757), .Z(n47754) );
  NANDN U57179 ( .A(n47757), .B(n47756), .Z(n47752) );
  AND U57180 ( .A(n47758), .B(n47759), .Z(n47713) );
  NAND U57181 ( .A(n47760), .B(n47761), .Z(n47759) );
  OR U57182 ( .A(n47762), .B(n47763), .Z(n47760) );
  NANDN U57183 ( .A(n47764), .B(n47762), .Z(n47758) );
  XNOR U57184 ( .A(n47739), .B(n47765), .Z(N61165) );
  XOR U57185 ( .A(n47741), .B(n47742), .Z(n47765) );
  XNOR U57186 ( .A(n47755), .B(n47766), .Z(n47742) );
  XOR U57187 ( .A(n47756), .B(n47757), .Z(n47766) );
  XOR U57188 ( .A(n47762), .B(n47767), .Z(n47757) );
  XOR U57189 ( .A(n47761), .B(n47764), .Z(n47767) );
  IV U57190 ( .A(n47763), .Z(n47764) );
  NAND U57191 ( .A(n47768), .B(n47769), .Z(n47763) );
  OR U57192 ( .A(n47770), .B(n47771), .Z(n47769) );
  OR U57193 ( .A(n47772), .B(n47773), .Z(n47768) );
  NAND U57194 ( .A(n47774), .B(n47775), .Z(n47761) );
  OR U57195 ( .A(n47776), .B(n47777), .Z(n47775) );
  OR U57196 ( .A(n47778), .B(n47779), .Z(n47774) );
  NOR U57197 ( .A(n47780), .B(n47781), .Z(n47762) );
  ANDN U57198 ( .B(n47782), .A(n47783), .Z(n47756) );
  XNOR U57199 ( .A(n47749), .B(n47784), .Z(n47755) );
  XNOR U57200 ( .A(n47748), .B(n47750), .Z(n47784) );
  NAND U57201 ( .A(n47785), .B(n47786), .Z(n47750) );
  OR U57202 ( .A(n47787), .B(n47788), .Z(n47786) );
  OR U57203 ( .A(n47789), .B(n47790), .Z(n47785) );
  NAND U57204 ( .A(n47791), .B(n47792), .Z(n47748) );
  OR U57205 ( .A(n47793), .B(n47794), .Z(n47792) );
  OR U57206 ( .A(n47795), .B(n47796), .Z(n47791) );
  ANDN U57207 ( .B(n47797), .A(n47798), .Z(n47749) );
  IV U57208 ( .A(n47799), .Z(n47797) );
  ANDN U57209 ( .B(n47800), .A(n47801), .Z(n47741) );
  XOR U57210 ( .A(n47727), .B(n47802), .Z(n47739) );
  XOR U57211 ( .A(n47728), .B(n47729), .Z(n47802) );
  XOR U57212 ( .A(n47734), .B(n47803), .Z(n47729) );
  XOR U57213 ( .A(n47733), .B(n47736), .Z(n47803) );
  IV U57214 ( .A(n47735), .Z(n47736) );
  NAND U57215 ( .A(n47804), .B(n47805), .Z(n47735) );
  OR U57216 ( .A(n47806), .B(n47807), .Z(n47805) );
  OR U57217 ( .A(n47808), .B(n47809), .Z(n47804) );
  NAND U57218 ( .A(n47810), .B(n47811), .Z(n47733) );
  OR U57219 ( .A(n47812), .B(n47813), .Z(n47811) );
  OR U57220 ( .A(n47814), .B(n47815), .Z(n47810) );
  NOR U57221 ( .A(n47816), .B(n47817), .Z(n47734) );
  ANDN U57222 ( .B(n47818), .A(n47819), .Z(n47728) );
  IV U57223 ( .A(n47820), .Z(n47818) );
  XNOR U57224 ( .A(n47721), .B(n47821), .Z(n47727) );
  XNOR U57225 ( .A(n47720), .B(n47722), .Z(n47821) );
  NAND U57226 ( .A(n47822), .B(n47823), .Z(n47722) );
  OR U57227 ( .A(n47824), .B(n47825), .Z(n47823) );
  OR U57228 ( .A(n47826), .B(n47827), .Z(n47822) );
  NAND U57229 ( .A(n47828), .B(n47829), .Z(n47720) );
  OR U57230 ( .A(n47830), .B(n47831), .Z(n47829) );
  OR U57231 ( .A(n47832), .B(n47833), .Z(n47828) );
  ANDN U57232 ( .B(n47834), .A(n47835), .Z(n47721) );
  IV U57233 ( .A(n47836), .Z(n47834) );
  XNOR U57234 ( .A(n47801), .B(n47800), .Z(N61164) );
  XOR U57235 ( .A(n47820), .B(n47819), .Z(n47800) );
  XNOR U57236 ( .A(n47835), .B(n47836), .Z(n47819) );
  XNOR U57237 ( .A(n47830), .B(n47831), .Z(n47836) );
  XNOR U57238 ( .A(n47832), .B(n47833), .Z(n47831) );
  XNOR U57239 ( .A(y[1069]), .B(x[1069]), .Z(n47833) );
  XNOR U57240 ( .A(y[1070]), .B(x[1070]), .Z(n47832) );
  XNOR U57241 ( .A(y[1068]), .B(x[1068]), .Z(n47830) );
  XNOR U57242 ( .A(n47824), .B(n47825), .Z(n47835) );
  XNOR U57243 ( .A(y[1065]), .B(x[1065]), .Z(n47825) );
  XNOR U57244 ( .A(n47826), .B(n47827), .Z(n47824) );
  XNOR U57245 ( .A(y[1066]), .B(x[1066]), .Z(n47827) );
  XNOR U57246 ( .A(y[1067]), .B(x[1067]), .Z(n47826) );
  XNOR U57247 ( .A(n47817), .B(n47816), .Z(n47820) );
  XNOR U57248 ( .A(n47812), .B(n47813), .Z(n47816) );
  XNOR U57249 ( .A(y[1062]), .B(x[1062]), .Z(n47813) );
  XNOR U57250 ( .A(n47814), .B(n47815), .Z(n47812) );
  XNOR U57251 ( .A(y[1063]), .B(x[1063]), .Z(n47815) );
  XNOR U57252 ( .A(y[1064]), .B(x[1064]), .Z(n47814) );
  XNOR U57253 ( .A(n47806), .B(n47807), .Z(n47817) );
  XNOR U57254 ( .A(y[1059]), .B(x[1059]), .Z(n47807) );
  XNOR U57255 ( .A(n47808), .B(n47809), .Z(n47806) );
  XNOR U57256 ( .A(y[1060]), .B(x[1060]), .Z(n47809) );
  XNOR U57257 ( .A(y[1061]), .B(x[1061]), .Z(n47808) );
  XOR U57258 ( .A(n47782), .B(n47783), .Z(n47801) );
  XNOR U57259 ( .A(n47798), .B(n47799), .Z(n47783) );
  XNOR U57260 ( .A(n47793), .B(n47794), .Z(n47799) );
  XNOR U57261 ( .A(n47795), .B(n47796), .Z(n47794) );
  XNOR U57262 ( .A(y[1057]), .B(x[1057]), .Z(n47796) );
  XNOR U57263 ( .A(y[1058]), .B(x[1058]), .Z(n47795) );
  XNOR U57264 ( .A(y[1056]), .B(x[1056]), .Z(n47793) );
  XNOR U57265 ( .A(n47787), .B(n47788), .Z(n47798) );
  XNOR U57266 ( .A(y[1053]), .B(x[1053]), .Z(n47788) );
  XNOR U57267 ( .A(n47789), .B(n47790), .Z(n47787) );
  XNOR U57268 ( .A(y[1054]), .B(x[1054]), .Z(n47790) );
  XNOR U57269 ( .A(y[1055]), .B(x[1055]), .Z(n47789) );
  XOR U57270 ( .A(n47781), .B(n47780), .Z(n47782) );
  XNOR U57271 ( .A(n47776), .B(n47777), .Z(n47780) );
  XNOR U57272 ( .A(y[1050]), .B(x[1050]), .Z(n47777) );
  XNOR U57273 ( .A(n47778), .B(n47779), .Z(n47776) );
  XNOR U57274 ( .A(y[1051]), .B(x[1051]), .Z(n47779) );
  XNOR U57275 ( .A(y[1052]), .B(x[1052]), .Z(n47778) );
  XNOR U57276 ( .A(n47770), .B(n47771), .Z(n47781) );
  XNOR U57277 ( .A(y[1047]), .B(x[1047]), .Z(n47771) );
  XNOR U57278 ( .A(n47772), .B(n47773), .Z(n47770) );
  XNOR U57279 ( .A(y[1048]), .B(x[1048]), .Z(n47773) );
  XNOR U57280 ( .A(y[1049]), .B(x[1049]), .Z(n47772) );
  NAND U57281 ( .A(n47837), .B(n47838), .Z(N61155) );
  NANDN U57282 ( .A(n47839), .B(n47840), .Z(n47838) );
  OR U57283 ( .A(n47841), .B(n47842), .Z(n47840) );
  NAND U57284 ( .A(n47841), .B(n47842), .Z(n47837) );
  XOR U57285 ( .A(n47841), .B(n47843), .Z(N61154) );
  XNOR U57286 ( .A(n47839), .B(n47842), .Z(n47843) );
  AND U57287 ( .A(n47844), .B(n47845), .Z(n47842) );
  NANDN U57288 ( .A(n47846), .B(n47847), .Z(n47845) );
  NANDN U57289 ( .A(n47848), .B(n47849), .Z(n47847) );
  NANDN U57290 ( .A(n47849), .B(n47848), .Z(n47844) );
  NAND U57291 ( .A(n47850), .B(n47851), .Z(n47839) );
  NANDN U57292 ( .A(n47852), .B(n47853), .Z(n47851) );
  OR U57293 ( .A(n47854), .B(n47855), .Z(n47853) );
  NAND U57294 ( .A(n47855), .B(n47854), .Z(n47850) );
  AND U57295 ( .A(n47856), .B(n47857), .Z(n47841) );
  NANDN U57296 ( .A(n47858), .B(n47859), .Z(n47857) );
  NANDN U57297 ( .A(n47860), .B(n47861), .Z(n47859) );
  NANDN U57298 ( .A(n47861), .B(n47860), .Z(n47856) );
  XOR U57299 ( .A(n47855), .B(n47862), .Z(N61153) );
  XOR U57300 ( .A(n47852), .B(n47854), .Z(n47862) );
  XNOR U57301 ( .A(n47848), .B(n47863), .Z(n47854) );
  XNOR U57302 ( .A(n47846), .B(n47849), .Z(n47863) );
  NAND U57303 ( .A(n47864), .B(n47865), .Z(n47849) );
  NAND U57304 ( .A(n47866), .B(n47867), .Z(n47865) );
  OR U57305 ( .A(n47868), .B(n47869), .Z(n47866) );
  NANDN U57306 ( .A(n47870), .B(n47868), .Z(n47864) );
  IV U57307 ( .A(n47869), .Z(n47870) );
  NAND U57308 ( .A(n47871), .B(n47872), .Z(n47846) );
  NAND U57309 ( .A(n47873), .B(n47874), .Z(n47872) );
  NANDN U57310 ( .A(n47875), .B(n47876), .Z(n47873) );
  NANDN U57311 ( .A(n47876), .B(n47875), .Z(n47871) );
  AND U57312 ( .A(n47877), .B(n47878), .Z(n47848) );
  NAND U57313 ( .A(n47879), .B(n47880), .Z(n47878) );
  OR U57314 ( .A(n47881), .B(n47882), .Z(n47879) );
  NANDN U57315 ( .A(n47883), .B(n47881), .Z(n47877) );
  NAND U57316 ( .A(n47884), .B(n47885), .Z(n47852) );
  NANDN U57317 ( .A(n47886), .B(n47887), .Z(n47885) );
  OR U57318 ( .A(n47888), .B(n47889), .Z(n47887) );
  NANDN U57319 ( .A(n47890), .B(n47888), .Z(n47884) );
  IV U57320 ( .A(n47889), .Z(n47890) );
  XNOR U57321 ( .A(n47860), .B(n47891), .Z(n47855) );
  XNOR U57322 ( .A(n47858), .B(n47861), .Z(n47891) );
  NAND U57323 ( .A(n47892), .B(n47893), .Z(n47861) );
  NAND U57324 ( .A(n47894), .B(n47895), .Z(n47893) );
  OR U57325 ( .A(n47896), .B(n47897), .Z(n47894) );
  NANDN U57326 ( .A(n47898), .B(n47896), .Z(n47892) );
  IV U57327 ( .A(n47897), .Z(n47898) );
  NAND U57328 ( .A(n47899), .B(n47900), .Z(n47858) );
  NAND U57329 ( .A(n47901), .B(n47902), .Z(n47900) );
  NANDN U57330 ( .A(n47903), .B(n47904), .Z(n47901) );
  NANDN U57331 ( .A(n47904), .B(n47903), .Z(n47899) );
  AND U57332 ( .A(n47905), .B(n47906), .Z(n47860) );
  NAND U57333 ( .A(n47907), .B(n47908), .Z(n47906) );
  OR U57334 ( .A(n47909), .B(n47910), .Z(n47907) );
  NANDN U57335 ( .A(n47911), .B(n47909), .Z(n47905) );
  XNOR U57336 ( .A(n47886), .B(n47912), .Z(N61152) );
  XOR U57337 ( .A(n47888), .B(n47889), .Z(n47912) );
  XNOR U57338 ( .A(n47902), .B(n47913), .Z(n47889) );
  XOR U57339 ( .A(n47903), .B(n47904), .Z(n47913) );
  XOR U57340 ( .A(n47909), .B(n47914), .Z(n47904) );
  XOR U57341 ( .A(n47908), .B(n47911), .Z(n47914) );
  IV U57342 ( .A(n47910), .Z(n47911) );
  NAND U57343 ( .A(n47915), .B(n47916), .Z(n47910) );
  OR U57344 ( .A(n47917), .B(n47918), .Z(n47916) );
  OR U57345 ( .A(n47919), .B(n47920), .Z(n47915) );
  NAND U57346 ( .A(n47921), .B(n47922), .Z(n47908) );
  OR U57347 ( .A(n47923), .B(n47924), .Z(n47922) );
  OR U57348 ( .A(n47925), .B(n47926), .Z(n47921) );
  NOR U57349 ( .A(n47927), .B(n47928), .Z(n47909) );
  ANDN U57350 ( .B(n47929), .A(n47930), .Z(n47903) );
  XNOR U57351 ( .A(n47896), .B(n47931), .Z(n47902) );
  XNOR U57352 ( .A(n47895), .B(n47897), .Z(n47931) );
  NAND U57353 ( .A(n47932), .B(n47933), .Z(n47897) );
  OR U57354 ( .A(n47934), .B(n47935), .Z(n47933) );
  OR U57355 ( .A(n47936), .B(n47937), .Z(n47932) );
  NAND U57356 ( .A(n47938), .B(n47939), .Z(n47895) );
  OR U57357 ( .A(n47940), .B(n47941), .Z(n47939) );
  OR U57358 ( .A(n47942), .B(n47943), .Z(n47938) );
  ANDN U57359 ( .B(n47944), .A(n47945), .Z(n47896) );
  IV U57360 ( .A(n47946), .Z(n47944) );
  ANDN U57361 ( .B(n47947), .A(n47948), .Z(n47888) );
  XOR U57362 ( .A(n47874), .B(n47949), .Z(n47886) );
  XOR U57363 ( .A(n47875), .B(n47876), .Z(n47949) );
  XOR U57364 ( .A(n47881), .B(n47950), .Z(n47876) );
  XOR U57365 ( .A(n47880), .B(n47883), .Z(n47950) );
  IV U57366 ( .A(n47882), .Z(n47883) );
  NAND U57367 ( .A(n47951), .B(n47952), .Z(n47882) );
  OR U57368 ( .A(n47953), .B(n47954), .Z(n47952) );
  OR U57369 ( .A(n47955), .B(n47956), .Z(n47951) );
  NAND U57370 ( .A(n47957), .B(n47958), .Z(n47880) );
  OR U57371 ( .A(n47959), .B(n47960), .Z(n47958) );
  OR U57372 ( .A(n47961), .B(n47962), .Z(n47957) );
  NOR U57373 ( .A(n47963), .B(n47964), .Z(n47881) );
  ANDN U57374 ( .B(n47965), .A(n47966), .Z(n47875) );
  IV U57375 ( .A(n47967), .Z(n47965) );
  XNOR U57376 ( .A(n47868), .B(n47968), .Z(n47874) );
  XNOR U57377 ( .A(n47867), .B(n47869), .Z(n47968) );
  NAND U57378 ( .A(n47969), .B(n47970), .Z(n47869) );
  OR U57379 ( .A(n47971), .B(n47972), .Z(n47970) );
  OR U57380 ( .A(n47973), .B(n47974), .Z(n47969) );
  NAND U57381 ( .A(n47975), .B(n47976), .Z(n47867) );
  OR U57382 ( .A(n47977), .B(n47978), .Z(n47976) );
  OR U57383 ( .A(n47979), .B(n47980), .Z(n47975) );
  ANDN U57384 ( .B(n47981), .A(n47982), .Z(n47868) );
  IV U57385 ( .A(n47983), .Z(n47981) );
  XNOR U57386 ( .A(n47948), .B(n47947), .Z(N61151) );
  XOR U57387 ( .A(n47967), .B(n47966), .Z(n47947) );
  XNOR U57388 ( .A(n47982), .B(n47983), .Z(n47966) );
  XNOR U57389 ( .A(n47977), .B(n47978), .Z(n47983) );
  XNOR U57390 ( .A(n47979), .B(n47980), .Z(n47978) );
  XNOR U57391 ( .A(y[1045]), .B(x[1045]), .Z(n47980) );
  XNOR U57392 ( .A(y[1046]), .B(x[1046]), .Z(n47979) );
  XNOR U57393 ( .A(y[1044]), .B(x[1044]), .Z(n47977) );
  XNOR U57394 ( .A(n47971), .B(n47972), .Z(n47982) );
  XNOR U57395 ( .A(y[1041]), .B(x[1041]), .Z(n47972) );
  XNOR U57396 ( .A(n47973), .B(n47974), .Z(n47971) );
  XNOR U57397 ( .A(y[1042]), .B(x[1042]), .Z(n47974) );
  XNOR U57398 ( .A(y[1043]), .B(x[1043]), .Z(n47973) );
  XNOR U57399 ( .A(n47964), .B(n47963), .Z(n47967) );
  XNOR U57400 ( .A(n47959), .B(n47960), .Z(n47963) );
  XNOR U57401 ( .A(y[1038]), .B(x[1038]), .Z(n47960) );
  XNOR U57402 ( .A(n47961), .B(n47962), .Z(n47959) );
  XNOR U57403 ( .A(y[1039]), .B(x[1039]), .Z(n47962) );
  XNOR U57404 ( .A(y[1040]), .B(x[1040]), .Z(n47961) );
  XNOR U57405 ( .A(n47953), .B(n47954), .Z(n47964) );
  XNOR U57406 ( .A(y[1035]), .B(x[1035]), .Z(n47954) );
  XNOR U57407 ( .A(n47955), .B(n47956), .Z(n47953) );
  XNOR U57408 ( .A(y[1036]), .B(x[1036]), .Z(n47956) );
  XNOR U57409 ( .A(y[1037]), .B(x[1037]), .Z(n47955) );
  XOR U57410 ( .A(n47929), .B(n47930), .Z(n47948) );
  XNOR U57411 ( .A(n47945), .B(n47946), .Z(n47930) );
  XNOR U57412 ( .A(n47940), .B(n47941), .Z(n47946) );
  XNOR U57413 ( .A(n47942), .B(n47943), .Z(n47941) );
  XNOR U57414 ( .A(y[1033]), .B(x[1033]), .Z(n47943) );
  XNOR U57415 ( .A(y[1034]), .B(x[1034]), .Z(n47942) );
  XNOR U57416 ( .A(y[1032]), .B(x[1032]), .Z(n47940) );
  XNOR U57417 ( .A(n47934), .B(n47935), .Z(n47945) );
  XNOR U57418 ( .A(y[1029]), .B(x[1029]), .Z(n47935) );
  XNOR U57419 ( .A(n47936), .B(n47937), .Z(n47934) );
  XNOR U57420 ( .A(y[1030]), .B(x[1030]), .Z(n47937) );
  XNOR U57421 ( .A(y[1031]), .B(x[1031]), .Z(n47936) );
  XOR U57422 ( .A(n47928), .B(n47927), .Z(n47929) );
  XNOR U57423 ( .A(n47923), .B(n47924), .Z(n47927) );
  XNOR U57424 ( .A(y[1026]), .B(x[1026]), .Z(n47924) );
  XNOR U57425 ( .A(n47925), .B(n47926), .Z(n47923) );
  XNOR U57426 ( .A(y[1027]), .B(x[1027]), .Z(n47926) );
  XNOR U57427 ( .A(y[1028]), .B(x[1028]), .Z(n47925) );
  XNOR U57428 ( .A(n47917), .B(n47918), .Z(n47928) );
  XNOR U57429 ( .A(y[1023]), .B(x[1023]), .Z(n47918) );
  XNOR U57430 ( .A(n47919), .B(n47920), .Z(n47917) );
  XNOR U57431 ( .A(y[1024]), .B(x[1024]), .Z(n47920) );
  XNOR U57432 ( .A(y[1025]), .B(x[1025]), .Z(n47919) );
  NAND U57433 ( .A(n47984), .B(n47985), .Z(N61142) );
  NANDN U57434 ( .A(n47986), .B(n47987), .Z(n47985) );
  OR U57435 ( .A(n47988), .B(n47989), .Z(n47987) );
  NAND U57436 ( .A(n47988), .B(n47989), .Z(n47984) );
  XOR U57437 ( .A(n47988), .B(n47990), .Z(N61141) );
  XNOR U57438 ( .A(n47986), .B(n47989), .Z(n47990) );
  AND U57439 ( .A(n47991), .B(n47992), .Z(n47989) );
  NANDN U57440 ( .A(n47993), .B(n47994), .Z(n47992) );
  NANDN U57441 ( .A(n47995), .B(n47996), .Z(n47994) );
  NANDN U57442 ( .A(n47996), .B(n47995), .Z(n47991) );
  NAND U57443 ( .A(n47997), .B(n47998), .Z(n47986) );
  NANDN U57444 ( .A(n47999), .B(n48000), .Z(n47998) );
  OR U57445 ( .A(n48001), .B(n48002), .Z(n48000) );
  NAND U57446 ( .A(n48002), .B(n48001), .Z(n47997) );
  AND U57447 ( .A(n48003), .B(n48004), .Z(n47988) );
  NANDN U57448 ( .A(n48005), .B(n48006), .Z(n48004) );
  NANDN U57449 ( .A(n48007), .B(n48008), .Z(n48006) );
  NANDN U57450 ( .A(n48008), .B(n48007), .Z(n48003) );
  XOR U57451 ( .A(n48002), .B(n48009), .Z(N61140) );
  XOR U57452 ( .A(n47999), .B(n48001), .Z(n48009) );
  XNOR U57453 ( .A(n47995), .B(n48010), .Z(n48001) );
  XNOR U57454 ( .A(n47993), .B(n47996), .Z(n48010) );
  NAND U57455 ( .A(n48011), .B(n48012), .Z(n47996) );
  NAND U57456 ( .A(n48013), .B(n48014), .Z(n48012) );
  OR U57457 ( .A(n48015), .B(n48016), .Z(n48013) );
  NANDN U57458 ( .A(n48017), .B(n48015), .Z(n48011) );
  IV U57459 ( .A(n48016), .Z(n48017) );
  NAND U57460 ( .A(n48018), .B(n48019), .Z(n47993) );
  NAND U57461 ( .A(n48020), .B(n48021), .Z(n48019) );
  NANDN U57462 ( .A(n48022), .B(n48023), .Z(n48020) );
  NANDN U57463 ( .A(n48023), .B(n48022), .Z(n48018) );
  AND U57464 ( .A(n48024), .B(n48025), .Z(n47995) );
  NAND U57465 ( .A(n48026), .B(n48027), .Z(n48025) );
  OR U57466 ( .A(n48028), .B(n48029), .Z(n48026) );
  NANDN U57467 ( .A(n48030), .B(n48028), .Z(n48024) );
  NAND U57468 ( .A(n48031), .B(n48032), .Z(n47999) );
  NANDN U57469 ( .A(n48033), .B(n48034), .Z(n48032) );
  OR U57470 ( .A(n48035), .B(n48036), .Z(n48034) );
  NANDN U57471 ( .A(n48037), .B(n48035), .Z(n48031) );
  IV U57472 ( .A(n48036), .Z(n48037) );
  XNOR U57473 ( .A(n48007), .B(n48038), .Z(n48002) );
  XNOR U57474 ( .A(n48005), .B(n48008), .Z(n48038) );
  NAND U57475 ( .A(n48039), .B(n48040), .Z(n48008) );
  NAND U57476 ( .A(n48041), .B(n48042), .Z(n48040) );
  OR U57477 ( .A(n48043), .B(n48044), .Z(n48041) );
  NANDN U57478 ( .A(n48045), .B(n48043), .Z(n48039) );
  IV U57479 ( .A(n48044), .Z(n48045) );
  NAND U57480 ( .A(n48046), .B(n48047), .Z(n48005) );
  NAND U57481 ( .A(n48048), .B(n48049), .Z(n48047) );
  NANDN U57482 ( .A(n48050), .B(n48051), .Z(n48048) );
  NANDN U57483 ( .A(n48051), .B(n48050), .Z(n48046) );
  AND U57484 ( .A(n48052), .B(n48053), .Z(n48007) );
  NAND U57485 ( .A(n48054), .B(n48055), .Z(n48053) );
  OR U57486 ( .A(n48056), .B(n48057), .Z(n48054) );
  NANDN U57487 ( .A(n48058), .B(n48056), .Z(n48052) );
  XNOR U57488 ( .A(n48033), .B(n48059), .Z(N61139) );
  XOR U57489 ( .A(n48035), .B(n48036), .Z(n48059) );
  XNOR U57490 ( .A(n48049), .B(n48060), .Z(n48036) );
  XOR U57491 ( .A(n48050), .B(n48051), .Z(n48060) );
  XOR U57492 ( .A(n48056), .B(n48061), .Z(n48051) );
  XOR U57493 ( .A(n48055), .B(n48058), .Z(n48061) );
  IV U57494 ( .A(n48057), .Z(n48058) );
  NAND U57495 ( .A(n48062), .B(n48063), .Z(n48057) );
  OR U57496 ( .A(n48064), .B(n48065), .Z(n48063) );
  OR U57497 ( .A(n48066), .B(n48067), .Z(n48062) );
  NAND U57498 ( .A(n48068), .B(n48069), .Z(n48055) );
  OR U57499 ( .A(n48070), .B(n48071), .Z(n48069) );
  OR U57500 ( .A(n48072), .B(n48073), .Z(n48068) );
  NOR U57501 ( .A(n48074), .B(n48075), .Z(n48056) );
  ANDN U57502 ( .B(n48076), .A(n48077), .Z(n48050) );
  XNOR U57503 ( .A(n48043), .B(n48078), .Z(n48049) );
  XNOR U57504 ( .A(n48042), .B(n48044), .Z(n48078) );
  NAND U57505 ( .A(n48079), .B(n48080), .Z(n48044) );
  OR U57506 ( .A(n48081), .B(n48082), .Z(n48080) );
  OR U57507 ( .A(n48083), .B(n48084), .Z(n48079) );
  NAND U57508 ( .A(n48085), .B(n48086), .Z(n48042) );
  OR U57509 ( .A(n48087), .B(n48088), .Z(n48086) );
  OR U57510 ( .A(n48089), .B(n48090), .Z(n48085) );
  ANDN U57511 ( .B(n48091), .A(n48092), .Z(n48043) );
  IV U57512 ( .A(n48093), .Z(n48091) );
  ANDN U57513 ( .B(n48094), .A(n48095), .Z(n48035) );
  XOR U57514 ( .A(n48021), .B(n48096), .Z(n48033) );
  XOR U57515 ( .A(n48022), .B(n48023), .Z(n48096) );
  XOR U57516 ( .A(n48028), .B(n48097), .Z(n48023) );
  XOR U57517 ( .A(n48027), .B(n48030), .Z(n48097) );
  IV U57518 ( .A(n48029), .Z(n48030) );
  NAND U57519 ( .A(n48098), .B(n48099), .Z(n48029) );
  OR U57520 ( .A(n48100), .B(n48101), .Z(n48099) );
  OR U57521 ( .A(n48102), .B(n48103), .Z(n48098) );
  NAND U57522 ( .A(n48104), .B(n48105), .Z(n48027) );
  OR U57523 ( .A(n48106), .B(n48107), .Z(n48105) );
  OR U57524 ( .A(n48108), .B(n48109), .Z(n48104) );
  NOR U57525 ( .A(n48110), .B(n48111), .Z(n48028) );
  ANDN U57526 ( .B(n48112), .A(n48113), .Z(n48022) );
  IV U57527 ( .A(n48114), .Z(n48112) );
  XNOR U57528 ( .A(n48015), .B(n48115), .Z(n48021) );
  XNOR U57529 ( .A(n48014), .B(n48016), .Z(n48115) );
  NAND U57530 ( .A(n48116), .B(n48117), .Z(n48016) );
  OR U57531 ( .A(n48118), .B(n48119), .Z(n48117) );
  OR U57532 ( .A(n48120), .B(n48121), .Z(n48116) );
  NAND U57533 ( .A(n48122), .B(n48123), .Z(n48014) );
  OR U57534 ( .A(n48124), .B(n48125), .Z(n48123) );
  OR U57535 ( .A(n48126), .B(n48127), .Z(n48122) );
  ANDN U57536 ( .B(n48128), .A(n48129), .Z(n48015) );
  IV U57537 ( .A(n48130), .Z(n48128) );
  XNOR U57538 ( .A(n48095), .B(n48094), .Z(N61138) );
  XOR U57539 ( .A(n48114), .B(n48113), .Z(n48094) );
  XNOR U57540 ( .A(n48129), .B(n48130), .Z(n48113) );
  XNOR U57541 ( .A(n48124), .B(n48125), .Z(n48130) );
  XNOR U57542 ( .A(n48126), .B(n48127), .Z(n48125) );
  XNOR U57543 ( .A(y[1021]), .B(x[1021]), .Z(n48127) );
  XNOR U57544 ( .A(y[1022]), .B(x[1022]), .Z(n48126) );
  XNOR U57545 ( .A(y[1020]), .B(x[1020]), .Z(n48124) );
  XNOR U57546 ( .A(n48118), .B(n48119), .Z(n48129) );
  XNOR U57547 ( .A(y[1017]), .B(x[1017]), .Z(n48119) );
  XNOR U57548 ( .A(n48120), .B(n48121), .Z(n48118) );
  XNOR U57549 ( .A(y[1018]), .B(x[1018]), .Z(n48121) );
  XNOR U57550 ( .A(y[1019]), .B(x[1019]), .Z(n48120) );
  XNOR U57551 ( .A(n48111), .B(n48110), .Z(n48114) );
  XNOR U57552 ( .A(n48106), .B(n48107), .Z(n48110) );
  XNOR U57553 ( .A(y[1014]), .B(x[1014]), .Z(n48107) );
  XNOR U57554 ( .A(n48108), .B(n48109), .Z(n48106) );
  XNOR U57555 ( .A(y[1015]), .B(x[1015]), .Z(n48109) );
  XNOR U57556 ( .A(y[1016]), .B(x[1016]), .Z(n48108) );
  XNOR U57557 ( .A(n48100), .B(n48101), .Z(n48111) );
  XNOR U57558 ( .A(y[1011]), .B(x[1011]), .Z(n48101) );
  XNOR U57559 ( .A(n48102), .B(n48103), .Z(n48100) );
  XNOR U57560 ( .A(y[1012]), .B(x[1012]), .Z(n48103) );
  XNOR U57561 ( .A(y[1013]), .B(x[1013]), .Z(n48102) );
  XOR U57562 ( .A(n48076), .B(n48077), .Z(n48095) );
  XNOR U57563 ( .A(n48092), .B(n48093), .Z(n48077) );
  XNOR U57564 ( .A(n48087), .B(n48088), .Z(n48093) );
  XNOR U57565 ( .A(n48089), .B(n48090), .Z(n48088) );
  XNOR U57566 ( .A(y[1009]), .B(x[1009]), .Z(n48090) );
  XNOR U57567 ( .A(y[1010]), .B(x[1010]), .Z(n48089) );
  XNOR U57568 ( .A(y[1008]), .B(x[1008]), .Z(n48087) );
  XNOR U57569 ( .A(n48081), .B(n48082), .Z(n48092) );
  XNOR U57570 ( .A(y[1005]), .B(x[1005]), .Z(n48082) );
  XNOR U57571 ( .A(n48083), .B(n48084), .Z(n48081) );
  XNOR U57572 ( .A(y[1006]), .B(x[1006]), .Z(n48084) );
  XNOR U57573 ( .A(y[1007]), .B(x[1007]), .Z(n48083) );
  XOR U57574 ( .A(n48075), .B(n48074), .Z(n48076) );
  XNOR U57575 ( .A(n48070), .B(n48071), .Z(n48074) );
  XNOR U57576 ( .A(y[1002]), .B(x[1002]), .Z(n48071) );
  XNOR U57577 ( .A(n48072), .B(n48073), .Z(n48070) );
  XNOR U57578 ( .A(y[1003]), .B(x[1003]), .Z(n48073) );
  XNOR U57579 ( .A(y[1004]), .B(x[1004]), .Z(n48072) );
  XNOR U57580 ( .A(n48064), .B(n48065), .Z(n48075) );
  XNOR U57581 ( .A(y[999]), .B(x[999]), .Z(n48065) );
  XNOR U57582 ( .A(n48066), .B(n48067), .Z(n48064) );
  XNOR U57583 ( .A(y[1000]), .B(x[1000]), .Z(n48067) );
  XNOR U57584 ( .A(y[1001]), .B(x[1001]), .Z(n48066) );
  NAND U57585 ( .A(n48131), .B(n48132), .Z(N61129) );
  NANDN U57586 ( .A(n48133), .B(n48134), .Z(n48132) );
  OR U57587 ( .A(n48135), .B(n48136), .Z(n48134) );
  NAND U57588 ( .A(n48135), .B(n48136), .Z(n48131) );
  XOR U57589 ( .A(n48135), .B(n48137), .Z(N61128) );
  XNOR U57590 ( .A(n48133), .B(n48136), .Z(n48137) );
  AND U57591 ( .A(n48138), .B(n48139), .Z(n48136) );
  NANDN U57592 ( .A(n48140), .B(n48141), .Z(n48139) );
  NANDN U57593 ( .A(n48142), .B(n48143), .Z(n48141) );
  NANDN U57594 ( .A(n48143), .B(n48142), .Z(n48138) );
  NAND U57595 ( .A(n48144), .B(n48145), .Z(n48133) );
  NANDN U57596 ( .A(n48146), .B(n48147), .Z(n48145) );
  OR U57597 ( .A(n48148), .B(n48149), .Z(n48147) );
  NAND U57598 ( .A(n48149), .B(n48148), .Z(n48144) );
  AND U57599 ( .A(n48150), .B(n48151), .Z(n48135) );
  NANDN U57600 ( .A(n48152), .B(n48153), .Z(n48151) );
  NANDN U57601 ( .A(n48154), .B(n48155), .Z(n48153) );
  NANDN U57602 ( .A(n48155), .B(n48154), .Z(n48150) );
  XOR U57603 ( .A(n48149), .B(n48156), .Z(N61127) );
  XOR U57604 ( .A(n48146), .B(n48148), .Z(n48156) );
  XNOR U57605 ( .A(n48142), .B(n48157), .Z(n48148) );
  XNOR U57606 ( .A(n48140), .B(n48143), .Z(n48157) );
  NAND U57607 ( .A(n48158), .B(n48159), .Z(n48143) );
  NAND U57608 ( .A(n48160), .B(n48161), .Z(n48159) );
  OR U57609 ( .A(n48162), .B(n48163), .Z(n48160) );
  NANDN U57610 ( .A(n48164), .B(n48162), .Z(n48158) );
  IV U57611 ( .A(n48163), .Z(n48164) );
  NAND U57612 ( .A(n48165), .B(n48166), .Z(n48140) );
  NAND U57613 ( .A(n48167), .B(n48168), .Z(n48166) );
  NANDN U57614 ( .A(n48169), .B(n48170), .Z(n48167) );
  NANDN U57615 ( .A(n48170), .B(n48169), .Z(n48165) );
  AND U57616 ( .A(n48171), .B(n48172), .Z(n48142) );
  NAND U57617 ( .A(n48173), .B(n48174), .Z(n48172) );
  OR U57618 ( .A(n48175), .B(n48176), .Z(n48173) );
  NANDN U57619 ( .A(n48177), .B(n48175), .Z(n48171) );
  NAND U57620 ( .A(n48178), .B(n48179), .Z(n48146) );
  NANDN U57621 ( .A(n48180), .B(n48181), .Z(n48179) );
  OR U57622 ( .A(n48182), .B(n48183), .Z(n48181) );
  NANDN U57623 ( .A(n48184), .B(n48182), .Z(n48178) );
  IV U57624 ( .A(n48183), .Z(n48184) );
  XNOR U57625 ( .A(n48154), .B(n48185), .Z(n48149) );
  XNOR U57626 ( .A(n48152), .B(n48155), .Z(n48185) );
  NAND U57627 ( .A(n48186), .B(n48187), .Z(n48155) );
  NAND U57628 ( .A(n48188), .B(n48189), .Z(n48187) );
  OR U57629 ( .A(n48190), .B(n48191), .Z(n48188) );
  NANDN U57630 ( .A(n48192), .B(n48190), .Z(n48186) );
  IV U57631 ( .A(n48191), .Z(n48192) );
  NAND U57632 ( .A(n48193), .B(n48194), .Z(n48152) );
  NAND U57633 ( .A(n48195), .B(n48196), .Z(n48194) );
  NANDN U57634 ( .A(n48197), .B(n48198), .Z(n48195) );
  NANDN U57635 ( .A(n48198), .B(n48197), .Z(n48193) );
  AND U57636 ( .A(n48199), .B(n48200), .Z(n48154) );
  NAND U57637 ( .A(n48201), .B(n48202), .Z(n48200) );
  OR U57638 ( .A(n48203), .B(n48204), .Z(n48201) );
  NANDN U57639 ( .A(n48205), .B(n48203), .Z(n48199) );
  XNOR U57640 ( .A(n48180), .B(n48206), .Z(N61126) );
  XOR U57641 ( .A(n48182), .B(n48183), .Z(n48206) );
  XNOR U57642 ( .A(n48196), .B(n48207), .Z(n48183) );
  XOR U57643 ( .A(n48197), .B(n48198), .Z(n48207) );
  XOR U57644 ( .A(n48203), .B(n48208), .Z(n48198) );
  XOR U57645 ( .A(n48202), .B(n48205), .Z(n48208) );
  IV U57646 ( .A(n48204), .Z(n48205) );
  NAND U57647 ( .A(n48209), .B(n48210), .Z(n48204) );
  OR U57648 ( .A(n48211), .B(n48212), .Z(n48210) );
  OR U57649 ( .A(n48213), .B(n48214), .Z(n48209) );
  NAND U57650 ( .A(n48215), .B(n48216), .Z(n48202) );
  OR U57651 ( .A(n48217), .B(n48218), .Z(n48216) );
  OR U57652 ( .A(n48219), .B(n48220), .Z(n48215) );
  NOR U57653 ( .A(n48221), .B(n48222), .Z(n48203) );
  ANDN U57654 ( .B(n48223), .A(n48224), .Z(n48197) );
  XNOR U57655 ( .A(n48190), .B(n48225), .Z(n48196) );
  XNOR U57656 ( .A(n48189), .B(n48191), .Z(n48225) );
  NAND U57657 ( .A(n48226), .B(n48227), .Z(n48191) );
  OR U57658 ( .A(n48228), .B(n48229), .Z(n48227) );
  OR U57659 ( .A(n48230), .B(n48231), .Z(n48226) );
  NAND U57660 ( .A(n48232), .B(n48233), .Z(n48189) );
  OR U57661 ( .A(n48234), .B(n48235), .Z(n48233) );
  OR U57662 ( .A(n48236), .B(n48237), .Z(n48232) );
  ANDN U57663 ( .B(n48238), .A(n48239), .Z(n48190) );
  IV U57664 ( .A(n48240), .Z(n48238) );
  ANDN U57665 ( .B(n48241), .A(n48242), .Z(n48182) );
  XOR U57666 ( .A(n48168), .B(n48243), .Z(n48180) );
  XOR U57667 ( .A(n48169), .B(n48170), .Z(n48243) );
  XOR U57668 ( .A(n48175), .B(n48244), .Z(n48170) );
  XOR U57669 ( .A(n48174), .B(n48177), .Z(n48244) );
  IV U57670 ( .A(n48176), .Z(n48177) );
  NAND U57671 ( .A(n48245), .B(n48246), .Z(n48176) );
  OR U57672 ( .A(n48247), .B(n48248), .Z(n48246) );
  OR U57673 ( .A(n48249), .B(n48250), .Z(n48245) );
  NAND U57674 ( .A(n48251), .B(n48252), .Z(n48174) );
  OR U57675 ( .A(n48253), .B(n48254), .Z(n48252) );
  OR U57676 ( .A(n48255), .B(n48256), .Z(n48251) );
  NOR U57677 ( .A(n48257), .B(n48258), .Z(n48175) );
  ANDN U57678 ( .B(n48259), .A(n48260), .Z(n48169) );
  IV U57679 ( .A(n48261), .Z(n48259) );
  XNOR U57680 ( .A(n48162), .B(n48262), .Z(n48168) );
  XNOR U57681 ( .A(n48161), .B(n48163), .Z(n48262) );
  NAND U57682 ( .A(n48263), .B(n48264), .Z(n48163) );
  OR U57683 ( .A(n48265), .B(n48266), .Z(n48264) );
  OR U57684 ( .A(n48267), .B(n48268), .Z(n48263) );
  NAND U57685 ( .A(n48269), .B(n48270), .Z(n48161) );
  OR U57686 ( .A(n48271), .B(n48272), .Z(n48270) );
  OR U57687 ( .A(n48273), .B(n48274), .Z(n48269) );
  ANDN U57688 ( .B(n48275), .A(n48276), .Z(n48162) );
  IV U57689 ( .A(n48277), .Z(n48275) );
  XNOR U57690 ( .A(n48242), .B(n48241), .Z(N61125) );
  XOR U57691 ( .A(n48261), .B(n48260), .Z(n48241) );
  XNOR U57692 ( .A(n48276), .B(n48277), .Z(n48260) );
  XNOR U57693 ( .A(n48271), .B(n48272), .Z(n48277) );
  XNOR U57694 ( .A(n48273), .B(n48274), .Z(n48272) );
  XNOR U57695 ( .A(y[997]), .B(x[997]), .Z(n48274) );
  XNOR U57696 ( .A(y[998]), .B(x[998]), .Z(n48273) );
  XNOR U57697 ( .A(y[996]), .B(x[996]), .Z(n48271) );
  XNOR U57698 ( .A(n48265), .B(n48266), .Z(n48276) );
  XNOR U57699 ( .A(y[993]), .B(x[993]), .Z(n48266) );
  XNOR U57700 ( .A(n48267), .B(n48268), .Z(n48265) );
  XNOR U57701 ( .A(y[994]), .B(x[994]), .Z(n48268) );
  XNOR U57702 ( .A(y[995]), .B(x[995]), .Z(n48267) );
  XNOR U57703 ( .A(n48258), .B(n48257), .Z(n48261) );
  XNOR U57704 ( .A(n48253), .B(n48254), .Z(n48257) );
  XNOR U57705 ( .A(y[990]), .B(x[990]), .Z(n48254) );
  XNOR U57706 ( .A(n48255), .B(n48256), .Z(n48253) );
  XNOR U57707 ( .A(y[991]), .B(x[991]), .Z(n48256) );
  XNOR U57708 ( .A(y[992]), .B(x[992]), .Z(n48255) );
  XNOR U57709 ( .A(n48247), .B(n48248), .Z(n48258) );
  XNOR U57710 ( .A(y[987]), .B(x[987]), .Z(n48248) );
  XNOR U57711 ( .A(n48249), .B(n48250), .Z(n48247) );
  XNOR U57712 ( .A(y[988]), .B(x[988]), .Z(n48250) );
  XNOR U57713 ( .A(y[989]), .B(x[989]), .Z(n48249) );
  XOR U57714 ( .A(n48223), .B(n48224), .Z(n48242) );
  XNOR U57715 ( .A(n48239), .B(n48240), .Z(n48224) );
  XNOR U57716 ( .A(n48234), .B(n48235), .Z(n48240) );
  XNOR U57717 ( .A(n48236), .B(n48237), .Z(n48235) );
  XNOR U57718 ( .A(y[985]), .B(x[985]), .Z(n48237) );
  XNOR U57719 ( .A(y[986]), .B(x[986]), .Z(n48236) );
  XNOR U57720 ( .A(y[984]), .B(x[984]), .Z(n48234) );
  XNOR U57721 ( .A(n48228), .B(n48229), .Z(n48239) );
  XNOR U57722 ( .A(y[981]), .B(x[981]), .Z(n48229) );
  XNOR U57723 ( .A(n48230), .B(n48231), .Z(n48228) );
  XNOR U57724 ( .A(y[982]), .B(x[982]), .Z(n48231) );
  XNOR U57725 ( .A(y[983]), .B(x[983]), .Z(n48230) );
  XOR U57726 ( .A(n48222), .B(n48221), .Z(n48223) );
  XNOR U57727 ( .A(n48217), .B(n48218), .Z(n48221) );
  XNOR U57728 ( .A(y[978]), .B(x[978]), .Z(n48218) );
  XNOR U57729 ( .A(n48219), .B(n48220), .Z(n48217) );
  XNOR U57730 ( .A(y[979]), .B(x[979]), .Z(n48220) );
  XNOR U57731 ( .A(y[980]), .B(x[980]), .Z(n48219) );
  XNOR U57732 ( .A(n48211), .B(n48212), .Z(n48222) );
  XNOR U57733 ( .A(y[975]), .B(x[975]), .Z(n48212) );
  XNOR U57734 ( .A(n48213), .B(n48214), .Z(n48211) );
  XNOR U57735 ( .A(y[976]), .B(x[976]), .Z(n48214) );
  XNOR U57736 ( .A(y[977]), .B(x[977]), .Z(n48213) );
  NAND U57737 ( .A(n48278), .B(n48279), .Z(N61116) );
  NANDN U57738 ( .A(n48280), .B(n48281), .Z(n48279) );
  OR U57739 ( .A(n48282), .B(n48283), .Z(n48281) );
  NAND U57740 ( .A(n48282), .B(n48283), .Z(n48278) );
  XOR U57741 ( .A(n48282), .B(n48284), .Z(N61115) );
  XNOR U57742 ( .A(n48280), .B(n48283), .Z(n48284) );
  AND U57743 ( .A(n48285), .B(n48286), .Z(n48283) );
  NANDN U57744 ( .A(n48287), .B(n48288), .Z(n48286) );
  NANDN U57745 ( .A(n48289), .B(n48290), .Z(n48288) );
  NANDN U57746 ( .A(n48290), .B(n48289), .Z(n48285) );
  NAND U57747 ( .A(n48291), .B(n48292), .Z(n48280) );
  NANDN U57748 ( .A(n48293), .B(n48294), .Z(n48292) );
  OR U57749 ( .A(n48295), .B(n48296), .Z(n48294) );
  NAND U57750 ( .A(n48296), .B(n48295), .Z(n48291) );
  AND U57751 ( .A(n48297), .B(n48298), .Z(n48282) );
  NANDN U57752 ( .A(n48299), .B(n48300), .Z(n48298) );
  NANDN U57753 ( .A(n48301), .B(n48302), .Z(n48300) );
  NANDN U57754 ( .A(n48302), .B(n48301), .Z(n48297) );
  XOR U57755 ( .A(n48296), .B(n48303), .Z(N61114) );
  XOR U57756 ( .A(n48293), .B(n48295), .Z(n48303) );
  XNOR U57757 ( .A(n48289), .B(n48304), .Z(n48295) );
  XNOR U57758 ( .A(n48287), .B(n48290), .Z(n48304) );
  NAND U57759 ( .A(n48305), .B(n48306), .Z(n48290) );
  NAND U57760 ( .A(n48307), .B(n48308), .Z(n48306) );
  OR U57761 ( .A(n48309), .B(n48310), .Z(n48307) );
  NANDN U57762 ( .A(n48311), .B(n48309), .Z(n48305) );
  IV U57763 ( .A(n48310), .Z(n48311) );
  NAND U57764 ( .A(n48312), .B(n48313), .Z(n48287) );
  NAND U57765 ( .A(n48314), .B(n48315), .Z(n48313) );
  NANDN U57766 ( .A(n48316), .B(n48317), .Z(n48314) );
  NANDN U57767 ( .A(n48317), .B(n48316), .Z(n48312) );
  AND U57768 ( .A(n48318), .B(n48319), .Z(n48289) );
  NAND U57769 ( .A(n48320), .B(n48321), .Z(n48319) );
  OR U57770 ( .A(n48322), .B(n48323), .Z(n48320) );
  NANDN U57771 ( .A(n48324), .B(n48322), .Z(n48318) );
  NAND U57772 ( .A(n48325), .B(n48326), .Z(n48293) );
  NANDN U57773 ( .A(n48327), .B(n48328), .Z(n48326) );
  OR U57774 ( .A(n48329), .B(n48330), .Z(n48328) );
  NANDN U57775 ( .A(n48331), .B(n48329), .Z(n48325) );
  IV U57776 ( .A(n48330), .Z(n48331) );
  XNOR U57777 ( .A(n48301), .B(n48332), .Z(n48296) );
  XNOR U57778 ( .A(n48299), .B(n48302), .Z(n48332) );
  NAND U57779 ( .A(n48333), .B(n48334), .Z(n48302) );
  NAND U57780 ( .A(n48335), .B(n48336), .Z(n48334) );
  OR U57781 ( .A(n48337), .B(n48338), .Z(n48335) );
  NANDN U57782 ( .A(n48339), .B(n48337), .Z(n48333) );
  IV U57783 ( .A(n48338), .Z(n48339) );
  NAND U57784 ( .A(n48340), .B(n48341), .Z(n48299) );
  NAND U57785 ( .A(n48342), .B(n48343), .Z(n48341) );
  NANDN U57786 ( .A(n48344), .B(n48345), .Z(n48342) );
  NANDN U57787 ( .A(n48345), .B(n48344), .Z(n48340) );
  AND U57788 ( .A(n48346), .B(n48347), .Z(n48301) );
  NAND U57789 ( .A(n48348), .B(n48349), .Z(n48347) );
  OR U57790 ( .A(n48350), .B(n48351), .Z(n48348) );
  NANDN U57791 ( .A(n48352), .B(n48350), .Z(n48346) );
  XNOR U57792 ( .A(n48327), .B(n48353), .Z(N61113) );
  XOR U57793 ( .A(n48329), .B(n48330), .Z(n48353) );
  XNOR U57794 ( .A(n48343), .B(n48354), .Z(n48330) );
  XOR U57795 ( .A(n48344), .B(n48345), .Z(n48354) );
  XOR U57796 ( .A(n48350), .B(n48355), .Z(n48345) );
  XOR U57797 ( .A(n48349), .B(n48352), .Z(n48355) );
  IV U57798 ( .A(n48351), .Z(n48352) );
  NAND U57799 ( .A(n48356), .B(n48357), .Z(n48351) );
  OR U57800 ( .A(n48358), .B(n48359), .Z(n48357) );
  OR U57801 ( .A(n48360), .B(n48361), .Z(n48356) );
  NAND U57802 ( .A(n48362), .B(n48363), .Z(n48349) );
  OR U57803 ( .A(n48364), .B(n48365), .Z(n48363) );
  OR U57804 ( .A(n48366), .B(n48367), .Z(n48362) );
  NOR U57805 ( .A(n48368), .B(n48369), .Z(n48350) );
  ANDN U57806 ( .B(n48370), .A(n48371), .Z(n48344) );
  XNOR U57807 ( .A(n48337), .B(n48372), .Z(n48343) );
  XNOR U57808 ( .A(n48336), .B(n48338), .Z(n48372) );
  NAND U57809 ( .A(n48373), .B(n48374), .Z(n48338) );
  OR U57810 ( .A(n48375), .B(n48376), .Z(n48374) );
  OR U57811 ( .A(n48377), .B(n48378), .Z(n48373) );
  NAND U57812 ( .A(n48379), .B(n48380), .Z(n48336) );
  OR U57813 ( .A(n48381), .B(n48382), .Z(n48380) );
  OR U57814 ( .A(n48383), .B(n48384), .Z(n48379) );
  ANDN U57815 ( .B(n48385), .A(n48386), .Z(n48337) );
  IV U57816 ( .A(n48387), .Z(n48385) );
  ANDN U57817 ( .B(n48388), .A(n48389), .Z(n48329) );
  XOR U57818 ( .A(n48315), .B(n48390), .Z(n48327) );
  XOR U57819 ( .A(n48316), .B(n48317), .Z(n48390) );
  XOR U57820 ( .A(n48322), .B(n48391), .Z(n48317) );
  XOR U57821 ( .A(n48321), .B(n48324), .Z(n48391) );
  IV U57822 ( .A(n48323), .Z(n48324) );
  NAND U57823 ( .A(n48392), .B(n48393), .Z(n48323) );
  OR U57824 ( .A(n48394), .B(n48395), .Z(n48393) );
  OR U57825 ( .A(n48396), .B(n48397), .Z(n48392) );
  NAND U57826 ( .A(n48398), .B(n48399), .Z(n48321) );
  OR U57827 ( .A(n48400), .B(n48401), .Z(n48399) );
  OR U57828 ( .A(n48402), .B(n48403), .Z(n48398) );
  NOR U57829 ( .A(n48404), .B(n48405), .Z(n48322) );
  ANDN U57830 ( .B(n48406), .A(n48407), .Z(n48316) );
  IV U57831 ( .A(n48408), .Z(n48406) );
  XNOR U57832 ( .A(n48309), .B(n48409), .Z(n48315) );
  XNOR U57833 ( .A(n48308), .B(n48310), .Z(n48409) );
  NAND U57834 ( .A(n48410), .B(n48411), .Z(n48310) );
  OR U57835 ( .A(n48412), .B(n48413), .Z(n48411) );
  OR U57836 ( .A(n48414), .B(n48415), .Z(n48410) );
  NAND U57837 ( .A(n48416), .B(n48417), .Z(n48308) );
  OR U57838 ( .A(n48418), .B(n48419), .Z(n48417) );
  OR U57839 ( .A(n48420), .B(n48421), .Z(n48416) );
  ANDN U57840 ( .B(n48422), .A(n48423), .Z(n48309) );
  IV U57841 ( .A(n48424), .Z(n48422) );
  XNOR U57842 ( .A(n48389), .B(n48388), .Z(N61112) );
  XOR U57843 ( .A(n48408), .B(n48407), .Z(n48388) );
  XNOR U57844 ( .A(n48423), .B(n48424), .Z(n48407) );
  XNOR U57845 ( .A(n48418), .B(n48419), .Z(n48424) );
  XNOR U57846 ( .A(n48420), .B(n48421), .Z(n48419) );
  XNOR U57847 ( .A(y[973]), .B(x[973]), .Z(n48421) );
  XNOR U57848 ( .A(y[974]), .B(x[974]), .Z(n48420) );
  XNOR U57849 ( .A(y[972]), .B(x[972]), .Z(n48418) );
  XNOR U57850 ( .A(n48412), .B(n48413), .Z(n48423) );
  XNOR U57851 ( .A(y[969]), .B(x[969]), .Z(n48413) );
  XNOR U57852 ( .A(n48414), .B(n48415), .Z(n48412) );
  XNOR U57853 ( .A(y[970]), .B(x[970]), .Z(n48415) );
  XNOR U57854 ( .A(y[971]), .B(x[971]), .Z(n48414) );
  XNOR U57855 ( .A(n48405), .B(n48404), .Z(n48408) );
  XNOR U57856 ( .A(n48400), .B(n48401), .Z(n48404) );
  XNOR U57857 ( .A(y[966]), .B(x[966]), .Z(n48401) );
  XNOR U57858 ( .A(n48402), .B(n48403), .Z(n48400) );
  XNOR U57859 ( .A(y[967]), .B(x[967]), .Z(n48403) );
  XNOR U57860 ( .A(y[968]), .B(x[968]), .Z(n48402) );
  XNOR U57861 ( .A(n48394), .B(n48395), .Z(n48405) );
  XNOR U57862 ( .A(y[963]), .B(x[963]), .Z(n48395) );
  XNOR U57863 ( .A(n48396), .B(n48397), .Z(n48394) );
  XNOR U57864 ( .A(y[964]), .B(x[964]), .Z(n48397) );
  XNOR U57865 ( .A(y[965]), .B(x[965]), .Z(n48396) );
  XOR U57866 ( .A(n48370), .B(n48371), .Z(n48389) );
  XNOR U57867 ( .A(n48386), .B(n48387), .Z(n48371) );
  XNOR U57868 ( .A(n48381), .B(n48382), .Z(n48387) );
  XNOR U57869 ( .A(n48383), .B(n48384), .Z(n48382) );
  XNOR U57870 ( .A(y[961]), .B(x[961]), .Z(n48384) );
  XNOR U57871 ( .A(y[962]), .B(x[962]), .Z(n48383) );
  XNOR U57872 ( .A(y[960]), .B(x[960]), .Z(n48381) );
  XNOR U57873 ( .A(n48375), .B(n48376), .Z(n48386) );
  XNOR U57874 ( .A(y[957]), .B(x[957]), .Z(n48376) );
  XNOR U57875 ( .A(n48377), .B(n48378), .Z(n48375) );
  XNOR U57876 ( .A(y[958]), .B(x[958]), .Z(n48378) );
  XNOR U57877 ( .A(y[959]), .B(x[959]), .Z(n48377) );
  XOR U57878 ( .A(n48369), .B(n48368), .Z(n48370) );
  XNOR U57879 ( .A(n48364), .B(n48365), .Z(n48368) );
  XNOR U57880 ( .A(y[954]), .B(x[954]), .Z(n48365) );
  XNOR U57881 ( .A(n48366), .B(n48367), .Z(n48364) );
  XNOR U57882 ( .A(y[955]), .B(x[955]), .Z(n48367) );
  XNOR U57883 ( .A(y[956]), .B(x[956]), .Z(n48366) );
  XNOR U57884 ( .A(n48358), .B(n48359), .Z(n48369) );
  XNOR U57885 ( .A(y[951]), .B(x[951]), .Z(n48359) );
  XNOR U57886 ( .A(n48360), .B(n48361), .Z(n48358) );
  XNOR U57887 ( .A(y[952]), .B(x[952]), .Z(n48361) );
  XNOR U57888 ( .A(y[953]), .B(x[953]), .Z(n48360) );
  NAND U57889 ( .A(n48425), .B(n48426), .Z(N61103) );
  NANDN U57890 ( .A(n48427), .B(n48428), .Z(n48426) );
  OR U57891 ( .A(n48429), .B(n48430), .Z(n48428) );
  NAND U57892 ( .A(n48429), .B(n48430), .Z(n48425) );
  XOR U57893 ( .A(n48429), .B(n48431), .Z(N61102) );
  XNOR U57894 ( .A(n48427), .B(n48430), .Z(n48431) );
  AND U57895 ( .A(n48432), .B(n48433), .Z(n48430) );
  NANDN U57896 ( .A(n48434), .B(n48435), .Z(n48433) );
  NANDN U57897 ( .A(n48436), .B(n48437), .Z(n48435) );
  NANDN U57898 ( .A(n48437), .B(n48436), .Z(n48432) );
  NAND U57899 ( .A(n48438), .B(n48439), .Z(n48427) );
  NANDN U57900 ( .A(n48440), .B(n48441), .Z(n48439) );
  OR U57901 ( .A(n48442), .B(n48443), .Z(n48441) );
  NAND U57902 ( .A(n48443), .B(n48442), .Z(n48438) );
  AND U57903 ( .A(n48444), .B(n48445), .Z(n48429) );
  NANDN U57904 ( .A(n48446), .B(n48447), .Z(n48445) );
  NANDN U57905 ( .A(n48448), .B(n48449), .Z(n48447) );
  NANDN U57906 ( .A(n48449), .B(n48448), .Z(n48444) );
  XOR U57907 ( .A(n48443), .B(n48450), .Z(N61101) );
  XOR U57908 ( .A(n48440), .B(n48442), .Z(n48450) );
  XNOR U57909 ( .A(n48436), .B(n48451), .Z(n48442) );
  XNOR U57910 ( .A(n48434), .B(n48437), .Z(n48451) );
  NAND U57911 ( .A(n48452), .B(n48453), .Z(n48437) );
  NAND U57912 ( .A(n48454), .B(n48455), .Z(n48453) );
  OR U57913 ( .A(n48456), .B(n48457), .Z(n48454) );
  NANDN U57914 ( .A(n48458), .B(n48456), .Z(n48452) );
  IV U57915 ( .A(n48457), .Z(n48458) );
  NAND U57916 ( .A(n48459), .B(n48460), .Z(n48434) );
  NAND U57917 ( .A(n48461), .B(n48462), .Z(n48460) );
  NANDN U57918 ( .A(n48463), .B(n48464), .Z(n48461) );
  NANDN U57919 ( .A(n48464), .B(n48463), .Z(n48459) );
  AND U57920 ( .A(n48465), .B(n48466), .Z(n48436) );
  NAND U57921 ( .A(n48467), .B(n48468), .Z(n48466) );
  OR U57922 ( .A(n48469), .B(n48470), .Z(n48467) );
  NANDN U57923 ( .A(n48471), .B(n48469), .Z(n48465) );
  NAND U57924 ( .A(n48472), .B(n48473), .Z(n48440) );
  NANDN U57925 ( .A(n48474), .B(n48475), .Z(n48473) );
  OR U57926 ( .A(n48476), .B(n48477), .Z(n48475) );
  NANDN U57927 ( .A(n48478), .B(n48476), .Z(n48472) );
  IV U57928 ( .A(n48477), .Z(n48478) );
  XNOR U57929 ( .A(n48448), .B(n48479), .Z(n48443) );
  XNOR U57930 ( .A(n48446), .B(n48449), .Z(n48479) );
  NAND U57931 ( .A(n48480), .B(n48481), .Z(n48449) );
  NAND U57932 ( .A(n48482), .B(n48483), .Z(n48481) );
  OR U57933 ( .A(n48484), .B(n48485), .Z(n48482) );
  NANDN U57934 ( .A(n48486), .B(n48484), .Z(n48480) );
  IV U57935 ( .A(n48485), .Z(n48486) );
  NAND U57936 ( .A(n48487), .B(n48488), .Z(n48446) );
  NAND U57937 ( .A(n48489), .B(n48490), .Z(n48488) );
  NANDN U57938 ( .A(n48491), .B(n48492), .Z(n48489) );
  NANDN U57939 ( .A(n48492), .B(n48491), .Z(n48487) );
  AND U57940 ( .A(n48493), .B(n48494), .Z(n48448) );
  NAND U57941 ( .A(n48495), .B(n48496), .Z(n48494) );
  OR U57942 ( .A(n48497), .B(n48498), .Z(n48495) );
  NANDN U57943 ( .A(n48499), .B(n48497), .Z(n48493) );
  XNOR U57944 ( .A(n48474), .B(n48500), .Z(N61100) );
  XOR U57945 ( .A(n48476), .B(n48477), .Z(n48500) );
  XNOR U57946 ( .A(n48490), .B(n48501), .Z(n48477) );
  XOR U57947 ( .A(n48491), .B(n48492), .Z(n48501) );
  XOR U57948 ( .A(n48497), .B(n48502), .Z(n48492) );
  XOR U57949 ( .A(n48496), .B(n48499), .Z(n48502) );
  IV U57950 ( .A(n48498), .Z(n48499) );
  NAND U57951 ( .A(n48503), .B(n48504), .Z(n48498) );
  OR U57952 ( .A(n48505), .B(n48506), .Z(n48504) );
  OR U57953 ( .A(n48507), .B(n48508), .Z(n48503) );
  NAND U57954 ( .A(n48509), .B(n48510), .Z(n48496) );
  OR U57955 ( .A(n48511), .B(n48512), .Z(n48510) );
  OR U57956 ( .A(n48513), .B(n48514), .Z(n48509) );
  NOR U57957 ( .A(n48515), .B(n48516), .Z(n48497) );
  ANDN U57958 ( .B(n48517), .A(n48518), .Z(n48491) );
  XNOR U57959 ( .A(n48484), .B(n48519), .Z(n48490) );
  XNOR U57960 ( .A(n48483), .B(n48485), .Z(n48519) );
  NAND U57961 ( .A(n48520), .B(n48521), .Z(n48485) );
  OR U57962 ( .A(n48522), .B(n48523), .Z(n48521) );
  OR U57963 ( .A(n48524), .B(n48525), .Z(n48520) );
  NAND U57964 ( .A(n48526), .B(n48527), .Z(n48483) );
  OR U57965 ( .A(n48528), .B(n48529), .Z(n48527) );
  OR U57966 ( .A(n48530), .B(n48531), .Z(n48526) );
  ANDN U57967 ( .B(n48532), .A(n48533), .Z(n48484) );
  IV U57968 ( .A(n48534), .Z(n48532) );
  ANDN U57969 ( .B(n48535), .A(n48536), .Z(n48476) );
  XOR U57970 ( .A(n48462), .B(n48537), .Z(n48474) );
  XOR U57971 ( .A(n48463), .B(n48464), .Z(n48537) );
  XOR U57972 ( .A(n48469), .B(n48538), .Z(n48464) );
  XOR U57973 ( .A(n48468), .B(n48471), .Z(n48538) );
  IV U57974 ( .A(n48470), .Z(n48471) );
  NAND U57975 ( .A(n48539), .B(n48540), .Z(n48470) );
  OR U57976 ( .A(n48541), .B(n48542), .Z(n48540) );
  OR U57977 ( .A(n48543), .B(n48544), .Z(n48539) );
  NAND U57978 ( .A(n48545), .B(n48546), .Z(n48468) );
  OR U57979 ( .A(n48547), .B(n48548), .Z(n48546) );
  OR U57980 ( .A(n48549), .B(n48550), .Z(n48545) );
  NOR U57981 ( .A(n48551), .B(n48552), .Z(n48469) );
  ANDN U57982 ( .B(n48553), .A(n48554), .Z(n48463) );
  IV U57983 ( .A(n48555), .Z(n48553) );
  XNOR U57984 ( .A(n48456), .B(n48556), .Z(n48462) );
  XNOR U57985 ( .A(n48455), .B(n48457), .Z(n48556) );
  NAND U57986 ( .A(n48557), .B(n48558), .Z(n48457) );
  OR U57987 ( .A(n48559), .B(n48560), .Z(n48558) );
  OR U57988 ( .A(n48561), .B(n48562), .Z(n48557) );
  NAND U57989 ( .A(n48563), .B(n48564), .Z(n48455) );
  OR U57990 ( .A(n48565), .B(n48566), .Z(n48564) );
  OR U57991 ( .A(n48567), .B(n48568), .Z(n48563) );
  ANDN U57992 ( .B(n48569), .A(n48570), .Z(n48456) );
  IV U57993 ( .A(n48571), .Z(n48569) );
  XNOR U57994 ( .A(n48536), .B(n48535), .Z(N61099) );
  XOR U57995 ( .A(n48555), .B(n48554), .Z(n48535) );
  XNOR U57996 ( .A(n48570), .B(n48571), .Z(n48554) );
  XNOR U57997 ( .A(n48565), .B(n48566), .Z(n48571) );
  XNOR U57998 ( .A(n48567), .B(n48568), .Z(n48566) );
  XNOR U57999 ( .A(y[949]), .B(x[949]), .Z(n48568) );
  XNOR U58000 ( .A(y[950]), .B(x[950]), .Z(n48567) );
  XNOR U58001 ( .A(y[948]), .B(x[948]), .Z(n48565) );
  XNOR U58002 ( .A(n48559), .B(n48560), .Z(n48570) );
  XNOR U58003 ( .A(y[945]), .B(x[945]), .Z(n48560) );
  XNOR U58004 ( .A(n48561), .B(n48562), .Z(n48559) );
  XNOR U58005 ( .A(y[946]), .B(x[946]), .Z(n48562) );
  XNOR U58006 ( .A(y[947]), .B(x[947]), .Z(n48561) );
  XNOR U58007 ( .A(n48552), .B(n48551), .Z(n48555) );
  XNOR U58008 ( .A(n48547), .B(n48548), .Z(n48551) );
  XNOR U58009 ( .A(y[942]), .B(x[942]), .Z(n48548) );
  XNOR U58010 ( .A(n48549), .B(n48550), .Z(n48547) );
  XNOR U58011 ( .A(y[943]), .B(x[943]), .Z(n48550) );
  XNOR U58012 ( .A(y[944]), .B(x[944]), .Z(n48549) );
  XNOR U58013 ( .A(n48541), .B(n48542), .Z(n48552) );
  XNOR U58014 ( .A(y[939]), .B(x[939]), .Z(n48542) );
  XNOR U58015 ( .A(n48543), .B(n48544), .Z(n48541) );
  XNOR U58016 ( .A(y[940]), .B(x[940]), .Z(n48544) );
  XNOR U58017 ( .A(y[941]), .B(x[941]), .Z(n48543) );
  XOR U58018 ( .A(n48517), .B(n48518), .Z(n48536) );
  XNOR U58019 ( .A(n48533), .B(n48534), .Z(n48518) );
  XNOR U58020 ( .A(n48528), .B(n48529), .Z(n48534) );
  XNOR U58021 ( .A(n48530), .B(n48531), .Z(n48529) );
  XNOR U58022 ( .A(y[937]), .B(x[937]), .Z(n48531) );
  XNOR U58023 ( .A(y[938]), .B(x[938]), .Z(n48530) );
  XNOR U58024 ( .A(y[936]), .B(x[936]), .Z(n48528) );
  XNOR U58025 ( .A(n48522), .B(n48523), .Z(n48533) );
  XNOR U58026 ( .A(y[933]), .B(x[933]), .Z(n48523) );
  XNOR U58027 ( .A(n48524), .B(n48525), .Z(n48522) );
  XNOR U58028 ( .A(y[934]), .B(x[934]), .Z(n48525) );
  XNOR U58029 ( .A(y[935]), .B(x[935]), .Z(n48524) );
  XOR U58030 ( .A(n48516), .B(n48515), .Z(n48517) );
  XNOR U58031 ( .A(n48511), .B(n48512), .Z(n48515) );
  XNOR U58032 ( .A(y[930]), .B(x[930]), .Z(n48512) );
  XNOR U58033 ( .A(n48513), .B(n48514), .Z(n48511) );
  XNOR U58034 ( .A(y[931]), .B(x[931]), .Z(n48514) );
  XNOR U58035 ( .A(y[932]), .B(x[932]), .Z(n48513) );
  XNOR U58036 ( .A(n48505), .B(n48506), .Z(n48516) );
  XNOR U58037 ( .A(y[927]), .B(x[927]), .Z(n48506) );
  XNOR U58038 ( .A(n48507), .B(n48508), .Z(n48505) );
  XNOR U58039 ( .A(y[928]), .B(x[928]), .Z(n48508) );
  XNOR U58040 ( .A(y[929]), .B(x[929]), .Z(n48507) );
  NAND U58041 ( .A(n48572), .B(n48573), .Z(N61090) );
  NANDN U58042 ( .A(n48574), .B(n48575), .Z(n48573) );
  OR U58043 ( .A(n48576), .B(n48577), .Z(n48575) );
  NAND U58044 ( .A(n48576), .B(n48577), .Z(n48572) );
  XOR U58045 ( .A(n48576), .B(n48578), .Z(N61089) );
  XNOR U58046 ( .A(n48574), .B(n48577), .Z(n48578) );
  AND U58047 ( .A(n48579), .B(n48580), .Z(n48577) );
  NANDN U58048 ( .A(n48581), .B(n48582), .Z(n48580) );
  NANDN U58049 ( .A(n48583), .B(n48584), .Z(n48582) );
  NANDN U58050 ( .A(n48584), .B(n48583), .Z(n48579) );
  NAND U58051 ( .A(n48585), .B(n48586), .Z(n48574) );
  NANDN U58052 ( .A(n48587), .B(n48588), .Z(n48586) );
  OR U58053 ( .A(n48589), .B(n48590), .Z(n48588) );
  NAND U58054 ( .A(n48590), .B(n48589), .Z(n48585) );
  AND U58055 ( .A(n48591), .B(n48592), .Z(n48576) );
  NANDN U58056 ( .A(n48593), .B(n48594), .Z(n48592) );
  NANDN U58057 ( .A(n48595), .B(n48596), .Z(n48594) );
  NANDN U58058 ( .A(n48596), .B(n48595), .Z(n48591) );
  XOR U58059 ( .A(n48590), .B(n48597), .Z(N61088) );
  XOR U58060 ( .A(n48587), .B(n48589), .Z(n48597) );
  XNOR U58061 ( .A(n48583), .B(n48598), .Z(n48589) );
  XNOR U58062 ( .A(n48581), .B(n48584), .Z(n48598) );
  NAND U58063 ( .A(n48599), .B(n48600), .Z(n48584) );
  NAND U58064 ( .A(n48601), .B(n48602), .Z(n48600) );
  OR U58065 ( .A(n48603), .B(n48604), .Z(n48601) );
  NANDN U58066 ( .A(n48605), .B(n48603), .Z(n48599) );
  IV U58067 ( .A(n48604), .Z(n48605) );
  NAND U58068 ( .A(n48606), .B(n48607), .Z(n48581) );
  NAND U58069 ( .A(n48608), .B(n48609), .Z(n48607) );
  NANDN U58070 ( .A(n48610), .B(n48611), .Z(n48608) );
  NANDN U58071 ( .A(n48611), .B(n48610), .Z(n48606) );
  AND U58072 ( .A(n48612), .B(n48613), .Z(n48583) );
  NAND U58073 ( .A(n48614), .B(n48615), .Z(n48613) );
  OR U58074 ( .A(n48616), .B(n48617), .Z(n48614) );
  NANDN U58075 ( .A(n48618), .B(n48616), .Z(n48612) );
  NAND U58076 ( .A(n48619), .B(n48620), .Z(n48587) );
  NANDN U58077 ( .A(n48621), .B(n48622), .Z(n48620) );
  OR U58078 ( .A(n48623), .B(n48624), .Z(n48622) );
  NANDN U58079 ( .A(n48625), .B(n48623), .Z(n48619) );
  IV U58080 ( .A(n48624), .Z(n48625) );
  XNOR U58081 ( .A(n48595), .B(n48626), .Z(n48590) );
  XNOR U58082 ( .A(n48593), .B(n48596), .Z(n48626) );
  NAND U58083 ( .A(n48627), .B(n48628), .Z(n48596) );
  NAND U58084 ( .A(n48629), .B(n48630), .Z(n48628) );
  OR U58085 ( .A(n48631), .B(n48632), .Z(n48629) );
  NANDN U58086 ( .A(n48633), .B(n48631), .Z(n48627) );
  IV U58087 ( .A(n48632), .Z(n48633) );
  NAND U58088 ( .A(n48634), .B(n48635), .Z(n48593) );
  NAND U58089 ( .A(n48636), .B(n48637), .Z(n48635) );
  NANDN U58090 ( .A(n48638), .B(n48639), .Z(n48636) );
  NANDN U58091 ( .A(n48639), .B(n48638), .Z(n48634) );
  AND U58092 ( .A(n48640), .B(n48641), .Z(n48595) );
  NAND U58093 ( .A(n48642), .B(n48643), .Z(n48641) );
  OR U58094 ( .A(n48644), .B(n48645), .Z(n48642) );
  NANDN U58095 ( .A(n48646), .B(n48644), .Z(n48640) );
  XNOR U58096 ( .A(n48621), .B(n48647), .Z(N61087) );
  XOR U58097 ( .A(n48623), .B(n48624), .Z(n48647) );
  XNOR U58098 ( .A(n48637), .B(n48648), .Z(n48624) );
  XOR U58099 ( .A(n48638), .B(n48639), .Z(n48648) );
  XOR U58100 ( .A(n48644), .B(n48649), .Z(n48639) );
  XOR U58101 ( .A(n48643), .B(n48646), .Z(n48649) );
  IV U58102 ( .A(n48645), .Z(n48646) );
  NAND U58103 ( .A(n48650), .B(n48651), .Z(n48645) );
  OR U58104 ( .A(n48652), .B(n48653), .Z(n48651) );
  OR U58105 ( .A(n48654), .B(n48655), .Z(n48650) );
  NAND U58106 ( .A(n48656), .B(n48657), .Z(n48643) );
  OR U58107 ( .A(n48658), .B(n48659), .Z(n48657) );
  OR U58108 ( .A(n48660), .B(n48661), .Z(n48656) );
  NOR U58109 ( .A(n48662), .B(n48663), .Z(n48644) );
  ANDN U58110 ( .B(n48664), .A(n48665), .Z(n48638) );
  XNOR U58111 ( .A(n48631), .B(n48666), .Z(n48637) );
  XNOR U58112 ( .A(n48630), .B(n48632), .Z(n48666) );
  NAND U58113 ( .A(n48667), .B(n48668), .Z(n48632) );
  OR U58114 ( .A(n48669), .B(n48670), .Z(n48668) );
  OR U58115 ( .A(n48671), .B(n48672), .Z(n48667) );
  NAND U58116 ( .A(n48673), .B(n48674), .Z(n48630) );
  OR U58117 ( .A(n48675), .B(n48676), .Z(n48674) );
  OR U58118 ( .A(n48677), .B(n48678), .Z(n48673) );
  ANDN U58119 ( .B(n48679), .A(n48680), .Z(n48631) );
  IV U58120 ( .A(n48681), .Z(n48679) );
  ANDN U58121 ( .B(n48682), .A(n48683), .Z(n48623) );
  XOR U58122 ( .A(n48609), .B(n48684), .Z(n48621) );
  XOR U58123 ( .A(n48610), .B(n48611), .Z(n48684) );
  XOR U58124 ( .A(n48616), .B(n48685), .Z(n48611) );
  XOR U58125 ( .A(n48615), .B(n48618), .Z(n48685) );
  IV U58126 ( .A(n48617), .Z(n48618) );
  NAND U58127 ( .A(n48686), .B(n48687), .Z(n48617) );
  OR U58128 ( .A(n48688), .B(n48689), .Z(n48687) );
  OR U58129 ( .A(n48690), .B(n48691), .Z(n48686) );
  NAND U58130 ( .A(n48692), .B(n48693), .Z(n48615) );
  OR U58131 ( .A(n48694), .B(n48695), .Z(n48693) );
  OR U58132 ( .A(n48696), .B(n48697), .Z(n48692) );
  NOR U58133 ( .A(n48698), .B(n48699), .Z(n48616) );
  ANDN U58134 ( .B(n48700), .A(n48701), .Z(n48610) );
  IV U58135 ( .A(n48702), .Z(n48700) );
  XNOR U58136 ( .A(n48603), .B(n48703), .Z(n48609) );
  XNOR U58137 ( .A(n48602), .B(n48604), .Z(n48703) );
  NAND U58138 ( .A(n48704), .B(n48705), .Z(n48604) );
  OR U58139 ( .A(n48706), .B(n48707), .Z(n48705) );
  OR U58140 ( .A(n48708), .B(n48709), .Z(n48704) );
  NAND U58141 ( .A(n48710), .B(n48711), .Z(n48602) );
  OR U58142 ( .A(n48712), .B(n48713), .Z(n48711) );
  OR U58143 ( .A(n48714), .B(n48715), .Z(n48710) );
  ANDN U58144 ( .B(n48716), .A(n48717), .Z(n48603) );
  IV U58145 ( .A(n48718), .Z(n48716) );
  XNOR U58146 ( .A(n48683), .B(n48682), .Z(N61086) );
  XOR U58147 ( .A(n48702), .B(n48701), .Z(n48682) );
  XNOR U58148 ( .A(n48717), .B(n48718), .Z(n48701) );
  XNOR U58149 ( .A(n48712), .B(n48713), .Z(n48718) );
  XNOR U58150 ( .A(n48714), .B(n48715), .Z(n48713) );
  XNOR U58151 ( .A(y[925]), .B(x[925]), .Z(n48715) );
  XNOR U58152 ( .A(y[926]), .B(x[926]), .Z(n48714) );
  XNOR U58153 ( .A(y[924]), .B(x[924]), .Z(n48712) );
  XNOR U58154 ( .A(n48706), .B(n48707), .Z(n48717) );
  XNOR U58155 ( .A(y[921]), .B(x[921]), .Z(n48707) );
  XNOR U58156 ( .A(n48708), .B(n48709), .Z(n48706) );
  XNOR U58157 ( .A(y[922]), .B(x[922]), .Z(n48709) );
  XNOR U58158 ( .A(y[923]), .B(x[923]), .Z(n48708) );
  XNOR U58159 ( .A(n48699), .B(n48698), .Z(n48702) );
  XNOR U58160 ( .A(n48694), .B(n48695), .Z(n48698) );
  XNOR U58161 ( .A(y[918]), .B(x[918]), .Z(n48695) );
  XNOR U58162 ( .A(n48696), .B(n48697), .Z(n48694) );
  XNOR U58163 ( .A(y[919]), .B(x[919]), .Z(n48697) );
  XNOR U58164 ( .A(y[920]), .B(x[920]), .Z(n48696) );
  XNOR U58165 ( .A(n48688), .B(n48689), .Z(n48699) );
  XNOR U58166 ( .A(y[915]), .B(x[915]), .Z(n48689) );
  XNOR U58167 ( .A(n48690), .B(n48691), .Z(n48688) );
  XNOR U58168 ( .A(y[916]), .B(x[916]), .Z(n48691) );
  XNOR U58169 ( .A(y[917]), .B(x[917]), .Z(n48690) );
  XOR U58170 ( .A(n48664), .B(n48665), .Z(n48683) );
  XNOR U58171 ( .A(n48680), .B(n48681), .Z(n48665) );
  XNOR U58172 ( .A(n48675), .B(n48676), .Z(n48681) );
  XNOR U58173 ( .A(n48677), .B(n48678), .Z(n48676) );
  XNOR U58174 ( .A(y[913]), .B(x[913]), .Z(n48678) );
  XNOR U58175 ( .A(y[914]), .B(x[914]), .Z(n48677) );
  XNOR U58176 ( .A(y[912]), .B(x[912]), .Z(n48675) );
  XNOR U58177 ( .A(n48669), .B(n48670), .Z(n48680) );
  XNOR U58178 ( .A(y[909]), .B(x[909]), .Z(n48670) );
  XNOR U58179 ( .A(n48671), .B(n48672), .Z(n48669) );
  XNOR U58180 ( .A(y[910]), .B(x[910]), .Z(n48672) );
  XNOR U58181 ( .A(y[911]), .B(x[911]), .Z(n48671) );
  XOR U58182 ( .A(n48663), .B(n48662), .Z(n48664) );
  XNOR U58183 ( .A(n48658), .B(n48659), .Z(n48662) );
  XNOR U58184 ( .A(y[906]), .B(x[906]), .Z(n48659) );
  XNOR U58185 ( .A(n48660), .B(n48661), .Z(n48658) );
  XNOR U58186 ( .A(y[907]), .B(x[907]), .Z(n48661) );
  XNOR U58187 ( .A(y[908]), .B(x[908]), .Z(n48660) );
  XNOR U58188 ( .A(n48652), .B(n48653), .Z(n48663) );
  XNOR U58189 ( .A(y[903]), .B(x[903]), .Z(n48653) );
  XNOR U58190 ( .A(n48654), .B(n48655), .Z(n48652) );
  XNOR U58191 ( .A(y[904]), .B(x[904]), .Z(n48655) );
  XNOR U58192 ( .A(y[905]), .B(x[905]), .Z(n48654) );
  NAND U58193 ( .A(n48719), .B(n48720), .Z(N61077) );
  NANDN U58194 ( .A(n48721), .B(n48722), .Z(n48720) );
  OR U58195 ( .A(n48723), .B(n48724), .Z(n48722) );
  NAND U58196 ( .A(n48723), .B(n48724), .Z(n48719) );
  XOR U58197 ( .A(n48723), .B(n48725), .Z(N61076) );
  XNOR U58198 ( .A(n48721), .B(n48724), .Z(n48725) );
  AND U58199 ( .A(n48726), .B(n48727), .Z(n48724) );
  NANDN U58200 ( .A(n48728), .B(n48729), .Z(n48727) );
  NANDN U58201 ( .A(n48730), .B(n48731), .Z(n48729) );
  NANDN U58202 ( .A(n48731), .B(n48730), .Z(n48726) );
  NAND U58203 ( .A(n48732), .B(n48733), .Z(n48721) );
  NANDN U58204 ( .A(n48734), .B(n48735), .Z(n48733) );
  OR U58205 ( .A(n48736), .B(n48737), .Z(n48735) );
  NAND U58206 ( .A(n48737), .B(n48736), .Z(n48732) );
  AND U58207 ( .A(n48738), .B(n48739), .Z(n48723) );
  NANDN U58208 ( .A(n48740), .B(n48741), .Z(n48739) );
  NANDN U58209 ( .A(n48742), .B(n48743), .Z(n48741) );
  NANDN U58210 ( .A(n48743), .B(n48742), .Z(n48738) );
  XOR U58211 ( .A(n48737), .B(n48744), .Z(N61075) );
  XOR U58212 ( .A(n48734), .B(n48736), .Z(n48744) );
  XNOR U58213 ( .A(n48730), .B(n48745), .Z(n48736) );
  XNOR U58214 ( .A(n48728), .B(n48731), .Z(n48745) );
  NAND U58215 ( .A(n48746), .B(n48747), .Z(n48731) );
  NAND U58216 ( .A(n48748), .B(n48749), .Z(n48747) );
  OR U58217 ( .A(n48750), .B(n48751), .Z(n48748) );
  NANDN U58218 ( .A(n48752), .B(n48750), .Z(n48746) );
  IV U58219 ( .A(n48751), .Z(n48752) );
  NAND U58220 ( .A(n48753), .B(n48754), .Z(n48728) );
  NAND U58221 ( .A(n48755), .B(n48756), .Z(n48754) );
  NANDN U58222 ( .A(n48757), .B(n48758), .Z(n48755) );
  NANDN U58223 ( .A(n48758), .B(n48757), .Z(n48753) );
  AND U58224 ( .A(n48759), .B(n48760), .Z(n48730) );
  NAND U58225 ( .A(n48761), .B(n48762), .Z(n48760) );
  OR U58226 ( .A(n48763), .B(n48764), .Z(n48761) );
  NANDN U58227 ( .A(n48765), .B(n48763), .Z(n48759) );
  NAND U58228 ( .A(n48766), .B(n48767), .Z(n48734) );
  NANDN U58229 ( .A(n48768), .B(n48769), .Z(n48767) );
  OR U58230 ( .A(n48770), .B(n48771), .Z(n48769) );
  NANDN U58231 ( .A(n48772), .B(n48770), .Z(n48766) );
  IV U58232 ( .A(n48771), .Z(n48772) );
  XNOR U58233 ( .A(n48742), .B(n48773), .Z(n48737) );
  XNOR U58234 ( .A(n48740), .B(n48743), .Z(n48773) );
  NAND U58235 ( .A(n48774), .B(n48775), .Z(n48743) );
  NAND U58236 ( .A(n48776), .B(n48777), .Z(n48775) );
  OR U58237 ( .A(n48778), .B(n48779), .Z(n48776) );
  NANDN U58238 ( .A(n48780), .B(n48778), .Z(n48774) );
  IV U58239 ( .A(n48779), .Z(n48780) );
  NAND U58240 ( .A(n48781), .B(n48782), .Z(n48740) );
  NAND U58241 ( .A(n48783), .B(n48784), .Z(n48782) );
  NANDN U58242 ( .A(n48785), .B(n48786), .Z(n48783) );
  NANDN U58243 ( .A(n48786), .B(n48785), .Z(n48781) );
  AND U58244 ( .A(n48787), .B(n48788), .Z(n48742) );
  NAND U58245 ( .A(n48789), .B(n48790), .Z(n48788) );
  OR U58246 ( .A(n48791), .B(n48792), .Z(n48789) );
  NANDN U58247 ( .A(n48793), .B(n48791), .Z(n48787) );
  XNOR U58248 ( .A(n48768), .B(n48794), .Z(N61074) );
  XOR U58249 ( .A(n48770), .B(n48771), .Z(n48794) );
  XNOR U58250 ( .A(n48784), .B(n48795), .Z(n48771) );
  XOR U58251 ( .A(n48785), .B(n48786), .Z(n48795) );
  XOR U58252 ( .A(n48791), .B(n48796), .Z(n48786) );
  XOR U58253 ( .A(n48790), .B(n48793), .Z(n48796) );
  IV U58254 ( .A(n48792), .Z(n48793) );
  NAND U58255 ( .A(n48797), .B(n48798), .Z(n48792) );
  OR U58256 ( .A(n48799), .B(n48800), .Z(n48798) );
  OR U58257 ( .A(n48801), .B(n48802), .Z(n48797) );
  NAND U58258 ( .A(n48803), .B(n48804), .Z(n48790) );
  OR U58259 ( .A(n48805), .B(n48806), .Z(n48804) );
  OR U58260 ( .A(n48807), .B(n48808), .Z(n48803) );
  NOR U58261 ( .A(n48809), .B(n48810), .Z(n48791) );
  ANDN U58262 ( .B(n48811), .A(n48812), .Z(n48785) );
  XNOR U58263 ( .A(n48778), .B(n48813), .Z(n48784) );
  XNOR U58264 ( .A(n48777), .B(n48779), .Z(n48813) );
  NAND U58265 ( .A(n48814), .B(n48815), .Z(n48779) );
  OR U58266 ( .A(n48816), .B(n48817), .Z(n48815) );
  OR U58267 ( .A(n48818), .B(n48819), .Z(n48814) );
  NAND U58268 ( .A(n48820), .B(n48821), .Z(n48777) );
  OR U58269 ( .A(n48822), .B(n48823), .Z(n48821) );
  OR U58270 ( .A(n48824), .B(n48825), .Z(n48820) );
  ANDN U58271 ( .B(n48826), .A(n48827), .Z(n48778) );
  IV U58272 ( .A(n48828), .Z(n48826) );
  ANDN U58273 ( .B(n48829), .A(n48830), .Z(n48770) );
  XOR U58274 ( .A(n48756), .B(n48831), .Z(n48768) );
  XOR U58275 ( .A(n48757), .B(n48758), .Z(n48831) );
  XOR U58276 ( .A(n48763), .B(n48832), .Z(n48758) );
  XOR U58277 ( .A(n48762), .B(n48765), .Z(n48832) );
  IV U58278 ( .A(n48764), .Z(n48765) );
  NAND U58279 ( .A(n48833), .B(n48834), .Z(n48764) );
  OR U58280 ( .A(n48835), .B(n48836), .Z(n48834) );
  OR U58281 ( .A(n48837), .B(n48838), .Z(n48833) );
  NAND U58282 ( .A(n48839), .B(n48840), .Z(n48762) );
  OR U58283 ( .A(n48841), .B(n48842), .Z(n48840) );
  OR U58284 ( .A(n48843), .B(n48844), .Z(n48839) );
  NOR U58285 ( .A(n48845), .B(n48846), .Z(n48763) );
  ANDN U58286 ( .B(n48847), .A(n48848), .Z(n48757) );
  IV U58287 ( .A(n48849), .Z(n48847) );
  XNOR U58288 ( .A(n48750), .B(n48850), .Z(n48756) );
  XNOR U58289 ( .A(n48749), .B(n48751), .Z(n48850) );
  NAND U58290 ( .A(n48851), .B(n48852), .Z(n48751) );
  OR U58291 ( .A(n48853), .B(n48854), .Z(n48852) );
  OR U58292 ( .A(n48855), .B(n48856), .Z(n48851) );
  NAND U58293 ( .A(n48857), .B(n48858), .Z(n48749) );
  OR U58294 ( .A(n48859), .B(n48860), .Z(n48858) );
  OR U58295 ( .A(n48861), .B(n48862), .Z(n48857) );
  ANDN U58296 ( .B(n48863), .A(n48864), .Z(n48750) );
  IV U58297 ( .A(n48865), .Z(n48863) );
  XNOR U58298 ( .A(n48830), .B(n48829), .Z(N61073) );
  XOR U58299 ( .A(n48849), .B(n48848), .Z(n48829) );
  XNOR U58300 ( .A(n48864), .B(n48865), .Z(n48848) );
  XNOR U58301 ( .A(n48859), .B(n48860), .Z(n48865) );
  XNOR U58302 ( .A(n48861), .B(n48862), .Z(n48860) );
  XNOR U58303 ( .A(y[901]), .B(x[901]), .Z(n48862) );
  XNOR U58304 ( .A(y[902]), .B(x[902]), .Z(n48861) );
  XNOR U58305 ( .A(y[900]), .B(x[900]), .Z(n48859) );
  XNOR U58306 ( .A(n48853), .B(n48854), .Z(n48864) );
  XNOR U58307 ( .A(y[897]), .B(x[897]), .Z(n48854) );
  XNOR U58308 ( .A(n48855), .B(n48856), .Z(n48853) );
  XNOR U58309 ( .A(y[898]), .B(x[898]), .Z(n48856) );
  XNOR U58310 ( .A(y[899]), .B(x[899]), .Z(n48855) );
  XNOR U58311 ( .A(n48846), .B(n48845), .Z(n48849) );
  XNOR U58312 ( .A(n48841), .B(n48842), .Z(n48845) );
  XNOR U58313 ( .A(y[894]), .B(x[894]), .Z(n48842) );
  XNOR U58314 ( .A(n48843), .B(n48844), .Z(n48841) );
  XNOR U58315 ( .A(y[895]), .B(x[895]), .Z(n48844) );
  XNOR U58316 ( .A(y[896]), .B(x[896]), .Z(n48843) );
  XNOR U58317 ( .A(n48835), .B(n48836), .Z(n48846) );
  XNOR U58318 ( .A(y[891]), .B(x[891]), .Z(n48836) );
  XNOR U58319 ( .A(n48837), .B(n48838), .Z(n48835) );
  XNOR U58320 ( .A(y[892]), .B(x[892]), .Z(n48838) );
  XNOR U58321 ( .A(y[893]), .B(x[893]), .Z(n48837) );
  XOR U58322 ( .A(n48811), .B(n48812), .Z(n48830) );
  XNOR U58323 ( .A(n48827), .B(n48828), .Z(n48812) );
  XNOR U58324 ( .A(n48822), .B(n48823), .Z(n48828) );
  XNOR U58325 ( .A(n48824), .B(n48825), .Z(n48823) );
  XNOR U58326 ( .A(y[889]), .B(x[889]), .Z(n48825) );
  XNOR U58327 ( .A(y[890]), .B(x[890]), .Z(n48824) );
  XNOR U58328 ( .A(y[888]), .B(x[888]), .Z(n48822) );
  XNOR U58329 ( .A(n48816), .B(n48817), .Z(n48827) );
  XNOR U58330 ( .A(y[885]), .B(x[885]), .Z(n48817) );
  XNOR U58331 ( .A(n48818), .B(n48819), .Z(n48816) );
  XNOR U58332 ( .A(y[886]), .B(x[886]), .Z(n48819) );
  XNOR U58333 ( .A(y[887]), .B(x[887]), .Z(n48818) );
  XOR U58334 ( .A(n48810), .B(n48809), .Z(n48811) );
  XNOR U58335 ( .A(n48805), .B(n48806), .Z(n48809) );
  XNOR U58336 ( .A(y[882]), .B(x[882]), .Z(n48806) );
  XNOR U58337 ( .A(n48807), .B(n48808), .Z(n48805) );
  XNOR U58338 ( .A(y[883]), .B(x[883]), .Z(n48808) );
  XNOR U58339 ( .A(y[884]), .B(x[884]), .Z(n48807) );
  XNOR U58340 ( .A(n48799), .B(n48800), .Z(n48810) );
  XNOR U58341 ( .A(y[879]), .B(x[879]), .Z(n48800) );
  XNOR U58342 ( .A(n48801), .B(n48802), .Z(n48799) );
  XNOR U58343 ( .A(y[880]), .B(x[880]), .Z(n48802) );
  XNOR U58344 ( .A(y[881]), .B(x[881]), .Z(n48801) );
  NAND U58345 ( .A(n48866), .B(n48867), .Z(N61064) );
  NANDN U58346 ( .A(n48868), .B(n48869), .Z(n48867) );
  OR U58347 ( .A(n48870), .B(n48871), .Z(n48869) );
  NAND U58348 ( .A(n48870), .B(n48871), .Z(n48866) );
  XOR U58349 ( .A(n48870), .B(n48872), .Z(N61063) );
  XNOR U58350 ( .A(n48868), .B(n48871), .Z(n48872) );
  AND U58351 ( .A(n48873), .B(n48874), .Z(n48871) );
  NANDN U58352 ( .A(n48875), .B(n48876), .Z(n48874) );
  NANDN U58353 ( .A(n48877), .B(n48878), .Z(n48876) );
  NANDN U58354 ( .A(n48878), .B(n48877), .Z(n48873) );
  NAND U58355 ( .A(n48879), .B(n48880), .Z(n48868) );
  NANDN U58356 ( .A(n48881), .B(n48882), .Z(n48880) );
  OR U58357 ( .A(n48883), .B(n48884), .Z(n48882) );
  NAND U58358 ( .A(n48884), .B(n48883), .Z(n48879) );
  AND U58359 ( .A(n48885), .B(n48886), .Z(n48870) );
  NANDN U58360 ( .A(n48887), .B(n48888), .Z(n48886) );
  NANDN U58361 ( .A(n48889), .B(n48890), .Z(n48888) );
  NANDN U58362 ( .A(n48890), .B(n48889), .Z(n48885) );
  XOR U58363 ( .A(n48884), .B(n48891), .Z(N61062) );
  XOR U58364 ( .A(n48881), .B(n48883), .Z(n48891) );
  XNOR U58365 ( .A(n48877), .B(n48892), .Z(n48883) );
  XNOR U58366 ( .A(n48875), .B(n48878), .Z(n48892) );
  NAND U58367 ( .A(n48893), .B(n48894), .Z(n48878) );
  NAND U58368 ( .A(n48895), .B(n48896), .Z(n48894) );
  OR U58369 ( .A(n48897), .B(n48898), .Z(n48895) );
  NANDN U58370 ( .A(n48899), .B(n48897), .Z(n48893) );
  IV U58371 ( .A(n48898), .Z(n48899) );
  NAND U58372 ( .A(n48900), .B(n48901), .Z(n48875) );
  NAND U58373 ( .A(n48902), .B(n48903), .Z(n48901) );
  NANDN U58374 ( .A(n48904), .B(n48905), .Z(n48902) );
  NANDN U58375 ( .A(n48905), .B(n48904), .Z(n48900) );
  AND U58376 ( .A(n48906), .B(n48907), .Z(n48877) );
  NAND U58377 ( .A(n48908), .B(n48909), .Z(n48907) );
  OR U58378 ( .A(n48910), .B(n48911), .Z(n48908) );
  NANDN U58379 ( .A(n48912), .B(n48910), .Z(n48906) );
  NAND U58380 ( .A(n48913), .B(n48914), .Z(n48881) );
  NANDN U58381 ( .A(n48915), .B(n48916), .Z(n48914) );
  OR U58382 ( .A(n48917), .B(n48918), .Z(n48916) );
  NANDN U58383 ( .A(n48919), .B(n48917), .Z(n48913) );
  IV U58384 ( .A(n48918), .Z(n48919) );
  XNOR U58385 ( .A(n48889), .B(n48920), .Z(n48884) );
  XNOR U58386 ( .A(n48887), .B(n48890), .Z(n48920) );
  NAND U58387 ( .A(n48921), .B(n48922), .Z(n48890) );
  NAND U58388 ( .A(n48923), .B(n48924), .Z(n48922) );
  OR U58389 ( .A(n48925), .B(n48926), .Z(n48923) );
  NANDN U58390 ( .A(n48927), .B(n48925), .Z(n48921) );
  IV U58391 ( .A(n48926), .Z(n48927) );
  NAND U58392 ( .A(n48928), .B(n48929), .Z(n48887) );
  NAND U58393 ( .A(n48930), .B(n48931), .Z(n48929) );
  NANDN U58394 ( .A(n48932), .B(n48933), .Z(n48930) );
  NANDN U58395 ( .A(n48933), .B(n48932), .Z(n48928) );
  AND U58396 ( .A(n48934), .B(n48935), .Z(n48889) );
  NAND U58397 ( .A(n48936), .B(n48937), .Z(n48935) );
  OR U58398 ( .A(n48938), .B(n48939), .Z(n48936) );
  NANDN U58399 ( .A(n48940), .B(n48938), .Z(n48934) );
  XNOR U58400 ( .A(n48915), .B(n48941), .Z(N61061) );
  XOR U58401 ( .A(n48917), .B(n48918), .Z(n48941) );
  XNOR U58402 ( .A(n48931), .B(n48942), .Z(n48918) );
  XOR U58403 ( .A(n48932), .B(n48933), .Z(n48942) );
  XOR U58404 ( .A(n48938), .B(n48943), .Z(n48933) );
  XOR U58405 ( .A(n48937), .B(n48940), .Z(n48943) );
  IV U58406 ( .A(n48939), .Z(n48940) );
  NAND U58407 ( .A(n48944), .B(n48945), .Z(n48939) );
  OR U58408 ( .A(n48946), .B(n48947), .Z(n48945) );
  OR U58409 ( .A(n48948), .B(n48949), .Z(n48944) );
  NAND U58410 ( .A(n48950), .B(n48951), .Z(n48937) );
  OR U58411 ( .A(n48952), .B(n48953), .Z(n48951) );
  OR U58412 ( .A(n48954), .B(n48955), .Z(n48950) );
  NOR U58413 ( .A(n48956), .B(n48957), .Z(n48938) );
  ANDN U58414 ( .B(n48958), .A(n48959), .Z(n48932) );
  XNOR U58415 ( .A(n48925), .B(n48960), .Z(n48931) );
  XNOR U58416 ( .A(n48924), .B(n48926), .Z(n48960) );
  NAND U58417 ( .A(n48961), .B(n48962), .Z(n48926) );
  OR U58418 ( .A(n48963), .B(n48964), .Z(n48962) );
  OR U58419 ( .A(n48965), .B(n48966), .Z(n48961) );
  NAND U58420 ( .A(n48967), .B(n48968), .Z(n48924) );
  OR U58421 ( .A(n48969), .B(n48970), .Z(n48968) );
  OR U58422 ( .A(n48971), .B(n48972), .Z(n48967) );
  ANDN U58423 ( .B(n48973), .A(n48974), .Z(n48925) );
  IV U58424 ( .A(n48975), .Z(n48973) );
  ANDN U58425 ( .B(n48976), .A(n48977), .Z(n48917) );
  XOR U58426 ( .A(n48903), .B(n48978), .Z(n48915) );
  XOR U58427 ( .A(n48904), .B(n48905), .Z(n48978) );
  XOR U58428 ( .A(n48910), .B(n48979), .Z(n48905) );
  XOR U58429 ( .A(n48909), .B(n48912), .Z(n48979) );
  IV U58430 ( .A(n48911), .Z(n48912) );
  NAND U58431 ( .A(n48980), .B(n48981), .Z(n48911) );
  OR U58432 ( .A(n48982), .B(n48983), .Z(n48981) );
  OR U58433 ( .A(n48984), .B(n48985), .Z(n48980) );
  NAND U58434 ( .A(n48986), .B(n48987), .Z(n48909) );
  OR U58435 ( .A(n48988), .B(n48989), .Z(n48987) );
  OR U58436 ( .A(n48990), .B(n48991), .Z(n48986) );
  NOR U58437 ( .A(n48992), .B(n48993), .Z(n48910) );
  ANDN U58438 ( .B(n48994), .A(n48995), .Z(n48904) );
  IV U58439 ( .A(n48996), .Z(n48994) );
  XNOR U58440 ( .A(n48897), .B(n48997), .Z(n48903) );
  XNOR U58441 ( .A(n48896), .B(n48898), .Z(n48997) );
  NAND U58442 ( .A(n48998), .B(n48999), .Z(n48898) );
  OR U58443 ( .A(n49000), .B(n49001), .Z(n48999) );
  OR U58444 ( .A(n49002), .B(n49003), .Z(n48998) );
  NAND U58445 ( .A(n49004), .B(n49005), .Z(n48896) );
  OR U58446 ( .A(n49006), .B(n49007), .Z(n49005) );
  OR U58447 ( .A(n49008), .B(n49009), .Z(n49004) );
  ANDN U58448 ( .B(n49010), .A(n49011), .Z(n48897) );
  IV U58449 ( .A(n49012), .Z(n49010) );
  XNOR U58450 ( .A(n48977), .B(n48976), .Z(N61060) );
  XOR U58451 ( .A(n48996), .B(n48995), .Z(n48976) );
  XNOR U58452 ( .A(n49011), .B(n49012), .Z(n48995) );
  XNOR U58453 ( .A(n49006), .B(n49007), .Z(n49012) );
  XNOR U58454 ( .A(n49008), .B(n49009), .Z(n49007) );
  XNOR U58455 ( .A(y[877]), .B(x[877]), .Z(n49009) );
  XNOR U58456 ( .A(y[878]), .B(x[878]), .Z(n49008) );
  XNOR U58457 ( .A(y[876]), .B(x[876]), .Z(n49006) );
  XNOR U58458 ( .A(n49000), .B(n49001), .Z(n49011) );
  XNOR U58459 ( .A(y[873]), .B(x[873]), .Z(n49001) );
  XNOR U58460 ( .A(n49002), .B(n49003), .Z(n49000) );
  XNOR U58461 ( .A(y[874]), .B(x[874]), .Z(n49003) );
  XNOR U58462 ( .A(y[875]), .B(x[875]), .Z(n49002) );
  XNOR U58463 ( .A(n48993), .B(n48992), .Z(n48996) );
  XNOR U58464 ( .A(n48988), .B(n48989), .Z(n48992) );
  XNOR U58465 ( .A(y[870]), .B(x[870]), .Z(n48989) );
  XNOR U58466 ( .A(n48990), .B(n48991), .Z(n48988) );
  XNOR U58467 ( .A(y[871]), .B(x[871]), .Z(n48991) );
  XNOR U58468 ( .A(y[872]), .B(x[872]), .Z(n48990) );
  XNOR U58469 ( .A(n48982), .B(n48983), .Z(n48993) );
  XNOR U58470 ( .A(y[867]), .B(x[867]), .Z(n48983) );
  XNOR U58471 ( .A(n48984), .B(n48985), .Z(n48982) );
  XNOR U58472 ( .A(y[868]), .B(x[868]), .Z(n48985) );
  XNOR U58473 ( .A(y[869]), .B(x[869]), .Z(n48984) );
  XOR U58474 ( .A(n48958), .B(n48959), .Z(n48977) );
  XNOR U58475 ( .A(n48974), .B(n48975), .Z(n48959) );
  XNOR U58476 ( .A(n48969), .B(n48970), .Z(n48975) );
  XNOR U58477 ( .A(n48971), .B(n48972), .Z(n48970) );
  XNOR U58478 ( .A(y[865]), .B(x[865]), .Z(n48972) );
  XNOR U58479 ( .A(y[866]), .B(x[866]), .Z(n48971) );
  XNOR U58480 ( .A(y[864]), .B(x[864]), .Z(n48969) );
  XNOR U58481 ( .A(n48963), .B(n48964), .Z(n48974) );
  XNOR U58482 ( .A(y[861]), .B(x[861]), .Z(n48964) );
  XNOR U58483 ( .A(n48965), .B(n48966), .Z(n48963) );
  XNOR U58484 ( .A(y[862]), .B(x[862]), .Z(n48966) );
  XNOR U58485 ( .A(y[863]), .B(x[863]), .Z(n48965) );
  XOR U58486 ( .A(n48957), .B(n48956), .Z(n48958) );
  XNOR U58487 ( .A(n48952), .B(n48953), .Z(n48956) );
  XNOR U58488 ( .A(y[858]), .B(x[858]), .Z(n48953) );
  XNOR U58489 ( .A(n48954), .B(n48955), .Z(n48952) );
  XNOR U58490 ( .A(y[859]), .B(x[859]), .Z(n48955) );
  XNOR U58491 ( .A(y[860]), .B(x[860]), .Z(n48954) );
  XNOR U58492 ( .A(n48946), .B(n48947), .Z(n48957) );
  XNOR U58493 ( .A(y[855]), .B(x[855]), .Z(n48947) );
  XNOR U58494 ( .A(n48948), .B(n48949), .Z(n48946) );
  XNOR U58495 ( .A(y[856]), .B(x[856]), .Z(n48949) );
  XNOR U58496 ( .A(y[857]), .B(x[857]), .Z(n48948) );
  NAND U58497 ( .A(n49013), .B(n49014), .Z(N61051) );
  NANDN U58498 ( .A(n49015), .B(n49016), .Z(n49014) );
  OR U58499 ( .A(n49017), .B(n49018), .Z(n49016) );
  NAND U58500 ( .A(n49017), .B(n49018), .Z(n49013) );
  XOR U58501 ( .A(n49017), .B(n49019), .Z(N61050) );
  XNOR U58502 ( .A(n49015), .B(n49018), .Z(n49019) );
  AND U58503 ( .A(n49020), .B(n49021), .Z(n49018) );
  NANDN U58504 ( .A(n49022), .B(n49023), .Z(n49021) );
  NANDN U58505 ( .A(n49024), .B(n49025), .Z(n49023) );
  NANDN U58506 ( .A(n49025), .B(n49024), .Z(n49020) );
  NAND U58507 ( .A(n49026), .B(n49027), .Z(n49015) );
  NANDN U58508 ( .A(n49028), .B(n49029), .Z(n49027) );
  OR U58509 ( .A(n49030), .B(n49031), .Z(n49029) );
  NAND U58510 ( .A(n49031), .B(n49030), .Z(n49026) );
  AND U58511 ( .A(n49032), .B(n49033), .Z(n49017) );
  NANDN U58512 ( .A(n49034), .B(n49035), .Z(n49033) );
  NANDN U58513 ( .A(n49036), .B(n49037), .Z(n49035) );
  NANDN U58514 ( .A(n49037), .B(n49036), .Z(n49032) );
  XOR U58515 ( .A(n49031), .B(n49038), .Z(N61049) );
  XOR U58516 ( .A(n49028), .B(n49030), .Z(n49038) );
  XNOR U58517 ( .A(n49024), .B(n49039), .Z(n49030) );
  XNOR U58518 ( .A(n49022), .B(n49025), .Z(n49039) );
  NAND U58519 ( .A(n49040), .B(n49041), .Z(n49025) );
  NAND U58520 ( .A(n49042), .B(n49043), .Z(n49041) );
  OR U58521 ( .A(n49044), .B(n49045), .Z(n49042) );
  NANDN U58522 ( .A(n49046), .B(n49044), .Z(n49040) );
  IV U58523 ( .A(n49045), .Z(n49046) );
  NAND U58524 ( .A(n49047), .B(n49048), .Z(n49022) );
  NAND U58525 ( .A(n49049), .B(n49050), .Z(n49048) );
  NANDN U58526 ( .A(n49051), .B(n49052), .Z(n49049) );
  NANDN U58527 ( .A(n49052), .B(n49051), .Z(n49047) );
  AND U58528 ( .A(n49053), .B(n49054), .Z(n49024) );
  NAND U58529 ( .A(n49055), .B(n49056), .Z(n49054) );
  OR U58530 ( .A(n49057), .B(n49058), .Z(n49055) );
  NANDN U58531 ( .A(n49059), .B(n49057), .Z(n49053) );
  NAND U58532 ( .A(n49060), .B(n49061), .Z(n49028) );
  NANDN U58533 ( .A(n49062), .B(n49063), .Z(n49061) );
  OR U58534 ( .A(n49064), .B(n49065), .Z(n49063) );
  NANDN U58535 ( .A(n49066), .B(n49064), .Z(n49060) );
  IV U58536 ( .A(n49065), .Z(n49066) );
  XNOR U58537 ( .A(n49036), .B(n49067), .Z(n49031) );
  XNOR U58538 ( .A(n49034), .B(n49037), .Z(n49067) );
  NAND U58539 ( .A(n49068), .B(n49069), .Z(n49037) );
  NAND U58540 ( .A(n49070), .B(n49071), .Z(n49069) );
  OR U58541 ( .A(n49072), .B(n49073), .Z(n49070) );
  NANDN U58542 ( .A(n49074), .B(n49072), .Z(n49068) );
  IV U58543 ( .A(n49073), .Z(n49074) );
  NAND U58544 ( .A(n49075), .B(n49076), .Z(n49034) );
  NAND U58545 ( .A(n49077), .B(n49078), .Z(n49076) );
  NANDN U58546 ( .A(n49079), .B(n49080), .Z(n49077) );
  NANDN U58547 ( .A(n49080), .B(n49079), .Z(n49075) );
  AND U58548 ( .A(n49081), .B(n49082), .Z(n49036) );
  NAND U58549 ( .A(n49083), .B(n49084), .Z(n49082) );
  OR U58550 ( .A(n49085), .B(n49086), .Z(n49083) );
  NANDN U58551 ( .A(n49087), .B(n49085), .Z(n49081) );
  XNOR U58552 ( .A(n49062), .B(n49088), .Z(N61048) );
  XOR U58553 ( .A(n49064), .B(n49065), .Z(n49088) );
  XNOR U58554 ( .A(n49078), .B(n49089), .Z(n49065) );
  XOR U58555 ( .A(n49079), .B(n49080), .Z(n49089) );
  XOR U58556 ( .A(n49085), .B(n49090), .Z(n49080) );
  XOR U58557 ( .A(n49084), .B(n49087), .Z(n49090) );
  IV U58558 ( .A(n49086), .Z(n49087) );
  NAND U58559 ( .A(n49091), .B(n49092), .Z(n49086) );
  OR U58560 ( .A(n49093), .B(n49094), .Z(n49092) );
  OR U58561 ( .A(n49095), .B(n49096), .Z(n49091) );
  NAND U58562 ( .A(n49097), .B(n49098), .Z(n49084) );
  OR U58563 ( .A(n49099), .B(n49100), .Z(n49098) );
  OR U58564 ( .A(n49101), .B(n49102), .Z(n49097) );
  NOR U58565 ( .A(n49103), .B(n49104), .Z(n49085) );
  ANDN U58566 ( .B(n49105), .A(n49106), .Z(n49079) );
  XNOR U58567 ( .A(n49072), .B(n49107), .Z(n49078) );
  XNOR U58568 ( .A(n49071), .B(n49073), .Z(n49107) );
  NAND U58569 ( .A(n49108), .B(n49109), .Z(n49073) );
  OR U58570 ( .A(n49110), .B(n49111), .Z(n49109) );
  OR U58571 ( .A(n49112), .B(n49113), .Z(n49108) );
  NAND U58572 ( .A(n49114), .B(n49115), .Z(n49071) );
  OR U58573 ( .A(n49116), .B(n49117), .Z(n49115) );
  OR U58574 ( .A(n49118), .B(n49119), .Z(n49114) );
  ANDN U58575 ( .B(n49120), .A(n49121), .Z(n49072) );
  IV U58576 ( .A(n49122), .Z(n49120) );
  ANDN U58577 ( .B(n49123), .A(n49124), .Z(n49064) );
  XOR U58578 ( .A(n49050), .B(n49125), .Z(n49062) );
  XOR U58579 ( .A(n49051), .B(n49052), .Z(n49125) );
  XOR U58580 ( .A(n49057), .B(n49126), .Z(n49052) );
  XOR U58581 ( .A(n49056), .B(n49059), .Z(n49126) );
  IV U58582 ( .A(n49058), .Z(n49059) );
  NAND U58583 ( .A(n49127), .B(n49128), .Z(n49058) );
  OR U58584 ( .A(n49129), .B(n49130), .Z(n49128) );
  OR U58585 ( .A(n49131), .B(n49132), .Z(n49127) );
  NAND U58586 ( .A(n49133), .B(n49134), .Z(n49056) );
  OR U58587 ( .A(n49135), .B(n49136), .Z(n49134) );
  OR U58588 ( .A(n49137), .B(n49138), .Z(n49133) );
  NOR U58589 ( .A(n49139), .B(n49140), .Z(n49057) );
  ANDN U58590 ( .B(n49141), .A(n49142), .Z(n49051) );
  IV U58591 ( .A(n49143), .Z(n49141) );
  XNOR U58592 ( .A(n49044), .B(n49144), .Z(n49050) );
  XNOR U58593 ( .A(n49043), .B(n49045), .Z(n49144) );
  NAND U58594 ( .A(n49145), .B(n49146), .Z(n49045) );
  OR U58595 ( .A(n49147), .B(n49148), .Z(n49146) );
  OR U58596 ( .A(n49149), .B(n49150), .Z(n49145) );
  NAND U58597 ( .A(n49151), .B(n49152), .Z(n49043) );
  OR U58598 ( .A(n49153), .B(n49154), .Z(n49152) );
  OR U58599 ( .A(n49155), .B(n49156), .Z(n49151) );
  ANDN U58600 ( .B(n49157), .A(n49158), .Z(n49044) );
  IV U58601 ( .A(n49159), .Z(n49157) );
  XNOR U58602 ( .A(n49124), .B(n49123), .Z(N61047) );
  XOR U58603 ( .A(n49143), .B(n49142), .Z(n49123) );
  XNOR U58604 ( .A(n49158), .B(n49159), .Z(n49142) );
  XNOR U58605 ( .A(n49153), .B(n49154), .Z(n49159) );
  XNOR U58606 ( .A(n49155), .B(n49156), .Z(n49154) );
  XNOR U58607 ( .A(y[853]), .B(x[853]), .Z(n49156) );
  XNOR U58608 ( .A(y[854]), .B(x[854]), .Z(n49155) );
  XNOR U58609 ( .A(y[852]), .B(x[852]), .Z(n49153) );
  XNOR U58610 ( .A(n49147), .B(n49148), .Z(n49158) );
  XNOR U58611 ( .A(y[849]), .B(x[849]), .Z(n49148) );
  XNOR U58612 ( .A(n49149), .B(n49150), .Z(n49147) );
  XNOR U58613 ( .A(y[850]), .B(x[850]), .Z(n49150) );
  XNOR U58614 ( .A(y[851]), .B(x[851]), .Z(n49149) );
  XNOR U58615 ( .A(n49140), .B(n49139), .Z(n49143) );
  XNOR U58616 ( .A(n49135), .B(n49136), .Z(n49139) );
  XNOR U58617 ( .A(y[846]), .B(x[846]), .Z(n49136) );
  XNOR U58618 ( .A(n49137), .B(n49138), .Z(n49135) );
  XNOR U58619 ( .A(y[847]), .B(x[847]), .Z(n49138) );
  XNOR U58620 ( .A(y[848]), .B(x[848]), .Z(n49137) );
  XNOR U58621 ( .A(n49129), .B(n49130), .Z(n49140) );
  XNOR U58622 ( .A(y[843]), .B(x[843]), .Z(n49130) );
  XNOR U58623 ( .A(n49131), .B(n49132), .Z(n49129) );
  XNOR U58624 ( .A(y[844]), .B(x[844]), .Z(n49132) );
  XNOR U58625 ( .A(y[845]), .B(x[845]), .Z(n49131) );
  XOR U58626 ( .A(n49105), .B(n49106), .Z(n49124) );
  XNOR U58627 ( .A(n49121), .B(n49122), .Z(n49106) );
  XNOR U58628 ( .A(n49116), .B(n49117), .Z(n49122) );
  XNOR U58629 ( .A(n49118), .B(n49119), .Z(n49117) );
  XNOR U58630 ( .A(y[841]), .B(x[841]), .Z(n49119) );
  XNOR U58631 ( .A(y[842]), .B(x[842]), .Z(n49118) );
  XNOR U58632 ( .A(y[840]), .B(x[840]), .Z(n49116) );
  XNOR U58633 ( .A(n49110), .B(n49111), .Z(n49121) );
  XNOR U58634 ( .A(y[837]), .B(x[837]), .Z(n49111) );
  XNOR U58635 ( .A(n49112), .B(n49113), .Z(n49110) );
  XNOR U58636 ( .A(y[838]), .B(x[838]), .Z(n49113) );
  XNOR U58637 ( .A(y[839]), .B(x[839]), .Z(n49112) );
  XOR U58638 ( .A(n49104), .B(n49103), .Z(n49105) );
  XNOR U58639 ( .A(n49099), .B(n49100), .Z(n49103) );
  XNOR U58640 ( .A(y[834]), .B(x[834]), .Z(n49100) );
  XNOR U58641 ( .A(n49101), .B(n49102), .Z(n49099) );
  XNOR U58642 ( .A(y[835]), .B(x[835]), .Z(n49102) );
  XNOR U58643 ( .A(y[836]), .B(x[836]), .Z(n49101) );
  XNOR U58644 ( .A(n49093), .B(n49094), .Z(n49104) );
  XNOR U58645 ( .A(y[831]), .B(x[831]), .Z(n49094) );
  XNOR U58646 ( .A(n49095), .B(n49096), .Z(n49093) );
  XNOR U58647 ( .A(y[832]), .B(x[832]), .Z(n49096) );
  XNOR U58648 ( .A(y[833]), .B(x[833]), .Z(n49095) );
  NAND U58649 ( .A(n49160), .B(n49161), .Z(N61038) );
  NANDN U58650 ( .A(n49162), .B(n49163), .Z(n49161) );
  OR U58651 ( .A(n49164), .B(n49165), .Z(n49163) );
  NAND U58652 ( .A(n49164), .B(n49165), .Z(n49160) );
  XOR U58653 ( .A(n49164), .B(n49166), .Z(N61037) );
  XNOR U58654 ( .A(n49162), .B(n49165), .Z(n49166) );
  AND U58655 ( .A(n49167), .B(n49168), .Z(n49165) );
  NANDN U58656 ( .A(n49169), .B(n49170), .Z(n49168) );
  NANDN U58657 ( .A(n49171), .B(n49172), .Z(n49170) );
  NANDN U58658 ( .A(n49172), .B(n49171), .Z(n49167) );
  NAND U58659 ( .A(n49173), .B(n49174), .Z(n49162) );
  NANDN U58660 ( .A(n49175), .B(n49176), .Z(n49174) );
  OR U58661 ( .A(n49177), .B(n49178), .Z(n49176) );
  NAND U58662 ( .A(n49178), .B(n49177), .Z(n49173) );
  AND U58663 ( .A(n49179), .B(n49180), .Z(n49164) );
  NANDN U58664 ( .A(n49181), .B(n49182), .Z(n49180) );
  NANDN U58665 ( .A(n49183), .B(n49184), .Z(n49182) );
  NANDN U58666 ( .A(n49184), .B(n49183), .Z(n49179) );
  XOR U58667 ( .A(n49178), .B(n49185), .Z(N61036) );
  XOR U58668 ( .A(n49175), .B(n49177), .Z(n49185) );
  XNOR U58669 ( .A(n49171), .B(n49186), .Z(n49177) );
  XNOR U58670 ( .A(n49169), .B(n49172), .Z(n49186) );
  NAND U58671 ( .A(n49187), .B(n49188), .Z(n49172) );
  NAND U58672 ( .A(n49189), .B(n49190), .Z(n49188) );
  OR U58673 ( .A(n49191), .B(n49192), .Z(n49189) );
  NANDN U58674 ( .A(n49193), .B(n49191), .Z(n49187) );
  IV U58675 ( .A(n49192), .Z(n49193) );
  NAND U58676 ( .A(n49194), .B(n49195), .Z(n49169) );
  NAND U58677 ( .A(n49196), .B(n49197), .Z(n49195) );
  NANDN U58678 ( .A(n49198), .B(n49199), .Z(n49196) );
  NANDN U58679 ( .A(n49199), .B(n49198), .Z(n49194) );
  AND U58680 ( .A(n49200), .B(n49201), .Z(n49171) );
  NAND U58681 ( .A(n49202), .B(n49203), .Z(n49201) );
  OR U58682 ( .A(n49204), .B(n49205), .Z(n49202) );
  NANDN U58683 ( .A(n49206), .B(n49204), .Z(n49200) );
  NAND U58684 ( .A(n49207), .B(n49208), .Z(n49175) );
  NANDN U58685 ( .A(n49209), .B(n49210), .Z(n49208) );
  OR U58686 ( .A(n49211), .B(n49212), .Z(n49210) );
  NANDN U58687 ( .A(n49213), .B(n49211), .Z(n49207) );
  IV U58688 ( .A(n49212), .Z(n49213) );
  XNOR U58689 ( .A(n49183), .B(n49214), .Z(n49178) );
  XNOR U58690 ( .A(n49181), .B(n49184), .Z(n49214) );
  NAND U58691 ( .A(n49215), .B(n49216), .Z(n49184) );
  NAND U58692 ( .A(n49217), .B(n49218), .Z(n49216) );
  OR U58693 ( .A(n49219), .B(n49220), .Z(n49217) );
  NANDN U58694 ( .A(n49221), .B(n49219), .Z(n49215) );
  IV U58695 ( .A(n49220), .Z(n49221) );
  NAND U58696 ( .A(n49222), .B(n49223), .Z(n49181) );
  NAND U58697 ( .A(n49224), .B(n49225), .Z(n49223) );
  NANDN U58698 ( .A(n49226), .B(n49227), .Z(n49224) );
  NANDN U58699 ( .A(n49227), .B(n49226), .Z(n49222) );
  AND U58700 ( .A(n49228), .B(n49229), .Z(n49183) );
  NAND U58701 ( .A(n49230), .B(n49231), .Z(n49229) );
  OR U58702 ( .A(n49232), .B(n49233), .Z(n49230) );
  NANDN U58703 ( .A(n49234), .B(n49232), .Z(n49228) );
  XNOR U58704 ( .A(n49209), .B(n49235), .Z(N61035) );
  XOR U58705 ( .A(n49211), .B(n49212), .Z(n49235) );
  XNOR U58706 ( .A(n49225), .B(n49236), .Z(n49212) );
  XOR U58707 ( .A(n49226), .B(n49227), .Z(n49236) );
  XOR U58708 ( .A(n49232), .B(n49237), .Z(n49227) );
  XOR U58709 ( .A(n49231), .B(n49234), .Z(n49237) );
  IV U58710 ( .A(n49233), .Z(n49234) );
  NAND U58711 ( .A(n49238), .B(n49239), .Z(n49233) );
  OR U58712 ( .A(n49240), .B(n49241), .Z(n49239) );
  OR U58713 ( .A(n49242), .B(n49243), .Z(n49238) );
  NAND U58714 ( .A(n49244), .B(n49245), .Z(n49231) );
  OR U58715 ( .A(n49246), .B(n49247), .Z(n49245) );
  OR U58716 ( .A(n49248), .B(n49249), .Z(n49244) );
  NOR U58717 ( .A(n49250), .B(n49251), .Z(n49232) );
  ANDN U58718 ( .B(n49252), .A(n49253), .Z(n49226) );
  XNOR U58719 ( .A(n49219), .B(n49254), .Z(n49225) );
  XNOR U58720 ( .A(n49218), .B(n49220), .Z(n49254) );
  NAND U58721 ( .A(n49255), .B(n49256), .Z(n49220) );
  OR U58722 ( .A(n49257), .B(n49258), .Z(n49256) );
  OR U58723 ( .A(n49259), .B(n49260), .Z(n49255) );
  NAND U58724 ( .A(n49261), .B(n49262), .Z(n49218) );
  OR U58725 ( .A(n49263), .B(n49264), .Z(n49262) );
  OR U58726 ( .A(n49265), .B(n49266), .Z(n49261) );
  ANDN U58727 ( .B(n49267), .A(n49268), .Z(n49219) );
  IV U58728 ( .A(n49269), .Z(n49267) );
  ANDN U58729 ( .B(n49270), .A(n49271), .Z(n49211) );
  XOR U58730 ( .A(n49197), .B(n49272), .Z(n49209) );
  XOR U58731 ( .A(n49198), .B(n49199), .Z(n49272) );
  XOR U58732 ( .A(n49204), .B(n49273), .Z(n49199) );
  XOR U58733 ( .A(n49203), .B(n49206), .Z(n49273) );
  IV U58734 ( .A(n49205), .Z(n49206) );
  NAND U58735 ( .A(n49274), .B(n49275), .Z(n49205) );
  OR U58736 ( .A(n49276), .B(n49277), .Z(n49275) );
  OR U58737 ( .A(n49278), .B(n49279), .Z(n49274) );
  NAND U58738 ( .A(n49280), .B(n49281), .Z(n49203) );
  OR U58739 ( .A(n49282), .B(n49283), .Z(n49281) );
  OR U58740 ( .A(n49284), .B(n49285), .Z(n49280) );
  NOR U58741 ( .A(n49286), .B(n49287), .Z(n49204) );
  ANDN U58742 ( .B(n49288), .A(n49289), .Z(n49198) );
  IV U58743 ( .A(n49290), .Z(n49288) );
  XNOR U58744 ( .A(n49191), .B(n49291), .Z(n49197) );
  XNOR U58745 ( .A(n49190), .B(n49192), .Z(n49291) );
  NAND U58746 ( .A(n49292), .B(n49293), .Z(n49192) );
  OR U58747 ( .A(n49294), .B(n49295), .Z(n49293) );
  OR U58748 ( .A(n49296), .B(n49297), .Z(n49292) );
  NAND U58749 ( .A(n49298), .B(n49299), .Z(n49190) );
  OR U58750 ( .A(n49300), .B(n49301), .Z(n49299) );
  OR U58751 ( .A(n49302), .B(n49303), .Z(n49298) );
  ANDN U58752 ( .B(n49304), .A(n49305), .Z(n49191) );
  IV U58753 ( .A(n49306), .Z(n49304) );
  XNOR U58754 ( .A(n49271), .B(n49270), .Z(N61034) );
  XOR U58755 ( .A(n49290), .B(n49289), .Z(n49270) );
  XNOR U58756 ( .A(n49305), .B(n49306), .Z(n49289) );
  XNOR U58757 ( .A(n49300), .B(n49301), .Z(n49306) );
  XNOR U58758 ( .A(n49302), .B(n49303), .Z(n49301) );
  XNOR U58759 ( .A(y[829]), .B(x[829]), .Z(n49303) );
  XNOR U58760 ( .A(y[830]), .B(x[830]), .Z(n49302) );
  XNOR U58761 ( .A(y[828]), .B(x[828]), .Z(n49300) );
  XNOR U58762 ( .A(n49294), .B(n49295), .Z(n49305) );
  XNOR U58763 ( .A(y[825]), .B(x[825]), .Z(n49295) );
  XNOR U58764 ( .A(n49296), .B(n49297), .Z(n49294) );
  XNOR U58765 ( .A(y[826]), .B(x[826]), .Z(n49297) );
  XNOR U58766 ( .A(y[827]), .B(x[827]), .Z(n49296) );
  XNOR U58767 ( .A(n49287), .B(n49286), .Z(n49290) );
  XNOR U58768 ( .A(n49282), .B(n49283), .Z(n49286) );
  XNOR U58769 ( .A(y[822]), .B(x[822]), .Z(n49283) );
  XNOR U58770 ( .A(n49284), .B(n49285), .Z(n49282) );
  XNOR U58771 ( .A(y[823]), .B(x[823]), .Z(n49285) );
  XNOR U58772 ( .A(y[824]), .B(x[824]), .Z(n49284) );
  XNOR U58773 ( .A(n49276), .B(n49277), .Z(n49287) );
  XNOR U58774 ( .A(y[819]), .B(x[819]), .Z(n49277) );
  XNOR U58775 ( .A(n49278), .B(n49279), .Z(n49276) );
  XNOR U58776 ( .A(y[820]), .B(x[820]), .Z(n49279) );
  XNOR U58777 ( .A(y[821]), .B(x[821]), .Z(n49278) );
  XOR U58778 ( .A(n49252), .B(n49253), .Z(n49271) );
  XNOR U58779 ( .A(n49268), .B(n49269), .Z(n49253) );
  XNOR U58780 ( .A(n49263), .B(n49264), .Z(n49269) );
  XNOR U58781 ( .A(n49265), .B(n49266), .Z(n49264) );
  XNOR U58782 ( .A(y[817]), .B(x[817]), .Z(n49266) );
  XNOR U58783 ( .A(y[818]), .B(x[818]), .Z(n49265) );
  XNOR U58784 ( .A(y[816]), .B(x[816]), .Z(n49263) );
  XNOR U58785 ( .A(n49257), .B(n49258), .Z(n49268) );
  XNOR U58786 ( .A(y[813]), .B(x[813]), .Z(n49258) );
  XNOR U58787 ( .A(n49259), .B(n49260), .Z(n49257) );
  XNOR U58788 ( .A(y[814]), .B(x[814]), .Z(n49260) );
  XNOR U58789 ( .A(y[815]), .B(x[815]), .Z(n49259) );
  XOR U58790 ( .A(n49251), .B(n49250), .Z(n49252) );
  XNOR U58791 ( .A(n49246), .B(n49247), .Z(n49250) );
  XNOR U58792 ( .A(y[810]), .B(x[810]), .Z(n49247) );
  XNOR U58793 ( .A(n49248), .B(n49249), .Z(n49246) );
  XNOR U58794 ( .A(y[811]), .B(x[811]), .Z(n49249) );
  XNOR U58795 ( .A(y[812]), .B(x[812]), .Z(n49248) );
  XNOR U58796 ( .A(n49240), .B(n49241), .Z(n49251) );
  XNOR U58797 ( .A(y[807]), .B(x[807]), .Z(n49241) );
  XNOR U58798 ( .A(n49242), .B(n49243), .Z(n49240) );
  XNOR U58799 ( .A(y[808]), .B(x[808]), .Z(n49243) );
  XNOR U58800 ( .A(y[809]), .B(x[809]), .Z(n49242) );
  NAND U58801 ( .A(n49307), .B(n49308), .Z(N61025) );
  NANDN U58802 ( .A(n49309), .B(n49310), .Z(n49308) );
  OR U58803 ( .A(n49311), .B(n49312), .Z(n49310) );
  NAND U58804 ( .A(n49311), .B(n49312), .Z(n49307) );
  XOR U58805 ( .A(n49311), .B(n49313), .Z(N61024) );
  XNOR U58806 ( .A(n49309), .B(n49312), .Z(n49313) );
  AND U58807 ( .A(n49314), .B(n49315), .Z(n49312) );
  NANDN U58808 ( .A(n49316), .B(n49317), .Z(n49315) );
  NANDN U58809 ( .A(n49318), .B(n49319), .Z(n49317) );
  NANDN U58810 ( .A(n49319), .B(n49318), .Z(n49314) );
  NAND U58811 ( .A(n49320), .B(n49321), .Z(n49309) );
  NANDN U58812 ( .A(n49322), .B(n49323), .Z(n49321) );
  OR U58813 ( .A(n49324), .B(n49325), .Z(n49323) );
  NAND U58814 ( .A(n49325), .B(n49324), .Z(n49320) );
  AND U58815 ( .A(n49326), .B(n49327), .Z(n49311) );
  NANDN U58816 ( .A(n49328), .B(n49329), .Z(n49327) );
  NANDN U58817 ( .A(n49330), .B(n49331), .Z(n49329) );
  NANDN U58818 ( .A(n49331), .B(n49330), .Z(n49326) );
  XOR U58819 ( .A(n49325), .B(n49332), .Z(N61023) );
  XOR U58820 ( .A(n49322), .B(n49324), .Z(n49332) );
  XNOR U58821 ( .A(n49318), .B(n49333), .Z(n49324) );
  XNOR U58822 ( .A(n49316), .B(n49319), .Z(n49333) );
  NAND U58823 ( .A(n49334), .B(n49335), .Z(n49319) );
  NAND U58824 ( .A(n49336), .B(n49337), .Z(n49335) );
  OR U58825 ( .A(n49338), .B(n49339), .Z(n49336) );
  NANDN U58826 ( .A(n49340), .B(n49338), .Z(n49334) );
  IV U58827 ( .A(n49339), .Z(n49340) );
  NAND U58828 ( .A(n49341), .B(n49342), .Z(n49316) );
  NAND U58829 ( .A(n49343), .B(n49344), .Z(n49342) );
  NANDN U58830 ( .A(n49345), .B(n49346), .Z(n49343) );
  NANDN U58831 ( .A(n49346), .B(n49345), .Z(n49341) );
  AND U58832 ( .A(n49347), .B(n49348), .Z(n49318) );
  NAND U58833 ( .A(n49349), .B(n49350), .Z(n49348) );
  OR U58834 ( .A(n49351), .B(n49352), .Z(n49349) );
  NANDN U58835 ( .A(n49353), .B(n49351), .Z(n49347) );
  NAND U58836 ( .A(n49354), .B(n49355), .Z(n49322) );
  NANDN U58837 ( .A(n49356), .B(n49357), .Z(n49355) );
  OR U58838 ( .A(n49358), .B(n49359), .Z(n49357) );
  NANDN U58839 ( .A(n49360), .B(n49358), .Z(n49354) );
  IV U58840 ( .A(n49359), .Z(n49360) );
  XNOR U58841 ( .A(n49330), .B(n49361), .Z(n49325) );
  XNOR U58842 ( .A(n49328), .B(n49331), .Z(n49361) );
  NAND U58843 ( .A(n49362), .B(n49363), .Z(n49331) );
  NAND U58844 ( .A(n49364), .B(n49365), .Z(n49363) );
  OR U58845 ( .A(n49366), .B(n49367), .Z(n49364) );
  NANDN U58846 ( .A(n49368), .B(n49366), .Z(n49362) );
  IV U58847 ( .A(n49367), .Z(n49368) );
  NAND U58848 ( .A(n49369), .B(n49370), .Z(n49328) );
  NAND U58849 ( .A(n49371), .B(n49372), .Z(n49370) );
  NANDN U58850 ( .A(n49373), .B(n49374), .Z(n49371) );
  NANDN U58851 ( .A(n49374), .B(n49373), .Z(n49369) );
  AND U58852 ( .A(n49375), .B(n49376), .Z(n49330) );
  NAND U58853 ( .A(n49377), .B(n49378), .Z(n49376) );
  OR U58854 ( .A(n49379), .B(n49380), .Z(n49377) );
  NANDN U58855 ( .A(n49381), .B(n49379), .Z(n49375) );
  XNOR U58856 ( .A(n49356), .B(n49382), .Z(N61022) );
  XOR U58857 ( .A(n49358), .B(n49359), .Z(n49382) );
  XNOR U58858 ( .A(n49372), .B(n49383), .Z(n49359) );
  XOR U58859 ( .A(n49373), .B(n49374), .Z(n49383) );
  XOR U58860 ( .A(n49379), .B(n49384), .Z(n49374) );
  XOR U58861 ( .A(n49378), .B(n49381), .Z(n49384) );
  IV U58862 ( .A(n49380), .Z(n49381) );
  NAND U58863 ( .A(n49385), .B(n49386), .Z(n49380) );
  OR U58864 ( .A(n49387), .B(n49388), .Z(n49386) );
  OR U58865 ( .A(n49389), .B(n49390), .Z(n49385) );
  NAND U58866 ( .A(n49391), .B(n49392), .Z(n49378) );
  OR U58867 ( .A(n49393), .B(n49394), .Z(n49392) );
  OR U58868 ( .A(n49395), .B(n49396), .Z(n49391) );
  NOR U58869 ( .A(n49397), .B(n49398), .Z(n49379) );
  ANDN U58870 ( .B(n49399), .A(n49400), .Z(n49373) );
  XNOR U58871 ( .A(n49366), .B(n49401), .Z(n49372) );
  XNOR U58872 ( .A(n49365), .B(n49367), .Z(n49401) );
  NAND U58873 ( .A(n49402), .B(n49403), .Z(n49367) );
  OR U58874 ( .A(n49404), .B(n49405), .Z(n49403) );
  OR U58875 ( .A(n49406), .B(n49407), .Z(n49402) );
  NAND U58876 ( .A(n49408), .B(n49409), .Z(n49365) );
  OR U58877 ( .A(n49410), .B(n49411), .Z(n49409) );
  OR U58878 ( .A(n49412), .B(n49413), .Z(n49408) );
  ANDN U58879 ( .B(n49414), .A(n49415), .Z(n49366) );
  IV U58880 ( .A(n49416), .Z(n49414) );
  ANDN U58881 ( .B(n49417), .A(n49418), .Z(n49358) );
  XOR U58882 ( .A(n49344), .B(n49419), .Z(n49356) );
  XOR U58883 ( .A(n49345), .B(n49346), .Z(n49419) );
  XOR U58884 ( .A(n49351), .B(n49420), .Z(n49346) );
  XOR U58885 ( .A(n49350), .B(n49353), .Z(n49420) );
  IV U58886 ( .A(n49352), .Z(n49353) );
  NAND U58887 ( .A(n49421), .B(n49422), .Z(n49352) );
  OR U58888 ( .A(n49423), .B(n49424), .Z(n49422) );
  OR U58889 ( .A(n49425), .B(n49426), .Z(n49421) );
  NAND U58890 ( .A(n49427), .B(n49428), .Z(n49350) );
  OR U58891 ( .A(n49429), .B(n49430), .Z(n49428) );
  OR U58892 ( .A(n49431), .B(n49432), .Z(n49427) );
  NOR U58893 ( .A(n49433), .B(n49434), .Z(n49351) );
  ANDN U58894 ( .B(n49435), .A(n49436), .Z(n49345) );
  IV U58895 ( .A(n49437), .Z(n49435) );
  XNOR U58896 ( .A(n49338), .B(n49438), .Z(n49344) );
  XNOR U58897 ( .A(n49337), .B(n49339), .Z(n49438) );
  NAND U58898 ( .A(n49439), .B(n49440), .Z(n49339) );
  OR U58899 ( .A(n49441), .B(n49442), .Z(n49440) );
  OR U58900 ( .A(n49443), .B(n49444), .Z(n49439) );
  NAND U58901 ( .A(n49445), .B(n49446), .Z(n49337) );
  OR U58902 ( .A(n49447), .B(n49448), .Z(n49446) );
  OR U58903 ( .A(n49449), .B(n49450), .Z(n49445) );
  ANDN U58904 ( .B(n49451), .A(n49452), .Z(n49338) );
  IV U58905 ( .A(n49453), .Z(n49451) );
  XNOR U58906 ( .A(n49418), .B(n49417), .Z(N61021) );
  XOR U58907 ( .A(n49437), .B(n49436), .Z(n49417) );
  XNOR U58908 ( .A(n49452), .B(n49453), .Z(n49436) );
  XNOR U58909 ( .A(n49447), .B(n49448), .Z(n49453) );
  XNOR U58910 ( .A(n49449), .B(n49450), .Z(n49448) );
  XNOR U58911 ( .A(y[805]), .B(x[805]), .Z(n49450) );
  XNOR U58912 ( .A(y[806]), .B(x[806]), .Z(n49449) );
  XNOR U58913 ( .A(y[804]), .B(x[804]), .Z(n49447) );
  XNOR U58914 ( .A(n49441), .B(n49442), .Z(n49452) );
  XNOR U58915 ( .A(y[801]), .B(x[801]), .Z(n49442) );
  XNOR U58916 ( .A(n49443), .B(n49444), .Z(n49441) );
  XNOR U58917 ( .A(y[802]), .B(x[802]), .Z(n49444) );
  XNOR U58918 ( .A(y[803]), .B(x[803]), .Z(n49443) );
  XNOR U58919 ( .A(n49434), .B(n49433), .Z(n49437) );
  XNOR U58920 ( .A(n49429), .B(n49430), .Z(n49433) );
  XNOR U58921 ( .A(y[798]), .B(x[798]), .Z(n49430) );
  XNOR U58922 ( .A(n49431), .B(n49432), .Z(n49429) );
  XNOR U58923 ( .A(y[799]), .B(x[799]), .Z(n49432) );
  XNOR U58924 ( .A(y[800]), .B(x[800]), .Z(n49431) );
  XNOR U58925 ( .A(n49423), .B(n49424), .Z(n49434) );
  XNOR U58926 ( .A(y[795]), .B(x[795]), .Z(n49424) );
  XNOR U58927 ( .A(n49425), .B(n49426), .Z(n49423) );
  XNOR U58928 ( .A(y[796]), .B(x[796]), .Z(n49426) );
  XNOR U58929 ( .A(y[797]), .B(x[797]), .Z(n49425) );
  XOR U58930 ( .A(n49399), .B(n49400), .Z(n49418) );
  XNOR U58931 ( .A(n49415), .B(n49416), .Z(n49400) );
  XNOR U58932 ( .A(n49410), .B(n49411), .Z(n49416) );
  XNOR U58933 ( .A(n49412), .B(n49413), .Z(n49411) );
  XNOR U58934 ( .A(y[793]), .B(x[793]), .Z(n49413) );
  XNOR U58935 ( .A(y[794]), .B(x[794]), .Z(n49412) );
  XNOR U58936 ( .A(y[792]), .B(x[792]), .Z(n49410) );
  XNOR U58937 ( .A(n49404), .B(n49405), .Z(n49415) );
  XNOR U58938 ( .A(y[789]), .B(x[789]), .Z(n49405) );
  XNOR U58939 ( .A(n49406), .B(n49407), .Z(n49404) );
  XNOR U58940 ( .A(y[790]), .B(x[790]), .Z(n49407) );
  XNOR U58941 ( .A(y[791]), .B(x[791]), .Z(n49406) );
  XOR U58942 ( .A(n49398), .B(n49397), .Z(n49399) );
  XNOR U58943 ( .A(n49393), .B(n49394), .Z(n49397) );
  XNOR U58944 ( .A(y[786]), .B(x[786]), .Z(n49394) );
  XNOR U58945 ( .A(n49395), .B(n49396), .Z(n49393) );
  XNOR U58946 ( .A(y[787]), .B(x[787]), .Z(n49396) );
  XNOR U58947 ( .A(y[788]), .B(x[788]), .Z(n49395) );
  XNOR U58948 ( .A(n49387), .B(n49388), .Z(n49398) );
  XNOR U58949 ( .A(y[783]), .B(x[783]), .Z(n49388) );
  XNOR U58950 ( .A(n49389), .B(n49390), .Z(n49387) );
  XNOR U58951 ( .A(y[784]), .B(x[784]), .Z(n49390) );
  XNOR U58952 ( .A(y[785]), .B(x[785]), .Z(n49389) );
  NAND U58953 ( .A(n49454), .B(n49455), .Z(N61012) );
  NANDN U58954 ( .A(n49456), .B(n49457), .Z(n49455) );
  OR U58955 ( .A(n49458), .B(n49459), .Z(n49457) );
  NAND U58956 ( .A(n49458), .B(n49459), .Z(n49454) );
  XOR U58957 ( .A(n49458), .B(n49460), .Z(N61011) );
  XNOR U58958 ( .A(n49456), .B(n49459), .Z(n49460) );
  AND U58959 ( .A(n49461), .B(n49462), .Z(n49459) );
  NANDN U58960 ( .A(n49463), .B(n49464), .Z(n49462) );
  NANDN U58961 ( .A(n49465), .B(n49466), .Z(n49464) );
  NANDN U58962 ( .A(n49466), .B(n49465), .Z(n49461) );
  NAND U58963 ( .A(n49467), .B(n49468), .Z(n49456) );
  NANDN U58964 ( .A(n49469), .B(n49470), .Z(n49468) );
  OR U58965 ( .A(n49471), .B(n49472), .Z(n49470) );
  NAND U58966 ( .A(n49472), .B(n49471), .Z(n49467) );
  AND U58967 ( .A(n49473), .B(n49474), .Z(n49458) );
  NANDN U58968 ( .A(n49475), .B(n49476), .Z(n49474) );
  NANDN U58969 ( .A(n49477), .B(n49478), .Z(n49476) );
  NANDN U58970 ( .A(n49478), .B(n49477), .Z(n49473) );
  XOR U58971 ( .A(n49472), .B(n49479), .Z(N61010) );
  XOR U58972 ( .A(n49469), .B(n49471), .Z(n49479) );
  XNOR U58973 ( .A(n49465), .B(n49480), .Z(n49471) );
  XNOR U58974 ( .A(n49463), .B(n49466), .Z(n49480) );
  NAND U58975 ( .A(n49481), .B(n49482), .Z(n49466) );
  NAND U58976 ( .A(n49483), .B(n49484), .Z(n49482) );
  OR U58977 ( .A(n49485), .B(n49486), .Z(n49483) );
  NANDN U58978 ( .A(n49487), .B(n49485), .Z(n49481) );
  IV U58979 ( .A(n49486), .Z(n49487) );
  NAND U58980 ( .A(n49488), .B(n49489), .Z(n49463) );
  NAND U58981 ( .A(n49490), .B(n49491), .Z(n49489) );
  NANDN U58982 ( .A(n49492), .B(n49493), .Z(n49490) );
  NANDN U58983 ( .A(n49493), .B(n49492), .Z(n49488) );
  AND U58984 ( .A(n49494), .B(n49495), .Z(n49465) );
  NAND U58985 ( .A(n49496), .B(n49497), .Z(n49495) );
  OR U58986 ( .A(n49498), .B(n49499), .Z(n49496) );
  NANDN U58987 ( .A(n49500), .B(n49498), .Z(n49494) );
  NAND U58988 ( .A(n49501), .B(n49502), .Z(n49469) );
  NANDN U58989 ( .A(n49503), .B(n49504), .Z(n49502) );
  OR U58990 ( .A(n49505), .B(n49506), .Z(n49504) );
  NANDN U58991 ( .A(n49507), .B(n49505), .Z(n49501) );
  IV U58992 ( .A(n49506), .Z(n49507) );
  XNOR U58993 ( .A(n49477), .B(n49508), .Z(n49472) );
  XNOR U58994 ( .A(n49475), .B(n49478), .Z(n49508) );
  NAND U58995 ( .A(n49509), .B(n49510), .Z(n49478) );
  NAND U58996 ( .A(n49511), .B(n49512), .Z(n49510) );
  OR U58997 ( .A(n49513), .B(n49514), .Z(n49511) );
  NANDN U58998 ( .A(n49515), .B(n49513), .Z(n49509) );
  IV U58999 ( .A(n49514), .Z(n49515) );
  NAND U59000 ( .A(n49516), .B(n49517), .Z(n49475) );
  NAND U59001 ( .A(n49518), .B(n49519), .Z(n49517) );
  NANDN U59002 ( .A(n49520), .B(n49521), .Z(n49518) );
  NANDN U59003 ( .A(n49521), .B(n49520), .Z(n49516) );
  AND U59004 ( .A(n49522), .B(n49523), .Z(n49477) );
  NAND U59005 ( .A(n49524), .B(n49525), .Z(n49523) );
  OR U59006 ( .A(n49526), .B(n49527), .Z(n49524) );
  NANDN U59007 ( .A(n49528), .B(n49526), .Z(n49522) );
  XNOR U59008 ( .A(n49503), .B(n49529), .Z(N61009) );
  XOR U59009 ( .A(n49505), .B(n49506), .Z(n49529) );
  XNOR U59010 ( .A(n49519), .B(n49530), .Z(n49506) );
  XOR U59011 ( .A(n49520), .B(n49521), .Z(n49530) );
  XOR U59012 ( .A(n49526), .B(n49531), .Z(n49521) );
  XOR U59013 ( .A(n49525), .B(n49528), .Z(n49531) );
  IV U59014 ( .A(n49527), .Z(n49528) );
  NAND U59015 ( .A(n49532), .B(n49533), .Z(n49527) );
  OR U59016 ( .A(n49534), .B(n49535), .Z(n49533) );
  OR U59017 ( .A(n49536), .B(n49537), .Z(n49532) );
  NAND U59018 ( .A(n49538), .B(n49539), .Z(n49525) );
  OR U59019 ( .A(n49540), .B(n49541), .Z(n49539) );
  OR U59020 ( .A(n49542), .B(n49543), .Z(n49538) );
  NOR U59021 ( .A(n49544), .B(n49545), .Z(n49526) );
  ANDN U59022 ( .B(n49546), .A(n49547), .Z(n49520) );
  XNOR U59023 ( .A(n49513), .B(n49548), .Z(n49519) );
  XNOR U59024 ( .A(n49512), .B(n49514), .Z(n49548) );
  NAND U59025 ( .A(n49549), .B(n49550), .Z(n49514) );
  OR U59026 ( .A(n49551), .B(n49552), .Z(n49550) );
  OR U59027 ( .A(n49553), .B(n49554), .Z(n49549) );
  NAND U59028 ( .A(n49555), .B(n49556), .Z(n49512) );
  OR U59029 ( .A(n49557), .B(n49558), .Z(n49556) );
  OR U59030 ( .A(n49559), .B(n49560), .Z(n49555) );
  ANDN U59031 ( .B(n49561), .A(n49562), .Z(n49513) );
  IV U59032 ( .A(n49563), .Z(n49561) );
  ANDN U59033 ( .B(n49564), .A(n49565), .Z(n49505) );
  XOR U59034 ( .A(n49491), .B(n49566), .Z(n49503) );
  XOR U59035 ( .A(n49492), .B(n49493), .Z(n49566) );
  XOR U59036 ( .A(n49498), .B(n49567), .Z(n49493) );
  XOR U59037 ( .A(n49497), .B(n49500), .Z(n49567) );
  IV U59038 ( .A(n49499), .Z(n49500) );
  NAND U59039 ( .A(n49568), .B(n49569), .Z(n49499) );
  OR U59040 ( .A(n49570), .B(n49571), .Z(n49569) );
  OR U59041 ( .A(n49572), .B(n49573), .Z(n49568) );
  NAND U59042 ( .A(n49574), .B(n49575), .Z(n49497) );
  OR U59043 ( .A(n49576), .B(n49577), .Z(n49575) );
  OR U59044 ( .A(n49578), .B(n49579), .Z(n49574) );
  NOR U59045 ( .A(n49580), .B(n49581), .Z(n49498) );
  ANDN U59046 ( .B(n49582), .A(n49583), .Z(n49492) );
  IV U59047 ( .A(n49584), .Z(n49582) );
  XNOR U59048 ( .A(n49485), .B(n49585), .Z(n49491) );
  XNOR U59049 ( .A(n49484), .B(n49486), .Z(n49585) );
  NAND U59050 ( .A(n49586), .B(n49587), .Z(n49486) );
  OR U59051 ( .A(n49588), .B(n49589), .Z(n49587) );
  OR U59052 ( .A(n49590), .B(n49591), .Z(n49586) );
  NAND U59053 ( .A(n49592), .B(n49593), .Z(n49484) );
  OR U59054 ( .A(n49594), .B(n49595), .Z(n49593) );
  OR U59055 ( .A(n49596), .B(n49597), .Z(n49592) );
  ANDN U59056 ( .B(n49598), .A(n49599), .Z(n49485) );
  IV U59057 ( .A(n49600), .Z(n49598) );
  XNOR U59058 ( .A(n49565), .B(n49564), .Z(N61008) );
  XOR U59059 ( .A(n49584), .B(n49583), .Z(n49564) );
  XNOR U59060 ( .A(n49599), .B(n49600), .Z(n49583) );
  XNOR U59061 ( .A(n49594), .B(n49595), .Z(n49600) );
  XNOR U59062 ( .A(n49596), .B(n49597), .Z(n49595) );
  XNOR U59063 ( .A(y[781]), .B(x[781]), .Z(n49597) );
  XNOR U59064 ( .A(y[782]), .B(x[782]), .Z(n49596) );
  XNOR U59065 ( .A(y[780]), .B(x[780]), .Z(n49594) );
  XNOR U59066 ( .A(n49588), .B(n49589), .Z(n49599) );
  XNOR U59067 ( .A(y[777]), .B(x[777]), .Z(n49589) );
  XNOR U59068 ( .A(n49590), .B(n49591), .Z(n49588) );
  XNOR U59069 ( .A(y[778]), .B(x[778]), .Z(n49591) );
  XNOR U59070 ( .A(y[779]), .B(x[779]), .Z(n49590) );
  XNOR U59071 ( .A(n49581), .B(n49580), .Z(n49584) );
  XNOR U59072 ( .A(n49576), .B(n49577), .Z(n49580) );
  XNOR U59073 ( .A(y[774]), .B(x[774]), .Z(n49577) );
  XNOR U59074 ( .A(n49578), .B(n49579), .Z(n49576) );
  XNOR U59075 ( .A(y[775]), .B(x[775]), .Z(n49579) );
  XNOR U59076 ( .A(y[776]), .B(x[776]), .Z(n49578) );
  XNOR U59077 ( .A(n49570), .B(n49571), .Z(n49581) );
  XNOR U59078 ( .A(y[771]), .B(x[771]), .Z(n49571) );
  XNOR U59079 ( .A(n49572), .B(n49573), .Z(n49570) );
  XNOR U59080 ( .A(y[772]), .B(x[772]), .Z(n49573) );
  XNOR U59081 ( .A(y[773]), .B(x[773]), .Z(n49572) );
  XOR U59082 ( .A(n49546), .B(n49547), .Z(n49565) );
  XNOR U59083 ( .A(n49562), .B(n49563), .Z(n49547) );
  XNOR U59084 ( .A(n49557), .B(n49558), .Z(n49563) );
  XNOR U59085 ( .A(n49559), .B(n49560), .Z(n49558) );
  XNOR U59086 ( .A(y[769]), .B(x[769]), .Z(n49560) );
  XNOR U59087 ( .A(y[770]), .B(x[770]), .Z(n49559) );
  XNOR U59088 ( .A(y[768]), .B(x[768]), .Z(n49557) );
  XNOR U59089 ( .A(n49551), .B(n49552), .Z(n49562) );
  XNOR U59090 ( .A(y[765]), .B(x[765]), .Z(n49552) );
  XNOR U59091 ( .A(n49553), .B(n49554), .Z(n49551) );
  XNOR U59092 ( .A(y[766]), .B(x[766]), .Z(n49554) );
  XNOR U59093 ( .A(y[767]), .B(x[767]), .Z(n49553) );
  XOR U59094 ( .A(n49545), .B(n49544), .Z(n49546) );
  XNOR U59095 ( .A(n49540), .B(n49541), .Z(n49544) );
  XNOR U59096 ( .A(y[762]), .B(x[762]), .Z(n49541) );
  XNOR U59097 ( .A(n49542), .B(n49543), .Z(n49540) );
  XNOR U59098 ( .A(y[763]), .B(x[763]), .Z(n49543) );
  XNOR U59099 ( .A(y[764]), .B(x[764]), .Z(n49542) );
  XNOR U59100 ( .A(n49534), .B(n49535), .Z(n49545) );
  XNOR U59101 ( .A(y[759]), .B(x[759]), .Z(n49535) );
  XNOR U59102 ( .A(n49536), .B(n49537), .Z(n49534) );
  XNOR U59103 ( .A(y[760]), .B(x[760]), .Z(n49537) );
  XNOR U59104 ( .A(y[761]), .B(x[761]), .Z(n49536) );
  NAND U59105 ( .A(n49601), .B(n49602), .Z(N60999) );
  NANDN U59106 ( .A(n49603), .B(n49604), .Z(n49602) );
  OR U59107 ( .A(n49605), .B(n49606), .Z(n49604) );
  NAND U59108 ( .A(n49605), .B(n49606), .Z(n49601) );
  XOR U59109 ( .A(n49605), .B(n49607), .Z(N60998) );
  XNOR U59110 ( .A(n49603), .B(n49606), .Z(n49607) );
  AND U59111 ( .A(n49608), .B(n49609), .Z(n49606) );
  NANDN U59112 ( .A(n49610), .B(n49611), .Z(n49609) );
  NANDN U59113 ( .A(n49612), .B(n49613), .Z(n49611) );
  NANDN U59114 ( .A(n49613), .B(n49612), .Z(n49608) );
  NAND U59115 ( .A(n49614), .B(n49615), .Z(n49603) );
  NANDN U59116 ( .A(n49616), .B(n49617), .Z(n49615) );
  OR U59117 ( .A(n49618), .B(n49619), .Z(n49617) );
  NAND U59118 ( .A(n49619), .B(n49618), .Z(n49614) );
  AND U59119 ( .A(n49620), .B(n49621), .Z(n49605) );
  NANDN U59120 ( .A(n49622), .B(n49623), .Z(n49621) );
  NANDN U59121 ( .A(n49624), .B(n49625), .Z(n49623) );
  NANDN U59122 ( .A(n49625), .B(n49624), .Z(n49620) );
  XOR U59123 ( .A(n49619), .B(n49626), .Z(N60997) );
  XOR U59124 ( .A(n49616), .B(n49618), .Z(n49626) );
  XNOR U59125 ( .A(n49612), .B(n49627), .Z(n49618) );
  XNOR U59126 ( .A(n49610), .B(n49613), .Z(n49627) );
  NAND U59127 ( .A(n49628), .B(n49629), .Z(n49613) );
  NAND U59128 ( .A(n49630), .B(n49631), .Z(n49629) );
  OR U59129 ( .A(n49632), .B(n49633), .Z(n49630) );
  NANDN U59130 ( .A(n49634), .B(n49632), .Z(n49628) );
  IV U59131 ( .A(n49633), .Z(n49634) );
  NAND U59132 ( .A(n49635), .B(n49636), .Z(n49610) );
  NAND U59133 ( .A(n49637), .B(n49638), .Z(n49636) );
  NANDN U59134 ( .A(n49639), .B(n49640), .Z(n49637) );
  NANDN U59135 ( .A(n49640), .B(n49639), .Z(n49635) );
  AND U59136 ( .A(n49641), .B(n49642), .Z(n49612) );
  NAND U59137 ( .A(n49643), .B(n49644), .Z(n49642) );
  OR U59138 ( .A(n49645), .B(n49646), .Z(n49643) );
  NANDN U59139 ( .A(n49647), .B(n49645), .Z(n49641) );
  NAND U59140 ( .A(n49648), .B(n49649), .Z(n49616) );
  NANDN U59141 ( .A(n49650), .B(n49651), .Z(n49649) );
  OR U59142 ( .A(n49652), .B(n49653), .Z(n49651) );
  NANDN U59143 ( .A(n49654), .B(n49652), .Z(n49648) );
  IV U59144 ( .A(n49653), .Z(n49654) );
  XNOR U59145 ( .A(n49624), .B(n49655), .Z(n49619) );
  XNOR U59146 ( .A(n49622), .B(n49625), .Z(n49655) );
  NAND U59147 ( .A(n49656), .B(n49657), .Z(n49625) );
  NAND U59148 ( .A(n49658), .B(n49659), .Z(n49657) );
  OR U59149 ( .A(n49660), .B(n49661), .Z(n49658) );
  NANDN U59150 ( .A(n49662), .B(n49660), .Z(n49656) );
  IV U59151 ( .A(n49661), .Z(n49662) );
  NAND U59152 ( .A(n49663), .B(n49664), .Z(n49622) );
  NAND U59153 ( .A(n49665), .B(n49666), .Z(n49664) );
  NANDN U59154 ( .A(n49667), .B(n49668), .Z(n49665) );
  NANDN U59155 ( .A(n49668), .B(n49667), .Z(n49663) );
  AND U59156 ( .A(n49669), .B(n49670), .Z(n49624) );
  NAND U59157 ( .A(n49671), .B(n49672), .Z(n49670) );
  OR U59158 ( .A(n49673), .B(n49674), .Z(n49671) );
  NANDN U59159 ( .A(n49675), .B(n49673), .Z(n49669) );
  XNOR U59160 ( .A(n49650), .B(n49676), .Z(N60996) );
  XOR U59161 ( .A(n49652), .B(n49653), .Z(n49676) );
  XNOR U59162 ( .A(n49666), .B(n49677), .Z(n49653) );
  XOR U59163 ( .A(n49667), .B(n49668), .Z(n49677) );
  XOR U59164 ( .A(n49673), .B(n49678), .Z(n49668) );
  XOR U59165 ( .A(n49672), .B(n49675), .Z(n49678) );
  IV U59166 ( .A(n49674), .Z(n49675) );
  NAND U59167 ( .A(n49679), .B(n49680), .Z(n49674) );
  OR U59168 ( .A(n49681), .B(n49682), .Z(n49680) );
  OR U59169 ( .A(n49683), .B(n49684), .Z(n49679) );
  NAND U59170 ( .A(n49685), .B(n49686), .Z(n49672) );
  OR U59171 ( .A(n49687), .B(n49688), .Z(n49686) );
  OR U59172 ( .A(n49689), .B(n49690), .Z(n49685) );
  NOR U59173 ( .A(n49691), .B(n49692), .Z(n49673) );
  ANDN U59174 ( .B(n49693), .A(n49694), .Z(n49667) );
  XNOR U59175 ( .A(n49660), .B(n49695), .Z(n49666) );
  XNOR U59176 ( .A(n49659), .B(n49661), .Z(n49695) );
  NAND U59177 ( .A(n49696), .B(n49697), .Z(n49661) );
  OR U59178 ( .A(n49698), .B(n49699), .Z(n49697) );
  OR U59179 ( .A(n49700), .B(n49701), .Z(n49696) );
  NAND U59180 ( .A(n49702), .B(n49703), .Z(n49659) );
  OR U59181 ( .A(n49704), .B(n49705), .Z(n49703) );
  OR U59182 ( .A(n49706), .B(n49707), .Z(n49702) );
  ANDN U59183 ( .B(n49708), .A(n49709), .Z(n49660) );
  IV U59184 ( .A(n49710), .Z(n49708) );
  ANDN U59185 ( .B(n49711), .A(n49712), .Z(n49652) );
  XOR U59186 ( .A(n49638), .B(n49713), .Z(n49650) );
  XOR U59187 ( .A(n49639), .B(n49640), .Z(n49713) );
  XOR U59188 ( .A(n49645), .B(n49714), .Z(n49640) );
  XOR U59189 ( .A(n49644), .B(n49647), .Z(n49714) );
  IV U59190 ( .A(n49646), .Z(n49647) );
  NAND U59191 ( .A(n49715), .B(n49716), .Z(n49646) );
  OR U59192 ( .A(n49717), .B(n49718), .Z(n49716) );
  OR U59193 ( .A(n49719), .B(n49720), .Z(n49715) );
  NAND U59194 ( .A(n49721), .B(n49722), .Z(n49644) );
  OR U59195 ( .A(n49723), .B(n49724), .Z(n49722) );
  OR U59196 ( .A(n49725), .B(n49726), .Z(n49721) );
  NOR U59197 ( .A(n49727), .B(n49728), .Z(n49645) );
  ANDN U59198 ( .B(n49729), .A(n49730), .Z(n49639) );
  IV U59199 ( .A(n49731), .Z(n49729) );
  XNOR U59200 ( .A(n49632), .B(n49732), .Z(n49638) );
  XNOR U59201 ( .A(n49631), .B(n49633), .Z(n49732) );
  NAND U59202 ( .A(n49733), .B(n49734), .Z(n49633) );
  OR U59203 ( .A(n49735), .B(n49736), .Z(n49734) );
  OR U59204 ( .A(n49737), .B(n49738), .Z(n49733) );
  NAND U59205 ( .A(n49739), .B(n49740), .Z(n49631) );
  OR U59206 ( .A(n49741), .B(n49742), .Z(n49740) );
  OR U59207 ( .A(n49743), .B(n49744), .Z(n49739) );
  ANDN U59208 ( .B(n49745), .A(n49746), .Z(n49632) );
  IV U59209 ( .A(n49747), .Z(n49745) );
  XNOR U59210 ( .A(n49712), .B(n49711), .Z(N60995) );
  XOR U59211 ( .A(n49731), .B(n49730), .Z(n49711) );
  XNOR U59212 ( .A(n49746), .B(n49747), .Z(n49730) );
  XNOR U59213 ( .A(n49741), .B(n49742), .Z(n49747) );
  XNOR U59214 ( .A(n49743), .B(n49744), .Z(n49742) );
  XNOR U59215 ( .A(y[757]), .B(x[757]), .Z(n49744) );
  XNOR U59216 ( .A(y[758]), .B(x[758]), .Z(n49743) );
  XNOR U59217 ( .A(y[756]), .B(x[756]), .Z(n49741) );
  XNOR U59218 ( .A(n49735), .B(n49736), .Z(n49746) );
  XNOR U59219 ( .A(y[753]), .B(x[753]), .Z(n49736) );
  XNOR U59220 ( .A(n49737), .B(n49738), .Z(n49735) );
  XNOR U59221 ( .A(y[754]), .B(x[754]), .Z(n49738) );
  XNOR U59222 ( .A(y[755]), .B(x[755]), .Z(n49737) );
  XNOR U59223 ( .A(n49728), .B(n49727), .Z(n49731) );
  XNOR U59224 ( .A(n49723), .B(n49724), .Z(n49727) );
  XNOR U59225 ( .A(y[750]), .B(x[750]), .Z(n49724) );
  XNOR U59226 ( .A(n49725), .B(n49726), .Z(n49723) );
  XNOR U59227 ( .A(y[751]), .B(x[751]), .Z(n49726) );
  XNOR U59228 ( .A(y[752]), .B(x[752]), .Z(n49725) );
  XNOR U59229 ( .A(n49717), .B(n49718), .Z(n49728) );
  XNOR U59230 ( .A(y[747]), .B(x[747]), .Z(n49718) );
  XNOR U59231 ( .A(n49719), .B(n49720), .Z(n49717) );
  XNOR U59232 ( .A(y[748]), .B(x[748]), .Z(n49720) );
  XNOR U59233 ( .A(y[749]), .B(x[749]), .Z(n49719) );
  XOR U59234 ( .A(n49693), .B(n49694), .Z(n49712) );
  XNOR U59235 ( .A(n49709), .B(n49710), .Z(n49694) );
  XNOR U59236 ( .A(n49704), .B(n49705), .Z(n49710) );
  XNOR U59237 ( .A(n49706), .B(n49707), .Z(n49705) );
  XNOR U59238 ( .A(y[745]), .B(x[745]), .Z(n49707) );
  XNOR U59239 ( .A(y[746]), .B(x[746]), .Z(n49706) );
  XNOR U59240 ( .A(y[744]), .B(x[744]), .Z(n49704) );
  XNOR U59241 ( .A(n49698), .B(n49699), .Z(n49709) );
  XNOR U59242 ( .A(y[741]), .B(x[741]), .Z(n49699) );
  XNOR U59243 ( .A(n49700), .B(n49701), .Z(n49698) );
  XNOR U59244 ( .A(y[742]), .B(x[742]), .Z(n49701) );
  XNOR U59245 ( .A(y[743]), .B(x[743]), .Z(n49700) );
  XOR U59246 ( .A(n49692), .B(n49691), .Z(n49693) );
  XNOR U59247 ( .A(n49687), .B(n49688), .Z(n49691) );
  XNOR U59248 ( .A(y[738]), .B(x[738]), .Z(n49688) );
  XNOR U59249 ( .A(n49689), .B(n49690), .Z(n49687) );
  XNOR U59250 ( .A(y[739]), .B(x[739]), .Z(n49690) );
  XNOR U59251 ( .A(y[740]), .B(x[740]), .Z(n49689) );
  XNOR U59252 ( .A(n49681), .B(n49682), .Z(n49692) );
  XNOR U59253 ( .A(y[735]), .B(x[735]), .Z(n49682) );
  XNOR U59254 ( .A(n49683), .B(n49684), .Z(n49681) );
  XNOR U59255 ( .A(y[736]), .B(x[736]), .Z(n49684) );
  XNOR U59256 ( .A(y[737]), .B(x[737]), .Z(n49683) );
  NAND U59257 ( .A(n49748), .B(n49749), .Z(N60986) );
  NANDN U59258 ( .A(n49750), .B(n49751), .Z(n49749) );
  OR U59259 ( .A(n49752), .B(n49753), .Z(n49751) );
  NAND U59260 ( .A(n49752), .B(n49753), .Z(n49748) );
  XOR U59261 ( .A(n49752), .B(n49754), .Z(N60985) );
  XNOR U59262 ( .A(n49750), .B(n49753), .Z(n49754) );
  AND U59263 ( .A(n49755), .B(n49756), .Z(n49753) );
  NANDN U59264 ( .A(n49757), .B(n49758), .Z(n49756) );
  NANDN U59265 ( .A(n49759), .B(n49760), .Z(n49758) );
  NANDN U59266 ( .A(n49760), .B(n49759), .Z(n49755) );
  NAND U59267 ( .A(n49761), .B(n49762), .Z(n49750) );
  NANDN U59268 ( .A(n49763), .B(n49764), .Z(n49762) );
  OR U59269 ( .A(n49765), .B(n49766), .Z(n49764) );
  NAND U59270 ( .A(n49766), .B(n49765), .Z(n49761) );
  AND U59271 ( .A(n49767), .B(n49768), .Z(n49752) );
  NANDN U59272 ( .A(n49769), .B(n49770), .Z(n49768) );
  NANDN U59273 ( .A(n49771), .B(n49772), .Z(n49770) );
  NANDN U59274 ( .A(n49772), .B(n49771), .Z(n49767) );
  XOR U59275 ( .A(n49766), .B(n49773), .Z(N60984) );
  XOR U59276 ( .A(n49763), .B(n49765), .Z(n49773) );
  XNOR U59277 ( .A(n49759), .B(n49774), .Z(n49765) );
  XNOR U59278 ( .A(n49757), .B(n49760), .Z(n49774) );
  NAND U59279 ( .A(n49775), .B(n49776), .Z(n49760) );
  NAND U59280 ( .A(n49777), .B(n49778), .Z(n49776) );
  OR U59281 ( .A(n49779), .B(n49780), .Z(n49777) );
  NANDN U59282 ( .A(n49781), .B(n49779), .Z(n49775) );
  IV U59283 ( .A(n49780), .Z(n49781) );
  NAND U59284 ( .A(n49782), .B(n49783), .Z(n49757) );
  NAND U59285 ( .A(n49784), .B(n49785), .Z(n49783) );
  NANDN U59286 ( .A(n49786), .B(n49787), .Z(n49784) );
  NANDN U59287 ( .A(n49787), .B(n49786), .Z(n49782) );
  AND U59288 ( .A(n49788), .B(n49789), .Z(n49759) );
  NAND U59289 ( .A(n49790), .B(n49791), .Z(n49789) );
  OR U59290 ( .A(n49792), .B(n49793), .Z(n49790) );
  NANDN U59291 ( .A(n49794), .B(n49792), .Z(n49788) );
  NAND U59292 ( .A(n49795), .B(n49796), .Z(n49763) );
  NANDN U59293 ( .A(n49797), .B(n49798), .Z(n49796) );
  OR U59294 ( .A(n49799), .B(n49800), .Z(n49798) );
  NANDN U59295 ( .A(n49801), .B(n49799), .Z(n49795) );
  IV U59296 ( .A(n49800), .Z(n49801) );
  XNOR U59297 ( .A(n49771), .B(n49802), .Z(n49766) );
  XNOR U59298 ( .A(n49769), .B(n49772), .Z(n49802) );
  NAND U59299 ( .A(n49803), .B(n49804), .Z(n49772) );
  NAND U59300 ( .A(n49805), .B(n49806), .Z(n49804) );
  OR U59301 ( .A(n49807), .B(n49808), .Z(n49805) );
  NANDN U59302 ( .A(n49809), .B(n49807), .Z(n49803) );
  IV U59303 ( .A(n49808), .Z(n49809) );
  NAND U59304 ( .A(n49810), .B(n49811), .Z(n49769) );
  NAND U59305 ( .A(n49812), .B(n49813), .Z(n49811) );
  NANDN U59306 ( .A(n49814), .B(n49815), .Z(n49812) );
  NANDN U59307 ( .A(n49815), .B(n49814), .Z(n49810) );
  AND U59308 ( .A(n49816), .B(n49817), .Z(n49771) );
  NAND U59309 ( .A(n49818), .B(n49819), .Z(n49817) );
  OR U59310 ( .A(n49820), .B(n49821), .Z(n49818) );
  NANDN U59311 ( .A(n49822), .B(n49820), .Z(n49816) );
  XNOR U59312 ( .A(n49797), .B(n49823), .Z(N60983) );
  XOR U59313 ( .A(n49799), .B(n49800), .Z(n49823) );
  XNOR U59314 ( .A(n49813), .B(n49824), .Z(n49800) );
  XOR U59315 ( .A(n49814), .B(n49815), .Z(n49824) );
  XOR U59316 ( .A(n49820), .B(n49825), .Z(n49815) );
  XOR U59317 ( .A(n49819), .B(n49822), .Z(n49825) );
  IV U59318 ( .A(n49821), .Z(n49822) );
  NAND U59319 ( .A(n49826), .B(n49827), .Z(n49821) );
  OR U59320 ( .A(n49828), .B(n49829), .Z(n49827) );
  OR U59321 ( .A(n49830), .B(n49831), .Z(n49826) );
  NAND U59322 ( .A(n49832), .B(n49833), .Z(n49819) );
  OR U59323 ( .A(n49834), .B(n49835), .Z(n49833) );
  OR U59324 ( .A(n49836), .B(n49837), .Z(n49832) );
  NOR U59325 ( .A(n49838), .B(n49839), .Z(n49820) );
  ANDN U59326 ( .B(n49840), .A(n49841), .Z(n49814) );
  XNOR U59327 ( .A(n49807), .B(n49842), .Z(n49813) );
  XNOR U59328 ( .A(n49806), .B(n49808), .Z(n49842) );
  NAND U59329 ( .A(n49843), .B(n49844), .Z(n49808) );
  OR U59330 ( .A(n49845), .B(n49846), .Z(n49844) );
  OR U59331 ( .A(n49847), .B(n49848), .Z(n49843) );
  NAND U59332 ( .A(n49849), .B(n49850), .Z(n49806) );
  OR U59333 ( .A(n49851), .B(n49852), .Z(n49850) );
  OR U59334 ( .A(n49853), .B(n49854), .Z(n49849) );
  ANDN U59335 ( .B(n49855), .A(n49856), .Z(n49807) );
  IV U59336 ( .A(n49857), .Z(n49855) );
  ANDN U59337 ( .B(n49858), .A(n49859), .Z(n49799) );
  XOR U59338 ( .A(n49785), .B(n49860), .Z(n49797) );
  XOR U59339 ( .A(n49786), .B(n49787), .Z(n49860) );
  XOR U59340 ( .A(n49792), .B(n49861), .Z(n49787) );
  XOR U59341 ( .A(n49791), .B(n49794), .Z(n49861) );
  IV U59342 ( .A(n49793), .Z(n49794) );
  NAND U59343 ( .A(n49862), .B(n49863), .Z(n49793) );
  OR U59344 ( .A(n49864), .B(n49865), .Z(n49863) );
  OR U59345 ( .A(n49866), .B(n49867), .Z(n49862) );
  NAND U59346 ( .A(n49868), .B(n49869), .Z(n49791) );
  OR U59347 ( .A(n49870), .B(n49871), .Z(n49869) );
  OR U59348 ( .A(n49872), .B(n49873), .Z(n49868) );
  NOR U59349 ( .A(n49874), .B(n49875), .Z(n49792) );
  ANDN U59350 ( .B(n49876), .A(n49877), .Z(n49786) );
  IV U59351 ( .A(n49878), .Z(n49876) );
  XNOR U59352 ( .A(n49779), .B(n49879), .Z(n49785) );
  XNOR U59353 ( .A(n49778), .B(n49780), .Z(n49879) );
  NAND U59354 ( .A(n49880), .B(n49881), .Z(n49780) );
  OR U59355 ( .A(n49882), .B(n49883), .Z(n49881) );
  OR U59356 ( .A(n49884), .B(n49885), .Z(n49880) );
  NAND U59357 ( .A(n49886), .B(n49887), .Z(n49778) );
  OR U59358 ( .A(n49888), .B(n49889), .Z(n49887) );
  OR U59359 ( .A(n49890), .B(n49891), .Z(n49886) );
  ANDN U59360 ( .B(n49892), .A(n49893), .Z(n49779) );
  IV U59361 ( .A(n49894), .Z(n49892) );
  XNOR U59362 ( .A(n49859), .B(n49858), .Z(N60982) );
  XOR U59363 ( .A(n49878), .B(n49877), .Z(n49858) );
  XNOR U59364 ( .A(n49893), .B(n49894), .Z(n49877) );
  XNOR U59365 ( .A(n49888), .B(n49889), .Z(n49894) );
  XNOR U59366 ( .A(n49890), .B(n49891), .Z(n49889) );
  XNOR U59367 ( .A(y[733]), .B(x[733]), .Z(n49891) );
  XNOR U59368 ( .A(y[734]), .B(x[734]), .Z(n49890) );
  XNOR U59369 ( .A(y[732]), .B(x[732]), .Z(n49888) );
  XNOR U59370 ( .A(n49882), .B(n49883), .Z(n49893) );
  XNOR U59371 ( .A(y[729]), .B(x[729]), .Z(n49883) );
  XNOR U59372 ( .A(n49884), .B(n49885), .Z(n49882) );
  XNOR U59373 ( .A(y[730]), .B(x[730]), .Z(n49885) );
  XNOR U59374 ( .A(y[731]), .B(x[731]), .Z(n49884) );
  XNOR U59375 ( .A(n49875), .B(n49874), .Z(n49878) );
  XNOR U59376 ( .A(n49870), .B(n49871), .Z(n49874) );
  XNOR U59377 ( .A(y[726]), .B(x[726]), .Z(n49871) );
  XNOR U59378 ( .A(n49872), .B(n49873), .Z(n49870) );
  XNOR U59379 ( .A(y[727]), .B(x[727]), .Z(n49873) );
  XNOR U59380 ( .A(y[728]), .B(x[728]), .Z(n49872) );
  XNOR U59381 ( .A(n49864), .B(n49865), .Z(n49875) );
  XNOR U59382 ( .A(y[723]), .B(x[723]), .Z(n49865) );
  XNOR U59383 ( .A(n49866), .B(n49867), .Z(n49864) );
  XNOR U59384 ( .A(y[724]), .B(x[724]), .Z(n49867) );
  XNOR U59385 ( .A(y[725]), .B(x[725]), .Z(n49866) );
  XOR U59386 ( .A(n49840), .B(n49841), .Z(n49859) );
  XNOR U59387 ( .A(n49856), .B(n49857), .Z(n49841) );
  XNOR U59388 ( .A(n49851), .B(n49852), .Z(n49857) );
  XNOR U59389 ( .A(n49853), .B(n49854), .Z(n49852) );
  XNOR U59390 ( .A(y[721]), .B(x[721]), .Z(n49854) );
  XNOR U59391 ( .A(y[722]), .B(x[722]), .Z(n49853) );
  XNOR U59392 ( .A(y[720]), .B(x[720]), .Z(n49851) );
  XNOR U59393 ( .A(n49845), .B(n49846), .Z(n49856) );
  XNOR U59394 ( .A(y[717]), .B(x[717]), .Z(n49846) );
  XNOR U59395 ( .A(n49847), .B(n49848), .Z(n49845) );
  XNOR U59396 ( .A(y[718]), .B(x[718]), .Z(n49848) );
  XNOR U59397 ( .A(y[719]), .B(x[719]), .Z(n49847) );
  XOR U59398 ( .A(n49839), .B(n49838), .Z(n49840) );
  XNOR U59399 ( .A(n49834), .B(n49835), .Z(n49838) );
  XNOR U59400 ( .A(y[714]), .B(x[714]), .Z(n49835) );
  XNOR U59401 ( .A(n49836), .B(n49837), .Z(n49834) );
  XNOR U59402 ( .A(y[715]), .B(x[715]), .Z(n49837) );
  XNOR U59403 ( .A(y[716]), .B(x[716]), .Z(n49836) );
  XNOR U59404 ( .A(n49828), .B(n49829), .Z(n49839) );
  XNOR U59405 ( .A(y[711]), .B(x[711]), .Z(n49829) );
  XNOR U59406 ( .A(n49830), .B(n49831), .Z(n49828) );
  XNOR U59407 ( .A(y[712]), .B(x[712]), .Z(n49831) );
  XNOR U59408 ( .A(y[713]), .B(x[713]), .Z(n49830) );
  NAND U59409 ( .A(n49895), .B(n49896), .Z(N60973) );
  NANDN U59410 ( .A(n49897), .B(n49898), .Z(n49896) );
  OR U59411 ( .A(n49899), .B(n49900), .Z(n49898) );
  NAND U59412 ( .A(n49899), .B(n49900), .Z(n49895) );
  XOR U59413 ( .A(n49899), .B(n49901), .Z(N60972) );
  XNOR U59414 ( .A(n49897), .B(n49900), .Z(n49901) );
  AND U59415 ( .A(n49902), .B(n49903), .Z(n49900) );
  NANDN U59416 ( .A(n49904), .B(n49905), .Z(n49903) );
  NANDN U59417 ( .A(n49906), .B(n49907), .Z(n49905) );
  NANDN U59418 ( .A(n49907), .B(n49906), .Z(n49902) );
  NAND U59419 ( .A(n49908), .B(n49909), .Z(n49897) );
  NANDN U59420 ( .A(n49910), .B(n49911), .Z(n49909) );
  OR U59421 ( .A(n49912), .B(n49913), .Z(n49911) );
  NAND U59422 ( .A(n49913), .B(n49912), .Z(n49908) );
  AND U59423 ( .A(n49914), .B(n49915), .Z(n49899) );
  NANDN U59424 ( .A(n49916), .B(n49917), .Z(n49915) );
  NANDN U59425 ( .A(n49918), .B(n49919), .Z(n49917) );
  NANDN U59426 ( .A(n49919), .B(n49918), .Z(n49914) );
  XOR U59427 ( .A(n49913), .B(n49920), .Z(N60971) );
  XOR U59428 ( .A(n49910), .B(n49912), .Z(n49920) );
  XNOR U59429 ( .A(n49906), .B(n49921), .Z(n49912) );
  XNOR U59430 ( .A(n49904), .B(n49907), .Z(n49921) );
  NAND U59431 ( .A(n49922), .B(n49923), .Z(n49907) );
  NAND U59432 ( .A(n49924), .B(n49925), .Z(n49923) );
  OR U59433 ( .A(n49926), .B(n49927), .Z(n49924) );
  NANDN U59434 ( .A(n49928), .B(n49926), .Z(n49922) );
  IV U59435 ( .A(n49927), .Z(n49928) );
  NAND U59436 ( .A(n49929), .B(n49930), .Z(n49904) );
  NAND U59437 ( .A(n49931), .B(n49932), .Z(n49930) );
  NANDN U59438 ( .A(n49933), .B(n49934), .Z(n49931) );
  NANDN U59439 ( .A(n49934), .B(n49933), .Z(n49929) );
  AND U59440 ( .A(n49935), .B(n49936), .Z(n49906) );
  NAND U59441 ( .A(n49937), .B(n49938), .Z(n49936) );
  OR U59442 ( .A(n49939), .B(n49940), .Z(n49937) );
  NANDN U59443 ( .A(n49941), .B(n49939), .Z(n49935) );
  NAND U59444 ( .A(n49942), .B(n49943), .Z(n49910) );
  NANDN U59445 ( .A(n49944), .B(n49945), .Z(n49943) );
  OR U59446 ( .A(n49946), .B(n49947), .Z(n49945) );
  NANDN U59447 ( .A(n49948), .B(n49946), .Z(n49942) );
  IV U59448 ( .A(n49947), .Z(n49948) );
  XNOR U59449 ( .A(n49918), .B(n49949), .Z(n49913) );
  XNOR U59450 ( .A(n49916), .B(n49919), .Z(n49949) );
  NAND U59451 ( .A(n49950), .B(n49951), .Z(n49919) );
  NAND U59452 ( .A(n49952), .B(n49953), .Z(n49951) );
  OR U59453 ( .A(n49954), .B(n49955), .Z(n49952) );
  NANDN U59454 ( .A(n49956), .B(n49954), .Z(n49950) );
  IV U59455 ( .A(n49955), .Z(n49956) );
  NAND U59456 ( .A(n49957), .B(n49958), .Z(n49916) );
  NAND U59457 ( .A(n49959), .B(n49960), .Z(n49958) );
  NANDN U59458 ( .A(n49961), .B(n49962), .Z(n49959) );
  NANDN U59459 ( .A(n49962), .B(n49961), .Z(n49957) );
  AND U59460 ( .A(n49963), .B(n49964), .Z(n49918) );
  NAND U59461 ( .A(n49965), .B(n49966), .Z(n49964) );
  OR U59462 ( .A(n49967), .B(n49968), .Z(n49965) );
  NANDN U59463 ( .A(n49969), .B(n49967), .Z(n49963) );
  XNOR U59464 ( .A(n49944), .B(n49970), .Z(N60970) );
  XOR U59465 ( .A(n49946), .B(n49947), .Z(n49970) );
  XNOR U59466 ( .A(n49960), .B(n49971), .Z(n49947) );
  XOR U59467 ( .A(n49961), .B(n49962), .Z(n49971) );
  XOR U59468 ( .A(n49967), .B(n49972), .Z(n49962) );
  XOR U59469 ( .A(n49966), .B(n49969), .Z(n49972) );
  IV U59470 ( .A(n49968), .Z(n49969) );
  NAND U59471 ( .A(n49973), .B(n49974), .Z(n49968) );
  OR U59472 ( .A(n49975), .B(n49976), .Z(n49974) );
  OR U59473 ( .A(n49977), .B(n49978), .Z(n49973) );
  NAND U59474 ( .A(n49979), .B(n49980), .Z(n49966) );
  OR U59475 ( .A(n49981), .B(n49982), .Z(n49980) );
  OR U59476 ( .A(n49983), .B(n49984), .Z(n49979) );
  NOR U59477 ( .A(n49985), .B(n49986), .Z(n49967) );
  ANDN U59478 ( .B(n49987), .A(n49988), .Z(n49961) );
  XNOR U59479 ( .A(n49954), .B(n49989), .Z(n49960) );
  XNOR U59480 ( .A(n49953), .B(n49955), .Z(n49989) );
  NAND U59481 ( .A(n49990), .B(n49991), .Z(n49955) );
  OR U59482 ( .A(n49992), .B(n49993), .Z(n49991) );
  OR U59483 ( .A(n49994), .B(n49995), .Z(n49990) );
  NAND U59484 ( .A(n49996), .B(n49997), .Z(n49953) );
  OR U59485 ( .A(n49998), .B(n49999), .Z(n49997) );
  OR U59486 ( .A(n50000), .B(n50001), .Z(n49996) );
  ANDN U59487 ( .B(n50002), .A(n50003), .Z(n49954) );
  IV U59488 ( .A(n50004), .Z(n50002) );
  ANDN U59489 ( .B(n50005), .A(n50006), .Z(n49946) );
  XOR U59490 ( .A(n49932), .B(n50007), .Z(n49944) );
  XOR U59491 ( .A(n49933), .B(n49934), .Z(n50007) );
  XOR U59492 ( .A(n49939), .B(n50008), .Z(n49934) );
  XOR U59493 ( .A(n49938), .B(n49941), .Z(n50008) );
  IV U59494 ( .A(n49940), .Z(n49941) );
  NAND U59495 ( .A(n50009), .B(n50010), .Z(n49940) );
  OR U59496 ( .A(n50011), .B(n50012), .Z(n50010) );
  OR U59497 ( .A(n50013), .B(n50014), .Z(n50009) );
  NAND U59498 ( .A(n50015), .B(n50016), .Z(n49938) );
  OR U59499 ( .A(n50017), .B(n50018), .Z(n50016) );
  OR U59500 ( .A(n50019), .B(n50020), .Z(n50015) );
  NOR U59501 ( .A(n50021), .B(n50022), .Z(n49939) );
  ANDN U59502 ( .B(n50023), .A(n50024), .Z(n49933) );
  IV U59503 ( .A(n50025), .Z(n50023) );
  XNOR U59504 ( .A(n49926), .B(n50026), .Z(n49932) );
  XNOR U59505 ( .A(n49925), .B(n49927), .Z(n50026) );
  NAND U59506 ( .A(n50027), .B(n50028), .Z(n49927) );
  OR U59507 ( .A(n50029), .B(n50030), .Z(n50028) );
  OR U59508 ( .A(n50031), .B(n50032), .Z(n50027) );
  NAND U59509 ( .A(n50033), .B(n50034), .Z(n49925) );
  OR U59510 ( .A(n50035), .B(n50036), .Z(n50034) );
  OR U59511 ( .A(n50037), .B(n50038), .Z(n50033) );
  ANDN U59512 ( .B(n50039), .A(n50040), .Z(n49926) );
  IV U59513 ( .A(n50041), .Z(n50039) );
  XNOR U59514 ( .A(n50006), .B(n50005), .Z(N60969) );
  XOR U59515 ( .A(n50025), .B(n50024), .Z(n50005) );
  XNOR U59516 ( .A(n50040), .B(n50041), .Z(n50024) );
  XNOR U59517 ( .A(n50035), .B(n50036), .Z(n50041) );
  XNOR U59518 ( .A(n50037), .B(n50038), .Z(n50036) );
  XNOR U59519 ( .A(y[709]), .B(x[709]), .Z(n50038) );
  XNOR U59520 ( .A(y[710]), .B(x[710]), .Z(n50037) );
  XNOR U59521 ( .A(y[708]), .B(x[708]), .Z(n50035) );
  XNOR U59522 ( .A(n50029), .B(n50030), .Z(n50040) );
  XNOR U59523 ( .A(y[705]), .B(x[705]), .Z(n50030) );
  XNOR U59524 ( .A(n50031), .B(n50032), .Z(n50029) );
  XNOR U59525 ( .A(y[706]), .B(x[706]), .Z(n50032) );
  XNOR U59526 ( .A(y[707]), .B(x[707]), .Z(n50031) );
  XNOR U59527 ( .A(n50022), .B(n50021), .Z(n50025) );
  XNOR U59528 ( .A(n50017), .B(n50018), .Z(n50021) );
  XNOR U59529 ( .A(y[702]), .B(x[702]), .Z(n50018) );
  XNOR U59530 ( .A(n50019), .B(n50020), .Z(n50017) );
  XNOR U59531 ( .A(y[703]), .B(x[703]), .Z(n50020) );
  XNOR U59532 ( .A(y[704]), .B(x[704]), .Z(n50019) );
  XNOR U59533 ( .A(n50011), .B(n50012), .Z(n50022) );
  XNOR U59534 ( .A(y[699]), .B(x[699]), .Z(n50012) );
  XNOR U59535 ( .A(n50013), .B(n50014), .Z(n50011) );
  XNOR U59536 ( .A(y[700]), .B(x[700]), .Z(n50014) );
  XNOR U59537 ( .A(y[701]), .B(x[701]), .Z(n50013) );
  XOR U59538 ( .A(n49987), .B(n49988), .Z(n50006) );
  XNOR U59539 ( .A(n50003), .B(n50004), .Z(n49988) );
  XNOR U59540 ( .A(n49998), .B(n49999), .Z(n50004) );
  XNOR U59541 ( .A(n50000), .B(n50001), .Z(n49999) );
  XNOR U59542 ( .A(y[697]), .B(x[697]), .Z(n50001) );
  XNOR U59543 ( .A(y[698]), .B(x[698]), .Z(n50000) );
  XNOR U59544 ( .A(y[696]), .B(x[696]), .Z(n49998) );
  XNOR U59545 ( .A(n49992), .B(n49993), .Z(n50003) );
  XNOR U59546 ( .A(y[693]), .B(x[693]), .Z(n49993) );
  XNOR U59547 ( .A(n49994), .B(n49995), .Z(n49992) );
  XNOR U59548 ( .A(y[694]), .B(x[694]), .Z(n49995) );
  XNOR U59549 ( .A(y[695]), .B(x[695]), .Z(n49994) );
  XOR U59550 ( .A(n49986), .B(n49985), .Z(n49987) );
  XNOR U59551 ( .A(n49981), .B(n49982), .Z(n49985) );
  XNOR U59552 ( .A(y[690]), .B(x[690]), .Z(n49982) );
  XNOR U59553 ( .A(n49983), .B(n49984), .Z(n49981) );
  XNOR U59554 ( .A(y[691]), .B(x[691]), .Z(n49984) );
  XNOR U59555 ( .A(y[692]), .B(x[692]), .Z(n49983) );
  XNOR U59556 ( .A(n49975), .B(n49976), .Z(n49986) );
  XNOR U59557 ( .A(y[687]), .B(x[687]), .Z(n49976) );
  XNOR U59558 ( .A(n49977), .B(n49978), .Z(n49975) );
  XNOR U59559 ( .A(y[688]), .B(x[688]), .Z(n49978) );
  XNOR U59560 ( .A(y[689]), .B(x[689]), .Z(n49977) );
  NAND U59561 ( .A(n50042), .B(n50043), .Z(N60960) );
  NANDN U59562 ( .A(n50044), .B(n50045), .Z(n50043) );
  OR U59563 ( .A(n50046), .B(n50047), .Z(n50045) );
  NAND U59564 ( .A(n50046), .B(n50047), .Z(n50042) );
  XOR U59565 ( .A(n50046), .B(n50048), .Z(N60959) );
  XNOR U59566 ( .A(n50044), .B(n50047), .Z(n50048) );
  AND U59567 ( .A(n50049), .B(n50050), .Z(n50047) );
  NANDN U59568 ( .A(n50051), .B(n50052), .Z(n50050) );
  NANDN U59569 ( .A(n50053), .B(n50054), .Z(n50052) );
  NANDN U59570 ( .A(n50054), .B(n50053), .Z(n50049) );
  NAND U59571 ( .A(n50055), .B(n50056), .Z(n50044) );
  NANDN U59572 ( .A(n50057), .B(n50058), .Z(n50056) );
  OR U59573 ( .A(n50059), .B(n50060), .Z(n50058) );
  NAND U59574 ( .A(n50060), .B(n50059), .Z(n50055) );
  AND U59575 ( .A(n50061), .B(n50062), .Z(n50046) );
  NANDN U59576 ( .A(n50063), .B(n50064), .Z(n50062) );
  NANDN U59577 ( .A(n50065), .B(n50066), .Z(n50064) );
  NANDN U59578 ( .A(n50066), .B(n50065), .Z(n50061) );
  XOR U59579 ( .A(n50060), .B(n50067), .Z(N60958) );
  XOR U59580 ( .A(n50057), .B(n50059), .Z(n50067) );
  XNOR U59581 ( .A(n50053), .B(n50068), .Z(n50059) );
  XNOR U59582 ( .A(n50051), .B(n50054), .Z(n50068) );
  NAND U59583 ( .A(n50069), .B(n50070), .Z(n50054) );
  NAND U59584 ( .A(n50071), .B(n50072), .Z(n50070) );
  OR U59585 ( .A(n50073), .B(n50074), .Z(n50071) );
  NANDN U59586 ( .A(n50075), .B(n50073), .Z(n50069) );
  IV U59587 ( .A(n50074), .Z(n50075) );
  NAND U59588 ( .A(n50076), .B(n50077), .Z(n50051) );
  NAND U59589 ( .A(n50078), .B(n50079), .Z(n50077) );
  NANDN U59590 ( .A(n50080), .B(n50081), .Z(n50078) );
  NANDN U59591 ( .A(n50081), .B(n50080), .Z(n50076) );
  AND U59592 ( .A(n50082), .B(n50083), .Z(n50053) );
  NAND U59593 ( .A(n50084), .B(n50085), .Z(n50083) );
  OR U59594 ( .A(n50086), .B(n50087), .Z(n50084) );
  NANDN U59595 ( .A(n50088), .B(n50086), .Z(n50082) );
  NAND U59596 ( .A(n50089), .B(n50090), .Z(n50057) );
  NANDN U59597 ( .A(n50091), .B(n50092), .Z(n50090) );
  OR U59598 ( .A(n50093), .B(n50094), .Z(n50092) );
  NANDN U59599 ( .A(n50095), .B(n50093), .Z(n50089) );
  IV U59600 ( .A(n50094), .Z(n50095) );
  XNOR U59601 ( .A(n50065), .B(n50096), .Z(n50060) );
  XNOR U59602 ( .A(n50063), .B(n50066), .Z(n50096) );
  NAND U59603 ( .A(n50097), .B(n50098), .Z(n50066) );
  NAND U59604 ( .A(n50099), .B(n50100), .Z(n50098) );
  OR U59605 ( .A(n50101), .B(n50102), .Z(n50099) );
  NANDN U59606 ( .A(n50103), .B(n50101), .Z(n50097) );
  IV U59607 ( .A(n50102), .Z(n50103) );
  NAND U59608 ( .A(n50104), .B(n50105), .Z(n50063) );
  NAND U59609 ( .A(n50106), .B(n50107), .Z(n50105) );
  NANDN U59610 ( .A(n50108), .B(n50109), .Z(n50106) );
  NANDN U59611 ( .A(n50109), .B(n50108), .Z(n50104) );
  AND U59612 ( .A(n50110), .B(n50111), .Z(n50065) );
  NAND U59613 ( .A(n50112), .B(n50113), .Z(n50111) );
  OR U59614 ( .A(n50114), .B(n50115), .Z(n50112) );
  NANDN U59615 ( .A(n50116), .B(n50114), .Z(n50110) );
  XNOR U59616 ( .A(n50091), .B(n50117), .Z(N60957) );
  XOR U59617 ( .A(n50093), .B(n50094), .Z(n50117) );
  XNOR U59618 ( .A(n50107), .B(n50118), .Z(n50094) );
  XOR U59619 ( .A(n50108), .B(n50109), .Z(n50118) );
  XOR U59620 ( .A(n50114), .B(n50119), .Z(n50109) );
  XOR U59621 ( .A(n50113), .B(n50116), .Z(n50119) );
  IV U59622 ( .A(n50115), .Z(n50116) );
  NAND U59623 ( .A(n50120), .B(n50121), .Z(n50115) );
  OR U59624 ( .A(n50122), .B(n50123), .Z(n50121) );
  OR U59625 ( .A(n50124), .B(n50125), .Z(n50120) );
  NAND U59626 ( .A(n50126), .B(n50127), .Z(n50113) );
  OR U59627 ( .A(n50128), .B(n50129), .Z(n50127) );
  OR U59628 ( .A(n50130), .B(n50131), .Z(n50126) );
  NOR U59629 ( .A(n50132), .B(n50133), .Z(n50114) );
  ANDN U59630 ( .B(n50134), .A(n50135), .Z(n50108) );
  XNOR U59631 ( .A(n50101), .B(n50136), .Z(n50107) );
  XNOR U59632 ( .A(n50100), .B(n50102), .Z(n50136) );
  NAND U59633 ( .A(n50137), .B(n50138), .Z(n50102) );
  OR U59634 ( .A(n50139), .B(n50140), .Z(n50138) );
  OR U59635 ( .A(n50141), .B(n50142), .Z(n50137) );
  NAND U59636 ( .A(n50143), .B(n50144), .Z(n50100) );
  OR U59637 ( .A(n50145), .B(n50146), .Z(n50144) );
  OR U59638 ( .A(n50147), .B(n50148), .Z(n50143) );
  ANDN U59639 ( .B(n50149), .A(n50150), .Z(n50101) );
  IV U59640 ( .A(n50151), .Z(n50149) );
  ANDN U59641 ( .B(n50152), .A(n50153), .Z(n50093) );
  XOR U59642 ( .A(n50079), .B(n50154), .Z(n50091) );
  XOR U59643 ( .A(n50080), .B(n50081), .Z(n50154) );
  XOR U59644 ( .A(n50086), .B(n50155), .Z(n50081) );
  XOR U59645 ( .A(n50085), .B(n50088), .Z(n50155) );
  IV U59646 ( .A(n50087), .Z(n50088) );
  NAND U59647 ( .A(n50156), .B(n50157), .Z(n50087) );
  OR U59648 ( .A(n50158), .B(n50159), .Z(n50157) );
  OR U59649 ( .A(n50160), .B(n50161), .Z(n50156) );
  NAND U59650 ( .A(n50162), .B(n50163), .Z(n50085) );
  OR U59651 ( .A(n50164), .B(n50165), .Z(n50163) );
  OR U59652 ( .A(n50166), .B(n50167), .Z(n50162) );
  NOR U59653 ( .A(n50168), .B(n50169), .Z(n50086) );
  ANDN U59654 ( .B(n50170), .A(n50171), .Z(n50080) );
  IV U59655 ( .A(n50172), .Z(n50170) );
  XNOR U59656 ( .A(n50073), .B(n50173), .Z(n50079) );
  XNOR U59657 ( .A(n50072), .B(n50074), .Z(n50173) );
  NAND U59658 ( .A(n50174), .B(n50175), .Z(n50074) );
  OR U59659 ( .A(n50176), .B(n50177), .Z(n50175) );
  OR U59660 ( .A(n50178), .B(n50179), .Z(n50174) );
  NAND U59661 ( .A(n50180), .B(n50181), .Z(n50072) );
  OR U59662 ( .A(n50182), .B(n50183), .Z(n50181) );
  OR U59663 ( .A(n50184), .B(n50185), .Z(n50180) );
  ANDN U59664 ( .B(n50186), .A(n50187), .Z(n50073) );
  IV U59665 ( .A(n50188), .Z(n50186) );
  XNOR U59666 ( .A(n50153), .B(n50152), .Z(N60956) );
  XOR U59667 ( .A(n50172), .B(n50171), .Z(n50152) );
  XNOR U59668 ( .A(n50187), .B(n50188), .Z(n50171) );
  XNOR U59669 ( .A(n50182), .B(n50183), .Z(n50188) );
  XNOR U59670 ( .A(n50184), .B(n50185), .Z(n50183) );
  XNOR U59671 ( .A(y[685]), .B(x[685]), .Z(n50185) );
  XNOR U59672 ( .A(y[686]), .B(x[686]), .Z(n50184) );
  XNOR U59673 ( .A(y[684]), .B(x[684]), .Z(n50182) );
  XNOR U59674 ( .A(n50176), .B(n50177), .Z(n50187) );
  XNOR U59675 ( .A(y[681]), .B(x[681]), .Z(n50177) );
  XNOR U59676 ( .A(n50178), .B(n50179), .Z(n50176) );
  XNOR U59677 ( .A(y[682]), .B(x[682]), .Z(n50179) );
  XNOR U59678 ( .A(y[683]), .B(x[683]), .Z(n50178) );
  XNOR U59679 ( .A(n50169), .B(n50168), .Z(n50172) );
  XNOR U59680 ( .A(n50164), .B(n50165), .Z(n50168) );
  XNOR U59681 ( .A(y[678]), .B(x[678]), .Z(n50165) );
  XNOR U59682 ( .A(n50166), .B(n50167), .Z(n50164) );
  XNOR U59683 ( .A(y[679]), .B(x[679]), .Z(n50167) );
  XNOR U59684 ( .A(y[680]), .B(x[680]), .Z(n50166) );
  XNOR U59685 ( .A(n50158), .B(n50159), .Z(n50169) );
  XNOR U59686 ( .A(y[675]), .B(x[675]), .Z(n50159) );
  XNOR U59687 ( .A(n50160), .B(n50161), .Z(n50158) );
  XNOR U59688 ( .A(y[676]), .B(x[676]), .Z(n50161) );
  XNOR U59689 ( .A(y[677]), .B(x[677]), .Z(n50160) );
  XOR U59690 ( .A(n50134), .B(n50135), .Z(n50153) );
  XNOR U59691 ( .A(n50150), .B(n50151), .Z(n50135) );
  XNOR U59692 ( .A(n50145), .B(n50146), .Z(n50151) );
  XNOR U59693 ( .A(n50147), .B(n50148), .Z(n50146) );
  XNOR U59694 ( .A(y[673]), .B(x[673]), .Z(n50148) );
  XNOR U59695 ( .A(y[674]), .B(x[674]), .Z(n50147) );
  XNOR U59696 ( .A(y[672]), .B(x[672]), .Z(n50145) );
  XNOR U59697 ( .A(n50139), .B(n50140), .Z(n50150) );
  XNOR U59698 ( .A(y[669]), .B(x[669]), .Z(n50140) );
  XNOR U59699 ( .A(n50141), .B(n50142), .Z(n50139) );
  XNOR U59700 ( .A(y[670]), .B(x[670]), .Z(n50142) );
  XNOR U59701 ( .A(y[671]), .B(x[671]), .Z(n50141) );
  XOR U59702 ( .A(n50133), .B(n50132), .Z(n50134) );
  XNOR U59703 ( .A(n50128), .B(n50129), .Z(n50132) );
  XNOR U59704 ( .A(y[666]), .B(x[666]), .Z(n50129) );
  XNOR U59705 ( .A(n50130), .B(n50131), .Z(n50128) );
  XNOR U59706 ( .A(y[667]), .B(x[667]), .Z(n50131) );
  XNOR U59707 ( .A(y[668]), .B(x[668]), .Z(n50130) );
  XNOR U59708 ( .A(n50122), .B(n50123), .Z(n50133) );
  XNOR U59709 ( .A(y[663]), .B(x[663]), .Z(n50123) );
  XNOR U59710 ( .A(n50124), .B(n50125), .Z(n50122) );
  XNOR U59711 ( .A(y[664]), .B(x[664]), .Z(n50125) );
  XNOR U59712 ( .A(y[665]), .B(x[665]), .Z(n50124) );
  NAND U59713 ( .A(n50189), .B(n50190), .Z(N60947) );
  NANDN U59714 ( .A(n50191), .B(n50192), .Z(n50190) );
  OR U59715 ( .A(n50193), .B(n50194), .Z(n50192) );
  NAND U59716 ( .A(n50193), .B(n50194), .Z(n50189) );
  XOR U59717 ( .A(n50193), .B(n50195), .Z(N60946) );
  XNOR U59718 ( .A(n50191), .B(n50194), .Z(n50195) );
  AND U59719 ( .A(n50196), .B(n50197), .Z(n50194) );
  NANDN U59720 ( .A(n50198), .B(n50199), .Z(n50197) );
  NANDN U59721 ( .A(n50200), .B(n50201), .Z(n50199) );
  NANDN U59722 ( .A(n50201), .B(n50200), .Z(n50196) );
  NAND U59723 ( .A(n50202), .B(n50203), .Z(n50191) );
  NANDN U59724 ( .A(n50204), .B(n50205), .Z(n50203) );
  OR U59725 ( .A(n50206), .B(n50207), .Z(n50205) );
  NAND U59726 ( .A(n50207), .B(n50206), .Z(n50202) );
  AND U59727 ( .A(n50208), .B(n50209), .Z(n50193) );
  NANDN U59728 ( .A(n50210), .B(n50211), .Z(n50209) );
  NANDN U59729 ( .A(n50212), .B(n50213), .Z(n50211) );
  NANDN U59730 ( .A(n50213), .B(n50212), .Z(n50208) );
  XOR U59731 ( .A(n50207), .B(n50214), .Z(N60945) );
  XOR U59732 ( .A(n50204), .B(n50206), .Z(n50214) );
  XNOR U59733 ( .A(n50200), .B(n50215), .Z(n50206) );
  XNOR U59734 ( .A(n50198), .B(n50201), .Z(n50215) );
  NAND U59735 ( .A(n50216), .B(n50217), .Z(n50201) );
  NAND U59736 ( .A(n50218), .B(n50219), .Z(n50217) );
  OR U59737 ( .A(n50220), .B(n50221), .Z(n50218) );
  NANDN U59738 ( .A(n50222), .B(n50220), .Z(n50216) );
  IV U59739 ( .A(n50221), .Z(n50222) );
  NAND U59740 ( .A(n50223), .B(n50224), .Z(n50198) );
  NAND U59741 ( .A(n50225), .B(n50226), .Z(n50224) );
  NANDN U59742 ( .A(n50227), .B(n50228), .Z(n50225) );
  NANDN U59743 ( .A(n50228), .B(n50227), .Z(n50223) );
  AND U59744 ( .A(n50229), .B(n50230), .Z(n50200) );
  NAND U59745 ( .A(n50231), .B(n50232), .Z(n50230) );
  OR U59746 ( .A(n50233), .B(n50234), .Z(n50231) );
  NANDN U59747 ( .A(n50235), .B(n50233), .Z(n50229) );
  NAND U59748 ( .A(n50236), .B(n50237), .Z(n50204) );
  NANDN U59749 ( .A(n50238), .B(n50239), .Z(n50237) );
  OR U59750 ( .A(n50240), .B(n50241), .Z(n50239) );
  NANDN U59751 ( .A(n50242), .B(n50240), .Z(n50236) );
  IV U59752 ( .A(n50241), .Z(n50242) );
  XNOR U59753 ( .A(n50212), .B(n50243), .Z(n50207) );
  XNOR U59754 ( .A(n50210), .B(n50213), .Z(n50243) );
  NAND U59755 ( .A(n50244), .B(n50245), .Z(n50213) );
  NAND U59756 ( .A(n50246), .B(n50247), .Z(n50245) );
  OR U59757 ( .A(n50248), .B(n50249), .Z(n50246) );
  NANDN U59758 ( .A(n50250), .B(n50248), .Z(n50244) );
  IV U59759 ( .A(n50249), .Z(n50250) );
  NAND U59760 ( .A(n50251), .B(n50252), .Z(n50210) );
  NAND U59761 ( .A(n50253), .B(n50254), .Z(n50252) );
  NANDN U59762 ( .A(n50255), .B(n50256), .Z(n50253) );
  NANDN U59763 ( .A(n50256), .B(n50255), .Z(n50251) );
  AND U59764 ( .A(n50257), .B(n50258), .Z(n50212) );
  NAND U59765 ( .A(n50259), .B(n50260), .Z(n50258) );
  OR U59766 ( .A(n50261), .B(n50262), .Z(n50259) );
  NANDN U59767 ( .A(n50263), .B(n50261), .Z(n50257) );
  XNOR U59768 ( .A(n50238), .B(n50264), .Z(N60944) );
  XOR U59769 ( .A(n50240), .B(n50241), .Z(n50264) );
  XNOR U59770 ( .A(n50254), .B(n50265), .Z(n50241) );
  XOR U59771 ( .A(n50255), .B(n50256), .Z(n50265) );
  XOR U59772 ( .A(n50261), .B(n50266), .Z(n50256) );
  XOR U59773 ( .A(n50260), .B(n50263), .Z(n50266) );
  IV U59774 ( .A(n50262), .Z(n50263) );
  NAND U59775 ( .A(n50267), .B(n50268), .Z(n50262) );
  OR U59776 ( .A(n50269), .B(n50270), .Z(n50268) );
  OR U59777 ( .A(n50271), .B(n50272), .Z(n50267) );
  NAND U59778 ( .A(n50273), .B(n50274), .Z(n50260) );
  OR U59779 ( .A(n50275), .B(n50276), .Z(n50274) );
  OR U59780 ( .A(n50277), .B(n50278), .Z(n50273) );
  NOR U59781 ( .A(n50279), .B(n50280), .Z(n50261) );
  ANDN U59782 ( .B(n50281), .A(n50282), .Z(n50255) );
  XNOR U59783 ( .A(n50248), .B(n50283), .Z(n50254) );
  XNOR U59784 ( .A(n50247), .B(n50249), .Z(n50283) );
  NAND U59785 ( .A(n50284), .B(n50285), .Z(n50249) );
  OR U59786 ( .A(n50286), .B(n50287), .Z(n50285) );
  OR U59787 ( .A(n50288), .B(n50289), .Z(n50284) );
  NAND U59788 ( .A(n50290), .B(n50291), .Z(n50247) );
  OR U59789 ( .A(n50292), .B(n50293), .Z(n50291) );
  OR U59790 ( .A(n50294), .B(n50295), .Z(n50290) );
  ANDN U59791 ( .B(n50296), .A(n50297), .Z(n50248) );
  IV U59792 ( .A(n50298), .Z(n50296) );
  ANDN U59793 ( .B(n50299), .A(n50300), .Z(n50240) );
  XOR U59794 ( .A(n50226), .B(n50301), .Z(n50238) );
  XOR U59795 ( .A(n50227), .B(n50228), .Z(n50301) );
  XOR U59796 ( .A(n50233), .B(n50302), .Z(n50228) );
  XOR U59797 ( .A(n50232), .B(n50235), .Z(n50302) );
  IV U59798 ( .A(n50234), .Z(n50235) );
  NAND U59799 ( .A(n50303), .B(n50304), .Z(n50234) );
  OR U59800 ( .A(n50305), .B(n50306), .Z(n50304) );
  OR U59801 ( .A(n50307), .B(n50308), .Z(n50303) );
  NAND U59802 ( .A(n50309), .B(n50310), .Z(n50232) );
  OR U59803 ( .A(n50311), .B(n50312), .Z(n50310) );
  OR U59804 ( .A(n50313), .B(n50314), .Z(n50309) );
  NOR U59805 ( .A(n50315), .B(n50316), .Z(n50233) );
  ANDN U59806 ( .B(n50317), .A(n50318), .Z(n50227) );
  IV U59807 ( .A(n50319), .Z(n50317) );
  XNOR U59808 ( .A(n50220), .B(n50320), .Z(n50226) );
  XNOR U59809 ( .A(n50219), .B(n50221), .Z(n50320) );
  NAND U59810 ( .A(n50321), .B(n50322), .Z(n50221) );
  OR U59811 ( .A(n50323), .B(n50324), .Z(n50322) );
  OR U59812 ( .A(n50325), .B(n50326), .Z(n50321) );
  NAND U59813 ( .A(n50327), .B(n50328), .Z(n50219) );
  OR U59814 ( .A(n50329), .B(n50330), .Z(n50328) );
  OR U59815 ( .A(n50331), .B(n50332), .Z(n50327) );
  ANDN U59816 ( .B(n50333), .A(n50334), .Z(n50220) );
  IV U59817 ( .A(n50335), .Z(n50333) );
  XNOR U59818 ( .A(n50300), .B(n50299), .Z(N60943) );
  XOR U59819 ( .A(n50319), .B(n50318), .Z(n50299) );
  XNOR U59820 ( .A(n50334), .B(n50335), .Z(n50318) );
  XNOR U59821 ( .A(n50329), .B(n50330), .Z(n50335) );
  XNOR U59822 ( .A(n50331), .B(n50332), .Z(n50330) );
  XNOR U59823 ( .A(y[661]), .B(x[661]), .Z(n50332) );
  XNOR U59824 ( .A(y[662]), .B(x[662]), .Z(n50331) );
  XNOR U59825 ( .A(y[660]), .B(x[660]), .Z(n50329) );
  XNOR U59826 ( .A(n50323), .B(n50324), .Z(n50334) );
  XNOR U59827 ( .A(y[657]), .B(x[657]), .Z(n50324) );
  XNOR U59828 ( .A(n50325), .B(n50326), .Z(n50323) );
  XNOR U59829 ( .A(y[658]), .B(x[658]), .Z(n50326) );
  XNOR U59830 ( .A(y[659]), .B(x[659]), .Z(n50325) );
  XNOR U59831 ( .A(n50316), .B(n50315), .Z(n50319) );
  XNOR U59832 ( .A(n50311), .B(n50312), .Z(n50315) );
  XNOR U59833 ( .A(y[654]), .B(x[654]), .Z(n50312) );
  XNOR U59834 ( .A(n50313), .B(n50314), .Z(n50311) );
  XNOR U59835 ( .A(y[655]), .B(x[655]), .Z(n50314) );
  XNOR U59836 ( .A(y[656]), .B(x[656]), .Z(n50313) );
  XNOR U59837 ( .A(n50305), .B(n50306), .Z(n50316) );
  XNOR U59838 ( .A(y[651]), .B(x[651]), .Z(n50306) );
  XNOR U59839 ( .A(n50307), .B(n50308), .Z(n50305) );
  XNOR U59840 ( .A(y[652]), .B(x[652]), .Z(n50308) );
  XNOR U59841 ( .A(y[653]), .B(x[653]), .Z(n50307) );
  XOR U59842 ( .A(n50281), .B(n50282), .Z(n50300) );
  XNOR U59843 ( .A(n50297), .B(n50298), .Z(n50282) );
  XNOR U59844 ( .A(n50292), .B(n50293), .Z(n50298) );
  XNOR U59845 ( .A(n50294), .B(n50295), .Z(n50293) );
  XNOR U59846 ( .A(y[649]), .B(x[649]), .Z(n50295) );
  XNOR U59847 ( .A(y[650]), .B(x[650]), .Z(n50294) );
  XNOR U59848 ( .A(y[648]), .B(x[648]), .Z(n50292) );
  XNOR U59849 ( .A(n50286), .B(n50287), .Z(n50297) );
  XNOR U59850 ( .A(y[645]), .B(x[645]), .Z(n50287) );
  XNOR U59851 ( .A(n50288), .B(n50289), .Z(n50286) );
  XNOR U59852 ( .A(y[646]), .B(x[646]), .Z(n50289) );
  XNOR U59853 ( .A(y[647]), .B(x[647]), .Z(n50288) );
  XOR U59854 ( .A(n50280), .B(n50279), .Z(n50281) );
  XNOR U59855 ( .A(n50275), .B(n50276), .Z(n50279) );
  XNOR U59856 ( .A(y[642]), .B(x[642]), .Z(n50276) );
  XNOR U59857 ( .A(n50277), .B(n50278), .Z(n50275) );
  XNOR U59858 ( .A(y[643]), .B(x[643]), .Z(n50278) );
  XNOR U59859 ( .A(y[644]), .B(x[644]), .Z(n50277) );
  XNOR U59860 ( .A(n50269), .B(n50270), .Z(n50280) );
  XNOR U59861 ( .A(y[639]), .B(x[639]), .Z(n50270) );
  XNOR U59862 ( .A(n50271), .B(n50272), .Z(n50269) );
  XNOR U59863 ( .A(y[640]), .B(x[640]), .Z(n50272) );
  XNOR U59864 ( .A(y[641]), .B(x[641]), .Z(n50271) );
  NAND U59865 ( .A(n50336), .B(n50337), .Z(N60934) );
  NANDN U59866 ( .A(n50338), .B(n50339), .Z(n50337) );
  OR U59867 ( .A(n50340), .B(n50341), .Z(n50339) );
  NAND U59868 ( .A(n50340), .B(n50341), .Z(n50336) );
  XOR U59869 ( .A(n50340), .B(n50342), .Z(N60933) );
  XNOR U59870 ( .A(n50338), .B(n50341), .Z(n50342) );
  AND U59871 ( .A(n50343), .B(n50344), .Z(n50341) );
  NANDN U59872 ( .A(n50345), .B(n50346), .Z(n50344) );
  NANDN U59873 ( .A(n50347), .B(n50348), .Z(n50346) );
  NANDN U59874 ( .A(n50348), .B(n50347), .Z(n50343) );
  NAND U59875 ( .A(n50349), .B(n50350), .Z(n50338) );
  NANDN U59876 ( .A(n50351), .B(n50352), .Z(n50350) );
  OR U59877 ( .A(n50353), .B(n50354), .Z(n50352) );
  NAND U59878 ( .A(n50354), .B(n50353), .Z(n50349) );
  AND U59879 ( .A(n50355), .B(n50356), .Z(n50340) );
  NANDN U59880 ( .A(n50357), .B(n50358), .Z(n50356) );
  NANDN U59881 ( .A(n50359), .B(n50360), .Z(n50358) );
  NANDN U59882 ( .A(n50360), .B(n50359), .Z(n50355) );
  XOR U59883 ( .A(n50354), .B(n50361), .Z(N60932) );
  XOR U59884 ( .A(n50351), .B(n50353), .Z(n50361) );
  XNOR U59885 ( .A(n50347), .B(n50362), .Z(n50353) );
  XNOR U59886 ( .A(n50345), .B(n50348), .Z(n50362) );
  NAND U59887 ( .A(n50363), .B(n50364), .Z(n50348) );
  NAND U59888 ( .A(n50365), .B(n50366), .Z(n50364) );
  OR U59889 ( .A(n50367), .B(n50368), .Z(n50365) );
  NANDN U59890 ( .A(n50369), .B(n50367), .Z(n50363) );
  IV U59891 ( .A(n50368), .Z(n50369) );
  NAND U59892 ( .A(n50370), .B(n50371), .Z(n50345) );
  NAND U59893 ( .A(n50372), .B(n50373), .Z(n50371) );
  NANDN U59894 ( .A(n50374), .B(n50375), .Z(n50372) );
  NANDN U59895 ( .A(n50375), .B(n50374), .Z(n50370) );
  AND U59896 ( .A(n50376), .B(n50377), .Z(n50347) );
  NAND U59897 ( .A(n50378), .B(n50379), .Z(n50377) );
  OR U59898 ( .A(n50380), .B(n50381), .Z(n50378) );
  NANDN U59899 ( .A(n50382), .B(n50380), .Z(n50376) );
  NAND U59900 ( .A(n50383), .B(n50384), .Z(n50351) );
  NANDN U59901 ( .A(n50385), .B(n50386), .Z(n50384) );
  OR U59902 ( .A(n50387), .B(n50388), .Z(n50386) );
  NANDN U59903 ( .A(n50389), .B(n50387), .Z(n50383) );
  IV U59904 ( .A(n50388), .Z(n50389) );
  XNOR U59905 ( .A(n50359), .B(n50390), .Z(n50354) );
  XNOR U59906 ( .A(n50357), .B(n50360), .Z(n50390) );
  NAND U59907 ( .A(n50391), .B(n50392), .Z(n50360) );
  NAND U59908 ( .A(n50393), .B(n50394), .Z(n50392) );
  OR U59909 ( .A(n50395), .B(n50396), .Z(n50393) );
  NANDN U59910 ( .A(n50397), .B(n50395), .Z(n50391) );
  IV U59911 ( .A(n50396), .Z(n50397) );
  NAND U59912 ( .A(n50398), .B(n50399), .Z(n50357) );
  NAND U59913 ( .A(n50400), .B(n50401), .Z(n50399) );
  NANDN U59914 ( .A(n50402), .B(n50403), .Z(n50400) );
  NANDN U59915 ( .A(n50403), .B(n50402), .Z(n50398) );
  AND U59916 ( .A(n50404), .B(n50405), .Z(n50359) );
  NAND U59917 ( .A(n50406), .B(n50407), .Z(n50405) );
  OR U59918 ( .A(n50408), .B(n50409), .Z(n50406) );
  NANDN U59919 ( .A(n50410), .B(n50408), .Z(n50404) );
  XNOR U59920 ( .A(n50385), .B(n50411), .Z(N60931) );
  XOR U59921 ( .A(n50387), .B(n50388), .Z(n50411) );
  XNOR U59922 ( .A(n50401), .B(n50412), .Z(n50388) );
  XOR U59923 ( .A(n50402), .B(n50403), .Z(n50412) );
  XOR U59924 ( .A(n50408), .B(n50413), .Z(n50403) );
  XOR U59925 ( .A(n50407), .B(n50410), .Z(n50413) );
  IV U59926 ( .A(n50409), .Z(n50410) );
  NAND U59927 ( .A(n50414), .B(n50415), .Z(n50409) );
  OR U59928 ( .A(n50416), .B(n50417), .Z(n50415) );
  OR U59929 ( .A(n50418), .B(n50419), .Z(n50414) );
  NAND U59930 ( .A(n50420), .B(n50421), .Z(n50407) );
  OR U59931 ( .A(n50422), .B(n50423), .Z(n50421) );
  OR U59932 ( .A(n50424), .B(n50425), .Z(n50420) );
  NOR U59933 ( .A(n50426), .B(n50427), .Z(n50408) );
  ANDN U59934 ( .B(n50428), .A(n50429), .Z(n50402) );
  XNOR U59935 ( .A(n50395), .B(n50430), .Z(n50401) );
  XNOR U59936 ( .A(n50394), .B(n50396), .Z(n50430) );
  NAND U59937 ( .A(n50431), .B(n50432), .Z(n50396) );
  OR U59938 ( .A(n50433), .B(n50434), .Z(n50432) );
  OR U59939 ( .A(n50435), .B(n50436), .Z(n50431) );
  NAND U59940 ( .A(n50437), .B(n50438), .Z(n50394) );
  OR U59941 ( .A(n50439), .B(n50440), .Z(n50438) );
  OR U59942 ( .A(n50441), .B(n50442), .Z(n50437) );
  ANDN U59943 ( .B(n50443), .A(n50444), .Z(n50395) );
  IV U59944 ( .A(n50445), .Z(n50443) );
  ANDN U59945 ( .B(n50446), .A(n50447), .Z(n50387) );
  XOR U59946 ( .A(n50373), .B(n50448), .Z(n50385) );
  XOR U59947 ( .A(n50374), .B(n50375), .Z(n50448) );
  XOR U59948 ( .A(n50380), .B(n50449), .Z(n50375) );
  XOR U59949 ( .A(n50379), .B(n50382), .Z(n50449) );
  IV U59950 ( .A(n50381), .Z(n50382) );
  NAND U59951 ( .A(n50450), .B(n50451), .Z(n50381) );
  OR U59952 ( .A(n50452), .B(n50453), .Z(n50451) );
  OR U59953 ( .A(n50454), .B(n50455), .Z(n50450) );
  NAND U59954 ( .A(n50456), .B(n50457), .Z(n50379) );
  OR U59955 ( .A(n50458), .B(n50459), .Z(n50457) );
  OR U59956 ( .A(n50460), .B(n50461), .Z(n50456) );
  NOR U59957 ( .A(n50462), .B(n50463), .Z(n50380) );
  ANDN U59958 ( .B(n50464), .A(n50465), .Z(n50374) );
  IV U59959 ( .A(n50466), .Z(n50464) );
  XNOR U59960 ( .A(n50367), .B(n50467), .Z(n50373) );
  XNOR U59961 ( .A(n50366), .B(n50368), .Z(n50467) );
  NAND U59962 ( .A(n50468), .B(n50469), .Z(n50368) );
  OR U59963 ( .A(n50470), .B(n50471), .Z(n50469) );
  OR U59964 ( .A(n50472), .B(n50473), .Z(n50468) );
  NAND U59965 ( .A(n50474), .B(n50475), .Z(n50366) );
  OR U59966 ( .A(n50476), .B(n50477), .Z(n50475) );
  OR U59967 ( .A(n50478), .B(n50479), .Z(n50474) );
  ANDN U59968 ( .B(n50480), .A(n50481), .Z(n50367) );
  IV U59969 ( .A(n50482), .Z(n50480) );
  XNOR U59970 ( .A(n50447), .B(n50446), .Z(N60930) );
  XOR U59971 ( .A(n50466), .B(n50465), .Z(n50446) );
  XNOR U59972 ( .A(n50481), .B(n50482), .Z(n50465) );
  XNOR U59973 ( .A(n50476), .B(n50477), .Z(n50482) );
  XNOR U59974 ( .A(n50478), .B(n50479), .Z(n50477) );
  XNOR U59975 ( .A(y[637]), .B(x[637]), .Z(n50479) );
  XNOR U59976 ( .A(y[638]), .B(x[638]), .Z(n50478) );
  XNOR U59977 ( .A(y[636]), .B(x[636]), .Z(n50476) );
  XNOR U59978 ( .A(n50470), .B(n50471), .Z(n50481) );
  XNOR U59979 ( .A(y[633]), .B(x[633]), .Z(n50471) );
  XNOR U59980 ( .A(n50472), .B(n50473), .Z(n50470) );
  XNOR U59981 ( .A(y[634]), .B(x[634]), .Z(n50473) );
  XNOR U59982 ( .A(y[635]), .B(x[635]), .Z(n50472) );
  XNOR U59983 ( .A(n50463), .B(n50462), .Z(n50466) );
  XNOR U59984 ( .A(n50458), .B(n50459), .Z(n50462) );
  XNOR U59985 ( .A(y[630]), .B(x[630]), .Z(n50459) );
  XNOR U59986 ( .A(n50460), .B(n50461), .Z(n50458) );
  XNOR U59987 ( .A(y[631]), .B(x[631]), .Z(n50461) );
  XNOR U59988 ( .A(y[632]), .B(x[632]), .Z(n50460) );
  XNOR U59989 ( .A(n50452), .B(n50453), .Z(n50463) );
  XNOR U59990 ( .A(y[627]), .B(x[627]), .Z(n50453) );
  XNOR U59991 ( .A(n50454), .B(n50455), .Z(n50452) );
  XNOR U59992 ( .A(y[628]), .B(x[628]), .Z(n50455) );
  XNOR U59993 ( .A(y[629]), .B(x[629]), .Z(n50454) );
  XOR U59994 ( .A(n50428), .B(n50429), .Z(n50447) );
  XNOR U59995 ( .A(n50444), .B(n50445), .Z(n50429) );
  XNOR U59996 ( .A(n50439), .B(n50440), .Z(n50445) );
  XNOR U59997 ( .A(n50441), .B(n50442), .Z(n50440) );
  XNOR U59998 ( .A(y[625]), .B(x[625]), .Z(n50442) );
  XNOR U59999 ( .A(y[626]), .B(x[626]), .Z(n50441) );
  XNOR U60000 ( .A(y[624]), .B(x[624]), .Z(n50439) );
  XNOR U60001 ( .A(n50433), .B(n50434), .Z(n50444) );
  XNOR U60002 ( .A(y[621]), .B(x[621]), .Z(n50434) );
  XNOR U60003 ( .A(n50435), .B(n50436), .Z(n50433) );
  XNOR U60004 ( .A(y[622]), .B(x[622]), .Z(n50436) );
  XNOR U60005 ( .A(y[623]), .B(x[623]), .Z(n50435) );
  XOR U60006 ( .A(n50427), .B(n50426), .Z(n50428) );
  XNOR U60007 ( .A(n50422), .B(n50423), .Z(n50426) );
  XNOR U60008 ( .A(y[618]), .B(x[618]), .Z(n50423) );
  XNOR U60009 ( .A(n50424), .B(n50425), .Z(n50422) );
  XNOR U60010 ( .A(y[619]), .B(x[619]), .Z(n50425) );
  XNOR U60011 ( .A(y[620]), .B(x[620]), .Z(n50424) );
  XNOR U60012 ( .A(n50416), .B(n50417), .Z(n50427) );
  XNOR U60013 ( .A(y[615]), .B(x[615]), .Z(n50417) );
  XNOR U60014 ( .A(n50418), .B(n50419), .Z(n50416) );
  XNOR U60015 ( .A(y[616]), .B(x[616]), .Z(n50419) );
  XNOR U60016 ( .A(y[617]), .B(x[617]), .Z(n50418) );
  NAND U60017 ( .A(n50483), .B(n50484), .Z(N60921) );
  NANDN U60018 ( .A(n50485), .B(n50486), .Z(n50484) );
  OR U60019 ( .A(n50487), .B(n50488), .Z(n50486) );
  NAND U60020 ( .A(n50487), .B(n50488), .Z(n50483) );
  XOR U60021 ( .A(n50487), .B(n50489), .Z(N60920) );
  XNOR U60022 ( .A(n50485), .B(n50488), .Z(n50489) );
  AND U60023 ( .A(n50490), .B(n50491), .Z(n50488) );
  NANDN U60024 ( .A(n50492), .B(n50493), .Z(n50491) );
  NANDN U60025 ( .A(n50494), .B(n50495), .Z(n50493) );
  NANDN U60026 ( .A(n50495), .B(n50494), .Z(n50490) );
  NAND U60027 ( .A(n50496), .B(n50497), .Z(n50485) );
  NANDN U60028 ( .A(n50498), .B(n50499), .Z(n50497) );
  OR U60029 ( .A(n50500), .B(n50501), .Z(n50499) );
  NAND U60030 ( .A(n50501), .B(n50500), .Z(n50496) );
  AND U60031 ( .A(n50502), .B(n50503), .Z(n50487) );
  NANDN U60032 ( .A(n50504), .B(n50505), .Z(n50503) );
  NANDN U60033 ( .A(n50506), .B(n50507), .Z(n50505) );
  NANDN U60034 ( .A(n50507), .B(n50506), .Z(n50502) );
  XOR U60035 ( .A(n50501), .B(n50508), .Z(N60919) );
  XOR U60036 ( .A(n50498), .B(n50500), .Z(n50508) );
  XNOR U60037 ( .A(n50494), .B(n50509), .Z(n50500) );
  XNOR U60038 ( .A(n50492), .B(n50495), .Z(n50509) );
  NAND U60039 ( .A(n50510), .B(n50511), .Z(n50495) );
  NAND U60040 ( .A(n50512), .B(n50513), .Z(n50511) );
  OR U60041 ( .A(n50514), .B(n50515), .Z(n50512) );
  NANDN U60042 ( .A(n50516), .B(n50514), .Z(n50510) );
  IV U60043 ( .A(n50515), .Z(n50516) );
  NAND U60044 ( .A(n50517), .B(n50518), .Z(n50492) );
  NAND U60045 ( .A(n50519), .B(n50520), .Z(n50518) );
  NANDN U60046 ( .A(n50521), .B(n50522), .Z(n50519) );
  NANDN U60047 ( .A(n50522), .B(n50521), .Z(n50517) );
  AND U60048 ( .A(n50523), .B(n50524), .Z(n50494) );
  NAND U60049 ( .A(n50525), .B(n50526), .Z(n50524) );
  OR U60050 ( .A(n50527), .B(n50528), .Z(n50525) );
  NANDN U60051 ( .A(n50529), .B(n50527), .Z(n50523) );
  NAND U60052 ( .A(n50530), .B(n50531), .Z(n50498) );
  NANDN U60053 ( .A(n50532), .B(n50533), .Z(n50531) );
  OR U60054 ( .A(n50534), .B(n50535), .Z(n50533) );
  NANDN U60055 ( .A(n50536), .B(n50534), .Z(n50530) );
  IV U60056 ( .A(n50535), .Z(n50536) );
  XNOR U60057 ( .A(n50506), .B(n50537), .Z(n50501) );
  XNOR U60058 ( .A(n50504), .B(n50507), .Z(n50537) );
  NAND U60059 ( .A(n50538), .B(n50539), .Z(n50507) );
  NAND U60060 ( .A(n50540), .B(n50541), .Z(n50539) );
  OR U60061 ( .A(n50542), .B(n50543), .Z(n50540) );
  NANDN U60062 ( .A(n50544), .B(n50542), .Z(n50538) );
  IV U60063 ( .A(n50543), .Z(n50544) );
  NAND U60064 ( .A(n50545), .B(n50546), .Z(n50504) );
  NAND U60065 ( .A(n50547), .B(n50548), .Z(n50546) );
  NANDN U60066 ( .A(n50549), .B(n50550), .Z(n50547) );
  NANDN U60067 ( .A(n50550), .B(n50549), .Z(n50545) );
  AND U60068 ( .A(n50551), .B(n50552), .Z(n50506) );
  NAND U60069 ( .A(n50553), .B(n50554), .Z(n50552) );
  OR U60070 ( .A(n50555), .B(n50556), .Z(n50553) );
  NANDN U60071 ( .A(n50557), .B(n50555), .Z(n50551) );
  XNOR U60072 ( .A(n50532), .B(n50558), .Z(N60918) );
  XOR U60073 ( .A(n50534), .B(n50535), .Z(n50558) );
  XNOR U60074 ( .A(n50548), .B(n50559), .Z(n50535) );
  XOR U60075 ( .A(n50549), .B(n50550), .Z(n50559) );
  XOR U60076 ( .A(n50555), .B(n50560), .Z(n50550) );
  XOR U60077 ( .A(n50554), .B(n50557), .Z(n50560) );
  IV U60078 ( .A(n50556), .Z(n50557) );
  NAND U60079 ( .A(n50561), .B(n50562), .Z(n50556) );
  OR U60080 ( .A(n50563), .B(n50564), .Z(n50562) );
  OR U60081 ( .A(n50565), .B(n50566), .Z(n50561) );
  NAND U60082 ( .A(n50567), .B(n50568), .Z(n50554) );
  OR U60083 ( .A(n50569), .B(n50570), .Z(n50568) );
  OR U60084 ( .A(n50571), .B(n50572), .Z(n50567) );
  NOR U60085 ( .A(n50573), .B(n50574), .Z(n50555) );
  ANDN U60086 ( .B(n50575), .A(n50576), .Z(n50549) );
  XNOR U60087 ( .A(n50542), .B(n50577), .Z(n50548) );
  XNOR U60088 ( .A(n50541), .B(n50543), .Z(n50577) );
  NAND U60089 ( .A(n50578), .B(n50579), .Z(n50543) );
  OR U60090 ( .A(n50580), .B(n50581), .Z(n50579) );
  OR U60091 ( .A(n50582), .B(n50583), .Z(n50578) );
  NAND U60092 ( .A(n50584), .B(n50585), .Z(n50541) );
  OR U60093 ( .A(n50586), .B(n50587), .Z(n50585) );
  OR U60094 ( .A(n50588), .B(n50589), .Z(n50584) );
  ANDN U60095 ( .B(n50590), .A(n50591), .Z(n50542) );
  IV U60096 ( .A(n50592), .Z(n50590) );
  ANDN U60097 ( .B(n50593), .A(n50594), .Z(n50534) );
  XOR U60098 ( .A(n50520), .B(n50595), .Z(n50532) );
  XOR U60099 ( .A(n50521), .B(n50522), .Z(n50595) );
  XOR U60100 ( .A(n50527), .B(n50596), .Z(n50522) );
  XOR U60101 ( .A(n50526), .B(n50529), .Z(n50596) );
  IV U60102 ( .A(n50528), .Z(n50529) );
  NAND U60103 ( .A(n50597), .B(n50598), .Z(n50528) );
  OR U60104 ( .A(n50599), .B(n50600), .Z(n50598) );
  OR U60105 ( .A(n50601), .B(n50602), .Z(n50597) );
  NAND U60106 ( .A(n50603), .B(n50604), .Z(n50526) );
  OR U60107 ( .A(n50605), .B(n50606), .Z(n50604) );
  OR U60108 ( .A(n50607), .B(n50608), .Z(n50603) );
  NOR U60109 ( .A(n50609), .B(n50610), .Z(n50527) );
  ANDN U60110 ( .B(n50611), .A(n50612), .Z(n50521) );
  IV U60111 ( .A(n50613), .Z(n50611) );
  XNOR U60112 ( .A(n50514), .B(n50614), .Z(n50520) );
  XNOR U60113 ( .A(n50513), .B(n50515), .Z(n50614) );
  NAND U60114 ( .A(n50615), .B(n50616), .Z(n50515) );
  OR U60115 ( .A(n50617), .B(n50618), .Z(n50616) );
  OR U60116 ( .A(n50619), .B(n50620), .Z(n50615) );
  NAND U60117 ( .A(n50621), .B(n50622), .Z(n50513) );
  OR U60118 ( .A(n50623), .B(n50624), .Z(n50622) );
  OR U60119 ( .A(n50625), .B(n50626), .Z(n50621) );
  ANDN U60120 ( .B(n50627), .A(n50628), .Z(n50514) );
  IV U60121 ( .A(n50629), .Z(n50627) );
  XNOR U60122 ( .A(n50594), .B(n50593), .Z(N60917) );
  XOR U60123 ( .A(n50613), .B(n50612), .Z(n50593) );
  XNOR U60124 ( .A(n50628), .B(n50629), .Z(n50612) );
  XNOR U60125 ( .A(n50623), .B(n50624), .Z(n50629) );
  XNOR U60126 ( .A(n50625), .B(n50626), .Z(n50624) );
  XNOR U60127 ( .A(y[613]), .B(x[613]), .Z(n50626) );
  XNOR U60128 ( .A(y[614]), .B(x[614]), .Z(n50625) );
  XNOR U60129 ( .A(y[612]), .B(x[612]), .Z(n50623) );
  XNOR U60130 ( .A(n50617), .B(n50618), .Z(n50628) );
  XNOR U60131 ( .A(y[609]), .B(x[609]), .Z(n50618) );
  XNOR U60132 ( .A(n50619), .B(n50620), .Z(n50617) );
  XNOR U60133 ( .A(y[610]), .B(x[610]), .Z(n50620) );
  XNOR U60134 ( .A(y[611]), .B(x[611]), .Z(n50619) );
  XNOR U60135 ( .A(n50610), .B(n50609), .Z(n50613) );
  XNOR U60136 ( .A(n50605), .B(n50606), .Z(n50609) );
  XNOR U60137 ( .A(y[606]), .B(x[606]), .Z(n50606) );
  XNOR U60138 ( .A(n50607), .B(n50608), .Z(n50605) );
  XNOR U60139 ( .A(y[607]), .B(x[607]), .Z(n50608) );
  XNOR U60140 ( .A(y[608]), .B(x[608]), .Z(n50607) );
  XNOR U60141 ( .A(n50599), .B(n50600), .Z(n50610) );
  XNOR U60142 ( .A(y[603]), .B(x[603]), .Z(n50600) );
  XNOR U60143 ( .A(n50601), .B(n50602), .Z(n50599) );
  XNOR U60144 ( .A(y[604]), .B(x[604]), .Z(n50602) );
  XNOR U60145 ( .A(y[605]), .B(x[605]), .Z(n50601) );
  XOR U60146 ( .A(n50575), .B(n50576), .Z(n50594) );
  XNOR U60147 ( .A(n50591), .B(n50592), .Z(n50576) );
  XNOR U60148 ( .A(n50586), .B(n50587), .Z(n50592) );
  XNOR U60149 ( .A(n50588), .B(n50589), .Z(n50587) );
  XNOR U60150 ( .A(y[601]), .B(x[601]), .Z(n50589) );
  XNOR U60151 ( .A(y[602]), .B(x[602]), .Z(n50588) );
  XNOR U60152 ( .A(y[600]), .B(x[600]), .Z(n50586) );
  XNOR U60153 ( .A(n50580), .B(n50581), .Z(n50591) );
  XNOR U60154 ( .A(y[597]), .B(x[597]), .Z(n50581) );
  XNOR U60155 ( .A(n50582), .B(n50583), .Z(n50580) );
  XNOR U60156 ( .A(y[598]), .B(x[598]), .Z(n50583) );
  XNOR U60157 ( .A(y[599]), .B(x[599]), .Z(n50582) );
  XOR U60158 ( .A(n50574), .B(n50573), .Z(n50575) );
  XNOR U60159 ( .A(n50569), .B(n50570), .Z(n50573) );
  XNOR U60160 ( .A(y[594]), .B(x[594]), .Z(n50570) );
  XNOR U60161 ( .A(n50571), .B(n50572), .Z(n50569) );
  XNOR U60162 ( .A(y[595]), .B(x[595]), .Z(n50572) );
  XNOR U60163 ( .A(y[596]), .B(x[596]), .Z(n50571) );
  XNOR U60164 ( .A(n50563), .B(n50564), .Z(n50574) );
  XNOR U60165 ( .A(y[591]), .B(x[591]), .Z(n50564) );
  XNOR U60166 ( .A(n50565), .B(n50566), .Z(n50563) );
  XNOR U60167 ( .A(y[592]), .B(x[592]), .Z(n50566) );
  XNOR U60168 ( .A(y[593]), .B(x[593]), .Z(n50565) );
  NAND U60169 ( .A(n50630), .B(n50631), .Z(N60908) );
  NANDN U60170 ( .A(n50632), .B(n50633), .Z(n50631) );
  OR U60171 ( .A(n50634), .B(n50635), .Z(n50633) );
  NAND U60172 ( .A(n50634), .B(n50635), .Z(n50630) );
  XOR U60173 ( .A(n50634), .B(n50636), .Z(N60907) );
  XNOR U60174 ( .A(n50632), .B(n50635), .Z(n50636) );
  AND U60175 ( .A(n50637), .B(n50638), .Z(n50635) );
  NANDN U60176 ( .A(n50639), .B(n50640), .Z(n50638) );
  NANDN U60177 ( .A(n50641), .B(n50642), .Z(n50640) );
  NANDN U60178 ( .A(n50642), .B(n50641), .Z(n50637) );
  NAND U60179 ( .A(n50643), .B(n50644), .Z(n50632) );
  NANDN U60180 ( .A(n50645), .B(n50646), .Z(n50644) );
  OR U60181 ( .A(n50647), .B(n50648), .Z(n50646) );
  NAND U60182 ( .A(n50648), .B(n50647), .Z(n50643) );
  AND U60183 ( .A(n50649), .B(n50650), .Z(n50634) );
  NANDN U60184 ( .A(n50651), .B(n50652), .Z(n50650) );
  NANDN U60185 ( .A(n50653), .B(n50654), .Z(n50652) );
  NANDN U60186 ( .A(n50654), .B(n50653), .Z(n50649) );
  XOR U60187 ( .A(n50648), .B(n50655), .Z(N60906) );
  XOR U60188 ( .A(n50645), .B(n50647), .Z(n50655) );
  XNOR U60189 ( .A(n50641), .B(n50656), .Z(n50647) );
  XNOR U60190 ( .A(n50639), .B(n50642), .Z(n50656) );
  NAND U60191 ( .A(n50657), .B(n50658), .Z(n50642) );
  NAND U60192 ( .A(n50659), .B(n50660), .Z(n50658) );
  OR U60193 ( .A(n50661), .B(n50662), .Z(n50659) );
  NANDN U60194 ( .A(n50663), .B(n50661), .Z(n50657) );
  IV U60195 ( .A(n50662), .Z(n50663) );
  NAND U60196 ( .A(n50664), .B(n50665), .Z(n50639) );
  NAND U60197 ( .A(n50666), .B(n50667), .Z(n50665) );
  NANDN U60198 ( .A(n50668), .B(n50669), .Z(n50666) );
  NANDN U60199 ( .A(n50669), .B(n50668), .Z(n50664) );
  AND U60200 ( .A(n50670), .B(n50671), .Z(n50641) );
  NAND U60201 ( .A(n50672), .B(n50673), .Z(n50671) );
  OR U60202 ( .A(n50674), .B(n50675), .Z(n50672) );
  NANDN U60203 ( .A(n50676), .B(n50674), .Z(n50670) );
  NAND U60204 ( .A(n50677), .B(n50678), .Z(n50645) );
  NANDN U60205 ( .A(n50679), .B(n50680), .Z(n50678) );
  OR U60206 ( .A(n50681), .B(n50682), .Z(n50680) );
  NANDN U60207 ( .A(n50683), .B(n50681), .Z(n50677) );
  IV U60208 ( .A(n50682), .Z(n50683) );
  XNOR U60209 ( .A(n50653), .B(n50684), .Z(n50648) );
  XNOR U60210 ( .A(n50651), .B(n50654), .Z(n50684) );
  NAND U60211 ( .A(n50685), .B(n50686), .Z(n50654) );
  NAND U60212 ( .A(n50687), .B(n50688), .Z(n50686) );
  OR U60213 ( .A(n50689), .B(n50690), .Z(n50687) );
  NANDN U60214 ( .A(n50691), .B(n50689), .Z(n50685) );
  IV U60215 ( .A(n50690), .Z(n50691) );
  NAND U60216 ( .A(n50692), .B(n50693), .Z(n50651) );
  NAND U60217 ( .A(n50694), .B(n50695), .Z(n50693) );
  NANDN U60218 ( .A(n50696), .B(n50697), .Z(n50694) );
  NANDN U60219 ( .A(n50697), .B(n50696), .Z(n50692) );
  AND U60220 ( .A(n50698), .B(n50699), .Z(n50653) );
  NAND U60221 ( .A(n50700), .B(n50701), .Z(n50699) );
  OR U60222 ( .A(n50702), .B(n50703), .Z(n50700) );
  NANDN U60223 ( .A(n50704), .B(n50702), .Z(n50698) );
  XNOR U60224 ( .A(n50679), .B(n50705), .Z(N60905) );
  XOR U60225 ( .A(n50681), .B(n50682), .Z(n50705) );
  XNOR U60226 ( .A(n50695), .B(n50706), .Z(n50682) );
  XOR U60227 ( .A(n50696), .B(n50697), .Z(n50706) );
  XOR U60228 ( .A(n50702), .B(n50707), .Z(n50697) );
  XOR U60229 ( .A(n50701), .B(n50704), .Z(n50707) );
  IV U60230 ( .A(n50703), .Z(n50704) );
  NAND U60231 ( .A(n50708), .B(n50709), .Z(n50703) );
  OR U60232 ( .A(n50710), .B(n50711), .Z(n50709) );
  OR U60233 ( .A(n50712), .B(n50713), .Z(n50708) );
  NAND U60234 ( .A(n50714), .B(n50715), .Z(n50701) );
  OR U60235 ( .A(n50716), .B(n50717), .Z(n50715) );
  OR U60236 ( .A(n50718), .B(n50719), .Z(n50714) );
  NOR U60237 ( .A(n50720), .B(n50721), .Z(n50702) );
  ANDN U60238 ( .B(n50722), .A(n50723), .Z(n50696) );
  XNOR U60239 ( .A(n50689), .B(n50724), .Z(n50695) );
  XNOR U60240 ( .A(n50688), .B(n50690), .Z(n50724) );
  NAND U60241 ( .A(n50725), .B(n50726), .Z(n50690) );
  OR U60242 ( .A(n50727), .B(n50728), .Z(n50726) );
  OR U60243 ( .A(n50729), .B(n50730), .Z(n50725) );
  NAND U60244 ( .A(n50731), .B(n50732), .Z(n50688) );
  OR U60245 ( .A(n50733), .B(n50734), .Z(n50732) );
  OR U60246 ( .A(n50735), .B(n50736), .Z(n50731) );
  ANDN U60247 ( .B(n50737), .A(n50738), .Z(n50689) );
  IV U60248 ( .A(n50739), .Z(n50737) );
  ANDN U60249 ( .B(n50740), .A(n50741), .Z(n50681) );
  XOR U60250 ( .A(n50667), .B(n50742), .Z(n50679) );
  XOR U60251 ( .A(n50668), .B(n50669), .Z(n50742) );
  XOR U60252 ( .A(n50674), .B(n50743), .Z(n50669) );
  XOR U60253 ( .A(n50673), .B(n50676), .Z(n50743) );
  IV U60254 ( .A(n50675), .Z(n50676) );
  NAND U60255 ( .A(n50744), .B(n50745), .Z(n50675) );
  OR U60256 ( .A(n50746), .B(n50747), .Z(n50745) );
  OR U60257 ( .A(n50748), .B(n50749), .Z(n50744) );
  NAND U60258 ( .A(n50750), .B(n50751), .Z(n50673) );
  OR U60259 ( .A(n50752), .B(n50753), .Z(n50751) );
  OR U60260 ( .A(n50754), .B(n50755), .Z(n50750) );
  NOR U60261 ( .A(n50756), .B(n50757), .Z(n50674) );
  ANDN U60262 ( .B(n50758), .A(n50759), .Z(n50668) );
  IV U60263 ( .A(n50760), .Z(n50758) );
  XNOR U60264 ( .A(n50661), .B(n50761), .Z(n50667) );
  XNOR U60265 ( .A(n50660), .B(n50662), .Z(n50761) );
  NAND U60266 ( .A(n50762), .B(n50763), .Z(n50662) );
  OR U60267 ( .A(n50764), .B(n50765), .Z(n50763) );
  OR U60268 ( .A(n50766), .B(n50767), .Z(n50762) );
  NAND U60269 ( .A(n50768), .B(n50769), .Z(n50660) );
  OR U60270 ( .A(n50770), .B(n50771), .Z(n50769) );
  OR U60271 ( .A(n50772), .B(n50773), .Z(n50768) );
  ANDN U60272 ( .B(n50774), .A(n50775), .Z(n50661) );
  IV U60273 ( .A(n50776), .Z(n50774) );
  XNOR U60274 ( .A(n50741), .B(n50740), .Z(N60904) );
  XOR U60275 ( .A(n50760), .B(n50759), .Z(n50740) );
  XNOR U60276 ( .A(n50775), .B(n50776), .Z(n50759) );
  XNOR U60277 ( .A(n50770), .B(n50771), .Z(n50776) );
  XNOR U60278 ( .A(n50772), .B(n50773), .Z(n50771) );
  XNOR U60279 ( .A(y[589]), .B(x[589]), .Z(n50773) );
  XNOR U60280 ( .A(y[590]), .B(x[590]), .Z(n50772) );
  XNOR U60281 ( .A(y[588]), .B(x[588]), .Z(n50770) );
  XNOR U60282 ( .A(n50764), .B(n50765), .Z(n50775) );
  XNOR U60283 ( .A(y[585]), .B(x[585]), .Z(n50765) );
  XNOR U60284 ( .A(n50766), .B(n50767), .Z(n50764) );
  XNOR U60285 ( .A(y[586]), .B(x[586]), .Z(n50767) );
  XNOR U60286 ( .A(y[587]), .B(x[587]), .Z(n50766) );
  XNOR U60287 ( .A(n50757), .B(n50756), .Z(n50760) );
  XNOR U60288 ( .A(n50752), .B(n50753), .Z(n50756) );
  XNOR U60289 ( .A(y[582]), .B(x[582]), .Z(n50753) );
  XNOR U60290 ( .A(n50754), .B(n50755), .Z(n50752) );
  XNOR U60291 ( .A(y[583]), .B(x[583]), .Z(n50755) );
  XNOR U60292 ( .A(y[584]), .B(x[584]), .Z(n50754) );
  XNOR U60293 ( .A(n50746), .B(n50747), .Z(n50757) );
  XNOR U60294 ( .A(y[579]), .B(x[579]), .Z(n50747) );
  XNOR U60295 ( .A(n50748), .B(n50749), .Z(n50746) );
  XNOR U60296 ( .A(y[580]), .B(x[580]), .Z(n50749) );
  XNOR U60297 ( .A(y[581]), .B(x[581]), .Z(n50748) );
  XOR U60298 ( .A(n50722), .B(n50723), .Z(n50741) );
  XNOR U60299 ( .A(n50738), .B(n50739), .Z(n50723) );
  XNOR U60300 ( .A(n50733), .B(n50734), .Z(n50739) );
  XNOR U60301 ( .A(n50735), .B(n50736), .Z(n50734) );
  XNOR U60302 ( .A(y[577]), .B(x[577]), .Z(n50736) );
  XNOR U60303 ( .A(y[578]), .B(x[578]), .Z(n50735) );
  XNOR U60304 ( .A(y[576]), .B(x[576]), .Z(n50733) );
  XNOR U60305 ( .A(n50727), .B(n50728), .Z(n50738) );
  XNOR U60306 ( .A(y[573]), .B(x[573]), .Z(n50728) );
  XNOR U60307 ( .A(n50729), .B(n50730), .Z(n50727) );
  XNOR U60308 ( .A(y[574]), .B(x[574]), .Z(n50730) );
  XNOR U60309 ( .A(y[575]), .B(x[575]), .Z(n50729) );
  XOR U60310 ( .A(n50721), .B(n50720), .Z(n50722) );
  XNOR U60311 ( .A(n50716), .B(n50717), .Z(n50720) );
  XNOR U60312 ( .A(y[570]), .B(x[570]), .Z(n50717) );
  XNOR U60313 ( .A(n50718), .B(n50719), .Z(n50716) );
  XNOR U60314 ( .A(y[571]), .B(x[571]), .Z(n50719) );
  XNOR U60315 ( .A(y[572]), .B(x[572]), .Z(n50718) );
  XNOR U60316 ( .A(n50710), .B(n50711), .Z(n50721) );
  XNOR U60317 ( .A(y[567]), .B(x[567]), .Z(n50711) );
  XNOR U60318 ( .A(n50712), .B(n50713), .Z(n50710) );
  XNOR U60319 ( .A(y[568]), .B(x[568]), .Z(n50713) );
  XNOR U60320 ( .A(y[569]), .B(x[569]), .Z(n50712) );
  NAND U60321 ( .A(n50777), .B(n50778), .Z(N60895) );
  NANDN U60322 ( .A(n50779), .B(n50780), .Z(n50778) );
  OR U60323 ( .A(n50781), .B(n50782), .Z(n50780) );
  NAND U60324 ( .A(n50781), .B(n50782), .Z(n50777) );
  XOR U60325 ( .A(n50781), .B(n50783), .Z(N60894) );
  XNOR U60326 ( .A(n50779), .B(n50782), .Z(n50783) );
  AND U60327 ( .A(n50784), .B(n50785), .Z(n50782) );
  NANDN U60328 ( .A(n50786), .B(n50787), .Z(n50785) );
  NANDN U60329 ( .A(n50788), .B(n50789), .Z(n50787) );
  NANDN U60330 ( .A(n50789), .B(n50788), .Z(n50784) );
  NAND U60331 ( .A(n50790), .B(n50791), .Z(n50779) );
  NANDN U60332 ( .A(n50792), .B(n50793), .Z(n50791) );
  OR U60333 ( .A(n50794), .B(n50795), .Z(n50793) );
  NAND U60334 ( .A(n50795), .B(n50794), .Z(n50790) );
  AND U60335 ( .A(n50796), .B(n50797), .Z(n50781) );
  NANDN U60336 ( .A(n50798), .B(n50799), .Z(n50797) );
  NANDN U60337 ( .A(n50800), .B(n50801), .Z(n50799) );
  NANDN U60338 ( .A(n50801), .B(n50800), .Z(n50796) );
  XOR U60339 ( .A(n50795), .B(n50802), .Z(N60893) );
  XOR U60340 ( .A(n50792), .B(n50794), .Z(n50802) );
  XNOR U60341 ( .A(n50788), .B(n50803), .Z(n50794) );
  XNOR U60342 ( .A(n50786), .B(n50789), .Z(n50803) );
  NAND U60343 ( .A(n50804), .B(n50805), .Z(n50789) );
  NAND U60344 ( .A(n50806), .B(n50807), .Z(n50805) );
  OR U60345 ( .A(n50808), .B(n50809), .Z(n50806) );
  NANDN U60346 ( .A(n50810), .B(n50808), .Z(n50804) );
  IV U60347 ( .A(n50809), .Z(n50810) );
  NAND U60348 ( .A(n50811), .B(n50812), .Z(n50786) );
  NAND U60349 ( .A(n50813), .B(n50814), .Z(n50812) );
  NANDN U60350 ( .A(n50815), .B(n50816), .Z(n50813) );
  NANDN U60351 ( .A(n50816), .B(n50815), .Z(n50811) );
  AND U60352 ( .A(n50817), .B(n50818), .Z(n50788) );
  NAND U60353 ( .A(n50819), .B(n50820), .Z(n50818) );
  OR U60354 ( .A(n50821), .B(n50822), .Z(n50819) );
  NANDN U60355 ( .A(n50823), .B(n50821), .Z(n50817) );
  NAND U60356 ( .A(n50824), .B(n50825), .Z(n50792) );
  NANDN U60357 ( .A(n50826), .B(n50827), .Z(n50825) );
  OR U60358 ( .A(n50828), .B(n50829), .Z(n50827) );
  NANDN U60359 ( .A(n50830), .B(n50828), .Z(n50824) );
  IV U60360 ( .A(n50829), .Z(n50830) );
  XNOR U60361 ( .A(n50800), .B(n50831), .Z(n50795) );
  XNOR U60362 ( .A(n50798), .B(n50801), .Z(n50831) );
  NAND U60363 ( .A(n50832), .B(n50833), .Z(n50801) );
  NAND U60364 ( .A(n50834), .B(n50835), .Z(n50833) );
  OR U60365 ( .A(n50836), .B(n50837), .Z(n50834) );
  NANDN U60366 ( .A(n50838), .B(n50836), .Z(n50832) );
  IV U60367 ( .A(n50837), .Z(n50838) );
  NAND U60368 ( .A(n50839), .B(n50840), .Z(n50798) );
  NAND U60369 ( .A(n50841), .B(n50842), .Z(n50840) );
  NANDN U60370 ( .A(n50843), .B(n50844), .Z(n50841) );
  NANDN U60371 ( .A(n50844), .B(n50843), .Z(n50839) );
  AND U60372 ( .A(n50845), .B(n50846), .Z(n50800) );
  NAND U60373 ( .A(n50847), .B(n50848), .Z(n50846) );
  OR U60374 ( .A(n50849), .B(n50850), .Z(n50847) );
  NANDN U60375 ( .A(n50851), .B(n50849), .Z(n50845) );
  XNOR U60376 ( .A(n50826), .B(n50852), .Z(N60892) );
  XOR U60377 ( .A(n50828), .B(n50829), .Z(n50852) );
  XNOR U60378 ( .A(n50842), .B(n50853), .Z(n50829) );
  XOR U60379 ( .A(n50843), .B(n50844), .Z(n50853) );
  XOR U60380 ( .A(n50849), .B(n50854), .Z(n50844) );
  XOR U60381 ( .A(n50848), .B(n50851), .Z(n50854) );
  IV U60382 ( .A(n50850), .Z(n50851) );
  NAND U60383 ( .A(n50855), .B(n50856), .Z(n50850) );
  OR U60384 ( .A(n50857), .B(n50858), .Z(n50856) );
  OR U60385 ( .A(n50859), .B(n50860), .Z(n50855) );
  NAND U60386 ( .A(n50861), .B(n50862), .Z(n50848) );
  OR U60387 ( .A(n50863), .B(n50864), .Z(n50862) );
  OR U60388 ( .A(n50865), .B(n50866), .Z(n50861) );
  NOR U60389 ( .A(n50867), .B(n50868), .Z(n50849) );
  ANDN U60390 ( .B(n50869), .A(n50870), .Z(n50843) );
  XNOR U60391 ( .A(n50836), .B(n50871), .Z(n50842) );
  XNOR U60392 ( .A(n50835), .B(n50837), .Z(n50871) );
  NAND U60393 ( .A(n50872), .B(n50873), .Z(n50837) );
  OR U60394 ( .A(n50874), .B(n50875), .Z(n50873) );
  OR U60395 ( .A(n50876), .B(n50877), .Z(n50872) );
  NAND U60396 ( .A(n50878), .B(n50879), .Z(n50835) );
  OR U60397 ( .A(n50880), .B(n50881), .Z(n50879) );
  OR U60398 ( .A(n50882), .B(n50883), .Z(n50878) );
  ANDN U60399 ( .B(n50884), .A(n50885), .Z(n50836) );
  IV U60400 ( .A(n50886), .Z(n50884) );
  ANDN U60401 ( .B(n50887), .A(n50888), .Z(n50828) );
  XOR U60402 ( .A(n50814), .B(n50889), .Z(n50826) );
  XOR U60403 ( .A(n50815), .B(n50816), .Z(n50889) );
  XOR U60404 ( .A(n50821), .B(n50890), .Z(n50816) );
  XOR U60405 ( .A(n50820), .B(n50823), .Z(n50890) );
  IV U60406 ( .A(n50822), .Z(n50823) );
  NAND U60407 ( .A(n50891), .B(n50892), .Z(n50822) );
  OR U60408 ( .A(n50893), .B(n50894), .Z(n50892) );
  OR U60409 ( .A(n50895), .B(n50896), .Z(n50891) );
  NAND U60410 ( .A(n50897), .B(n50898), .Z(n50820) );
  OR U60411 ( .A(n50899), .B(n50900), .Z(n50898) );
  OR U60412 ( .A(n50901), .B(n50902), .Z(n50897) );
  NOR U60413 ( .A(n50903), .B(n50904), .Z(n50821) );
  ANDN U60414 ( .B(n50905), .A(n50906), .Z(n50815) );
  IV U60415 ( .A(n50907), .Z(n50905) );
  XNOR U60416 ( .A(n50808), .B(n50908), .Z(n50814) );
  XNOR U60417 ( .A(n50807), .B(n50809), .Z(n50908) );
  NAND U60418 ( .A(n50909), .B(n50910), .Z(n50809) );
  OR U60419 ( .A(n50911), .B(n50912), .Z(n50910) );
  OR U60420 ( .A(n50913), .B(n50914), .Z(n50909) );
  NAND U60421 ( .A(n50915), .B(n50916), .Z(n50807) );
  OR U60422 ( .A(n50917), .B(n50918), .Z(n50916) );
  OR U60423 ( .A(n50919), .B(n50920), .Z(n50915) );
  ANDN U60424 ( .B(n50921), .A(n50922), .Z(n50808) );
  IV U60425 ( .A(n50923), .Z(n50921) );
  XNOR U60426 ( .A(n50888), .B(n50887), .Z(N60891) );
  XOR U60427 ( .A(n50907), .B(n50906), .Z(n50887) );
  XNOR U60428 ( .A(n50922), .B(n50923), .Z(n50906) );
  XNOR U60429 ( .A(n50917), .B(n50918), .Z(n50923) );
  XNOR U60430 ( .A(n50919), .B(n50920), .Z(n50918) );
  XNOR U60431 ( .A(y[565]), .B(x[565]), .Z(n50920) );
  XNOR U60432 ( .A(y[566]), .B(x[566]), .Z(n50919) );
  XNOR U60433 ( .A(y[564]), .B(x[564]), .Z(n50917) );
  XNOR U60434 ( .A(n50911), .B(n50912), .Z(n50922) );
  XNOR U60435 ( .A(y[561]), .B(x[561]), .Z(n50912) );
  XNOR U60436 ( .A(n50913), .B(n50914), .Z(n50911) );
  XNOR U60437 ( .A(y[562]), .B(x[562]), .Z(n50914) );
  XNOR U60438 ( .A(y[563]), .B(x[563]), .Z(n50913) );
  XNOR U60439 ( .A(n50904), .B(n50903), .Z(n50907) );
  XNOR U60440 ( .A(n50899), .B(n50900), .Z(n50903) );
  XNOR U60441 ( .A(y[558]), .B(x[558]), .Z(n50900) );
  XNOR U60442 ( .A(n50901), .B(n50902), .Z(n50899) );
  XNOR U60443 ( .A(y[559]), .B(x[559]), .Z(n50902) );
  XNOR U60444 ( .A(y[560]), .B(x[560]), .Z(n50901) );
  XNOR U60445 ( .A(n50893), .B(n50894), .Z(n50904) );
  XNOR U60446 ( .A(y[555]), .B(x[555]), .Z(n50894) );
  XNOR U60447 ( .A(n50895), .B(n50896), .Z(n50893) );
  XNOR U60448 ( .A(y[556]), .B(x[556]), .Z(n50896) );
  XNOR U60449 ( .A(y[557]), .B(x[557]), .Z(n50895) );
  XOR U60450 ( .A(n50869), .B(n50870), .Z(n50888) );
  XNOR U60451 ( .A(n50885), .B(n50886), .Z(n50870) );
  XNOR U60452 ( .A(n50880), .B(n50881), .Z(n50886) );
  XNOR U60453 ( .A(n50882), .B(n50883), .Z(n50881) );
  XNOR U60454 ( .A(y[553]), .B(x[553]), .Z(n50883) );
  XNOR U60455 ( .A(y[554]), .B(x[554]), .Z(n50882) );
  XNOR U60456 ( .A(y[552]), .B(x[552]), .Z(n50880) );
  XNOR U60457 ( .A(n50874), .B(n50875), .Z(n50885) );
  XNOR U60458 ( .A(y[549]), .B(x[549]), .Z(n50875) );
  XNOR U60459 ( .A(n50876), .B(n50877), .Z(n50874) );
  XNOR U60460 ( .A(y[550]), .B(x[550]), .Z(n50877) );
  XNOR U60461 ( .A(y[551]), .B(x[551]), .Z(n50876) );
  XOR U60462 ( .A(n50868), .B(n50867), .Z(n50869) );
  XNOR U60463 ( .A(n50863), .B(n50864), .Z(n50867) );
  XNOR U60464 ( .A(y[546]), .B(x[546]), .Z(n50864) );
  XNOR U60465 ( .A(n50865), .B(n50866), .Z(n50863) );
  XNOR U60466 ( .A(y[547]), .B(x[547]), .Z(n50866) );
  XNOR U60467 ( .A(y[548]), .B(x[548]), .Z(n50865) );
  XNOR U60468 ( .A(n50857), .B(n50858), .Z(n50868) );
  XNOR U60469 ( .A(y[543]), .B(x[543]), .Z(n50858) );
  XNOR U60470 ( .A(n50859), .B(n50860), .Z(n50857) );
  XNOR U60471 ( .A(y[544]), .B(x[544]), .Z(n50860) );
  XNOR U60472 ( .A(y[545]), .B(x[545]), .Z(n50859) );
  NAND U60473 ( .A(n50924), .B(n50925), .Z(N60882) );
  NANDN U60474 ( .A(n50926), .B(n50927), .Z(n50925) );
  OR U60475 ( .A(n50928), .B(n50929), .Z(n50927) );
  NAND U60476 ( .A(n50928), .B(n50929), .Z(n50924) );
  XOR U60477 ( .A(n50928), .B(n50930), .Z(N60881) );
  XNOR U60478 ( .A(n50926), .B(n50929), .Z(n50930) );
  AND U60479 ( .A(n50931), .B(n50932), .Z(n50929) );
  NANDN U60480 ( .A(n50933), .B(n50934), .Z(n50932) );
  NANDN U60481 ( .A(n50935), .B(n50936), .Z(n50934) );
  NANDN U60482 ( .A(n50936), .B(n50935), .Z(n50931) );
  NAND U60483 ( .A(n50937), .B(n50938), .Z(n50926) );
  NANDN U60484 ( .A(n50939), .B(n50940), .Z(n50938) );
  OR U60485 ( .A(n50941), .B(n50942), .Z(n50940) );
  NAND U60486 ( .A(n50942), .B(n50941), .Z(n50937) );
  AND U60487 ( .A(n50943), .B(n50944), .Z(n50928) );
  NANDN U60488 ( .A(n50945), .B(n50946), .Z(n50944) );
  NANDN U60489 ( .A(n50947), .B(n50948), .Z(n50946) );
  NANDN U60490 ( .A(n50948), .B(n50947), .Z(n50943) );
  XOR U60491 ( .A(n50942), .B(n50949), .Z(N60880) );
  XOR U60492 ( .A(n50939), .B(n50941), .Z(n50949) );
  XNOR U60493 ( .A(n50935), .B(n50950), .Z(n50941) );
  XNOR U60494 ( .A(n50933), .B(n50936), .Z(n50950) );
  NAND U60495 ( .A(n50951), .B(n50952), .Z(n50936) );
  NAND U60496 ( .A(n50953), .B(n50954), .Z(n50952) );
  OR U60497 ( .A(n50955), .B(n50956), .Z(n50953) );
  NANDN U60498 ( .A(n50957), .B(n50955), .Z(n50951) );
  IV U60499 ( .A(n50956), .Z(n50957) );
  NAND U60500 ( .A(n50958), .B(n50959), .Z(n50933) );
  NAND U60501 ( .A(n50960), .B(n50961), .Z(n50959) );
  NANDN U60502 ( .A(n50962), .B(n50963), .Z(n50960) );
  NANDN U60503 ( .A(n50963), .B(n50962), .Z(n50958) );
  AND U60504 ( .A(n50964), .B(n50965), .Z(n50935) );
  NAND U60505 ( .A(n50966), .B(n50967), .Z(n50965) );
  OR U60506 ( .A(n50968), .B(n50969), .Z(n50966) );
  NANDN U60507 ( .A(n50970), .B(n50968), .Z(n50964) );
  NAND U60508 ( .A(n50971), .B(n50972), .Z(n50939) );
  NANDN U60509 ( .A(n50973), .B(n50974), .Z(n50972) );
  OR U60510 ( .A(n50975), .B(n50976), .Z(n50974) );
  NANDN U60511 ( .A(n50977), .B(n50975), .Z(n50971) );
  IV U60512 ( .A(n50976), .Z(n50977) );
  XNOR U60513 ( .A(n50947), .B(n50978), .Z(n50942) );
  XNOR U60514 ( .A(n50945), .B(n50948), .Z(n50978) );
  NAND U60515 ( .A(n50979), .B(n50980), .Z(n50948) );
  NAND U60516 ( .A(n50981), .B(n50982), .Z(n50980) );
  OR U60517 ( .A(n50983), .B(n50984), .Z(n50981) );
  NANDN U60518 ( .A(n50985), .B(n50983), .Z(n50979) );
  IV U60519 ( .A(n50984), .Z(n50985) );
  NAND U60520 ( .A(n50986), .B(n50987), .Z(n50945) );
  NAND U60521 ( .A(n50988), .B(n50989), .Z(n50987) );
  NANDN U60522 ( .A(n50990), .B(n50991), .Z(n50988) );
  NANDN U60523 ( .A(n50991), .B(n50990), .Z(n50986) );
  AND U60524 ( .A(n50992), .B(n50993), .Z(n50947) );
  NAND U60525 ( .A(n50994), .B(n50995), .Z(n50993) );
  OR U60526 ( .A(n50996), .B(n50997), .Z(n50994) );
  NANDN U60527 ( .A(n50998), .B(n50996), .Z(n50992) );
  XNOR U60528 ( .A(n50973), .B(n50999), .Z(N60879) );
  XOR U60529 ( .A(n50975), .B(n50976), .Z(n50999) );
  XNOR U60530 ( .A(n50989), .B(n51000), .Z(n50976) );
  XOR U60531 ( .A(n50990), .B(n50991), .Z(n51000) );
  XOR U60532 ( .A(n50996), .B(n51001), .Z(n50991) );
  XOR U60533 ( .A(n50995), .B(n50998), .Z(n51001) );
  IV U60534 ( .A(n50997), .Z(n50998) );
  NAND U60535 ( .A(n51002), .B(n51003), .Z(n50997) );
  OR U60536 ( .A(n51004), .B(n51005), .Z(n51003) );
  OR U60537 ( .A(n51006), .B(n51007), .Z(n51002) );
  NAND U60538 ( .A(n51008), .B(n51009), .Z(n50995) );
  OR U60539 ( .A(n51010), .B(n51011), .Z(n51009) );
  OR U60540 ( .A(n51012), .B(n51013), .Z(n51008) );
  NOR U60541 ( .A(n51014), .B(n51015), .Z(n50996) );
  ANDN U60542 ( .B(n51016), .A(n51017), .Z(n50990) );
  XNOR U60543 ( .A(n50983), .B(n51018), .Z(n50989) );
  XNOR U60544 ( .A(n50982), .B(n50984), .Z(n51018) );
  NAND U60545 ( .A(n51019), .B(n51020), .Z(n50984) );
  OR U60546 ( .A(n51021), .B(n51022), .Z(n51020) );
  OR U60547 ( .A(n51023), .B(n51024), .Z(n51019) );
  NAND U60548 ( .A(n51025), .B(n51026), .Z(n50982) );
  OR U60549 ( .A(n51027), .B(n51028), .Z(n51026) );
  OR U60550 ( .A(n51029), .B(n51030), .Z(n51025) );
  ANDN U60551 ( .B(n51031), .A(n51032), .Z(n50983) );
  IV U60552 ( .A(n51033), .Z(n51031) );
  ANDN U60553 ( .B(n51034), .A(n51035), .Z(n50975) );
  XOR U60554 ( .A(n50961), .B(n51036), .Z(n50973) );
  XOR U60555 ( .A(n50962), .B(n50963), .Z(n51036) );
  XOR U60556 ( .A(n50968), .B(n51037), .Z(n50963) );
  XOR U60557 ( .A(n50967), .B(n50970), .Z(n51037) );
  IV U60558 ( .A(n50969), .Z(n50970) );
  NAND U60559 ( .A(n51038), .B(n51039), .Z(n50969) );
  OR U60560 ( .A(n51040), .B(n51041), .Z(n51039) );
  OR U60561 ( .A(n51042), .B(n51043), .Z(n51038) );
  NAND U60562 ( .A(n51044), .B(n51045), .Z(n50967) );
  OR U60563 ( .A(n51046), .B(n51047), .Z(n51045) );
  OR U60564 ( .A(n51048), .B(n51049), .Z(n51044) );
  NOR U60565 ( .A(n51050), .B(n51051), .Z(n50968) );
  ANDN U60566 ( .B(n51052), .A(n51053), .Z(n50962) );
  IV U60567 ( .A(n51054), .Z(n51052) );
  XNOR U60568 ( .A(n50955), .B(n51055), .Z(n50961) );
  XNOR U60569 ( .A(n50954), .B(n50956), .Z(n51055) );
  NAND U60570 ( .A(n51056), .B(n51057), .Z(n50956) );
  OR U60571 ( .A(n51058), .B(n51059), .Z(n51057) );
  OR U60572 ( .A(n51060), .B(n51061), .Z(n51056) );
  NAND U60573 ( .A(n51062), .B(n51063), .Z(n50954) );
  OR U60574 ( .A(n51064), .B(n51065), .Z(n51063) );
  OR U60575 ( .A(n51066), .B(n51067), .Z(n51062) );
  ANDN U60576 ( .B(n51068), .A(n51069), .Z(n50955) );
  IV U60577 ( .A(n51070), .Z(n51068) );
  XNOR U60578 ( .A(n51035), .B(n51034), .Z(N60878) );
  XOR U60579 ( .A(n51054), .B(n51053), .Z(n51034) );
  XNOR U60580 ( .A(n51069), .B(n51070), .Z(n51053) );
  XNOR U60581 ( .A(n51064), .B(n51065), .Z(n51070) );
  XNOR U60582 ( .A(n51066), .B(n51067), .Z(n51065) );
  XNOR U60583 ( .A(y[541]), .B(x[541]), .Z(n51067) );
  XNOR U60584 ( .A(y[542]), .B(x[542]), .Z(n51066) );
  XNOR U60585 ( .A(y[540]), .B(x[540]), .Z(n51064) );
  XNOR U60586 ( .A(n51058), .B(n51059), .Z(n51069) );
  XNOR U60587 ( .A(y[537]), .B(x[537]), .Z(n51059) );
  XNOR U60588 ( .A(n51060), .B(n51061), .Z(n51058) );
  XNOR U60589 ( .A(y[538]), .B(x[538]), .Z(n51061) );
  XNOR U60590 ( .A(y[539]), .B(x[539]), .Z(n51060) );
  XNOR U60591 ( .A(n51051), .B(n51050), .Z(n51054) );
  XNOR U60592 ( .A(n51046), .B(n51047), .Z(n51050) );
  XNOR U60593 ( .A(y[534]), .B(x[534]), .Z(n51047) );
  XNOR U60594 ( .A(n51048), .B(n51049), .Z(n51046) );
  XNOR U60595 ( .A(y[535]), .B(x[535]), .Z(n51049) );
  XNOR U60596 ( .A(y[536]), .B(x[536]), .Z(n51048) );
  XNOR U60597 ( .A(n51040), .B(n51041), .Z(n51051) );
  XNOR U60598 ( .A(y[531]), .B(x[531]), .Z(n51041) );
  XNOR U60599 ( .A(n51042), .B(n51043), .Z(n51040) );
  XNOR U60600 ( .A(y[532]), .B(x[532]), .Z(n51043) );
  XNOR U60601 ( .A(y[533]), .B(x[533]), .Z(n51042) );
  XOR U60602 ( .A(n51016), .B(n51017), .Z(n51035) );
  XNOR U60603 ( .A(n51032), .B(n51033), .Z(n51017) );
  XNOR U60604 ( .A(n51027), .B(n51028), .Z(n51033) );
  XNOR U60605 ( .A(n51029), .B(n51030), .Z(n51028) );
  XNOR U60606 ( .A(y[529]), .B(x[529]), .Z(n51030) );
  XNOR U60607 ( .A(y[530]), .B(x[530]), .Z(n51029) );
  XNOR U60608 ( .A(y[528]), .B(x[528]), .Z(n51027) );
  XNOR U60609 ( .A(n51021), .B(n51022), .Z(n51032) );
  XNOR U60610 ( .A(y[525]), .B(x[525]), .Z(n51022) );
  XNOR U60611 ( .A(n51023), .B(n51024), .Z(n51021) );
  XNOR U60612 ( .A(y[526]), .B(x[526]), .Z(n51024) );
  XNOR U60613 ( .A(y[527]), .B(x[527]), .Z(n51023) );
  XOR U60614 ( .A(n51015), .B(n51014), .Z(n51016) );
  XNOR U60615 ( .A(n51010), .B(n51011), .Z(n51014) );
  XNOR U60616 ( .A(y[522]), .B(x[522]), .Z(n51011) );
  XNOR U60617 ( .A(n51012), .B(n51013), .Z(n51010) );
  XNOR U60618 ( .A(y[523]), .B(x[523]), .Z(n51013) );
  XNOR U60619 ( .A(y[524]), .B(x[524]), .Z(n51012) );
  XNOR U60620 ( .A(n51004), .B(n51005), .Z(n51015) );
  XNOR U60621 ( .A(y[519]), .B(x[519]), .Z(n51005) );
  XNOR U60622 ( .A(n51006), .B(n51007), .Z(n51004) );
  XNOR U60623 ( .A(y[520]), .B(x[520]), .Z(n51007) );
  XNOR U60624 ( .A(y[521]), .B(x[521]), .Z(n51006) );
  NAND U60625 ( .A(n51071), .B(n51072), .Z(N60869) );
  NANDN U60626 ( .A(n51073), .B(n51074), .Z(n51072) );
  OR U60627 ( .A(n51075), .B(n51076), .Z(n51074) );
  NAND U60628 ( .A(n51075), .B(n51076), .Z(n51071) );
  XOR U60629 ( .A(n51075), .B(n51077), .Z(N60868) );
  XNOR U60630 ( .A(n51073), .B(n51076), .Z(n51077) );
  AND U60631 ( .A(n51078), .B(n51079), .Z(n51076) );
  NANDN U60632 ( .A(n51080), .B(n51081), .Z(n51079) );
  NANDN U60633 ( .A(n51082), .B(n51083), .Z(n51081) );
  NANDN U60634 ( .A(n51083), .B(n51082), .Z(n51078) );
  NAND U60635 ( .A(n51084), .B(n51085), .Z(n51073) );
  NANDN U60636 ( .A(n51086), .B(n51087), .Z(n51085) );
  OR U60637 ( .A(n51088), .B(n51089), .Z(n51087) );
  NAND U60638 ( .A(n51089), .B(n51088), .Z(n51084) );
  AND U60639 ( .A(n51090), .B(n51091), .Z(n51075) );
  NANDN U60640 ( .A(n51092), .B(n51093), .Z(n51091) );
  NANDN U60641 ( .A(n51094), .B(n51095), .Z(n51093) );
  NANDN U60642 ( .A(n51095), .B(n51094), .Z(n51090) );
  XOR U60643 ( .A(n51089), .B(n51096), .Z(N60867) );
  XOR U60644 ( .A(n51086), .B(n51088), .Z(n51096) );
  XNOR U60645 ( .A(n51082), .B(n51097), .Z(n51088) );
  XNOR U60646 ( .A(n51080), .B(n51083), .Z(n51097) );
  NAND U60647 ( .A(n51098), .B(n51099), .Z(n51083) );
  NAND U60648 ( .A(n51100), .B(n51101), .Z(n51099) );
  OR U60649 ( .A(n51102), .B(n51103), .Z(n51100) );
  NANDN U60650 ( .A(n51104), .B(n51102), .Z(n51098) );
  IV U60651 ( .A(n51103), .Z(n51104) );
  NAND U60652 ( .A(n51105), .B(n51106), .Z(n51080) );
  NAND U60653 ( .A(n51107), .B(n51108), .Z(n51106) );
  NANDN U60654 ( .A(n51109), .B(n51110), .Z(n51107) );
  NANDN U60655 ( .A(n51110), .B(n51109), .Z(n51105) );
  AND U60656 ( .A(n51111), .B(n51112), .Z(n51082) );
  NAND U60657 ( .A(n51113), .B(n51114), .Z(n51112) );
  OR U60658 ( .A(n51115), .B(n51116), .Z(n51113) );
  NANDN U60659 ( .A(n51117), .B(n51115), .Z(n51111) );
  NAND U60660 ( .A(n51118), .B(n51119), .Z(n51086) );
  NANDN U60661 ( .A(n51120), .B(n51121), .Z(n51119) );
  OR U60662 ( .A(n51122), .B(n51123), .Z(n51121) );
  NANDN U60663 ( .A(n51124), .B(n51122), .Z(n51118) );
  IV U60664 ( .A(n51123), .Z(n51124) );
  XNOR U60665 ( .A(n51094), .B(n51125), .Z(n51089) );
  XNOR U60666 ( .A(n51092), .B(n51095), .Z(n51125) );
  NAND U60667 ( .A(n51126), .B(n51127), .Z(n51095) );
  NAND U60668 ( .A(n51128), .B(n51129), .Z(n51127) );
  OR U60669 ( .A(n51130), .B(n51131), .Z(n51128) );
  NANDN U60670 ( .A(n51132), .B(n51130), .Z(n51126) );
  IV U60671 ( .A(n51131), .Z(n51132) );
  NAND U60672 ( .A(n51133), .B(n51134), .Z(n51092) );
  NAND U60673 ( .A(n51135), .B(n51136), .Z(n51134) );
  NANDN U60674 ( .A(n51137), .B(n51138), .Z(n51135) );
  NANDN U60675 ( .A(n51138), .B(n51137), .Z(n51133) );
  AND U60676 ( .A(n51139), .B(n51140), .Z(n51094) );
  NAND U60677 ( .A(n51141), .B(n51142), .Z(n51140) );
  OR U60678 ( .A(n51143), .B(n51144), .Z(n51141) );
  NANDN U60679 ( .A(n51145), .B(n51143), .Z(n51139) );
  XNOR U60680 ( .A(n51120), .B(n51146), .Z(N60866) );
  XOR U60681 ( .A(n51122), .B(n51123), .Z(n51146) );
  XNOR U60682 ( .A(n51136), .B(n51147), .Z(n51123) );
  XOR U60683 ( .A(n51137), .B(n51138), .Z(n51147) );
  XOR U60684 ( .A(n51143), .B(n51148), .Z(n51138) );
  XOR U60685 ( .A(n51142), .B(n51145), .Z(n51148) );
  IV U60686 ( .A(n51144), .Z(n51145) );
  NAND U60687 ( .A(n51149), .B(n51150), .Z(n51144) );
  OR U60688 ( .A(n51151), .B(n51152), .Z(n51150) );
  OR U60689 ( .A(n51153), .B(n51154), .Z(n51149) );
  NAND U60690 ( .A(n51155), .B(n51156), .Z(n51142) );
  OR U60691 ( .A(n51157), .B(n51158), .Z(n51156) );
  OR U60692 ( .A(n51159), .B(n51160), .Z(n51155) );
  NOR U60693 ( .A(n51161), .B(n51162), .Z(n51143) );
  ANDN U60694 ( .B(n51163), .A(n51164), .Z(n51137) );
  XNOR U60695 ( .A(n51130), .B(n51165), .Z(n51136) );
  XNOR U60696 ( .A(n51129), .B(n51131), .Z(n51165) );
  NAND U60697 ( .A(n51166), .B(n51167), .Z(n51131) );
  OR U60698 ( .A(n51168), .B(n51169), .Z(n51167) );
  OR U60699 ( .A(n51170), .B(n51171), .Z(n51166) );
  NAND U60700 ( .A(n51172), .B(n51173), .Z(n51129) );
  OR U60701 ( .A(n51174), .B(n51175), .Z(n51173) );
  OR U60702 ( .A(n51176), .B(n51177), .Z(n51172) );
  ANDN U60703 ( .B(n51178), .A(n51179), .Z(n51130) );
  IV U60704 ( .A(n51180), .Z(n51178) );
  ANDN U60705 ( .B(n51181), .A(n51182), .Z(n51122) );
  XOR U60706 ( .A(n51108), .B(n51183), .Z(n51120) );
  XOR U60707 ( .A(n51109), .B(n51110), .Z(n51183) );
  XOR U60708 ( .A(n51115), .B(n51184), .Z(n51110) );
  XOR U60709 ( .A(n51114), .B(n51117), .Z(n51184) );
  IV U60710 ( .A(n51116), .Z(n51117) );
  NAND U60711 ( .A(n51185), .B(n51186), .Z(n51116) );
  OR U60712 ( .A(n51187), .B(n51188), .Z(n51186) );
  OR U60713 ( .A(n51189), .B(n51190), .Z(n51185) );
  NAND U60714 ( .A(n51191), .B(n51192), .Z(n51114) );
  OR U60715 ( .A(n51193), .B(n51194), .Z(n51192) );
  OR U60716 ( .A(n51195), .B(n51196), .Z(n51191) );
  NOR U60717 ( .A(n51197), .B(n51198), .Z(n51115) );
  ANDN U60718 ( .B(n51199), .A(n51200), .Z(n51109) );
  IV U60719 ( .A(n51201), .Z(n51199) );
  XNOR U60720 ( .A(n51102), .B(n51202), .Z(n51108) );
  XNOR U60721 ( .A(n51101), .B(n51103), .Z(n51202) );
  NAND U60722 ( .A(n51203), .B(n51204), .Z(n51103) );
  OR U60723 ( .A(n51205), .B(n51206), .Z(n51204) );
  OR U60724 ( .A(n51207), .B(n51208), .Z(n51203) );
  NAND U60725 ( .A(n51209), .B(n51210), .Z(n51101) );
  OR U60726 ( .A(n51211), .B(n51212), .Z(n51210) );
  OR U60727 ( .A(n51213), .B(n51214), .Z(n51209) );
  ANDN U60728 ( .B(n51215), .A(n51216), .Z(n51102) );
  IV U60729 ( .A(n51217), .Z(n51215) );
  XNOR U60730 ( .A(n51182), .B(n51181), .Z(N60865) );
  XOR U60731 ( .A(n51201), .B(n51200), .Z(n51181) );
  XNOR U60732 ( .A(n51216), .B(n51217), .Z(n51200) );
  XNOR U60733 ( .A(n51211), .B(n51212), .Z(n51217) );
  XNOR U60734 ( .A(n51213), .B(n51214), .Z(n51212) );
  XNOR U60735 ( .A(y[517]), .B(x[517]), .Z(n51214) );
  XNOR U60736 ( .A(y[518]), .B(x[518]), .Z(n51213) );
  XNOR U60737 ( .A(y[516]), .B(x[516]), .Z(n51211) );
  XNOR U60738 ( .A(n51205), .B(n51206), .Z(n51216) );
  XNOR U60739 ( .A(y[513]), .B(x[513]), .Z(n51206) );
  XNOR U60740 ( .A(n51207), .B(n51208), .Z(n51205) );
  XNOR U60741 ( .A(y[514]), .B(x[514]), .Z(n51208) );
  XNOR U60742 ( .A(y[515]), .B(x[515]), .Z(n51207) );
  XNOR U60743 ( .A(n51198), .B(n51197), .Z(n51201) );
  XNOR U60744 ( .A(n51193), .B(n51194), .Z(n51197) );
  XNOR U60745 ( .A(y[510]), .B(x[510]), .Z(n51194) );
  XNOR U60746 ( .A(n51195), .B(n51196), .Z(n51193) );
  XNOR U60747 ( .A(y[511]), .B(x[511]), .Z(n51196) );
  XNOR U60748 ( .A(y[512]), .B(x[512]), .Z(n51195) );
  XNOR U60749 ( .A(n51187), .B(n51188), .Z(n51198) );
  XNOR U60750 ( .A(y[507]), .B(x[507]), .Z(n51188) );
  XNOR U60751 ( .A(n51189), .B(n51190), .Z(n51187) );
  XNOR U60752 ( .A(y[508]), .B(x[508]), .Z(n51190) );
  XNOR U60753 ( .A(y[509]), .B(x[509]), .Z(n51189) );
  XOR U60754 ( .A(n51163), .B(n51164), .Z(n51182) );
  XNOR U60755 ( .A(n51179), .B(n51180), .Z(n51164) );
  XNOR U60756 ( .A(n51174), .B(n51175), .Z(n51180) );
  XNOR U60757 ( .A(n51176), .B(n51177), .Z(n51175) );
  XNOR U60758 ( .A(y[505]), .B(x[505]), .Z(n51177) );
  XNOR U60759 ( .A(y[506]), .B(x[506]), .Z(n51176) );
  XNOR U60760 ( .A(y[504]), .B(x[504]), .Z(n51174) );
  XNOR U60761 ( .A(n51168), .B(n51169), .Z(n51179) );
  XNOR U60762 ( .A(y[501]), .B(x[501]), .Z(n51169) );
  XNOR U60763 ( .A(n51170), .B(n51171), .Z(n51168) );
  XNOR U60764 ( .A(y[502]), .B(x[502]), .Z(n51171) );
  XNOR U60765 ( .A(y[503]), .B(x[503]), .Z(n51170) );
  XOR U60766 ( .A(n51162), .B(n51161), .Z(n51163) );
  XNOR U60767 ( .A(n51157), .B(n51158), .Z(n51161) );
  XNOR U60768 ( .A(y[498]), .B(x[498]), .Z(n51158) );
  XNOR U60769 ( .A(n51159), .B(n51160), .Z(n51157) );
  XNOR U60770 ( .A(y[499]), .B(x[499]), .Z(n51160) );
  XNOR U60771 ( .A(y[500]), .B(x[500]), .Z(n51159) );
  XNOR U60772 ( .A(n51151), .B(n51152), .Z(n51162) );
  XNOR U60773 ( .A(y[495]), .B(x[495]), .Z(n51152) );
  XNOR U60774 ( .A(n51153), .B(n51154), .Z(n51151) );
  XNOR U60775 ( .A(y[496]), .B(x[496]), .Z(n51154) );
  XNOR U60776 ( .A(y[497]), .B(x[497]), .Z(n51153) );
  NAND U60777 ( .A(n51218), .B(n51219), .Z(N60856) );
  NANDN U60778 ( .A(n51220), .B(n51221), .Z(n51219) );
  OR U60779 ( .A(n51222), .B(n51223), .Z(n51221) );
  NAND U60780 ( .A(n51222), .B(n51223), .Z(n51218) );
  XOR U60781 ( .A(n51222), .B(n51224), .Z(N60855) );
  XNOR U60782 ( .A(n51220), .B(n51223), .Z(n51224) );
  AND U60783 ( .A(n51225), .B(n51226), .Z(n51223) );
  NANDN U60784 ( .A(n51227), .B(n51228), .Z(n51226) );
  NANDN U60785 ( .A(n51229), .B(n51230), .Z(n51228) );
  NANDN U60786 ( .A(n51230), .B(n51229), .Z(n51225) );
  NAND U60787 ( .A(n51231), .B(n51232), .Z(n51220) );
  NANDN U60788 ( .A(n51233), .B(n51234), .Z(n51232) );
  OR U60789 ( .A(n51235), .B(n51236), .Z(n51234) );
  NAND U60790 ( .A(n51236), .B(n51235), .Z(n51231) );
  AND U60791 ( .A(n51237), .B(n51238), .Z(n51222) );
  NANDN U60792 ( .A(n51239), .B(n51240), .Z(n51238) );
  NANDN U60793 ( .A(n51241), .B(n51242), .Z(n51240) );
  NANDN U60794 ( .A(n51242), .B(n51241), .Z(n51237) );
  XOR U60795 ( .A(n51236), .B(n51243), .Z(N60854) );
  XOR U60796 ( .A(n51233), .B(n51235), .Z(n51243) );
  XNOR U60797 ( .A(n51229), .B(n51244), .Z(n51235) );
  XNOR U60798 ( .A(n51227), .B(n51230), .Z(n51244) );
  NAND U60799 ( .A(n51245), .B(n51246), .Z(n51230) );
  NAND U60800 ( .A(n51247), .B(n51248), .Z(n51246) );
  OR U60801 ( .A(n51249), .B(n51250), .Z(n51247) );
  NANDN U60802 ( .A(n51251), .B(n51249), .Z(n51245) );
  IV U60803 ( .A(n51250), .Z(n51251) );
  NAND U60804 ( .A(n51252), .B(n51253), .Z(n51227) );
  NAND U60805 ( .A(n51254), .B(n51255), .Z(n51253) );
  NANDN U60806 ( .A(n51256), .B(n51257), .Z(n51254) );
  NANDN U60807 ( .A(n51257), .B(n51256), .Z(n51252) );
  AND U60808 ( .A(n51258), .B(n51259), .Z(n51229) );
  NAND U60809 ( .A(n51260), .B(n51261), .Z(n51259) );
  OR U60810 ( .A(n51262), .B(n51263), .Z(n51260) );
  NANDN U60811 ( .A(n51264), .B(n51262), .Z(n51258) );
  NAND U60812 ( .A(n51265), .B(n51266), .Z(n51233) );
  NANDN U60813 ( .A(n51267), .B(n51268), .Z(n51266) );
  OR U60814 ( .A(n51269), .B(n51270), .Z(n51268) );
  NANDN U60815 ( .A(n51271), .B(n51269), .Z(n51265) );
  IV U60816 ( .A(n51270), .Z(n51271) );
  XNOR U60817 ( .A(n51241), .B(n51272), .Z(n51236) );
  XNOR U60818 ( .A(n51239), .B(n51242), .Z(n51272) );
  NAND U60819 ( .A(n51273), .B(n51274), .Z(n51242) );
  NAND U60820 ( .A(n51275), .B(n51276), .Z(n51274) );
  OR U60821 ( .A(n51277), .B(n51278), .Z(n51275) );
  NANDN U60822 ( .A(n51279), .B(n51277), .Z(n51273) );
  IV U60823 ( .A(n51278), .Z(n51279) );
  NAND U60824 ( .A(n51280), .B(n51281), .Z(n51239) );
  NAND U60825 ( .A(n51282), .B(n51283), .Z(n51281) );
  NANDN U60826 ( .A(n51284), .B(n51285), .Z(n51282) );
  NANDN U60827 ( .A(n51285), .B(n51284), .Z(n51280) );
  AND U60828 ( .A(n51286), .B(n51287), .Z(n51241) );
  NAND U60829 ( .A(n51288), .B(n51289), .Z(n51287) );
  OR U60830 ( .A(n51290), .B(n51291), .Z(n51288) );
  NANDN U60831 ( .A(n51292), .B(n51290), .Z(n51286) );
  XNOR U60832 ( .A(n51267), .B(n51293), .Z(N60853) );
  XOR U60833 ( .A(n51269), .B(n51270), .Z(n51293) );
  XNOR U60834 ( .A(n51283), .B(n51294), .Z(n51270) );
  XOR U60835 ( .A(n51284), .B(n51285), .Z(n51294) );
  XOR U60836 ( .A(n51290), .B(n51295), .Z(n51285) );
  XOR U60837 ( .A(n51289), .B(n51292), .Z(n51295) );
  IV U60838 ( .A(n51291), .Z(n51292) );
  NAND U60839 ( .A(n51296), .B(n51297), .Z(n51291) );
  OR U60840 ( .A(n51298), .B(n51299), .Z(n51297) );
  OR U60841 ( .A(n51300), .B(n51301), .Z(n51296) );
  NAND U60842 ( .A(n51302), .B(n51303), .Z(n51289) );
  OR U60843 ( .A(n51304), .B(n51305), .Z(n51303) );
  OR U60844 ( .A(n51306), .B(n51307), .Z(n51302) );
  NOR U60845 ( .A(n51308), .B(n51309), .Z(n51290) );
  ANDN U60846 ( .B(n51310), .A(n51311), .Z(n51284) );
  XNOR U60847 ( .A(n51277), .B(n51312), .Z(n51283) );
  XNOR U60848 ( .A(n51276), .B(n51278), .Z(n51312) );
  NAND U60849 ( .A(n51313), .B(n51314), .Z(n51278) );
  OR U60850 ( .A(n51315), .B(n51316), .Z(n51314) );
  OR U60851 ( .A(n51317), .B(n51318), .Z(n51313) );
  NAND U60852 ( .A(n51319), .B(n51320), .Z(n51276) );
  OR U60853 ( .A(n51321), .B(n51322), .Z(n51320) );
  OR U60854 ( .A(n51323), .B(n51324), .Z(n51319) );
  ANDN U60855 ( .B(n51325), .A(n51326), .Z(n51277) );
  IV U60856 ( .A(n51327), .Z(n51325) );
  ANDN U60857 ( .B(n51328), .A(n51329), .Z(n51269) );
  XOR U60858 ( .A(n51255), .B(n51330), .Z(n51267) );
  XOR U60859 ( .A(n51256), .B(n51257), .Z(n51330) );
  XOR U60860 ( .A(n51262), .B(n51331), .Z(n51257) );
  XOR U60861 ( .A(n51261), .B(n51264), .Z(n51331) );
  IV U60862 ( .A(n51263), .Z(n51264) );
  NAND U60863 ( .A(n51332), .B(n51333), .Z(n51263) );
  OR U60864 ( .A(n51334), .B(n51335), .Z(n51333) );
  OR U60865 ( .A(n51336), .B(n51337), .Z(n51332) );
  NAND U60866 ( .A(n51338), .B(n51339), .Z(n51261) );
  OR U60867 ( .A(n51340), .B(n51341), .Z(n51339) );
  OR U60868 ( .A(n51342), .B(n51343), .Z(n51338) );
  NOR U60869 ( .A(n51344), .B(n51345), .Z(n51262) );
  ANDN U60870 ( .B(n51346), .A(n51347), .Z(n51256) );
  IV U60871 ( .A(n51348), .Z(n51346) );
  XNOR U60872 ( .A(n51249), .B(n51349), .Z(n51255) );
  XNOR U60873 ( .A(n51248), .B(n51250), .Z(n51349) );
  NAND U60874 ( .A(n51350), .B(n51351), .Z(n51250) );
  OR U60875 ( .A(n51352), .B(n51353), .Z(n51351) );
  OR U60876 ( .A(n51354), .B(n51355), .Z(n51350) );
  NAND U60877 ( .A(n51356), .B(n51357), .Z(n51248) );
  OR U60878 ( .A(n51358), .B(n51359), .Z(n51357) );
  OR U60879 ( .A(n51360), .B(n51361), .Z(n51356) );
  ANDN U60880 ( .B(n51362), .A(n51363), .Z(n51249) );
  IV U60881 ( .A(n51364), .Z(n51362) );
  XNOR U60882 ( .A(n51329), .B(n51328), .Z(N60852) );
  XOR U60883 ( .A(n51348), .B(n51347), .Z(n51328) );
  XNOR U60884 ( .A(n51363), .B(n51364), .Z(n51347) );
  XNOR U60885 ( .A(n51358), .B(n51359), .Z(n51364) );
  XNOR U60886 ( .A(n51360), .B(n51361), .Z(n51359) );
  XNOR U60887 ( .A(y[493]), .B(x[493]), .Z(n51361) );
  XNOR U60888 ( .A(y[494]), .B(x[494]), .Z(n51360) );
  XNOR U60889 ( .A(y[492]), .B(x[492]), .Z(n51358) );
  XNOR U60890 ( .A(n51352), .B(n51353), .Z(n51363) );
  XNOR U60891 ( .A(y[489]), .B(x[489]), .Z(n51353) );
  XNOR U60892 ( .A(n51354), .B(n51355), .Z(n51352) );
  XNOR U60893 ( .A(y[490]), .B(x[490]), .Z(n51355) );
  XNOR U60894 ( .A(y[491]), .B(x[491]), .Z(n51354) );
  XNOR U60895 ( .A(n51345), .B(n51344), .Z(n51348) );
  XNOR U60896 ( .A(n51340), .B(n51341), .Z(n51344) );
  XNOR U60897 ( .A(y[486]), .B(x[486]), .Z(n51341) );
  XNOR U60898 ( .A(n51342), .B(n51343), .Z(n51340) );
  XNOR U60899 ( .A(y[487]), .B(x[487]), .Z(n51343) );
  XNOR U60900 ( .A(y[488]), .B(x[488]), .Z(n51342) );
  XNOR U60901 ( .A(n51334), .B(n51335), .Z(n51345) );
  XNOR U60902 ( .A(y[483]), .B(x[483]), .Z(n51335) );
  XNOR U60903 ( .A(n51336), .B(n51337), .Z(n51334) );
  XNOR U60904 ( .A(y[484]), .B(x[484]), .Z(n51337) );
  XNOR U60905 ( .A(y[485]), .B(x[485]), .Z(n51336) );
  XOR U60906 ( .A(n51310), .B(n51311), .Z(n51329) );
  XNOR U60907 ( .A(n51326), .B(n51327), .Z(n51311) );
  XNOR U60908 ( .A(n51321), .B(n51322), .Z(n51327) );
  XNOR U60909 ( .A(n51323), .B(n51324), .Z(n51322) );
  XNOR U60910 ( .A(y[481]), .B(x[481]), .Z(n51324) );
  XNOR U60911 ( .A(y[482]), .B(x[482]), .Z(n51323) );
  XNOR U60912 ( .A(y[480]), .B(x[480]), .Z(n51321) );
  XNOR U60913 ( .A(n51315), .B(n51316), .Z(n51326) );
  XNOR U60914 ( .A(y[477]), .B(x[477]), .Z(n51316) );
  XNOR U60915 ( .A(n51317), .B(n51318), .Z(n51315) );
  XNOR U60916 ( .A(y[478]), .B(x[478]), .Z(n51318) );
  XNOR U60917 ( .A(y[479]), .B(x[479]), .Z(n51317) );
  XOR U60918 ( .A(n51309), .B(n51308), .Z(n51310) );
  XNOR U60919 ( .A(n51304), .B(n51305), .Z(n51308) );
  XNOR U60920 ( .A(y[474]), .B(x[474]), .Z(n51305) );
  XNOR U60921 ( .A(n51306), .B(n51307), .Z(n51304) );
  XNOR U60922 ( .A(y[475]), .B(x[475]), .Z(n51307) );
  XNOR U60923 ( .A(y[476]), .B(x[476]), .Z(n51306) );
  XNOR U60924 ( .A(n51298), .B(n51299), .Z(n51309) );
  XNOR U60925 ( .A(y[471]), .B(x[471]), .Z(n51299) );
  XNOR U60926 ( .A(n51300), .B(n51301), .Z(n51298) );
  XNOR U60927 ( .A(y[472]), .B(x[472]), .Z(n51301) );
  XNOR U60928 ( .A(y[473]), .B(x[473]), .Z(n51300) );
  NAND U60929 ( .A(n51365), .B(n51366), .Z(N60843) );
  NANDN U60930 ( .A(n51367), .B(n51368), .Z(n51366) );
  OR U60931 ( .A(n51369), .B(n51370), .Z(n51368) );
  NAND U60932 ( .A(n51369), .B(n51370), .Z(n51365) );
  XOR U60933 ( .A(n51369), .B(n51371), .Z(N60842) );
  XNOR U60934 ( .A(n51367), .B(n51370), .Z(n51371) );
  AND U60935 ( .A(n51372), .B(n51373), .Z(n51370) );
  NANDN U60936 ( .A(n51374), .B(n51375), .Z(n51373) );
  NANDN U60937 ( .A(n51376), .B(n51377), .Z(n51375) );
  NANDN U60938 ( .A(n51377), .B(n51376), .Z(n51372) );
  NAND U60939 ( .A(n51378), .B(n51379), .Z(n51367) );
  NANDN U60940 ( .A(n51380), .B(n51381), .Z(n51379) );
  OR U60941 ( .A(n51382), .B(n51383), .Z(n51381) );
  NAND U60942 ( .A(n51383), .B(n51382), .Z(n51378) );
  AND U60943 ( .A(n51384), .B(n51385), .Z(n51369) );
  NANDN U60944 ( .A(n51386), .B(n51387), .Z(n51385) );
  NANDN U60945 ( .A(n51388), .B(n51389), .Z(n51387) );
  NANDN U60946 ( .A(n51389), .B(n51388), .Z(n51384) );
  XOR U60947 ( .A(n51383), .B(n51390), .Z(N60841) );
  XOR U60948 ( .A(n51380), .B(n51382), .Z(n51390) );
  XNOR U60949 ( .A(n51376), .B(n51391), .Z(n51382) );
  XNOR U60950 ( .A(n51374), .B(n51377), .Z(n51391) );
  NAND U60951 ( .A(n51392), .B(n51393), .Z(n51377) );
  NAND U60952 ( .A(n51394), .B(n51395), .Z(n51393) );
  OR U60953 ( .A(n51396), .B(n51397), .Z(n51394) );
  NANDN U60954 ( .A(n51398), .B(n51396), .Z(n51392) );
  IV U60955 ( .A(n51397), .Z(n51398) );
  NAND U60956 ( .A(n51399), .B(n51400), .Z(n51374) );
  NAND U60957 ( .A(n51401), .B(n51402), .Z(n51400) );
  NANDN U60958 ( .A(n51403), .B(n51404), .Z(n51401) );
  NANDN U60959 ( .A(n51404), .B(n51403), .Z(n51399) );
  AND U60960 ( .A(n51405), .B(n51406), .Z(n51376) );
  NAND U60961 ( .A(n51407), .B(n51408), .Z(n51406) );
  OR U60962 ( .A(n51409), .B(n51410), .Z(n51407) );
  NANDN U60963 ( .A(n51411), .B(n51409), .Z(n51405) );
  NAND U60964 ( .A(n51412), .B(n51413), .Z(n51380) );
  NANDN U60965 ( .A(n51414), .B(n51415), .Z(n51413) );
  OR U60966 ( .A(n51416), .B(n51417), .Z(n51415) );
  NANDN U60967 ( .A(n51418), .B(n51416), .Z(n51412) );
  IV U60968 ( .A(n51417), .Z(n51418) );
  XNOR U60969 ( .A(n51388), .B(n51419), .Z(n51383) );
  XNOR U60970 ( .A(n51386), .B(n51389), .Z(n51419) );
  NAND U60971 ( .A(n51420), .B(n51421), .Z(n51389) );
  NAND U60972 ( .A(n51422), .B(n51423), .Z(n51421) );
  OR U60973 ( .A(n51424), .B(n51425), .Z(n51422) );
  NANDN U60974 ( .A(n51426), .B(n51424), .Z(n51420) );
  IV U60975 ( .A(n51425), .Z(n51426) );
  NAND U60976 ( .A(n51427), .B(n51428), .Z(n51386) );
  NAND U60977 ( .A(n51429), .B(n51430), .Z(n51428) );
  NANDN U60978 ( .A(n51431), .B(n51432), .Z(n51429) );
  NANDN U60979 ( .A(n51432), .B(n51431), .Z(n51427) );
  AND U60980 ( .A(n51433), .B(n51434), .Z(n51388) );
  NAND U60981 ( .A(n51435), .B(n51436), .Z(n51434) );
  OR U60982 ( .A(n51437), .B(n51438), .Z(n51435) );
  NANDN U60983 ( .A(n51439), .B(n51437), .Z(n51433) );
  XNOR U60984 ( .A(n51414), .B(n51440), .Z(N60840) );
  XOR U60985 ( .A(n51416), .B(n51417), .Z(n51440) );
  XNOR U60986 ( .A(n51430), .B(n51441), .Z(n51417) );
  XOR U60987 ( .A(n51431), .B(n51432), .Z(n51441) );
  XOR U60988 ( .A(n51437), .B(n51442), .Z(n51432) );
  XOR U60989 ( .A(n51436), .B(n51439), .Z(n51442) );
  IV U60990 ( .A(n51438), .Z(n51439) );
  NAND U60991 ( .A(n51443), .B(n51444), .Z(n51438) );
  OR U60992 ( .A(n51445), .B(n51446), .Z(n51444) );
  OR U60993 ( .A(n51447), .B(n51448), .Z(n51443) );
  NAND U60994 ( .A(n51449), .B(n51450), .Z(n51436) );
  OR U60995 ( .A(n51451), .B(n51452), .Z(n51450) );
  OR U60996 ( .A(n51453), .B(n51454), .Z(n51449) );
  NOR U60997 ( .A(n51455), .B(n51456), .Z(n51437) );
  ANDN U60998 ( .B(n51457), .A(n51458), .Z(n51431) );
  XNOR U60999 ( .A(n51424), .B(n51459), .Z(n51430) );
  XNOR U61000 ( .A(n51423), .B(n51425), .Z(n51459) );
  NAND U61001 ( .A(n51460), .B(n51461), .Z(n51425) );
  OR U61002 ( .A(n51462), .B(n51463), .Z(n51461) );
  OR U61003 ( .A(n51464), .B(n51465), .Z(n51460) );
  NAND U61004 ( .A(n51466), .B(n51467), .Z(n51423) );
  OR U61005 ( .A(n51468), .B(n51469), .Z(n51467) );
  OR U61006 ( .A(n51470), .B(n51471), .Z(n51466) );
  ANDN U61007 ( .B(n51472), .A(n51473), .Z(n51424) );
  IV U61008 ( .A(n51474), .Z(n51472) );
  ANDN U61009 ( .B(n51475), .A(n51476), .Z(n51416) );
  XOR U61010 ( .A(n51402), .B(n51477), .Z(n51414) );
  XOR U61011 ( .A(n51403), .B(n51404), .Z(n51477) );
  XOR U61012 ( .A(n51409), .B(n51478), .Z(n51404) );
  XOR U61013 ( .A(n51408), .B(n51411), .Z(n51478) );
  IV U61014 ( .A(n51410), .Z(n51411) );
  NAND U61015 ( .A(n51479), .B(n51480), .Z(n51410) );
  OR U61016 ( .A(n51481), .B(n51482), .Z(n51480) );
  OR U61017 ( .A(n51483), .B(n51484), .Z(n51479) );
  NAND U61018 ( .A(n51485), .B(n51486), .Z(n51408) );
  OR U61019 ( .A(n51487), .B(n51488), .Z(n51486) );
  OR U61020 ( .A(n51489), .B(n51490), .Z(n51485) );
  NOR U61021 ( .A(n51491), .B(n51492), .Z(n51409) );
  ANDN U61022 ( .B(n51493), .A(n51494), .Z(n51403) );
  IV U61023 ( .A(n51495), .Z(n51493) );
  XNOR U61024 ( .A(n51396), .B(n51496), .Z(n51402) );
  XNOR U61025 ( .A(n51395), .B(n51397), .Z(n51496) );
  NAND U61026 ( .A(n51497), .B(n51498), .Z(n51397) );
  OR U61027 ( .A(n51499), .B(n51500), .Z(n51498) );
  OR U61028 ( .A(n51501), .B(n51502), .Z(n51497) );
  NAND U61029 ( .A(n51503), .B(n51504), .Z(n51395) );
  OR U61030 ( .A(n51505), .B(n51506), .Z(n51504) );
  OR U61031 ( .A(n51507), .B(n51508), .Z(n51503) );
  ANDN U61032 ( .B(n51509), .A(n51510), .Z(n51396) );
  IV U61033 ( .A(n51511), .Z(n51509) );
  XNOR U61034 ( .A(n51476), .B(n51475), .Z(N60839) );
  XOR U61035 ( .A(n51495), .B(n51494), .Z(n51475) );
  XNOR U61036 ( .A(n51510), .B(n51511), .Z(n51494) );
  XNOR U61037 ( .A(n51505), .B(n51506), .Z(n51511) );
  XNOR U61038 ( .A(n51507), .B(n51508), .Z(n51506) );
  XNOR U61039 ( .A(y[469]), .B(x[469]), .Z(n51508) );
  XNOR U61040 ( .A(y[470]), .B(x[470]), .Z(n51507) );
  XNOR U61041 ( .A(y[468]), .B(x[468]), .Z(n51505) );
  XNOR U61042 ( .A(n51499), .B(n51500), .Z(n51510) );
  XNOR U61043 ( .A(y[465]), .B(x[465]), .Z(n51500) );
  XNOR U61044 ( .A(n51501), .B(n51502), .Z(n51499) );
  XNOR U61045 ( .A(y[466]), .B(x[466]), .Z(n51502) );
  XNOR U61046 ( .A(y[467]), .B(x[467]), .Z(n51501) );
  XNOR U61047 ( .A(n51492), .B(n51491), .Z(n51495) );
  XNOR U61048 ( .A(n51487), .B(n51488), .Z(n51491) );
  XNOR U61049 ( .A(y[462]), .B(x[462]), .Z(n51488) );
  XNOR U61050 ( .A(n51489), .B(n51490), .Z(n51487) );
  XNOR U61051 ( .A(y[463]), .B(x[463]), .Z(n51490) );
  XNOR U61052 ( .A(y[464]), .B(x[464]), .Z(n51489) );
  XNOR U61053 ( .A(n51481), .B(n51482), .Z(n51492) );
  XNOR U61054 ( .A(y[459]), .B(x[459]), .Z(n51482) );
  XNOR U61055 ( .A(n51483), .B(n51484), .Z(n51481) );
  XNOR U61056 ( .A(y[460]), .B(x[460]), .Z(n51484) );
  XNOR U61057 ( .A(y[461]), .B(x[461]), .Z(n51483) );
  XOR U61058 ( .A(n51457), .B(n51458), .Z(n51476) );
  XNOR U61059 ( .A(n51473), .B(n51474), .Z(n51458) );
  XNOR U61060 ( .A(n51468), .B(n51469), .Z(n51474) );
  XNOR U61061 ( .A(n51470), .B(n51471), .Z(n51469) );
  XNOR U61062 ( .A(y[457]), .B(x[457]), .Z(n51471) );
  XNOR U61063 ( .A(y[458]), .B(x[458]), .Z(n51470) );
  XNOR U61064 ( .A(y[456]), .B(x[456]), .Z(n51468) );
  XNOR U61065 ( .A(n51462), .B(n51463), .Z(n51473) );
  XNOR U61066 ( .A(y[453]), .B(x[453]), .Z(n51463) );
  XNOR U61067 ( .A(n51464), .B(n51465), .Z(n51462) );
  XNOR U61068 ( .A(y[454]), .B(x[454]), .Z(n51465) );
  XNOR U61069 ( .A(y[455]), .B(x[455]), .Z(n51464) );
  XOR U61070 ( .A(n51456), .B(n51455), .Z(n51457) );
  XNOR U61071 ( .A(n51451), .B(n51452), .Z(n51455) );
  XNOR U61072 ( .A(y[450]), .B(x[450]), .Z(n51452) );
  XNOR U61073 ( .A(n51453), .B(n51454), .Z(n51451) );
  XNOR U61074 ( .A(y[451]), .B(x[451]), .Z(n51454) );
  XNOR U61075 ( .A(y[452]), .B(x[452]), .Z(n51453) );
  XNOR U61076 ( .A(n51445), .B(n51446), .Z(n51456) );
  XNOR U61077 ( .A(y[447]), .B(x[447]), .Z(n51446) );
  XNOR U61078 ( .A(n51447), .B(n51448), .Z(n51445) );
  XNOR U61079 ( .A(y[448]), .B(x[448]), .Z(n51448) );
  XNOR U61080 ( .A(y[449]), .B(x[449]), .Z(n51447) );
  NAND U61081 ( .A(n51512), .B(n51513), .Z(N60830) );
  NANDN U61082 ( .A(n51514), .B(n51515), .Z(n51513) );
  OR U61083 ( .A(n51516), .B(n51517), .Z(n51515) );
  NAND U61084 ( .A(n51516), .B(n51517), .Z(n51512) );
  XOR U61085 ( .A(n51516), .B(n51518), .Z(N60829) );
  XNOR U61086 ( .A(n51514), .B(n51517), .Z(n51518) );
  AND U61087 ( .A(n51519), .B(n51520), .Z(n51517) );
  NANDN U61088 ( .A(n51521), .B(n51522), .Z(n51520) );
  NANDN U61089 ( .A(n51523), .B(n51524), .Z(n51522) );
  NANDN U61090 ( .A(n51524), .B(n51523), .Z(n51519) );
  NAND U61091 ( .A(n51525), .B(n51526), .Z(n51514) );
  NANDN U61092 ( .A(n51527), .B(n51528), .Z(n51526) );
  OR U61093 ( .A(n51529), .B(n51530), .Z(n51528) );
  NAND U61094 ( .A(n51530), .B(n51529), .Z(n51525) );
  AND U61095 ( .A(n51531), .B(n51532), .Z(n51516) );
  NANDN U61096 ( .A(n51533), .B(n51534), .Z(n51532) );
  NANDN U61097 ( .A(n51535), .B(n51536), .Z(n51534) );
  NANDN U61098 ( .A(n51536), .B(n51535), .Z(n51531) );
  XOR U61099 ( .A(n51530), .B(n51537), .Z(N60828) );
  XOR U61100 ( .A(n51527), .B(n51529), .Z(n51537) );
  XNOR U61101 ( .A(n51523), .B(n51538), .Z(n51529) );
  XNOR U61102 ( .A(n51521), .B(n51524), .Z(n51538) );
  NAND U61103 ( .A(n51539), .B(n51540), .Z(n51524) );
  NAND U61104 ( .A(n51541), .B(n51542), .Z(n51540) );
  OR U61105 ( .A(n51543), .B(n51544), .Z(n51541) );
  NANDN U61106 ( .A(n51545), .B(n51543), .Z(n51539) );
  IV U61107 ( .A(n51544), .Z(n51545) );
  NAND U61108 ( .A(n51546), .B(n51547), .Z(n51521) );
  NAND U61109 ( .A(n51548), .B(n51549), .Z(n51547) );
  NANDN U61110 ( .A(n51550), .B(n51551), .Z(n51548) );
  NANDN U61111 ( .A(n51551), .B(n51550), .Z(n51546) );
  AND U61112 ( .A(n51552), .B(n51553), .Z(n51523) );
  NAND U61113 ( .A(n51554), .B(n51555), .Z(n51553) );
  OR U61114 ( .A(n51556), .B(n51557), .Z(n51554) );
  NANDN U61115 ( .A(n51558), .B(n51556), .Z(n51552) );
  NAND U61116 ( .A(n51559), .B(n51560), .Z(n51527) );
  NANDN U61117 ( .A(n51561), .B(n51562), .Z(n51560) );
  OR U61118 ( .A(n51563), .B(n51564), .Z(n51562) );
  NANDN U61119 ( .A(n51565), .B(n51563), .Z(n51559) );
  IV U61120 ( .A(n51564), .Z(n51565) );
  XNOR U61121 ( .A(n51535), .B(n51566), .Z(n51530) );
  XNOR U61122 ( .A(n51533), .B(n51536), .Z(n51566) );
  NAND U61123 ( .A(n51567), .B(n51568), .Z(n51536) );
  NAND U61124 ( .A(n51569), .B(n51570), .Z(n51568) );
  OR U61125 ( .A(n51571), .B(n51572), .Z(n51569) );
  NANDN U61126 ( .A(n51573), .B(n51571), .Z(n51567) );
  IV U61127 ( .A(n51572), .Z(n51573) );
  NAND U61128 ( .A(n51574), .B(n51575), .Z(n51533) );
  NAND U61129 ( .A(n51576), .B(n51577), .Z(n51575) );
  NANDN U61130 ( .A(n51578), .B(n51579), .Z(n51576) );
  NANDN U61131 ( .A(n51579), .B(n51578), .Z(n51574) );
  AND U61132 ( .A(n51580), .B(n51581), .Z(n51535) );
  NAND U61133 ( .A(n51582), .B(n51583), .Z(n51581) );
  OR U61134 ( .A(n51584), .B(n51585), .Z(n51582) );
  NANDN U61135 ( .A(n51586), .B(n51584), .Z(n51580) );
  XNOR U61136 ( .A(n51561), .B(n51587), .Z(N60827) );
  XOR U61137 ( .A(n51563), .B(n51564), .Z(n51587) );
  XNOR U61138 ( .A(n51577), .B(n51588), .Z(n51564) );
  XOR U61139 ( .A(n51578), .B(n51579), .Z(n51588) );
  XOR U61140 ( .A(n51584), .B(n51589), .Z(n51579) );
  XOR U61141 ( .A(n51583), .B(n51586), .Z(n51589) );
  IV U61142 ( .A(n51585), .Z(n51586) );
  NAND U61143 ( .A(n51590), .B(n51591), .Z(n51585) );
  OR U61144 ( .A(n51592), .B(n51593), .Z(n51591) );
  OR U61145 ( .A(n51594), .B(n51595), .Z(n51590) );
  NAND U61146 ( .A(n51596), .B(n51597), .Z(n51583) );
  OR U61147 ( .A(n51598), .B(n51599), .Z(n51597) );
  OR U61148 ( .A(n51600), .B(n51601), .Z(n51596) );
  NOR U61149 ( .A(n51602), .B(n51603), .Z(n51584) );
  ANDN U61150 ( .B(n51604), .A(n51605), .Z(n51578) );
  XNOR U61151 ( .A(n51571), .B(n51606), .Z(n51577) );
  XNOR U61152 ( .A(n51570), .B(n51572), .Z(n51606) );
  NAND U61153 ( .A(n51607), .B(n51608), .Z(n51572) );
  OR U61154 ( .A(n51609), .B(n51610), .Z(n51608) );
  OR U61155 ( .A(n51611), .B(n51612), .Z(n51607) );
  NAND U61156 ( .A(n51613), .B(n51614), .Z(n51570) );
  OR U61157 ( .A(n51615), .B(n51616), .Z(n51614) );
  OR U61158 ( .A(n51617), .B(n51618), .Z(n51613) );
  ANDN U61159 ( .B(n51619), .A(n51620), .Z(n51571) );
  IV U61160 ( .A(n51621), .Z(n51619) );
  ANDN U61161 ( .B(n51622), .A(n51623), .Z(n51563) );
  XOR U61162 ( .A(n51549), .B(n51624), .Z(n51561) );
  XOR U61163 ( .A(n51550), .B(n51551), .Z(n51624) );
  XOR U61164 ( .A(n51556), .B(n51625), .Z(n51551) );
  XOR U61165 ( .A(n51555), .B(n51558), .Z(n51625) );
  IV U61166 ( .A(n51557), .Z(n51558) );
  NAND U61167 ( .A(n51626), .B(n51627), .Z(n51557) );
  OR U61168 ( .A(n51628), .B(n51629), .Z(n51627) );
  OR U61169 ( .A(n51630), .B(n51631), .Z(n51626) );
  NAND U61170 ( .A(n51632), .B(n51633), .Z(n51555) );
  OR U61171 ( .A(n51634), .B(n51635), .Z(n51633) );
  OR U61172 ( .A(n51636), .B(n51637), .Z(n51632) );
  NOR U61173 ( .A(n51638), .B(n51639), .Z(n51556) );
  ANDN U61174 ( .B(n51640), .A(n51641), .Z(n51550) );
  IV U61175 ( .A(n51642), .Z(n51640) );
  XNOR U61176 ( .A(n51543), .B(n51643), .Z(n51549) );
  XNOR U61177 ( .A(n51542), .B(n51544), .Z(n51643) );
  NAND U61178 ( .A(n51644), .B(n51645), .Z(n51544) );
  OR U61179 ( .A(n51646), .B(n51647), .Z(n51645) );
  OR U61180 ( .A(n51648), .B(n51649), .Z(n51644) );
  NAND U61181 ( .A(n51650), .B(n51651), .Z(n51542) );
  OR U61182 ( .A(n51652), .B(n51653), .Z(n51651) );
  OR U61183 ( .A(n51654), .B(n51655), .Z(n51650) );
  ANDN U61184 ( .B(n51656), .A(n51657), .Z(n51543) );
  IV U61185 ( .A(n51658), .Z(n51656) );
  XNOR U61186 ( .A(n51623), .B(n51622), .Z(N60826) );
  XOR U61187 ( .A(n51642), .B(n51641), .Z(n51622) );
  XNOR U61188 ( .A(n51657), .B(n51658), .Z(n51641) );
  XNOR U61189 ( .A(n51652), .B(n51653), .Z(n51658) );
  XNOR U61190 ( .A(n51654), .B(n51655), .Z(n51653) );
  XNOR U61191 ( .A(y[445]), .B(x[445]), .Z(n51655) );
  XNOR U61192 ( .A(y[446]), .B(x[446]), .Z(n51654) );
  XNOR U61193 ( .A(y[444]), .B(x[444]), .Z(n51652) );
  XNOR U61194 ( .A(n51646), .B(n51647), .Z(n51657) );
  XNOR U61195 ( .A(y[441]), .B(x[441]), .Z(n51647) );
  XNOR U61196 ( .A(n51648), .B(n51649), .Z(n51646) );
  XNOR U61197 ( .A(y[442]), .B(x[442]), .Z(n51649) );
  XNOR U61198 ( .A(y[443]), .B(x[443]), .Z(n51648) );
  XNOR U61199 ( .A(n51639), .B(n51638), .Z(n51642) );
  XNOR U61200 ( .A(n51634), .B(n51635), .Z(n51638) );
  XNOR U61201 ( .A(y[438]), .B(x[438]), .Z(n51635) );
  XNOR U61202 ( .A(n51636), .B(n51637), .Z(n51634) );
  XNOR U61203 ( .A(y[439]), .B(x[439]), .Z(n51637) );
  XNOR U61204 ( .A(y[440]), .B(x[440]), .Z(n51636) );
  XNOR U61205 ( .A(n51628), .B(n51629), .Z(n51639) );
  XNOR U61206 ( .A(y[435]), .B(x[435]), .Z(n51629) );
  XNOR U61207 ( .A(n51630), .B(n51631), .Z(n51628) );
  XNOR U61208 ( .A(y[436]), .B(x[436]), .Z(n51631) );
  XNOR U61209 ( .A(y[437]), .B(x[437]), .Z(n51630) );
  XOR U61210 ( .A(n51604), .B(n51605), .Z(n51623) );
  XNOR U61211 ( .A(n51620), .B(n51621), .Z(n51605) );
  XNOR U61212 ( .A(n51615), .B(n51616), .Z(n51621) );
  XNOR U61213 ( .A(n51617), .B(n51618), .Z(n51616) );
  XNOR U61214 ( .A(y[433]), .B(x[433]), .Z(n51618) );
  XNOR U61215 ( .A(y[434]), .B(x[434]), .Z(n51617) );
  XNOR U61216 ( .A(y[432]), .B(x[432]), .Z(n51615) );
  XNOR U61217 ( .A(n51609), .B(n51610), .Z(n51620) );
  XNOR U61218 ( .A(y[429]), .B(x[429]), .Z(n51610) );
  XNOR U61219 ( .A(n51611), .B(n51612), .Z(n51609) );
  XNOR U61220 ( .A(y[430]), .B(x[430]), .Z(n51612) );
  XNOR U61221 ( .A(y[431]), .B(x[431]), .Z(n51611) );
  XOR U61222 ( .A(n51603), .B(n51602), .Z(n51604) );
  XNOR U61223 ( .A(n51598), .B(n51599), .Z(n51602) );
  XNOR U61224 ( .A(y[426]), .B(x[426]), .Z(n51599) );
  XNOR U61225 ( .A(n51600), .B(n51601), .Z(n51598) );
  XNOR U61226 ( .A(y[427]), .B(x[427]), .Z(n51601) );
  XNOR U61227 ( .A(y[428]), .B(x[428]), .Z(n51600) );
  XNOR U61228 ( .A(n51592), .B(n51593), .Z(n51603) );
  XNOR U61229 ( .A(y[423]), .B(x[423]), .Z(n51593) );
  XNOR U61230 ( .A(n51594), .B(n51595), .Z(n51592) );
  XNOR U61231 ( .A(y[424]), .B(x[424]), .Z(n51595) );
  XNOR U61232 ( .A(y[425]), .B(x[425]), .Z(n51594) );
  NAND U61233 ( .A(n51659), .B(n51660), .Z(N60817) );
  NANDN U61234 ( .A(n51661), .B(n51662), .Z(n51660) );
  OR U61235 ( .A(n51663), .B(n51664), .Z(n51662) );
  NAND U61236 ( .A(n51663), .B(n51664), .Z(n51659) );
  XOR U61237 ( .A(n51663), .B(n51665), .Z(N60816) );
  XNOR U61238 ( .A(n51661), .B(n51664), .Z(n51665) );
  AND U61239 ( .A(n51666), .B(n51667), .Z(n51664) );
  NANDN U61240 ( .A(n51668), .B(n51669), .Z(n51667) );
  NANDN U61241 ( .A(n51670), .B(n51671), .Z(n51669) );
  NANDN U61242 ( .A(n51671), .B(n51670), .Z(n51666) );
  NAND U61243 ( .A(n51672), .B(n51673), .Z(n51661) );
  NANDN U61244 ( .A(n51674), .B(n51675), .Z(n51673) );
  OR U61245 ( .A(n51676), .B(n51677), .Z(n51675) );
  NAND U61246 ( .A(n51677), .B(n51676), .Z(n51672) );
  AND U61247 ( .A(n51678), .B(n51679), .Z(n51663) );
  NANDN U61248 ( .A(n51680), .B(n51681), .Z(n51679) );
  NANDN U61249 ( .A(n51682), .B(n51683), .Z(n51681) );
  NANDN U61250 ( .A(n51683), .B(n51682), .Z(n51678) );
  XOR U61251 ( .A(n51677), .B(n51684), .Z(N60815) );
  XOR U61252 ( .A(n51674), .B(n51676), .Z(n51684) );
  XNOR U61253 ( .A(n51670), .B(n51685), .Z(n51676) );
  XNOR U61254 ( .A(n51668), .B(n51671), .Z(n51685) );
  NAND U61255 ( .A(n51686), .B(n51687), .Z(n51671) );
  NAND U61256 ( .A(n51688), .B(n51689), .Z(n51687) );
  OR U61257 ( .A(n51690), .B(n51691), .Z(n51688) );
  NANDN U61258 ( .A(n51692), .B(n51690), .Z(n51686) );
  IV U61259 ( .A(n51691), .Z(n51692) );
  NAND U61260 ( .A(n51693), .B(n51694), .Z(n51668) );
  NAND U61261 ( .A(n51695), .B(n51696), .Z(n51694) );
  NANDN U61262 ( .A(n51697), .B(n51698), .Z(n51695) );
  NANDN U61263 ( .A(n51698), .B(n51697), .Z(n51693) );
  AND U61264 ( .A(n51699), .B(n51700), .Z(n51670) );
  NAND U61265 ( .A(n51701), .B(n51702), .Z(n51700) );
  OR U61266 ( .A(n51703), .B(n51704), .Z(n51701) );
  NANDN U61267 ( .A(n51705), .B(n51703), .Z(n51699) );
  NAND U61268 ( .A(n51706), .B(n51707), .Z(n51674) );
  NANDN U61269 ( .A(n51708), .B(n51709), .Z(n51707) );
  OR U61270 ( .A(n51710), .B(n51711), .Z(n51709) );
  NANDN U61271 ( .A(n51712), .B(n51710), .Z(n51706) );
  IV U61272 ( .A(n51711), .Z(n51712) );
  XNOR U61273 ( .A(n51682), .B(n51713), .Z(n51677) );
  XNOR U61274 ( .A(n51680), .B(n51683), .Z(n51713) );
  NAND U61275 ( .A(n51714), .B(n51715), .Z(n51683) );
  NAND U61276 ( .A(n51716), .B(n51717), .Z(n51715) );
  OR U61277 ( .A(n51718), .B(n51719), .Z(n51716) );
  NANDN U61278 ( .A(n51720), .B(n51718), .Z(n51714) );
  IV U61279 ( .A(n51719), .Z(n51720) );
  NAND U61280 ( .A(n51721), .B(n51722), .Z(n51680) );
  NAND U61281 ( .A(n51723), .B(n51724), .Z(n51722) );
  NANDN U61282 ( .A(n51725), .B(n51726), .Z(n51723) );
  NANDN U61283 ( .A(n51726), .B(n51725), .Z(n51721) );
  AND U61284 ( .A(n51727), .B(n51728), .Z(n51682) );
  NAND U61285 ( .A(n51729), .B(n51730), .Z(n51728) );
  OR U61286 ( .A(n51731), .B(n51732), .Z(n51729) );
  NANDN U61287 ( .A(n51733), .B(n51731), .Z(n51727) );
  XNOR U61288 ( .A(n51708), .B(n51734), .Z(N60814) );
  XOR U61289 ( .A(n51710), .B(n51711), .Z(n51734) );
  XNOR U61290 ( .A(n51724), .B(n51735), .Z(n51711) );
  XOR U61291 ( .A(n51725), .B(n51726), .Z(n51735) );
  XOR U61292 ( .A(n51731), .B(n51736), .Z(n51726) );
  XOR U61293 ( .A(n51730), .B(n51733), .Z(n51736) );
  IV U61294 ( .A(n51732), .Z(n51733) );
  NAND U61295 ( .A(n51737), .B(n51738), .Z(n51732) );
  OR U61296 ( .A(n51739), .B(n51740), .Z(n51738) );
  OR U61297 ( .A(n51741), .B(n51742), .Z(n51737) );
  NAND U61298 ( .A(n51743), .B(n51744), .Z(n51730) );
  OR U61299 ( .A(n51745), .B(n51746), .Z(n51744) );
  OR U61300 ( .A(n51747), .B(n51748), .Z(n51743) );
  NOR U61301 ( .A(n51749), .B(n51750), .Z(n51731) );
  ANDN U61302 ( .B(n51751), .A(n51752), .Z(n51725) );
  XNOR U61303 ( .A(n51718), .B(n51753), .Z(n51724) );
  XNOR U61304 ( .A(n51717), .B(n51719), .Z(n51753) );
  NAND U61305 ( .A(n51754), .B(n51755), .Z(n51719) );
  OR U61306 ( .A(n51756), .B(n51757), .Z(n51755) );
  OR U61307 ( .A(n51758), .B(n51759), .Z(n51754) );
  NAND U61308 ( .A(n51760), .B(n51761), .Z(n51717) );
  OR U61309 ( .A(n51762), .B(n51763), .Z(n51761) );
  OR U61310 ( .A(n51764), .B(n51765), .Z(n51760) );
  ANDN U61311 ( .B(n51766), .A(n51767), .Z(n51718) );
  IV U61312 ( .A(n51768), .Z(n51766) );
  ANDN U61313 ( .B(n51769), .A(n51770), .Z(n51710) );
  XOR U61314 ( .A(n51696), .B(n51771), .Z(n51708) );
  XOR U61315 ( .A(n51697), .B(n51698), .Z(n51771) );
  XOR U61316 ( .A(n51703), .B(n51772), .Z(n51698) );
  XOR U61317 ( .A(n51702), .B(n51705), .Z(n51772) );
  IV U61318 ( .A(n51704), .Z(n51705) );
  NAND U61319 ( .A(n51773), .B(n51774), .Z(n51704) );
  OR U61320 ( .A(n51775), .B(n51776), .Z(n51774) );
  OR U61321 ( .A(n51777), .B(n51778), .Z(n51773) );
  NAND U61322 ( .A(n51779), .B(n51780), .Z(n51702) );
  OR U61323 ( .A(n51781), .B(n51782), .Z(n51780) );
  OR U61324 ( .A(n51783), .B(n51784), .Z(n51779) );
  NOR U61325 ( .A(n51785), .B(n51786), .Z(n51703) );
  ANDN U61326 ( .B(n51787), .A(n51788), .Z(n51697) );
  IV U61327 ( .A(n51789), .Z(n51787) );
  XNOR U61328 ( .A(n51690), .B(n51790), .Z(n51696) );
  XNOR U61329 ( .A(n51689), .B(n51691), .Z(n51790) );
  NAND U61330 ( .A(n51791), .B(n51792), .Z(n51691) );
  OR U61331 ( .A(n51793), .B(n51794), .Z(n51792) );
  OR U61332 ( .A(n51795), .B(n51796), .Z(n51791) );
  NAND U61333 ( .A(n51797), .B(n51798), .Z(n51689) );
  OR U61334 ( .A(n51799), .B(n51800), .Z(n51798) );
  OR U61335 ( .A(n51801), .B(n51802), .Z(n51797) );
  ANDN U61336 ( .B(n51803), .A(n51804), .Z(n51690) );
  IV U61337 ( .A(n51805), .Z(n51803) );
  XNOR U61338 ( .A(n51770), .B(n51769), .Z(N60813) );
  XOR U61339 ( .A(n51789), .B(n51788), .Z(n51769) );
  XNOR U61340 ( .A(n51804), .B(n51805), .Z(n51788) );
  XNOR U61341 ( .A(n51799), .B(n51800), .Z(n51805) );
  XNOR U61342 ( .A(n51801), .B(n51802), .Z(n51800) );
  XNOR U61343 ( .A(y[421]), .B(x[421]), .Z(n51802) );
  XNOR U61344 ( .A(y[422]), .B(x[422]), .Z(n51801) );
  XNOR U61345 ( .A(y[420]), .B(x[420]), .Z(n51799) );
  XNOR U61346 ( .A(n51793), .B(n51794), .Z(n51804) );
  XNOR U61347 ( .A(y[417]), .B(x[417]), .Z(n51794) );
  XNOR U61348 ( .A(n51795), .B(n51796), .Z(n51793) );
  XNOR U61349 ( .A(y[418]), .B(x[418]), .Z(n51796) );
  XNOR U61350 ( .A(y[419]), .B(x[419]), .Z(n51795) );
  XNOR U61351 ( .A(n51786), .B(n51785), .Z(n51789) );
  XNOR U61352 ( .A(n51781), .B(n51782), .Z(n51785) );
  XNOR U61353 ( .A(y[414]), .B(x[414]), .Z(n51782) );
  XNOR U61354 ( .A(n51783), .B(n51784), .Z(n51781) );
  XNOR U61355 ( .A(y[415]), .B(x[415]), .Z(n51784) );
  XNOR U61356 ( .A(y[416]), .B(x[416]), .Z(n51783) );
  XNOR U61357 ( .A(n51775), .B(n51776), .Z(n51786) );
  XNOR U61358 ( .A(y[411]), .B(x[411]), .Z(n51776) );
  XNOR U61359 ( .A(n51777), .B(n51778), .Z(n51775) );
  XNOR U61360 ( .A(y[412]), .B(x[412]), .Z(n51778) );
  XNOR U61361 ( .A(y[413]), .B(x[413]), .Z(n51777) );
  XOR U61362 ( .A(n51751), .B(n51752), .Z(n51770) );
  XNOR U61363 ( .A(n51767), .B(n51768), .Z(n51752) );
  XNOR U61364 ( .A(n51762), .B(n51763), .Z(n51768) );
  XNOR U61365 ( .A(n51764), .B(n51765), .Z(n51763) );
  XNOR U61366 ( .A(y[409]), .B(x[409]), .Z(n51765) );
  XNOR U61367 ( .A(y[410]), .B(x[410]), .Z(n51764) );
  XNOR U61368 ( .A(y[408]), .B(x[408]), .Z(n51762) );
  XNOR U61369 ( .A(n51756), .B(n51757), .Z(n51767) );
  XNOR U61370 ( .A(y[405]), .B(x[405]), .Z(n51757) );
  XNOR U61371 ( .A(n51758), .B(n51759), .Z(n51756) );
  XNOR U61372 ( .A(y[406]), .B(x[406]), .Z(n51759) );
  XNOR U61373 ( .A(y[407]), .B(x[407]), .Z(n51758) );
  XOR U61374 ( .A(n51750), .B(n51749), .Z(n51751) );
  XNOR U61375 ( .A(n51745), .B(n51746), .Z(n51749) );
  XNOR U61376 ( .A(y[402]), .B(x[402]), .Z(n51746) );
  XNOR U61377 ( .A(n51747), .B(n51748), .Z(n51745) );
  XNOR U61378 ( .A(y[403]), .B(x[403]), .Z(n51748) );
  XNOR U61379 ( .A(y[404]), .B(x[404]), .Z(n51747) );
  XNOR U61380 ( .A(n51739), .B(n51740), .Z(n51750) );
  XNOR U61381 ( .A(y[399]), .B(x[399]), .Z(n51740) );
  XNOR U61382 ( .A(n51741), .B(n51742), .Z(n51739) );
  XNOR U61383 ( .A(y[400]), .B(x[400]), .Z(n51742) );
  XNOR U61384 ( .A(y[401]), .B(x[401]), .Z(n51741) );
  NAND U61385 ( .A(n51806), .B(n51807), .Z(N60804) );
  NANDN U61386 ( .A(n51808), .B(n51809), .Z(n51807) );
  OR U61387 ( .A(n51810), .B(n51811), .Z(n51809) );
  NAND U61388 ( .A(n51810), .B(n51811), .Z(n51806) );
  XOR U61389 ( .A(n51810), .B(n51812), .Z(N60803) );
  XNOR U61390 ( .A(n51808), .B(n51811), .Z(n51812) );
  AND U61391 ( .A(n51813), .B(n51814), .Z(n51811) );
  NANDN U61392 ( .A(n51815), .B(n51816), .Z(n51814) );
  NANDN U61393 ( .A(n51817), .B(n51818), .Z(n51816) );
  NANDN U61394 ( .A(n51818), .B(n51817), .Z(n51813) );
  NAND U61395 ( .A(n51819), .B(n51820), .Z(n51808) );
  NANDN U61396 ( .A(n51821), .B(n51822), .Z(n51820) );
  OR U61397 ( .A(n51823), .B(n51824), .Z(n51822) );
  NAND U61398 ( .A(n51824), .B(n51823), .Z(n51819) );
  AND U61399 ( .A(n51825), .B(n51826), .Z(n51810) );
  NANDN U61400 ( .A(n51827), .B(n51828), .Z(n51826) );
  NANDN U61401 ( .A(n51829), .B(n51830), .Z(n51828) );
  NANDN U61402 ( .A(n51830), .B(n51829), .Z(n51825) );
  XOR U61403 ( .A(n51824), .B(n51831), .Z(N60802) );
  XOR U61404 ( .A(n51821), .B(n51823), .Z(n51831) );
  XNOR U61405 ( .A(n51817), .B(n51832), .Z(n51823) );
  XNOR U61406 ( .A(n51815), .B(n51818), .Z(n51832) );
  NAND U61407 ( .A(n51833), .B(n51834), .Z(n51818) );
  NAND U61408 ( .A(n51835), .B(n51836), .Z(n51834) );
  OR U61409 ( .A(n51837), .B(n51838), .Z(n51835) );
  NANDN U61410 ( .A(n51839), .B(n51837), .Z(n51833) );
  IV U61411 ( .A(n51838), .Z(n51839) );
  NAND U61412 ( .A(n51840), .B(n51841), .Z(n51815) );
  NAND U61413 ( .A(n51842), .B(n51843), .Z(n51841) );
  NANDN U61414 ( .A(n51844), .B(n51845), .Z(n51842) );
  NANDN U61415 ( .A(n51845), .B(n51844), .Z(n51840) );
  AND U61416 ( .A(n51846), .B(n51847), .Z(n51817) );
  NAND U61417 ( .A(n51848), .B(n51849), .Z(n51847) );
  OR U61418 ( .A(n51850), .B(n51851), .Z(n51848) );
  NANDN U61419 ( .A(n51852), .B(n51850), .Z(n51846) );
  NAND U61420 ( .A(n51853), .B(n51854), .Z(n51821) );
  NANDN U61421 ( .A(n51855), .B(n51856), .Z(n51854) );
  OR U61422 ( .A(n51857), .B(n51858), .Z(n51856) );
  NANDN U61423 ( .A(n51859), .B(n51857), .Z(n51853) );
  IV U61424 ( .A(n51858), .Z(n51859) );
  XNOR U61425 ( .A(n51829), .B(n51860), .Z(n51824) );
  XNOR U61426 ( .A(n51827), .B(n51830), .Z(n51860) );
  NAND U61427 ( .A(n51861), .B(n51862), .Z(n51830) );
  NAND U61428 ( .A(n51863), .B(n51864), .Z(n51862) );
  OR U61429 ( .A(n51865), .B(n51866), .Z(n51863) );
  NANDN U61430 ( .A(n51867), .B(n51865), .Z(n51861) );
  IV U61431 ( .A(n51866), .Z(n51867) );
  NAND U61432 ( .A(n51868), .B(n51869), .Z(n51827) );
  NAND U61433 ( .A(n51870), .B(n51871), .Z(n51869) );
  NANDN U61434 ( .A(n51872), .B(n51873), .Z(n51870) );
  NANDN U61435 ( .A(n51873), .B(n51872), .Z(n51868) );
  AND U61436 ( .A(n51874), .B(n51875), .Z(n51829) );
  NAND U61437 ( .A(n51876), .B(n51877), .Z(n51875) );
  OR U61438 ( .A(n51878), .B(n51879), .Z(n51876) );
  NANDN U61439 ( .A(n51880), .B(n51878), .Z(n51874) );
  XNOR U61440 ( .A(n51855), .B(n51881), .Z(N60801) );
  XOR U61441 ( .A(n51857), .B(n51858), .Z(n51881) );
  XNOR U61442 ( .A(n51871), .B(n51882), .Z(n51858) );
  XOR U61443 ( .A(n51872), .B(n51873), .Z(n51882) );
  XOR U61444 ( .A(n51878), .B(n51883), .Z(n51873) );
  XOR U61445 ( .A(n51877), .B(n51880), .Z(n51883) );
  IV U61446 ( .A(n51879), .Z(n51880) );
  NAND U61447 ( .A(n51884), .B(n51885), .Z(n51879) );
  OR U61448 ( .A(n51886), .B(n51887), .Z(n51885) );
  OR U61449 ( .A(n51888), .B(n51889), .Z(n51884) );
  NAND U61450 ( .A(n51890), .B(n51891), .Z(n51877) );
  OR U61451 ( .A(n51892), .B(n51893), .Z(n51891) );
  OR U61452 ( .A(n51894), .B(n51895), .Z(n51890) );
  NOR U61453 ( .A(n51896), .B(n51897), .Z(n51878) );
  ANDN U61454 ( .B(n51898), .A(n51899), .Z(n51872) );
  XNOR U61455 ( .A(n51865), .B(n51900), .Z(n51871) );
  XNOR U61456 ( .A(n51864), .B(n51866), .Z(n51900) );
  NAND U61457 ( .A(n51901), .B(n51902), .Z(n51866) );
  OR U61458 ( .A(n51903), .B(n51904), .Z(n51902) );
  OR U61459 ( .A(n51905), .B(n51906), .Z(n51901) );
  NAND U61460 ( .A(n51907), .B(n51908), .Z(n51864) );
  OR U61461 ( .A(n51909), .B(n51910), .Z(n51908) );
  OR U61462 ( .A(n51911), .B(n51912), .Z(n51907) );
  ANDN U61463 ( .B(n51913), .A(n51914), .Z(n51865) );
  IV U61464 ( .A(n51915), .Z(n51913) );
  ANDN U61465 ( .B(n51916), .A(n51917), .Z(n51857) );
  XOR U61466 ( .A(n51843), .B(n51918), .Z(n51855) );
  XOR U61467 ( .A(n51844), .B(n51845), .Z(n51918) );
  XOR U61468 ( .A(n51850), .B(n51919), .Z(n51845) );
  XOR U61469 ( .A(n51849), .B(n51852), .Z(n51919) );
  IV U61470 ( .A(n51851), .Z(n51852) );
  NAND U61471 ( .A(n51920), .B(n51921), .Z(n51851) );
  OR U61472 ( .A(n51922), .B(n51923), .Z(n51921) );
  OR U61473 ( .A(n51924), .B(n51925), .Z(n51920) );
  NAND U61474 ( .A(n51926), .B(n51927), .Z(n51849) );
  OR U61475 ( .A(n51928), .B(n51929), .Z(n51927) );
  OR U61476 ( .A(n51930), .B(n51931), .Z(n51926) );
  NOR U61477 ( .A(n51932), .B(n51933), .Z(n51850) );
  ANDN U61478 ( .B(n51934), .A(n51935), .Z(n51844) );
  IV U61479 ( .A(n51936), .Z(n51934) );
  XNOR U61480 ( .A(n51837), .B(n51937), .Z(n51843) );
  XNOR U61481 ( .A(n51836), .B(n51838), .Z(n51937) );
  NAND U61482 ( .A(n51938), .B(n51939), .Z(n51838) );
  OR U61483 ( .A(n51940), .B(n51941), .Z(n51939) );
  OR U61484 ( .A(n51942), .B(n51943), .Z(n51938) );
  NAND U61485 ( .A(n51944), .B(n51945), .Z(n51836) );
  OR U61486 ( .A(n51946), .B(n51947), .Z(n51945) );
  OR U61487 ( .A(n51948), .B(n51949), .Z(n51944) );
  ANDN U61488 ( .B(n51950), .A(n51951), .Z(n51837) );
  IV U61489 ( .A(n51952), .Z(n51950) );
  XNOR U61490 ( .A(n51917), .B(n51916), .Z(N60800) );
  XOR U61491 ( .A(n51936), .B(n51935), .Z(n51916) );
  XNOR U61492 ( .A(n51951), .B(n51952), .Z(n51935) );
  XNOR U61493 ( .A(n51946), .B(n51947), .Z(n51952) );
  XNOR U61494 ( .A(n51948), .B(n51949), .Z(n51947) );
  XNOR U61495 ( .A(y[397]), .B(x[397]), .Z(n51949) );
  XNOR U61496 ( .A(y[398]), .B(x[398]), .Z(n51948) );
  XNOR U61497 ( .A(y[396]), .B(x[396]), .Z(n51946) );
  XNOR U61498 ( .A(n51940), .B(n51941), .Z(n51951) );
  XNOR U61499 ( .A(y[393]), .B(x[393]), .Z(n51941) );
  XNOR U61500 ( .A(n51942), .B(n51943), .Z(n51940) );
  XNOR U61501 ( .A(y[394]), .B(x[394]), .Z(n51943) );
  XNOR U61502 ( .A(y[395]), .B(x[395]), .Z(n51942) );
  XNOR U61503 ( .A(n51933), .B(n51932), .Z(n51936) );
  XNOR U61504 ( .A(n51928), .B(n51929), .Z(n51932) );
  XNOR U61505 ( .A(y[390]), .B(x[390]), .Z(n51929) );
  XNOR U61506 ( .A(n51930), .B(n51931), .Z(n51928) );
  XNOR U61507 ( .A(y[391]), .B(x[391]), .Z(n51931) );
  XNOR U61508 ( .A(y[392]), .B(x[392]), .Z(n51930) );
  XNOR U61509 ( .A(n51922), .B(n51923), .Z(n51933) );
  XNOR U61510 ( .A(y[387]), .B(x[387]), .Z(n51923) );
  XNOR U61511 ( .A(n51924), .B(n51925), .Z(n51922) );
  XNOR U61512 ( .A(y[388]), .B(x[388]), .Z(n51925) );
  XNOR U61513 ( .A(y[389]), .B(x[389]), .Z(n51924) );
  XOR U61514 ( .A(n51898), .B(n51899), .Z(n51917) );
  XNOR U61515 ( .A(n51914), .B(n51915), .Z(n51899) );
  XNOR U61516 ( .A(n51909), .B(n51910), .Z(n51915) );
  XNOR U61517 ( .A(n51911), .B(n51912), .Z(n51910) );
  XNOR U61518 ( .A(y[385]), .B(x[385]), .Z(n51912) );
  XNOR U61519 ( .A(y[386]), .B(x[386]), .Z(n51911) );
  XNOR U61520 ( .A(y[384]), .B(x[384]), .Z(n51909) );
  XNOR U61521 ( .A(n51903), .B(n51904), .Z(n51914) );
  XNOR U61522 ( .A(y[381]), .B(x[381]), .Z(n51904) );
  XNOR U61523 ( .A(n51905), .B(n51906), .Z(n51903) );
  XNOR U61524 ( .A(y[382]), .B(x[382]), .Z(n51906) );
  XNOR U61525 ( .A(y[383]), .B(x[383]), .Z(n51905) );
  XOR U61526 ( .A(n51897), .B(n51896), .Z(n51898) );
  XNOR U61527 ( .A(n51892), .B(n51893), .Z(n51896) );
  XNOR U61528 ( .A(y[378]), .B(x[378]), .Z(n51893) );
  XNOR U61529 ( .A(n51894), .B(n51895), .Z(n51892) );
  XNOR U61530 ( .A(y[379]), .B(x[379]), .Z(n51895) );
  XNOR U61531 ( .A(y[380]), .B(x[380]), .Z(n51894) );
  XNOR U61532 ( .A(n51886), .B(n51887), .Z(n51897) );
  XNOR U61533 ( .A(y[375]), .B(x[375]), .Z(n51887) );
  XNOR U61534 ( .A(n51888), .B(n51889), .Z(n51886) );
  XNOR U61535 ( .A(y[376]), .B(x[376]), .Z(n51889) );
  XNOR U61536 ( .A(y[377]), .B(x[377]), .Z(n51888) );
  NAND U61537 ( .A(n51953), .B(n51954), .Z(N60791) );
  NANDN U61538 ( .A(n51955), .B(n51956), .Z(n51954) );
  OR U61539 ( .A(n51957), .B(n51958), .Z(n51956) );
  NAND U61540 ( .A(n51957), .B(n51958), .Z(n51953) );
  XOR U61541 ( .A(n51957), .B(n51959), .Z(N60790) );
  XNOR U61542 ( .A(n51955), .B(n51958), .Z(n51959) );
  AND U61543 ( .A(n51960), .B(n51961), .Z(n51958) );
  NANDN U61544 ( .A(n51962), .B(n51963), .Z(n51961) );
  NANDN U61545 ( .A(n51964), .B(n51965), .Z(n51963) );
  NANDN U61546 ( .A(n51965), .B(n51964), .Z(n51960) );
  NAND U61547 ( .A(n51966), .B(n51967), .Z(n51955) );
  NANDN U61548 ( .A(n51968), .B(n51969), .Z(n51967) );
  OR U61549 ( .A(n51970), .B(n51971), .Z(n51969) );
  NAND U61550 ( .A(n51971), .B(n51970), .Z(n51966) );
  AND U61551 ( .A(n51972), .B(n51973), .Z(n51957) );
  NANDN U61552 ( .A(n51974), .B(n51975), .Z(n51973) );
  NANDN U61553 ( .A(n51976), .B(n51977), .Z(n51975) );
  NANDN U61554 ( .A(n51977), .B(n51976), .Z(n51972) );
  XOR U61555 ( .A(n51971), .B(n51978), .Z(N60789) );
  XOR U61556 ( .A(n51968), .B(n51970), .Z(n51978) );
  XNOR U61557 ( .A(n51964), .B(n51979), .Z(n51970) );
  XNOR U61558 ( .A(n51962), .B(n51965), .Z(n51979) );
  NAND U61559 ( .A(n51980), .B(n51981), .Z(n51965) );
  NAND U61560 ( .A(n51982), .B(n51983), .Z(n51981) );
  OR U61561 ( .A(n51984), .B(n51985), .Z(n51982) );
  NANDN U61562 ( .A(n51986), .B(n51984), .Z(n51980) );
  IV U61563 ( .A(n51985), .Z(n51986) );
  NAND U61564 ( .A(n51987), .B(n51988), .Z(n51962) );
  NAND U61565 ( .A(n51989), .B(n51990), .Z(n51988) );
  NANDN U61566 ( .A(n51991), .B(n51992), .Z(n51989) );
  NANDN U61567 ( .A(n51992), .B(n51991), .Z(n51987) );
  AND U61568 ( .A(n51993), .B(n51994), .Z(n51964) );
  NAND U61569 ( .A(n51995), .B(n51996), .Z(n51994) );
  OR U61570 ( .A(n51997), .B(n51998), .Z(n51995) );
  NANDN U61571 ( .A(n51999), .B(n51997), .Z(n51993) );
  NAND U61572 ( .A(n52000), .B(n52001), .Z(n51968) );
  NANDN U61573 ( .A(n52002), .B(n52003), .Z(n52001) );
  OR U61574 ( .A(n52004), .B(n52005), .Z(n52003) );
  NANDN U61575 ( .A(n52006), .B(n52004), .Z(n52000) );
  IV U61576 ( .A(n52005), .Z(n52006) );
  XNOR U61577 ( .A(n51976), .B(n52007), .Z(n51971) );
  XNOR U61578 ( .A(n51974), .B(n51977), .Z(n52007) );
  NAND U61579 ( .A(n52008), .B(n52009), .Z(n51977) );
  NAND U61580 ( .A(n52010), .B(n52011), .Z(n52009) );
  OR U61581 ( .A(n52012), .B(n52013), .Z(n52010) );
  NANDN U61582 ( .A(n52014), .B(n52012), .Z(n52008) );
  IV U61583 ( .A(n52013), .Z(n52014) );
  NAND U61584 ( .A(n52015), .B(n52016), .Z(n51974) );
  NAND U61585 ( .A(n52017), .B(n52018), .Z(n52016) );
  NANDN U61586 ( .A(n52019), .B(n52020), .Z(n52017) );
  NANDN U61587 ( .A(n52020), .B(n52019), .Z(n52015) );
  AND U61588 ( .A(n52021), .B(n52022), .Z(n51976) );
  NAND U61589 ( .A(n52023), .B(n52024), .Z(n52022) );
  OR U61590 ( .A(n52025), .B(n52026), .Z(n52023) );
  NANDN U61591 ( .A(n52027), .B(n52025), .Z(n52021) );
  XNOR U61592 ( .A(n52002), .B(n52028), .Z(N60788) );
  XOR U61593 ( .A(n52004), .B(n52005), .Z(n52028) );
  XNOR U61594 ( .A(n52018), .B(n52029), .Z(n52005) );
  XOR U61595 ( .A(n52019), .B(n52020), .Z(n52029) );
  XOR U61596 ( .A(n52025), .B(n52030), .Z(n52020) );
  XOR U61597 ( .A(n52024), .B(n52027), .Z(n52030) );
  IV U61598 ( .A(n52026), .Z(n52027) );
  NAND U61599 ( .A(n52031), .B(n52032), .Z(n52026) );
  OR U61600 ( .A(n52033), .B(n52034), .Z(n52032) );
  OR U61601 ( .A(n52035), .B(n52036), .Z(n52031) );
  NAND U61602 ( .A(n52037), .B(n52038), .Z(n52024) );
  OR U61603 ( .A(n52039), .B(n52040), .Z(n52038) );
  OR U61604 ( .A(n52041), .B(n52042), .Z(n52037) );
  NOR U61605 ( .A(n52043), .B(n52044), .Z(n52025) );
  ANDN U61606 ( .B(n52045), .A(n52046), .Z(n52019) );
  XNOR U61607 ( .A(n52012), .B(n52047), .Z(n52018) );
  XNOR U61608 ( .A(n52011), .B(n52013), .Z(n52047) );
  NAND U61609 ( .A(n52048), .B(n52049), .Z(n52013) );
  OR U61610 ( .A(n52050), .B(n52051), .Z(n52049) );
  OR U61611 ( .A(n52052), .B(n52053), .Z(n52048) );
  NAND U61612 ( .A(n52054), .B(n52055), .Z(n52011) );
  OR U61613 ( .A(n52056), .B(n52057), .Z(n52055) );
  OR U61614 ( .A(n52058), .B(n52059), .Z(n52054) );
  ANDN U61615 ( .B(n52060), .A(n52061), .Z(n52012) );
  IV U61616 ( .A(n52062), .Z(n52060) );
  ANDN U61617 ( .B(n52063), .A(n52064), .Z(n52004) );
  XOR U61618 ( .A(n51990), .B(n52065), .Z(n52002) );
  XOR U61619 ( .A(n51991), .B(n51992), .Z(n52065) );
  XOR U61620 ( .A(n51997), .B(n52066), .Z(n51992) );
  XOR U61621 ( .A(n51996), .B(n51999), .Z(n52066) );
  IV U61622 ( .A(n51998), .Z(n51999) );
  NAND U61623 ( .A(n52067), .B(n52068), .Z(n51998) );
  OR U61624 ( .A(n52069), .B(n52070), .Z(n52068) );
  OR U61625 ( .A(n52071), .B(n52072), .Z(n52067) );
  NAND U61626 ( .A(n52073), .B(n52074), .Z(n51996) );
  OR U61627 ( .A(n52075), .B(n52076), .Z(n52074) );
  OR U61628 ( .A(n52077), .B(n52078), .Z(n52073) );
  NOR U61629 ( .A(n52079), .B(n52080), .Z(n51997) );
  ANDN U61630 ( .B(n52081), .A(n52082), .Z(n51991) );
  IV U61631 ( .A(n52083), .Z(n52081) );
  XNOR U61632 ( .A(n51984), .B(n52084), .Z(n51990) );
  XNOR U61633 ( .A(n51983), .B(n51985), .Z(n52084) );
  NAND U61634 ( .A(n52085), .B(n52086), .Z(n51985) );
  OR U61635 ( .A(n52087), .B(n52088), .Z(n52086) );
  OR U61636 ( .A(n52089), .B(n52090), .Z(n52085) );
  NAND U61637 ( .A(n52091), .B(n52092), .Z(n51983) );
  OR U61638 ( .A(n52093), .B(n52094), .Z(n52092) );
  OR U61639 ( .A(n52095), .B(n52096), .Z(n52091) );
  ANDN U61640 ( .B(n52097), .A(n52098), .Z(n51984) );
  IV U61641 ( .A(n52099), .Z(n52097) );
  XNOR U61642 ( .A(n52064), .B(n52063), .Z(N60787) );
  XOR U61643 ( .A(n52083), .B(n52082), .Z(n52063) );
  XNOR U61644 ( .A(n52098), .B(n52099), .Z(n52082) );
  XNOR U61645 ( .A(n52093), .B(n52094), .Z(n52099) );
  XNOR U61646 ( .A(n52095), .B(n52096), .Z(n52094) );
  XNOR U61647 ( .A(y[373]), .B(x[373]), .Z(n52096) );
  XNOR U61648 ( .A(y[374]), .B(x[374]), .Z(n52095) );
  XNOR U61649 ( .A(y[372]), .B(x[372]), .Z(n52093) );
  XNOR U61650 ( .A(n52087), .B(n52088), .Z(n52098) );
  XNOR U61651 ( .A(y[369]), .B(x[369]), .Z(n52088) );
  XNOR U61652 ( .A(n52089), .B(n52090), .Z(n52087) );
  XNOR U61653 ( .A(y[370]), .B(x[370]), .Z(n52090) );
  XNOR U61654 ( .A(y[371]), .B(x[371]), .Z(n52089) );
  XNOR U61655 ( .A(n52080), .B(n52079), .Z(n52083) );
  XNOR U61656 ( .A(n52075), .B(n52076), .Z(n52079) );
  XNOR U61657 ( .A(y[366]), .B(x[366]), .Z(n52076) );
  XNOR U61658 ( .A(n52077), .B(n52078), .Z(n52075) );
  XNOR U61659 ( .A(y[367]), .B(x[367]), .Z(n52078) );
  XNOR U61660 ( .A(y[368]), .B(x[368]), .Z(n52077) );
  XNOR U61661 ( .A(n52069), .B(n52070), .Z(n52080) );
  XNOR U61662 ( .A(y[363]), .B(x[363]), .Z(n52070) );
  XNOR U61663 ( .A(n52071), .B(n52072), .Z(n52069) );
  XNOR U61664 ( .A(y[364]), .B(x[364]), .Z(n52072) );
  XNOR U61665 ( .A(y[365]), .B(x[365]), .Z(n52071) );
  XOR U61666 ( .A(n52045), .B(n52046), .Z(n52064) );
  XNOR U61667 ( .A(n52061), .B(n52062), .Z(n52046) );
  XNOR U61668 ( .A(n52056), .B(n52057), .Z(n52062) );
  XNOR U61669 ( .A(n52058), .B(n52059), .Z(n52057) );
  XNOR U61670 ( .A(y[361]), .B(x[361]), .Z(n52059) );
  XNOR U61671 ( .A(y[362]), .B(x[362]), .Z(n52058) );
  XNOR U61672 ( .A(y[360]), .B(x[360]), .Z(n52056) );
  XNOR U61673 ( .A(n52050), .B(n52051), .Z(n52061) );
  XNOR U61674 ( .A(y[357]), .B(x[357]), .Z(n52051) );
  XNOR U61675 ( .A(n52052), .B(n52053), .Z(n52050) );
  XNOR U61676 ( .A(y[358]), .B(x[358]), .Z(n52053) );
  XNOR U61677 ( .A(y[359]), .B(x[359]), .Z(n52052) );
  XOR U61678 ( .A(n52044), .B(n52043), .Z(n52045) );
  XNOR U61679 ( .A(n52039), .B(n52040), .Z(n52043) );
  XNOR U61680 ( .A(y[354]), .B(x[354]), .Z(n52040) );
  XNOR U61681 ( .A(n52041), .B(n52042), .Z(n52039) );
  XNOR U61682 ( .A(y[355]), .B(x[355]), .Z(n52042) );
  XNOR U61683 ( .A(y[356]), .B(x[356]), .Z(n52041) );
  XNOR U61684 ( .A(n52033), .B(n52034), .Z(n52044) );
  XNOR U61685 ( .A(y[351]), .B(x[351]), .Z(n52034) );
  XNOR U61686 ( .A(n52035), .B(n52036), .Z(n52033) );
  XNOR U61687 ( .A(y[352]), .B(x[352]), .Z(n52036) );
  XNOR U61688 ( .A(y[353]), .B(x[353]), .Z(n52035) );
  NAND U61689 ( .A(n52100), .B(n52101), .Z(N60778) );
  NANDN U61690 ( .A(n52102), .B(n52103), .Z(n52101) );
  OR U61691 ( .A(n52104), .B(n52105), .Z(n52103) );
  NAND U61692 ( .A(n52104), .B(n52105), .Z(n52100) );
  XOR U61693 ( .A(n52104), .B(n52106), .Z(N60777) );
  XNOR U61694 ( .A(n52102), .B(n52105), .Z(n52106) );
  AND U61695 ( .A(n52107), .B(n52108), .Z(n52105) );
  NANDN U61696 ( .A(n52109), .B(n52110), .Z(n52108) );
  NANDN U61697 ( .A(n52111), .B(n52112), .Z(n52110) );
  NANDN U61698 ( .A(n52112), .B(n52111), .Z(n52107) );
  NAND U61699 ( .A(n52113), .B(n52114), .Z(n52102) );
  NANDN U61700 ( .A(n52115), .B(n52116), .Z(n52114) );
  OR U61701 ( .A(n52117), .B(n52118), .Z(n52116) );
  NAND U61702 ( .A(n52118), .B(n52117), .Z(n52113) );
  AND U61703 ( .A(n52119), .B(n52120), .Z(n52104) );
  NANDN U61704 ( .A(n52121), .B(n52122), .Z(n52120) );
  NANDN U61705 ( .A(n52123), .B(n52124), .Z(n52122) );
  NANDN U61706 ( .A(n52124), .B(n52123), .Z(n52119) );
  XOR U61707 ( .A(n52118), .B(n52125), .Z(N60776) );
  XOR U61708 ( .A(n52115), .B(n52117), .Z(n52125) );
  XNOR U61709 ( .A(n52111), .B(n52126), .Z(n52117) );
  XNOR U61710 ( .A(n52109), .B(n52112), .Z(n52126) );
  NAND U61711 ( .A(n52127), .B(n52128), .Z(n52112) );
  NAND U61712 ( .A(n52129), .B(n52130), .Z(n52128) );
  OR U61713 ( .A(n52131), .B(n52132), .Z(n52129) );
  NANDN U61714 ( .A(n52133), .B(n52131), .Z(n52127) );
  IV U61715 ( .A(n52132), .Z(n52133) );
  NAND U61716 ( .A(n52134), .B(n52135), .Z(n52109) );
  NAND U61717 ( .A(n52136), .B(n52137), .Z(n52135) );
  NANDN U61718 ( .A(n52138), .B(n52139), .Z(n52136) );
  NANDN U61719 ( .A(n52139), .B(n52138), .Z(n52134) );
  AND U61720 ( .A(n52140), .B(n52141), .Z(n52111) );
  NAND U61721 ( .A(n52142), .B(n52143), .Z(n52141) );
  OR U61722 ( .A(n52144), .B(n52145), .Z(n52142) );
  NANDN U61723 ( .A(n52146), .B(n52144), .Z(n52140) );
  NAND U61724 ( .A(n52147), .B(n52148), .Z(n52115) );
  NANDN U61725 ( .A(n52149), .B(n52150), .Z(n52148) );
  OR U61726 ( .A(n52151), .B(n52152), .Z(n52150) );
  NANDN U61727 ( .A(n52153), .B(n52151), .Z(n52147) );
  IV U61728 ( .A(n52152), .Z(n52153) );
  XNOR U61729 ( .A(n52123), .B(n52154), .Z(n52118) );
  XNOR U61730 ( .A(n52121), .B(n52124), .Z(n52154) );
  NAND U61731 ( .A(n52155), .B(n52156), .Z(n52124) );
  NAND U61732 ( .A(n52157), .B(n52158), .Z(n52156) );
  OR U61733 ( .A(n52159), .B(n52160), .Z(n52157) );
  NANDN U61734 ( .A(n52161), .B(n52159), .Z(n52155) );
  IV U61735 ( .A(n52160), .Z(n52161) );
  NAND U61736 ( .A(n52162), .B(n52163), .Z(n52121) );
  NAND U61737 ( .A(n52164), .B(n52165), .Z(n52163) );
  NANDN U61738 ( .A(n52166), .B(n52167), .Z(n52164) );
  NANDN U61739 ( .A(n52167), .B(n52166), .Z(n52162) );
  AND U61740 ( .A(n52168), .B(n52169), .Z(n52123) );
  NAND U61741 ( .A(n52170), .B(n52171), .Z(n52169) );
  OR U61742 ( .A(n52172), .B(n52173), .Z(n52170) );
  NANDN U61743 ( .A(n52174), .B(n52172), .Z(n52168) );
  XNOR U61744 ( .A(n52149), .B(n52175), .Z(N60775) );
  XOR U61745 ( .A(n52151), .B(n52152), .Z(n52175) );
  XNOR U61746 ( .A(n52165), .B(n52176), .Z(n52152) );
  XOR U61747 ( .A(n52166), .B(n52167), .Z(n52176) );
  XOR U61748 ( .A(n52172), .B(n52177), .Z(n52167) );
  XOR U61749 ( .A(n52171), .B(n52174), .Z(n52177) );
  IV U61750 ( .A(n52173), .Z(n52174) );
  NAND U61751 ( .A(n52178), .B(n52179), .Z(n52173) );
  OR U61752 ( .A(n52180), .B(n52181), .Z(n52179) );
  OR U61753 ( .A(n52182), .B(n52183), .Z(n52178) );
  NAND U61754 ( .A(n52184), .B(n52185), .Z(n52171) );
  OR U61755 ( .A(n52186), .B(n52187), .Z(n52185) );
  OR U61756 ( .A(n52188), .B(n52189), .Z(n52184) );
  NOR U61757 ( .A(n52190), .B(n52191), .Z(n52172) );
  ANDN U61758 ( .B(n52192), .A(n52193), .Z(n52166) );
  XNOR U61759 ( .A(n52159), .B(n52194), .Z(n52165) );
  XNOR U61760 ( .A(n52158), .B(n52160), .Z(n52194) );
  NAND U61761 ( .A(n52195), .B(n52196), .Z(n52160) );
  OR U61762 ( .A(n52197), .B(n52198), .Z(n52196) );
  OR U61763 ( .A(n52199), .B(n52200), .Z(n52195) );
  NAND U61764 ( .A(n52201), .B(n52202), .Z(n52158) );
  OR U61765 ( .A(n52203), .B(n52204), .Z(n52202) );
  OR U61766 ( .A(n52205), .B(n52206), .Z(n52201) );
  ANDN U61767 ( .B(n52207), .A(n52208), .Z(n52159) );
  IV U61768 ( .A(n52209), .Z(n52207) );
  ANDN U61769 ( .B(n52210), .A(n52211), .Z(n52151) );
  XOR U61770 ( .A(n52137), .B(n52212), .Z(n52149) );
  XOR U61771 ( .A(n52138), .B(n52139), .Z(n52212) );
  XOR U61772 ( .A(n52144), .B(n52213), .Z(n52139) );
  XOR U61773 ( .A(n52143), .B(n52146), .Z(n52213) );
  IV U61774 ( .A(n52145), .Z(n52146) );
  NAND U61775 ( .A(n52214), .B(n52215), .Z(n52145) );
  OR U61776 ( .A(n52216), .B(n52217), .Z(n52215) );
  OR U61777 ( .A(n52218), .B(n52219), .Z(n52214) );
  NAND U61778 ( .A(n52220), .B(n52221), .Z(n52143) );
  OR U61779 ( .A(n52222), .B(n52223), .Z(n52221) );
  OR U61780 ( .A(n52224), .B(n52225), .Z(n52220) );
  NOR U61781 ( .A(n52226), .B(n52227), .Z(n52144) );
  ANDN U61782 ( .B(n52228), .A(n52229), .Z(n52138) );
  IV U61783 ( .A(n52230), .Z(n52228) );
  XNOR U61784 ( .A(n52131), .B(n52231), .Z(n52137) );
  XNOR U61785 ( .A(n52130), .B(n52132), .Z(n52231) );
  NAND U61786 ( .A(n52232), .B(n52233), .Z(n52132) );
  OR U61787 ( .A(n52234), .B(n52235), .Z(n52233) );
  OR U61788 ( .A(n52236), .B(n52237), .Z(n52232) );
  NAND U61789 ( .A(n52238), .B(n52239), .Z(n52130) );
  OR U61790 ( .A(n52240), .B(n52241), .Z(n52239) );
  OR U61791 ( .A(n52242), .B(n52243), .Z(n52238) );
  ANDN U61792 ( .B(n52244), .A(n52245), .Z(n52131) );
  IV U61793 ( .A(n52246), .Z(n52244) );
  XNOR U61794 ( .A(n52211), .B(n52210), .Z(N60774) );
  XOR U61795 ( .A(n52230), .B(n52229), .Z(n52210) );
  XNOR U61796 ( .A(n52245), .B(n52246), .Z(n52229) );
  XNOR U61797 ( .A(n52240), .B(n52241), .Z(n52246) );
  XNOR U61798 ( .A(n52242), .B(n52243), .Z(n52241) );
  XNOR U61799 ( .A(y[349]), .B(x[349]), .Z(n52243) );
  XNOR U61800 ( .A(y[350]), .B(x[350]), .Z(n52242) );
  XNOR U61801 ( .A(y[348]), .B(x[348]), .Z(n52240) );
  XNOR U61802 ( .A(n52234), .B(n52235), .Z(n52245) );
  XNOR U61803 ( .A(y[345]), .B(x[345]), .Z(n52235) );
  XNOR U61804 ( .A(n52236), .B(n52237), .Z(n52234) );
  XNOR U61805 ( .A(y[346]), .B(x[346]), .Z(n52237) );
  XNOR U61806 ( .A(y[347]), .B(x[347]), .Z(n52236) );
  XNOR U61807 ( .A(n52227), .B(n52226), .Z(n52230) );
  XNOR U61808 ( .A(n52222), .B(n52223), .Z(n52226) );
  XNOR U61809 ( .A(y[342]), .B(x[342]), .Z(n52223) );
  XNOR U61810 ( .A(n52224), .B(n52225), .Z(n52222) );
  XNOR U61811 ( .A(y[343]), .B(x[343]), .Z(n52225) );
  XNOR U61812 ( .A(y[344]), .B(x[344]), .Z(n52224) );
  XNOR U61813 ( .A(n52216), .B(n52217), .Z(n52227) );
  XNOR U61814 ( .A(y[339]), .B(x[339]), .Z(n52217) );
  XNOR U61815 ( .A(n52218), .B(n52219), .Z(n52216) );
  XNOR U61816 ( .A(y[340]), .B(x[340]), .Z(n52219) );
  XNOR U61817 ( .A(y[341]), .B(x[341]), .Z(n52218) );
  XOR U61818 ( .A(n52192), .B(n52193), .Z(n52211) );
  XNOR U61819 ( .A(n52208), .B(n52209), .Z(n52193) );
  XNOR U61820 ( .A(n52203), .B(n52204), .Z(n52209) );
  XNOR U61821 ( .A(n52205), .B(n52206), .Z(n52204) );
  XNOR U61822 ( .A(y[337]), .B(x[337]), .Z(n52206) );
  XNOR U61823 ( .A(y[338]), .B(x[338]), .Z(n52205) );
  XNOR U61824 ( .A(y[336]), .B(x[336]), .Z(n52203) );
  XNOR U61825 ( .A(n52197), .B(n52198), .Z(n52208) );
  XNOR U61826 ( .A(y[333]), .B(x[333]), .Z(n52198) );
  XNOR U61827 ( .A(n52199), .B(n52200), .Z(n52197) );
  XNOR U61828 ( .A(y[334]), .B(x[334]), .Z(n52200) );
  XNOR U61829 ( .A(y[335]), .B(x[335]), .Z(n52199) );
  XOR U61830 ( .A(n52191), .B(n52190), .Z(n52192) );
  XNOR U61831 ( .A(n52186), .B(n52187), .Z(n52190) );
  XNOR U61832 ( .A(y[330]), .B(x[330]), .Z(n52187) );
  XNOR U61833 ( .A(n52188), .B(n52189), .Z(n52186) );
  XNOR U61834 ( .A(y[331]), .B(x[331]), .Z(n52189) );
  XNOR U61835 ( .A(y[332]), .B(x[332]), .Z(n52188) );
  XNOR U61836 ( .A(n52180), .B(n52181), .Z(n52191) );
  XNOR U61837 ( .A(y[327]), .B(x[327]), .Z(n52181) );
  XNOR U61838 ( .A(n52182), .B(n52183), .Z(n52180) );
  XNOR U61839 ( .A(y[328]), .B(x[328]), .Z(n52183) );
  XNOR U61840 ( .A(y[329]), .B(x[329]), .Z(n52182) );
  NAND U61841 ( .A(n52247), .B(n52248), .Z(N60765) );
  NANDN U61842 ( .A(n52249), .B(n52250), .Z(n52248) );
  OR U61843 ( .A(n52251), .B(n52252), .Z(n52250) );
  NAND U61844 ( .A(n52251), .B(n52252), .Z(n52247) );
  XOR U61845 ( .A(n52251), .B(n52253), .Z(N60764) );
  XNOR U61846 ( .A(n52249), .B(n52252), .Z(n52253) );
  AND U61847 ( .A(n52254), .B(n52255), .Z(n52252) );
  NANDN U61848 ( .A(n52256), .B(n52257), .Z(n52255) );
  NANDN U61849 ( .A(n52258), .B(n52259), .Z(n52257) );
  NANDN U61850 ( .A(n52259), .B(n52258), .Z(n52254) );
  NAND U61851 ( .A(n52260), .B(n52261), .Z(n52249) );
  NANDN U61852 ( .A(n52262), .B(n52263), .Z(n52261) );
  OR U61853 ( .A(n52264), .B(n52265), .Z(n52263) );
  NAND U61854 ( .A(n52265), .B(n52264), .Z(n52260) );
  AND U61855 ( .A(n52266), .B(n52267), .Z(n52251) );
  NANDN U61856 ( .A(n52268), .B(n52269), .Z(n52267) );
  NANDN U61857 ( .A(n52270), .B(n52271), .Z(n52269) );
  NANDN U61858 ( .A(n52271), .B(n52270), .Z(n52266) );
  XOR U61859 ( .A(n52265), .B(n52272), .Z(N60763) );
  XOR U61860 ( .A(n52262), .B(n52264), .Z(n52272) );
  XNOR U61861 ( .A(n52258), .B(n52273), .Z(n52264) );
  XNOR U61862 ( .A(n52256), .B(n52259), .Z(n52273) );
  NAND U61863 ( .A(n52274), .B(n52275), .Z(n52259) );
  NAND U61864 ( .A(n52276), .B(n52277), .Z(n52275) );
  OR U61865 ( .A(n52278), .B(n52279), .Z(n52276) );
  NANDN U61866 ( .A(n52280), .B(n52278), .Z(n52274) );
  IV U61867 ( .A(n52279), .Z(n52280) );
  NAND U61868 ( .A(n52281), .B(n52282), .Z(n52256) );
  NAND U61869 ( .A(n52283), .B(n52284), .Z(n52282) );
  NANDN U61870 ( .A(n52285), .B(n52286), .Z(n52283) );
  NANDN U61871 ( .A(n52286), .B(n52285), .Z(n52281) );
  AND U61872 ( .A(n52287), .B(n52288), .Z(n52258) );
  NAND U61873 ( .A(n52289), .B(n52290), .Z(n52288) );
  OR U61874 ( .A(n52291), .B(n52292), .Z(n52289) );
  NANDN U61875 ( .A(n52293), .B(n52291), .Z(n52287) );
  NAND U61876 ( .A(n52294), .B(n52295), .Z(n52262) );
  NANDN U61877 ( .A(n52296), .B(n52297), .Z(n52295) );
  OR U61878 ( .A(n52298), .B(n52299), .Z(n52297) );
  NANDN U61879 ( .A(n52300), .B(n52298), .Z(n52294) );
  IV U61880 ( .A(n52299), .Z(n52300) );
  XNOR U61881 ( .A(n52270), .B(n52301), .Z(n52265) );
  XNOR U61882 ( .A(n52268), .B(n52271), .Z(n52301) );
  NAND U61883 ( .A(n52302), .B(n52303), .Z(n52271) );
  NAND U61884 ( .A(n52304), .B(n52305), .Z(n52303) );
  OR U61885 ( .A(n52306), .B(n52307), .Z(n52304) );
  NANDN U61886 ( .A(n52308), .B(n52306), .Z(n52302) );
  IV U61887 ( .A(n52307), .Z(n52308) );
  NAND U61888 ( .A(n52309), .B(n52310), .Z(n52268) );
  NAND U61889 ( .A(n52311), .B(n52312), .Z(n52310) );
  NANDN U61890 ( .A(n52313), .B(n52314), .Z(n52311) );
  NANDN U61891 ( .A(n52314), .B(n52313), .Z(n52309) );
  AND U61892 ( .A(n52315), .B(n52316), .Z(n52270) );
  NAND U61893 ( .A(n52317), .B(n52318), .Z(n52316) );
  OR U61894 ( .A(n52319), .B(n52320), .Z(n52317) );
  NANDN U61895 ( .A(n52321), .B(n52319), .Z(n52315) );
  XNOR U61896 ( .A(n52296), .B(n52322), .Z(N60762) );
  XOR U61897 ( .A(n52298), .B(n52299), .Z(n52322) );
  XNOR U61898 ( .A(n52312), .B(n52323), .Z(n52299) );
  XOR U61899 ( .A(n52313), .B(n52314), .Z(n52323) );
  XOR U61900 ( .A(n52319), .B(n52324), .Z(n52314) );
  XOR U61901 ( .A(n52318), .B(n52321), .Z(n52324) );
  IV U61902 ( .A(n52320), .Z(n52321) );
  NAND U61903 ( .A(n52325), .B(n52326), .Z(n52320) );
  OR U61904 ( .A(n52327), .B(n52328), .Z(n52326) );
  OR U61905 ( .A(n52329), .B(n52330), .Z(n52325) );
  NAND U61906 ( .A(n52331), .B(n52332), .Z(n52318) );
  OR U61907 ( .A(n52333), .B(n52334), .Z(n52332) );
  OR U61908 ( .A(n52335), .B(n52336), .Z(n52331) );
  NOR U61909 ( .A(n52337), .B(n52338), .Z(n52319) );
  ANDN U61910 ( .B(n52339), .A(n52340), .Z(n52313) );
  XNOR U61911 ( .A(n52306), .B(n52341), .Z(n52312) );
  XNOR U61912 ( .A(n52305), .B(n52307), .Z(n52341) );
  NAND U61913 ( .A(n52342), .B(n52343), .Z(n52307) );
  OR U61914 ( .A(n52344), .B(n52345), .Z(n52343) );
  OR U61915 ( .A(n52346), .B(n52347), .Z(n52342) );
  NAND U61916 ( .A(n52348), .B(n52349), .Z(n52305) );
  OR U61917 ( .A(n52350), .B(n52351), .Z(n52349) );
  OR U61918 ( .A(n52352), .B(n52353), .Z(n52348) );
  ANDN U61919 ( .B(n52354), .A(n52355), .Z(n52306) );
  IV U61920 ( .A(n52356), .Z(n52354) );
  ANDN U61921 ( .B(n52357), .A(n52358), .Z(n52298) );
  XOR U61922 ( .A(n52284), .B(n52359), .Z(n52296) );
  XOR U61923 ( .A(n52285), .B(n52286), .Z(n52359) );
  XOR U61924 ( .A(n52291), .B(n52360), .Z(n52286) );
  XOR U61925 ( .A(n52290), .B(n52293), .Z(n52360) );
  IV U61926 ( .A(n52292), .Z(n52293) );
  NAND U61927 ( .A(n52361), .B(n52362), .Z(n52292) );
  OR U61928 ( .A(n52363), .B(n52364), .Z(n52362) );
  OR U61929 ( .A(n52365), .B(n52366), .Z(n52361) );
  NAND U61930 ( .A(n52367), .B(n52368), .Z(n52290) );
  OR U61931 ( .A(n52369), .B(n52370), .Z(n52368) );
  OR U61932 ( .A(n52371), .B(n52372), .Z(n52367) );
  NOR U61933 ( .A(n52373), .B(n52374), .Z(n52291) );
  ANDN U61934 ( .B(n52375), .A(n52376), .Z(n52285) );
  IV U61935 ( .A(n52377), .Z(n52375) );
  XNOR U61936 ( .A(n52278), .B(n52378), .Z(n52284) );
  XNOR U61937 ( .A(n52277), .B(n52279), .Z(n52378) );
  NAND U61938 ( .A(n52379), .B(n52380), .Z(n52279) );
  OR U61939 ( .A(n52381), .B(n52382), .Z(n52380) );
  OR U61940 ( .A(n52383), .B(n52384), .Z(n52379) );
  NAND U61941 ( .A(n52385), .B(n52386), .Z(n52277) );
  OR U61942 ( .A(n52387), .B(n52388), .Z(n52386) );
  OR U61943 ( .A(n52389), .B(n52390), .Z(n52385) );
  ANDN U61944 ( .B(n52391), .A(n52392), .Z(n52278) );
  IV U61945 ( .A(n52393), .Z(n52391) );
  XNOR U61946 ( .A(n52358), .B(n52357), .Z(N60761) );
  XOR U61947 ( .A(n52377), .B(n52376), .Z(n52357) );
  XNOR U61948 ( .A(n52392), .B(n52393), .Z(n52376) );
  XNOR U61949 ( .A(n52387), .B(n52388), .Z(n52393) );
  XNOR U61950 ( .A(n52389), .B(n52390), .Z(n52388) );
  XNOR U61951 ( .A(y[325]), .B(x[325]), .Z(n52390) );
  XNOR U61952 ( .A(y[326]), .B(x[326]), .Z(n52389) );
  XNOR U61953 ( .A(y[324]), .B(x[324]), .Z(n52387) );
  XNOR U61954 ( .A(n52381), .B(n52382), .Z(n52392) );
  XNOR U61955 ( .A(y[321]), .B(x[321]), .Z(n52382) );
  XNOR U61956 ( .A(n52383), .B(n52384), .Z(n52381) );
  XNOR U61957 ( .A(y[322]), .B(x[322]), .Z(n52384) );
  XNOR U61958 ( .A(y[323]), .B(x[323]), .Z(n52383) );
  XNOR U61959 ( .A(n52374), .B(n52373), .Z(n52377) );
  XNOR U61960 ( .A(n52369), .B(n52370), .Z(n52373) );
  XNOR U61961 ( .A(y[318]), .B(x[318]), .Z(n52370) );
  XNOR U61962 ( .A(n52371), .B(n52372), .Z(n52369) );
  XNOR U61963 ( .A(y[319]), .B(x[319]), .Z(n52372) );
  XNOR U61964 ( .A(y[320]), .B(x[320]), .Z(n52371) );
  XNOR U61965 ( .A(n52363), .B(n52364), .Z(n52374) );
  XNOR U61966 ( .A(y[315]), .B(x[315]), .Z(n52364) );
  XNOR U61967 ( .A(n52365), .B(n52366), .Z(n52363) );
  XNOR U61968 ( .A(y[316]), .B(x[316]), .Z(n52366) );
  XNOR U61969 ( .A(y[317]), .B(x[317]), .Z(n52365) );
  XOR U61970 ( .A(n52339), .B(n52340), .Z(n52358) );
  XNOR U61971 ( .A(n52355), .B(n52356), .Z(n52340) );
  XNOR U61972 ( .A(n52350), .B(n52351), .Z(n52356) );
  XNOR U61973 ( .A(n52352), .B(n52353), .Z(n52351) );
  XNOR U61974 ( .A(y[313]), .B(x[313]), .Z(n52353) );
  XNOR U61975 ( .A(y[314]), .B(x[314]), .Z(n52352) );
  XNOR U61976 ( .A(y[312]), .B(x[312]), .Z(n52350) );
  XNOR U61977 ( .A(n52344), .B(n52345), .Z(n52355) );
  XNOR U61978 ( .A(y[309]), .B(x[309]), .Z(n52345) );
  XNOR U61979 ( .A(n52346), .B(n52347), .Z(n52344) );
  XNOR U61980 ( .A(y[310]), .B(x[310]), .Z(n52347) );
  XNOR U61981 ( .A(y[311]), .B(x[311]), .Z(n52346) );
  XOR U61982 ( .A(n52338), .B(n52337), .Z(n52339) );
  XNOR U61983 ( .A(n52333), .B(n52334), .Z(n52337) );
  XNOR U61984 ( .A(y[306]), .B(x[306]), .Z(n52334) );
  XNOR U61985 ( .A(n52335), .B(n52336), .Z(n52333) );
  XNOR U61986 ( .A(y[307]), .B(x[307]), .Z(n52336) );
  XNOR U61987 ( .A(y[308]), .B(x[308]), .Z(n52335) );
  XNOR U61988 ( .A(n52327), .B(n52328), .Z(n52338) );
  XNOR U61989 ( .A(y[303]), .B(x[303]), .Z(n52328) );
  XNOR U61990 ( .A(n52329), .B(n52330), .Z(n52327) );
  XNOR U61991 ( .A(y[304]), .B(x[304]), .Z(n52330) );
  XNOR U61992 ( .A(y[305]), .B(x[305]), .Z(n52329) );
  NAND U61993 ( .A(n52394), .B(n52395), .Z(N60752) );
  NANDN U61994 ( .A(n52396), .B(n52397), .Z(n52395) );
  OR U61995 ( .A(n52398), .B(n52399), .Z(n52397) );
  NAND U61996 ( .A(n52398), .B(n52399), .Z(n52394) );
  XOR U61997 ( .A(n52398), .B(n52400), .Z(N60751) );
  XNOR U61998 ( .A(n52396), .B(n52399), .Z(n52400) );
  AND U61999 ( .A(n52401), .B(n52402), .Z(n52399) );
  NANDN U62000 ( .A(n52403), .B(n52404), .Z(n52402) );
  NANDN U62001 ( .A(n52405), .B(n52406), .Z(n52404) );
  NANDN U62002 ( .A(n52406), .B(n52405), .Z(n52401) );
  NAND U62003 ( .A(n52407), .B(n52408), .Z(n52396) );
  NANDN U62004 ( .A(n52409), .B(n52410), .Z(n52408) );
  OR U62005 ( .A(n52411), .B(n52412), .Z(n52410) );
  NAND U62006 ( .A(n52412), .B(n52411), .Z(n52407) );
  AND U62007 ( .A(n52413), .B(n52414), .Z(n52398) );
  NANDN U62008 ( .A(n52415), .B(n52416), .Z(n52414) );
  NANDN U62009 ( .A(n52417), .B(n52418), .Z(n52416) );
  NANDN U62010 ( .A(n52418), .B(n52417), .Z(n52413) );
  XOR U62011 ( .A(n52412), .B(n52419), .Z(N60750) );
  XOR U62012 ( .A(n52409), .B(n52411), .Z(n52419) );
  XNOR U62013 ( .A(n52405), .B(n52420), .Z(n52411) );
  XNOR U62014 ( .A(n52403), .B(n52406), .Z(n52420) );
  NAND U62015 ( .A(n52421), .B(n52422), .Z(n52406) );
  NAND U62016 ( .A(n52423), .B(n52424), .Z(n52422) );
  OR U62017 ( .A(n52425), .B(n52426), .Z(n52423) );
  NANDN U62018 ( .A(n52427), .B(n52425), .Z(n52421) );
  IV U62019 ( .A(n52426), .Z(n52427) );
  NAND U62020 ( .A(n52428), .B(n52429), .Z(n52403) );
  NAND U62021 ( .A(n52430), .B(n52431), .Z(n52429) );
  NANDN U62022 ( .A(n52432), .B(n52433), .Z(n52430) );
  NANDN U62023 ( .A(n52433), .B(n52432), .Z(n52428) );
  AND U62024 ( .A(n52434), .B(n52435), .Z(n52405) );
  NAND U62025 ( .A(n52436), .B(n52437), .Z(n52435) );
  OR U62026 ( .A(n52438), .B(n52439), .Z(n52436) );
  NANDN U62027 ( .A(n52440), .B(n52438), .Z(n52434) );
  NAND U62028 ( .A(n52441), .B(n52442), .Z(n52409) );
  NANDN U62029 ( .A(n52443), .B(n52444), .Z(n52442) );
  OR U62030 ( .A(n52445), .B(n52446), .Z(n52444) );
  NANDN U62031 ( .A(n52447), .B(n52445), .Z(n52441) );
  IV U62032 ( .A(n52446), .Z(n52447) );
  XNOR U62033 ( .A(n52417), .B(n52448), .Z(n52412) );
  XNOR U62034 ( .A(n52415), .B(n52418), .Z(n52448) );
  NAND U62035 ( .A(n52449), .B(n52450), .Z(n52418) );
  NAND U62036 ( .A(n52451), .B(n52452), .Z(n52450) );
  OR U62037 ( .A(n52453), .B(n52454), .Z(n52451) );
  NANDN U62038 ( .A(n52455), .B(n52453), .Z(n52449) );
  IV U62039 ( .A(n52454), .Z(n52455) );
  NAND U62040 ( .A(n52456), .B(n52457), .Z(n52415) );
  NAND U62041 ( .A(n52458), .B(n52459), .Z(n52457) );
  NANDN U62042 ( .A(n52460), .B(n52461), .Z(n52458) );
  NANDN U62043 ( .A(n52461), .B(n52460), .Z(n52456) );
  AND U62044 ( .A(n52462), .B(n52463), .Z(n52417) );
  NAND U62045 ( .A(n52464), .B(n52465), .Z(n52463) );
  OR U62046 ( .A(n52466), .B(n52467), .Z(n52464) );
  NANDN U62047 ( .A(n52468), .B(n52466), .Z(n52462) );
  XNOR U62048 ( .A(n52443), .B(n52469), .Z(N60749) );
  XOR U62049 ( .A(n52445), .B(n52446), .Z(n52469) );
  XNOR U62050 ( .A(n52459), .B(n52470), .Z(n52446) );
  XOR U62051 ( .A(n52460), .B(n52461), .Z(n52470) );
  XOR U62052 ( .A(n52466), .B(n52471), .Z(n52461) );
  XOR U62053 ( .A(n52465), .B(n52468), .Z(n52471) );
  IV U62054 ( .A(n52467), .Z(n52468) );
  NAND U62055 ( .A(n52472), .B(n52473), .Z(n52467) );
  OR U62056 ( .A(n52474), .B(n52475), .Z(n52473) );
  OR U62057 ( .A(n52476), .B(n52477), .Z(n52472) );
  NAND U62058 ( .A(n52478), .B(n52479), .Z(n52465) );
  OR U62059 ( .A(n52480), .B(n52481), .Z(n52479) );
  OR U62060 ( .A(n52482), .B(n52483), .Z(n52478) );
  NOR U62061 ( .A(n52484), .B(n52485), .Z(n52466) );
  ANDN U62062 ( .B(n52486), .A(n52487), .Z(n52460) );
  XNOR U62063 ( .A(n52453), .B(n52488), .Z(n52459) );
  XNOR U62064 ( .A(n52452), .B(n52454), .Z(n52488) );
  NAND U62065 ( .A(n52489), .B(n52490), .Z(n52454) );
  OR U62066 ( .A(n52491), .B(n52492), .Z(n52490) );
  OR U62067 ( .A(n52493), .B(n52494), .Z(n52489) );
  NAND U62068 ( .A(n52495), .B(n52496), .Z(n52452) );
  OR U62069 ( .A(n52497), .B(n52498), .Z(n52496) );
  OR U62070 ( .A(n52499), .B(n52500), .Z(n52495) );
  ANDN U62071 ( .B(n52501), .A(n52502), .Z(n52453) );
  IV U62072 ( .A(n52503), .Z(n52501) );
  ANDN U62073 ( .B(n52504), .A(n52505), .Z(n52445) );
  XOR U62074 ( .A(n52431), .B(n52506), .Z(n52443) );
  XOR U62075 ( .A(n52432), .B(n52433), .Z(n52506) );
  XOR U62076 ( .A(n52438), .B(n52507), .Z(n52433) );
  XOR U62077 ( .A(n52437), .B(n52440), .Z(n52507) );
  IV U62078 ( .A(n52439), .Z(n52440) );
  NAND U62079 ( .A(n52508), .B(n52509), .Z(n52439) );
  OR U62080 ( .A(n52510), .B(n52511), .Z(n52509) );
  OR U62081 ( .A(n52512), .B(n52513), .Z(n52508) );
  NAND U62082 ( .A(n52514), .B(n52515), .Z(n52437) );
  OR U62083 ( .A(n52516), .B(n52517), .Z(n52515) );
  OR U62084 ( .A(n52518), .B(n52519), .Z(n52514) );
  NOR U62085 ( .A(n52520), .B(n52521), .Z(n52438) );
  ANDN U62086 ( .B(n52522), .A(n52523), .Z(n52432) );
  IV U62087 ( .A(n52524), .Z(n52522) );
  XNOR U62088 ( .A(n52425), .B(n52525), .Z(n52431) );
  XNOR U62089 ( .A(n52424), .B(n52426), .Z(n52525) );
  NAND U62090 ( .A(n52526), .B(n52527), .Z(n52426) );
  OR U62091 ( .A(n52528), .B(n52529), .Z(n52527) );
  OR U62092 ( .A(n52530), .B(n52531), .Z(n52526) );
  NAND U62093 ( .A(n52532), .B(n52533), .Z(n52424) );
  OR U62094 ( .A(n52534), .B(n52535), .Z(n52533) );
  OR U62095 ( .A(n52536), .B(n52537), .Z(n52532) );
  ANDN U62096 ( .B(n52538), .A(n52539), .Z(n52425) );
  IV U62097 ( .A(n52540), .Z(n52538) );
  XNOR U62098 ( .A(n52505), .B(n52504), .Z(N60748) );
  XOR U62099 ( .A(n52524), .B(n52523), .Z(n52504) );
  XNOR U62100 ( .A(n52539), .B(n52540), .Z(n52523) );
  XNOR U62101 ( .A(n52534), .B(n52535), .Z(n52540) );
  XNOR U62102 ( .A(n52536), .B(n52537), .Z(n52535) );
  XNOR U62103 ( .A(y[301]), .B(x[301]), .Z(n52537) );
  XNOR U62104 ( .A(y[302]), .B(x[302]), .Z(n52536) );
  XNOR U62105 ( .A(y[300]), .B(x[300]), .Z(n52534) );
  XNOR U62106 ( .A(n52528), .B(n52529), .Z(n52539) );
  XNOR U62107 ( .A(y[297]), .B(x[297]), .Z(n52529) );
  XNOR U62108 ( .A(n52530), .B(n52531), .Z(n52528) );
  XNOR U62109 ( .A(y[298]), .B(x[298]), .Z(n52531) );
  XNOR U62110 ( .A(y[299]), .B(x[299]), .Z(n52530) );
  XNOR U62111 ( .A(n52521), .B(n52520), .Z(n52524) );
  XNOR U62112 ( .A(n52516), .B(n52517), .Z(n52520) );
  XNOR U62113 ( .A(y[294]), .B(x[294]), .Z(n52517) );
  XNOR U62114 ( .A(n52518), .B(n52519), .Z(n52516) );
  XNOR U62115 ( .A(y[295]), .B(x[295]), .Z(n52519) );
  XNOR U62116 ( .A(y[296]), .B(x[296]), .Z(n52518) );
  XNOR U62117 ( .A(n52510), .B(n52511), .Z(n52521) );
  XNOR U62118 ( .A(y[291]), .B(x[291]), .Z(n52511) );
  XNOR U62119 ( .A(n52512), .B(n52513), .Z(n52510) );
  XNOR U62120 ( .A(y[292]), .B(x[292]), .Z(n52513) );
  XNOR U62121 ( .A(y[293]), .B(x[293]), .Z(n52512) );
  XOR U62122 ( .A(n52486), .B(n52487), .Z(n52505) );
  XNOR U62123 ( .A(n52502), .B(n52503), .Z(n52487) );
  XNOR U62124 ( .A(n52497), .B(n52498), .Z(n52503) );
  XNOR U62125 ( .A(n52499), .B(n52500), .Z(n52498) );
  XNOR U62126 ( .A(y[289]), .B(x[289]), .Z(n52500) );
  XNOR U62127 ( .A(y[290]), .B(x[290]), .Z(n52499) );
  XNOR U62128 ( .A(y[288]), .B(x[288]), .Z(n52497) );
  XNOR U62129 ( .A(n52491), .B(n52492), .Z(n52502) );
  XNOR U62130 ( .A(y[285]), .B(x[285]), .Z(n52492) );
  XNOR U62131 ( .A(n52493), .B(n52494), .Z(n52491) );
  XNOR U62132 ( .A(y[286]), .B(x[286]), .Z(n52494) );
  XNOR U62133 ( .A(y[287]), .B(x[287]), .Z(n52493) );
  XOR U62134 ( .A(n52485), .B(n52484), .Z(n52486) );
  XNOR U62135 ( .A(n52480), .B(n52481), .Z(n52484) );
  XNOR U62136 ( .A(y[282]), .B(x[282]), .Z(n52481) );
  XNOR U62137 ( .A(n52482), .B(n52483), .Z(n52480) );
  XNOR U62138 ( .A(y[283]), .B(x[283]), .Z(n52483) );
  XNOR U62139 ( .A(y[284]), .B(x[284]), .Z(n52482) );
  XNOR U62140 ( .A(n52474), .B(n52475), .Z(n52485) );
  XNOR U62141 ( .A(y[279]), .B(x[279]), .Z(n52475) );
  XNOR U62142 ( .A(n52476), .B(n52477), .Z(n52474) );
  XNOR U62143 ( .A(y[280]), .B(x[280]), .Z(n52477) );
  XNOR U62144 ( .A(y[281]), .B(x[281]), .Z(n52476) );
  NAND U62145 ( .A(n52541), .B(n52542), .Z(N60739) );
  NANDN U62146 ( .A(n52543), .B(n52544), .Z(n52542) );
  OR U62147 ( .A(n52545), .B(n52546), .Z(n52544) );
  NAND U62148 ( .A(n52545), .B(n52546), .Z(n52541) );
  XOR U62149 ( .A(n52545), .B(n52547), .Z(N60738) );
  XNOR U62150 ( .A(n52543), .B(n52546), .Z(n52547) );
  AND U62151 ( .A(n52548), .B(n52549), .Z(n52546) );
  NANDN U62152 ( .A(n52550), .B(n52551), .Z(n52549) );
  NANDN U62153 ( .A(n52552), .B(n52553), .Z(n52551) );
  NANDN U62154 ( .A(n52553), .B(n52552), .Z(n52548) );
  NAND U62155 ( .A(n52554), .B(n52555), .Z(n52543) );
  NANDN U62156 ( .A(n52556), .B(n52557), .Z(n52555) );
  OR U62157 ( .A(n52558), .B(n52559), .Z(n52557) );
  NAND U62158 ( .A(n52559), .B(n52558), .Z(n52554) );
  AND U62159 ( .A(n52560), .B(n52561), .Z(n52545) );
  NANDN U62160 ( .A(n52562), .B(n52563), .Z(n52561) );
  NANDN U62161 ( .A(n52564), .B(n52565), .Z(n52563) );
  NANDN U62162 ( .A(n52565), .B(n52564), .Z(n52560) );
  XOR U62163 ( .A(n52559), .B(n52566), .Z(N60737) );
  XOR U62164 ( .A(n52556), .B(n52558), .Z(n52566) );
  XNOR U62165 ( .A(n52552), .B(n52567), .Z(n52558) );
  XNOR U62166 ( .A(n52550), .B(n52553), .Z(n52567) );
  NAND U62167 ( .A(n52568), .B(n52569), .Z(n52553) );
  NAND U62168 ( .A(n52570), .B(n52571), .Z(n52569) );
  OR U62169 ( .A(n52572), .B(n52573), .Z(n52570) );
  NANDN U62170 ( .A(n52574), .B(n52572), .Z(n52568) );
  IV U62171 ( .A(n52573), .Z(n52574) );
  NAND U62172 ( .A(n52575), .B(n52576), .Z(n52550) );
  NAND U62173 ( .A(n52577), .B(n52578), .Z(n52576) );
  NANDN U62174 ( .A(n52579), .B(n52580), .Z(n52577) );
  NANDN U62175 ( .A(n52580), .B(n52579), .Z(n52575) );
  AND U62176 ( .A(n52581), .B(n52582), .Z(n52552) );
  NAND U62177 ( .A(n52583), .B(n52584), .Z(n52582) );
  OR U62178 ( .A(n52585), .B(n52586), .Z(n52583) );
  NANDN U62179 ( .A(n52587), .B(n52585), .Z(n52581) );
  NAND U62180 ( .A(n52588), .B(n52589), .Z(n52556) );
  NANDN U62181 ( .A(n52590), .B(n52591), .Z(n52589) );
  OR U62182 ( .A(n52592), .B(n52593), .Z(n52591) );
  NANDN U62183 ( .A(n52594), .B(n52592), .Z(n52588) );
  IV U62184 ( .A(n52593), .Z(n52594) );
  XNOR U62185 ( .A(n52564), .B(n52595), .Z(n52559) );
  XNOR U62186 ( .A(n52562), .B(n52565), .Z(n52595) );
  NAND U62187 ( .A(n52596), .B(n52597), .Z(n52565) );
  NAND U62188 ( .A(n52598), .B(n52599), .Z(n52597) );
  OR U62189 ( .A(n52600), .B(n52601), .Z(n52598) );
  NANDN U62190 ( .A(n52602), .B(n52600), .Z(n52596) );
  IV U62191 ( .A(n52601), .Z(n52602) );
  NAND U62192 ( .A(n52603), .B(n52604), .Z(n52562) );
  NAND U62193 ( .A(n52605), .B(n52606), .Z(n52604) );
  NANDN U62194 ( .A(n52607), .B(n52608), .Z(n52605) );
  NANDN U62195 ( .A(n52608), .B(n52607), .Z(n52603) );
  AND U62196 ( .A(n52609), .B(n52610), .Z(n52564) );
  NAND U62197 ( .A(n52611), .B(n52612), .Z(n52610) );
  OR U62198 ( .A(n52613), .B(n52614), .Z(n52611) );
  NANDN U62199 ( .A(n52615), .B(n52613), .Z(n52609) );
  XNOR U62200 ( .A(n52590), .B(n52616), .Z(N60736) );
  XOR U62201 ( .A(n52592), .B(n52593), .Z(n52616) );
  XNOR U62202 ( .A(n52606), .B(n52617), .Z(n52593) );
  XOR U62203 ( .A(n52607), .B(n52608), .Z(n52617) );
  XOR U62204 ( .A(n52613), .B(n52618), .Z(n52608) );
  XOR U62205 ( .A(n52612), .B(n52615), .Z(n52618) );
  IV U62206 ( .A(n52614), .Z(n52615) );
  NAND U62207 ( .A(n52619), .B(n52620), .Z(n52614) );
  OR U62208 ( .A(n52621), .B(n52622), .Z(n52620) );
  OR U62209 ( .A(n52623), .B(n52624), .Z(n52619) );
  NAND U62210 ( .A(n52625), .B(n52626), .Z(n52612) );
  OR U62211 ( .A(n52627), .B(n52628), .Z(n52626) );
  OR U62212 ( .A(n52629), .B(n52630), .Z(n52625) );
  NOR U62213 ( .A(n52631), .B(n52632), .Z(n52613) );
  ANDN U62214 ( .B(n52633), .A(n52634), .Z(n52607) );
  XNOR U62215 ( .A(n52600), .B(n52635), .Z(n52606) );
  XNOR U62216 ( .A(n52599), .B(n52601), .Z(n52635) );
  NAND U62217 ( .A(n52636), .B(n52637), .Z(n52601) );
  OR U62218 ( .A(n52638), .B(n52639), .Z(n52637) );
  OR U62219 ( .A(n52640), .B(n52641), .Z(n52636) );
  NAND U62220 ( .A(n52642), .B(n52643), .Z(n52599) );
  OR U62221 ( .A(n52644), .B(n52645), .Z(n52643) );
  OR U62222 ( .A(n52646), .B(n52647), .Z(n52642) );
  ANDN U62223 ( .B(n52648), .A(n52649), .Z(n52600) );
  IV U62224 ( .A(n52650), .Z(n52648) );
  ANDN U62225 ( .B(n52651), .A(n52652), .Z(n52592) );
  XOR U62226 ( .A(n52578), .B(n52653), .Z(n52590) );
  XOR U62227 ( .A(n52579), .B(n52580), .Z(n52653) );
  XOR U62228 ( .A(n52585), .B(n52654), .Z(n52580) );
  XOR U62229 ( .A(n52584), .B(n52587), .Z(n52654) );
  IV U62230 ( .A(n52586), .Z(n52587) );
  NAND U62231 ( .A(n52655), .B(n52656), .Z(n52586) );
  OR U62232 ( .A(n52657), .B(n52658), .Z(n52656) );
  OR U62233 ( .A(n52659), .B(n52660), .Z(n52655) );
  NAND U62234 ( .A(n52661), .B(n52662), .Z(n52584) );
  OR U62235 ( .A(n52663), .B(n52664), .Z(n52662) );
  OR U62236 ( .A(n52665), .B(n52666), .Z(n52661) );
  NOR U62237 ( .A(n52667), .B(n52668), .Z(n52585) );
  ANDN U62238 ( .B(n52669), .A(n52670), .Z(n52579) );
  IV U62239 ( .A(n52671), .Z(n52669) );
  XNOR U62240 ( .A(n52572), .B(n52672), .Z(n52578) );
  XNOR U62241 ( .A(n52571), .B(n52573), .Z(n52672) );
  NAND U62242 ( .A(n52673), .B(n52674), .Z(n52573) );
  OR U62243 ( .A(n52675), .B(n52676), .Z(n52674) );
  OR U62244 ( .A(n52677), .B(n52678), .Z(n52673) );
  NAND U62245 ( .A(n52679), .B(n52680), .Z(n52571) );
  OR U62246 ( .A(n52681), .B(n52682), .Z(n52680) );
  OR U62247 ( .A(n52683), .B(n52684), .Z(n52679) );
  ANDN U62248 ( .B(n52685), .A(n52686), .Z(n52572) );
  IV U62249 ( .A(n52687), .Z(n52685) );
  XNOR U62250 ( .A(n52652), .B(n52651), .Z(N60735) );
  XOR U62251 ( .A(n52671), .B(n52670), .Z(n52651) );
  XNOR U62252 ( .A(n52686), .B(n52687), .Z(n52670) );
  XNOR U62253 ( .A(n52681), .B(n52682), .Z(n52687) );
  XNOR U62254 ( .A(n52683), .B(n52684), .Z(n52682) );
  XNOR U62255 ( .A(y[277]), .B(x[277]), .Z(n52684) );
  XNOR U62256 ( .A(y[278]), .B(x[278]), .Z(n52683) );
  XNOR U62257 ( .A(y[276]), .B(x[276]), .Z(n52681) );
  XNOR U62258 ( .A(n52675), .B(n52676), .Z(n52686) );
  XNOR U62259 ( .A(y[273]), .B(x[273]), .Z(n52676) );
  XNOR U62260 ( .A(n52677), .B(n52678), .Z(n52675) );
  XNOR U62261 ( .A(y[274]), .B(x[274]), .Z(n52678) );
  XNOR U62262 ( .A(y[275]), .B(x[275]), .Z(n52677) );
  XNOR U62263 ( .A(n52668), .B(n52667), .Z(n52671) );
  XNOR U62264 ( .A(n52663), .B(n52664), .Z(n52667) );
  XNOR U62265 ( .A(y[270]), .B(x[270]), .Z(n52664) );
  XNOR U62266 ( .A(n52665), .B(n52666), .Z(n52663) );
  XNOR U62267 ( .A(y[271]), .B(x[271]), .Z(n52666) );
  XNOR U62268 ( .A(y[272]), .B(x[272]), .Z(n52665) );
  XNOR U62269 ( .A(n52657), .B(n52658), .Z(n52668) );
  XNOR U62270 ( .A(y[267]), .B(x[267]), .Z(n52658) );
  XNOR U62271 ( .A(n52659), .B(n52660), .Z(n52657) );
  XNOR U62272 ( .A(y[268]), .B(x[268]), .Z(n52660) );
  XNOR U62273 ( .A(y[269]), .B(x[269]), .Z(n52659) );
  XOR U62274 ( .A(n52633), .B(n52634), .Z(n52652) );
  XNOR U62275 ( .A(n52649), .B(n52650), .Z(n52634) );
  XNOR U62276 ( .A(n52644), .B(n52645), .Z(n52650) );
  XNOR U62277 ( .A(n52646), .B(n52647), .Z(n52645) );
  XNOR U62278 ( .A(y[265]), .B(x[265]), .Z(n52647) );
  XNOR U62279 ( .A(y[266]), .B(x[266]), .Z(n52646) );
  XNOR U62280 ( .A(y[264]), .B(x[264]), .Z(n52644) );
  XNOR U62281 ( .A(n52638), .B(n52639), .Z(n52649) );
  XNOR U62282 ( .A(y[261]), .B(x[261]), .Z(n52639) );
  XNOR U62283 ( .A(n52640), .B(n52641), .Z(n52638) );
  XNOR U62284 ( .A(y[262]), .B(x[262]), .Z(n52641) );
  XNOR U62285 ( .A(y[263]), .B(x[263]), .Z(n52640) );
  XOR U62286 ( .A(n52632), .B(n52631), .Z(n52633) );
  XNOR U62287 ( .A(n52627), .B(n52628), .Z(n52631) );
  XNOR U62288 ( .A(y[258]), .B(x[258]), .Z(n52628) );
  XNOR U62289 ( .A(n52629), .B(n52630), .Z(n52627) );
  XNOR U62290 ( .A(y[259]), .B(x[259]), .Z(n52630) );
  XNOR U62291 ( .A(y[260]), .B(x[260]), .Z(n52629) );
  XNOR U62292 ( .A(n52621), .B(n52622), .Z(n52632) );
  XNOR U62293 ( .A(y[255]), .B(x[255]), .Z(n52622) );
  XNOR U62294 ( .A(n52623), .B(n52624), .Z(n52621) );
  XNOR U62295 ( .A(y[256]), .B(x[256]), .Z(n52624) );
  XNOR U62296 ( .A(y[257]), .B(x[257]), .Z(n52623) );
  NAND U62297 ( .A(n52688), .B(n52689), .Z(N60726) );
  NANDN U62298 ( .A(n52690), .B(n52691), .Z(n52689) );
  OR U62299 ( .A(n52692), .B(n52693), .Z(n52691) );
  NAND U62300 ( .A(n52692), .B(n52693), .Z(n52688) );
  XOR U62301 ( .A(n52692), .B(n52694), .Z(N60725) );
  XNOR U62302 ( .A(n52690), .B(n52693), .Z(n52694) );
  AND U62303 ( .A(n52695), .B(n52696), .Z(n52693) );
  NANDN U62304 ( .A(n52697), .B(n52698), .Z(n52696) );
  NANDN U62305 ( .A(n52699), .B(n52700), .Z(n52698) );
  NANDN U62306 ( .A(n52700), .B(n52699), .Z(n52695) );
  NAND U62307 ( .A(n52701), .B(n52702), .Z(n52690) );
  NANDN U62308 ( .A(n52703), .B(n52704), .Z(n52702) );
  OR U62309 ( .A(n52705), .B(n52706), .Z(n52704) );
  NAND U62310 ( .A(n52706), .B(n52705), .Z(n52701) );
  AND U62311 ( .A(n52707), .B(n52708), .Z(n52692) );
  NANDN U62312 ( .A(n52709), .B(n52710), .Z(n52708) );
  NANDN U62313 ( .A(n52711), .B(n52712), .Z(n52710) );
  NANDN U62314 ( .A(n52712), .B(n52711), .Z(n52707) );
  XOR U62315 ( .A(n52706), .B(n52713), .Z(N60724) );
  XOR U62316 ( .A(n52703), .B(n52705), .Z(n52713) );
  XNOR U62317 ( .A(n52699), .B(n52714), .Z(n52705) );
  XNOR U62318 ( .A(n52697), .B(n52700), .Z(n52714) );
  NAND U62319 ( .A(n52715), .B(n52716), .Z(n52700) );
  NAND U62320 ( .A(n52717), .B(n52718), .Z(n52716) );
  OR U62321 ( .A(n52719), .B(n52720), .Z(n52717) );
  NANDN U62322 ( .A(n52721), .B(n52719), .Z(n52715) );
  IV U62323 ( .A(n52720), .Z(n52721) );
  NAND U62324 ( .A(n52722), .B(n52723), .Z(n52697) );
  NAND U62325 ( .A(n52724), .B(n52725), .Z(n52723) );
  NANDN U62326 ( .A(n52726), .B(n52727), .Z(n52724) );
  NANDN U62327 ( .A(n52727), .B(n52726), .Z(n52722) );
  AND U62328 ( .A(n52728), .B(n52729), .Z(n52699) );
  NAND U62329 ( .A(n52730), .B(n52731), .Z(n52729) );
  OR U62330 ( .A(n52732), .B(n52733), .Z(n52730) );
  NANDN U62331 ( .A(n52734), .B(n52732), .Z(n52728) );
  NAND U62332 ( .A(n52735), .B(n52736), .Z(n52703) );
  NANDN U62333 ( .A(n52737), .B(n52738), .Z(n52736) );
  OR U62334 ( .A(n52739), .B(n52740), .Z(n52738) );
  NANDN U62335 ( .A(n52741), .B(n52739), .Z(n52735) );
  IV U62336 ( .A(n52740), .Z(n52741) );
  XNOR U62337 ( .A(n52711), .B(n52742), .Z(n52706) );
  XNOR U62338 ( .A(n52709), .B(n52712), .Z(n52742) );
  NAND U62339 ( .A(n52743), .B(n52744), .Z(n52712) );
  NAND U62340 ( .A(n52745), .B(n52746), .Z(n52744) );
  OR U62341 ( .A(n52747), .B(n52748), .Z(n52745) );
  NANDN U62342 ( .A(n52749), .B(n52747), .Z(n52743) );
  IV U62343 ( .A(n52748), .Z(n52749) );
  NAND U62344 ( .A(n52750), .B(n52751), .Z(n52709) );
  NAND U62345 ( .A(n52752), .B(n52753), .Z(n52751) );
  NANDN U62346 ( .A(n52754), .B(n52755), .Z(n52752) );
  NANDN U62347 ( .A(n52755), .B(n52754), .Z(n52750) );
  AND U62348 ( .A(n52756), .B(n52757), .Z(n52711) );
  NAND U62349 ( .A(n52758), .B(n52759), .Z(n52757) );
  OR U62350 ( .A(n52760), .B(n52761), .Z(n52758) );
  NANDN U62351 ( .A(n52762), .B(n52760), .Z(n52756) );
  XNOR U62352 ( .A(n52737), .B(n52763), .Z(N60723) );
  XOR U62353 ( .A(n52739), .B(n52740), .Z(n52763) );
  XNOR U62354 ( .A(n52753), .B(n52764), .Z(n52740) );
  XOR U62355 ( .A(n52754), .B(n52755), .Z(n52764) );
  XOR U62356 ( .A(n52760), .B(n52765), .Z(n52755) );
  XOR U62357 ( .A(n52759), .B(n52762), .Z(n52765) );
  IV U62358 ( .A(n52761), .Z(n52762) );
  NAND U62359 ( .A(n52766), .B(n52767), .Z(n52761) );
  OR U62360 ( .A(n52768), .B(n52769), .Z(n52767) );
  OR U62361 ( .A(n52770), .B(n52771), .Z(n52766) );
  NAND U62362 ( .A(n52772), .B(n52773), .Z(n52759) );
  OR U62363 ( .A(n52774), .B(n52775), .Z(n52773) );
  OR U62364 ( .A(n52776), .B(n52777), .Z(n52772) );
  NOR U62365 ( .A(n52778), .B(n52779), .Z(n52760) );
  ANDN U62366 ( .B(n52780), .A(n52781), .Z(n52754) );
  XNOR U62367 ( .A(n52747), .B(n52782), .Z(n52753) );
  XNOR U62368 ( .A(n52746), .B(n52748), .Z(n52782) );
  NAND U62369 ( .A(n52783), .B(n52784), .Z(n52748) );
  OR U62370 ( .A(n52785), .B(n52786), .Z(n52784) );
  OR U62371 ( .A(n52787), .B(n52788), .Z(n52783) );
  NAND U62372 ( .A(n52789), .B(n52790), .Z(n52746) );
  OR U62373 ( .A(n52791), .B(n52792), .Z(n52790) );
  OR U62374 ( .A(n52793), .B(n52794), .Z(n52789) );
  ANDN U62375 ( .B(n52795), .A(n52796), .Z(n52747) );
  IV U62376 ( .A(n52797), .Z(n52795) );
  ANDN U62377 ( .B(n52798), .A(n52799), .Z(n52739) );
  XOR U62378 ( .A(n52725), .B(n52800), .Z(n52737) );
  XOR U62379 ( .A(n52726), .B(n52727), .Z(n52800) );
  XOR U62380 ( .A(n52732), .B(n52801), .Z(n52727) );
  XOR U62381 ( .A(n52731), .B(n52734), .Z(n52801) );
  IV U62382 ( .A(n52733), .Z(n52734) );
  NAND U62383 ( .A(n52802), .B(n52803), .Z(n52733) );
  OR U62384 ( .A(n52804), .B(n52805), .Z(n52803) );
  OR U62385 ( .A(n52806), .B(n52807), .Z(n52802) );
  NAND U62386 ( .A(n52808), .B(n52809), .Z(n52731) );
  OR U62387 ( .A(n52810), .B(n52811), .Z(n52809) );
  OR U62388 ( .A(n52812), .B(n52813), .Z(n52808) );
  NOR U62389 ( .A(n52814), .B(n52815), .Z(n52732) );
  ANDN U62390 ( .B(n52816), .A(n52817), .Z(n52726) );
  IV U62391 ( .A(n52818), .Z(n52816) );
  XNOR U62392 ( .A(n52719), .B(n52819), .Z(n52725) );
  XNOR U62393 ( .A(n52718), .B(n52720), .Z(n52819) );
  NAND U62394 ( .A(n52820), .B(n52821), .Z(n52720) );
  OR U62395 ( .A(n52822), .B(n52823), .Z(n52821) );
  OR U62396 ( .A(n52824), .B(n52825), .Z(n52820) );
  NAND U62397 ( .A(n52826), .B(n52827), .Z(n52718) );
  OR U62398 ( .A(n52828), .B(n52829), .Z(n52827) );
  OR U62399 ( .A(n52830), .B(n52831), .Z(n52826) );
  ANDN U62400 ( .B(n52832), .A(n52833), .Z(n52719) );
  IV U62401 ( .A(n52834), .Z(n52832) );
  XNOR U62402 ( .A(n52799), .B(n52798), .Z(N60722) );
  XOR U62403 ( .A(n52818), .B(n52817), .Z(n52798) );
  XNOR U62404 ( .A(n52833), .B(n52834), .Z(n52817) );
  XNOR U62405 ( .A(n52828), .B(n52829), .Z(n52834) );
  XNOR U62406 ( .A(n52830), .B(n52831), .Z(n52829) );
  XNOR U62407 ( .A(y[253]), .B(x[253]), .Z(n52831) );
  XNOR U62408 ( .A(y[254]), .B(x[254]), .Z(n52830) );
  XNOR U62409 ( .A(y[252]), .B(x[252]), .Z(n52828) );
  XNOR U62410 ( .A(n52822), .B(n52823), .Z(n52833) );
  XNOR U62411 ( .A(y[249]), .B(x[249]), .Z(n52823) );
  XNOR U62412 ( .A(n52824), .B(n52825), .Z(n52822) );
  XNOR U62413 ( .A(y[250]), .B(x[250]), .Z(n52825) );
  XNOR U62414 ( .A(y[251]), .B(x[251]), .Z(n52824) );
  XNOR U62415 ( .A(n52815), .B(n52814), .Z(n52818) );
  XNOR U62416 ( .A(n52810), .B(n52811), .Z(n52814) );
  XNOR U62417 ( .A(y[246]), .B(x[246]), .Z(n52811) );
  XNOR U62418 ( .A(n52812), .B(n52813), .Z(n52810) );
  XNOR U62419 ( .A(y[247]), .B(x[247]), .Z(n52813) );
  XNOR U62420 ( .A(y[248]), .B(x[248]), .Z(n52812) );
  XNOR U62421 ( .A(n52804), .B(n52805), .Z(n52815) );
  XNOR U62422 ( .A(y[243]), .B(x[243]), .Z(n52805) );
  XNOR U62423 ( .A(n52806), .B(n52807), .Z(n52804) );
  XNOR U62424 ( .A(y[244]), .B(x[244]), .Z(n52807) );
  XNOR U62425 ( .A(y[245]), .B(x[245]), .Z(n52806) );
  XOR U62426 ( .A(n52780), .B(n52781), .Z(n52799) );
  XNOR U62427 ( .A(n52796), .B(n52797), .Z(n52781) );
  XNOR U62428 ( .A(n52791), .B(n52792), .Z(n52797) );
  XNOR U62429 ( .A(n52793), .B(n52794), .Z(n52792) );
  XNOR U62430 ( .A(y[241]), .B(x[241]), .Z(n52794) );
  XNOR U62431 ( .A(y[242]), .B(x[242]), .Z(n52793) );
  XNOR U62432 ( .A(y[240]), .B(x[240]), .Z(n52791) );
  XNOR U62433 ( .A(n52785), .B(n52786), .Z(n52796) );
  XNOR U62434 ( .A(y[237]), .B(x[237]), .Z(n52786) );
  XNOR U62435 ( .A(n52787), .B(n52788), .Z(n52785) );
  XNOR U62436 ( .A(y[238]), .B(x[238]), .Z(n52788) );
  XNOR U62437 ( .A(y[239]), .B(x[239]), .Z(n52787) );
  XOR U62438 ( .A(n52779), .B(n52778), .Z(n52780) );
  XNOR U62439 ( .A(n52774), .B(n52775), .Z(n52778) );
  XNOR U62440 ( .A(y[234]), .B(x[234]), .Z(n52775) );
  XNOR U62441 ( .A(n52776), .B(n52777), .Z(n52774) );
  XNOR U62442 ( .A(y[235]), .B(x[235]), .Z(n52777) );
  XNOR U62443 ( .A(y[236]), .B(x[236]), .Z(n52776) );
  XNOR U62444 ( .A(n52768), .B(n52769), .Z(n52779) );
  XNOR U62445 ( .A(y[231]), .B(x[231]), .Z(n52769) );
  XNOR U62446 ( .A(n52770), .B(n52771), .Z(n52768) );
  XNOR U62447 ( .A(y[232]), .B(x[232]), .Z(n52771) );
  XNOR U62448 ( .A(y[233]), .B(x[233]), .Z(n52770) );
  NAND U62449 ( .A(n52835), .B(n52836), .Z(N60713) );
  NANDN U62450 ( .A(n52837), .B(n52838), .Z(n52836) );
  OR U62451 ( .A(n52839), .B(n52840), .Z(n52838) );
  NAND U62452 ( .A(n52839), .B(n52840), .Z(n52835) );
  XOR U62453 ( .A(n52839), .B(n52841), .Z(N60712) );
  XNOR U62454 ( .A(n52837), .B(n52840), .Z(n52841) );
  AND U62455 ( .A(n52842), .B(n52843), .Z(n52840) );
  NANDN U62456 ( .A(n52844), .B(n52845), .Z(n52843) );
  NANDN U62457 ( .A(n52846), .B(n52847), .Z(n52845) );
  NANDN U62458 ( .A(n52847), .B(n52846), .Z(n52842) );
  NAND U62459 ( .A(n52848), .B(n52849), .Z(n52837) );
  NANDN U62460 ( .A(n52850), .B(n52851), .Z(n52849) );
  OR U62461 ( .A(n52852), .B(n52853), .Z(n52851) );
  NAND U62462 ( .A(n52853), .B(n52852), .Z(n52848) );
  AND U62463 ( .A(n52854), .B(n52855), .Z(n52839) );
  NANDN U62464 ( .A(n52856), .B(n52857), .Z(n52855) );
  NANDN U62465 ( .A(n52858), .B(n52859), .Z(n52857) );
  NANDN U62466 ( .A(n52859), .B(n52858), .Z(n52854) );
  XOR U62467 ( .A(n52853), .B(n52860), .Z(N60711) );
  XOR U62468 ( .A(n52850), .B(n52852), .Z(n52860) );
  XNOR U62469 ( .A(n52846), .B(n52861), .Z(n52852) );
  XNOR U62470 ( .A(n52844), .B(n52847), .Z(n52861) );
  NAND U62471 ( .A(n52862), .B(n52863), .Z(n52847) );
  NAND U62472 ( .A(n52864), .B(n52865), .Z(n52863) );
  OR U62473 ( .A(n52866), .B(n52867), .Z(n52864) );
  NANDN U62474 ( .A(n52868), .B(n52866), .Z(n52862) );
  IV U62475 ( .A(n52867), .Z(n52868) );
  NAND U62476 ( .A(n52869), .B(n52870), .Z(n52844) );
  NAND U62477 ( .A(n52871), .B(n52872), .Z(n52870) );
  NANDN U62478 ( .A(n52873), .B(n52874), .Z(n52871) );
  NANDN U62479 ( .A(n52874), .B(n52873), .Z(n52869) );
  AND U62480 ( .A(n52875), .B(n52876), .Z(n52846) );
  NAND U62481 ( .A(n52877), .B(n52878), .Z(n52876) );
  OR U62482 ( .A(n52879), .B(n52880), .Z(n52877) );
  NANDN U62483 ( .A(n52881), .B(n52879), .Z(n52875) );
  NAND U62484 ( .A(n52882), .B(n52883), .Z(n52850) );
  NANDN U62485 ( .A(n52884), .B(n52885), .Z(n52883) );
  OR U62486 ( .A(n52886), .B(n52887), .Z(n52885) );
  NANDN U62487 ( .A(n52888), .B(n52886), .Z(n52882) );
  IV U62488 ( .A(n52887), .Z(n52888) );
  XNOR U62489 ( .A(n52858), .B(n52889), .Z(n52853) );
  XNOR U62490 ( .A(n52856), .B(n52859), .Z(n52889) );
  NAND U62491 ( .A(n52890), .B(n52891), .Z(n52859) );
  NAND U62492 ( .A(n52892), .B(n52893), .Z(n52891) );
  OR U62493 ( .A(n52894), .B(n52895), .Z(n52892) );
  NANDN U62494 ( .A(n52896), .B(n52894), .Z(n52890) );
  IV U62495 ( .A(n52895), .Z(n52896) );
  NAND U62496 ( .A(n52897), .B(n52898), .Z(n52856) );
  NAND U62497 ( .A(n52899), .B(n52900), .Z(n52898) );
  NANDN U62498 ( .A(n52901), .B(n52902), .Z(n52899) );
  NANDN U62499 ( .A(n52902), .B(n52901), .Z(n52897) );
  AND U62500 ( .A(n52903), .B(n52904), .Z(n52858) );
  NAND U62501 ( .A(n52905), .B(n52906), .Z(n52904) );
  OR U62502 ( .A(n52907), .B(n52908), .Z(n52905) );
  NANDN U62503 ( .A(n52909), .B(n52907), .Z(n52903) );
  XNOR U62504 ( .A(n52884), .B(n52910), .Z(N60710) );
  XOR U62505 ( .A(n52886), .B(n52887), .Z(n52910) );
  XNOR U62506 ( .A(n52900), .B(n52911), .Z(n52887) );
  XOR U62507 ( .A(n52901), .B(n52902), .Z(n52911) );
  XOR U62508 ( .A(n52907), .B(n52912), .Z(n52902) );
  XOR U62509 ( .A(n52906), .B(n52909), .Z(n52912) );
  IV U62510 ( .A(n52908), .Z(n52909) );
  NAND U62511 ( .A(n52913), .B(n52914), .Z(n52908) );
  OR U62512 ( .A(n52915), .B(n52916), .Z(n52914) );
  OR U62513 ( .A(n52917), .B(n52918), .Z(n52913) );
  NAND U62514 ( .A(n52919), .B(n52920), .Z(n52906) );
  OR U62515 ( .A(n52921), .B(n52922), .Z(n52920) );
  OR U62516 ( .A(n52923), .B(n52924), .Z(n52919) );
  NOR U62517 ( .A(n52925), .B(n52926), .Z(n52907) );
  ANDN U62518 ( .B(n52927), .A(n52928), .Z(n52901) );
  XNOR U62519 ( .A(n52894), .B(n52929), .Z(n52900) );
  XNOR U62520 ( .A(n52893), .B(n52895), .Z(n52929) );
  NAND U62521 ( .A(n52930), .B(n52931), .Z(n52895) );
  OR U62522 ( .A(n52932), .B(n52933), .Z(n52931) );
  OR U62523 ( .A(n52934), .B(n52935), .Z(n52930) );
  NAND U62524 ( .A(n52936), .B(n52937), .Z(n52893) );
  OR U62525 ( .A(n52938), .B(n52939), .Z(n52937) );
  OR U62526 ( .A(n52940), .B(n52941), .Z(n52936) );
  ANDN U62527 ( .B(n52942), .A(n52943), .Z(n52894) );
  IV U62528 ( .A(n52944), .Z(n52942) );
  ANDN U62529 ( .B(n52945), .A(n52946), .Z(n52886) );
  XOR U62530 ( .A(n52872), .B(n52947), .Z(n52884) );
  XOR U62531 ( .A(n52873), .B(n52874), .Z(n52947) );
  XOR U62532 ( .A(n52879), .B(n52948), .Z(n52874) );
  XOR U62533 ( .A(n52878), .B(n52881), .Z(n52948) );
  IV U62534 ( .A(n52880), .Z(n52881) );
  NAND U62535 ( .A(n52949), .B(n52950), .Z(n52880) );
  OR U62536 ( .A(n52951), .B(n52952), .Z(n52950) );
  OR U62537 ( .A(n52953), .B(n52954), .Z(n52949) );
  NAND U62538 ( .A(n52955), .B(n52956), .Z(n52878) );
  OR U62539 ( .A(n52957), .B(n52958), .Z(n52956) );
  OR U62540 ( .A(n52959), .B(n52960), .Z(n52955) );
  NOR U62541 ( .A(n52961), .B(n52962), .Z(n52879) );
  ANDN U62542 ( .B(n52963), .A(n52964), .Z(n52873) );
  IV U62543 ( .A(n52965), .Z(n52963) );
  XNOR U62544 ( .A(n52866), .B(n52966), .Z(n52872) );
  XNOR U62545 ( .A(n52865), .B(n52867), .Z(n52966) );
  NAND U62546 ( .A(n52967), .B(n52968), .Z(n52867) );
  OR U62547 ( .A(n52969), .B(n52970), .Z(n52968) );
  OR U62548 ( .A(n52971), .B(n52972), .Z(n52967) );
  NAND U62549 ( .A(n52973), .B(n52974), .Z(n52865) );
  OR U62550 ( .A(n52975), .B(n52976), .Z(n52974) );
  OR U62551 ( .A(n52977), .B(n52978), .Z(n52973) );
  ANDN U62552 ( .B(n52979), .A(n52980), .Z(n52866) );
  IV U62553 ( .A(n52981), .Z(n52979) );
  XNOR U62554 ( .A(n52946), .B(n52945), .Z(N60709) );
  XOR U62555 ( .A(n52965), .B(n52964), .Z(n52945) );
  XNOR U62556 ( .A(n52980), .B(n52981), .Z(n52964) );
  XNOR U62557 ( .A(n52975), .B(n52976), .Z(n52981) );
  XNOR U62558 ( .A(n52977), .B(n52978), .Z(n52976) );
  XNOR U62559 ( .A(y[229]), .B(x[229]), .Z(n52978) );
  XNOR U62560 ( .A(y[230]), .B(x[230]), .Z(n52977) );
  XNOR U62561 ( .A(y[228]), .B(x[228]), .Z(n52975) );
  XNOR U62562 ( .A(n52969), .B(n52970), .Z(n52980) );
  XNOR U62563 ( .A(y[225]), .B(x[225]), .Z(n52970) );
  XNOR U62564 ( .A(n52971), .B(n52972), .Z(n52969) );
  XNOR U62565 ( .A(y[226]), .B(x[226]), .Z(n52972) );
  XNOR U62566 ( .A(y[227]), .B(x[227]), .Z(n52971) );
  XNOR U62567 ( .A(n52962), .B(n52961), .Z(n52965) );
  XNOR U62568 ( .A(n52957), .B(n52958), .Z(n52961) );
  XNOR U62569 ( .A(y[222]), .B(x[222]), .Z(n52958) );
  XNOR U62570 ( .A(n52959), .B(n52960), .Z(n52957) );
  XNOR U62571 ( .A(y[223]), .B(x[223]), .Z(n52960) );
  XNOR U62572 ( .A(y[224]), .B(x[224]), .Z(n52959) );
  XNOR U62573 ( .A(n52951), .B(n52952), .Z(n52962) );
  XNOR U62574 ( .A(y[219]), .B(x[219]), .Z(n52952) );
  XNOR U62575 ( .A(n52953), .B(n52954), .Z(n52951) );
  XNOR U62576 ( .A(y[220]), .B(x[220]), .Z(n52954) );
  XNOR U62577 ( .A(y[221]), .B(x[221]), .Z(n52953) );
  XOR U62578 ( .A(n52927), .B(n52928), .Z(n52946) );
  XNOR U62579 ( .A(n52943), .B(n52944), .Z(n52928) );
  XNOR U62580 ( .A(n52938), .B(n52939), .Z(n52944) );
  XNOR U62581 ( .A(n52940), .B(n52941), .Z(n52939) );
  XNOR U62582 ( .A(y[217]), .B(x[217]), .Z(n52941) );
  XNOR U62583 ( .A(y[218]), .B(x[218]), .Z(n52940) );
  XNOR U62584 ( .A(y[216]), .B(x[216]), .Z(n52938) );
  XNOR U62585 ( .A(n52932), .B(n52933), .Z(n52943) );
  XNOR U62586 ( .A(y[213]), .B(x[213]), .Z(n52933) );
  XNOR U62587 ( .A(n52934), .B(n52935), .Z(n52932) );
  XNOR U62588 ( .A(y[214]), .B(x[214]), .Z(n52935) );
  XNOR U62589 ( .A(y[215]), .B(x[215]), .Z(n52934) );
  XOR U62590 ( .A(n52926), .B(n52925), .Z(n52927) );
  XNOR U62591 ( .A(n52921), .B(n52922), .Z(n52925) );
  XNOR U62592 ( .A(y[210]), .B(x[210]), .Z(n52922) );
  XNOR U62593 ( .A(n52923), .B(n52924), .Z(n52921) );
  XNOR U62594 ( .A(y[211]), .B(x[211]), .Z(n52924) );
  XNOR U62595 ( .A(y[212]), .B(x[212]), .Z(n52923) );
  XNOR U62596 ( .A(n52915), .B(n52916), .Z(n52926) );
  XNOR U62597 ( .A(y[207]), .B(x[207]), .Z(n52916) );
  XNOR U62598 ( .A(n52917), .B(n52918), .Z(n52915) );
  XNOR U62599 ( .A(y[208]), .B(x[208]), .Z(n52918) );
  XNOR U62600 ( .A(y[209]), .B(x[209]), .Z(n52917) );
  NAND U62601 ( .A(n52982), .B(n52983), .Z(N60700) );
  NANDN U62602 ( .A(n52984), .B(n52985), .Z(n52983) );
  OR U62603 ( .A(n52986), .B(n52987), .Z(n52985) );
  NAND U62604 ( .A(n52986), .B(n52987), .Z(n52982) );
  XOR U62605 ( .A(n52986), .B(n52988), .Z(N60699) );
  XNOR U62606 ( .A(n52984), .B(n52987), .Z(n52988) );
  AND U62607 ( .A(n52989), .B(n52990), .Z(n52987) );
  NANDN U62608 ( .A(n52991), .B(n52992), .Z(n52990) );
  NANDN U62609 ( .A(n52993), .B(n52994), .Z(n52992) );
  NANDN U62610 ( .A(n52994), .B(n52993), .Z(n52989) );
  NAND U62611 ( .A(n52995), .B(n52996), .Z(n52984) );
  NANDN U62612 ( .A(n52997), .B(n52998), .Z(n52996) );
  OR U62613 ( .A(n52999), .B(n53000), .Z(n52998) );
  NAND U62614 ( .A(n53000), .B(n52999), .Z(n52995) );
  AND U62615 ( .A(n53001), .B(n53002), .Z(n52986) );
  NANDN U62616 ( .A(n53003), .B(n53004), .Z(n53002) );
  NANDN U62617 ( .A(n53005), .B(n53006), .Z(n53004) );
  NANDN U62618 ( .A(n53006), .B(n53005), .Z(n53001) );
  XOR U62619 ( .A(n53000), .B(n53007), .Z(N60698) );
  XOR U62620 ( .A(n52997), .B(n52999), .Z(n53007) );
  XNOR U62621 ( .A(n52993), .B(n53008), .Z(n52999) );
  XNOR U62622 ( .A(n52991), .B(n52994), .Z(n53008) );
  NAND U62623 ( .A(n53009), .B(n53010), .Z(n52994) );
  NAND U62624 ( .A(n53011), .B(n53012), .Z(n53010) );
  OR U62625 ( .A(n53013), .B(n53014), .Z(n53011) );
  NANDN U62626 ( .A(n53015), .B(n53013), .Z(n53009) );
  IV U62627 ( .A(n53014), .Z(n53015) );
  NAND U62628 ( .A(n53016), .B(n53017), .Z(n52991) );
  NAND U62629 ( .A(n53018), .B(n53019), .Z(n53017) );
  NANDN U62630 ( .A(n53020), .B(n53021), .Z(n53018) );
  NANDN U62631 ( .A(n53021), .B(n53020), .Z(n53016) );
  AND U62632 ( .A(n53022), .B(n53023), .Z(n52993) );
  NAND U62633 ( .A(n53024), .B(n53025), .Z(n53023) );
  OR U62634 ( .A(n53026), .B(n53027), .Z(n53024) );
  NANDN U62635 ( .A(n53028), .B(n53026), .Z(n53022) );
  NAND U62636 ( .A(n53029), .B(n53030), .Z(n52997) );
  NANDN U62637 ( .A(n53031), .B(n53032), .Z(n53030) );
  OR U62638 ( .A(n53033), .B(n53034), .Z(n53032) );
  NANDN U62639 ( .A(n53035), .B(n53033), .Z(n53029) );
  IV U62640 ( .A(n53034), .Z(n53035) );
  XNOR U62641 ( .A(n53005), .B(n53036), .Z(n53000) );
  XNOR U62642 ( .A(n53003), .B(n53006), .Z(n53036) );
  NAND U62643 ( .A(n53037), .B(n53038), .Z(n53006) );
  NAND U62644 ( .A(n53039), .B(n53040), .Z(n53038) );
  OR U62645 ( .A(n53041), .B(n53042), .Z(n53039) );
  NANDN U62646 ( .A(n53043), .B(n53041), .Z(n53037) );
  IV U62647 ( .A(n53042), .Z(n53043) );
  NAND U62648 ( .A(n53044), .B(n53045), .Z(n53003) );
  NAND U62649 ( .A(n53046), .B(n53047), .Z(n53045) );
  NANDN U62650 ( .A(n53048), .B(n53049), .Z(n53046) );
  NANDN U62651 ( .A(n53049), .B(n53048), .Z(n53044) );
  AND U62652 ( .A(n53050), .B(n53051), .Z(n53005) );
  NAND U62653 ( .A(n53052), .B(n53053), .Z(n53051) );
  OR U62654 ( .A(n53054), .B(n53055), .Z(n53052) );
  NANDN U62655 ( .A(n53056), .B(n53054), .Z(n53050) );
  XNOR U62656 ( .A(n53031), .B(n53057), .Z(N60697) );
  XOR U62657 ( .A(n53033), .B(n53034), .Z(n53057) );
  XNOR U62658 ( .A(n53047), .B(n53058), .Z(n53034) );
  XOR U62659 ( .A(n53048), .B(n53049), .Z(n53058) );
  XOR U62660 ( .A(n53054), .B(n53059), .Z(n53049) );
  XOR U62661 ( .A(n53053), .B(n53056), .Z(n53059) );
  IV U62662 ( .A(n53055), .Z(n53056) );
  NAND U62663 ( .A(n53060), .B(n53061), .Z(n53055) );
  OR U62664 ( .A(n53062), .B(n53063), .Z(n53061) );
  OR U62665 ( .A(n53064), .B(n53065), .Z(n53060) );
  NAND U62666 ( .A(n53066), .B(n53067), .Z(n53053) );
  OR U62667 ( .A(n53068), .B(n53069), .Z(n53067) );
  OR U62668 ( .A(n53070), .B(n53071), .Z(n53066) );
  NOR U62669 ( .A(n53072), .B(n53073), .Z(n53054) );
  ANDN U62670 ( .B(n53074), .A(n53075), .Z(n53048) );
  XNOR U62671 ( .A(n53041), .B(n53076), .Z(n53047) );
  XNOR U62672 ( .A(n53040), .B(n53042), .Z(n53076) );
  NAND U62673 ( .A(n53077), .B(n53078), .Z(n53042) );
  OR U62674 ( .A(n53079), .B(n53080), .Z(n53078) );
  OR U62675 ( .A(n53081), .B(n53082), .Z(n53077) );
  NAND U62676 ( .A(n53083), .B(n53084), .Z(n53040) );
  OR U62677 ( .A(n53085), .B(n53086), .Z(n53084) );
  OR U62678 ( .A(n53087), .B(n53088), .Z(n53083) );
  ANDN U62679 ( .B(n53089), .A(n53090), .Z(n53041) );
  IV U62680 ( .A(n53091), .Z(n53089) );
  ANDN U62681 ( .B(n53092), .A(n53093), .Z(n53033) );
  XOR U62682 ( .A(n53019), .B(n53094), .Z(n53031) );
  XOR U62683 ( .A(n53020), .B(n53021), .Z(n53094) );
  XOR U62684 ( .A(n53026), .B(n53095), .Z(n53021) );
  XOR U62685 ( .A(n53025), .B(n53028), .Z(n53095) );
  IV U62686 ( .A(n53027), .Z(n53028) );
  NAND U62687 ( .A(n53096), .B(n53097), .Z(n53027) );
  OR U62688 ( .A(n53098), .B(n53099), .Z(n53097) );
  OR U62689 ( .A(n53100), .B(n53101), .Z(n53096) );
  NAND U62690 ( .A(n53102), .B(n53103), .Z(n53025) );
  OR U62691 ( .A(n53104), .B(n53105), .Z(n53103) );
  OR U62692 ( .A(n53106), .B(n53107), .Z(n53102) );
  NOR U62693 ( .A(n53108), .B(n53109), .Z(n53026) );
  ANDN U62694 ( .B(n53110), .A(n53111), .Z(n53020) );
  IV U62695 ( .A(n53112), .Z(n53110) );
  XNOR U62696 ( .A(n53013), .B(n53113), .Z(n53019) );
  XNOR U62697 ( .A(n53012), .B(n53014), .Z(n53113) );
  NAND U62698 ( .A(n53114), .B(n53115), .Z(n53014) );
  OR U62699 ( .A(n53116), .B(n53117), .Z(n53115) );
  OR U62700 ( .A(n53118), .B(n53119), .Z(n53114) );
  NAND U62701 ( .A(n53120), .B(n53121), .Z(n53012) );
  OR U62702 ( .A(n53122), .B(n53123), .Z(n53121) );
  OR U62703 ( .A(n53124), .B(n53125), .Z(n53120) );
  ANDN U62704 ( .B(n53126), .A(n53127), .Z(n53013) );
  IV U62705 ( .A(n53128), .Z(n53126) );
  XNOR U62706 ( .A(n53093), .B(n53092), .Z(N60696) );
  XOR U62707 ( .A(n53112), .B(n53111), .Z(n53092) );
  XNOR U62708 ( .A(n53127), .B(n53128), .Z(n53111) );
  XNOR U62709 ( .A(n53122), .B(n53123), .Z(n53128) );
  XNOR U62710 ( .A(n53124), .B(n53125), .Z(n53123) );
  XNOR U62711 ( .A(y[205]), .B(x[205]), .Z(n53125) );
  XNOR U62712 ( .A(y[206]), .B(x[206]), .Z(n53124) );
  XNOR U62713 ( .A(y[204]), .B(x[204]), .Z(n53122) );
  XNOR U62714 ( .A(n53116), .B(n53117), .Z(n53127) );
  XNOR U62715 ( .A(y[201]), .B(x[201]), .Z(n53117) );
  XNOR U62716 ( .A(n53118), .B(n53119), .Z(n53116) );
  XNOR U62717 ( .A(y[202]), .B(x[202]), .Z(n53119) );
  XNOR U62718 ( .A(y[203]), .B(x[203]), .Z(n53118) );
  XNOR U62719 ( .A(n53109), .B(n53108), .Z(n53112) );
  XNOR U62720 ( .A(n53104), .B(n53105), .Z(n53108) );
  XNOR U62721 ( .A(y[198]), .B(x[198]), .Z(n53105) );
  XNOR U62722 ( .A(n53106), .B(n53107), .Z(n53104) );
  XNOR U62723 ( .A(y[199]), .B(x[199]), .Z(n53107) );
  XNOR U62724 ( .A(y[200]), .B(x[200]), .Z(n53106) );
  XNOR U62725 ( .A(n53098), .B(n53099), .Z(n53109) );
  XNOR U62726 ( .A(y[195]), .B(x[195]), .Z(n53099) );
  XNOR U62727 ( .A(n53100), .B(n53101), .Z(n53098) );
  XNOR U62728 ( .A(y[196]), .B(x[196]), .Z(n53101) );
  XNOR U62729 ( .A(y[197]), .B(x[197]), .Z(n53100) );
  XOR U62730 ( .A(n53074), .B(n53075), .Z(n53093) );
  XNOR U62731 ( .A(n53090), .B(n53091), .Z(n53075) );
  XNOR U62732 ( .A(n53085), .B(n53086), .Z(n53091) );
  XNOR U62733 ( .A(n53087), .B(n53088), .Z(n53086) );
  XNOR U62734 ( .A(y[193]), .B(x[193]), .Z(n53088) );
  XNOR U62735 ( .A(y[194]), .B(x[194]), .Z(n53087) );
  XNOR U62736 ( .A(y[192]), .B(x[192]), .Z(n53085) );
  XNOR U62737 ( .A(n53079), .B(n53080), .Z(n53090) );
  XNOR U62738 ( .A(y[189]), .B(x[189]), .Z(n53080) );
  XNOR U62739 ( .A(n53081), .B(n53082), .Z(n53079) );
  XNOR U62740 ( .A(y[190]), .B(x[190]), .Z(n53082) );
  XNOR U62741 ( .A(y[191]), .B(x[191]), .Z(n53081) );
  XOR U62742 ( .A(n53073), .B(n53072), .Z(n53074) );
  XNOR U62743 ( .A(n53068), .B(n53069), .Z(n53072) );
  XNOR U62744 ( .A(y[186]), .B(x[186]), .Z(n53069) );
  XNOR U62745 ( .A(n53070), .B(n53071), .Z(n53068) );
  XNOR U62746 ( .A(y[187]), .B(x[187]), .Z(n53071) );
  XNOR U62747 ( .A(y[188]), .B(x[188]), .Z(n53070) );
  XNOR U62748 ( .A(n53062), .B(n53063), .Z(n53073) );
  XNOR U62749 ( .A(y[183]), .B(x[183]), .Z(n53063) );
  XNOR U62750 ( .A(n53064), .B(n53065), .Z(n53062) );
  XNOR U62751 ( .A(y[184]), .B(x[184]), .Z(n53065) );
  XNOR U62752 ( .A(y[185]), .B(x[185]), .Z(n53064) );
  NAND U62753 ( .A(n53129), .B(n53130), .Z(N60687) );
  NANDN U62754 ( .A(n53131), .B(n53132), .Z(n53130) );
  OR U62755 ( .A(n53133), .B(n53134), .Z(n53132) );
  NAND U62756 ( .A(n53133), .B(n53134), .Z(n53129) );
  XOR U62757 ( .A(n53133), .B(n53135), .Z(N60686) );
  XNOR U62758 ( .A(n53131), .B(n53134), .Z(n53135) );
  AND U62759 ( .A(n53136), .B(n53137), .Z(n53134) );
  NANDN U62760 ( .A(n53138), .B(n53139), .Z(n53137) );
  NANDN U62761 ( .A(n53140), .B(n53141), .Z(n53139) );
  NANDN U62762 ( .A(n53141), .B(n53140), .Z(n53136) );
  NAND U62763 ( .A(n53142), .B(n53143), .Z(n53131) );
  NANDN U62764 ( .A(n53144), .B(n53145), .Z(n53143) );
  OR U62765 ( .A(n53146), .B(n53147), .Z(n53145) );
  NAND U62766 ( .A(n53147), .B(n53146), .Z(n53142) );
  AND U62767 ( .A(n53148), .B(n53149), .Z(n53133) );
  NANDN U62768 ( .A(n53150), .B(n53151), .Z(n53149) );
  NANDN U62769 ( .A(n53152), .B(n53153), .Z(n53151) );
  NANDN U62770 ( .A(n53153), .B(n53152), .Z(n53148) );
  XOR U62771 ( .A(n53147), .B(n53154), .Z(N60685) );
  XOR U62772 ( .A(n53144), .B(n53146), .Z(n53154) );
  XNOR U62773 ( .A(n53140), .B(n53155), .Z(n53146) );
  XNOR U62774 ( .A(n53138), .B(n53141), .Z(n53155) );
  NAND U62775 ( .A(n53156), .B(n53157), .Z(n53141) );
  NAND U62776 ( .A(n53158), .B(n53159), .Z(n53157) );
  OR U62777 ( .A(n53160), .B(n53161), .Z(n53158) );
  NANDN U62778 ( .A(n53162), .B(n53160), .Z(n53156) );
  IV U62779 ( .A(n53161), .Z(n53162) );
  NAND U62780 ( .A(n53163), .B(n53164), .Z(n53138) );
  NAND U62781 ( .A(n53165), .B(n53166), .Z(n53164) );
  NANDN U62782 ( .A(n53167), .B(n53168), .Z(n53165) );
  NANDN U62783 ( .A(n53168), .B(n53167), .Z(n53163) );
  AND U62784 ( .A(n53169), .B(n53170), .Z(n53140) );
  NAND U62785 ( .A(n53171), .B(n53172), .Z(n53170) );
  OR U62786 ( .A(n53173), .B(n53174), .Z(n53171) );
  NANDN U62787 ( .A(n53175), .B(n53173), .Z(n53169) );
  NAND U62788 ( .A(n53176), .B(n53177), .Z(n53144) );
  NANDN U62789 ( .A(n53178), .B(n53179), .Z(n53177) );
  OR U62790 ( .A(n53180), .B(n53181), .Z(n53179) );
  NANDN U62791 ( .A(n53182), .B(n53180), .Z(n53176) );
  IV U62792 ( .A(n53181), .Z(n53182) );
  XNOR U62793 ( .A(n53152), .B(n53183), .Z(n53147) );
  XNOR U62794 ( .A(n53150), .B(n53153), .Z(n53183) );
  NAND U62795 ( .A(n53184), .B(n53185), .Z(n53153) );
  NAND U62796 ( .A(n53186), .B(n53187), .Z(n53185) );
  OR U62797 ( .A(n53188), .B(n53189), .Z(n53186) );
  NANDN U62798 ( .A(n53190), .B(n53188), .Z(n53184) );
  IV U62799 ( .A(n53189), .Z(n53190) );
  NAND U62800 ( .A(n53191), .B(n53192), .Z(n53150) );
  NAND U62801 ( .A(n53193), .B(n53194), .Z(n53192) );
  NANDN U62802 ( .A(n53195), .B(n53196), .Z(n53193) );
  NANDN U62803 ( .A(n53196), .B(n53195), .Z(n53191) );
  AND U62804 ( .A(n53197), .B(n53198), .Z(n53152) );
  NAND U62805 ( .A(n53199), .B(n53200), .Z(n53198) );
  OR U62806 ( .A(n53201), .B(n53202), .Z(n53199) );
  NANDN U62807 ( .A(n53203), .B(n53201), .Z(n53197) );
  XNOR U62808 ( .A(n53178), .B(n53204), .Z(N60684) );
  XOR U62809 ( .A(n53180), .B(n53181), .Z(n53204) );
  XNOR U62810 ( .A(n53194), .B(n53205), .Z(n53181) );
  XOR U62811 ( .A(n53195), .B(n53196), .Z(n53205) );
  XOR U62812 ( .A(n53201), .B(n53206), .Z(n53196) );
  XOR U62813 ( .A(n53200), .B(n53203), .Z(n53206) );
  IV U62814 ( .A(n53202), .Z(n53203) );
  NAND U62815 ( .A(n53207), .B(n53208), .Z(n53202) );
  OR U62816 ( .A(n53209), .B(n53210), .Z(n53208) );
  OR U62817 ( .A(n53211), .B(n53212), .Z(n53207) );
  NAND U62818 ( .A(n53213), .B(n53214), .Z(n53200) );
  OR U62819 ( .A(n53215), .B(n53216), .Z(n53214) );
  OR U62820 ( .A(n53217), .B(n53218), .Z(n53213) );
  NOR U62821 ( .A(n53219), .B(n53220), .Z(n53201) );
  ANDN U62822 ( .B(n53221), .A(n53222), .Z(n53195) );
  XNOR U62823 ( .A(n53188), .B(n53223), .Z(n53194) );
  XNOR U62824 ( .A(n53187), .B(n53189), .Z(n53223) );
  NAND U62825 ( .A(n53224), .B(n53225), .Z(n53189) );
  OR U62826 ( .A(n53226), .B(n53227), .Z(n53225) );
  OR U62827 ( .A(n53228), .B(n53229), .Z(n53224) );
  NAND U62828 ( .A(n53230), .B(n53231), .Z(n53187) );
  OR U62829 ( .A(n53232), .B(n53233), .Z(n53231) );
  OR U62830 ( .A(n53234), .B(n53235), .Z(n53230) );
  ANDN U62831 ( .B(n53236), .A(n53237), .Z(n53188) );
  IV U62832 ( .A(n53238), .Z(n53236) );
  ANDN U62833 ( .B(n53239), .A(n53240), .Z(n53180) );
  XOR U62834 ( .A(n53166), .B(n53241), .Z(n53178) );
  XOR U62835 ( .A(n53167), .B(n53168), .Z(n53241) );
  XOR U62836 ( .A(n53173), .B(n53242), .Z(n53168) );
  XOR U62837 ( .A(n53172), .B(n53175), .Z(n53242) );
  IV U62838 ( .A(n53174), .Z(n53175) );
  NAND U62839 ( .A(n53243), .B(n53244), .Z(n53174) );
  OR U62840 ( .A(n53245), .B(n53246), .Z(n53244) );
  OR U62841 ( .A(n53247), .B(n53248), .Z(n53243) );
  NAND U62842 ( .A(n53249), .B(n53250), .Z(n53172) );
  OR U62843 ( .A(n53251), .B(n53252), .Z(n53250) );
  OR U62844 ( .A(n53253), .B(n53254), .Z(n53249) );
  NOR U62845 ( .A(n53255), .B(n53256), .Z(n53173) );
  ANDN U62846 ( .B(n53257), .A(n53258), .Z(n53167) );
  IV U62847 ( .A(n53259), .Z(n53257) );
  XNOR U62848 ( .A(n53160), .B(n53260), .Z(n53166) );
  XNOR U62849 ( .A(n53159), .B(n53161), .Z(n53260) );
  NAND U62850 ( .A(n53261), .B(n53262), .Z(n53161) );
  OR U62851 ( .A(n53263), .B(n53264), .Z(n53262) );
  OR U62852 ( .A(n53265), .B(n53266), .Z(n53261) );
  NAND U62853 ( .A(n53267), .B(n53268), .Z(n53159) );
  OR U62854 ( .A(n53269), .B(n53270), .Z(n53268) );
  OR U62855 ( .A(n53271), .B(n53272), .Z(n53267) );
  ANDN U62856 ( .B(n53273), .A(n53274), .Z(n53160) );
  IV U62857 ( .A(n53275), .Z(n53273) );
  XNOR U62858 ( .A(n53240), .B(n53239), .Z(N60683) );
  XOR U62859 ( .A(n53259), .B(n53258), .Z(n53239) );
  XNOR U62860 ( .A(n53274), .B(n53275), .Z(n53258) );
  XNOR U62861 ( .A(n53269), .B(n53270), .Z(n53275) );
  XNOR U62862 ( .A(n53271), .B(n53272), .Z(n53270) );
  XNOR U62863 ( .A(y[181]), .B(x[181]), .Z(n53272) );
  XNOR U62864 ( .A(y[182]), .B(x[182]), .Z(n53271) );
  XNOR U62865 ( .A(y[180]), .B(x[180]), .Z(n53269) );
  XNOR U62866 ( .A(n53263), .B(n53264), .Z(n53274) );
  XNOR U62867 ( .A(y[177]), .B(x[177]), .Z(n53264) );
  XNOR U62868 ( .A(n53265), .B(n53266), .Z(n53263) );
  XNOR U62869 ( .A(y[178]), .B(x[178]), .Z(n53266) );
  XNOR U62870 ( .A(y[179]), .B(x[179]), .Z(n53265) );
  XNOR U62871 ( .A(n53256), .B(n53255), .Z(n53259) );
  XNOR U62872 ( .A(n53251), .B(n53252), .Z(n53255) );
  XNOR U62873 ( .A(y[174]), .B(x[174]), .Z(n53252) );
  XNOR U62874 ( .A(n53253), .B(n53254), .Z(n53251) );
  XNOR U62875 ( .A(y[175]), .B(x[175]), .Z(n53254) );
  XNOR U62876 ( .A(y[176]), .B(x[176]), .Z(n53253) );
  XNOR U62877 ( .A(n53245), .B(n53246), .Z(n53256) );
  XNOR U62878 ( .A(y[171]), .B(x[171]), .Z(n53246) );
  XNOR U62879 ( .A(n53247), .B(n53248), .Z(n53245) );
  XNOR U62880 ( .A(y[172]), .B(x[172]), .Z(n53248) );
  XNOR U62881 ( .A(y[173]), .B(x[173]), .Z(n53247) );
  XOR U62882 ( .A(n53221), .B(n53222), .Z(n53240) );
  XNOR U62883 ( .A(n53237), .B(n53238), .Z(n53222) );
  XNOR U62884 ( .A(n53232), .B(n53233), .Z(n53238) );
  XNOR U62885 ( .A(n53234), .B(n53235), .Z(n53233) );
  XNOR U62886 ( .A(y[169]), .B(x[169]), .Z(n53235) );
  XNOR U62887 ( .A(y[170]), .B(x[170]), .Z(n53234) );
  XNOR U62888 ( .A(y[168]), .B(x[168]), .Z(n53232) );
  XNOR U62889 ( .A(n53226), .B(n53227), .Z(n53237) );
  XNOR U62890 ( .A(y[165]), .B(x[165]), .Z(n53227) );
  XNOR U62891 ( .A(n53228), .B(n53229), .Z(n53226) );
  XNOR U62892 ( .A(y[166]), .B(x[166]), .Z(n53229) );
  XNOR U62893 ( .A(y[167]), .B(x[167]), .Z(n53228) );
  XOR U62894 ( .A(n53220), .B(n53219), .Z(n53221) );
  XNOR U62895 ( .A(n53215), .B(n53216), .Z(n53219) );
  XNOR U62896 ( .A(y[162]), .B(x[162]), .Z(n53216) );
  XNOR U62897 ( .A(n53217), .B(n53218), .Z(n53215) );
  XNOR U62898 ( .A(y[163]), .B(x[163]), .Z(n53218) );
  XNOR U62899 ( .A(y[164]), .B(x[164]), .Z(n53217) );
  XNOR U62900 ( .A(n53209), .B(n53210), .Z(n53220) );
  XNOR U62901 ( .A(y[159]), .B(x[159]), .Z(n53210) );
  XNOR U62902 ( .A(n53211), .B(n53212), .Z(n53209) );
  XNOR U62903 ( .A(y[160]), .B(x[160]), .Z(n53212) );
  XNOR U62904 ( .A(y[161]), .B(x[161]), .Z(n53211) );
  NAND U62905 ( .A(n53276), .B(n53277), .Z(N60674) );
  NANDN U62906 ( .A(n53278), .B(n53279), .Z(n53277) );
  OR U62907 ( .A(n53280), .B(n53281), .Z(n53279) );
  NAND U62908 ( .A(n53280), .B(n53281), .Z(n53276) );
  XOR U62909 ( .A(n53280), .B(n53282), .Z(N60673) );
  XNOR U62910 ( .A(n53278), .B(n53281), .Z(n53282) );
  AND U62911 ( .A(n53283), .B(n53284), .Z(n53281) );
  NANDN U62912 ( .A(n53285), .B(n53286), .Z(n53284) );
  NANDN U62913 ( .A(n53287), .B(n53288), .Z(n53286) );
  NANDN U62914 ( .A(n53288), .B(n53287), .Z(n53283) );
  NAND U62915 ( .A(n53289), .B(n53290), .Z(n53278) );
  NANDN U62916 ( .A(n53291), .B(n53292), .Z(n53290) );
  OR U62917 ( .A(n53293), .B(n53294), .Z(n53292) );
  NAND U62918 ( .A(n53294), .B(n53293), .Z(n53289) );
  AND U62919 ( .A(n53295), .B(n53296), .Z(n53280) );
  NANDN U62920 ( .A(n53297), .B(n53298), .Z(n53296) );
  NANDN U62921 ( .A(n53299), .B(n53300), .Z(n53298) );
  NANDN U62922 ( .A(n53300), .B(n53299), .Z(n53295) );
  XOR U62923 ( .A(n53294), .B(n53301), .Z(N60672) );
  XOR U62924 ( .A(n53291), .B(n53293), .Z(n53301) );
  XNOR U62925 ( .A(n53287), .B(n53302), .Z(n53293) );
  XNOR U62926 ( .A(n53285), .B(n53288), .Z(n53302) );
  NAND U62927 ( .A(n53303), .B(n53304), .Z(n53288) );
  NAND U62928 ( .A(n53305), .B(n53306), .Z(n53304) );
  OR U62929 ( .A(n53307), .B(n53308), .Z(n53305) );
  NANDN U62930 ( .A(n53309), .B(n53307), .Z(n53303) );
  IV U62931 ( .A(n53308), .Z(n53309) );
  NAND U62932 ( .A(n53310), .B(n53311), .Z(n53285) );
  NAND U62933 ( .A(n53312), .B(n53313), .Z(n53311) );
  NANDN U62934 ( .A(n53314), .B(n53315), .Z(n53312) );
  NANDN U62935 ( .A(n53315), .B(n53314), .Z(n53310) );
  AND U62936 ( .A(n53316), .B(n53317), .Z(n53287) );
  NAND U62937 ( .A(n53318), .B(n53319), .Z(n53317) );
  OR U62938 ( .A(n53320), .B(n53321), .Z(n53318) );
  NANDN U62939 ( .A(n53322), .B(n53320), .Z(n53316) );
  NAND U62940 ( .A(n53323), .B(n53324), .Z(n53291) );
  NANDN U62941 ( .A(n53325), .B(n53326), .Z(n53324) );
  OR U62942 ( .A(n53327), .B(n53328), .Z(n53326) );
  NANDN U62943 ( .A(n53329), .B(n53327), .Z(n53323) );
  IV U62944 ( .A(n53328), .Z(n53329) );
  XNOR U62945 ( .A(n53299), .B(n53330), .Z(n53294) );
  XNOR U62946 ( .A(n53297), .B(n53300), .Z(n53330) );
  NAND U62947 ( .A(n53331), .B(n53332), .Z(n53300) );
  NAND U62948 ( .A(n53333), .B(n53334), .Z(n53332) );
  OR U62949 ( .A(n53335), .B(n53336), .Z(n53333) );
  NANDN U62950 ( .A(n53337), .B(n53335), .Z(n53331) );
  IV U62951 ( .A(n53336), .Z(n53337) );
  NAND U62952 ( .A(n53338), .B(n53339), .Z(n53297) );
  NAND U62953 ( .A(n53340), .B(n53341), .Z(n53339) );
  NANDN U62954 ( .A(n53342), .B(n53343), .Z(n53340) );
  NANDN U62955 ( .A(n53343), .B(n53342), .Z(n53338) );
  AND U62956 ( .A(n53344), .B(n53345), .Z(n53299) );
  NAND U62957 ( .A(n53346), .B(n53347), .Z(n53345) );
  OR U62958 ( .A(n53348), .B(n53349), .Z(n53346) );
  NANDN U62959 ( .A(n53350), .B(n53348), .Z(n53344) );
  XNOR U62960 ( .A(n53325), .B(n53351), .Z(N60671) );
  XOR U62961 ( .A(n53327), .B(n53328), .Z(n53351) );
  XNOR U62962 ( .A(n53341), .B(n53352), .Z(n53328) );
  XOR U62963 ( .A(n53342), .B(n53343), .Z(n53352) );
  XOR U62964 ( .A(n53348), .B(n53353), .Z(n53343) );
  XOR U62965 ( .A(n53347), .B(n53350), .Z(n53353) );
  IV U62966 ( .A(n53349), .Z(n53350) );
  NAND U62967 ( .A(n53354), .B(n53355), .Z(n53349) );
  OR U62968 ( .A(n53356), .B(n53357), .Z(n53355) );
  OR U62969 ( .A(n53358), .B(n53359), .Z(n53354) );
  NAND U62970 ( .A(n53360), .B(n53361), .Z(n53347) );
  OR U62971 ( .A(n53362), .B(n53363), .Z(n53361) );
  OR U62972 ( .A(n53364), .B(n53365), .Z(n53360) );
  NOR U62973 ( .A(n53366), .B(n53367), .Z(n53348) );
  ANDN U62974 ( .B(n53368), .A(n53369), .Z(n53342) );
  XNOR U62975 ( .A(n53335), .B(n53370), .Z(n53341) );
  XNOR U62976 ( .A(n53334), .B(n53336), .Z(n53370) );
  NAND U62977 ( .A(n53371), .B(n53372), .Z(n53336) );
  OR U62978 ( .A(n53373), .B(n53374), .Z(n53372) );
  OR U62979 ( .A(n53375), .B(n53376), .Z(n53371) );
  NAND U62980 ( .A(n53377), .B(n53378), .Z(n53334) );
  OR U62981 ( .A(n53379), .B(n53380), .Z(n53378) );
  OR U62982 ( .A(n53381), .B(n53382), .Z(n53377) );
  ANDN U62983 ( .B(n53383), .A(n53384), .Z(n53335) );
  IV U62984 ( .A(n53385), .Z(n53383) );
  ANDN U62985 ( .B(n53386), .A(n53387), .Z(n53327) );
  XOR U62986 ( .A(n53313), .B(n53388), .Z(n53325) );
  XOR U62987 ( .A(n53314), .B(n53315), .Z(n53388) );
  XOR U62988 ( .A(n53320), .B(n53389), .Z(n53315) );
  XOR U62989 ( .A(n53319), .B(n53322), .Z(n53389) );
  IV U62990 ( .A(n53321), .Z(n53322) );
  NAND U62991 ( .A(n53390), .B(n53391), .Z(n53321) );
  OR U62992 ( .A(n53392), .B(n53393), .Z(n53391) );
  OR U62993 ( .A(n53394), .B(n53395), .Z(n53390) );
  NAND U62994 ( .A(n53396), .B(n53397), .Z(n53319) );
  OR U62995 ( .A(n53398), .B(n53399), .Z(n53397) );
  OR U62996 ( .A(n53400), .B(n53401), .Z(n53396) );
  NOR U62997 ( .A(n53402), .B(n53403), .Z(n53320) );
  ANDN U62998 ( .B(n53404), .A(n53405), .Z(n53314) );
  IV U62999 ( .A(n53406), .Z(n53404) );
  XNOR U63000 ( .A(n53307), .B(n53407), .Z(n53313) );
  XNOR U63001 ( .A(n53306), .B(n53308), .Z(n53407) );
  NAND U63002 ( .A(n53408), .B(n53409), .Z(n53308) );
  OR U63003 ( .A(n53410), .B(n53411), .Z(n53409) );
  OR U63004 ( .A(n53412), .B(n53413), .Z(n53408) );
  NAND U63005 ( .A(n53414), .B(n53415), .Z(n53306) );
  OR U63006 ( .A(n53416), .B(n53417), .Z(n53415) );
  OR U63007 ( .A(n53418), .B(n53419), .Z(n53414) );
  ANDN U63008 ( .B(n53420), .A(n53421), .Z(n53307) );
  IV U63009 ( .A(n53422), .Z(n53420) );
  XNOR U63010 ( .A(n53387), .B(n53386), .Z(N60670) );
  XOR U63011 ( .A(n53406), .B(n53405), .Z(n53386) );
  XNOR U63012 ( .A(n53421), .B(n53422), .Z(n53405) );
  XNOR U63013 ( .A(n53416), .B(n53417), .Z(n53422) );
  XNOR U63014 ( .A(n53418), .B(n53419), .Z(n53417) );
  XNOR U63015 ( .A(y[157]), .B(x[157]), .Z(n53419) );
  XNOR U63016 ( .A(y[158]), .B(x[158]), .Z(n53418) );
  XNOR U63017 ( .A(y[156]), .B(x[156]), .Z(n53416) );
  XNOR U63018 ( .A(n53410), .B(n53411), .Z(n53421) );
  XNOR U63019 ( .A(y[153]), .B(x[153]), .Z(n53411) );
  XNOR U63020 ( .A(n53412), .B(n53413), .Z(n53410) );
  XNOR U63021 ( .A(y[154]), .B(x[154]), .Z(n53413) );
  XNOR U63022 ( .A(y[155]), .B(x[155]), .Z(n53412) );
  XNOR U63023 ( .A(n53403), .B(n53402), .Z(n53406) );
  XNOR U63024 ( .A(n53398), .B(n53399), .Z(n53402) );
  XNOR U63025 ( .A(y[150]), .B(x[150]), .Z(n53399) );
  XNOR U63026 ( .A(n53400), .B(n53401), .Z(n53398) );
  XNOR U63027 ( .A(y[151]), .B(x[151]), .Z(n53401) );
  XNOR U63028 ( .A(y[152]), .B(x[152]), .Z(n53400) );
  XNOR U63029 ( .A(n53392), .B(n53393), .Z(n53403) );
  XNOR U63030 ( .A(y[147]), .B(x[147]), .Z(n53393) );
  XNOR U63031 ( .A(n53394), .B(n53395), .Z(n53392) );
  XNOR U63032 ( .A(y[148]), .B(x[148]), .Z(n53395) );
  XNOR U63033 ( .A(y[149]), .B(x[149]), .Z(n53394) );
  XOR U63034 ( .A(n53368), .B(n53369), .Z(n53387) );
  XNOR U63035 ( .A(n53384), .B(n53385), .Z(n53369) );
  XNOR U63036 ( .A(n53379), .B(n53380), .Z(n53385) );
  XNOR U63037 ( .A(n53381), .B(n53382), .Z(n53380) );
  XNOR U63038 ( .A(y[145]), .B(x[145]), .Z(n53382) );
  XNOR U63039 ( .A(y[146]), .B(x[146]), .Z(n53381) );
  XNOR U63040 ( .A(y[144]), .B(x[144]), .Z(n53379) );
  XNOR U63041 ( .A(n53373), .B(n53374), .Z(n53384) );
  XNOR U63042 ( .A(y[141]), .B(x[141]), .Z(n53374) );
  XNOR U63043 ( .A(n53375), .B(n53376), .Z(n53373) );
  XNOR U63044 ( .A(y[142]), .B(x[142]), .Z(n53376) );
  XNOR U63045 ( .A(y[143]), .B(x[143]), .Z(n53375) );
  XOR U63046 ( .A(n53367), .B(n53366), .Z(n53368) );
  XNOR U63047 ( .A(n53362), .B(n53363), .Z(n53366) );
  XNOR U63048 ( .A(y[138]), .B(x[138]), .Z(n53363) );
  XNOR U63049 ( .A(n53364), .B(n53365), .Z(n53362) );
  XNOR U63050 ( .A(y[139]), .B(x[139]), .Z(n53365) );
  XNOR U63051 ( .A(y[140]), .B(x[140]), .Z(n53364) );
  XNOR U63052 ( .A(n53356), .B(n53357), .Z(n53367) );
  XNOR U63053 ( .A(y[135]), .B(x[135]), .Z(n53357) );
  XNOR U63054 ( .A(n53358), .B(n53359), .Z(n53356) );
  XNOR U63055 ( .A(y[136]), .B(x[136]), .Z(n53359) );
  XNOR U63056 ( .A(y[137]), .B(x[137]), .Z(n53358) );
  NAND U63057 ( .A(n53423), .B(n53424), .Z(N60661) );
  NANDN U63058 ( .A(n53425), .B(n53426), .Z(n53424) );
  OR U63059 ( .A(n53427), .B(n53428), .Z(n53426) );
  NAND U63060 ( .A(n53427), .B(n53428), .Z(n53423) );
  XOR U63061 ( .A(n53427), .B(n53429), .Z(N60660) );
  XNOR U63062 ( .A(n53425), .B(n53428), .Z(n53429) );
  AND U63063 ( .A(n53430), .B(n53431), .Z(n53428) );
  NANDN U63064 ( .A(n53432), .B(n53433), .Z(n53431) );
  NANDN U63065 ( .A(n53434), .B(n53435), .Z(n53433) );
  NANDN U63066 ( .A(n53435), .B(n53434), .Z(n53430) );
  NAND U63067 ( .A(n53436), .B(n53437), .Z(n53425) );
  NANDN U63068 ( .A(n53438), .B(n53439), .Z(n53437) );
  OR U63069 ( .A(n53440), .B(n53441), .Z(n53439) );
  NAND U63070 ( .A(n53441), .B(n53440), .Z(n53436) );
  AND U63071 ( .A(n53442), .B(n53443), .Z(n53427) );
  NANDN U63072 ( .A(n53444), .B(n53445), .Z(n53443) );
  NANDN U63073 ( .A(n53446), .B(n53447), .Z(n53445) );
  NANDN U63074 ( .A(n53447), .B(n53446), .Z(n53442) );
  XOR U63075 ( .A(n53441), .B(n53448), .Z(N60659) );
  XOR U63076 ( .A(n53438), .B(n53440), .Z(n53448) );
  XNOR U63077 ( .A(n53434), .B(n53449), .Z(n53440) );
  XNOR U63078 ( .A(n53432), .B(n53435), .Z(n53449) );
  NAND U63079 ( .A(n53450), .B(n53451), .Z(n53435) );
  NAND U63080 ( .A(n53452), .B(n53453), .Z(n53451) );
  OR U63081 ( .A(n53454), .B(n53455), .Z(n53452) );
  NANDN U63082 ( .A(n53456), .B(n53454), .Z(n53450) );
  IV U63083 ( .A(n53455), .Z(n53456) );
  NAND U63084 ( .A(n53457), .B(n53458), .Z(n53432) );
  NAND U63085 ( .A(n53459), .B(n53460), .Z(n53458) );
  NANDN U63086 ( .A(n53461), .B(n53462), .Z(n53459) );
  NANDN U63087 ( .A(n53462), .B(n53461), .Z(n53457) );
  AND U63088 ( .A(n53463), .B(n53464), .Z(n53434) );
  NAND U63089 ( .A(n53465), .B(n53466), .Z(n53464) );
  OR U63090 ( .A(n53467), .B(n53468), .Z(n53465) );
  NANDN U63091 ( .A(n53469), .B(n53467), .Z(n53463) );
  NAND U63092 ( .A(n53470), .B(n53471), .Z(n53438) );
  NANDN U63093 ( .A(n53472), .B(n53473), .Z(n53471) );
  OR U63094 ( .A(n53474), .B(n53475), .Z(n53473) );
  NANDN U63095 ( .A(n53476), .B(n53474), .Z(n53470) );
  IV U63096 ( .A(n53475), .Z(n53476) );
  XNOR U63097 ( .A(n53446), .B(n53477), .Z(n53441) );
  XNOR U63098 ( .A(n53444), .B(n53447), .Z(n53477) );
  NAND U63099 ( .A(n53478), .B(n53479), .Z(n53447) );
  NAND U63100 ( .A(n53480), .B(n53481), .Z(n53479) );
  OR U63101 ( .A(n53482), .B(n53483), .Z(n53480) );
  NANDN U63102 ( .A(n53484), .B(n53482), .Z(n53478) );
  IV U63103 ( .A(n53483), .Z(n53484) );
  NAND U63104 ( .A(n53485), .B(n53486), .Z(n53444) );
  NAND U63105 ( .A(n53487), .B(n53488), .Z(n53486) );
  NANDN U63106 ( .A(n53489), .B(n53490), .Z(n53487) );
  NANDN U63107 ( .A(n53490), .B(n53489), .Z(n53485) );
  AND U63108 ( .A(n53491), .B(n53492), .Z(n53446) );
  NAND U63109 ( .A(n53493), .B(n53494), .Z(n53492) );
  OR U63110 ( .A(n53495), .B(n53496), .Z(n53493) );
  NANDN U63111 ( .A(n53497), .B(n53495), .Z(n53491) );
  XNOR U63112 ( .A(n53472), .B(n53498), .Z(N60658) );
  XOR U63113 ( .A(n53474), .B(n53475), .Z(n53498) );
  XNOR U63114 ( .A(n53488), .B(n53499), .Z(n53475) );
  XOR U63115 ( .A(n53489), .B(n53490), .Z(n53499) );
  XOR U63116 ( .A(n53495), .B(n53500), .Z(n53490) );
  XOR U63117 ( .A(n53494), .B(n53497), .Z(n53500) );
  IV U63118 ( .A(n53496), .Z(n53497) );
  NAND U63119 ( .A(n53501), .B(n53502), .Z(n53496) );
  OR U63120 ( .A(n53503), .B(n53504), .Z(n53502) );
  OR U63121 ( .A(n53505), .B(n53506), .Z(n53501) );
  NAND U63122 ( .A(n53507), .B(n53508), .Z(n53494) );
  OR U63123 ( .A(n53509), .B(n53510), .Z(n53508) );
  OR U63124 ( .A(n53511), .B(n53512), .Z(n53507) );
  NOR U63125 ( .A(n53513), .B(n53514), .Z(n53495) );
  ANDN U63126 ( .B(n53515), .A(n53516), .Z(n53489) );
  XNOR U63127 ( .A(n53482), .B(n53517), .Z(n53488) );
  XNOR U63128 ( .A(n53481), .B(n53483), .Z(n53517) );
  NAND U63129 ( .A(n53518), .B(n53519), .Z(n53483) );
  OR U63130 ( .A(n53520), .B(n53521), .Z(n53519) );
  OR U63131 ( .A(n53522), .B(n53523), .Z(n53518) );
  NAND U63132 ( .A(n53524), .B(n53525), .Z(n53481) );
  OR U63133 ( .A(n53526), .B(n53527), .Z(n53525) );
  OR U63134 ( .A(n53528), .B(n53529), .Z(n53524) );
  ANDN U63135 ( .B(n53530), .A(n53531), .Z(n53482) );
  IV U63136 ( .A(n53532), .Z(n53530) );
  ANDN U63137 ( .B(n53533), .A(n53534), .Z(n53474) );
  XOR U63138 ( .A(n53460), .B(n53535), .Z(n53472) );
  XOR U63139 ( .A(n53461), .B(n53462), .Z(n53535) );
  XOR U63140 ( .A(n53467), .B(n53536), .Z(n53462) );
  XOR U63141 ( .A(n53466), .B(n53469), .Z(n53536) );
  IV U63142 ( .A(n53468), .Z(n53469) );
  NAND U63143 ( .A(n53537), .B(n53538), .Z(n53468) );
  OR U63144 ( .A(n53539), .B(n53540), .Z(n53538) );
  OR U63145 ( .A(n53541), .B(n53542), .Z(n53537) );
  NAND U63146 ( .A(n53543), .B(n53544), .Z(n53466) );
  OR U63147 ( .A(n53545), .B(n53546), .Z(n53544) );
  OR U63148 ( .A(n53547), .B(n53548), .Z(n53543) );
  NOR U63149 ( .A(n53549), .B(n53550), .Z(n53467) );
  ANDN U63150 ( .B(n53551), .A(n53552), .Z(n53461) );
  IV U63151 ( .A(n53553), .Z(n53551) );
  XNOR U63152 ( .A(n53454), .B(n53554), .Z(n53460) );
  XNOR U63153 ( .A(n53453), .B(n53455), .Z(n53554) );
  NAND U63154 ( .A(n53555), .B(n53556), .Z(n53455) );
  OR U63155 ( .A(n53557), .B(n53558), .Z(n53556) );
  OR U63156 ( .A(n53559), .B(n53560), .Z(n53555) );
  NAND U63157 ( .A(n53561), .B(n53562), .Z(n53453) );
  OR U63158 ( .A(n53563), .B(n53564), .Z(n53562) );
  OR U63159 ( .A(n53565), .B(n53566), .Z(n53561) );
  ANDN U63160 ( .B(n53567), .A(n53568), .Z(n53454) );
  IV U63161 ( .A(n53569), .Z(n53567) );
  XNOR U63162 ( .A(n53534), .B(n53533), .Z(N60657) );
  XOR U63163 ( .A(n53553), .B(n53552), .Z(n53533) );
  XNOR U63164 ( .A(n53568), .B(n53569), .Z(n53552) );
  XNOR U63165 ( .A(n53563), .B(n53564), .Z(n53569) );
  XNOR U63166 ( .A(n53565), .B(n53566), .Z(n53564) );
  XNOR U63167 ( .A(y[133]), .B(x[133]), .Z(n53566) );
  XNOR U63168 ( .A(y[134]), .B(x[134]), .Z(n53565) );
  XNOR U63169 ( .A(y[132]), .B(x[132]), .Z(n53563) );
  XNOR U63170 ( .A(n53557), .B(n53558), .Z(n53568) );
  XNOR U63171 ( .A(y[129]), .B(x[129]), .Z(n53558) );
  XNOR U63172 ( .A(n53559), .B(n53560), .Z(n53557) );
  XNOR U63173 ( .A(y[130]), .B(x[130]), .Z(n53560) );
  XNOR U63174 ( .A(y[131]), .B(x[131]), .Z(n53559) );
  XNOR U63175 ( .A(n53550), .B(n53549), .Z(n53553) );
  XNOR U63176 ( .A(n53545), .B(n53546), .Z(n53549) );
  XNOR U63177 ( .A(y[126]), .B(x[126]), .Z(n53546) );
  XNOR U63178 ( .A(n53547), .B(n53548), .Z(n53545) );
  XNOR U63179 ( .A(y[127]), .B(x[127]), .Z(n53548) );
  XNOR U63180 ( .A(y[128]), .B(x[128]), .Z(n53547) );
  XNOR U63181 ( .A(n53539), .B(n53540), .Z(n53550) );
  XNOR U63182 ( .A(y[123]), .B(x[123]), .Z(n53540) );
  XNOR U63183 ( .A(n53541), .B(n53542), .Z(n53539) );
  XNOR U63184 ( .A(y[124]), .B(x[124]), .Z(n53542) );
  XNOR U63185 ( .A(y[125]), .B(x[125]), .Z(n53541) );
  XOR U63186 ( .A(n53515), .B(n53516), .Z(n53534) );
  XNOR U63187 ( .A(n53531), .B(n53532), .Z(n53516) );
  XNOR U63188 ( .A(n53526), .B(n53527), .Z(n53532) );
  XNOR U63189 ( .A(n53528), .B(n53529), .Z(n53527) );
  XNOR U63190 ( .A(y[121]), .B(x[121]), .Z(n53529) );
  XNOR U63191 ( .A(y[122]), .B(x[122]), .Z(n53528) );
  XNOR U63192 ( .A(y[120]), .B(x[120]), .Z(n53526) );
  XNOR U63193 ( .A(n53520), .B(n53521), .Z(n53531) );
  XNOR U63194 ( .A(y[117]), .B(x[117]), .Z(n53521) );
  XNOR U63195 ( .A(n53522), .B(n53523), .Z(n53520) );
  XNOR U63196 ( .A(y[118]), .B(x[118]), .Z(n53523) );
  XNOR U63197 ( .A(y[119]), .B(x[119]), .Z(n53522) );
  XOR U63198 ( .A(n53514), .B(n53513), .Z(n53515) );
  XNOR U63199 ( .A(n53509), .B(n53510), .Z(n53513) );
  XNOR U63200 ( .A(y[114]), .B(x[114]), .Z(n53510) );
  XNOR U63201 ( .A(n53511), .B(n53512), .Z(n53509) );
  XNOR U63202 ( .A(y[115]), .B(x[115]), .Z(n53512) );
  XNOR U63203 ( .A(y[116]), .B(x[116]), .Z(n53511) );
  XNOR U63204 ( .A(n53503), .B(n53504), .Z(n53514) );
  XNOR U63205 ( .A(y[111]), .B(x[111]), .Z(n53504) );
  XNOR U63206 ( .A(n53505), .B(n53506), .Z(n53503) );
  XNOR U63207 ( .A(y[112]), .B(x[112]), .Z(n53506) );
  XNOR U63208 ( .A(y[113]), .B(x[113]), .Z(n53505) );
  NAND U63209 ( .A(n53570), .B(n53571), .Z(N60648) );
  NANDN U63210 ( .A(n53572), .B(n53573), .Z(n53571) );
  OR U63211 ( .A(n53574), .B(n53575), .Z(n53573) );
  NAND U63212 ( .A(n53574), .B(n53575), .Z(n53570) );
  XOR U63213 ( .A(n53574), .B(n53576), .Z(N60647) );
  XNOR U63214 ( .A(n53572), .B(n53575), .Z(n53576) );
  AND U63215 ( .A(n53577), .B(n53578), .Z(n53575) );
  NANDN U63216 ( .A(n53579), .B(n53580), .Z(n53578) );
  NANDN U63217 ( .A(n53581), .B(n53582), .Z(n53580) );
  NANDN U63218 ( .A(n53582), .B(n53581), .Z(n53577) );
  NAND U63219 ( .A(n53583), .B(n53584), .Z(n53572) );
  NANDN U63220 ( .A(n53585), .B(n53586), .Z(n53584) );
  OR U63221 ( .A(n53587), .B(n53588), .Z(n53586) );
  NAND U63222 ( .A(n53588), .B(n53587), .Z(n53583) );
  AND U63223 ( .A(n53589), .B(n53590), .Z(n53574) );
  NANDN U63224 ( .A(n53591), .B(n53592), .Z(n53590) );
  NANDN U63225 ( .A(n53593), .B(n53594), .Z(n53592) );
  NANDN U63226 ( .A(n53594), .B(n53593), .Z(n53589) );
  XOR U63227 ( .A(n53588), .B(n53595), .Z(N60646) );
  XOR U63228 ( .A(n53585), .B(n53587), .Z(n53595) );
  XNOR U63229 ( .A(n53581), .B(n53596), .Z(n53587) );
  XNOR U63230 ( .A(n53579), .B(n53582), .Z(n53596) );
  NAND U63231 ( .A(n53597), .B(n53598), .Z(n53582) );
  NAND U63232 ( .A(n53599), .B(n53600), .Z(n53598) );
  OR U63233 ( .A(n53601), .B(n53602), .Z(n53599) );
  NANDN U63234 ( .A(n53603), .B(n53601), .Z(n53597) );
  IV U63235 ( .A(n53602), .Z(n53603) );
  NAND U63236 ( .A(n53604), .B(n53605), .Z(n53579) );
  NAND U63237 ( .A(n53606), .B(n53607), .Z(n53605) );
  NANDN U63238 ( .A(n53608), .B(n53609), .Z(n53606) );
  NANDN U63239 ( .A(n53609), .B(n53608), .Z(n53604) );
  AND U63240 ( .A(n53610), .B(n53611), .Z(n53581) );
  NAND U63241 ( .A(n53612), .B(n53613), .Z(n53611) );
  OR U63242 ( .A(n53614), .B(n53615), .Z(n53612) );
  NANDN U63243 ( .A(n53616), .B(n53614), .Z(n53610) );
  NAND U63244 ( .A(n53617), .B(n53618), .Z(n53585) );
  NANDN U63245 ( .A(n53619), .B(n53620), .Z(n53618) );
  OR U63246 ( .A(n53621), .B(n53622), .Z(n53620) );
  NANDN U63247 ( .A(n53623), .B(n53621), .Z(n53617) );
  IV U63248 ( .A(n53622), .Z(n53623) );
  XNOR U63249 ( .A(n53593), .B(n53624), .Z(n53588) );
  XNOR U63250 ( .A(n53591), .B(n53594), .Z(n53624) );
  NAND U63251 ( .A(n53625), .B(n53626), .Z(n53594) );
  NAND U63252 ( .A(n53627), .B(n53628), .Z(n53626) );
  OR U63253 ( .A(n53629), .B(n53630), .Z(n53627) );
  NANDN U63254 ( .A(n53631), .B(n53629), .Z(n53625) );
  IV U63255 ( .A(n53630), .Z(n53631) );
  NAND U63256 ( .A(n53632), .B(n53633), .Z(n53591) );
  NAND U63257 ( .A(n53634), .B(n53635), .Z(n53633) );
  NANDN U63258 ( .A(n53636), .B(n53637), .Z(n53634) );
  NANDN U63259 ( .A(n53637), .B(n53636), .Z(n53632) );
  AND U63260 ( .A(n53638), .B(n53639), .Z(n53593) );
  NAND U63261 ( .A(n53640), .B(n53641), .Z(n53639) );
  OR U63262 ( .A(n53642), .B(n53643), .Z(n53640) );
  NANDN U63263 ( .A(n53644), .B(n53642), .Z(n53638) );
  XNOR U63264 ( .A(n53619), .B(n53645), .Z(N60645) );
  XOR U63265 ( .A(n53621), .B(n53622), .Z(n53645) );
  XNOR U63266 ( .A(n53635), .B(n53646), .Z(n53622) );
  XOR U63267 ( .A(n53636), .B(n53637), .Z(n53646) );
  XOR U63268 ( .A(n53642), .B(n53647), .Z(n53637) );
  XOR U63269 ( .A(n53641), .B(n53644), .Z(n53647) );
  IV U63270 ( .A(n53643), .Z(n53644) );
  NAND U63271 ( .A(n53648), .B(n53649), .Z(n53643) );
  OR U63272 ( .A(n53650), .B(n53651), .Z(n53649) );
  OR U63273 ( .A(n53652), .B(n53653), .Z(n53648) );
  NAND U63274 ( .A(n53654), .B(n53655), .Z(n53641) );
  OR U63275 ( .A(n53656), .B(n53657), .Z(n53655) );
  OR U63276 ( .A(n53658), .B(n53659), .Z(n53654) );
  NOR U63277 ( .A(n53660), .B(n53661), .Z(n53642) );
  ANDN U63278 ( .B(n53662), .A(n53663), .Z(n53636) );
  XNOR U63279 ( .A(n53629), .B(n53664), .Z(n53635) );
  XNOR U63280 ( .A(n53628), .B(n53630), .Z(n53664) );
  NAND U63281 ( .A(n53665), .B(n53666), .Z(n53630) );
  OR U63282 ( .A(n53667), .B(n53668), .Z(n53666) );
  OR U63283 ( .A(n53669), .B(n53670), .Z(n53665) );
  NAND U63284 ( .A(n53671), .B(n53672), .Z(n53628) );
  OR U63285 ( .A(n53673), .B(n53674), .Z(n53672) );
  OR U63286 ( .A(n53675), .B(n53676), .Z(n53671) );
  ANDN U63287 ( .B(n53677), .A(n53678), .Z(n53629) );
  IV U63288 ( .A(n53679), .Z(n53677) );
  ANDN U63289 ( .B(n53680), .A(n53681), .Z(n53621) );
  XOR U63290 ( .A(n53607), .B(n53682), .Z(n53619) );
  XOR U63291 ( .A(n53608), .B(n53609), .Z(n53682) );
  XOR U63292 ( .A(n53614), .B(n53683), .Z(n53609) );
  XOR U63293 ( .A(n53613), .B(n53616), .Z(n53683) );
  IV U63294 ( .A(n53615), .Z(n53616) );
  NAND U63295 ( .A(n53684), .B(n53685), .Z(n53615) );
  OR U63296 ( .A(n53686), .B(n53687), .Z(n53685) );
  OR U63297 ( .A(n53688), .B(n53689), .Z(n53684) );
  NAND U63298 ( .A(n53690), .B(n53691), .Z(n53613) );
  OR U63299 ( .A(n53692), .B(n53693), .Z(n53691) );
  OR U63300 ( .A(n53694), .B(n53695), .Z(n53690) );
  NOR U63301 ( .A(n53696), .B(n53697), .Z(n53614) );
  ANDN U63302 ( .B(n53698), .A(n53699), .Z(n53608) );
  IV U63303 ( .A(n53700), .Z(n53698) );
  XNOR U63304 ( .A(n53601), .B(n53701), .Z(n53607) );
  XNOR U63305 ( .A(n53600), .B(n53602), .Z(n53701) );
  NAND U63306 ( .A(n53702), .B(n53703), .Z(n53602) );
  OR U63307 ( .A(n53704), .B(n53705), .Z(n53703) );
  OR U63308 ( .A(n53706), .B(n53707), .Z(n53702) );
  NAND U63309 ( .A(n53708), .B(n53709), .Z(n53600) );
  OR U63310 ( .A(n53710), .B(n53711), .Z(n53709) );
  OR U63311 ( .A(n53712), .B(n53713), .Z(n53708) );
  ANDN U63312 ( .B(n53714), .A(n53715), .Z(n53601) );
  IV U63313 ( .A(n53716), .Z(n53714) );
  XNOR U63314 ( .A(n53681), .B(n53680), .Z(N60644) );
  XOR U63315 ( .A(n53700), .B(n53699), .Z(n53680) );
  XNOR U63316 ( .A(n53715), .B(n53716), .Z(n53699) );
  XNOR U63317 ( .A(n53710), .B(n53711), .Z(n53716) );
  XNOR U63318 ( .A(n53712), .B(n53713), .Z(n53711) );
  XNOR U63319 ( .A(y[109]), .B(x[109]), .Z(n53713) );
  XNOR U63320 ( .A(y[110]), .B(x[110]), .Z(n53712) );
  XNOR U63321 ( .A(y[108]), .B(x[108]), .Z(n53710) );
  XNOR U63322 ( .A(n53704), .B(n53705), .Z(n53715) );
  XNOR U63323 ( .A(y[105]), .B(x[105]), .Z(n53705) );
  XNOR U63324 ( .A(n53706), .B(n53707), .Z(n53704) );
  XNOR U63325 ( .A(y[106]), .B(x[106]), .Z(n53707) );
  XNOR U63326 ( .A(y[107]), .B(x[107]), .Z(n53706) );
  XNOR U63327 ( .A(n53697), .B(n53696), .Z(n53700) );
  XNOR U63328 ( .A(n53692), .B(n53693), .Z(n53696) );
  XNOR U63329 ( .A(y[102]), .B(x[102]), .Z(n53693) );
  XNOR U63330 ( .A(n53694), .B(n53695), .Z(n53692) );
  XNOR U63331 ( .A(y[103]), .B(x[103]), .Z(n53695) );
  XNOR U63332 ( .A(y[104]), .B(x[104]), .Z(n53694) );
  XNOR U63333 ( .A(n53686), .B(n53687), .Z(n53697) );
  XNOR U63334 ( .A(y[99]), .B(x[99]), .Z(n53687) );
  XNOR U63335 ( .A(n53688), .B(n53689), .Z(n53686) );
  XNOR U63336 ( .A(y[100]), .B(x[100]), .Z(n53689) );
  XNOR U63337 ( .A(y[101]), .B(x[101]), .Z(n53688) );
  XOR U63338 ( .A(n53662), .B(n53663), .Z(n53681) );
  XNOR U63339 ( .A(n53678), .B(n53679), .Z(n53663) );
  XNOR U63340 ( .A(n53673), .B(n53674), .Z(n53679) );
  XNOR U63341 ( .A(n53675), .B(n53676), .Z(n53674) );
  XNOR U63342 ( .A(y[97]), .B(x[97]), .Z(n53676) );
  XNOR U63343 ( .A(y[98]), .B(x[98]), .Z(n53675) );
  XNOR U63344 ( .A(y[96]), .B(x[96]), .Z(n53673) );
  XNOR U63345 ( .A(n53667), .B(n53668), .Z(n53678) );
  XNOR U63346 ( .A(y[93]), .B(x[93]), .Z(n53668) );
  XNOR U63347 ( .A(n53669), .B(n53670), .Z(n53667) );
  XNOR U63348 ( .A(y[94]), .B(x[94]), .Z(n53670) );
  XNOR U63349 ( .A(y[95]), .B(x[95]), .Z(n53669) );
  XOR U63350 ( .A(n53661), .B(n53660), .Z(n53662) );
  XNOR U63351 ( .A(n53656), .B(n53657), .Z(n53660) );
  XNOR U63352 ( .A(y[90]), .B(x[90]), .Z(n53657) );
  XNOR U63353 ( .A(n53658), .B(n53659), .Z(n53656) );
  XNOR U63354 ( .A(y[91]), .B(x[91]), .Z(n53659) );
  XNOR U63355 ( .A(y[92]), .B(x[92]), .Z(n53658) );
  XNOR U63356 ( .A(n53650), .B(n53651), .Z(n53661) );
  XNOR U63357 ( .A(y[87]), .B(x[87]), .Z(n53651) );
  XNOR U63358 ( .A(n53652), .B(n53653), .Z(n53650) );
  XNOR U63359 ( .A(y[88]), .B(x[88]), .Z(n53653) );
  XNOR U63360 ( .A(y[89]), .B(x[89]), .Z(n53652) );
  NAND U63361 ( .A(n53717), .B(n53718), .Z(N60635) );
  NANDN U63362 ( .A(n53719), .B(n53720), .Z(n53718) );
  OR U63363 ( .A(n53721), .B(n53722), .Z(n53720) );
  NAND U63364 ( .A(n53721), .B(n53722), .Z(n53717) );
  XOR U63365 ( .A(n53721), .B(n53723), .Z(N60634) );
  XNOR U63366 ( .A(n53719), .B(n53722), .Z(n53723) );
  AND U63367 ( .A(n53724), .B(n53725), .Z(n53722) );
  NANDN U63368 ( .A(n53726), .B(n53727), .Z(n53725) );
  NANDN U63369 ( .A(n53728), .B(n53729), .Z(n53727) );
  NANDN U63370 ( .A(n53729), .B(n53728), .Z(n53724) );
  NAND U63371 ( .A(n53730), .B(n53731), .Z(n53719) );
  NANDN U63372 ( .A(n53732), .B(n53733), .Z(n53731) );
  OR U63373 ( .A(n53734), .B(n53735), .Z(n53733) );
  NAND U63374 ( .A(n53735), .B(n53734), .Z(n53730) );
  AND U63375 ( .A(n53736), .B(n53737), .Z(n53721) );
  NANDN U63376 ( .A(n53738), .B(n53739), .Z(n53737) );
  NANDN U63377 ( .A(n53740), .B(n53741), .Z(n53739) );
  NANDN U63378 ( .A(n53741), .B(n53740), .Z(n53736) );
  XOR U63379 ( .A(n53735), .B(n53742), .Z(N60633) );
  XOR U63380 ( .A(n53732), .B(n53734), .Z(n53742) );
  XNOR U63381 ( .A(n53728), .B(n53743), .Z(n53734) );
  XNOR U63382 ( .A(n53726), .B(n53729), .Z(n53743) );
  NAND U63383 ( .A(n53744), .B(n53745), .Z(n53729) );
  NAND U63384 ( .A(n53746), .B(n53747), .Z(n53745) );
  OR U63385 ( .A(n53748), .B(n53749), .Z(n53746) );
  NANDN U63386 ( .A(n53750), .B(n53748), .Z(n53744) );
  IV U63387 ( .A(n53749), .Z(n53750) );
  NAND U63388 ( .A(n53751), .B(n53752), .Z(n53726) );
  NAND U63389 ( .A(n53753), .B(n53754), .Z(n53752) );
  NANDN U63390 ( .A(n53755), .B(n53756), .Z(n53753) );
  NANDN U63391 ( .A(n53756), .B(n53755), .Z(n53751) );
  AND U63392 ( .A(n53757), .B(n53758), .Z(n53728) );
  NAND U63393 ( .A(n53759), .B(n53760), .Z(n53758) );
  OR U63394 ( .A(n53761), .B(n53762), .Z(n53759) );
  NANDN U63395 ( .A(n53763), .B(n53761), .Z(n53757) );
  NAND U63396 ( .A(n53764), .B(n53765), .Z(n53732) );
  NANDN U63397 ( .A(n53766), .B(n53767), .Z(n53765) );
  OR U63398 ( .A(n53768), .B(n53769), .Z(n53767) );
  NANDN U63399 ( .A(n53770), .B(n53768), .Z(n53764) );
  IV U63400 ( .A(n53769), .Z(n53770) );
  XNOR U63401 ( .A(n53740), .B(n53771), .Z(n53735) );
  XNOR U63402 ( .A(n53738), .B(n53741), .Z(n53771) );
  NAND U63403 ( .A(n53772), .B(n53773), .Z(n53741) );
  NAND U63404 ( .A(n53774), .B(n53775), .Z(n53773) );
  OR U63405 ( .A(n53776), .B(n53777), .Z(n53774) );
  NANDN U63406 ( .A(n53778), .B(n53776), .Z(n53772) );
  IV U63407 ( .A(n53777), .Z(n53778) );
  NAND U63408 ( .A(n53779), .B(n53780), .Z(n53738) );
  NAND U63409 ( .A(n53781), .B(n53782), .Z(n53780) );
  NANDN U63410 ( .A(n53783), .B(n53784), .Z(n53781) );
  NANDN U63411 ( .A(n53784), .B(n53783), .Z(n53779) );
  AND U63412 ( .A(n53785), .B(n53786), .Z(n53740) );
  NAND U63413 ( .A(n53787), .B(n53788), .Z(n53786) );
  OR U63414 ( .A(n53789), .B(n53790), .Z(n53787) );
  NANDN U63415 ( .A(n53791), .B(n53789), .Z(n53785) );
  XNOR U63416 ( .A(n53766), .B(n53792), .Z(N60632) );
  XOR U63417 ( .A(n53768), .B(n53769), .Z(n53792) );
  XNOR U63418 ( .A(n53782), .B(n53793), .Z(n53769) );
  XOR U63419 ( .A(n53783), .B(n53784), .Z(n53793) );
  XOR U63420 ( .A(n53789), .B(n53794), .Z(n53784) );
  XOR U63421 ( .A(n53788), .B(n53791), .Z(n53794) );
  IV U63422 ( .A(n53790), .Z(n53791) );
  NAND U63423 ( .A(n53795), .B(n53796), .Z(n53790) );
  OR U63424 ( .A(n53797), .B(n53798), .Z(n53796) );
  OR U63425 ( .A(n53799), .B(n53800), .Z(n53795) );
  NAND U63426 ( .A(n53801), .B(n53802), .Z(n53788) );
  OR U63427 ( .A(n53803), .B(n53804), .Z(n53802) );
  OR U63428 ( .A(n53805), .B(n53806), .Z(n53801) );
  NOR U63429 ( .A(n53807), .B(n53808), .Z(n53789) );
  ANDN U63430 ( .B(n53809), .A(n53810), .Z(n53783) );
  XNOR U63431 ( .A(n53776), .B(n53811), .Z(n53782) );
  XNOR U63432 ( .A(n53775), .B(n53777), .Z(n53811) );
  NAND U63433 ( .A(n53812), .B(n53813), .Z(n53777) );
  OR U63434 ( .A(n53814), .B(n53815), .Z(n53813) );
  OR U63435 ( .A(n53816), .B(n53817), .Z(n53812) );
  NAND U63436 ( .A(n53818), .B(n53819), .Z(n53775) );
  OR U63437 ( .A(n53820), .B(n53821), .Z(n53819) );
  OR U63438 ( .A(n53822), .B(n53823), .Z(n53818) );
  ANDN U63439 ( .B(n53824), .A(n53825), .Z(n53776) );
  IV U63440 ( .A(n53826), .Z(n53824) );
  ANDN U63441 ( .B(n53827), .A(n53828), .Z(n53768) );
  XOR U63442 ( .A(n53754), .B(n53829), .Z(n53766) );
  XOR U63443 ( .A(n53755), .B(n53756), .Z(n53829) );
  XOR U63444 ( .A(n53761), .B(n53830), .Z(n53756) );
  XOR U63445 ( .A(n53760), .B(n53763), .Z(n53830) );
  IV U63446 ( .A(n53762), .Z(n53763) );
  NAND U63447 ( .A(n53831), .B(n53832), .Z(n53762) );
  OR U63448 ( .A(n53833), .B(n53834), .Z(n53832) );
  OR U63449 ( .A(n53835), .B(n53836), .Z(n53831) );
  NAND U63450 ( .A(n53837), .B(n53838), .Z(n53760) );
  OR U63451 ( .A(n53839), .B(n53840), .Z(n53838) );
  OR U63452 ( .A(n53841), .B(n53842), .Z(n53837) );
  NOR U63453 ( .A(n53843), .B(n53844), .Z(n53761) );
  ANDN U63454 ( .B(n53845), .A(n53846), .Z(n53755) );
  IV U63455 ( .A(n53847), .Z(n53845) );
  XNOR U63456 ( .A(n53748), .B(n53848), .Z(n53754) );
  XNOR U63457 ( .A(n53747), .B(n53749), .Z(n53848) );
  NAND U63458 ( .A(n53849), .B(n53850), .Z(n53749) );
  OR U63459 ( .A(n53851), .B(n53852), .Z(n53850) );
  OR U63460 ( .A(n53853), .B(n53854), .Z(n53849) );
  NAND U63461 ( .A(n53855), .B(n53856), .Z(n53747) );
  OR U63462 ( .A(n53857), .B(n53858), .Z(n53856) );
  OR U63463 ( .A(n53859), .B(n53860), .Z(n53855) );
  ANDN U63464 ( .B(n53861), .A(n53862), .Z(n53748) );
  IV U63465 ( .A(n53863), .Z(n53861) );
  XNOR U63466 ( .A(n53828), .B(n53827), .Z(N60631) );
  XOR U63467 ( .A(n53847), .B(n53846), .Z(n53827) );
  XNOR U63468 ( .A(n53862), .B(n53863), .Z(n53846) );
  XNOR U63469 ( .A(n53857), .B(n53858), .Z(n53863) );
  XNOR U63470 ( .A(n53859), .B(n53860), .Z(n53858) );
  XNOR U63471 ( .A(y[85]), .B(x[85]), .Z(n53860) );
  XNOR U63472 ( .A(y[86]), .B(x[86]), .Z(n53859) );
  XNOR U63473 ( .A(y[84]), .B(x[84]), .Z(n53857) );
  XNOR U63474 ( .A(n53851), .B(n53852), .Z(n53862) );
  XNOR U63475 ( .A(y[81]), .B(x[81]), .Z(n53852) );
  XNOR U63476 ( .A(n53853), .B(n53854), .Z(n53851) );
  XNOR U63477 ( .A(y[82]), .B(x[82]), .Z(n53854) );
  XNOR U63478 ( .A(y[83]), .B(x[83]), .Z(n53853) );
  XNOR U63479 ( .A(n53844), .B(n53843), .Z(n53847) );
  XNOR U63480 ( .A(n53839), .B(n53840), .Z(n53843) );
  XNOR U63481 ( .A(y[78]), .B(x[78]), .Z(n53840) );
  XNOR U63482 ( .A(n53841), .B(n53842), .Z(n53839) );
  XNOR U63483 ( .A(y[79]), .B(x[79]), .Z(n53842) );
  XNOR U63484 ( .A(y[80]), .B(x[80]), .Z(n53841) );
  XNOR U63485 ( .A(n53833), .B(n53834), .Z(n53844) );
  XNOR U63486 ( .A(y[75]), .B(x[75]), .Z(n53834) );
  XNOR U63487 ( .A(n53835), .B(n53836), .Z(n53833) );
  XNOR U63488 ( .A(y[76]), .B(x[76]), .Z(n53836) );
  XNOR U63489 ( .A(y[77]), .B(x[77]), .Z(n53835) );
  XOR U63490 ( .A(n53809), .B(n53810), .Z(n53828) );
  XNOR U63491 ( .A(n53825), .B(n53826), .Z(n53810) );
  XNOR U63492 ( .A(n53820), .B(n53821), .Z(n53826) );
  XNOR U63493 ( .A(n53822), .B(n53823), .Z(n53821) );
  XNOR U63494 ( .A(y[73]), .B(x[73]), .Z(n53823) );
  XNOR U63495 ( .A(y[74]), .B(x[74]), .Z(n53822) );
  XNOR U63496 ( .A(y[72]), .B(x[72]), .Z(n53820) );
  XNOR U63497 ( .A(n53814), .B(n53815), .Z(n53825) );
  XNOR U63498 ( .A(y[69]), .B(x[69]), .Z(n53815) );
  XNOR U63499 ( .A(n53816), .B(n53817), .Z(n53814) );
  XNOR U63500 ( .A(y[70]), .B(x[70]), .Z(n53817) );
  XNOR U63501 ( .A(y[71]), .B(x[71]), .Z(n53816) );
  XOR U63502 ( .A(n53808), .B(n53807), .Z(n53809) );
  XNOR U63503 ( .A(n53803), .B(n53804), .Z(n53807) );
  XNOR U63504 ( .A(y[66]), .B(x[66]), .Z(n53804) );
  XNOR U63505 ( .A(n53805), .B(n53806), .Z(n53803) );
  XNOR U63506 ( .A(y[67]), .B(x[67]), .Z(n53806) );
  XNOR U63507 ( .A(y[68]), .B(x[68]), .Z(n53805) );
  XNOR U63508 ( .A(n53797), .B(n53798), .Z(n53808) );
  XNOR U63509 ( .A(y[63]), .B(x[63]), .Z(n53798) );
  XNOR U63510 ( .A(n53799), .B(n53800), .Z(n53797) );
  XNOR U63511 ( .A(y[64]), .B(x[64]), .Z(n53800) );
  XNOR U63512 ( .A(y[65]), .B(x[65]), .Z(n53799) );
  NAND U63513 ( .A(n53864), .B(n53865), .Z(N60622) );
  NANDN U63514 ( .A(n53866), .B(n53867), .Z(n53865) );
  OR U63515 ( .A(n53868), .B(n53869), .Z(n53867) );
  NAND U63516 ( .A(n53868), .B(n53869), .Z(n53864) );
  XOR U63517 ( .A(n53868), .B(n53870), .Z(N60621) );
  XNOR U63518 ( .A(n53866), .B(n53869), .Z(n53870) );
  AND U63519 ( .A(n53871), .B(n53872), .Z(n53869) );
  NANDN U63520 ( .A(n53873), .B(n53874), .Z(n53872) );
  NANDN U63521 ( .A(n53875), .B(n53876), .Z(n53874) );
  NANDN U63522 ( .A(n53876), .B(n53875), .Z(n53871) );
  NAND U63523 ( .A(n53877), .B(n53878), .Z(n53866) );
  NANDN U63524 ( .A(n53879), .B(n53880), .Z(n53878) );
  OR U63525 ( .A(n53881), .B(n53882), .Z(n53880) );
  NAND U63526 ( .A(n53882), .B(n53881), .Z(n53877) );
  AND U63527 ( .A(n53883), .B(n53884), .Z(n53868) );
  NANDN U63528 ( .A(n53885), .B(n53886), .Z(n53884) );
  NANDN U63529 ( .A(n53887), .B(n53888), .Z(n53886) );
  NANDN U63530 ( .A(n53888), .B(n53887), .Z(n53883) );
  XOR U63531 ( .A(n53882), .B(n53889), .Z(N60620) );
  XOR U63532 ( .A(n53879), .B(n53881), .Z(n53889) );
  XNOR U63533 ( .A(n53875), .B(n53890), .Z(n53881) );
  XNOR U63534 ( .A(n53873), .B(n53876), .Z(n53890) );
  NAND U63535 ( .A(n53891), .B(n53892), .Z(n53876) );
  NAND U63536 ( .A(n53893), .B(n53894), .Z(n53892) );
  OR U63537 ( .A(n53895), .B(n53896), .Z(n53893) );
  NANDN U63538 ( .A(n53897), .B(n53895), .Z(n53891) );
  IV U63539 ( .A(n53896), .Z(n53897) );
  NAND U63540 ( .A(n53898), .B(n53899), .Z(n53873) );
  NAND U63541 ( .A(n53900), .B(n53901), .Z(n53899) );
  NANDN U63542 ( .A(n53902), .B(n53903), .Z(n53900) );
  NANDN U63543 ( .A(n53903), .B(n53902), .Z(n53898) );
  AND U63544 ( .A(n53904), .B(n53905), .Z(n53875) );
  NAND U63545 ( .A(n53906), .B(n53907), .Z(n53905) );
  OR U63546 ( .A(n53908), .B(n53909), .Z(n53906) );
  NANDN U63547 ( .A(n53910), .B(n53908), .Z(n53904) );
  NAND U63548 ( .A(n53911), .B(n53912), .Z(n53879) );
  NANDN U63549 ( .A(n53913), .B(n53914), .Z(n53912) );
  OR U63550 ( .A(n53915), .B(n53916), .Z(n53914) );
  NANDN U63551 ( .A(n53917), .B(n53915), .Z(n53911) );
  IV U63552 ( .A(n53916), .Z(n53917) );
  XNOR U63553 ( .A(n53887), .B(n53918), .Z(n53882) );
  XNOR U63554 ( .A(n53885), .B(n53888), .Z(n53918) );
  NAND U63555 ( .A(n53919), .B(n53920), .Z(n53888) );
  NAND U63556 ( .A(n53921), .B(n53922), .Z(n53920) );
  OR U63557 ( .A(n53923), .B(n53924), .Z(n53921) );
  NANDN U63558 ( .A(n53925), .B(n53923), .Z(n53919) );
  IV U63559 ( .A(n53924), .Z(n53925) );
  NAND U63560 ( .A(n53926), .B(n53927), .Z(n53885) );
  NAND U63561 ( .A(n53928), .B(n53929), .Z(n53927) );
  NANDN U63562 ( .A(n53930), .B(n53931), .Z(n53928) );
  NANDN U63563 ( .A(n53931), .B(n53930), .Z(n53926) );
  AND U63564 ( .A(n53932), .B(n53933), .Z(n53887) );
  NAND U63565 ( .A(n53934), .B(n53935), .Z(n53933) );
  OR U63566 ( .A(n53936), .B(n53937), .Z(n53934) );
  NANDN U63567 ( .A(n53938), .B(n53936), .Z(n53932) );
  XNOR U63568 ( .A(n53913), .B(n53939), .Z(N60619) );
  XOR U63569 ( .A(n53915), .B(n53916), .Z(n53939) );
  XNOR U63570 ( .A(n53929), .B(n53940), .Z(n53916) );
  XOR U63571 ( .A(n53930), .B(n53931), .Z(n53940) );
  XOR U63572 ( .A(n53936), .B(n53941), .Z(n53931) );
  XOR U63573 ( .A(n53935), .B(n53938), .Z(n53941) );
  IV U63574 ( .A(n53937), .Z(n53938) );
  NAND U63575 ( .A(n53942), .B(n53943), .Z(n53937) );
  OR U63576 ( .A(n53944), .B(n53945), .Z(n53943) );
  OR U63577 ( .A(n53946), .B(n53947), .Z(n53942) );
  NAND U63578 ( .A(n53948), .B(n53949), .Z(n53935) );
  OR U63579 ( .A(n53950), .B(n53951), .Z(n53949) );
  OR U63580 ( .A(n53952), .B(n53953), .Z(n53948) );
  NOR U63581 ( .A(n53954), .B(n53955), .Z(n53936) );
  ANDN U63582 ( .B(n53956), .A(n53957), .Z(n53930) );
  XNOR U63583 ( .A(n53923), .B(n53958), .Z(n53929) );
  XNOR U63584 ( .A(n53922), .B(n53924), .Z(n53958) );
  NAND U63585 ( .A(n53959), .B(n53960), .Z(n53924) );
  OR U63586 ( .A(n53961), .B(n53962), .Z(n53960) );
  OR U63587 ( .A(n53963), .B(n53964), .Z(n53959) );
  NAND U63588 ( .A(n53965), .B(n53966), .Z(n53922) );
  OR U63589 ( .A(n53967), .B(n53968), .Z(n53966) );
  OR U63590 ( .A(n53969), .B(n53970), .Z(n53965) );
  ANDN U63591 ( .B(n53971), .A(n53972), .Z(n53923) );
  IV U63592 ( .A(n53973), .Z(n53971) );
  ANDN U63593 ( .B(n53974), .A(n53975), .Z(n53915) );
  XOR U63594 ( .A(n53901), .B(n53976), .Z(n53913) );
  XOR U63595 ( .A(n53902), .B(n53903), .Z(n53976) );
  XOR U63596 ( .A(n53908), .B(n53977), .Z(n53903) );
  XOR U63597 ( .A(n53907), .B(n53910), .Z(n53977) );
  IV U63598 ( .A(n53909), .Z(n53910) );
  NAND U63599 ( .A(n53978), .B(n53979), .Z(n53909) );
  OR U63600 ( .A(n53980), .B(n53981), .Z(n53979) );
  OR U63601 ( .A(n53982), .B(n53983), .Z(n53978) );
  NAND U63602 ( .A(n53984), .B(n53985), .Z(n53907) );
  OR U63603 ( .A(n53986), .B(n53987), .Z(n53985) );
  OR U63604 ( .A(n53988), .B(n53989), .Z(n53984) );
  NOR U63605 ( .A(n53990), .B(n53991), .Z(n53908) );
  ANDN U63606 ( .B(n53992), .A(n53993), .Z(n53902) );
  IV U63607 ( .A(n53994), .Z(n53992) );
  XNOR U63608 ( .A(n53895), .B(n53995), .Z(n53901) );
  XNOR U63609 ( .A(n53894), .B(n53896), .Z(n53995) );
  NAND U63610 ( .A(n53996), .B(n53997), .Z(n53896) );
  OR U63611 ( .A(n53998), .B(n53999), .Z(n53997) );
  OR U63612 ( .A(n54000), .B(n54001), .Z(n53996) );
  NAND U63613 ( .A(n54002), .B(n54003), .Z(n53894) );
  OR U63614 ( .A(n54004), .B(n54005), .Z(n54003) );
  OR U63615 ( .A(n54006), .B(n54007), .Z(n54002) );
  ANDN U63616 ( .B(n54008), .A(n54009), .Z(n53895) );
  IV U63617 ( .A(n54010), .Z(n54008) );
  XNOR U63618 ( .A(n53975), .B(n53974), .Z(N60618) );
  XOR U63619 ( .A(n53994), .B(n53993), .Z(n53974) );
  XNOR U63620 ( .A(n54009), .B(n54010), .Z(n53993) );
  XNOR U63621 ( .A(n54004), .B(n54005), .Z(n54010) );
  XNOR U63622 ( .A(n54006), .B(n54007), .Z(n54005) );
  XNOR U63623 ( .A(y[61]), .B(x[61]), .Z(n54007) );
  XNOR U63624 ( .A(y[62]), .B(x[62]), .Z(n54006) );
  XNOR U63625 ( .A(y[60]), .B(x[60]), .Z(n54004) );
  XNOR U63626 ( .A(n53998), .B(n53999), .Z(n54009) );
  XNOR U63627 ( .A(y[57]), .B(x[57]), .Z(n53999) );
  XNOR U63628 ( .A(n54000), .B(n54001), .Z(n53998) );
  XNOR U63629 ( .A(y[58]), .B(x[58]), .Z(n54001) );
  XNOR U63630 ( .A(y[59]), .B(x[59]), .Z(n54000) );
  XNOR U63631 ( .A(n53991), .B(n53990), .Z(n53994) );
  XNOR U63632 ( .A(n53986), .B(n53987), .Z(n53990) );
  XNOR U63633 ( .A(y[54]), .B(x[54]), .Z(n53987) );
  XNOR U63634 ( .A(n53988), .B(n53989), .Z(n53986) );
  XNOR U63635 ( .A(y[55]), .B(x[55]), .Z(n53989) );
  XNOR U63636 ( .A(y[56]), .B(x[56]), .Z(n53988) );
  XNOR U63637 ( .A(n53980), .B(n53981), .Z(n53991) );
  XNOR U63638 ( .A(y[51]), .B(x[51]), .Z(n53981) );
  XNOR U63639 ( .A(n53982), .B(n53983), .Z(n53980) );
  XNOR U63640 ( .A(y[52]), .B(x[52]), .Z(n53983) );
  XNOR U63641 ( .A(y[53]), .B(x[53]), .Z(n53982) );
  XOR U63642 ( .A(n53956), .B(n53957), .Z(n53975) );
  XNOR U63643 ( .A(n53972), .B(n53973), .Z(n53957) );
  XNOR U63644 ( .A(n53967), .B(n53968), .Z(n53973) );
  XNOR U63645 ( .A(n53969), .B(n53970), .Z(n53968) );
  XNOR U63646 ( .A(y[49]), .B(x[49]), .Z(n53970) );
  XNOR U63647 ( .A(y[50]), .B(x[50]), .Z(n53969) );
  XNOR U63648 ( .A(y[48]), .B(x[48]), .Z(n53967) );
  XNOR U63649 ( .A(n53961), .B(n53962), .Z(n53972) );
  XNOR U63650 ( .A(y[45]), .B(x[45]), .Z(n53962) );
  XNOR U63651 ( .A(n53963), .B(n53964), .Z(n53961) );
  XNOR U63652 ( .A(y[46]), .B(x[46]), .Z(n53964) );
  XNOR U63653 ( .A(y[47]), .B(x[47]), .Z(n53963) );
  XOR U63654 ( .A(n53955), .B(n53954), .Z(n53956) );
  XNOR U63655 ( .A(n53950), .B(n53951), .Z(n53954) );
  XNOR U63656 ( .A(y[42]), .B(x[42]), .Z(n53951) );
  XNOR U63657 ( .A(n53952), .B(n53953), .Z(n53950) );
  XNOR U63658 ( .A(y[43]), .B(x[43]), .Z(n53953) );
  XNOR U63659 ( .A(y[44]), .B(x[44]), .Z(n53952) );
  XNOR U63660 ( .A(n53944), .B(n53945), .Z(n53955) );
  XNOR U63661 ( .A(y[39]), .B(x[39]), .Z(n53945) );
  XNOR U63662 ( .A(n53946), .B(n53947), .Z(n53944) );
  XNOR U63663 ( .A(y[40]), .B(x[40]), .Z(n53947) );
  XNOR U63664 ( .A(y[41]), .B(x[41]), .Z(n53946) );
  NAND U63665 ( .A(n54011), .B(n54012), .Z(N60609) );
  NANDN U63666 ( .A(n54013), .B(n54014), .Z(n54012) );
  OR U63667 ( .A(n54015), .B(n54016), .Z(n54014) );
  NAND U63668 ( .A(n54015), .B(n54016), .Z(n54011) );
  XOR U63669 ( .A(n54015), .B(n54017), .Z(N60608) );
  XNOR U63670 ( .A(n54013), .B(n54016), .Z(n54017) );
  AND U63671 ( .A(n54018), .B(n54019), .Z(n54016) );
  NANDN U63672 ( .A(n54020), .B(n54021), .Z(n54019) );
  NANDN U63673 ( .A(n54022), .B(n54023), .Z(n54021) );
  NANDN U63674 ( .A(n54023), .B(n54022), .Z(n54018) );
  NAND U63675 ( .A(n54024), .B(n54025), .Z(n54013) );
  NANDN U63676 ( .A(n54026), .B(n54027), .Z(n54025) );
  OR U63677 ( .A(n54028), .B(n54029), .Z(n54027) );
  NAND U63678 ( .A(n54029), .B(n54028), .Z(n54024) );
  AND U63679 ( .A(n54030), .B(n54031), .Z(n54015) );
  NANDN U63680 ( .A(n54032), .B(n54033), .Z(n54031) );
  NANDN U63681 ( .A(n54034), .B(n54035), .Z(n54033) );
  NANDN U63682 ( .A(n54035), .B(n54034), .Z(n54030) );
  XOR U63683 ( .A(n54029), .B(n54036), .Z(N60607) );
  XOR U63684 ( .A(n54026), .B(n54028), .Z(n54036) );
  XNOR U63685 ( .A(n54022), .B(n54037), .Z(n54028) );
  XNOR U63686 ( .A(n54020), .B(n54023), .Z(n54037) );
  NAND U63687 ( .A(n54038), .B(n54039), .Z(n54023) );
  NAND U63688 ( .A(n54040), .B(n54041), .Z(n54039) );
  OR U63689 ( .A(n54042), .B(n54043), .Z(n54040) );
  NANDN U63690 ( .A(n54044), .B(n54042), .Z(n54038) );
  IV U63691 ( .A(n54043), .Z(n54044) );
  NAND U63692 ( .A(n54045), .B(n54046), .Z(n54020) );
  NAND U63693 ( .A(n54047), .B(n54048), .Z(n54046) );
  NANDN U63694 ( .A(n54049), .B(n54050), .Z(n54047) );
  NANDN U63695 ( .A(n54050), .B(n54049), .Z(n54045) );
  AND U63696 ( .A(n54051), .B(n54052), .Z(n54022) );
  NAND U63697 ( .A(n54053), .B(n54054), .Z(n54052) );
  OR U63698 ( .A(n54055), .B(n54056), .Z(n54053) );
  NANDN U63699 ( .A(n54057), .B(n54055), .Z(n54051) );
  NAND U63700 ( .A(n54058), .B(n54059), .Z(n54026) );
  NANDN U63701 ( .A(n54060), .B(n54061), .Z(n54059) );
  OR U63702 ( .A(n54062), .B(n54063), .Z(n54061) );
  NANDN U63703 ( .A(n54064), .B(n54062), .Z(n54058) );
  IV U63704 ( .A(n54063), .Z(n54064) );
  XNOR U63705 ( .A(n54034), .B(n54065), .Z(n54029) );
  XNOR U63706 ( .A(n54032), .B(n54035), .Z(n54065) );
  NAND U63707 ( .A(n54066), .B(n54067), .Z(n54035) );
  NAND U63708 ( .A(n54068), .B(n54069), .Z(n54067) );
  OR U63709 ( .A(n54070), .B(n54071), .Z(n54068) );
  NANDN U63710 ( .A(n54072), .B(n54070), .Z(n54066) );
  IV U63711 ( .A(n54071), .Z(n54072) );
  NAND U63712 ( .A(n54073), .B(n54074), .Z(n54032) );
  NAND U63713 ( .A(n54075), .B(n54076), .Z(n54074) );
  NANDN U63714 ( .A(n54077), .B(n54078), .Z(n54075) );
  NANDN U63715 ( .A(n54078), .B(n54077), .Z(n54073) );
  AND U63716 ( .A(n54079), .B(n54080), .Z(n54034) );
  NAND U63717 ( .A(n54081), .B(n54082), .Z(n54080) );
  OR U63718 ( .A(n54083), .B(n54084), .Z(n54081) );
  NANDN U63719 ( .A(n54085), .B(n54083), .Z(n54079) );
  XNOR U63720 ( .A(n54060), .B(n54086), .Z(N60606) );
  XOR U63721 ( .A(n54062), .B(n54063), .Z(n54086) );
  XNOR U63722 ( .A(n54076), .B(n54087), .Z(n54063) );
  XOR U63723 ( .A(n54077), .B(n54078), .Z(n54087) );
  XOR U63724 ( .A(n54083), .B(n54088), .Z(n54078) );
  XOR U63725 ( .A(n54082), .B(n54085), .Z(n54088) );
  IV U63726 ( .A(n54084), .Z(n54085) );
  NAND U63727 ( .A(n54089), .B(n54090), .Z(n54084) );
  OR U63728 ( .A(n54091), .B(n54092), .Z(n54090) );
  OR U63729 ( .A(n54093), .B(n54094), .Z(n54089) );
  NAND U63730 ( .A(n54095), .B(n54096), .Z(n54082) );
  OR U63731 ( .A(n54097), .B(n54098), .Z(n54096) );
  OR U63732 ( .A(n54099), .B(n54100), .Z(n54095) );
  NOR U63733 ( .A(n54101), .B(n54102), .Z(n54083) );
  ANDN U63734 ( .B(n54103), .A(n54104), .Z(n54077) );
  XNOR U63735 ( .A(n54070), .B(n54105), .Z(n54076) );
  XNOR U63736 ( .A(n54069), .B(n54071), .Z(n54105) );
  NAND U63737 ( .A(n54106), .B(n54107), .Z(n54071) );
  OR U63738 ( .A(n54108), .B(n54109), .Z(n54107) );
  OR U63739 ( .A(n54110), .B(n54111), .Z(n54106) );
  NAND U63740 ( .A(n54112), .B(n54113), .Z(n54069) );
  OR U63741 ( .A(n54114), .B(n54115), .Z(n54113) );
  OR U63742 ( .A(n54116), .B(n54117), .Z(n54112) );
  ANDN U63743 ( .B(n54118), .A(n54119), .Z(n54070) );
  IV U63744 ( .A(n54120), .Z(n54118) );
  ANDN U63745 ( .B(n54121), .A(n54122), .Z(n54062) );
  XOR U63746 ( .A(n54048), .B(n54123), .Z(n54060) );
  XOR U63747 ( .A(n54049), .B(n54050), .Z(n54123) );
  XOR U63748 ( .A(n54055), .B(n54124), .Z(n54050) );
  XOR U63749 ( .A(n54054), .B(n54057), .Z(n54124) );
  IV U63750 ( .A(n54056), .Z(n54057) );
  NAND U63751 ( .A(n54125), .B(n54126), .Z(n54056) );
  OR U63752 ( .A(n54127), .B(n54128), .Z(n54126) );
  OR U63753 ( .A(n54129), .B(n54130), .Z(n54125) );
  NAND U63754 ( .A(n54131), .B(n54132), .Z(n54054) );
  OR U63755 ( .A(n54133), .B(n54134), .Z(n54132) );
  OR U63756 ( .A(n54135), .B(n54136), .Z(n54131) );
  NOR U63757 ( .A(n54137), .B(n54138), .Z(n54055) );
  ANDN U63758 ( .B(n54139), .A(n54140), .Z(n54049) );
  IV U63759 ( .A(n54141), .Z(n54139) );
  XNOR U63760 ( .A(n54042), .B(n54142), .Z(n54048) );
  XNOR U63761 ( .A(n54041), .B(n54043), .Z(n54142) );
  NAND U63762 ( .A(n54143), .B(n54144), .Z(n54043) );
  OR U63763 ( .A(n54145), .B(n54146), .Z(n54144) );
  OR U63764 ( .A(n54147), .B(n54148), .Z(n54143) );
  NAND U63765 ( .A(n54149), .B(n54150), .Z(n54041) );
  OR U63766 ( .A(n54151), .B(n54152), .Z(n54150) );
  OR U63767 ( .A(n54153), .B(n54154), .Z(n54149) );
  ANDN U63768 ( .B(n54155), .A(n54156), .Z(n54042) );
  IV U63769 ( .A(n54157), .Z(n54155) );
  XNOR U63770 ( .A(n54122), .B(n54121), .Z(N60605) );
  XOR U63771 ( .A(n54141), .B(n54140), .Z(n54121) );
  XNOR U63772 ( .A(n54156), .B(n54157), .Z(n54140) );
  XNOR U63773 ( .A(n54151), .B(n54152), .Z(n54157) );
  XNOR U63774 ( .A(n54153), .B(n54154), .Z(n54152) );
  XNOR U63775 ( .A(y[37]), .B(x[37]), .Z(n54154) );
  XNOR U63776 ( .A(y[38]), .B(x[38]), .Z(n54153) );
  XNOR U63777 ( .A(y[36]), .B(x[36]), .Z(n54151) );
  XNOR U63778 ( .A(n54145), .B(n54146), .Z(n54156) );
  XNOR U63779 ( .A(y[33]), .B(x[33]), .Z(n54146) );
  XNOR U63780 ( .A(n54147), .B(n54148), .Z(n54145) );
  XNOR U63781 ( .A(y[34]), .B(x[34]), .Z(n54148) );
  XNOR U63782 ( .A(y[35]), .B(x[35]), .Z(n54147) );
  XNOR U63783 ( .A(n54138), .B(n54137), .Z(n54141) );
  XNOR U63784 ( .A(n54133), .B(n54134), .Z(n54137) );
  XNOR U63785 ( .A(y[30]), .B(x[30]), .Z(n54134) );
  XNOR U63786 ( .A(n54135), .B(n54136), .Z(n54133) );
  XNOR U63787 ( .A(y[31]), .B(x[31]), .Z(n54136) );
  XNOR U63788 ( .A(y[32]), .B(x[32]), .Z(n54135) );
  XNOR U63789 ( .A(n54127), .B(n54128), .Z(n54138) );
  XNOR U63790 ( .A(y[27]), .B(x[27]), .Z(n54128) );
  XNOR U63791 ( .A(n54129), .B(n54130), .Z(n54127) );
  XNOR U63792 ( .A(y[28]), .B(x[28]), .Z(n54130) );
  XNOR U63793 ( .A(y[29]), .B(x[29]), .Z(n54129) );
  XOR U63794 ( .A(n54103), .B(n54104), .Z(n54122) );
  XNOR U63795 ( .A(n54119), .B(n54120), .Z(n54104) );
  XNOR U63796 ( .A(n54114), .B(n54115), .Z(n54120) );
  XNOR U63797 ( .A(n54116), .B(n54117), .Z(n54115) );
  XNOR U63798 ( .A(y[25]), .B(x[25]), .Z(n54117) );
  XNOR U63799 ( .A(y[26]), .B(x[26]), .Z(n54116) );
  XNOR U63800 ( .A(y[24]), .B(x[24]), .Z(n54114) );
  XNOR U63801 ( .A(n54108), .B(n54109), .Z(n54119) );
  XNOR U63802 ( .A(y[21]), .B(x[21]), .Z(n54109) );
  XNOR U63803 ( .A(n54110), .B(n54111), .Z(n54108) );
  XNOR U63804 ( .A(y[22]), .B(x[22]), .Z(n54111) );
  XNOR U63805 ( .A(y[23]), .B(x[23]), .Z(n54110) );
  XOR U63806 ( .A(n54102), .B(n54101), .Z(n54103) );
  XNOR U63807 ( .A(n54097), .B(n54098), .Z(n54101) );
  XNOR U63808 ( .A(y[18]), .B(x[18]), .Z(n54098) );
  XNOR U63809 ( .A(n54099), .B(n54100), .Z(n54097) );
  XNOR U63810 ( .A(y[19]), .B(x[19]), .Z(n54100) );
  XNOR U63811 ( .A(y[20]), .B(x[20]), .Z(n54099) );
  XNOR U63812 ( .A(n54091), .B(n54092), .Z(n54102) );
  XNOR U63813 ( .A(y[15]), .B(x[15]), .Z(n54092) );
  XNOR U63814 ( .A(n54093), .B(n54094), .Z(n54091) );
  XNOR U63815 ( .A(y[16]), .B(x[16]), .Z(n54094) );
  XNOR U63816 ( .A(y[17]), .B(x[17]), .Z(n54093) );
  NAND U63817 ( .A(n54158), .B(n54159), .Z(N60596) );
  OR U63818 ( .A(n54160), .B(n54161), .Z(n54159) );
  OR U63819 ( .A(n54161), .B(n54162), .Z(n54158) );
  XNOR U63820 ( .A(n54162), .B(n54163), .Z(N60595) );
  XOR U63821 ( .A(n54160), .B(n54161), .Z(n54163) );
  NAND U63822 ( .A(n54164), .B(n54165), .Z(n54161) );
  NANDN U63823 ( .A(n54166), .B(n54167), .Z(n54165) );
  NANDN U63824 ( .A(n54168), .B(n54169), .Z(n54167) );
  NANDN U63825 ( .A(n54169), .B(n54168), .Z(n54164) );
  NAND U63826 ( .A(n54170), .B(n54171), .Z(n54160) );
  NANDN U63827 ( .A(n54172), .B(n54173), .Z(n54171) );
  OR U63828 ( .A(n54174), .B(n54175), .Z(n54173) );
  NANDN U63829 ( .A(n54176), .B(n54174), .Z(n54170) );
  IV U63830 ( .A(n54175), .Z(n54176) );
  NANDN U63831 ( .A(n54177), .B(n54178), .Z(n54162) );
  XOR U63832 ( .A(n54175), .B(n54179), .Z(N60594) );
  XOR U63833 ( .A(n54172), .B(n54174), .Z(n54179) );
  XNOR U63834 ( .A(n54168), .B(n54180), .Z(n54174) );
  XNOR U63835 ( .A(n54166), .B(n54169), .Z(n54180) );
  NAND U63836 ( .A(n54181), .B(n54182), .Z(n54169) );
  NAND U63837 ( .A(n54183), .B(n54184), .Z(n54182) );
  OR U63838 ( .A(n54185), .B(n54186), .Z(n54183) );
  NANDN U63839 ( .A(n54187), .B(n54185), .Z(n54181) );
  IV U63840 ( .A(n54186), .Z(n54187) );
  NAND U63841 ( .A(n54188), .B(n54189), .Z(n54166) );
  NAND U63842 ( .A(n54190), .B(n54191), .Z(n54189) );
  NANDN U63843 ( .A(n54192), .B(n54193), .Z(n54190) );
  NANDN U63844 ( .A(n54193), .B(n54192), .Z(n54188) );
  AND U63845 ( .A(n54194), .B(n54195), .Z(n54168) );
  NAND U63846 ( .A(n54196), .B(n54197), .Z(n54195) );
  NANDN U63847 ( .A(n54198), .B(n54199), .Z(n54194) );
  NAND U63848 ( .A(n54200), .B(n54201), .Z(n54172) );
  NANDN U63849 ( .A(n54202), .B(n54203), .Z(n54201) );
  OR U63850 ( .A(n54204), .B(n54205), .Z(n54203) );
  NAND U63851 ( .A(n54205), .B(n54204), .Z(n54200) );
  XOR U63852 ( .A(n54178), .B(n54177), .Z(n54175) );
  NANDN U63853 ( .A(n54206), .B(n54207), .Z(n54177) );
  NAND U63854 ( .A(n54208), .B(n54209), .Z(n54178) );
  NAND U63855 ( .A(n54210), .B(n54211), .Z(n54209) );
  NAND U63856 ( .A(n54212), .B(n54213), .Z(n54210) );
  OR U63857 ( .A(n54212), .B(n54213), .Z(n54208) );
  XNOR U63858 ( .A(n54202), .B(n54214), .Z(N60593) );
  XOR U63859 ( .A(n54204), .B(n54205), .Z(n54214) );
  XOR U63860 ( .A(n54211), .B(n54215), .Z(n54205) );
  XOR U63861 ( .A(n54213), .B(n54212), .Z(n54215) );
  NANDN U63862 ( .A(n54216), .B(n54217), .Z(n54212) );
  AND U63863 ( .A(n54218), .B(n54219), .Z(n54213) );
  OR U63864 ( .A(n54220), .B(n54221), .Z(n54219) );
  OR U63865 ( .A(n54222), .B(n54223), .Z(n54218) );
  XNOR U63866 ( .A(n54207), .B(n54206), .Z(n54211) );
  AND U63867 ( .A(n54224), .B(n54225), .Z(n54206) );
  OR U63868 ( .A(n54226), .B(n54227), .Z(n54225) );
  OR U63869 ( .A(n54228), .B(n54229), .Z(n54224) );
  NAND U63870 ( .A(n54230), .B(n54231), .Z(n54207) );
  OR U63871 ( .A(n54232), .B(n54233), .Z(n54230) );
  IV U63872 ( .A(n54234), .Z(n54233) );
  ANDN U63873 ( .B(n54235), .A(n54236), .Z(n54204) );
  XOR U63874 ( .A(n54191), .B(n54237), .Z(n54202) );
  XOR U63875 ( .A(n54192), .B(n54193), .Z(n54237) );
  XNOR U63876 ( .A(n54196), .B(n54197), .Z(n54193) );
  XNOR U63877 ( .A(n54199), .B(n54198), .Z(n54197) );
  AND U63878 ( .A(n54238), .B(n54239), .Z(n54198) );
  NANDN U63879 ( .A(n54240), .B(n54241), .Z(n54239) );
  OR U63880 ( .A(n54242), .B(n54243), .Z(n54238) );
  IV U63881 ( .A(n54244), .Z(n54243) );
  NAND U63882 ( .A(n54245), .B(n54246), .Z(n54199) );
  NANDN U63883 ( .A(n54247), .B(n54248), .Z(n54246) );
  OR U63884 ( .A(n54249), .B(n54250), .Z(n54245) );
  IV U63885 ( .A(n54251), .Z(n54250) );
  ANDN U63886 ( .B(n54252), .A(n54253), .Z(n54196) );
  NOR U63887 ( .A(n54254), .B(n54255), .Z(n54192) );
  XNOR U63888 ( .A(n54185), .B(n54256), .Z(n54191) );
  XNOR U63889 ( .A(n54184), .B(n54186), .Z(n54256) );
  NAND U63890 ( .A(n54257), .B(n54258), .Z(n54186) );
  OR U63891 ( .A(n54259), .B(n54260), .Z(n54258) );
  OR U63892 ( .A(n54261), .B(n54262), .Z(n54257) );
  NAND U63893 ( .A(n54263), .B(n54264), .Z(n54184) );
  OR U63894 ( .A(n54265), .B(n54266), .Z(n54264) );
  OR U63895 ( .A(n54267), .B(n54268), .Z(n54263) );
  ANDN U63896 ( .B(n54269), .A(n54270), .Z(n54185) );
  IV U63897 ( .A(n54271), .Z(n54269) );
  XNOR U63898 ( .A(n54236), .B(n54235), .Z(N60592) );
  XOR U63899 ( .A(n54255), .B(n54254), .Z(n54235) );
  XNOR U63900 ( .A(n54270), .B(n54271), .Z(n54254) );
  XNOR U63901 ( .A(n54265), .B(n54266), .Z(n54271) );
  XNOR U63902 ( .A(n54267), .B(n54268), .Z(n54266) );
  XNOR U63903 ( .A(y[13]), .B(x[13]), .Z(n54268) );
  XNOR U63904 ( .A(y[14]), .B(x[14]), .Z(n54267) );
  XNOR U63905 ( .A(y[12]), .B(x[12]), .Z(n54265) );
  XNOR U63906 ( .A(n54259), .B(n54260), .Z(n54270) );
  XNOR U63907 ( .A(y[9]), .B(x[9]), .Z(n54260) );
  XNOR U63908 ( .A(n54261), .B(n54262), .Z(n54259) );
  XNOR U63909 ( .A(y[10]), .B(x[10]), .Z(n54262) );
  XNOR U63910 ( .A(y[11]), .B(x[11]), .Z(n54261) );
  XOR U63911 ( .A(n54252), .B(n54253), .Z(n54255) );
  XOR U63912 ( .A(n54240), .B(n54241), .Z(n54253) );
  XNOR U63913 ( .A(n54242), .B(n54244), .Z(n54241) );
  XOR U63914 ( .A(y[4]), .B(x[4]), .Z(n54244) );
  XNOR U63915 ( .A(y[5]), .B(x[5]), .Z(n54242) );
  XNOR U63916 ( .A(y[3]), .B(x[3]), .Z(n54240) );
  XNOR U63917 ( .A(n54247), .B(n54248), .Z(n54252) );
  XNOR U63918 ( .A(n54249), .B(n54251), .Z(n54248) );
  XOR U63919 ( .A(y[7]), .B(x[7]), .Z(n54251) );
  XNOR U63920 ( .A(y[8]), .B(x[8]), .Z(n54249) );
  XNOR U63921 ( .A(y[6]), .B(x[6]), .Z(n54247) );
  XOR U63922 ( .A(n54216), .B(n54217), .Z(n54236) );
  XNOR U63923 ( .A(n54232), .B(n54234), .Z(n54217) );
  XOR U63924 ( .A(y[7998]), .B(x[7998]), .Z(n54234) );
  NAND U63925 ( .A(n54272), .B(n54231), .Z(n54232) );
  OR U63926 ( .A(n54273), .B(n54274), .Z(n54231) );
  NAND U63927 ( .A(n54274), .B(n54273), .Z(n54272) );
  XNOR U63928 ( .A(y[7999]), .B(x[7999]), .Z(n54273) );
  XOR U63929 ( .A(n54275), .B(n54226), .Z(n54274) );
  XNOR U63930 ( .A(y[0]), .B(x[0]), .Z(n54226) );
  IV U63931 ( .A(n54227), .Z(n54275) );
  XNOR U63932 ( .A(n54229), .B(n54228), .Z(n54227) );
  XNOR U63933 ( .A(y[1]), .B(x[1]), .Z(n54228) );
  XNOR U63934 ( .A(y[2]), .B(x[2]), .Z(n54229) );
  XNOR U63935 ( .A(n54220), .B(n54221), .Z(n54216) );
  XNOR U63936 ( .A(y[7995]), .B(x[7995]), .Z(n54221) );
  XNOR U63937 ( .A(n54222), .B(n54223), .Z(n54220) );
  XNOR U63938 ( .A(y[7996]), .B(x[7996]), .Z(n54223) );
  XNOR U63939 ( .A(y[7997]), .B(x[7997]), .Z(n54222) );
  NAND U63940 ( .A(n54276), .B(n54277), .Z(N60582) );
  NAND U63941 ( .A(n54278), .B(n54279), .Z(n54277) );
  OR U63942 ( .A(n54280), .B(n54281), .Z(n54278) );
  NANDN U63943 ( .A(n54282), .B(n54280), .Z(n54276) );
  XNOR U63944 ( .A(n54280), .B(n54283), .Z(N60581) );
  XOR U63945 ( .A(n54279), .B(n54282), .Z(n54283) );
  IV U63946 ( .A(n54281), .Z(n54282) );
  NAND U63947 ( .A(n54284), .B(n54285), .Z(n54281) );
  NAND U63948 ( .A(n54286), .B(n54287), .Z(n54285) );
  OR U63949 ( .A(n54288), .B(n54289), .Z(n54286) );
  NANDN U63950 ( .A(n54290), .B(n54288), .Z(n54284) );
  IV U63951 ( .A(n54289), .Z(n54290) );
  NAND U63952 ( .A(n54291), .B(n54292), .Z(n54279) );
  NAND U63953 ( .A(n54293), .B(n54294), .Z(n54292) );
  OR U63954 ( .A(n54295), .B(n54296), .Z(n54293) );
  NAND U63955 ( .A(n54296), .B(n54295), .Z(n54291) );
  NAND U63956 ( .A(n54297), .B(n54298), .Z(n54280) );
  NAND U63957 ( .A(n54299), .B(n54300), .Z(n54298) );
  OR U63958 ( .A(n54301), .B(n54302), .Z(n54299) );
  NANDN U63959 ( .A(n54303), .B(n54301), .Z(n54297) );
  XOR U63960 ( .A(n54294), .B(n54304), .Z(N60580) );
  XOR U63961 ( .A(n54295), .B(n54296), .Z(n54304) );
  XNOR U63962 ( .A(n54301), .B(n54305), .Z(n54296) );
  XOR U63963 ( .A(n54300), .B(n54303), .Z(n54305) );
  IV U63964 ( .A(n54302), .Z(n54303) );
  NAND U63965 ( .A(n54306), .B(n54307), .Z(n54302) );
  OR U63966 ( .A(n54308), .B(n54309), .Z(n54307) );
  OR U63967 ( .A(n54310), .B(n54311), .Z(n54306) );
  NAND U63968 ( .A(n54312), .B(n54313), .Z(n54300) );
  OR U63969 ( .A(n54314), .B(n54315), .Z(n54313) );
  OR U63970 ( .A(n54316), .B(n54317), .Z(n54312) );
  NOR U63971 ( .A(n54318), .B(n54319), .Z(n54301) );
  ANDN U63972 ( .B(n54320), .A(n54321), .Z(n54295) );
  XNOR U63973 ( .A(n54288), .B(n54322), .Z(n54294) );
  XNOR U63974 ( .A(n54287), .B(n54289), .Z(n54322) );
  NAND U63975 ( .A(n54323), .B(n54324), .Z(n54289) );
  OR U63976 ( .A(n54325), .B(n54326), .Z(n54324) );
  IV U63977 ( .A(n54327), .Z(n54326) );
  OR U63978 ( .A(n54328), .B(n54329), .Z(n54323) );
  NAND U63979 ( .A(n54330), .B(n54331), .Z(n54287) );
  OR U63980 ( .A(n54332), .B(n54333), .Z(n54331) );
  OR U63981 ( .A(n54334), .B(n54335), .Z(n54330) );
  AND U63982 ( .A(n54336), .B(n54337), .Z(n54288) );
  IV U63983 ( .A(n54338), .Z(n54337) );
  XNOR U63984 ( .A(n54321), .B(n54320), .Z(N60579) );
  XNOR U63985 ( .A(n54338), .B(n54336), .Z(n54320) );
  XOR U63986 ( .A(n54332), .B(n54333), .Z(n54336) );
  XNOR U63987 ( .A(n54334), .B(n54335), .Z(n54333) );
  XNOR U63988 ( .A(y[7993]), .B(x[7993]), .Z(n54335) );
  XNOR U63989 ( .A(y[7994]), .B(x[7994]), .Z(n54334) );
  XNOR U63990 ( .A(y[7992]), .B(x[7992]), .Z(n54332) );
  XOR U63991 ( .A(n54325), .B(n54327), .Z(n54338) );
  XOR U63992 ( .A(n54328), .B(n54329), .Z(n54327) );
  XNOR U63993 ( .A(y[7990]), .B(x[7990]), .Z(n54329) );
  XNOR U63994 ( .A(y[7991]), .B(x[7991]), .Z(n54328) );
  XNOR U63995 ( .A(y[7989]), .B(x[7989]), .Z(n54325) );
  XNOR U63996 ( .A(n54319), .B(n54318), .Z(n54321) );
  XNOR U63997 ( .A(n54314), .B(n54315), .Z(n54318) );
  XNOR U63998 ( .A(y[7986]), .B(x[7986]), .Z(n54315) );
  XNOR U63999 ( .A(n54316), .B(n54317), .Z(n54314) );
  XNOR U64000 ( .A(y[7987]), .B(x[7987]), .Z(n54317) );
  XNOR U64001 ( .A(y[7988]), .B(x[7988]), .Z(n54316) );
  XNOR U64002 ( .A(n54308), .B(n54309), .Z(n54319) );
  XNOR U64003 ( .A(y[7983]), .B(x[7983]), .Z(n54309) );
  XNOR U64004 ( .A(n54310), .B(n54311), .Z(n54308) );
  XNOR U64005 ( .A(y[7984]), .B(x[7984]), .Z(n54311) );
  XNOR U64006 ( .A(y[7985]), .B(x[7985]), .Z(n54310) );
endmodule

