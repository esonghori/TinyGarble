
module SubBytes ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962;

  XOR U2962 ( .A(n1048), .B(n1011), .Z(n1018) );
  XOR U2963 ( .A(n1690), .B(n1653), .Z(n1660) );
  XOR U2964 ( .A(n467), .B(n430), .Z(n437) );
  XOR U2965 ( .A(n923), .B(n886), .Z(n893) );
  XOR U2966 ( .A(n1565), .B(n1528), .Z(n1535) );
  XOR U2967 ( .A(n290), .B(n253), .Z(n260) );
  XOR U2968 ( .A(n800), .B(n738), .Z(n745) );
  XOR U2969 ( .A(n1442), .B(n1390), .Z(n1397) );
  XOR U2970 ( .A(n1304), .B(n1267), .Z(n1274) );
  XOR U2971 ( .A(n1939), .B(n1900), .Z(n1907) );
  XOR U2972 ( .A(n1427), .B(n775), .Z(n782) );
  XOR U2973 ( .A(n1181), .B(n1144), .Z(n1151) );
  XOR U2974 ( .A(n1814), .B(n1777), .Z(n1784) );
  XOR U2975 ( .A(n622), .B(n585), .Z(n592) );
  XNOR U2976 ( .A(n1011), .B(n1055), .Z(n1030) );
  XNOR U2977 ( .A(n1653), .B(n1697), .Z(n1672) );
  XNOR U2978 ( .A(n430), .B(n474), .Z(n449) );
  XNOR U2979 ( .A(n886), .B(n930), .Z(n905) );
  XNOR U2980 ( .A(n1528), .B(n1572), .Z(n1547) );
  XNOR U2981 ( .A(n253), .B(n297), .Z(n272) );
  XNOR U2982 ( .A(n738), .B(n807), .Z(n757) );
  XNOR U2983 ( .A(n1390), .B(n1449), .Z(n1409) );
  NOR U2984 ( .A(n654), .B(x[9]), .Z(n1) );
  XNOR U2985 ( .A(n329), .B(n328), .Z(n2) );
  XNOR U2986 ( .A(n1), .B(n2), .Z(n3) );
  XNOR U2987 ( .A(n312), .B(n3), .Z(n345) );
  XNOR U2988 ( .A(n1267), .B(n1311), .Z(n1286) );
  XNOR U2989 ( .A(n1900), .B(n1946), .Z(n1919) );
  XNOR U2990 ( .A(n775), .B(n1434), .Z(n794) );
  XNOR U2991 ( .A(n1144), .B(n1188), .Z(n1163) );
  XNOR U2992 ( .A(n1777), .B(n1821), .Z(n1796) );
  XNOR U2993 ( .A(n585), .B(n629), .Z(n604) );
  XOR U2994 ( .A(n163), .B(n134), .Z(n157) );
  XOR U2995 ( .A(n77), .B(n78), .Z(n129) );
  XNOR U2996 ( .A(x[9]), .B(n323), .Z(n318) );
  XOR U2997 ( .A(n1030), .B(n1014), .Z(n1016) );
  XOR U2998 ( .A(n1672), .B(n1656), .Z(n1658) );
  XOR U2999 ( .A(n449), .B(n433), .Z(n435) );
  XOR U3000 ( .A(n905), .B(n889), .Z(n891) );
  XOR U3001 ( .A(n1547), .B(n1531), .Z(n1533) );
  XOR U3002 ( .A(n272), .B(n256), .Z(n258) );
  XOR U3003 ( .A(n757), .B(n741), .Z(n743) );
  XOR U3004 ( .A(n1409), .B(n1393), .Z(n1395) );
  XOR U3005 ( .A(n116), .B(n119), .Z(n4) );
  NANDN U3006 ( .A(n116), .B(n121), .Z(n5) );
  OR U3007 ( .A(n121), .B(n4), .Z(n6) );
  NANDN U3008 ( .A(n117), .B(n6), .Z(n7) );
  NAND U3009 ( .A(n5), .B(n7), .Z(n169) );
  XOR U3010 ( .A(n643), .B(n508), .Z(n511) );
  XOR U3011 ( .A(n1286), .B(n1270), .Z(n1272) );
  XOR U3012 ( .A(n1919), .B(n1903), .Z(n1905) );
  XOR U3013 ( .A(n794), .B(n778), .Z(n780) );
  XOR U3014 ( .A(n1163), .B(n1147), .Z(n1149) );
  XOR U3015 ( .A(n1796), .B(n1780), .Z(n1782) );
  XOR U3016 ( .A(n604), .B(n588), .Z(n590) );
  XOR U3017 ( .A(x[3]), .B(x[1]), .Z(n10) );
  XNOR U3018 ( .A(x[0]), .B(x[6]), .Z(n9) );
  XOR U3019 ( .A(n9), .B(x[2]), .Z(n8) );
  XNOR U3020 ( .A(n10), .B(n8), .Z(n45) );
  XNOR U3021 ( .A(x[5]), .B(n9), .Z(n1432) );
  XOR U3022 ( .A(n1432), .B(x[4]), .Z(n787) );
  IV U3023 ( .A(n787), .Z(n19) );
  XNOR U3024 ( .A(x[7]), .B(x[4]), .Z(n13) );
  XNOR U3025 ( .A(n10), .B(n13), .Z(n73) );
  NOR U3026 ( .A(n19), .B(n73), .Z(n12) );
  XNOR U3027 ( .A(n1432), .B(x[7]), .Z(n1067) );
  XNOR U3028 ( .A(x[2]), .B(n1067), .Z(n28) );
  XNOR U3029 ( .A(x[1]), .B(n28), .Z(n23) );
  AND U3030 ( .A(x[0]), .B(n23), .Z(n11) );
  XNOR U3031 ( .A(n12), .B(n11), .Z(n16) );
  XNOR U3032 ( .A(n45), .B(n1067), .Z(n35) );
  IV U3033 ( .A(n45), .Z(n30) );
  XNOR U3034 ( .A(x[0]), .B(n30), .Z(n50) );
  IV U3035 ( .A(n13), .Z(n777) );
  AND U3036 ( .A(n50), .B(n777), .Z(n18) );
  IV U3037 ( .A(n1432), .Z(n37) );
  XNOR U3038 ( .A(n45), .B(n37), .Z(n67) );
  XOR U3039 ( .A(n67), .B(n73), .Z(n70) );
  XOR U3040 ( .A(x[2]), .B(x[4]), .Z(n779) );
  NAND U3041 ( .A(n70), .B(n779), .Z(n14) );
  XNOR U3042 ( .A(n18), .B(n14), .Z(n39) );
  XNOR U3043 ( .A(n35), .B(n39), .Z(n15) );
  XNOR U3044 ( .A(n16), .B(n15), .Z(n62) );
  XOR U3045 ( .A(x[2]), .B(x[7]), .Z(n793) );
  XNOR U3046 ( .A(x[0]), .B(n73), .Z(n74) );
  XNOR U3047 ( .A(n1432), .B(n74), .Z(n65) );
  NAND U3048 ( .A(n793), .B(n65), .Z(n17) );
  XNOR U3049 ( .A(n18), .B(n17), .Z(n31) );
  IV U3050 ( .A(n23), .Z(n776) );
  XNOR U3051 ( .A(n776), .B(n19), .Z(n783) );
  AND U3052 ( .A(n73), .B(n783), .Z(n21) );
  AND U3053 ( .A(x[0]), .B(n787), .Z(n20) );
  XNOR U3054 ( .A(n21), .B(n20), .Z(n22) );
  NANDN U3055 ( .A(n74), .B(n22), .Z(n26) );
  NAND U3056 ( .A(x[0]), .B(n73), .Z(n24) );
  OR U3057 ( .A(n24), .B(n23), .Z(n25) );
  NAND U3058 ( .A(n26), .B(n25), .Z(n27) );
  XNOR U3059 ( .A(n28), .B(n27), .Z(n29) );
  XNOR U3060 ( .A(n31), .B(n29), .Z(n51) );
  IV U3061 ( .A(n51), .Z(n58) );
  AND U3062 ( .A(n1067), .B(n30), .Z(n33) );
  XOR U3063 ( .A(x[1]), .B(x[7]), .Z(n1069) );
  AND U3064 ( .A(n67), .B(n1069), .Z(n36) );
  XNOR U3065 ( .A(n36), .B(n31), .Z(n32) );
  XNOR U3066 ( .A(n33), .B(n32), .Z(n57) );
  NANDN U3067 ( .A(n58), .B(n57), .Z(n34) );
  NAND U3068 ( .A(n62), .B(n34), .Z(n44) );
  XNOR U3069 ( .A(n36), .B(n35), .Z(n41) );
  ANDN U3070 ( .B(n37), .A(x[1]), .Z(n38) );
  XNOR U3071 ( .A(n39), .B(n38), .Z(n40) );
  XNOR U3072 ( .A(n41), .B(n40), .Z(n54) );
  XOR U3073 ( .A(n57), .B(n54), .Z(n42) );
  NAND U3074 ( .A(n58), .B(n42), .Z(n43) );
  NAND U3075 ( .A(n44), .B(n43), .Z(n1066) );
  ANDN U3076 ( .B(n45), .A(n1066), .Z(n69) );
  IV U3077 ( .A(n54), .Z(n60) );
  XOR U3078 ( .A(n62), .B(n58), .Z(n46) );
  NANDN U3079 ( .A(n60), .B(n46), .Z(n49) );
  NANDN U3080 ( .A(n58), .B(n60), .Z(n47) );
  NANDN U3081 ( .A(n57), .B(n47), .Z(n48) );
  NAND U3082 ( .A(n49), .B(n48), .Z(n1427) );
  XNOR U3083 ( .A(n1066), .B(n1427), .Z(n778) );
  AND U3084 ( .A(n50), .B(n778), .Z(n72) );
  OR U3085 ( .A(n57), .B(n54), .Z(n56) );
  ANDN U3086 ( .B(n57), .A(n51), .Z(n52) );
  XNOR U3087 ( .A(n52), .B(n62), .Z(n53) );
  NAND U3088 ( .A(n54), .B(n53), .Z(n55) );
  NAND U3089 ( .A(n56), .B(n55), .Z(n775) );
  NAND U3090 ( .A(n58), .B(n62), .Z(n64) );
  NAND U3091 ( .A(n58), .B(n57), .Z(n59) );
  XNOR U3092 ( .A(n60), .B(n59), .Z(n61) );
  NANDN U3093 ( .A(n62), .B(n61), .Z(n63) );
  NAND U3094 ( .A(n64), .B(n63), .Z(n1434) );
  NAND U3095 ( .A(n794), .B(n65), .Z(n66) );
  XNOR U3096 ( .A(n72), .B(n66), .Z(n1429) );
  XOR U3097 ( .A(n1066), .B(n1434), .Z(n1068) );
  AND U3098 ( .A(n67), .B(n1068), .Z(n789) );
  XNOR U3099 ( .A(n1429), .B(n789), .Z(n68) );
  XNOR U3100 ( .A(n69), .B(n68), .Z(n1437) );
  NAND U3101 ( .A(n780), .B(n70), .Z(n71) );
  XNOR U3102 ( .A(n72), .B(n71), .Z(n797) );
  AND U3103 ( .A(n73), .B(n782), .Z(n1428) );
  NANDN U3104 ( .A(n74), .B(n775), .Z(n75) );
  XNOR U3105 ( .A(n1428), .B(n75), .Z(n939) );
  XNOR U3106 ( .A(n797), .B(n939), .Z(n786) );
  XOR U3107 ( .A(n1437), .B(n786), .Z(z[0]) );
  XOR U3108 ( .A(x[99]), .B(x[97]), .Z(n76) );
  XNOR U3109 ( .A(n76), .B(x[98]), .Z(n77) );
  XNOR U3110 ( .A(x[101]), .B(n77), .Z(n114) );
  XOR U3111 ( .A(x[98]), .B(x[100]), .Z(n135) );
  XNOR U3112 ( .A(x[102]), .B(n77), .Z(n128) );
  XOR U3113 ( .A(x[103]), .B(x[100]), .Z(n133) );
  XOR U3114 ( .A(n76), .B(n133), .Z(n124) );
  XNOR U3115 ( .A(x[96]), .B(n124), .Z(n93) );
  IV U3116 ( .A(n93), .Z(n125) );
  XNOR U3117 ( .A(x[102]), .B(x[96]), .Z(n78) );
  XNOR U3118 ( .A(x[101]), .B(n78), .Z(n139) );
  XOR U3119 ( .A(n125), .B(n139), .Z(n127) );
  XOR U3120 ( .A(n128), .B(n127), .Z(n156) );
  AND U3121 ( .A(n135), .B(n156), .Z(n80) );
  AND U3122 ( .A(n128), .B(n133), .Z(n86) );
  IV U3123 ( .A(n139), .Z(n102) );
  XNOR U3124 ( .A(x[103]), .B(n102), .Z(n161) );
  XOR U3125 ( .A(n129), .B(n161), .Z(n84) );
  XNOR U3126 ( .A(n86), .B(n84), .Z(n79) );
  XNOR U3127 ( .A(n80), .B(n79), .Z(n103) );
  XOR U3128 ( .A(x[98]), .B(n161), .Z(n98) );
  XOR U3129 ( .A(x[97]), .B(n98), .Z(n150) );
  ANDN U3130 ( .B(x[96]), .A(n150), .Z(n82) );
  XNOR U3131 ( .A(x[100]), .B(n102), .Z(n170) );
  NANDN U3132 ( .A(n124), .B(n170), .Z(n81) );
  XNOR U3133 ( .A(n82), .B(n81), .Z(n83) );
  XOR U3134 ( .A(n103), .B(n83), .Z(n119) );
  XOR U3135 ( .A(x[97]), .B(x[103]), .Z(n138) );
  AND U3136 ( .A(n138), .B(n114), .Z(n104) );
  XOR U3137 ( .A(n84), .B(n104), .Z(n89) );
  XOR U3138 ( .A(x[98]), .B(x[103]), .Z(n162) );
  NAND U3139 ( .A(n162), .B(n127), .Z(n85) );
  XOR U3140 ( .A(n86), .B(n85), .Z(n99) );
  AND U3141 ( .A(n129), .B(n161), .Z(n87) );
  XOR U3142 ( .A(n99), .B(n87), .Z(n88) );
  XNOR U3143 ( .A(n89), .B(n88), .Z(n117) );
  XOR U3144 ( .A(n170), .B(n150), .Z(n152) );
  AND U3145 ( .A(n124), .B(n152), .Z(n91) );
  AND U3146 ( .A(x[96]), .B(n170), .Z(n90) );
  XNOR U3147 ( .A(n91), .B(n90), .Z(n92) );
  NANDN U3148 ( .A(n93), .B(n92), .Z(n96) );
  NAND U3149 ( .A(n124), .B(x[96]), .Z(n94) );
  NANDN U3150 ( .A(n94), .B(n150), .Z(n95) );
  NAND U3151 ( .A(n96), .B(n95), .Z(n97) );
  XNOR U3152 ( .A(n98), .B(n97), .Z(n100) );
  XNOR U3153 ( .A(n100), .B(n99), .Z(n116) );
  OR U3154 ( .A(n117), .B(n116), .Z(n101) );
  NANDN U3155 ( .A(n119), .B(n101), .Z(n109) );
  ANDN U3156 ( .B(n102), .A(x[97]), .Z(n106) );
  XNOR U3157 ( .A(n104), .B(n103), .Z(n105) );
  XNOR U3158 ( .A(n106), .B(n105), .Z(n121) );
  XOR U3159 ( .A(n117), .B(n121), .Z(n107) );
  NAND U3160 ( .A(n116), .B(n107), .Z(n108) );
  NAND U3161 ( .A(n109), .B(n108), .Z(n160) );
  OR U3162 ( .A(n119), .B(n116), .Z(n113) );
  ANDN U3163 ( .B(n116), .A(n117), .Z(n110) );
  XNOR U3164 ( .A(n110), .B(n121), .Z(n111) );
  NAND U3165 ( .A(n119), .B(n111), .Z(n112) );
  NAND U3166 ( .A(n113), .B(n112), .Z(n141) );
  XNOR U3167 ( .A(n160), .B(n141), .Z(n137) );
  AND U3168 ( .A(n114), .B(n137), .Z(n131) );
  NAND U3169 ( .A(n139), .B(n141), .Z(n115) );
  XNOR U3170 ( .A(n131), .B(n115), .Z(n172) );
  NANDN U3171 ( .A(n117), .B(n121), .Z(n123) );
  NANDN U3172 ( .A(n117), .B(n116), .Z(n118) );
  XOR U3173 ( .A(n119), .B(n118), .Z(n120) );
  NANDN U3174 ( .A(n121), .B(n120), .Z(n122) );
  NAND U3175 ( .A(n123), .B(n122), .Z(n149) );
  XOR U3176 ( .A(n169), .B(n149), .Z(n151) );
  AND U3177 ( .A(n124), .B(n151), .Z(n144) );
  NANDN U3178 ( .A(n149), .B(n125), .Z(n126) );
  XNOR U3179 ( .A(n144), .B(n126), .Z(n159) );
  XNOR U3180 ( .A(n172), .B(n159), .Z(z[98]) );
  XNOR U3181 ( .A(n149), .B(n141), .Z(n163) );
  AND U3182 ( .A(n127), .B(n163), .Z(n183) );
  XOR U3183 ( .A(n169), .B(n160), .Z(n134) );
  AND U3184 ( .A(n128), .B(n134), .Z(n181) );
  NANDN U3185 ( .A(n160), .B(n129), .Z(n130) );
  XNOR U3186 ( .A(n131), .B(n130), .Z(n145) );
  XNOR U3187 ( .A(n181), .B(n145), .Z(n132) );
  XNOR U3188 ( .A(n183), .B(n132), .Z(n1958) );
  XOR U3189 ( .A(n1958), .B(z[98]), .Z(z[100]) );
  AND U3190 ( .A(n133), .B(n134), .Z(n165) );
  NAND U3191 ( .A(n157), .B(n135), .Z(n136) );
  XNOR U3192 ( .A(n165), .B(n136), .Z(n153) );
  AND U3193 ( .A(n138), .B(n137), .Z(n166) );
  XOR U3194 ( .A(x[97]), .B(n139), .Z(n140) );
  NAND U3195 ( .A(n141), .B(n140), .Z(n142) );
  XNOR U3196 ( .A(n166), .B(n142), .Z(n147) );
  NANDN U3197 ( .A(n169), .B(x[96]), .Z(n143) );
  XNOR U3198 ( .A(n144), .B(n143), .Z(n180) );
  XNOR U3199 ( .A(n180), .B(n145), .Z(n146) );
  XNOR U3200 ( .A(n147), .B(n146), .Z(n148) );
  XNOR U3201 ( .A(n153), .B(n148), .Z(z[101]) );
  ANDN U3202 ( .B(n150), .A(n149), .Z(n155) );
  AND U3203 ( .A(n152), .B(n151), .Z(n171) );
  XNOR U3204 ( .A(n171), .B(n153), .Z(n154) );
  XNOR U3205 ( .A(n155), .B(n154), .Z(n1959) );
  NAND U3206 ( .A(n157), .B(n156), .Z(n158) );
  XNOR U3207 ( .A(n181), .B(n158), .Z(n175) );
  XNOR U3208 ( .A(n175), .B(n159), .Z(n1957) );
  XNOR U3209 ( .A(n1959), .B(n1957), .Z(n179) );
  ANDN U3210 ( .B(n161), .A(n160), .Z(n168) );
  NAND U3211 ( .A(n163), .B(n162), .Z(n164) );
  XNOR U3212 ( .A(n165), .B(n164), .Z(n176) );
  XNOR U3213 ( .A(n176), .B(n166), .Z(n167) );
  XNOR U3214 ( .A(n168), .B(n167), .Z(n1962) );
  XNOR U3215 ( .A(n179), .B(n1962), .Z(z[102]) );
  ANDN U3216 ( .B(n170), .A(n169), .Z(n174) );
  XNOR U3217 ( .A(n172), .B(n171), .Z(n173) );
  XNOR U3218 ( .A(n174), .B(n173), .Z(n178) );
  XNOR U3219 ( .A(n176), .B(n175), .Z(n177) );
  XNOR U3220 ( .A(n178), .B(n177), .Z(n1960) );
  XNOR U3221 ( .A(n1960), .B(n179), .Z(z[97]) );
  XNOR U3222 ( .A(n181), .B(n180), .Z(n182) );
  XNOR U3223 ( .A(n183), .B(n182), .Z(n184) );
  XOR U3224 ( .A(n184), .B(z[97]), .Z(z[103]) );
  XOR U3225 ( .A(x[107]), .B(x[105]), .Z(n187) );
  XNOR U3226 ( .A(x[104]), .B(x[110]), .Z(n186) );
  XOR U3227 ( .A(n186), .B(x[106]), .Z(n185) );
  XNOR U3228 ( .A(n187), .B(n185), .Z(n222) );
  XNOR U3229 ( .A(x[109]), .B(n186), .Z(n295) );
  XOR U3230 ( .A(n295), .B(x[108]), .Z(n265) );
  IV U3231 ( .A(n265), .Z(n196) );
  XNOR U3232 ( .A(x[111]), .B(x[108]), .Z(n190) );
  XNOR U3233 ( .A(n187), .B(n190), .Z(n250) );
  NOR U3234 ( .A(n196), .B(n250), .Z(n189) );
  XNOR U3235 ( .A(n295), .B(x[111]), .Z(n281) );
  XNOR U3236 ( .A(x[106]), .B(n281), .Z(n205) );
  XNOR U3237 ( .A(x[105]), .B(n205), .Z(n200) );
  AND U3238 ( .A(x[104]), .B(n200), .Z(n188) );
  XNOR U3239 ( .A(n189), .B(n188), .Z(n193) );
  XNOR U3240 ( .A(n222), .B(n281), .Z(n212) );
  IV U3241 ( .A(n222), .Z(n207) );
  XNOR U3242 ( .A(x[104]), .B(n207), .Z(n227) );
  IV U3243 ( .A(n190), .Z(n255) );
  AND U3244 ( .A(n227), .B(n255), .Z(n195) );
  IV U3245 ( .A(n295), .Z(n214) );
  XNOR U3246 ( .A(n222), .B(n214), .Z(n244) );
  XOR U3247 ( .A(n244), .B(n250), .Z(n247) );
  XOR U3248 ( .A(x[106]), .B(x[108]), .Z(n257) );
  NAND U3249 ( .A(n247), .B(n257), .Z(n191) );
  XNOR U3250 ( .A(n195), .B(n191), .Z(n216) );
  XNOR U3251 ( .A(n212), .B(n216), .Z(n192) );
  XNOR U3252 ( .A(n193), .B(n192), .Z(n239) );
  XOR U3253 ( .A(x[106]), .B(x[111]), .Z(n271) );
  XNOR U3254 ( .A(x[104]), .B(n250), .Z(n251) );
  XNOR U3255 ( .A(n295), .B(n251), .Z(n242) );
  NAND U3256 ( .A(n271), .B(n242), .Z(n194) );
  XNOR U3257 ( .A(n195), .B(n194), .Z(n208) );
  IV U3258 ( .A(n200), .Z(n254) );
  XNOR U3259 ( .A(n254), .B(n196), .Z(n261) );
  AND U3260 ( .A(n250), .B(n261), .Z(n198) );
  AND U3261 ( .A(x[104]), .B(n265), .Z(n197) );
  XNOR U3262 ( .A(n198), .B(n197), .Z(n199) );
  NANDN U3263 ( .A(n251), .B(n199), .Z(n203) );
  NAND U3264 ( .A(x[104]), .B(n250), .Z(n201) );
  OR U3265 ( .A(n201), .B(n200), .Z(n202) );
  NAND U3266 ( .A(n203), .B(n202), .Z(n204) );
  XNOR U3267 ( .A(n205), .B(n204), .Z(n206) );
  XNOR U3268 ( .A(n208), .B(n206), .Z(n228) );
  IV U3269 ( .A(n228), .Z(n235) );
  AND U3270 ( .A(n281), .B(n207), .Z(n210) );
  XOR U3271 ( .A(x[105]), .B(x[111]), .Z(n283) );
  AND U3272 ( .A(n244), .B(n283), .Z(n213) );
  XNOR U3273 ( .A(n213), .B(n208), .Z(n209) );
  XNOR U3274 ( .A(n210), .B(n209), .Z(n234) );
  NANDN U3275 ( .A(n235), .B(n234), .Z(n211) );
  NAND U3276 ( .A(n239), .B(n211), .Z(n221) );
  XNOR U3277 ( .A(n213), .B(n212), .Z(n218) );
  ANDN U3278 ( .B(n214), .A(x[105]), .Z(n215) );
  XNOR U3279 ( .A(n216), .B(n215), .Z(n217) );
  XNOR U3280 ( .A(n218), .B(n217), .Z(n231) );
  XOR U3281 ( .A(n234), .B(n231), .Z(n219) );
  NAND U3282 ( .A(n235), .B(n219), .Z(n220) );
  NAND U3283 ( .A(n221), .B(n220), .Z(n280) );
  ANDN U3284 ( .B(n222), .A(n280), .Z(n246) );
  IV U3285 ( .A(n231), .Z(n237) );
  XOR U3286 ( .A(n239), .B(n235), .Z(n223) );
  NANDN U3287 ( .A(n237), .B(n223), .Z(n226) );
  NANDN U3288 ( .A(n235), .B(n237), .Z(n224) );
  NANDN U3289 ( .A(n234), .B(n224), .Z(n225) );
  NAND U3290 ( .A(n226), .B(n225), .Z(n290) );
  XNOR U3291 ( .A(n280), .B(n290), .Z(n256) );
  AND U3292 ( .A(n227), .B(n256), .Z(n249) );
  OR U3293 ( .A(n234), .B(n231), .Z(n233) );
  ANDN U3294 ( .B(n234), .A(n228), .Z(n229) );
  XNOR U3295 ( .A(n229), .B(n239), .Z(n230) );
  NAND U3296 ( .A(n231), .B(n230), .Z(n232) );
  NAND U3297 ( .A(n233), .B(n232), .Z(n253) );
  NAND U3298 ( .A(n235), .B(n239), .Z(n241) );
  NAND U3299 ( .A(n235), .B(n234), .Z(n236) );
  XNOR U3300 ( .A(n237), .B(n236), .Z(n238) );
  NANDN U3301 ( .A(n239), .B(n238), .Z(n240) );
  NAND U3302 ( .A(n241), .B(n240), .Z(n297) );
  NAND U3303 ( .A(n272), .B(n242), .Z(n243) );
  XNOR U3304 ( .A(n249), .B(n243), .Z(n292) );
  XOR U3305 ( .A(n280), .B(n297), .Z(n282) );
  AND U3306 ( .A(n244), .B(n282), .Z(n267) );
  XNOR U3307 ( .A(n292), .B(n267), .Z(n245) );
  XNOR U3308 ( .A(n246), .B(n245), .Z(n300) );
  NAND U3309 ( .A(n258), .B(n247), .Z(n248) );
  XNOR U3310 ( .A(n249), .B(n248), .Z(n275) );
  AND U3311 ( .A(n250), .B(n260), .Z(n291) );
  NANDN U3312 ( .A(n251), .B(n253), .Z(n252) );
  XNOR U3313 ( .A(n291), .B(n252), .Z(n279) );
  XNOR U3314 ( .A(n275), .B(n279), .Z(n264) );
  XOR U3315 ( .A(n300), .B(n264), .Z(z[104]) );
  AND U3316 ( .A(n254), .B(n253), .Z(n263) );
  AND U3317 ( .A(n256), .B(n255), .Z(n274) );
  NAND U3318 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U3319 ( .A(n274), .B(n259), .Z(n301) );
  AND U3320 ( .A(n261), .B(n260), .Z(n268) );
  XNOR U3321 ( .A(n301), .B(n268), .Z(n262) );
  XNOR U3322 ( .A(n263), .B(n262), .Z(n288) );
  XNOR U3323 ( .A(n288), .B(n264), .Z(n360) );
  AND U3324 ( .A(n265), .B(n290), .Z(n270) );
  NANDN U3325 ( .A(n297), .B(n295), .Z(n266) );
  XNOR U3326 ( .A(n267), .B(n266), .Z(n278) );
  XNOR U3327 ( .A(n268), .B(n278), .Z(n269) );
  XNOR U3328 ( .A(n270), .B(n269), .Z(n277) );
  NAND U3329 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U3330 ( .A(n274), .B(n273), .Z(n284) );
  XNOR U3331 ( .A(n275), .B(n284), .Z(n276) );
  XNOR U3332 ( .A(n277), .B(n276), .Z(n287) );
  XNOR U3333 ( .A(n360), .B(n287), .Z(z[105]) );
  XNOR U3334 ( .A(n279), .B(n278), .Z(z[106]) );
  NOR U3335 ( .A(n281), .B(n280), .Z(n286) );
  AND U3336 ( .A(n283), .B(n282), .Z(n299) );
  XNOR U3337 ( .A(n284), .B(n299), .Z(n285) );
  XNOR U3338 ( .A(n286), .B(n285), .Z(n359) );
  XOR U3339 ( .A(n288), .B(n287), .Z(n289) );
  XNOR U3340 ( .A(n359), .B(n289), .Z(z[107]) );
  XOR U3341 ( .A(n300), .B(z[106]), .Z(z[108]) );
  AND U3342 ( .A(x[104]), .B(n290), .Z(n294) );
  XNOR U3343 ( .A(n292), .B(n291), .Z(n293) );
  XNOR U3344 ( .A(n294), .B(n293), .Z(n361) );
  XOR U3345 ( .A(n295), .B(x[105]), .Z(n296) );
  NANDN U3346 ( .A(n297), .B(n296), .Z(n298) );
  XNOR U3347 ( .A(n299), .B(n298), .Z(n303) );
  XNOR U3348 ( .A(n301), .B(n300), .Z(n302) );
  XNOR U3349 ( .A(n303), .B(n302), .Z(n304) );
  XNOR U3350 ( .A(n361), .B(n304), .Z(z[109]) );
  XOR U3351 ( .A(x[9]), .B(x[11]), .Z(n305) );
  XOR U3352 ( .A(x[15]), .B(x[12]), .Z(n486) );
  XOR U3353 ( .A(n305), .B(n486), .Z(n341) );
  XNOR U3354 ( .A(x[8]), .B(x[14]), .Z(n307) );
  XNOR U3355 ( .A(x[13]), .B(n307), .Z(n654) );
  XNOR U3356 ( .A(x[15]), .B(n654), .Z(n485) );
  XNOR U3357 ( .A(n305), .B(x[10]), .Z(n306) );
  XNOR U3358 ( .A(n307), .B(n306), .Z(n308) );
  AND U3359 ( .A(n485), .B(n308), .Z(n311) );
  IV U3360 ( .A(n308), .Z(n641) );
  XOR U3361 ( .A(n641), .B(n654), .Z(n357) );
  XOR U3362 ( .A(x[9]), .B(x[15]), .Z(n491) );
  AND U3363 ( .A(n357), .B(n491), .Z(n312) );
  XNOR U3364 ( .A(x[8]), .B(n308), .Z(n509) );
  AND U3365 ( .A(n486), .B(n509), .Z(n314) );
  XOR U3366 ( .A(x[15]), .B(x[10]), .Z(n488) );
  XNOR U3367 ( .A(n341), .B(x[8]), .Z(n342) );
  XNOR U3368 ( .A(n654), .B(n342), .Z(n642) );
  NAND U3369 ( .A(n488), .B(n642), .Z(n309) );
  XNOR U3370 ( .A(n314), .B(n309), .Z(n325) );
  XNOR U3371 ( .A(n312), .B(n325), .Z(n310) );
  XNOR U3372 ( .A(n311), .B(n310), .Z(n349) );
  XNOR U3373 ( .A(n641), .B(n485), .Z(n329) );
  XOR U3374 ( .A(x[12]), .B(x[10]), .Z(n496) );
  XOR U3375 ( .A(n341), .B(n357), .Z(n510) );
  NAND U3376 ( .A(n496), .B(n510), .Z(n313) );
  XNOR U3377 ( .A(n314), .B(n313), .Z(n328) );
  OR U3378 ( .A(n349), .B(n345), .Z(n335) );
  XNOR U3379 ( .A(x[10]), .B(n485), .Z(n323) );
  IV U3380 ( .A(n318), .Z(n495) );
  XNOR U3381 ( .A(x[12]), .B(n654), .Z(n503) );
  XNOR U3382 ( .A(n495), .B(n503), .Z(n500) );
  AND U3383 ( .A(n341), .B(n500), .Z(n316) );
  ANDN U3384 ( .B(x[8]), .A(n503), .Z(n315) );
  XNOR U3385 ( .A(n316), .B(n315), .Z(n317) );
  NANDN U3386 ( .A(n342), .B(n317), .Z(n321) );
  NAND U3387 ( .A(n341), .B(x[8]), .Z(n319) );
  OR U3388 ( .A(n319), .B(n318), .Z(n320) );
  NAND U3389 ( .A(n321), .B(n320), .Z(n322) );
  XNOR U3390 ( .A(n323), .B(n322), .Z(n324) );
  XNOR U3391 ( .A(n325), .B(n324), .Z(n336) );
  ANDN U3392 ( .B(n349), .A(n336), .Z(n332) );
  NOR U3393 ( .A(n503), .B(n341), .Z(n327) );
  ANDN U3394 ( .B(x[8]), .A(n495), .Z(n326) );
  XNOR U3395 ( .A(n327), .B(n326), .Z(n331) );
  XNOR U3396 ( .A(n329), .B(n328), .Z(n330) );
  XNOR U3397 ( .A(n331), .B(n330), .Z(n354) );
  XNOR U3398 ( .A(n332), .B(n354), .Z(n333) );
  NAND U3399 ( .A(n345), .B(n333), .Z(n334) );
  NAND U3400 ( .A(n335), .B(n334), .Z(n494) );
  IV U3401 ( .A(n494), .Z(n487) );
  IV U3402 ( .A(n345), .Z(n352) );
  IV U3403 ( .A(n336), .Z(n350) );
  XOR U3404 ( .A(n354), .B(n350), .Z(n337) );
  NANDN U3405 ( .A(n352), .B(n337), .Z(n340) );
  NANDN U3406 ( .A(n350), .B(n352), .Z(n338) );
  NANDN U3407 ( .A(n349), .B(n338), .Z(n339) );
  NAND U3408 ( .A(n340), .B(n339), .Z(n649) );
  XNOR U3409 ( .A(n487), .B(n649), .Z(n499) );
  AND U3410 ( .A(n341), .B(n499), .Z(n651) );
  NANDN U3411 ( .A(n342), .B(n494), .Z(n343) );
  XNOR U3412 ( .A(n651), .B(n343), .Z(n663) );
  NANDN U3413 ( .A(n350), .B(n349), .Z(n344) );
  NAND U3414 ( .A(n354), .B(n344), .Z(n348) );
  XOR U3415 ( .A(n349), .B(n345), .Z(n346) );
  NAND U3416 ( .A(n350), .B(n346), .Z(n347) );
  NAND U3417 ( .A(n348), .B(n347), .Z(n640) );
  NAND U3418 ( .A(n350), .B(n354), .Z(n356) );
  NAND U3419 ( .A(n350), .B(n349), .Z(n351) );
  XNOR U3420 ( .A(n352), .B(n351), .Z(n353) );
  NANDN U3421 ( .A(n354), .B(n353), .Z(n355) );
  NAND U3422 ( .A(n356), .B(n355), .Z(n656) );
  XOR U3423 ( .A(n640), .B(n656), .Z(n490) );
  AND U3424 ( .A(n357), .B(n490), .Z(n646) );
  NANDN U3425 ( .A(n656), .B(n654), .Z(n358) );
  XNOR U3426 ( .A(n646), .B(n358), .Z(n513) );
  XNOR U3427 ( .A(n663), .B(n513), .Z(z[10]) );
  XNOR U3428 ( .A(n360), .B(n359), .Z(z[110]) );
  XOR U3429 ( .A(n361), .B(z[105]), .Z(z[111]) );
  XOR U3430 ( .A(x[115]), .B(x[113]), .Z(n364) );
  XNOR U3431 ( .A(x[112]), .B(x[118]), .Z(n363) );
  XOR U3432 ( .A(n363), .B(x[114]), .Z(n362) );
  XNOR U3433 ( .A(n364), .B(n362), .Z(n399) );
  XNOR U3434 ( .A(x[117]), .B(n363), .Z(n472) );
  XOR U3435 ( .A(n472), .B(x[116]), .Z(n442) );
  IV U3436 ( .A(n442), .Z(n373) );
  XNOR U3437 ( .A(x[119]), .B(x[116]), .Z(n367) );
  XNOR U3438 ( .A(n364), .B(n367), .Z(n427) );
  NOR U3439 ( .A(n373), .B(n427), .Z(n366) );
  XNOR U3440 ( .A(n472), .B(x[119]), .Z(n458) );
  XNOR U3441 ( .A(x[114]), .B(n458), .Z(n382) );
  XNOR U3442 ( .A(x[113]), .B(n382), .Z(n377) );
  AND U3443 ( .A(x[112]), .B(n377), .Z(n365) );
  XNOR U3444 ( .A(n366), .B(n365), .Z(n370) );
  XNOR U3445 ( .A(n399), .B(n458), .Z(n389) );
  IV U3446 ( .A(n399), .Z(n384) );
  XNOR U3447 ( .A(x[112]), .B(n384), .Z(n404) );
  IV U3448 ( .A(n367), .Z(n432) );
  AND U3449 ( .A(n404), .B(n432), .Z(n372) );
  IV U3450 ( .A(n472), .Z(n391) );
  XNOR U3451 ( .A(n399), .B(n391), .Z(n421) );
  XOR U3452 ( .A(n421), .B(n427), .Z(n424) );
  XOR U3453 ( .A(x[114]), .B(x[116]), .Z(n434) );
  NAND U3454 ( .A(n424), .B(n434), .Z(n368) );
  XNOR U3455 ( .A(n372), .B(n368), .Z(n393) );
  XNOR U3456 ( .A(n389), .B(n393), .Z(n369) );
  XNOR U3457 ( .A(n370), .B(n369), .Z(n416) );
  XOR U3458 ( .A(x[114]), .B(x[119]), .Z(n448) );
  XNOR U3459 ( .A(x[112]), .B(n427), .Z(n428) );
  XNOR U3460 ( .A(n472), .B(n428), .Z(n419) );
  NAND U3461 ( .A(n448), .B(n419), .Z(n371) );
  XNOR U3462 ( .A(n372), .B(n371), .Z(n385) );
  IV U3463 ( .A(n377), .Z(n431) );
  XNOR U3464 ( .A(n431), .B(n373), .Z(n438) );
  AND U3465 ( .A(n427), .B(n438), .Z(n375) );
  AND U3466 ( .A(x[112]), .B(n442), .Z(n374) );
  XNOR U3467 ( .A(n375), .B(n374), .Z(n376) );
  NANDN U3468 ( .A(n428), .B(n376), .Z(n380) );
  NAND U3469 ( .A(x[112]), .B(n427), .Z(n378) );
  OR U3470 ( .A(n378), .B(n377), .Z(n379) );
  NAND U3471 ( .A(n380), .B(n379), .Z(n381) );
  XNOR U3472 ( .A(n382), .B(n381), .Z(n383) );
  XNOR U3473 ( .A(n385), .B(n383), .Z(n405) );
  IV U3474 ( .A(n405), .Z(n412) );
  AND U3475 ( .A(n458), .B(n384), .Z(n387) );
  XOR U3476 ( .A(x[113]), .B(x[119]), .Z(n460) );
  AND U3477 ( .A(n421), .B(n460), .Z(n390) );
  XNOR U3478 ( .A(n390), .B(n385), .Z(n386) );
  XNOR U3479 ( .A(n387), .B(n386), .Z(n411) );
  NANDN U3480 ( .A(n412), .B(n411), .Z(n388) );
  NAND U3481 ( .A(n416), .B(n388), .Z(n398) );
  XNOR U3482 ( .A(n390), .B(n389), .Z(n395) );
  ANDN U3483 ( .B(n391), .A(x[113]), .Z(n392) );
  XNOR U3484 ( .A(n393), .B(n392), .Z(n394) );
  XNOR U3485 ( .A(n395), .B(n394), .Z(n408) );
  XOR U3486 ( .A(n411), .B(n408), .Z(n396) );
  NAND U3487 ( .A(n412), .B(n396), .Z(n397) );
  NAND U3488 ( .A(n398), .B(n397), .Z(n457) );
  ANDN U3489 ( .B(n399), .A(n457), .Z(n423) );
  IV U3490 ( .A(n408), .Z(n414) );
  XOR U3491 ( .A(n416), .B(n412), .Z(n400) );
  NANDN U3492 ( .A(n414), .B(n400), .Z(n403) );
  NANDN U3493 ( .A(n412), .B(n414), .Z(n401) );
  NANDN U3494 ( .A(n411), .B(n401), .Z(n402) );
  NAND U3495 ( .A(n403), .B(n402), .Z(n467) );
  XNOR U3496 ( .A(n457), .B(n467), .Z(n433) );
  AND U3497 ( .A(n404), .B(n433), .Z(n426) );
  OR U3498 ( .A(n411), .B(n408), .Z(n410) );
  ANDN U3499 ( .B(n411), .A(n405), .Z(n406) );
  XNOR U3500 ( .A(n406), .B(n416), .Z(n407) );
  NAND U3501 ( .A(n408), .B(n407), .Z(n409) );
  NAND U3502 ( .A(n410), .B(n409), .Z(n430) );
  NAND U3503 ( .A(n412), .B(n416), .Z(n418) );
  NAND U3504 ( .A(n412), .B(n411), .Z(n413) );
  XNOR U3505 ( .A(n414), .B(n413), .Z(n415) );
  NANDN U3506 ( .A(n416), .B(n415), .Z(n417) );
  NAND U3507 ( .A(n418), .B(n417), .Z(n474) );
  NAND U3508 ( .A(n449), .B(n419), .Z(n420) );
  XNOR U3509 ( .A(n426), .B(n420), .Z(n469) );
  XOR U3510 ( .A(n457), .B(n474), .Z(n459) );
  AND U3511 ( .A(n421), .B(n459), .Z(n444) );
  XNOR U3512 ( .A(n469), .B(n444), .Z(n422) );
  XNOR U3513 ( .A(n423), .B(n422), .Z(n477) );
  NAND U3514 ( .A(n435), .B(n424), .Z(n425) );
  XNOR U3515 ( .A(n426), .B(n425), .Z(n452) );
  AND U3516 ( .A(n427), .B(n437), .Z(n468) );
  NANDN U3517 ( .A(n428), .B(n430), .Z(n429) );
  XNOR U3518 ( .A(n468), .B(n429), .Z(n456) );
  XNOR U3519 ( .A(n452), .B(n456), .Z(n441) );
  XOR U3520 ( .A(n477), .B(n441), .Z(z[112]) );
  AND U3521 ( .A(n431), .B(n430), .Z(n440) );
  AND U3522 ( .A(n433), .B(n432), .Z(n451) );
  NAND U3523 ( .A(n435), .B(n434), .Z(n436) );
  XNOR U3524 ( .A(n451), .B(n436), .Z(n478) );
  AND U3525 ( .A(n438), .B(n437), .Z(n445) );
  XNOR U3526 ( .A(n478), .B(n445), .Z(n439) );
  XNOR U3527 ( .A(n440), .B(n439), .Z(n465) );
  XNOR U3528 ( .A(n465), .B(n441), .Z(n483) );
  AND U3529 ( .A(n442), .B(n467), .Z(n447) );
  NANDN U3530 ( .A(n474), .B(n472), .Z(n443) );
  XNOR U3531 ( .A(n444), .B(n443), .Z(n455) );
  XNOR U3532 ( .A(n445), .B(n455), .Z(n446) );
  XNOR U3533 ( .A(n447), .B(n446), .Z(n454) );
  NAND U3534 ( .A(n449), .B(n448), .Z(n450) );
  XNOR U3535 ( .A(n451), .B(n450), .Z(n461) );
  XNOR U3536 ( .A(n452), .B(n461), .Z(n453) );
  XNOR U3537 ( .A(n454), .B(n453), .Z(n464) );
  XNOR U3538 ( .A(n483), .B(n464), .Z(z[113]) );
  XNOR U3539 ( .A(n456), .B(n455), .Z(z[114]) );
  NOR U3540 ( .A(n458), .B(n457), .Z(n463) );
  AND U3541 ( .A(n460), .B(n459), .Z(n476) );
  XNOR U3542 ( .A(n461), .B(n476), .Z(n462) );
  XNOR U3543 ( .A(n463), .B(n462), .Z(n482) );
  XOR U3544 ( .A(n465), .B(n464), .Z(n466) );
  XNOR U3545 ( .A(n482), .B(n466), .Z(z[115]) );
  XOR U3546 ( .A(n477), .B(z[114]), .Z(z[116]) );
  AND U3547 ( .A(x[112]), .B(n467), .Z(n471) );
  XNOR U3548 ( .A(n469), .B(n468), .Z(n470) );
  XNOR U3549 ( .A(n471), .B(n470), .Z(n484) );
  XOR U3550 ( .A(n472), .B(x[113]), .Z(n473) );
  NANDN U3551 ( .A(n474), .B(n473), .Z(n475) );
  XNOR U3552 ( .A(n476), .B(n475), .Z(n480) );
  XNOR U3553 ( .A(n478), .B(n477), .Z(n479) );
  XNOR U3554 ( .A(n480), .B(n479), .Z(n481) );
  XNOR U3555 ( .A(n484), .B(n481), .Z(z[117]) );
  XNOR U3556 ( .A(n483), .B(n482), .Z(z[118]) );
  XOR U3557 ( .A(n484), .B(z[113]), .Z(z[119]) );
  NOR U3558 ( .A(n485), .B(n640), .Z(n493) );
  XNOR U3559 ( .A(n640), .B(n649), .Z(n508) );
  AND U3560 ( .A(n486), .B(n508), .Z(n498) );
  XOR U3561 ( .A(n487), .B(n656), .Z(n643) );
  NAND U3562 ( .A(n643), .B(n488), .Z(n489) );
  XNOR U3563 ( .A(n498), .B(n489), .Z(n504) );
  AND U3564 ( .A(n491), .B(n490), .Z(n658) );
  XNOR U3565 ( .A(n504), .B(n658), .Z(n492) );
  XNOR U3566 ( .A(n493), .B(n492), .Z(n666) );
  AND U3567 ( .A(n495), .B(n494), .Z(n502) );
  NAND U3568 ( .A(n511), .B(n496), .Z(n497) );
  XNOR U3569 ( .A(n498), .B(n497), .Z(n659) );
  AND U3570 ( .A(n500), .B(n499), .Z(n505) );
  XNOR U3571 ( .A(n659), .B(n505), .Z(n501) );
  XNOR U3572 ( .A(n502), .B(n501), .Z(n665) );
  ANDN U3573 ( .B(n649), .A(n503), .Z(n507) );
  XNOR U3574 ( .A(n505), .B(n504), .Z(n506) );
  XNOR U3575 ( .A(n507), .B(n506), .Z(n515) );
  AND U3576 ( .A(n509), .B(n508), .Z(n645) );
  NAND U3577 ( .A(n511), .B(n510), .Z(n512) );
  XNOR U3578 ( .A(n645), .B(n512), .Z(n664) );
  XNOR U3579 ( .A(n664), .B(n513), .Z(n514) );
  XNOR U3580 ( .A(n515), .B(n514), .Z(n667) );
  XOR U3581 ( .A(n665), .B(n667), .Z(n516) );
  XNOR U3582 ( .A(n666), .B(n516), .Z(z[11]) );
  XOR U3583 ( .A(x[123]), .B(x[121]), .Z(n519) );
  XNOR U3584 ( .A(x[120]), .B(x[126]), .Z(n518) );
  XOR U3585 ( .A(n518), .B(x[122]), .Z(n517) );
  XNOR U3586 ( .A(n519), .B(n517), .Z(n554) );
  XNOR U3587 ( .A(x[125]), .B(n518), .Z(n627) );
  XOR U3588 ( .A(n627), .B(x[124]), .Z(n597) );
  IV U3589 ( .A(n597), .Z(n528) );
  XNOR U3590 ( .A(x[127]), .B(x[124]), .Z(n522) );
  XNOR U3591 ( .A(n519), .B(n522), .Z(n582) );
  NOR U3592 ( .A(n528), .B(n582), .Z(n521) );
  XNOR U3593 ( .A(n627), .B(x[127]), .Z(n613) );
  XNOR U3594 ( .A(x[122]), .B(n613), .Z(n537) );
  XNOR U3595 ( .A(x[121]), .B(n537), .Z(n532) );
  AND U3596 ( .A(x[120]), .B(n532), .Z(n520) );
  XNOR U3597 ( .A(n521), .B(n520), .Z(n525) );
  XNOR U3598 ( .A(n554), .B(n613), .Z(n544) );
  IV U3599 ( .A(n554), .Z(n539) );
  XNOR U3600 ( .A(x[120]), .B(n539), .Z(n559) );
  IV U3601 ( .A(n522), .Z(n587) );
  AND U3602 ( .A(n559), .B(n587), .Z(n527) );
  IV U3603 ( .A(n627), .Z(n546) );
  XNOR U3604 ( .A(n554), .B(n546), .Z(n576) );
  XOR U3605 ( .A(n576), .B(n582), .Z(n579) );
  XOR U3606 ( .A(x[122]), .B(x[124]), .Z(n589) );
  NAND U3607 ( .A(n579), .B(n589), .Z(n523) );
  XNOR U3608 ( .A(n527), .B(n523), .Z(n548) );
  XNOR U3609 ( .A(n544), .B(n548), .Z(n524) );
  XNOR U3610 ( .A(n525), .B(n524), .Z(n571) );
  XOR U3611 ( .A(x[122]), .B(x[127]), .Z(n603) );
  XNOR U3612 ( .A(x[120]), .B(n582), .Z(n583) );
  XNOR U3613 ( .A(n627), .B(n583), .Z(n574) );
  NAND U3614 ( .A(n603), .B(n574), .Z(n526) );
  XNOR U3615 ( .A(n527), .B(n526), .Z(n540) );
  IV U3616 ( .A(n532), .Z(n586) );
  XNOR U3617 ( .A(n586), .B(n528), .Z(n593) );
  AND U3618 ( .A(n582), .B(n593), .Z(n530) );
  AND U3619 ( .A(x[120]), .B(n597), .Z(n529) );
  XNOR U3620 ( .A(n530), .B(n529), .Z(n531) );
  NANDN U3621 ( .A(n583), .B(n531), .Z(n535) );
  NAND U3622 ( .A(x[120]), .B(n582), .Z(n533) );
  OR U3623 ( .A(n533), .B(n532), .Z(n534) );
  NAND U3624 ( .A(n535), .B(n534), .Z(n536) );
  XNOR U3625 ( .A(n537), .B(n536), .Z(n538) );
  XNOR U3626 ( .A(n540), .B(n538), .Z(n560) );
  IV U3627 ( .A(n560), .Z(n567) );
  AND U3628 ( .A(n613), .B(n539), .Z(n542) );
  XOR U3629 ( .A(x[121]), .B(x[127]), .Z(n615) );
  AND U3630 ( .A(n576), .B(n615), .Z(n545) );
  XNOR U3631 ( .A(n545), .B(n540), .Z(n541) );
  XNOR U3632 ( .A(n542), .B(n541), .Z(n566) );
  NANDN U3633 ( .A(n567), .B(n566), .Z(n543) );
  NAND U3634 ( .A(n571), .B(n543), .Z(n553) );
  XNOR U3635 ( .A(n545), .B(n544), .Z(n550) );
  ANDN U3636 ( .B(n546), .A(x[121]), .Z(n547) );
  XNOR U3637 ( .A(n548), .B(n547), .Z(n549) );
  XNOR U3638 ( .A(n550), .B(n549), .Z(n563) );
  XOR U3639 ( .A(n566), .B(n563), .Z(n551) );
  NAND U3640 ( .A(n567), .B(n551), .Z(n552) );
  NAND U3641 ( .A(n553), .B(n552), .Z(n612) );
  ANDN U3642 ( .B(n554), .A(n612), .Z(n578) );
  IV U3643 ( .A(n563), .Z(n569) );
  XOR U3644 ( .A(n571), .B(n567), .Z(n555) );
  NANDN U3645 ( .A(n569), .B(n555), .Z(n558) );
  NANDN U3646 ( .A(n567), .B(n569), .Z(n556) );
  NANDN U3647 ( .A(n566), .B(n556), .Z(n557) );
  NAND U3648 ( .A(n558), .B(n557), .Z(n622) );
  XNOR U3649 ( .A(n612), .B(n622), .Z(n588) );
  AND U3650 ( .A(n559), .B(n588), .Z(n581) );
  OR U3651 ( .A(n566), .B(n563), .Z(n565) );
  ANDN U3652 ( .B(n566), .A(n560), .Z(n561) );
  XNOR U3653 ( .A(n561), .B(n571), .Z(n562) );
  NAND U3654 ( .A(n563), .B(n562), .Z(n564) );
  NAND U3655 ( .A(n565), .B(n564), .Z(n585) );
  NAND U3656 ( .A(n567), .B(n571), .Z(n573) );
  NAND U3657 ( .A(n567), .B(n566), .Z(n568) );
  XNOR U3658 ( .A(n569), .B(n568), .Z(n570) );
  NANDN U3659 ( .A(n571), .B(n570), .Z(n572) );
  NAND U3660 ( .A(n573), .B(n572), .Z(n629) );
  NAND U3661 ( .A(n604), .B(n574), .Z(n575) );
  XNOR U3662 ( .A(n581), .B(n575), .Z(n624) );
  XOR U3663 ( .A(n612), .B(n629), .Z(n614) );
  AND U3664 ( .A(n576), .B(n614), .Z(n599) );
  XNOR U3665 ( .A(n624), .B(n599), .Z(n577) );
  XNOR U3666 ( .A(n578), .B(n577), .Z(n632) );
  NAND U3667 ( .A(n590), .B(n579), .Z(n580) );
  XNOR U3668 ( .A(n581), .B(n580), .Z(n607) );
  AND U3669 ( .A(n582), .B(n592), .Z(n623) );
  NANDN U3670 ( .A(n583), .B(n585), .Z(n584) );
  XNOR U3671 ( .A(n623), .B(n584), .Z(n611) );
  XNOR U3672 ( .A(n607), .B(n611), .Z(n596) );
  XOR U3673 ( .A(n632), .B(n596), .Z(z[120]) );
  AND U3674 ( .A(n586), .B(n585), .Z(n595) );
  AND U3675 ( .A(n588), .B(n587), .Z(n606) );
  NAND U3676 ( .A(n590), .B(n589), .Z(n591) );
  XNOR U3677 ( .A(n606), .B(n591), .Z(n633) );
  AND U3678 ( .A(n593), .B(n592), .Z(n600) );
  XNOR U3679 ( .A(n633), .B(n600), .Z(n594) );
  XNOR U3680 ( .A(n595), .B(n594), .Z(n620) );
  XNOR U3681 ( .A(n620), .B(n596), .Z(n638) );
  AND U3682 ( .A(n597), .B(n622), .Z(n602) );
  NANDN U3683 ( .A(n629), .B(n627), .Z(n598) );
  XNOR U3684 ( .A(n599), .B(n598), .Z(n610) );
  XNOR U3685 ( .A(n600), .B(n610), .Z(n601) );
  XNOR U3686 ( .A(n602), .B(n601), .Z(n609) );
  NAND U3687 ( .A(n604), .B(n603), .Z(n605) );
  XNOR U3688 ( .A(n606), .B(n605), .Z(n616) );
  XNOR U3689 ( .A(n607), .B(n616), .Z(n608) );
  XNOR U3690 ( .A(n609), .B(n608), .Z(n619) );
  XNOR U3691 ( .A(n638), .B(n619), .Z(z[121]) );
  XNOR U3692 ( .A(n611), .B(n610), .Z(z[122]) );
  NOR U3693 ( .A(n613), .B(n612), .Z(n618) );
  AND U3694 ( .A(n615), .B(n614), .Z(n631) );
  XNOR U3695 ( .A(n616), .B(n631), .Z(n617) );
  XNOR U3696 ( .A(n618), .B(n617), .Z(n637) );
  XOR U3697 ( .A(n620), .B(n619), .Z(n621) );
  XNOR U3698 ( .A(n637), .B(n621), .Z(z[123]) );
  XOR U3699 ( .A(n632), .B(z[122]), .Z(z[124]) );
  AND U3700 ( .A(x[120]), .B(n622), .Z(n626) );
  XNOR U3701 ( .A(n624), .B(n623), .Z(n625) );
  XNOR U3702 ( .A(n626), .B(n625), .Z(n639) );
  XOR U3703 ( .A(n627), .B(x[121]), .Z(n628) );
  NANDN U3704 ( .A(n629), .B(n628), .Z(n630) );
  XNOR U3705 ( .A(n631), .B(n630), .Z(n635) );
  XNOR U3706 ( .A(n633), .B(n632), .Z(n634) );
  XNOR U3707 ( .A(n635), .B(n634), .Z(n636) );
  XNOR U3708 ( .A(n639), .B(n636), .Z(z[125]) );
  XNOR U3709 ( .A(n638), .B(n637), .Z(z[126]) );
  XOR U3710 ( .A(n639), .B(z[121]), .Z(z[127]) );
  ANDN U3711 ( .B(n641), .A(n640), .Z(n648) );
  NAND U3712 ( .A(n643), .B(n642), .Z(n644) );
  XNOR U3713 ( .A(n645), .B(n644), .Z(n650) );
  XNOR U3714 ( .A(n650), .B(n646), .Z(n647) );
  XNOR U3715 ( .A(n648), .B(n647), .Z(n1926) );
  XOR U3716 ( .A(n1926), .B(z[10]), .Z(z[12]) );
  AND U3717 ( .A(x[8]), .B(n649), .Z(n653) );
  XNOR U3718 ( .A(n651), .B(n650), .Z(n652) );
  XNOR U3719 ( .A(n653), .B(n652), .Z(n669) );
  XOR U3720 ( .A(n654), .B(x[9]), .Z(n655) );
  NANDN U3721 ( .A(n656), .B(n655), .Z(n657) );
  XNOR U3722 ( .A(n658), .B(n657), .Z(n661) );
  XNOR U3723 ( .A(n659), .B(n1926), .Z(n660) );
  XNOR U3724 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U3725 ( .A(n669), .B(n662), .Z(z[13]) );
  XNOR U3726 ( .A(n664), .B(n663), .Z(n1925) );
  XNOR U3727 ( .A(n665), .B(n1925), .Z(n668) );
  XNOR U3728 ( .A(n668), .B(n666), .Z(z[14]) );
  XNOR U3729 ( .A(n668), .B(n667), .Z(z[9]) );
  XOR U3730 ( .A(n669), .B(z[9]), .Z(z[15]) );
  XOR U3731 ( .A(x[19]), .B(x[17]), .Z(n672) );
  XNOR U3732 ( .A(x[16]), .B(x[22]), .Z(n671) );
  XOR U3733 ( .A(n671), .B(x[18]), .Z(n670) );
  XNOR U3734 ( .A(n672), .B(n670), .Z(n707) );
  XNOR U3735 ( .A(x[21]), .B(n671), .Z(n805) );
  XOR U3736 ( .A(n805), .B(x[20]), .Z(n750) );
  IV U3737 ( .A(n750), .Z(n681) );
  XNOR U3738 ( .A(x[23]), .B(x[20]), .Z(n675) );
  XNOR U3739 ( .A(n672), .B(n675), .Z(n735) );
  NOR U3740 ( .A(n681), .B(n735), .Z(n674) );
  XNOR U3741 ( .A(n805), .B(x[23]), .Z(n766) );
  XNOR U3742 ( .A(x[18]), .B(n766), .Z(n690) );
  XNOR U3743 ( .A(x[17]), .B(n690), .Z(n685) );
  AND U3744 ( .A(x[16]), .B(n685), .Z(n673) );
  XNOR U3745 ( .A(n674), .B(n673), .Z(n678) );
  XNOR U3746 ( .A(n707), .B(n766), .Z(n697) );
  IV U3747 ( .A(n707), .Z(n692) );
  XNOR U3748 ( .A(x[16]), .B(n692), .Z(n712) );
  IV U3749 ( .A(n675), .Z(n740) );
  AND U3750 ( .A(n712), .B(n740), .Z(n680) );
  IV U3751 ( .A(n805), .Z(n699) );
  XNOR U3752 ( .A(n707), .B(n699), .Z(n729) );
  XOR U3753 ( .A(n729), .B(n735), .Z(n732) );
  XOR U3754 ( .A(x[18]), .B(x[20]), .Z(n742) );
  NAND U3755 ( .A(n732), .B(n742), .Z(n676) );
  XNOR U3756 ( .A(n680), .B(n676), .Z(n701) );
  XNOR U3757 ( .A(n697), .B(n701), .Z(n677) );
  XNOR U3758 ( .A(n678), .B(n677), .Z(n724) );
  XOR U3759 ( .A(x[18]), .B(x[23]), .Z(n756) );
  XNOR U3760 ( .A(x[16]), .B(n735), .Z(n736) );
  XNOR U3761 ( .A(n805), .B(n736), .Z(n727) );
  NAND U3762 ( .A(n756), .B(n727), .Z(n679) );
  XNOR U3763 ( .A(n680), .B(n679), .Z(n693) );
  IV U3764 ( .A(n685), .Z(n739) );
  XNOR U3765 ( .A(n739), .B(n681), .Z(n746) );
  AND U3766 ( .A(n735), .B(n746), .Z(n683) );
  AND U3767 ( .A(x[16]), .B(n750), .Z(n682) );
  XNOR U3768 ( .A(n683), .B(n682), .Z(n684) );
  NANDN U3769 ( .A(n736), .B(n684), .Z(n688) );
  NAND U3770 ( .A(x[16]), .B(n735), .Z(n686) );
  OR U3771 ( .A(n686), .B(n685), .Z(n687) );
  NAND U3772 ( .A(n688), .B(n687), .Z(n689) );
  XNOR U3773 ( .A(n690), .B(n689), .Z(n691) );
  XNOR U3774 ( .A(n693), .B(n691), .Z(n713) );
  IV U3775 ( .A(n713), .Z(n720) );
  AND U3776 ( .A(n766), .B(n692), .Z(n695) );
  XOR U3777 ( .A(x[17]), .B(x[23]), .Z(n768) );
  AND U3778 ( .A(n729), .B(n768), .Z(n698) );
  XNOR U3779 ( .A(n698), .B(n693), .Z(n694) );
  XNOR U3780 ( .A(n695), .B(n694), .Z(n719) );
  NANDN U3781 ( .A(n720), .B(n719), .Z(n696) );
  NAND U3782 ( .A(n724), .B(n696), .Z(n706) );
  XNOR U3783 ( .A(n698), .B(n697), .Z(n703) );
  ANDN U3784 ( .B(n699), .A(x[17]), .Z(n700) );
  XNOR U3785 ( .A(n701), .B(n700), .Z(n702) );
  XNOR U3786 ( .A(n703), .B(n702), .Z(n716) );
  XOR U3787 ( .A(n719), .B(n716), .Z(n704) );
  NAND U3788 ( .A(n720), .B(n704), .Z(n705) );
  NAND U3789 ( .A(n706), .B(n705), .Z(n765) );
  ANDN U3790 ( .B(n707), .A(n765), .Z(n731) );
  IV U3791 ( .A(n716), .Z(n722) );
  XOR U3792 ( .A(n724), .B(n720), .Z(n708) );
  NANDN U3793 ( .A(n722), .B(n708), .Z(n711) );
  NANDN U3794 ( .A(n720), .B(n722), .Z(n709) );
  NANDN U3795 ( .A(n719), .B(n709), .Z(n710) );
  NAND U3796 ( .A(n711), .B(n710), .Z(n800) );
  XNOR U3797 ( .A(n765), .B(n800), .Z(n741) );
  AND U3798 ( .A(n712), .B(n741), .Z(n734) );
  OR U3799 ( .A(n719), .B(n716), .Z(n718) );
  ANDN U3800 ( .B(n719), .A(n713), .Z(n714) );
  XNOR U3801 ( .A(n714), .B(n724), .Z(n715) );
  NAND U3802 ( .A(n716), .B(n715), .Z(n717) );
  NAND U3803 ( .A(n718), .B(n717), .Z(n738) );
  NAND U3804 ( .A(n720), .B(n724), .Z(n726) );
  NAND U3805 ( .A(n720), .B(n719), .Z(n721) );
  XNOR U3806 ( .A(n722), .B(n721), .Z(n723) );
  NANDN U3807 ( .A(n724), .B(n723), .Z(n725) );
  NAND U3808 ( .A(n726), .B(n725), .Z(n807) );
  NAND U3809 ( .A(n757), .B(n727), .Z(n728) );
  XNOR U3810 ( .A(n734), .B(n728), .Z(n802) );
  XOR U3811 ( .A(n765), .B(n807), .Z(n767) );
  AND U3812 ( .A(n729), .B(n767), .Z(n752) );
  XNOR U3813 ( .A(n802), .B(n752), .Z(n730) );
  XNOR U3814 ( .A(n731), .B(n730), .Z(n810) );
  NAND U3815 ( .A(n743), .B(n732), .Z(n733) );
  XNOR U3816 ( .A(n734), .B(n733), .Z(n760) );
  AND U3817 ( .A(n735), .B(n745), .Z(n801) );
  NANDN U3818 ( .A(n736), .B(n738), .Z(n737) );
  XNOR U3819 ( .A(n801), .B(n737), .Z(n764) );
  XNOR U3820 ( .A(n760), .B(n764), .Z(n749) );
  XOR U3821 ( .A(n810), .B(n749), .Z(z[16]) );
  AND U3822 ( .A(n739), .B(n738), .Z(n748) );
  AND U3823 ( .A(n741), .B(n740), .Z(n759) );
  NAND U3824 ( .A(n743), .B(n742), .Z(n744) );
  XNOR U3825 ( .A(n759), .B(n744), .Z(n811) );
  AND U3826 ( .A(n746), .B(n745), .Z(n753) );
  XNOR U3827 ( .A(n811), .B(n753), .Z(n747) );
  XNOR U3828 ( .A(n748), .B(n747), .Z(n773) );
  XNOR U3829 ( .A(n773), .B(n749), .Z(n816) );
  AND U3830 ( .A(n750), .B(n800), .Z(n755) );
  NANDN U3831 ( .A(n807), .B(n805), .Z(n751) );
  XNOR U3832 ( .A(n752), .B(n751), .Z(n763) );
  XNOR U3833 ( .A(n753), .B(n763), .Z(n754) );
  XNOR U3834 ( .A(n755), .B(n754), .Z(n762) );
  NAND U3835 ( .A(n757), .B(n756), .Z(n758) );
  XNOR U3836 ( .A(n759), .B(n758), .Z(n769) );
  XNOR U3837 ( .A(n760), .B(n769), .Z(n761) );
  XNOR U3838 ( .A(n762), .B(n761), .Z(n772) );
  XNOR U3839 ( .A(n816), .B(n772), .Z(z[17]) );
  XNOR U3840 ( .A(n764), .B(n763), .Z(z[18]) );
  NOR U3841 ( .A(n766), .B(n765), .Z(n771) );
  AND U3842 ( .A(n768), .B(n767), .Z(n809) );
  XNOR U3843 ( .A(n769), .B(n809), .Z(n770) );
  XNOR U3844 ( .A(n771), .B(n770), .Z(n815) );
  XOR U3845 ( .A(n773), .B(n772), .Z(n774) );
  XNOR U3846 ( .A(n815), .B(n774), .Z(z[19]) );
  AND U3847 ( .A(n776), .B(n775), .Z(n785) );
  AND U3848 ( .A(n778), .B(n777), .Z(n796) );
  NAND U3849 ( .A(n780), .B(n779), .Z(n781) );
  XNOR U3850 ( .A(n796), .B(n781), .Z(n1438) );
  AND U3851 ( .A(n783), .B(n782), .Z(n790) );
  XNOR U3852 ( .A(n1438), .B(n790), .Z(n784) );
  XNOR U3853 ( .A(n785), .B(n784), .Z(n1074) );
  XNOR U3854 ( .A(n1074), .B(n786), .Z(n1581) );
  AND U3855 ( .A(n787), .B(n1427), .Z(n792) );
  NANDN U3856 ( .A(n1434), .B(n1432), .Z(n788) );
  XNOR U3857 ( .A(n789), .B(n788), .Z(n938) );
  XNOR U3858 ( .A(n790), .B(n938), .Z(n791) );
  XNOR U3859 ( .A(n792), .B(n791), .Z(n799) );
  NAND U3860 ( .A(n794), .B(n793), .Z(n795) );
  XNOR U3861 ( .A(n796), .B(n795), .Z(n1070) );
  XNOR U3862 ( .A(n797), .B(n1070), .Z(n798) );
  XNOR U3863 ( .A(n799), .B(n798), .Z(n1073) );
  XNOR U3864 ( .A(n1581), .B(n1073), .Z(z[1]) );
  XOR U3865 ( .A(n810), .B(z[18]), .Z(z[20]) );
  AND U3866 ( .A(x[16]), .B(n800), .Z(n804) );
  XNOR U3867 ( .A(n802), .B(n801), .Z(n803) );
  XNOR U3868 ( .A(n804), .B(n803), .Z(n817) );
  XOR U3869 ( .A(n805), .B(x[17]), .Z(n806) );
  NANDN U3870 ( .A(n807), .B(n806), .Z(n808) );
  XNOR U3871 ( .A(n809), .B(n808), .Z(n813) );
  XNOR U3872 ( .A(n811), .B(n810), .Z(n812) );
  XNOR U3873 ( .A(n813), .B(n812), .Z(n814) );
  XNOR U3874 ( .A(n817), .B(n814), .Z(z[21]) );
  XNOR U3875 ( .A(n816), .B(n815), .Z(z[22]) );
  XOR U3876 ( .A(n817), .B(z[17]), .Z(z[23]) );
  XOR U3877 ( .A(x[27]), .B(x[25]), .Z(n820) );
  XNOR U3878 ( .A(x[24]), .B(x[30]), .Z(n819) );
  XOR U3879 ( .A(n819), .B(x[26]), .Z(n818) );
  XNOR U3880 ( .A(n820), .B(n818), .Z(n855) );
  XNOR U3881 ( .A(x[29]), .B(n819), .Z(n928) );
  XOR U3882 ( .A(n928), .B(x[28]), .Z(n898) );
  IV U3883 ( .A(n898), .Z(n829) );
  XNOR U3884 ( .A(x[31]), .B(x[28]), .Z(n823) );
  XNOR U3885 ( .A(n820), .B(n823), .Z(n883) );
  NOR U3886 ( .A(n829), .B(n883), .Z(n822) );
  XNOR U3887 ( .A(n928), .B(x[31]), .Z(n914) );
  XNOR U3888 ( .A(x[26]), .B(n914), .Z(n838) );
  XNOR U3889 ( .A(x[25]), .B(n838), .Z(n833) );
  AND U3890 ( .A(x[24]), .B(n833), .Z(n821) );
  XNOR U3891 ( .A(n822), .B(n821), .Z(n826) );
  XNOR U3892 ( .A(n855), .B(n914), .Z(n845) );
  IV U3893 ( .A(n855), .Z(n840) );
  XNOR U3894 ( .A(x[24]), .B(n840), .Z(n860) );
  IV U3895 ( .A(n823), .Z(n888) );
  AND U3896 ( .A(n860), .B(n888), .Z(n828) );
  IV U3897 ( .A(n928), .Z(n847) );
  XNOR U3898 ( .A(n855), .B(n847), .Z(n877) );
  XOR U3899 ( .A(n877), .B(n883), .Z(n880) );
  XOR U3900 ( .A(x[26]), .B(x[28]), .Z(n890) );
  NAND U3901 ( .A(n880), .B(n890), .Z(n824) );
  XNOR U3902 ( .A(n828), .B(n824), .Z(n849) );
  XNOR U3903 ( .A(n845), .B(n849), .Z(n825) );
  XNOR U3904 ( .A(n826), .B(n825), .Z(n872) );
  XOR U3905 ( .A(x[26]), .B(x[31]), .Z(n904) );
  XNOR U3906 ( .A(x[24]), .B(n883), .Z(n884) );
  XNOR U3907 ( .A(n928), .B(n884), .Z(n875) );
  NAND U3908 ( .A(n904), .B(n875), .Z(n827) );
  XNOR U3909 ( .A(n828), .B(n827), .Z(n841) );
  IV U3910 ( .A(n833), .Z(n887) );
  XNOR U3911 ( .A(n887), .B(n829), .Z(n894) );
  AND U3912 ( .A(n883), .B(n894), .Z(n831) );
  AND U3913 ( .A(x[24]), .B(n898), .Z(n830) );
  XNOR U3914 ( .A(n831), .B(n830), .Z(n832) );
  NANDN U3915 ( .A(n884), .B(n832), .Z(n836) );
  NAND U3916 ( .A(x[24]), .B(n883), .Z(n834) );
  OR U3917 ( .A(n834), .B(n833), .Z(n835) );
  NAND U3918 ( .A(n836), .B(n835), .Z(n837) );
  XNOR U3919 ( .A(n838), .B(n837), .Z(n839) );
  XNOR U3920 ( .A(n841), .B(n839), .Z(n861) );
  IV U3921 ( .A(n861), .Z(n868) );
  AND U3922 ( .A(n914), .B(n840), .Z(n843) );
  XOR U3923 ( .A(x[25]), .B(x[31]), .Z(n916) );
  AND U3924 ( .A(n877), .B(n916), .Z(n846) );
  XNOR U3925 ( .A(n846), .B(n841), .Z(n842) );
  XNOR U3926 ( .A(n843), .B(n842), .Z(n867) );
  NANDN U3927 ( .A(n868), .B(n867), .Z(n844) );
  NAND U3928 ( .A(n872), .B(n844), .Z(n854) );
  XNOR U3929 ( .A(n846), .B(n845), .Z(n851) );
  ANDN U3930 ( .B(n847), .A(x[25]), .Z(n848) );
  XNOR U3931 ( .A(n849), .B(n848), .Z(n850) );
  XNOR U3932 ( .A(n851), .B(n850), .Z(n864) );
  XOR U3933 ( .A(n867), .B(n864), .Z(n852) );
  NAND U3934 ( .A(n868), .B(n852), .Z(n853) );
  NAND U3935 ( .A(n854), .B(n853), .Z(n913) );
  ANDN U3936 ( .B(n855), .A(n913), .Z(n879) );
  IV U3937 ( .A(n864), .Z(n870) );
  XOR U3938 ( .A(n872), .B(n868), .Z(n856) );
  NANDN U3939 ( .A(n870), .B(n856), .Z(n859) );
  NANDN U3940 ( .A(n868), .B(n870), .Z(n857) );
  NANDN U3941 ( .A(n867), .B(n857), .Z(n858) );
  NAND U3942 ( .A(n859), .B(n858), .Z(n923) );
  XNOR U3943 ( .A(n913), .B(n923), .Z(n889) );
  AND U3944 ( .A(n860), .B(n889), .Z(n882) );
  OR U3945 ( .A(n867), .B(n864), .Z(n866) );
  ANDN U3946 ( .B(n867), .A(n861), .Z(n862) );
  XNOR U3947 ( .A(n862), .B(n872), .Z(n863) );
  NAND U3948 ( .A(n864), .B(n863), .Z(n865) );
  NAND U3949 ( .A(n866), .B(n865), .Z(n886) );
  NAND U3950 ( .A(n868), .B(n872), .Z(n874) );
  NAND U3951 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U3952 ( .A(n870), .B(n869), .Z(n871) );
  NANDN U3953 ( .A(n872), .B(n871), .Z(n873) );
  NAND U3954 ( .A(n874), .B(n873), .Z(n930) );
  NAND U3955 ( .A(n905), .B(n875), .Z(n876) );
  XNOR U3956 ( .A(n882), .B(n876), .Z(n925) );
  XOR U3957 ( .A(n913), .B(n930), .Z(n915) );
  AND U3958 ( .A(n877), .B(n915), .Z(n900) );
  XNOR U3959 ( .A(n925), .B(n900), .Z(n878) );
  XNOR U3960 ( .A(n879), .B(n878), .Z(n933) );
  NAND U3961 ( .A(n891), .B(n880), .Z(n881) );
  XNOR U3962 ( .A(n882), .B(n881), .Z(n908) );
  AND U3963 ( .A(n883), .B(n893), .Z(n924) );
  NANDN U3964 ( .A(n884), .B(n886), .Z(n885) );
  XNOR U3965 ( .A(n924), .B(n885), .Z(n912) );
  XNOR U3966 ( .A(n908), .B(n912), .Z(n897) );
  XOR U3967 ( .A(n933), .B(n897), .Z(z[24]) );
  AND U3968 ( .A(n887), .B(n886), .Z(n896) );
  AND U3969 ( .A(n889), .B(n888), .Z(n907) );
  NAND U3970 ( .A(n891), .B(n890), .Z(n892) );
  XNOR U3971 ( .A(n907), .B(n892), .Z(n934) );
  AND U3972 ( .A(n894), .B(n893), .Z(n901) );
  XNOR U3973 ( .A(n934), .B(n901), .Z(n895) );
  XNOR U3974 ( .A(n896), .B(n895), .Z(n921) );
  XNOR U3975 ( .A(n921), .B(n897), .Z(n941) );
  AND U3976 ( .A(n898), .B(n923), .Z(n903) );
  NANDN U3977 ( .A(n930), .B(n928), .Z(n899) );
  XNOR U3978 ( .A(n900), .B(n899), .Z(n911) );
  XNOR U3979 ( .A(n901), .B(n911), .Z(n902) );
  XNOR U3980 ( .A(n903), .B(n902), .Z(n910) );
  NAND U3981 ( .A(n905), .B(n904), .Z(n906) );
  XNOR U3982 ( .A(n907), .B(n906), .Z(n917) );
  XNOR U3983 ( .A(n908), .B(n917), .Z(n909) );
  XNOR U3984 ( .A(n910), .B(n909), .Z(n920) );
  XNOR U3985 ( .A(n941), .B(n920), .Z(z[25]) );
  XNOR U3986 ( .A(n912), .B(n911), .Z(z[26]) );
  NOR U3987 ( .A(n914), .B(n913), .Z(n919) );
  AND U3988 ( .A(n916), .B(n915), .Z(n932) );
  XNOR U3989 ( .A(n917), .B(n932), .Z(n918) );
  XNOR U3990 ( .A(n919), .B(n918), .Z(n940) );
  XOR U3991 ( .A(n921), .B(n920), .Z(n922) );
  XNOR U3992 ( .A(n940), .B(n922), .Z(z[27]) );
  XOR U3993 ( .A(n933), .B(z[26]), .Z(z[28]) );
  AND U3994 ( .A(x[24]), .B(n923), .Z(n927) );
  XNOR U3995 ( .A(n925), .B(n924), .Z(n926) );
  XNOR U3996 ( .A(n927), .B(n926), .Z(n942) );
  XOR U3997 ( .A(n928), .B(x[25]), .Z(n929) );
  NANDN U3998 ( .A(n930), .B(n929), .Z(n931) );
  XNOR U3999 ( .A(n932), .B(n931), .Z(n936) );
  XNOR U4000 ( .A(n934), .B(n933), .Z(n935) );
  XNOR U4001 ( .A(n936), .B(n935), .Z(n937) );
  XNOR U4002 ( .A(n942), .B(n937), .Z(z[29]) );
  XNOR U4003 ( .A(n939), .B(n938), .Z(z[2]) );
  XNOR U4004 ( .A(n941), .B(n940), .Z(z[30]) );
  XOR U4005 ( .A(n942), .B(z[25]), .Z(z[31]) );
  XOR U4006 ( .A(x[35]), .B(x[33]), .Z(n945) );
  XNOR U4007 ( .A(x[32]), .B(x[38]), .Z(n944) );
  XOR U4008 ( .A(n944), .B(x[34]), .Z(n943) );
  XNOR U4009 ( .A(n945), .B(n943), .Z(n980) );
  XNOR U4010 ( .A(x[37]), .B(n944), .Z(n1053) );
  XOR U4011 ( .A(n1053), .B(x[36]), .Z(n1023) );
  IV U4012 ( .A(n1023), .Z(n954) );
  XNOR U4013 ( .A(x[39]), .B(x[36]), .Z(n948) );
  XNOR U4014 ( .A(n945), .B(n948), .Z(n1008) );
  NOR U4015 ( .A(n954), .B(n1008), .Z(n947) );
  XNOR U4016 ( .A(n1053), .B(x[39]), .Z(n1039) );
  XNOR U4017 ( .A(x[34]), .B(n1039), .Z(n963) );
  XNOR U4018 ( .A(x[33]), .B(n963), .Z(n958) );
  AND U4019 ( .A(x[32]), .B(n958), .Z(n946) );
  XNOR U4020 ( .A(n947), .B(n946), .Z(n951) );
  XNOR U4021 ( .A(n980), .B(n1039), .Z(n970) );
  IV U4022 ( .A(n980), .Z(n965) );
  XNOR U4023 ( .A(x[32]), .B(n965), .Z(n985) );
  IV U4024 ( .A(n948), .Z(n1013) );
  AND U4025 ( .A(n985), .B(n1013), .Z(n953) );
  IV U4026 ( .A(n1053), .Z(n972) );
  XNOR U4027 ( .A(n980), .B(n972), .Z(n1002) );
  XOR U4028 ( .A(n1002), .B(n1008), .Z(n1005) );
  XOR U4029 ( .A(x[34]), .B(x[36]), .Z(n1015) );
  NAND U4030 ( .A(n1005), .B(n1015), .Z(n949) );
  XNOR U4031 ( .A(n953), .B(n949), .Z(n974) );
  XNOR U4032 ( .A(n970), .B(n974), .Z(n950) );
  XNOR U4033 ( .A(n951), .B(n950), .Z(n997) );
  XOR U4034 ( .A(x[34]), .B(x[39]), .Z(n1029) );
  XNOR U4035 ( .A(x[32]), .B(n1008), .Z(n1009) );
  XNOR U4036 ( .A(n1053), .B(n1009), .Z(n1000) );
  NAND U4037 ( .A(n1029), .B(n1000), .Z(n952) );
  XNOR U4038 ( .A(n953), .B(n952), .Z(n966) );
  IV U4039 ( .A(n958), .Z(n1012) );
  XNOR U4040 ( .A(n1012), .B(n954), .Z(n1019) );
  AND U4041 ( .A(n1008), .B(n1019), .Z(n956) );
  AND U4042 ( .A(x[32]), .B(n1023), .Z(n955) );
  XNOR U4043 ( .A(n956), .B(n955), .Z(n957) );
  NANDN U4044 ( .A(n1009), .B(n957), .Z(n961) );
  NAND U4045 ( .A(x[32]), .B(n1008), .Z(n959) );
  OR U4046 ( .A(n959), .B(n958), .Z(n960) );
  NAND U4047 ( .A(n961), .B(n960), .Z(n962) );
  XNOR U4048 ( .A(n963), .B(n962), .Z(n964) );
  XNOR U4049 ( .A(n966), .B(n964), .Z(n986) );
  IV U4050 ( .A(n986), .Z(n993) );
  AND U4051 ( .A(n1039), .B(n965), .Z(n968) );
  XOR U4052 ( .A(x[33]), .B(x[39]), .Z(n1041) );
  AND U4053 ( .A(n1002), .B(n1041), .Z(n971) );
  XNOR U4054 ( .A(n971), .B(n966), .Z(n967) );
  XNOR U4055 ( .A(n968), .B(n967), .Z(n992) );
  NANDN U4056 ( .A(n993), .B(n992), .Z(n969) );
  NAND U4057 ( .A(n997), .B(n969), .Z(n979) );
  XNOR U4058 ( .A(n971), .B(n970), .Z(n976) );
  ANDN U4059 ( .B(n972), .A(x[33]), .Z(n973) );
  XNOR U4060 ( .A(n974), .B(n973), .Z(n975) );
  XNOR U4061 ( .A(n976), .B(n975), .Z(n989) );
  XOR U4062 ( .A(n992), .B(n989), .Z(n977) );
  NAND U4063 ( .A(n993), .B(n977), .Z(n978) );
  NAND U4064 ( .A(n979), .B(n978), .Z(n1038) );
  ANDN U4065 ( .B(n980), .A(n1038), .Z(n1004) );
  IV U4066 ( .A(n989), .Z(n995) );
  XOR U4067 ( .A(n997), .B(n993), .Z(n981) );
  NANDN U4068 ( .A(n995), .B(n981), .Z(n984) );
  NANDN U4069 ( .A(n993), .B(n995), .Z(n982) );
  NANDN U4070 ( .A(n992), .B(n982), .Z(n983) );
  NAND U4071 ( .A(n984), .B(n983), .Z(n1048) );
  XNOR U4072 ( .A(n1038), .B(n1048), .Z(n1014) );
  AND U4073 ( .A(n985), .B(n1014), .Z(n1007) );
  OR U4074 ( .A(n992), .B(n989), .Z(n991) );
  ANDN U4075 ( .B(n992), .A(n986), .Z(n987) );
  XNOR U4076 ( .A(n987), .B(n997), .Z(n988) );
  NAND U4077 ( .A(n989), .B(n988), .Z(n990) );
  NAND U4078 ( .A(n991), .B(n990), .Z(n1011) );
  NAND U4079 ( .A(n993), .B(n997), .Z(n999) );
  NAND U4080 ( .A(n993), .B(n992), .Z(n994) );
  XNOR U4081 ( .A(n995), .B(n994), .Z(n996) );
  NANDN U4082 ( .A(n997), .B(n996), .Z(n998) );
  NAND U4083 ( .A(n999), .B(n998), .Z(n1055) );
  NAND U4084 ( .A(n1030), .B(n1000), .Z(n1001) );
  XNOR U4085 ( .A(n1007), .B(n1001), .Z(n1050) );
  XOR U4086 ( .A(n1038), .B(n1055), .Z(n1040) );
  AND U4087 ( .A(n1002), .B(n1040), .Z(n1025) );
  XNOR U4088 ( .A(n1050), .B(n1025), .Z(n1003) );
  XNOR U4089 ( .A(n1004), .B(n1003), .Z(n1058) );
  NAND U4090 ( .A(n1016), .B(n1005), .Z(n1006) );
  XNOR U4091 ( .A(n1007), .B(n1006), .Z(n1033) );
  AND U4092 ( .A(n1008), .B(n1018), .Z(n1049) );
  NANDN U4093 ( .A(n1009), .B(n1011), .Z(n1010) );
  XNOR U4094 ( .A(n1049), .B(n1010), .Z(n1037) );
  XNOR U4095 ( .A(n1033), .B(n1037), .Z(n1022) );
  XOR U4096 ( .A(n1058), .B(n1022), .Z(z[32]) );
  AND U4097 ( .A(n1012), .B(n1011), .Z(n1021) );
  AND U4098 ( .A(n1014), .B(n1013), .Z(n1032) );
  NAND U4099 ( .A(n1016), .B(n1015), .Z(n1017) );
  XNOR U4100 ( .A(n1032), .B(n1017), .Z(n1059) );
  AND U4101 ( .A(n1019), .B(n1018), .Z(n1026) );
  XNOR U4102 ( .A(n1059), .B(n1026), .Z(n1020) );
  XNOR U4103 ( .A(n1021), .B(n1020), .Z(n1046) );
  XNOR U4104 ( .A(n1046), .B(n1022), .Z(n1064) );
  AND U4105 ( .A(n1023), .B(n1048), .Z(n1028) );
  NANDN U4106 ( .A(n1055), .B(n1053), .Z(n1024) );
  XNOR U4107 ( .A(n1025), .B(n1024), .Z(n1036) );
  XNOR U4108 ( .A(n1026), .B(n1036), .Z(n1027) );
  XNOR U4109 ( .A(n1028), .B(n1027), .Z(n1035) );
  NAND U4110 ( .A(n1030), .B(n1029), .Z(n1031) );
  XNOR U4111 ( .A(n1032), .B(n1031), .Z(n1042) );
  XNOR U4112 ( .A(n1033), .B(n1042), .Z(n1034) );
  XNOR U4113 ( .A(n1035), .B(n1034), .Z(n1045) );
  XNOR U4114 ( .A(n1064), .B(n1045), .Z(z[33]) );
  XNOR U4115 ( .A(n1037), .B(n1036), .Z(z[34]) );
  NOR U4116 ( .A(n1039), .B(n1038), .Z(n1044) );
  AND U4117 ( .A(n1041), .B(n1040), .Z(n1057) );
  XNOR U4118 ( .A(n1042), .B(n1057), .Z(n1043) );
  XNOR U4119 ( .A(n1044), .B(n1043), .Z(n1063) );
  XOR U4120 ( .A(n1046), .B(n1045), .Z(n1047) );
  XNOR U4121 ( .A(n1063), .B(n1047), .Z(z[35]) );
  XOR U4122 ( .A(n1058), .B(z[34]), .Z(z[36]) );
  AND U4123 ( .A(x[32]), .B(n1048), .Z(n1052) );
  XNOR U4124 ( .A(n1050), .B(n1049), .Z(n1051) );
  XNOR U4125 ( .A(n1052), .B(n1051), .Z(n1065) );
  XOR U4126 ( .A(n1053), .B(x[33]), .Z(n1054) );
  NANDN U4127 ( .A(n1055), .B(n1054), .Z(n1056) );
  XNOR U4128 ( .A(n1057), .B(n1056), .Z(n1061) );
  XNOR U4129 ( .A(n1059), .B(n1058), .Z(n1060) );
  XNOR U4130 ( .A(n1061), .B(n1060), .Z(n1062) );
  XNOR U4131 ( .A(n1065), .B(n1062), .Z(z[37]) );
  XNOR U4132 ( .A(n1064), .B(n1063), .Z(z[38]) );
  XOR U4133 ( .A(n1065), .B(z[33]), .Z(z[39]) );
  NOR U4134 ( .A(n1067), .B(n1066), .Z(n1072) );
  AND U4135 ( .A(n1069), .B(n1068), .Z(n1436) );
  XNOR U4136 ( .A(n1070), .B(n1436), .Z(n1071) );
  XNOR U4137 ( .A(n1072), .B(n1071), .Z(n1580) );
  XOR U4138 ( .A(n1074), .B(n1073), .Z(n1075) );
  XNOR U4139 ( .A(n1580), .B(n1075), .Z(z[3]) );
  XOR U4140 ( .A(x[43]), .B(x[41]), .Z(n1078) );
  XNOR U4141 ( .A(x[40]), .B(x[46]), .Z(n1077) );
  XOR U4142 ( .A(n1077), .B(x[42]), .Z(n1076) );
  XNOR U4143 ( .A(n1078), .B(n1076), .Z(n1113) );
  XNOR U4144 ( .A(x[45]), .B(n1077), .Z(n1186) );
  XOR U4145 ( .A(n1186), .B(x[44]), .Z(n1156) );
  IV U4146 ( .A(n1156), .Z(n1087) );
  XNOR U4147 ( .A(x[47]), .B(x[44]), .Z(n1081) );
  XNOR U4148 ( .A(n1078), .B(n1081), .Z(n1141) );
  NOR U4149 ( .A(n1087), .B(n1141), .Z(n1080) );
  XNOR U4150 ( .A(n1186), .B(x[47]), .Z(n1172) );
  XNOR U4151 ( .A(x[42]), .B(n1172), .Z(n1096) );
  XNOR U4152 ( .A(x[41]), .B(n1096), .Z(n1091) );
  AND U4153 ( .A(x[40]), .B(n1091), .Z(n1079) );
  XNOR U4154 ( .A(n1080), .B(n1079), .Z(n1084) );
  XNOR U4155 ( .A(n1113), .B(n1172), .Z(n1103) );
  IV U4156 ( .A(n1113), .Z(n1098) );
  XNOR U4157 ( .A(x[40]), .B(n1098), .Z(n1118) );
  IV U4158 ( .A(n1081), .Z(n1146) );
  AND U4159 ( .A(n1118), .B(n1146), .Z(n1086) );
  IV U4160 ( .A(n1186), .Z(n1105) );
  XNOR U4161 ( .A(n1113), .B(n1105), .Z(n1135) );
  XOR U4162 ( .A(n1135), .B(n1141), .Z(n1138) );
  XOR U4163 ( .A(x[42]), .B(x[44]), .Z(n1148) );
  NAND U4164 ( .A(n1138), .B(n1148), .Z(n1082) );
  XNOR U4165 ( .A(n1086), .B(n1082), .Z(n1107) );
  XNOR U4166 ( .A(n1103), .B(n1107), .Z(n1083) );
  XNOR U4167 ( .A(n1084), .B(n1083), .Z(n1130) );
  XOR U4168 ( .A(x[42]), .B(x[47]), .Z(n1162) );
  XNOR U4169 ( .A(x[40]), .B(n1141), .Z(n1142) );
  XNOR U4170 ( .A(n1186), .B(n1142), .Z(n1133) );
  NAND U4171 ( .A(n1162), .B(n1133), .Z(n1085) );
  XNOR U4172 ( .A(n1086), .B(n1085), .Z(n1099) );
  IV U4173 ( .A(n1091), .Z(n1145) );
  XNOR U4174 ( .A(n1145), .B(n1087), .Z(n1152) );
  AND U4175 ( .A(n1141), .B(n1152), .Z(n1089) );
  AND U4176 ( .A(x[40]), .B(n1156), .Z(n1088) );
  XNOR U4177 ( .A(n1089), .B(n1088), .Z(n1090) );
  NANDN U4178 ( .A(n1142), .B(n1090), .Z(n1094) );
  NAND U4179 ( .A(x[40]), .B(n1141), .Z(n1092) );
  OR U4180 ( .A(n1092), .B(n1091), .Z(n1093) );
  NAND U4181 ( .A(n1094), .B(n1093), .Z(n1095) );
  XNOR U4182 ( .A(n1096), .B(n1095), .Z(n1097) );
  XNOR U4183 ( .A(n1099), .B(n1097), .Z(n1119) );
  IV U4184 ( .A(n1119), .Z(n1126) );
  AND U4185 ( .A(n1172), .B(n1098), .Z(n1101) );
  XOR U4186 ( .A(x[41]), .B(x[47]), .Z(n1174) );
  AND U4187 ( .A(n1135), .B(n1174), .Z(n1104) );
  XNOR U4188 ( .A(n1104), .B(n1099), .Z(n1100) );
  XNOR U4189 ( .A(n1101), .B(n1100), .Z(n1125) );
  NANDN U4190 ( .A(n1126), .B(n1125), .Z(n1102) );
  NAND U4191 ( .A(n1130), .B(n1102), .Z(n1112) );
  XNOR U4192 ( .A(n1104), .B(n1103), .Z(n1109) );
  ANDN U4193 ( .B(n1105), .A(x[41]), .Z(n1106) );
  XNOR U4194 ( .A(n1107), .B(n1106), .Z(n1108) );
  XNOR U4195 ( .A(n1109), .B(n1108), .Z(n1122) );
  XOR U4196 ( .A(n1125), .B(n1122), .Z(n1110) );
  NAND U4197 ( .A(n1126), .B(n1110), .Z(n1111) );
  NAND U4198 ( .A(n1112), .B(n1111), .Z(n1171) );
  ANDN U4199 ( .B(n1113), .A(n1171), .Z(n1137) );
  IV U4200 ( .A(n1122), .Z(n1128) );
  XOR U4201 ( .A(n1130), .B(n1126), .Z(n1114) );
  NANDN U4202 ( .A(n1128), .B(n1114), .Z(n1117) );
  NANDN U4203 ( .A(n1126), .B(n1128), .Z(n1115) );
  NANDN U4204 ( .A(n1125), .B(n1115), .Z(n1116) );
  NAND U4205 ( .A(n1117), .B(n1116), .Z(n1181) );
  XNOR U4206 ( .A(n1171), .B(n1181), .Z(n1147) );
  AND U4207 ( .A(n1118), .B(n1147), .Z(n1140) );
  OR U4208 ( .A(n1125), .B(n1122), .Z(n1124) );
  ANDN U4209 ( .B(n1125), .A(n1119), .Z(n1120) );
  XNOR U4210 ( .A(n1120), .B(n1130), .Z(n1121) );
  NAND U4211 ( .A(n1122), .B(n1121), .Z(n1123) );
  NAND U4212 ( .A(n1124), .B(n1123), .Z(n1144) );
  NAND U4213 ( .A(n1126), .B(n1130), .Z(n1132) );
  NAND U4214 ( .A(n1126), .B(n1125), .Z(n1127) );
  XNOR U4215 ( .A(n1128), .B(n1127), .Z(n1129) );
  NANDN U4216 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U4217 ( .A(n1132), .B(n1131), .Z(n1188) );
  NAND U4218 ( .A(n1163), .B(n1133), .Z(n1134) );
  XNOR U4219 ( .A(n1140), .B(n1134), .Z(n1183) );
  XOR U4220 ( .A(n1171), .B(n1188), .Z(n1173) );
  AND U4221 ( .A(n1135), .B(n1173), .Z(n1158) );
  XNOR U4222 ( .A(n1183), .B(n1158), .Z(n1136) );
  XNOR U4223 ( .A(n1137), .B(n1136), .Z(n1191) );
  NAND U4224 ( .A(n1149), .B(n1138), .Z(n1139) );
  XNOR U4225 ( .A(n1140), .B(n1139), .Z(n1166) );
  AND U4226 ( .A(n1141), .B(n1151), .Z(n1182) );
  NANDN U4227 ( .A(n1142), .B(n1144), .Z(n1143) );
  XNOR U4228 ( .A(n1182), .B(n1143), .Z(n1170) );
  XNOR U4229 ( .A(n1166), .B(n1170), .Z(n1155) );
  XOR U4230 ( .A(n1191), .B(n1155), .Z(z[40]) );
  AND U4231 ( .A(n1145), .B(n1144), .Z(n1154) );
  AND U4232 ( .A(n1147), .B(n1146), .Z(n1165) );
  NAND U4233 ( .A(n1149), .B(n1148), .Z(n1150) );
  XNOR U4234 ( .A(n1165), .B(n1150), .Z(n1192) );
  AND U4235 ( .A(n1152), .B(n1151), .Z(n1159) );
  XNOR U4236 ( .A(n1192), .B(n1159), .Z(n1153) );
  XNOR U4237 ( .A(n1154), .B(n1153), .Z(n1179) );
  XNOR U4238 ( .A(n1179), .B(n1155), .Z(n1197) );
  AND U4239 ( .A(n1156), .B(n1181), .Z(n1161) );
  NANDN U4240 ( .A(n1188), .B(n1186), .Z(n1157) );
  XNOR U4241 ( .A(n1158), .B(n1157), .Z(n1169) );
  XNOR U4242 ( .A(n1159), .B(n1169), .Z(n1160) );
  XNOR U4243 ( .A(n1161), .B(n1160), .Z(n1168) );
  NAND U4244 ( .A(n1163), .B(n1162), .Z(n1164) );
  XNOR U4245 ( .A(n1165), .B(n1164), .Z(n1175) );
  XNOR U4246 ( .A(n1166), .B(n1175), .Z(n1167) );
  XNOR U4247 ( .A(n1168), .B(n1167), .Z(n1178) );
  XNOR U4248 ( .A(n1197), .B(n1178), .Z(z[41]) );
  XNOR U4249 ( .A(n1170), .B(n1169), .Z(z[42]) );
  NOR U4250 ( .A(n1172), .B(n1171), .Z(n1177) );
  AND U4251 ( .A(n1174), .B(n1173), .Z(n1190) );
  XNOR U4252 ( .A(n1175), .B(n1190), .Z(n1176) );
  XNOR U4253 ( .A(n1177), .B(n1176), .Z(n1196) );
  XOR U4254 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U4255 ( .A(n1196), .B(n1180), .Z(z[43]) );
  XOR U4256 ( .A(n1191), .B(z[42]), .Z(z[44]) );
  AND U4257 ( .A(x[40]), .B(n1181), .Z(n1185) );
  XNOR U4258 ( .A(n1183), .B(n1182), .Z(n1184) );
  XNOR U4259 ( .A(n1185), .B(n1184), .Z(n1198) );
  XOR U4260 ( .A(n1186), .B(x[41]), .Z(n1187) );
  NANDN U4261 ( .A(n1188), .B(n1187), .Z(n1189) );
  XNOR U4262 ( .A(n1190), .B(n1189), .Z(n1194) );
  XNOR U4263 ( .A(n1192), .B(n1191), .Z(n1193) );
  XNOR U4264 ( .A(n1194), .B(n1193), .Z(n1195) );
  XNOR U4265 ( .A(n1198), .B(n1195), .Z(z[45]) );
  XNOR U4266 ( .A(n1197), .B(n1196), .Z(z[46]) );
  XOR U4267 ( .A(n1198), .B(z[41]), .Z(z[47]) );
  XOR U4268 ( .A(x[51]), .B(x[49]), .Z(n1201) );
  XNOR U4269 ( .A(x[48]), .B(x[54]), .Z(n1200) );
  XOR U4270 ( .A(n1200), .B(x[50]), .Z(n1199) );
  XNOR U4271 ( .A(n1201), .B(n1199), .Z(n1236) );
  XNOR U4272 ( .A(x[53]), .B(n1200), .Z(n1309) );
  XOR U4273 ( .A(n1309), .B(x[52]), .Z(n1279) );
  IV U4274 ( .A(n1279), .Z(n1210) );
  XNOR U4275 ( .A(x[55]), .B(x[52]), .Z(n1204) );
  XNOR U4276 ( .A(n1201), .B(n1204), .Z(n1264) );
  NOR U4277 ( .A(n1210), .B(n1264), .Z(n1203) );
  XNOR U4278 ( .A(n1309), .B(x[55]), .Z(n1295) );
  XNOR U4279 ( .A(x[50]), .B(n1295), .Z(n1219) );
  XNOR U4280 ( .A(x[49]), .B(n1219), .Z(n1214) );
  AND U4281 ( .A(x[48]), .B(n1214), .Z(n1202) );
  XNOR U4282 ( .A(n1203), .B(n1202), .Z(n1207) );
  XNOR U4283 ( .A(n1236), .B(n1295), .Z(n1226) );
  IV U4284 ( .A(n1236), .Z(n1221) );
  XNOR U4285 ( .A(x[48]), .B(n1221), .Z(n1241) );
  IV U4286 ( .A(n1204), .Z(n1269) );
  AND U4287 ( .A(n1241), .B(n1269), .Z(n1209) );
  IV U4288 ( .A(n1309), .Z(n1228) );
  XNOR U4289 ( .A(n1236), .B(n1228), .Z(n1258) );
  XOR U4290 ( .A(n1258), .B(n1264), .Z(n1261) );
  XOR U4291 ( .A(x[50]), .B(x[52]), .Z(n1271) );
  NAND U4292 ( .A(n1261), .B(n1271), .Z(n1205) );
  XNOR U4293 ( .A(n1209), .B(n1205), .Z(n1230) );
  XNOR U4294 ( .A(n1226), .B(n1230), .Z(n1206) );
  XNOR U4295 ( .A(n1207), .B(n1206), .Z(n1253) );
  XOR U4296 ( .A(x[50]), .B(x[55]), .Z(n1285) );
  XNOR U4297 ( .A(x[48]), .B(n1264), .Z(n1265) );
  XNOR U4298 ( .A(n1309), .B(n1265), .Z(n1256) );
  NAND U4299 ( .A(n1285), .B(n1256), .Z(n1208) );
  XNOR U4300 ( .A(n1209), .B(n1208), .Z(n1222) );
  IV U4301 ( .A(n1214), .Z(n1268) );
  XNOR U4302 ( .A(n1268), .B(n1210), .Z(n1275) );
  AND U4303 ( .A(n1264), .B(n1275), .Z(n1212) );
  AND U4304 ( .A(x[48]), .B(n1279), .Z(n1211) );
  XNOR U4305 ( .A(n1212), .B(n1211), .Z(n1213) );
  NANDN U4306 ( .A(n1265), .B(n1213), .Z(n1217) );
  NAND U4307 ( .A(x[48]), .B(n1264), .Z(n1215) );
  OR U4308 ( .A(n1215), .B(n1214), .Z(n1216) );
  NAND U4309 ( .A(n1217), .B(n1216), .Z(n1218) );
  XNOR U4310 ( .A(n1219), .B(n1218), .Z(n1220) );
  XNOR U4311 ( .A(n1222), .B(n1220), .Z(n1242) );
  IV U4312 ( .A(n1242), .Z(n1249) );
  AND U4313 ( .A(n1295), .B(n1221), .Z(n1224) );
  XOR U4314 ( .A(x[49]), .B(x[55]), .Z(n1297) );
  AND U4315 ( .A(n1258), .B(n1297), .Z(n1227) );
  XNOR U4316 ( .A(n1227), .B(n1222), .Z(n1223) );
  XNOR U4317 ( .A(n1224), .B(n1223), .Z(n1248) );
  NANDN U4318 ( .A(n1249), .B(n1248), .Z(n1225) );
  NAND U4319 ( .A(n1253), .B(n1225), .Z(n1235) );
  XNOR U4320 ( .A(n1227), .B(n1226), .Z(n1232) );
  ANDN U4321 ( .B(n1228), .A(x[49]), .Z(n1229) );
  XNOR U4322 ( .A(n1230), .B(n1229), .Z(n1231) );
  XNOR U4323 ( .A(n1232), .B(n1231), .Z(n1245) );
  XOR U4324 ( .A(n1248), .B(n1245), .Z(n1233) );
  NAND U4325 ( .A(n1249), .B(n1233), .Z(n1234) );
  NAND U4326 ( .A(n1235), .B(n1234), .Z(n1294) );
  ANDN U4327 ( .B(n1236), .A(n1294), .Z(n1260) );
  IV U4328 ( .A(n1245), .Z(n1251) );
  XOR U4329 ( .A(n1253), .B(n1249), .Z(n1237) );
  NANDN U4330 ( .A(n1251), .B(n1237), .Z(n1240) );
  NANDN U4331 ( .A(n1249), .B(n1251), .Z(n1238) );
  NANDN U4332 ( .A(n1248), .B(n1238), .Z(n1239) );
  NAND U4333 ( .A(n1240), .B(n1239), .Z(n1304) );
  XNOR U4334 ( .A(n1294), .B(n1304), .Z(n1270) );
  AND U4335 ( .A(n1241), .B(n1270), .Z(n1263) );
  OR U4336 ( .A(n1248), .B(n1245), .Z(n1247) );
  ANDN U4337 ( .B(n1248), .A(n1242), .Z(n1243) );
  XNOR U4338 ( .A(n1243), .B(n1253), .Z(n1244) );
  NAND U4339 ( .A(n1245), .B(n1244), .Z(n1246) );
  NAND U4340 ( .A(n1247), .B(n1246), .Z(n1267) );
  NAND U4341 ( .A(n1249), .B(n1253), .Z(n1255) );
  NAND U4342 ( .A(n1249), .B(n1248), .Z(n1250) );
  XNOR U4343 ( .A(n1251), .B(n1250), .Z(n1252) );
  NANDN U4344 ( .A(n1253), .B(n1252), .Z(n1254) );
  NAND U4345 ( .A(n1255), .B(n1254), .Z(n1311) );
  NAND U4346 ( .A(n1286), .B(n1256), .Z(n1257) );
  XNOR U4347 ( .A(n1263), .B(n1257), .Z(n1306) );
  XOR U4348 ( .A(n1294), .B(n1311), .Z(n1296) );
  AND U4349 ( .A(n1258), .B(n1296), .Z(n1281) );
  XNOR U4350 ( .A(n1306), .B(n1281), .Z(n1259) );
  XNOR U4351 ( .A(n1260), .B(n1259), .Z(n1314) );
  NAND U4352 ( .A(n1272), .B(n1261), .Z(n1262) );
  XNOR U4353 ( .A(n1263), .B(n1262), .Z(n1289) );
  AND U4354 ( .A(n1264), .B(n1274), .Z(n1305) );
  NANDN U4355 ( .A(n1265), .B(n1267), .Z(n1266) );
  XNOR U4356 ( .A(n1305), .B(n1266), .Z(n1293) );
  XNOR U4357 ( .A(n1289), .B(n1293), .Z(n1278) );
  XOR U4358 ( .A(n1314), .B(n1278), .Z(z[48]) );
  AND U4359 ( .A(n1268), .B(n1267), .Z(n1277) );
  AND U4360 ( .A(n1270), .B(n1269), .Z(n1288) );
  NAND U4361 ( .A(n1272), .B(n1271), .Z(n1273) );
  XNOR U4362 ( .A(n1288), .B(n1273), .Z(n1315) );
  AND U4363 ( .A(n1275), .B(n1274), .Z(n1282) );
  XNOR U4364 ( .A(n1315), .B(n1282), .Z(n1276) );
  XNOR U4365 ( .A(n1277), .B(n1276), .Z(n1302) );
  XNOR U4366 ( .A(n1302), .B(n1278), .Z(n1320) );
  AND U4367 ( .A(n1279), .B(n1304), .Z(n1284) );
  NANDN U4368 ( .A(n1311), .B(n1309), .Z(n1280) );
  XNOR U4369 ( .A(n1281), .B(n1280), .Z(n1292) );
  XNOR U4370 ( .A(n1282), .B(n1292), .Z(n1283) );
  XNOR U4371 ( .A(n1284), .B(n1283), .Z(n1291) );
  NAND U4372 ( .A(n1286), .B(n1285), .Z(n1287) );
  XNOR U4373 ( .A(n1288), .B(n1287), .Z(n1298) );
  XNOR U4374 ( .A(n1289), .B(n1298), .Z(n1290) );
  XNOR U4375 ( .A(n1291), .B(n1290), .Z(n1301) );
  XNOR U4376 ( .A(n1320), .B(n1301), .Z(z[49]) );
  XOR U4377 ( .A(n1437), .B(z[2]), .Z(z[4]) );
  XNOR U4378 ( .A(n1293), .B(n1292), .Z(z[50]) );
  NOR U4379 ( .A(n1295), .B(n1294), .Z(n1300) );
  AND U4380 ( .A(n1297), .B(n1296), .Z(n1313) );
  XNOR U4381 ( .A(n1298), .B(n1313), .Z(n1299) );
  XNOR U4382 ( .A(n1300), .B(n1299), .Z(n1319) );
  XOR U4383 ( .A(n1302), .B(n1301), .Z(n1303) );
  XNOR U4384 ( .A(n1319), .B(n1303), .Z(z[51]) );
  XOR U4385 ( .A(n1314), .B(z[50]), .Z(z[52]) );
  AND U4386 ( .A(x[48]), .B(n1304), .Z(n1308) );
  XNOR U4387 ( .A(n1306), .B(n1305), .Z(n1307) );
  XNOR U4388 ( .A(n1308), .B(n1307), .Z(n1321) );
  XOR U4389 ( .A(n1309), .B(x[49]), .Z(n1310) );
  NANDN U4390 ( .A(n1311), .B(n1310), .Z(n1312) );
  XNOR U4391 ( .A(n1313), .B(n1312), .Z(n1317) );
  XNOR U4392 ( .A(n1315), .B(n1314), .Z(n1316) );
  XNOR U4393 ( .A(n1317), .B(n1316), .Z(n1318) );
  XNOR U4394 ( .A(n1321), .B(n1318), .Z(z[53]) );
  XNOR U4395 ( .A(n1320), .B(n1319), .Z(z[54]) );
  XOR U4396 ( .A(n1321), .B(z[49]), .Z(z[55]) );
  XOR U4397 ( .A(x[59]), .B(x[57]), .Z(n1324) );
  XNOR U4398 ( .A(x[56]), .B(x[62]), .Z(n1323) );
  XOR U4399 ( .A(n1323), .B(x[58]), .Z(n1322) );
  XNOR U4400 ( .A(n1324), .B(n1322), .Z(n1359) );
  XNOR U4401 ( .A(x[61]), .B(n1323), .Z(n1447) );
  XOR U4402 ( .A(n1447), .B(x[60]), .Z(n1402) );
  IV U4403 ( .A(n1402), .Z(n1333) );
  XNOR U4404 ( .A(x[63]), .B(x[60]), .Z(n1327) );
  XNOR U4405 ( .A(n1324), .B(n1327), .Z(n1387) );
  NOR U4406 ( .A(n1333), .B(n1387), .Z(n1326) );
  XNOR U4407 ( .A(n1447), .B(x[63]), .Z(n1418) );
  XNOR U4408 ( .A(x[58]), .B(n1418), .Z(n1342) );
  XNOR U4409 ( .A(x[57]), .B(n1342), .Z(n1337) );
  AND U4410 ( .A(x[56]), .B(n1337), .Z(n1325) );
  XNOR U4411 ( .A(n1326), .B(n1325), .Z(n1330) );
  XNOR U4412 ( .A(n1359), .B(n1418), .Z(n1349) );
  IV U4413 ( .A(n1359), .Z(n1344) );
  XNOR U4414 ( .A(x[56]), .B(n1344), .Z(n1364) );
  IV U4415 ( .A(n1327), .Z(n1392) );
  AND U4416 ( .A(n1364), .B(n1392), .Z(n1332) );
  IV U4417 ( .A(n1447), .Z(n1351) );
  XNOR U4418 ( .A(n1359), .B(n1351), .Z(n1381) );
  XOR U4419 ( .A(n1381), .B(n1387), .Z(n1384) );
  XOR U4420 ( .A(x[58]), .B(x[60]), .Z(n1394) );
  NAND U4421 ( .A(n1384), .B(n1394), .Z(n1328) );
  XNOR U4422 ( .A(n1332), .B(n1328), .Z(n1353) );
  XNOR U4423 ( .A(n1349), .B(n1353), .Z(n1329) );
  XNOR U4424 ( .A(n1330), .B(n1329), .Z(n1376) );
  XOR U4425 ( .A(x[58]), .B(x[63]), .Z(n1408) );
  XNOR U4426 ( .A(x[56]), .B(n1387), .Z(n1388) );
  XNOR U4427 ( .A(n1447), .B(n1388), .Z(n1379) );
  NAND U4428 ( .A(n1408), .B(n1379), .Z(n1331) );
  XNOR U4429 ( .A(n1332), .B(n1331), .Z(n1345) );
  IV U4430 ( .A(n1337), .Z(n1391) );
  XNOR U4431 ( .A(n1391), .B(n1333), .Z(n1398) );
  AND U4432 ( .A(n1387), .B(n1398), .Z(n1335) );
  AND U4433 ( .A(x[56]), .B(n1402), .Z(n1334) );
  XNOR U4434 ( .A(n1335), .B(n1334), .Z(n1336) );
  NANDN U4435 ( .A(n1388), .B(n1336), .Z(n1340) );
  NAND U4436 ( .A(x[56]), .B(n1387), .Z(n1338) );
  OR U4437 ( .A(n1338), .B(n1337), .Z(n1339) );
  NAND U4438 ( .A(n1340), .B(n1339), .Z(n1341) );
  XNOR U4439 ( .A(n1342), .B(n1341), .Z(n1343) );
  XNOR U4440 ( .A(n1345), .B(n1343), .Z(n1365) );
  IV U4441 ( .A(n1365), .Z(n1372) );
  AND U4442 ( .A(n1418), .B(n1344), .Z(n1347) );
  XOR U4443 ( .A(x[57]), .B(x[63]), .Z(n1420) );
  AND U4444 ( .A(n1381), .B(n1420), .Z(n1350) );
  XNOR U4445 ( .A(n1350), .B(n1345), .Z(n1346) );
  XNOR U4446 ( .A(n1347), .B(n1346), .Z(n1371) );
  NANDN U4447 ( .A(n1372), .B(n1371), .Z(n1348) );
  NAND U4448 ( .A(n1376), .B(n1348), .Z(n1358) );
  XNOR U4449 ( .A(n1350), .B(n1349), .Z(n1355) );
  ANDN U4450 ( .B(n1351), .A(x[57]), .Z(n1352) );
  XNOR U4451 ( .A(n1353), .B(n1352), .Z(n1354) );
  XNOR U4452 ( .A(n1355), .B(n1354), .Z(n1368) );
  XOR U4453 ( .A(n1371), .B(n1368), .Z(n1356) );
  NAND U4454 ( .A(n1372), .B(n1356), .Z(n1357) );
  NAND U4455 ( .A(n1358), .B(n1357), .Z(n1417) );
  ANDN U4456 ( .B(n1359), .A(n1417), .Z(n1383) );
  IV U4457 ( .A(n1368), .Z(n1374) );
  XOR U4458 ( .A(n1376), .B(n1372), .Z(n1360) );
  NANDN U4459 ( .A(n1374), .B(n1360), .Z(n1363) );
  NANDN U4460 ( .A(n1372), .B(n1374), .Z(n1361) );
  NANDN U4461 ( .A(n1371), .B(n1361), .Z(n1362) );
  NAND U4462 ( .A(n1363), .B(n1362), .Z(n1442) );
  XNOR U4463 ( .A(n1417), .B(n1442), .Z(n1393) );
  AND U4464 ( .A(n1364), .B(n1393), .Z(n1386) );
  OR U4465 ( .A(n1371), .B(n1368), .Z(n1370) );
  ANDN U4466 ( .B(n1371), .A(n1365), .Z(n1366) );
  XNOR U4467 ( .A(n1366), .B(n1376), .Z(n1367) );
  NAND U4468 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U4469 ( .A(n1370), .B(n1369), .Z(n1390) );
  NAND U4470 ( .A(n1372), .B(n1376), .Z(n1378) );
  NAND U4471 ( .A(n1372), .B(n1371), .Z(n1373) );
  XNOR U4472 ( .A(n1374), .B(n1373), .Z(n1375) );
  NANDN U4473 ( .A(n1376), .B(n1375), .Z(n1377) );
  NAND U4474 ( .A(n1378), .B(n1377), .Z(n1449) );
  NAND U4475 ( .A(n1409), .B(n1379), .Z(n1380) );
  XNOR U4476 ( .A(n1386), .B(n1380), .Z(n1444) );
  XOR U4477 ( .A(n1417), .B(n1449), .Z(n1419) );
  AND U4478 ( .A(n1381), .B(n1419), .Z(n1404) );
  XNOR U4479 ( .A(n1444), .B(n1404), .Z(n1382) );
  XNOR U4480 ( .A(n1383), .B(n1382), .Z(n1452) );
  NAND U4481 ( .A(n1395), .B(n1384), .Z(n1385) );
  XNOR U4482 ( .A(n1386), .B(n1385), .Z(n1412) );
  AND U4483 ( .A(n1387), .B(n1397), .Z(n1443) );
  NANDN U4484 ( .A(n1388), .B(n1390), .Z(n1389) );
  XNOR U4485 ( .A(n1443), .B(n1389), .Z(n1416) );
  XNOR U4486 ( .A(n1412), .B(n1416), .Z(n1401) );
  XOR U4487 ( .A(n1452), .B(n1401), .Z(z[56]) );
  AND U4488 ( .A(n1391), .B(n1390), .Z(n1400) );
  AND U4489 ( .A(n1393), .B(n1392), .Z(n1411) );
  NAND U4490 ( .A(n1395), .B(n1394), .Z(n1396) );
  XNOR U4491 ( .A(n1411), .B(n1396), .Z(n1453) );
  AND U4492 ( .A(n1398), .B(n1397), .Z(n1405) );
  XNOR U4493 ( .A(n1453), .B(n1405), .Z(n1399) );
  XNOR U4494 ( .A(n1400), .B(n1399), .Z(n1425) );
  XNOR U4495 ( .A(n1425), .B(n1401), .Z(n1458) );
  AND U4496 ( .A(n1402), .B(n1442), .Z(n1407) );
  NANDN U4497 ( .A(n1449), .B(n1447), .Z(n1403) );
  XNOR U4498 ( .A(n1404), .B(n1403), .Z(n1415) );
  XNOR U4499 ( .A(n1405), .B(n1415), .Z(n1406) );
  XNOR U4500 ( .A(n1407), .B(n1406), .Z(n1414) );
  NAND U4501 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U4502 ( .A(n1411), .B(n1410), .Z(n1421) );
  XNOR U4503 ( .A(n1412), .B(n1421), .Z(n1413) );
  XNOR U4504 ( .A(n1414), .B(n1413), .Z(n1424) );
  XNOR U4505 ( .A(n1458), .B(n1424), .Z(z[57]) );
  XNOR U4506 ( .A(n1416), .B(n1415), .Z(z[58]) );
  NOR U4507 ( .A(n1418), .B(n1417), .Z(n1423) );
  AND U4508 ( .A(n1420), .B(n1419), .Z(n1451) );
  XNOR U4509 ( .A(n1421), .B(n1451), .Z(n1422) );
  XNOR U4510 ( .A(n1423), .B(n1422), .Z(n1457) );
  XOR U4511 ( .A(n1425), .B(n1424), .Z(n1426) );
  XNOR U4512 ( .A(n1457), .B(n1426), .Z(z[59]) );
  AND U4513 ( .A(x[0]), .B(n1427), .Z(n1431) );
  XNOR U4514 ( .A(n1429), .B(n1428), .Z(n1430) );
  XNOR U4515 ( .A(n1431), .B(n1430), .Z(n1708) );
  XOR U4516 ( .A(n1432), .B(x[1]), .Z(n1433) );
  NANDN U4517 ( .A(n1434), .B(n1433), .Z(n1435) );
  XNOR U4518 ( .A(n1436), .B(n1435), .Z(n1440) );
  XNOR U4519 ( .A(n1438), .B(n1437), .Z(n1439) );
  XNOR U4520 ( .A(n1440), .B(n1439), .Z(n1441) );
  XNOR U4521 ( .A(n1708), .B(n1441), .Z(z[5]) );
  XOR U4522 ( .A(n1452), .B(z[58]), .Z(z[60]) );
  AND U4523 ( .A(x[56]), .B(n1442), .Z(n1446) );
  XNOR U4524 ( .A(n1444), .B(n1443), .Z(n1445) );
  XNOR U4525 ( .A(n1446), .B(n1445), .Z(n1459) );
  XOR U4526 ( .A(n1447), .B(x[57]), .Z(n1448) );
  NANDN U4527 ( .A(n1449), .B(n1448), .Z(n1450) );
  XNOR U4528 ( .A(n1451), .B(n1450), .Z(n1455) );
  XNOR U4529 ( .A(n1453), .B(n1452), .Z(n1454) );
  XNOR U4530 ( .A(n1455), .B(n1454), .Z(n1456) );
  XNOR U4531 ( .A(n1459), .B(n1456), .Z(z[61]) );
  XNOR U4532 ( .A(n1458), .B(n1457), .Z(z[62]) );
  XOR U4533 ( .A(n1459), .B(z[57]), .Z(z[63]) );
  XOR U4534 ( .A(x[67]), .B(x[65]), .Z(n1462) );
  XNOR U4535 ( .A(x[64]), .B(x[70]), .Z(n1461) );
  XOR U4536 ( .A(n1461), .B(x[66]), .Z(n1460) );
  XNOR U4537 ( .A(n1462), .B(n1460), .Z(n1497) );
  XNOR U4538 ( .A(x[69]), .B(n1461), .Z(n1570) );
  XOR U4539 ( .A(n1570), .B(x[68]), .Z(n1540) );
  IV U4540 ( .A(n1540), .Z(n1471) );
  XNOR U4541 ( .A(x[71]), .B(x[68]), .Z(n1465) );
  XNOR U4542 ( .A(n1462), .B(n1465), .Z(n1525) );
  NOR U4543 ( .A(n1471), .B(n1525), .Z(n1464) );
  XNOR U4544 ( .A(n1570), .B(x[71]), .Z(n1556) );
  XNOR U4545 ( .A(x[66]), .B(n1556), .Z(n1480) );
  XNOR U4546 ( .A(x[65]), .B(n1480), .Z(n1475) );
  AND U4547 ( .A(x[64]), .B(n1475), .Z(n1463) );
  XNOR U4548 ( .A(n1464), .B(n1463), .Z(n1468) );
  XNOR U4549 ( .A(n1497), .B(n1556), .Z(n1487) );
  IV U4550 ( .A(n1497), .Z(n1482) );
  XNOR U4551 ( .A(x[64]), .B(n1482), .Z(n1502) );
  IV U4552 ( .A(n1465), .Z(n1530) );
  AND U4553 ( .A(n1502), .B(n1530), .Z(n1470) );
  IV U4554 ( .A(n1570), .Z(n1489) );
  XNOR U4555 ( .A(n1497), .B(n1489), .Z(n1519) );
  XOR U4556 ( .A(n1519), .B(n1525), .Z(n1522) );
  XOR U4557 ( .A(x[66]), .B(x[68]), .Z(n1532) );
  NAND U4558 ( .A(n1522), .B(n1532), .Z(n1466) );
  XNOR U4559 ( .A(n1470), .B(n1466), .Z(n1491) );
  XNOR U4560 ( .A(n1487), .B(n1491), .Z(n1467) );
  XNOR U4561 ( .A(n1468), .B(n1467), .Z(n1514) );
  XOR U4562 ( .A(x[66]), .B(x[71]), .Z(n1546) );
  XNOR U4563 ( .A(x[64]), .B(n1525), .Z(n1526) );
  XNOR U4564 ( .A(n1570), .B(n1526), .Z(n1517) );
  NAND U4565 ( .A(n1546), .B(n1517), .Z(n1469) );
  XNOR U4566 ( .A(n1470), .B(n1469), .Z(n1483) );
  IV U4567 ( .A(n1475), .Z(n1529) );
  XNOR U4568 ( .A(n1529), .B(n1471), .Z(n1536) );
  AND U4569 ( .A(n1525), .B(n1536), .Z(n1473) );
  AND U4570 ( .A(x[64]), .B(n1540), .Z(n1472) );
  XNOR U4571 ( .A(n1473), .B(n1472), .Z(n1474) );
  NANDN U4572 ( .A(n1526), .B(n1474), .Z(n1478) );
  NAND U4573 ( .A(x[64]), .B(n1525), .Z(n1476) );
  OR U4574 ( .A(n1476), .B(n1475), .Z(n1477) );
  NAND U4575 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U4576 ( .A(n1480), .B(n1479), .Z(n1481) );
  XNOR U4577 ( .A(n1483), .B(n1481), .Z(n1503) );
  IV U4578 ( .A(n1503), .Z(n1510) );
  AND U4579 ( .A(n1556), .B(n1482), .Z(n1485) );
  XOR U4580 ( .A(x[65]), .B(x[71]), .Z(n1558) );
  AND U4581 ( .A(n1519), .B(n1558), .Z(n1488) );
  XNOR U4582 ( .A(n1488), .B(n1483), .Z(n1484) );
  XNOR U4583 ( .A(n1485), .B(n1484), .Z(n1509) );
  NANDN U4584 ( .A(n1510), .B(n1509), .Z(n1486) );
  NAND U4585 ( .A(n1514), .B(n1486), .Z(n1496) );
  XNOR U4586 ( .A(n1488), .B(n1487), .Z(n1493) );
  ANDN U4587 ( .B(n1489), .A(x[65]), .Z(n1490) );
  XNOR U4588 ( .A(n1491), .B(n1490), .Z(n1492) );
  XNOR U4589 ( .A(n1493), .B(n1492), .Z(n1506) );
  XOR U4590 ( .A(n1509), .B(n1506), .Z(n1494) );
  NAND U4591 ( .A(n1510), .B(n1494), .Z(n1495) );
  NAND U4592 ( .A(n1496), .B(n1495), .Z(n1555) );
  ANDN U4593 ( .B(n1497), .A(n1555), .Z(n1521) );
  IV U4594 ( .A(n1506), .Z(n1512) );
  XOR U4595 ( .A(n1514), .B(n1510), .Z(n1498) );
  NANDN U4596 ( .A(n1512), .B(n1498), .Z(n1501) );
  NANDN U4597 ( .A(n1510), .B(n1512), .Z(n1499) );
  NANDN U4598 ( .A(n1509), .B(n1499), .Z(n1500) );
  NAND U4599 ( .A(n1501), .B(n1500), .Z(n1565) );
  XNOR U4600 ( .A(n1555), .B(n1565), .Z(n1531) );
  AND U4601 ( .A(n1502), .B(n1531), .Z(n1524) );
  OR U4602 ( .A(n1509), .B(n1506), .Z(n1508) );
  ANDN U4603 ( .B(n1509), .A(n1503), .Z(n1504) );
  XNOR U4604 ( .A(n1504), .B(n1514), .Z(n1505) );
  NAND U4605 ( .A(n1506), .B(n1505), .Z(n1507) );
  NAND U4606 ( .A(n1508), .B(n1507), .Z(n1528) );
  NAND U4607 ( .A(n1510), .B(n1514), .Z(n1516) );
  NAND U4608 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U4609 ( .A(n1512), .B(n1511), .Z(n1513) );
  NANDN U4610 ( .A(n1514), .B(n1513), .Z(n1515) );
  NAND U4611 ( .A(n1516), .B(n1515), .Z(n1572) );
  NAND U4612 ( .A(n1547), .B(n1517), .Z(n1518) );
  XNOR U4613 ( .A(n1524), .B(n1518), .Z(n1567) );
  XOR U4614 ( .A(n1555), .B(n1572), .Z(n1557) );
  AND U4615 ( .A(n1519), .B(n1557), .Z(n1542) );
  XNOR U4616 ( .A(n1567), .B(n1542), .Z(n1520) );
  XNOR U4617 ( .A(n1521), .B(n1520), .Z(n1575) );
  NAND U4618 ( .A(n1533), .B(n1522), .Z(n1523) );
  XNOR U4619 ( .A(n1524), .B(n1523), .Z(n1550) );
  AND U4620 ( .A(n1525), .B(n1535), .Z(n1566) );
  NANDN U4621 ( .A(n1526), .B(n1528), .Z(n1527) );
  XNOR U4622 ( .A(n1566), .B(n1527), .Z(n1554) );
  XNOR U4623 ( .A(n1550), .B(n1554), .Z(n1539) );
  XOR U4624 ( .A(n1575), .B(n1539), .Z(z[64]) );
  AND U4625 ( .A(n1529), .B(n1528), .Z(n1538) );
  AND U4626 ( .A(n1531), .B(n1530), .Z(n1549) );
  NAND U4627 ( .A(n1533), .B(n1532), .Z(n1534) );
  XNOR U4628 ( .A(n1549), .B(n1534), .Z(n1576) );
  AND U4629 ( .A(n1536), .B(n1535), .Z(n1543) );
  XNOR U4630 ( .A(n1576), .B(n1543), .Z(n1537) );
  XNOR U4631 ( .A(n1538), .B(n1537), .Z(n1563) );
  XNOR U4632 ( .A(n1563), .B(n1539), .Z(n1583) );
  AND U4633 ( .A(n1540), .B(n1565), .Z(n1545) );
  NANDN U4634 ( .A(n1572), .B(n1570), .Z(n1541) );
  XNOR U4635 ( .A(n1542), .B(n1541), .Z(n1553) );
  XNOR U4636 ( .A(n1543), .B(n1553), .Z(n1544) );
  XNOR U4637 ( .A(n1545), .B(n1544), .Z(n1552) );
  NAND U4638 ( .A(n1547), .B(n1546), .Z(n1548) );
  XNOR U4639 ( .A(n1549), .B(n1548), .Z(n1559) );
  XNOR U4640 ( .A(n1550), .B(n1559), .Z(n1551) );
  XNOR U4641 ( .A(n1552), .B(n1551), .Z(n1562) );
  XNOR U4642 ( .A(n1583), .B(n1562), .Z(z[65]) );
  XNOR U4643 ( .A(n1554), .B(n1553), .Z(z[66]) );
  NOR U4644 ( .A(n1556), .B(n1555), .Z(n1561) );
  AND U4645 ( .A(n1558), .B(n1557), .Z(n1574) );
  XNOR U4646 ( .A(n1559), .B(n1574), .Z(n1560) );
  XNOR U4647 ( .A(n1561), .B(n1560), .Z(n1582) );
  XOR U4648 ( .A(n1563), .B(n1562), .Z(n1564) );
  XNOR U4649 ( .A(n1582), .B(n1564), .Z(z[67]) );
  XOR U4650 ( .A(n1575), .B(z[66]), .Z(z[68]) );
  AND U4651 ( .A(x[64]), .B(n1565), .Z(n1569) );
  XNOR U4652 ( .A(n1567), .B(n1566), .Z(n1568) );
  XNOR U4653 ( .A(n1569), .B(n1568), .Z(n1584) );
  XOR U4654 ( .A(n1570), .B(x[65]), .Z(n1571) );
  NANDN U4655 ( .A(n1572), .B(n1571), .Z(n1573) );
  XNOR U4656 ( .A(n1574), .B(n1573), .Z(n1578) );
  XNOR U4657 ( .A(n1576), .B(n1575), .Z(n1577) );
  XNOR U4658 ( .A(n1578), .B(n1577), .Z(n1579) );
  XNOR U4659 ( .A(n1584), .B(n1579), .Z(z[69]) );
  XNOR U4660 ( .A(n1581), .B(n1580), .Z(z[6]) );
  XNOR U4661 ( .A(n1583), .B(n1582), .Z(z[70]) );
  XOR U4662 ( .A(n1584), .B(z[65]), .Z(z[71]) );
  XOR U4663 ( .A(x[75]), .B(x[73]), .Z(n1587) );
  XNOR U4664 ( .A(x[72]), .B(x[78]), .Z(n1586) );
  XOR U4665 ( .A(n1586), .B(x[74]), .Z(n1585) );
  XNOR U4666 ( .A(n1587), .B(n1585), .Z(n1622) );
  XNOR U4667 ( .A(x[77]), .B(n1586), .Z(n1695) );
  XOR U4668 ( .A(n1695), .B(x[76]), .Z(n1665) );
  IV U4669 ( .A(n1665), .Z(n1596) );
  XNOR U4670 ( .A(x[79]), .B(x[76]), .Z(n1590) );
  XNOR U4671 ( .A(n1587), .B(n1590), .Z(n1650) );
  NOR U4672 ( .A(n1596), .B(n1650), .Z(n1589) );
  XNOR U4673 ( .A(n1695), .B(x[79]), .Z(n1681) );
  XNOR U4674 ( .A(x[74]), .B(n1681), .Z(n1605) );
  XNOR U4675 ( .A(x[73]), .B(n1605), .Z(n1600) );
  AND U4676 ( .A(x[72]), .B(n1600), .Z(n1588) );
  XNOR U4677 ( .A(n1589), .B(n1588), .Z(n1593) );
  XNOR U4678 ( .A(n1622), .B(n1681), .Z(n1612) );
  IV U4679 ( .A(n1622), .Z(n1607) );
  XNOR U4680 ( .A(x[72]), .B(n1607), .Z(n1627) );
  IV U4681 ( .A(n1590), .Z(n1655) );
  AND U4682 ( .A(n1627), .B(n1655), .Z(n1595) );
  IV U4683 ( .A(n1695), .Z(n1614) );
  XNOR U4684 ( .A(n1622), .B(n1614), .Z(n1644) );
  XOR U4685 ( .A(n1644), .B(n1650), .Z(n1647) );
  XOR U4686 ( .A(x[74]), .B(x[76]), .Z(n1657) );
  NAND U4687 ( .A(n1647), .B(n1657), .Z(n1591) );
  XNOR U4688 ( .A(n1595), .B(n1591), .Z(n1616) );
  XNOR U4689 ( .A(n1612), .B(n1616), .Z(n1592) );
  XNOR U4690 ( .A(n1593), .B(n1592), .Z(n1639) );
  XOR U4691 ( .A(x[74]), .B(x[79]), .Z(n1671) );
  XNOR U4692 ( .A(x[72]), .B(n1650), .Z(n1651) );
  XNOR U4693 ( .A(n1695), .B(n1651), .Z(n1642) );
  NAND U4694 ( .A(n1671), .B(n1642), .Z(n1594) );
  XNOR U4695 ( .A(n1595), .B(n1594), .Z(n1608) );
  IV U4696 ( .A(n1600), .Z(n1654) );
  XNOR U4697 ( .A(n1654), .B(n1596), .Z(n1661) );
  AND U4698 ( .A(n1650), .B(n1661), .Z(n1598) );
  AND U4699 ( .A(x[72]), .B(n1665), .Z(n1597) );
  XNOR U4700 ( .A(n1598), .B(n1597), .Z(n1599) );
  NANDN U4701 ( .A(n1651), .B(n1599), .Z(n1603) );
  NAND U4702 ( .A(x[72]), .B(n1650), .Z(n1601) );
  OR U4703 ( .A(n1601), .B(n1600), .Z(n1602) );
  NAND U4704 ( .A(n1603), .B(n1602), .Z(n1604) );
  XNOR U4705 ( .A(n1605), .B(n1604), .Z(n1606) );
  XNOR U4706 ( .A(n1608), .B(n1606), .Z(n1628) );
  IV U4707 ( .A(n1628), .Z(n1635) );
  AND U4708 ( .A(n1681), .B(n1607), .Z(n1610) );
  XOR U4709 ( .A(x[73]), .B(x[79]), .Z(n1683) );
  AND U4710 ( .A(n1644), .B(n1683), .Z(n1613) );
  XNOR U4711 ( .A(n1613), .B(n1608), .Z(n1609) );
  XNOR U4712 ( .A(n1610), .B(n1609), .Z(n1634) );
  NANDN U4713 ( .A(n1635), .B(n1634), .Z(n1611) );
  NAND U4714 ( .A(n1639), .B(n1611), .Z(n1621) );
  XNOR U4715 ( .A(n1613), .B(n1612), .Z(n1618) );
  ANDN U4716 ( .B(n1614), .A(x[73]), .Z(n1615) );
  XNOR U4717 ( .A(n1616), .B(n1615), .Z(n1617) );
  XNOR U4718 ( .A(n1618), .B(n1617), .Z(n1631) );
  XOR U4719 ( .A(n1634), .B(n1631), .Z(n1619) );
  NAND U4720 ( .A(n1635), .B(n1619), .Z(n1620) );
  NAND U4721 ( .A(n1621), .B(n1620), .Z(n1680) );
  ANDN U4722 ( .B(n1622), .A(n1680), .Z(n1646) );
  IV U4723 ( .A(n1631), .Z(n1637) );
  XOR U4724 ( .A(n1639), .B(n1635), .Z(n1623) );
  NANDN U4725 ( .A(n1637), .B(n1623), .Z(n1626) );
  NANDN U4726 ( .A(n1635), .B(n1637), .Z(n1624) );
  NANDN U4727 ( .A(n1634), .B(n1624), .Z(n1625) );
  NAND U4728 ( .A(n1626), .B(n1625), .Z(n1690) );
  XNOR U4729 ( .A(n1680), .B(n1690), .Z(n1656) );
  AND U4730 ( .A(n1627), .B(n1656), .Z(n1649) );
  OR U4731 ( .A(n1634), .B(n1631), .Z(n1633) );
  ANDN U4732 ( .B(n1634), .A(n1628), .Z(n1629) );
  XNOR U4733 ( .A(n1629), .B(n1639), .Z(n1630) );
  NAND U4734 ( .A(n1631), .B(n1630), .Z(n1632) );
  NAND U4735 ( .A(n1633), .B(n1632), .Z(n1653) );
  NAND U4736 ( .A(n1635), .B(n1639), .Z(n1641) );
  NAND U4737 ( .A(n1635), .B(n1634), .Z(n1636) );
  XNOR U4738 ( .A(n1637), .B(n1636), .Z(n1638) );
  NANDN U4739 ( .A(n1639), .B(n1638), .Z(n1640) );
  NAND U4740 ( .A(n1641), .B(n1640), .Z(n1697) );
  NAND U4741 ( .A(n1672), .B(n1642), .Z(n1643) );
  XNOR U4742 ( .A(n1649), .B(n1643), .Z(n1692) );
  XOR U4743 ( .A(n1680), .B(n1697), .Z(n1682) );
  AND U4744 ( .A(n1644), .B(n1682), .Z(n1667) );
  XNOR U4745 ( .A(n1692), .B(n1667), .Z(n1645) );
  XNOR U4746 ( .A(n1646), .B(n1645), .Z(n1700) );
  NAND U4747 ( .A(n1658), .B(n1647), .Z(n1648) );
  XNOR U4748 ( .A(n1649), .B(n1648), .Z(n1675) );
  AND U4749 ( .A(n1650), .B(n1660), .Z(n1691) );
  NANDN U4750 ( .A(n1651), .B(n1653), .Z(n1652) );
  XNOR U4751 ( .A(n1691), .B(n1652), .Z(n1679) );
  XNOR U4752 ( .A(n1675), .B(n1679), .Z(n1664) );
  XOR U4753 ( .A(n1700), .B(n1664), .Z(z[72]) );
  AND U4754 ( .A(n1654), .B(n1653), .Z(n1663) );
  AND U4755 ( .A(n1656), .B(n1655), .Z(n1674) );
  NAND U4756 ( .A(n1658), .B(n1657), .Z(n1659) );
  XNOR U4757 ( .A(n1674), .B(n1659), .Z(n1701) );
  AND U4758 ( .A(n1661), .B(n1660), .Z(n1668) );
  XNOR U4759 ( .A(n1701), .B(n1668), .Z(n1662) );
  XNOR U4760 ( .A(n1663), .B(n1662), .Z(n1688) );
  XNOR U4761 ( .A(n1688), .B(n1664), .Z(n1706) );
  AND U4762 ( .A(n1665), .B(n1690), .Z(n1670) );
  NANDN U4763 ( .A(n1697), .B(n1695), .Z(n1666) );
  XNOR U4764 ( .A(n1667), .B(n1666), .Z(n1678) );
  XNOR U4765 ( .A(n1668), .B(n1678), .Z(n1669) );
  XNOR U4766 ( .A(n1670), .B(n1669), .Z(n1677) );
  NAND U4767 ( .A(n1672), .B(n1671), .Z(n1673) );
  XNOR U4768 ( .A(n1674), .B(n1673), .Z(n1684) );
  XNOR U4769 ( .A(n1675), .B(n1684), .Z(n1676) );
  XNOR U4770 ( .A(n1677), .B(n1676), .Z(n1687) );
  XNOR U4771 ( .A(n1706), .B(n1687), .Z(z[73]) );
  XNOR U4772 ( .A(n1679), .B(n1678), .Z(z[74]) );
  NOR U4773 ( .A(n1681), .B(n1680), .Z(n1686) );
  AND U4774 ( .A(n1683), .B(n1682), .Z(n1699) );
  XNOR U4775 ( .A(n1684), .B(n1699), .Z(n1685) );
  XNOR U4776 ( .A(n1686), .B(n1685), .Z(n1705) );
  XOR U4777 ( .A(n1688), .B(n1687), .Z(n1689) );
  XNOR U4778 ( .A(n1705), .B(n1689), .Z(z[75]) );
  XOR U4779 ( .A(n1700), .B(z[74]), .Z(z[76]) );
  AND U4780 ( .A(x[72]), .B(n1690), .Z(n1694) );
  XNOR U4781 ( .A(n1692), .B(n1691), .Z(n1693) );
  XNOR U4782 ( .A(n1694), .B(n1693), .Z(n1707) );
  XOR U4783 ( .A(n1695), .B(x[73]), .Z(n1696) );
  NANDN U4784 ( .A(n1697), .B(n1696), .Z(n1698) );
  XNOR U4785 ( .A(n1699), .B(n1698), .Z(n1703) );
  XNOR U4786 ( .A(n1701), .B(n1700), .Z(n1702) );
  XNOR U4787 ( .A(n1703), .B(n1702), .Z(n1704) );
  XNOR U4788 ( .A(n1707), .B(n1704), .Z(z[77]) );
  XNOR U4789 ( .A(n1706), .B(n1705), .Z(z[78]) );
  XOR U4790 ( .A(n1707), .B(z[73]), .Z(z[79]) );
  XOR U4791 ( .A(n1708), .B(z[1]), .Z(z[7]) );
  XOR U4792 ( .A(x[83]), .B(x[81]), .Z(n1711) );
  XNOR U4793 ( .A(x[80]), .B(x[86]), .Z(n1710) );
  XOR U4794 ( .A(n1710), .B(x[82]), .Z(n1709) );
  XNOR U4795 ( .A(n1711), .B(n1709), .Z(n1746) );
  XNOR U4796 ( .A(x[85]), .B(n1710), .Z(n1819) );
  XOR U4797 ( .A(n1819), .B(x[84]), .Z(n1789) );
  IV U4798 ( .A(n1789), .Z(n1720) );
  XNOR U4799 ( .A(x[87]), .B(x[84]), .Z(n1714) );
  XNOR U4800 ( .A(n1711), .B(n1714), .Z(n1774) );
  NOR U4801 ( .A(n1720), .B(n1774), .Z(n1713) );
  XNOR U4802 ( .A(n1819), .B(x[87]), .Z(n1805) );
  XNOR U4803 ( .A(x[82]), .B(n1805), .Z(n1729) );
  XNOR U4804 ( .A(x[81]), .B(n1729), .Z(n1724) );
  AND U4805 ( .A(x[80]), .B(n1724), .Z(n1712) );
  XNOR U4806 ( .A(n1713), .B(n1712), .Z(n1717) );
  XNOR U4807 ( .A(n1746), .B(n1805), .Z(n1736) );
  IV U4808 ( .A(n1746), .Z(n1731) );
  XNOR U4809 ( .A(x[80]), .B(n1731), .Z(n1751) );
  IV U4810 ( .A(n1714), .Z(n1779) );
  AND U4811 ( .A(n1751), .B(n1779), .Z(n1719) );
  IV U4812 ( .A(n1819), .Z(n1738) );
  XNOR U4813 ( .A(n1746), .B(n1738), .Z(n1768) );
  XOR U4814 ( .A(n1768), .B(n1774), .Z(n1771) );
  XOR U4815 ( .A(x[82]), .B(x[84]), .Z(n1781) );
  NAND U4816 ( .A(n1771), .B(n1781), .Z(n1715) );
  XNOR U4817 ( .A(n1719), .B(n1715), .Z(n1740) );
  XNOR U4818 ( .A(n1736), .B(n1740), .Z(n1716) );
  XNOR U4819 ( .A(n1717), .B(n1716), .Z(n1763) );
  XOR U4820 ( .A(x[82]), .B(x[87]), .Z(n1795) );
  XNOR U4821 ( .A(x[80]), .B(n1774), .Z(n1775) );
  XNOR U4822 ( .A(n1819), .B(n1775), .Z(n1766) );
  NAND U4823 ( .A(n1795), .B(n1766), .Z(n1718) );
  XNOR U4824 ( .A(n1719), .B(n1718), .Z(n1732) );
  IV U4825 ( .A(n1724), .Z(n1778) );
  XNOR U4826 ( .A(n1778), .B(n1720), .Z(n1785) );
  AND U4827 ( .A(n1774), .B(n1785), .Z(n1722) );
  AND U4828 ( .A(x[80]), .B(n1789), .Z(n1721) );
  XNOR U4829 ( .A(n1722), .B(n1721), .Z(n1723) );
  NANDN U4830 ( .A(n1775), .B(n1723), .Z(n1727) );
  NAND U4831 ( .A(x[80]), .B(n1774), .Z(n1725) );
  OR U4832 ( .A(n1725), .B(n1724), .Z(n1726) );
  NAND U4833 ( .A(n1727), .B(n1726), .Z(n1728) );
  XNOR U4834 ( .A(n1729), .B(n1728), .Z(n1730) );
  XNOR U4835 ( .A(n1732), .B(n1730), .Z(n1752) );
  IV U4836 ( .A(n1752), .Z(n1759) );
  AND U4837 ( .A(n1805), .B(n1731), .Z(n1734) );
  XOR U4838 ( .A(x[81]), .B(x[87]), .Z(n1807) );
  AND U4839 ( .A(n1768), .B(n1807), .Z(n1737) );
  XNOR U4840 ( .A(n1737), .B(n1732), .Z(n1733) );
  XNOR U4841 ( .A(n1734), .B(n1733), .Z(n1758) );
  NANDN U4842 ( .A(n1759), .B(n1758), .Z(n1735) );
  NAND U4843 ( .A(n1763), .B(n1735), .Z(n1745) );
  XNOR U4844 ( .A(n1737), .B(n1736), .Z(n1742) );
  ANDN U4845 ( .B(n1738), .A(x[81]), .Z(n1739) );
  XNOR U4846 ( .A(n1740), .B(n1739), .Z(n1741) );
  XNOR U4847 ( .A(n1742), .B(n1741), .Z(n1755) );
  XOR U4848 ( .A(n1758), .B(n1755), .Z(n1743) );
  NAND U4849 ( .A(n1759), .B(n1743), .Z(n1744) );
  NAND U4850 ( .A(n1745), .B(n1744), .Z(n1804) );
  ANDN U4851 ( .B(n1746), .A(n1804), .Z(n1770) );
  IV U4852 ( .A(n1755), .Z(n1761) );
  XOR U4853 ( .A(n1763), .B(n1759), .Z(n1747) );
  NANDN U4854 ( .A(n1761), .B(n1747), .Z(n1750) );
  NANDN U4855 ( .A(n1759), .B(n1761), .Z(n1748) );
  NANDN U4856 ( .A(n1758), .B(n1748), .Z(n1749) );
  NAND U4857 ( .A(n1750), .B(n1749), .Z(n1814) );
  XNOR U4858 ( .A(n1804), .B(n1814), .Z(n1780) );
  AND U4859 ( .A(n1751), .B(n1780), .Z(n1773) );
  OR U4860 ( .A(n1758), .B(n1755), .Z(n1757) );
  ANDN U4861 ( .B(n1758), .A(n1752), .Z(n1753) );
  XNOR U4862 ( .A(n1753), .B(n1763), .Z(n1754) );
  NAND U4863 ( .A(n1755), .B(n1754), .Z(n1756) );
  NAND U4864 ( .A(n1757), .B(n1756), .Z(n1777) );
  NAND U4865 ( .A(n1759), .B(n1763), .Z(n1765) );
  NAND U4866 ( .A(n1759), .B(n1758), .Z(n1760) );
  XNOR U4867 ( .A(n1761), .B(n1760), .Z(n1762) );
  NANDN U4868 ( .A(n1763), .B(n1762), .Z(n1764) );
  NAND U4869 ( .A(n1765), .B(n1764), .Z(n1821) );
  NAND U4870 ( .A(n1796), .B(n1766), .Z(n1767) );
  XNOR U4871 ( .A(n1773), .B(n1767), .Z(n1816) );
  XOR U4872 ( .A(n1804), .B(n1821), .Z(n1806) );
  AND U4873 ( .A(n1768), .B(n1806), .Z(n1791) );
  XNOR U4874 ( .A(n1816), .B(n1791), .Z(n1769) );
  XNOR U4875 ( .A(n1770), .B(n1769), .Z(n1824) );
  NAND U4876 ( .A(n1782), .B(n1771), .Z(n1772) );
  XNOR U4877 ( .A(n1773), .B(n1772), .Z(n1799) );
  AND U4878 ( .A(n1774), .B(n1784), .Z(n1815) );
  NANDN U4879 ( .A(n1775), .B(n1777), .Z(n1776) );
  XNOR U4880 ( .A(n1815), .B(n1776), .Z(n1803) );
  XNOR U4881 ( .A(n1799), .B(n1803), .Z(n1788) );
  XOR U4882 ( .A(n1824), .B(n1788), .Z(z[80]) );
  AND U4883 ( .A(n1778), .B(n1777), .Z(n1787) );
  AND U4884 ( .A(n1780), .B(n1779), .Z(n1798) );
  NAND U4885 ( .A(n1782), .B(n1781), .Z(n1783) );
  XNOR U4886 ( .A(n1798), .B(n1783), .Z(n1825) );
  AND U4887 ( .A(n1785), .B(n1784), .Z(n1792) );
  XNOR U4888 ( .A(n1825), .B(n1792), .Z(n1786) );
  XNOR U4889 ( .A(n1787), .B(n1786), .Z(n1812) );
  XNOR U4890 ( .A(n1812), .B(n1788), .Z(n1830) );
  AND U4891 ( .A(n1789), .B(n1814), .Z(n1794) );
  NANDN U4892 ( .A(n1821), .B(n1819), .Z(n1790) );
  XNOR U4893 ( .A(n1791), .B(n1790), .Z(n1802) );
  XNOR U4894 ( .A(n1792), .B(n1802), .Z(n1793) );
  XNOR U4895 ( .A(n1794), .B(n1793), .Z(n1801) );
  NAND U4896 ( .A(n1796), .B(n1795), .Z(n1797) );
  XNOR U4897 ( .A(n1798), .B(n1797), .Z(n1808) );
  XNOR U4898 ( .A(n1799), .B(n1808), .Z(n1800) );
  XNOR U4899 ( .A(n1801), .B(n1800), .Z(n1811) );
  XNOR U4900 ( .A(n1830), .B(n1811), .Z(z[81]) );
  XNOR U4901 ( .A(n1803), .B(n1802), .Z(z[82]) );
  NOR U4902 ( .A(n1805), .B(n1804), .Z(n1810) );
  AND U4903 ( .A(n1807), .B(n1806), .Z(n1823) );
  XNOR U4904 ( .A(n1808), .B(n1823), .Z(n1809) );
  XNOR U4905 ( .A(n1810), .B(n1809), .Z(n1829) );
  XOR U4906 ( .A(n1812), .B(n1811), .Z(n1813) );
  XNOR U4907 ( .A(n1829), .B(n1813), .Z(z[83]) );
  XOR U4908 ( .A(n1824), .B(z[82]), .Z(z[84]) );
  AND U4909 ( .A(x[80]), .B(n1814), .Z(n1818) );
  XNOR U4910 ( .A(n1816), .B(n1815), .Z(n1817) );
  XNOR U4911 ( .A(n1818), .B(n1817), .Z(n1831) );
  XOR U4912 ( .A(n1819), .B(x[81]), .Z(n1820) );
  NANDN U4913 ( .A(n1821), .B(n1820), .Z(n1822) );
  XNOR U4914 ( .A(n1823), .B(n1822), .Z(n1827) );
  XNOR U4915 ( .A(n1825), .B(n1824), .Z(n1826) );
  XNOR U4916 ( .A(n1827), .B(n1826), .Z(n1828) );
  XNOR U4917 ( .A(n1831), .B(n1828), .Z(z[85]) );
  XNOR U4918 ( .A(n1830), .B(n1829), .Z(z[86]) );
  XOR U4919 ( .A(n1831), .B(z[81]), .Z(z[87]) );
  XOR U4920 ( .A(x[91]), .B(x[89]), .Z(n1834) );
  XNOR U4921 ( .A(x[88]), .B(x[94]), .Z(n1833) );
  XOR U4922 ( .A(n1833), .B(x[90]), .Z(n1832) );
  XNOR U4923 ( .A(n1834), .B(n1832), .Z(n1869) );
  XNOR U4924 ( .A(x[93]), .B(n1833), .Z(n1944) );
  XOR U4925 ( .A(n1944), .B(x[92]), .Z(n1912) );
  IV U4926 ( .A(n1912), .Z(n1843) );
  XNOR U4927 ( .A(x[95]), .B(x[92]), .Z(n1837) );
  XNOR U4928 ( .A(n1834), .B(n1837), .Z(n1897) );
  NOR U4929 ( .A(n1843), .B(n1897), .Z(n1836) );
  XNOR U4930 ( .A(n1944), .B(x[95]), .Z(n1930) );
  XNOR U4931 ( .A(x[90]), .B(n1930), .Z(n1852) );
  XNOR U4932 ( .A(x[89]), .B(n1852), .Z(n1847) );
  AND U4933 ( .A(x[88]), .B(n1847), .Z(n1835) );
  XNOR U4934 ( .A(n1836), .B(n1835), .Z(n1840) );
  XNOR U4935 ( .A(n1869), .B(n1930), .Z(n1859) );
  IV U4936 ( .A(n1869), .Z(n1854) );
  XNOR U4937 ( .A(x[88]), .B(n1854), .Z(n1874) );
  IV U4938 ( .A(n1837), .Z(n1902) );
  AND U4939 ( .A(n1874), .B(n1902), .Z(n1842) );
  IV U4940 ( .A(n1944), .Z(n1861) );
  XNOR U4941 ( .A(n1869), .B(n1861), .Z(n1891) );
  XOR U4942 ( .A(n1891), .B(n1897), .Z(n1894) );
  XOR U4943 ( .A(x[90]), .B(x[92]), .Z(n1904) );
  NAND U4944 ( .A(n1894), .B(n1904), .Z(n1838) );
  XNOR U4945 ( .A(n1842), .B(n1838), .Z(n1863) );
  XNOR U4946 ( .A(n1859), .B(n1863), .Z(n1839) );
  XNOR U4947 ( .A(n1840), .B(n1839), .Z(n1886) );
  XOR U4948 ( .A(x[90]), .B(x[95]), .Z(n1918) );
  XNOR U4949 ( .A(x[88]), .B(n1897), .Z(n1898) );
  XNOR U4950 ( .A(n1944), .B(n1898), .Z(n1889) );
  NAND U4951 ( .A(n1918), .B(n1889), .Z(n1841) );
  XNOR U4952 ( .A(n1842), .B(n1841), .Z(n1855) );
  IV U4953 ( .A(n1847), .Z(n1901) );
  XNOR U4954 ( .A(n1901), .B(n1843), .Z(n1908) );
  AND U4955 ( .A(n1897), .B(n1908), .Z(n1845) );
  AND U4956 ( .A(x[88]), .B(n1912), .Z(n1844) );
  XNOR U4957 ( .A(n1845), .B(n1844), .Z(n1846) );
  NANDN U4958 ( .A(n1898), .B(n1846), .Z(n1850) );
  NAND U4959 ( .A(x[88]), .B(n1897), .Z(n1848) );
  OR U4960 ( .A(n1848), .B(n1847), .Z(n1849) );
  NAND U4961 ( .A(n1850), .B(n1849), .Z(n1851) );
  XNOR U4962 ( .A(n1852), .B(n1851), .Z(n1853) );
  XNOR U4963 ( .A(n1855), .B(n1853), .Z(n1875) );
  IV U4964 ( .A(n1875), .Z(n1882) );
  AND U4965 ( .A(n1930), .B(n1854), .Z(n1857) );
  XOR U4966 ( .A(x[89]), .B(x[95]), .Z(n1932) );
  AND U4967 ( .A(n1891), .B(n1932), .Z(n1860) );
  XNOR U4968 ( .A(n1860), .B(n1855), .Z(n1856) );
  XNOR U4969 ( .A(n1857), .B(n1856), .Z(n1881) );
  NANDN U4970 ( .A(n1882), .B(n1881), .Z(n1858) );
  NAND U4971 ( .A(n1886), .B(n1858), .Z(n1868) );
  XNOR U4972 ( .A(n1860), .B(n1859), .Z(n1865) );
  ANDN U4973 ( .B(n1861), .A(x[89]), .Z(n1862) );
  XNOR U4974 ( .A(n1863), .B(n1862), .Z(n1864) );
  XNOR U4975 ( .A(n1865), .B(n1864), .Z(n1878) );
  XOR U4976 ( .A(n1881), .B(n1878), .Z(n1866) );
  NAND U4977 ( .A(n1882), .B(n1866), .Z(n1867) );
  NAND U4978 ( .A(n1868), .B(n1867), .Z(n1929) );
  ANDN U4979 ( .B(n1869), .A(n1929), .Z(n1893) );
  IV U4980 ( .A(n1878), .Z(n1884) );
  XOR U4981 ( .A(n1886), .B(n1882), .Z(n1870) );
  NANDN U4982 ( .A(n1884), .B(n1870), .Z(n1873) );
  NANDN U4983 ( .A(n1882), .B(n1884), .Z(n1871) );
  NANDN U4984 ( .A(n1881), .B(n1871), .Z(n1872) );
  NAND U4985 ( .A(n1873), .B(n1872), .Z(n1939) );
  XNOR U4986 ( .A(n1929), .B(n1939), .Z(n1903) );
  AND U4987 ( .A(n1874), .B(n1903), .Z(n1896) );
  OR U4988 ( .A(n1881), .B(n1878), .Z(n1880) );
  ANDN U4989 ( .B(n1881), .A(n1875), .Z(n1876) );
  XNOR U4990 ( .A(n1876), .B(n1886), .Z(n1877) );
  NAND U4991 ( .A(n1878), .B(n1877), .Z(n1879) );
  NAND U4992 ( .A(n1880), .B(n1879), .Z(n1900) );
  NAND U4993 ( .A(n1882), .B(n1886), .Z(n1888) );
  NAND U4994 ( .A(n1882), .B(n1881), .Z(n1883) );
  XNOR U4995 ( .A(n1884), .B(n1883), .Z(n1885) );
  NANDN U4996 ( .A(n1886), .B(n1885), .Z(n1887) );
  NAND U4997 ( .A(n1888), .B(n1887), .Z(n1946) );
  NAND U4998 ( .A(n1919), .B(n1889), .Z(n1890) );
  XNOR U4999 ( .A(n1896), .B(n1890), .Z(n1941) );
  XOR U5000 ( .A(n1929), .B(n1946), .Z(n1931) );
  AND U5001 ( .A(n1891), .B(n1931), .Z(n1914) );
  XNOR U5002 ( .A(n1941), .B(n1914), .Z(n1892) );
  XNOR U5003 ( .A(n1893), .B(n1892), .Z(n1949) );
  NAND U5004 ( .A(n1905), .B(n1894), .Z(n1895) );
  XNOR U5005 ( .A(n1896), .B(n1895), .Z(n1922) );
  AND U5006 ( .A(n1897), .B(n1907), .Z(n1940) );
  NANDN U5007 ( .A(n1898), .B(n1900), .Z(n1899) );
  XNOR U5008 ( .A(n1940), .B(n1899), .Z(n1928) );
  XNOR U5009 ( .A(n1922), .B(n1928), .Z(n1911) );
  XOR U5010 ( .A(n1949), .B(n1911), .Z(z[88]) );
  AND U5011 ( .A(n1901), .B(n1900), .Z(n1910) );
  AND U5012 ( .A(n1903), .B(n1902), .Z(n1921) );
  NAND U5013 ( .A(n1905), .B(n1904), .Z(n1906) );
  XNOR U5014 ( .A(n1921), .B(n1906), .Z(n1950) );
  AND U5015 ( .A(n1908), .B(n1907), .Z(n1915) );
  XNOR U5016 ( .A(n1950), .B(n1915), .Z(n1909) );
  XNOR U5017 ( .A(n1910), .B(n1909), .Z(n1937) );
  XNOR U5018 ( .A(n1937), .B(n1911), .Z(n1955) );
  AND U5019 ( .A(n1912), .B(n1939), .Z(n1917) );
  NANDN U5020 ( .A(n1946), .B(n1944), .Z(n1913) );
  XNOR U5021 ( .A(n1914), .B(n1913), .Z(n1927) );
  XNOR U5022 ( .A(n1915), .B(n1927), .Z(n1916) );
  XNOR U5023 ( .A(n1917), .B(n1916), .Z(n1924) );
  NAND U5024 ( .A(n1919), .B(n1918), .Z(n1920) );
  XNOR U5025 ( .A(n1921), .B(n1920), .Z(n1933) );
  XNOR U5026 ( .A(n1922), .B(n1933), .Z(n1923) );
  XNOR U5027 ( .A(n1924), .B(n1923), .Z(n1936) );
  XNOR U5028 ( .A(n1955), .B(n1936), .Z(z[89]) );
  XOR U5029 ( .A(n1926), .B(n1925), .Z(z[8]) );
  XNOR U5030 ( .A(n1928), .B(n1927), .Z(z[90]) );
  NOR U5031 ( .A(n1930), .B(n1929), .Z(n1935) );
  AND U5032 ( .A(n1932), .B(n1931), .Z(n1948) );
  XNOR U5033 ( .A(n1933), .B(n1948), .Z(n1934) );
  XNOR U5034 ( .A(n1935), .B(n1934), .Z(n1954) );
  XOR U5035 ( .A(n1937), .B(n1936), .Z(n1938) );
  XNOR U5036 ( .A(n1954), .B(n1938), .Z(z[91]) );
  XOR U5037 ( .A(n1949), .B(z[90]), .Z(z[92]) );
  AND U5038 ( .A(x[88]), .B(n1939), .Z(n1943) );
  XNOR U5039 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U5040 ( .A(n1943), .B(n1942), .Z(n1956) );
  XOR U5041 ( .A(n1944), .B(x[89]), .Z(n1945) );
  NANDN U5042 ( .A(n1946), .B(n1945), .Z(n1947) );
  XNOR U5043 ( .A(n1948), .B(n1947), .Z(n1952) );
  XNOR U5044 ( .A(n1950), .B(n1949), .Z(n1951) );
  XNOR U5045 ( .A(n1952), .B(n1951), .Z(n1953) );
  XNOR U5046 ( .A(n1956), .B(n1953), .Z(z[93]) );
  XNOR U5047 ( .A(n1955), .B(n1954), .Z(z[94]) );
  XOR U5048 ( .A(n1956), .B(z[89]), .Z(z[95]) );
  XOR U5049 ( .A(n1958), .B(n1957), .Z(z[96]) );
  XOR U5050 ( .A(n1960), .B(n1959), .Z(n1961) );
  XNOR U5051 ( .A(n1962), .B(n1961), .Z(z[99]) );
endmodule


module aes_10 ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [127:0] key;
  output [127:0] out;
  input clk, rst;
  wire   init, \w0[0][127] , \w0[0][126] , \w0[0][125] , \w0[0][124] ,
         \w0[0][123] , \w0[0][122] , \w0[0][121] , \w0[0][120] , \w0[0][119] ,
         \w0[0][118] , \w0[0][117] , \w0[0][116] , \w0[0][115] , \w0[0][114] ,
         \w0[0][113] , \w0[0][112] , \w0[0][111] , \w0[0][110] , \w0[0][109] ,
         \w0[0][108] , \w0[0][107] , \w0[0][106] , \w0[0][105] , \w0[0][104] ,
         \w0[0][103] , \w0[0][102] , \w0[0][101] , \w0[0][100] , \w0[0][99] ,
         \w0[0][98] , \w0[0][97] , \w0[0][96] , \w0[0][95] , \w0[0][94] ,
         \w0[0][93] , \w0[0][92] , \w0[0][91] , \w0[0][90] , \w0[0][89] ,
         \w0[0][88] , \w0[0][87] , \w0[0][86] , \w0[0][85] , \w0[0][84] ,
         \w0[0][83] , \w0[0][82] , \w0[0][81] , \w0[0][80] , \w0[0][79] ,
         \w0[0][78] , \w0[0][77] , \w0[0][76] , \w0[0][75] , \w0[0][74] ,
         \w0[0][73] , \w0[0][72] , \w0[0][71] , \w0[0][70] , \w0[0][69] ,
         \w0[0][68] , \w0[0][67] , \w0[0][66] , \w0[0][65] , \w0[0][64] ,
         \w0[0][63] , \w0[0][62] , \w0[0][61] , \w0[0][60] , \w0[0][59] ,
         \w0[0][58] , \w0[0][57] , \w0[0][56] , \w0[0][55] , \w0[0][54] ,
         \w0[0][53] , \w0[0][52] , \w0[0][51] , \w0[0][50] , \w0[0][49] ,
         \w0[0][48] , \w0[0][47] , \w0[0][46] , \w0[0][45] , \w0[0][44] ,
         \w0[0][43] , \w0[0][42] , \w0[0][41] , \w0[0][40] , \w0[0][39] ,
         \w0[0][38] , \w0[0][37] , \w0[0][36] , \w0[0][35] , \w0[0][34] ,
         \w0[0][33] , \w0[0][32] , \w0[0][31] , \w0[0][30] , \w0[0][29] ,
         \w0[0][28] , \w0[0][27] , \w0[0][26] , \w0[0][25] , \w0[0][24] ,
         \w0[0][23] , \w0[0][22] , \w0[0][21] , \w0[0][20] , \w0[0][19] ,
         \w0[0][18] , \w0[0][17] , \w0[0][16] , \w0[0][15] , \w0[0][14] ,
         \w0[0][13] , \w0[0][12] , \w0[0][11] , \w0[0][10] , \w0[0][9] ,
         \w0[0][8] , \w0[0][7] , \w0[0][6] , \w0[0][5] , \w0[0][4] ,
         \w0[0][3] , \w0[0][2] , \w0[0][1] , \w0[0][0] , \w1[0][127] ,
         \w1[0][126] , \w1[0][125] , \w1[0][124] , \w1[0][123] , \w1[0][122] ,
         \w1[0][121] , \w1[0][120] , \w1[0][119] , \w1[0][118] , \w1[0][117] ,
         \w1[0][116] , \w1[0][115] , \w1[0][114] , \w1[0][113] , \w1[0][112] ,
         \w1[0][111] , \w1[0][110] , \w1[0][109] , \w1[0][108] , \w1[0][107] ,
         \w1[0][106] , \w1[0][105] , \w1[0][104] , \w1[0][103] , \w1[0][102] ,
         \w1[0][101] , \w1[0][100] , \w1[0][99] , \w1[0][98] , \w1[0][97] ,
         \w1[0][96] , \w1[0][95] , \w1[0][94] , \w1[0][93] , \w1[0][92] ,
         \w1[0][91] , \w1[0][90] , \w1[0][89] , \w1[0][88] , \w1[0][87] ,
         \w1[0][86] , \w1[0][85] , \w1[0][84] , \w1[0][83] , \w1[0][82] ,
         \w1[0][81] , \w1[0][80] , \w1[0][79] , \w1[0][78] , \w1[0][77] ,
         \w1[0][76] , \w1[0][75] , \w1[0][74] , \w1[0][73] , \w1[0][72] ,
         \w1[0][71] , \w1[0][70] , \w1[0][69] , \w1[0][68] , \w1[0][67] ,
         \w1[0][66] , \w1[0][65] , \w1[0][64] , \w1[0][63] , \w1[0][62] ,
         \w1[0][61] , \w1[0][60] , \w1[0][59] , \w1[0][58] , \w1[0][57] ,
         \w1[0][56] , \w1[0][55] , \w1[0][54] , \w1[0][53] , \w1[0][52] ,
         \w1[0][51] , \w1[0][50] , \w1[0][49] , \w1[0][48] , \w1[0][47] ,
         \w1[0][46] , \w1[0][45] , \w1[0][44] , \w1[0][43] , \w1[0][42] ,
         \w1[0][41] , \w1[0][40] , \w1[0][39] , \w1[0][38] , \w1[0][37] ,
         \w1[0][36] , \w1[0][35] , \w1[0][34] , \w1[0][33] , \w1[0][32] ,
         \w1[0][31] , \w1[0][30] , \w1[0][29] , \w1[0][28] , \w1[0][27] ,
         \w1[0][26] , \w1[0][25] , \w1[0][24] , \w1[0][23] , \w1[0][22] ,
         \w1[0][21] , \w1[0][20] , \w1[0][19] , \w1[0][18] , \w1[0][17] ,
         \w1[0][16] , \w1[0][15] , \w1[0][14] , \w1[0][13] , \w1[0][12] ,
         \w1[0][11] , \w1[0][10] , \w1[0][9] , \w1[0][8] , \w1[0][7] ,
         \w1[0][6] , \w1[0][5] , \w1[0][4] , \w1[0][3] , \w1[0][2] ,
         \w1[0][1] , \w1[0][0] , \w3[0][127] , \w3[0][126] , \w3[0][125] ,
         \w3[0][124] , \w3[0][123] , \w3[0][122] , \w3[0][121] , \w3[0][120] ,
         \w3[0][119] , \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] ,
         \w3[0][114] , \w3[0][113] , \w3[0][112] , \w3[0][111] , \w3[0][110] ,
         \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , \w3[0][105] ,
         \w3[0][104] , \w3[0][103] , \w3[0][102] , \w3[0][101] , \w3[0][100] ,
         \w3[0][99] , \w3[0][98] , \w3[0][97] , \w3[0][96] , \w3[0][95] ,
         \w3[0][94] , \w3[0][93] , \w3[0][92] , \w3[0][91] , \w3[0][90] ,
         \w3[0][89] , \w3[0][88] , \w3[0][87] , \w3[0][86] , \w3[0][85] ,
         \w3[0][84] , \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] ,
         \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , \w3[0][75] ,
         \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][71] , \w3[0][70] ,
         \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] ,
         \w3[0][64] , \w3[0][63] , \w3[0][62] , \w3[0][61] , \w3[0][60] ,
         \w3[0][59] , \w3[0][58] , \w3[0][57] , \w3[0][56] , \w3[0][55] ,
         \w3[0][54] , \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] ,
         \w3[0][49] , \w3[0][48] , \w3[0][47] , \w3[0][46] , \w3[0][45] ,
         \w3[0][44] , \w3[0][43] , \w3[0][42] , \w3[0][41] , \w3[0][40] ,
         \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] ,
         \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][31] , \w3[0][30] ,
         \w3[0][29] , \w3[0][28] , \w3[0][27] , \w3[0][26] , \w3[0][25] ,
         \w3[0][24] , \w3[0][23] , \w3[0][22] , \w3[0][21] , \w3[0][20] ,
         \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , \w3[0][15] ,
         \w3[0][14] , \w3[0][13] , \w3[0][12] , \w3[0][11] , \w3[0][10] ,
         \w3[0][9] , \w3[0][8] , \w3[0][7] , \w3[0][6] , \w3[0][5] ,
         \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512;
  wire   [127:0] state;

  SubBytes \SUBBYTES[0].a  ( .x({\w1[0][127] , \w1[0][126] , \w1[0][125] , 
        \w1[0][124] , \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] , 
        \w1[0][119] , \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] , 
        \w1[0][114] , \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] , 
        \w1[0][109] , \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] , 
        \w1[0][104] , \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] , 
        \w1[0][99] , \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] , 
        \w1[0][94] , \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] , 
        \w1[0][89] , \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] , 
        \w1[0][84] , \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] , 
        \w1[0][79] , \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] , 
        \w1[0][74] , \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] , 
        \w1[0][69] , \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] , 
        \w1[0][64] , \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] , 
        \w1[0][59] , \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] , 
        \w1[0][54] , \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] , 
        \w1[0][49] , \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] , 
        \w1[0][44] , \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] , 
        \w1[0][39] , \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] , 
        \w1[0][34] , \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] , 
        \w1[0][29] , \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] , 
        \w1[0][24] , \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] , 
        \w1[0][19] , \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] , 
        \w1[0][14] , \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] , 
        \w1[0][9] , \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] , \w1[0][4] , 
        \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] }), .z({\w3[0][127] , 
        \w3[0][126] , \w3[0][125] , \w3[0][124] , \w3[0][123] , \w3[0][122] , 
        \w3[0][121] , \w3[0][120] , \w3[0][23] , \w3[0][22] , \w3[0][21] , 
        \w3[0][20] , \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , 
        \w3[0][47] , \w3[0][46] , \w3[0][45] , \w3[0][44] , \w3[0][43] , 
        \w3[0][42] , \w3[0][41] , \w3[0][40] , \w3[0][71] , \w3[0][70] , 
        \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] , 
        \w3[0][64] , \w3[0][95] , \w3[0][94] , \w3[0][93] , \w3[0][92] , 
        \w3[0][91] , \w3[0][90] , \w3[0][89] , \w3[0][88] , \w3[0][119] , 
        \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] , \w3[0][114] , 
        \w3[0][113] , \w3[0][112] , \w3[0][15] , \w3[0][14] , \w3[0][13] , 
        \w3[0][12] , \w3[0][11] , \w3[0][10] , \w3[0][9] , \w3[0][8] , 
        \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] , 
        \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][63] , \w3[0][62] , 
        \w3[0][61] , \w3[0][60] , \w3[0][59] , \w3[0][58] , \w3[0][57] , 
        \w3[0][56] , \w3[0][87] , \w3[0][86] , \w3[0][85] , \w3[0][84] , 
        \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] , \w3[0][111] , 
        \w3[0][110] , \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , 
        \w3[0][105] , \w3[0][104] , \w3[0][7] , \w3[0][6] , \w3[0][5] , 
        \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , 
        \w3[0][31] , \w3[0][30] , \w3[0][29] , \w3[0][28] , \w3[0][27] , 
        \w3[0][26] , \w3[0][25] , \w3[0][24] , \w3[0][55] , \w3[0][54] , 
        \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] , \w3[0][49] , 
        \w3[0][48] , \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , 
        \w3[0][75] , \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][103] , 
        \w3[0][102] , \w3[0][101] , \w3[0][100] , \w3[0][99] , \w3[0][98] , 
        \w3[0][97] , \w3[0][96] }) );
  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \state_reg[127]  ( .D(\w0[0][127] ), .CLK(clk), .RST(rst), .Q(state[127]) );
  DFF \state_reg[126]  ( .D(\w0[0][126] ), .CLK(clk), .RST(rst), .Q(state[126]) );
  DFF \state_reg[125]  ( .D(\w0[0][125] ), .CLK(clk), .RST(rst), .Q(state[125]) );
  DFF \state_reg[124]  ( .D(\w0[0][124] ), .CLK(clk), .RST(rst), .Q(state[124]) );
  DFF \state_reg[123]  ( .D(\w0[0][123] ), .CLK(clk), .RST(rst), .Q(state[123]) );
  DFF \state_reg[122]  ( .D(\w0[0][122] ), .CLK(clk), .RST(rst), .Q(state[122]) );
  DFF \state_reg[121]  ( .D(\w0[0][121] ), .CLK(clk), .RST(rst), .Q(state[121]) );
  DFF \state_reg[120]  ( .D(\w0[0][120] ), .CLK(clk), .RST(rst), .Q(state[120]) );
  DFF \state_reg[119]  ( .D(\w0[0][119] ), .CLK(clk), .RST(rst), .Q(state[119]) );
  DFF \state_reg[118]  ( .D(\w0[0][118] ), .CLK(clk), .RST(rst), .Q(state[118]) );
  DFF \state_reg[117]  ( .D(\w0[0][117] ), .CLK(clk), .RST(rst), .Q(state[117]) );
  DFF \state_reg[116]  ( .D(\w0[0][116] ), .CLK(clk), .RST(rst), .Q(state[116]) );
  DFF \state_reg[115]  ( .D(\w0[0][115] ), .CLK(clk), .RST(rst), .Q(state[115]) );
  DFF \state_reg[114]  ( .D(\w0[0][114] ), .CLK(clk), .RST(rst), .Q(state[114]) );
  DFF \state_reg[113]  ( .D(\w0[0][113] ), .CLK(clk), .RST(rst), .Q(state[113]) );
  DFF \state_reg[112]  ( .D(\w0[0][112] ), .CLK(clk), .RST(rst), .Q(state[112]) );
  DFF \state_reg[111]  ( .D(\w0[0][111] ), .CLK(clk), .RST(rst), .Q(state[111]) );
  DFF \state_reg[110]  ( .D(\w0[0][110] ), .CLK(clk), .RST(rst), .Q(state[110]) );
  DFF \state_reg[109]  ( .D(\w0[0][109] ), .CLK(clk), .RST(rst), .Q(state[109]) );
  DFF \state_reg[108]  ( .D(\w0[0][108] ), .CLK(clk), .RST(rst), .Q(state[108]) );
  DFF \state_reg[107]  ( .D(\w0[0][107] ), .CLK(clk), .RST(rst), .Q(state[107]) );
  DFF \state_reg[106]  ( .D(\w0[0][106] ), .CLK(clk), .RST(rst), .Q(state[106]) );
  DFF \state_reg[105]  ( .D(\w0[0][105] ), .CLK(clk), .RST(rst), .Q(state[105]) );
  DFF \state_reg[104]  ( .D(\w0[0][104] ), .CLK(clk), .RST(rst), .Q(state[104]) );
  DFF \state_reg[103]  ( .D(\w0[0][103] ), .CLK(clk), .RST(rst), .Q(state[103]) );
  DFF \state_reg[102]  ( .D(\w0[0][102] ), .CLK(clk), .RST(rst), .Q(state[102]) );
  DFF \state_reg[101]  ( .D(\w0[0][101] ), .CLK(clk), .RST(rst), .Q(state[101]) );
  DFF \state_reg[100]  ( .D(\w0[0][100] ), .CLK(clk), .RST(rst), .Q(state[100]) );
  DFF \state_reg[99]  ( .D(\w0[0][99] ), .CLK(clk), .RST(rst), .Q(state[99])
         );
  DFF \state_reg[98]  ( .D(\w0[0][98] ), .CLK(clk), .RST(rst), .Q(state[98])
         );
  DFF \state_reg[97]  ( .D(\w0[0][97] ), .CLK(clk), .RST(rst), .Q(state[97])
         );
  DFF \state_reg[96]  ( .D(\w0[0][96] ), .CLK(clk), .RST(rst), .Q(state[96])
         );
  DFF \state_reg[95]  ( .D(\w0[0][95] ), .CLK(clk), .RST(rst), .Q(state[95])
         );
  DFF \state_reg[94]  ( .D(\w0[0][94] ), .CLK(clk), .RST(rst), .Q(state[94])
         );
  DFF \state_reg[93]  ( .D(\w0[0][93] ), .CLK(clk), .RST(rst), .Q(state[93])
         );
  DFF \state_reg[92]  ( .D(\w0[0][92] ), .CLK(clk), .RST(rst), .Q(state[92])
         );
  DFF \state_reg[91]  ( .D(\w0[0][91] ), .CLK(clk), .RST(rst), .Q(state[91])
         );
  DFF \state_reg[90]  ( .D(\w0[0][90] ), .CLK(clk), .RST(rst), .Q(state[90])
         );
  DFF \state_reg[89]  ( .D(\w0[0][89] ), .CLK(clk), .RST(rst), .Q(state[89])
         );
  DFF \state_reg[88]  ( .D(\w0[0][88] ), .CLK(clk), .RST(rst), .Q(state[88])
         );
  DFF \state_reg[87]  ( .D(\w0[0][87] ), .CLK(clk), .RST(rst), .Q(state[87])
         );
  DFF \state_reg[86]  ( .D(\w0[0][86] ), .CLK(clk), .RST(rst), .Q(state[86])
         );
  DFF \state_reg[85]  ( .D(\w0[0][85] ), .CLK(clk), .RST(rst), .Q(state[85])
         );
  DFF \state_reg[84]  ( .D(\w0[0][84] ), .CLK(clk), .RST(rst), .Q(state[84])
         );
  DFF \state_reg[83]  ( .D(\w0[0][83] ), .CLK(clk), .RST(rst), .Q(state[83])
         );
  DFF \state_reg[82]  ( .D(\w0[0][82] ), .CLK(clk), .RST(rst), .Q(state[82])
         );
  DFF \state_reg[81]  ( .D(\w0[0][81] ), .CLK(clk), .RST(rst), .Q(state[81])
         );
  DFF \state_reg[80]  ( .D(\w0[0][80] ), .CLK(clk), .RST(rst), .Q(state[80])
         );
  DFF \state_reg[79]  ( .D(\w0[0][79] ), .CLK(clk), .RST(rst), .Q(state[79])
         );
  DFF \state_reg[78]  ( .D(\w0[0][78] ), .CLK(clk), .RST(rst), .Q(state[78])
         );
  DFF \state_reg[77]  ( .D(\w0[0][77] ), .CLK(clk), .RST(rst), .Q(state[77])
         );
  DFF \state_reg[76]  ( .D(\w0[0][76] ), .CLK(clk), .RST(rst), .Q(state[76])
         );
  DFF \state_reg[75]  ( .D(\w0[0][75] ), .CLK(clk), .RST(rst), .Q(state[75])
         );
  DFF \state_reg[74]  ( .D(\w0[0][74] ), .CLK(clk), .RST(rst), .Q(state[74])
         );
  DFF \state_reg[73]  ( .D(\w0[0][73] ), .CLK(clk), .RST(rst), .Q(state[73])
         );
  DFF \state_reg[72]  ( .D(\w0[0][72] ), .CLK(clk), .RST(rst), .Q(state[72])
         );
  DFF \state_reg[71]  ( .D(\w0[0][71] ), .CLK(clk), .RST(rst), .Q(state[71])
         );
  DFF \state_reg[70]  ( .D(\w0[0][70] ), .CLK(clk), .RST(rst), .Q(state[70])
         );
  DFF \state_reg[69]  ( .D(\w0[0][69] ), .CLK(clk), .RST(rst), .Q(state[69])
         );
  DFF \state_reg[68]  ( .D(\w0[0][68] ), .CLK(clk), .RST(rst), .Q(state[68])
         );
  DFF \state_reg[67]  ( .D(\w0[0][67] ), .CLK(clk), .RST(rst), .Q(state[67])
         );
  DFF \state_reg[66]  ( .D(\w0[0][66] ), .CLK(clk), .RST(rst), .Q(state[66])
         );
  DFF \state_reg[65]  ( .D(\w0[0][65] ), .CLK(clk), .RST(rst), .Q(state[65])
         );
  DFF \state_reg[64]  ( .D(\w0[0][64] ), .CLK(clk), .RST(rst), .Q(state[64])
         );
  DFF \state_reg[63]  ( .D(\w0[0][63] ), .CLK(clk), .RST(rst), .Q(state[63])
         );
  DFF \state_reg[62]  ( .D(\w0[0][62] ), .CLK(clk), .RST(rst), .Q(state[62])
         );
  DFF \state_reg[61]  ( .D(\w0[0][61] ), .CLK(clk), .RST(rst), .Q(state[61])
         );
  DFF \state_reg[60]  ( .D(\w0[0][60] ), .CLK(clk), .RST(rst), .Q(state[60])
         );
  DFF \state_reg[59]  ( .D(\w0[0][59] ), .CLK(clk), .RST(rst), .Q(state[59])
         );
  DFF \state_reg[58]  ( .D(\w0[0][58] ), .CLK(clk), .RST(rst), .Q(state[58])
         );
  DFF \state_reg[57]  ( .D(\w0[0][57] ), .CLK(clk), .RST(rst), .Q(state[57])
         );
  DFF \state_reg[56]  ( .D(\w0[0][56] ), .CLK(clk), .RST(rst), .Q(state[56])
         );
  DFF \state_reg[55]  ( .D(\w0[0][55] ), .CLK(clk), .RST(rst), .Q(state[55])
         );
  DFF \state_reg[54]  ( .D(\w0[0][54] ), .CLK(clk), .RST(rst), .Q(state[54])
         );
  DFF \state_reg[53]  ( .D(\w0[0][53] ), .CLK(clk), .RST(rst), .Q(state[53])
         );
  DFF \state_reg[52]  ( .D(\w0[0][52] ), .CLK(clk), .RST(rst), .Q(state[52])
         );
  DFF \state_reg[51]  ( .D(\w0[0][51] ), .CLK(clk), .RST(rst), .Q(state[51])
         );
  DFF \state_reg[50]  ( .D(\w0[0][50] ), .CLK(clk), .RST(rst), .Q(state[50])
         );
  DFF \state_reg[49]  ( .D(\w0[0][49] ), .CLK(clk), .RST(rst), .Q(state[49])
         );
  DFF \state_reg[48]  ( .D(\w0[0][48] ), .CLK(clk), .RST(rst), .Q(state[48])
         );
  DFF \state_reg[47]  ( .D(\w0[0][47] ), .CLK(clk), .RST(rst), .Q(state[47])
         );
  DFF \state_reg[46]  ( .D(\w0[0][46] ), .CLK(clk), .RST(rst), .Q(state[46])
         );
  DFF \state_reg[45]  ( .D(\w0[0][45] ), .CLK(clk), .RST(rst), .Q(state[45])
         );
  DFF \state_reg[44]  ( .D(\w0[0][44] ), .CLK(clk), .RST(rst), .Q(state[44])
         );
  DFF \state_reg[43]  ( .D(\w0[0][43] ), .CLK(clk), .RST(rst), .Q(state[43])
         );
  DFF \state_reg[42]  ( .D(\w0[0][42] ), .CLK(clk), .RST(rst), .Q(state[42])
         );
  DFF \state_reg[41]  ( .D(\w0[0][41] ), .CLK(clk), .RST(rst), .Q(state[41])
         );
  DFF \state_reg[40]  ( .D(\w0[0][40] ), .CLK(clk), .RST(rst), .Q(state[40])
         );
  DFF \state_reg[39]  ( .D(\w0[0][39] ), .CLK(clk), .RST(rst), .Q(state[39])
         );
  DFF \state_reg[38]  ( .D(\w0[0][38] ), .CLK(clk), .RST(rst), .Q(state[38])
         );
  DFF \state_reg[37]  ( .D(\w0[0][37] ), .CLK(clk), .RST(rst), .Q(state[37])
         );
  DFF \state_reg[36]  ( .D(\w0[0][36] ), .CLK(clk), .RST(rst), .Q(state[36])
         );
  DFF \state_reg[35]  ( .D(\w0[0][35] ), .CLK(clk), .RST(rst), .Q(state[35])
         );
  DFF \state_reg[34]  ( .D(\w0[0][34] ), .CLK(clk), .RST(rst), .Q(state[34])
         );
  DFF \state_reg[33]  ( .D(\w0[0][33] ), .CLK(clk), .RST(rst), .Q(state[33])
         );
  DFF \state_reg[32]  ( .D(\w0[0][32] ), .CLK(clk), .RST(rst), .Q(state[32])
         );
  DFF \state_reg[31]  ( .D(\w0[0][31] ), .CLK(clk), .RST(rst), .Q(state[31])
         );
  DFF \state_reg[30]  ( .D(\w0[0][30] ), .CLK(clk), .RST(rst), .Q(state[30])
         );
  DFF \state_reg[29]  ( .D(\w0[0][29] ), .CLK(clk), .RST(rst), .Q(state[29])
         );
  DFF \state_reg[28]  ( .D(\w0[0][28] ), .CLK(clk), .RST(rst), .Q(state[28])
         );
  DFF \state_reg[27]  ( .D(\w0[0][27] ), .CLK(clk), .RST(rst), .Q(state[27])
         );
  DFF \state_reg[26]  ( .D(\w0[0][26] ), .CLK(clk), .RST(rst), .Q(state[26])
         );
  DFF \state_reg[25]  ( .D(\w0[0][25] ), .CLK(clk), .RST(rst), .Q(state[25])
         );
  DFF \state_reg[24]  ( .D(\w0[0][24] ), .CLK(clk), .RST(rst), .Q(state[24])
         );
  DFF \state_reg[23]  ( .D(\w0[0][23] ), .CLK(clk), .RST(rst), .Q(state[23])
         );
  DFF \state_reg[22]  ( .D(\w0[0][22] ), .CLK(clk), .RST(rst), .Q(state[22])
         );
  DFF \state_reg[21]  ( .D(\w0[0][21] ), .CLK(clk), .RST(rst), .Q(state[21])
         );
  DFF \state_reg[20]  ( .D(\w0[0][20] ), .CLK(clk), .RST(rst), .Q(state[20])
         );
  DFF \state_reg[19]  ( .D(\w0[0][19] ), .CLK(clk), .RST(rst), .Q(state[19])
         );
  DFF \state_reg[18]  ( .D(\w0[0][18] ), .CLK(clk), .RST(rst), .Q(state[18])
         );
  DFF \state_reg[17]  ( .D(\w0[0][17] ), .CLK(clk), .RST(rst), .Q(state[17])
         );
  DFF \state_reg[16]  ( .D(\w0[0][16] ), .CLK(clk), .RST(rst), .Q(state[16])
         );
  DFF \state_reg[15]  ( .D(\w0[0][15] ), .CLK(clk), .RST(rst), .Q(state[15])
         );
  DFF \state_reg[14]  ( .D(\w0[0][14] ), .CLK(clk), .RST(rst), .Q(state[14])
         );
  DFF \state_reg[13]  ( .D(\w0[0][13] ), .CLK(clk), .RST(rst), .Q(state[13])
         );
  DFF \state_reg[12]  ( .D(\w0[0][12] ), .CLK(clk), .RST(rst), .Q(state[12])
         );
  DFF \state_reg[11]  ( .D(\w0[0][11] ), .CLK(clk), .RST(rst), .Q(state[11])
         );
  DFF \state_reg[10]  ( .D(\w0[0][10] ), .CLK(clk), .RST(rst), .Q(state[10])
         );
  DFF \state_reg[9]  ( .D(\w0[0][9] ), .CLK(clk), .RST(rst), .Q(state[9]) );
  DFF \state_reg[8]  ( .D(\w0[0][8] ), .CLK(clk), .RST(rst), .Q(state[8]) );
  DFF \state_reg[7]  ( .D(\w0[0][7] ), .CLK(clk), .RST(rst), .Q(state[7]) );
  DFF \state_reg[6]  ( .D(\w0[0][6] ), .CLK(clk), .RST(rst), .Q(state[6]) );
  DFF \state_reg[5]  ( .D(\w0[0][5] ), .CLK(clk), .RST(rst), .Q(state[5]) );
  DFF \state_reg[4]  ( .D(\w0[0][4] ), .CLK(clk), .RST(rst), .Q(state[4]) );
  DFF \state_reg[3]  ( .D(\w0[0][3] ), .CLK(clk), .RST(rst), .Q(state[3]) );
  DFF \state_reg[2]  ( .D(\w0[0][2] ), .CLK(clk), .RST(rst), .Q(state[2]) );
  DFF \state_reg[1]  ( .D(\w0[0][1] ), .CLK(clk), .RST(rst), .Q(state[1]) );
  DFF \state_reg[0]  ( .D(\w0[0][0] ), .CLK(clk), .RST(rst), .Q(state[0]) );
  XOR U643 ( .A(key[0]), .B(\w3[0][0] ), .Z(out[0]) );
  XOR U644 ( .A(key[100]), .B(\w3[0][100] ), .Z(out[100]) );
  XOR U645 ( .A(key[101]), .B(\w3[0][101] ), .Z(out[101]) );
  XOR U646 ( .A(key[102]), .B(\w3[0][102] ), .Z(out[102]) );
  XOR U647 ( .A(key[103]), .B(\w3[0][103] ), .Z(out[103]) );
  XOR U648 ( .A(key[104]), .B(\w3[0][104] ), .Z(out[104]) );
  XOR U649 ( .A(key[105]), .B(\w3[0][105] ), .Z(out[105]) );
  XOR U650 ( .A(key[106]), .B(\w3[0][106] ), .Z(out[106]) );
  XOR U651 ( .A(key[107]), .B(\w3[0][107] ), .Z(out[107]) );
  XOR U652 ( .A(key[108]), .B(\w3[0][108] ), .Z(out[108]) );
  XOR U653 ( .A(key[109]), .B(\w3[0][109] ), .Z(out[109]) );
  XOR U654 ( .A(key[10]), .B(\w3[0][10] ), .Z(out[10]) );
  XOR U655 ( .A(key[110]), .B(\w3[0][110] ), .Z(out[110]) );
  XOR U656 ( .A(key[111]), .B(\w3[0][111] ), .Z(out[111]) );
  XOR U657 ( .A(key[112]), .B(\w3[0][112] ), .Z(out[112]) );
  XOR U658 ( .A(key[113]), .B(\w3[0][113] ), .Z(out[113]) );
  XOR U659 ( .A(key[114]), .B(\w3[0][114] ), .Z(out[114]) );
  XOR U660 ( .A(key[115]), .B(\w3[0][115] ), .Z(out[115]) );
  XOR U661 ( .A(key[116]), .B(\w3[0][116] ), .Z(out[116]) );
  XOR U662 ( .A(key[117]), .B(\w3[0][117] ), .Z(out[117]) );
  XOR U663 ( .A(key[118]), .B(\w3[0][118] ), .Z(out[118]) );
  XOR U664 ( .A(key[119]), .B(\w3[0][119] ), .Z(out[119]) );
  XOR U665 ( .A(key[11]), .B(\w3[0][11] ), .Z(out[11]) );
  XOR U666 ( .A(key[120]), .B(\w3[0][120] ), .Z(out[120]) );
  XOR U667 ( .A(key[121]), .B(\w3[0][121] ), .Z(out[121]) );
  XOR U668 ( .A(key[122]), .B(\w3[0][122] ), .Z(out[122]) );
  XOR U669 ( .A(key[123]), .B(\w3[0][123] ), .Z(out[123]) );
  XOR U670 ( .A(key[124]), .B(\w3[0][124] ), .Z(out[124]) );
  XOR U671 ( .A(key[125]), .B(\w3[0][125] ), .Z(out[125]) );
  XOR U672 ( .A(key[126]), .B(\w3[0][126] ), .Z(out[126]) );
  XOR U673 ( .A(key[127]), .B(\w3[0][127] ), .Z(out[127]) );
  XOR U674 ( .A(key[12]), .B(\w3[0][12] ), .Z(out[12]) );
  XOR U675 ( .A(key[13]), .B(\w3[0][13] ), .Z(out[13]) );
  XOR U676 ( .A(key[14]), .B(\w3[0][14] ), .Z(out[14]) );
  XOR U677 ( .A(key[15]), .B(\w3[0][15] ), .Z(out[15]) );
  XOR U678 ( .A(key[16]), .B(\w3[0][16] ), .Z(out[16]) );
  XOR U679 ( .A(key[17]), .B(\w3[0][17] ), .Z(out[17]) );
  XOR U680 ( .A(key[18]), .B(\w3[0][18] ), .Z(out[18]) );
  XOR U681 ( .A(key[19]), .B(\w3[0][19] ), .Z(out[19]) );
  XOR U682 ( .A(key[1]), .B(\w3[0][1] ), .Z(out[1]) );
  XOR U683 ( .A(key[20]), .B(\w3[0][20] ), .Z(out[20]) );
  XOR U684 ( .A(key[21]), .B(\w3[0][21] ), .Z(out[21]) );
  XOR U685 ( .A(key[22]), .B(\w3[0][22] ), .Z(out[22]) );
  XOR U686 ( .A(key[23]), .B(\w3[0][23] ), .Z(out[23]) );
  XOR U687 ( .A(key[24]), .B(\w3[0][24] ), .Z(out[24]) );
  XOR U688 ( .A(key[25]), .B(\w3[0][25] ), .Z(out[25]) );
  XOR U689 ( .A(key[26]), .B(\w3[0][26] ), .Z(out[26]) );
  XOR U690 ( .A(key[27]), .B(\w3[0][27] ), .Z(out[27]) );
  XOR U691 ( .A(key[28]), .B(\w3[0][28] ), .Z(out[28]) );
  XOR U692 ( .A(key[29]), .B(\w3[0][29] ), .Z(out[29]) );
  XOR U693 ( .A(key[2]), .B(\w3[0][2] ), .Z(out[2]) );
  XOR U694 ( .A(key[30]), .B(\w3[0][30] ), .Z(out[30]) );
  XOR U695 ( .A(key[31]), .B(\w3[0][31] ), .Z(out[31]) );
  XOR U696 ( .A(key[32]), .B(\w3[0][32] ), .Z(out[32]) );
  XOR U697 ( .A(key[33]), .B(\w3[0][33] ), .Z(out[33]) );
  XOR U698 ( .A(key[34]), .B(\w3[0][34] ), .Z(out[34]) );
  XOR U699 ( .A(key[35]), .B(\w3[0][35] ), .Z(out[35]) );
  XOR U700 ( .A(key[36]), .B(\w3[0][36] ), .Z(out[36]) );
  XOR U701 ( .A(key[37]), .B(\w3[0][37] ), .Z(out[37]) );
  XOR U702 ( .A(key[38]), .B(\w3[0][38] ), .Z(out[38]) );
  XOR U703 ( .A(key[39]), .B(\w3[0][39] ), .Z(out[39]) );
  XOR U704 ( .A(key[3]), .B(\w3[0][3] ), .Z(out[3]) );
  XOR U705 ( .A(key[40]), .B(\w3[0][40] ), .Z(out[40]) );
  XOR U706 ( .A(key[41]), .B(\w3[0][41] ), .Z(out[41]) );
  XOR U707 ( .A(key[42]), .B(\w3[0][42] ), .Z(out[42]) );
  XOR U708 ( .A(key[43]), .B(\w3[0][43] ), .Z(out[43]) );
  XOR U709 ( .A(key[44]), .B(\w3[0][44] ), .Z(out[44]) );
  XOR U710 ( .A(key[45]), .B(\w3[0][45] ), .Z(out[45]) );
  XOR U711 ( .A(key[46]), .B(\w3[0][46] ), .Z(out[46]) );
  XOR U712 ( .A(key[47]), .B(\w3[0][47] ), .Z(out[47]) );
  XOR U713 ( .A(key[48]), .B(\w3[0][48] ), .Z(out[48]) );
  XOR U714 ( .A(key[49]), .B(\w3[0][49] ), .Z(out[49]) );
  XOR U715 ( .A(key[4]), .B(\w3[0][4] ), .Z(out[4]) );
  XOR U716 ( .A(key[50]), .B(\w3[0][50] ), .Z(out[50]) );
  XOR U717 ( .A(key[51]), .B(\w3[0][51] ), .Z(out[51]) );
  XOR U718 ( .A(key[52]), .B(\w3[0][52] ), .Z(out[52]) );
  XOR U719 ( .A(key[53]), .B(\w3[0][53] ), .Z(out[53]) );
  XOR U720 ( .A(key[54]), .B(\w3[0][54] ), .Z(out[54]) );
  XOR U721 ( .A(key[55]), .B(\w3[0][55] ), .Z(out[55]) );
  XOR U722 ( .A(key[56]), .B(\w3[0][56] ), .Z(out[56]) );
  XOR U723 ( .A(key[57]), .B(\w3[0][57] ), .Z(out[57]) );
  XOR U724 ( .A(key[58]), .B(\w3[0][58] ), .Z(out[58]) );
  XOR U725 ( .A(key[59]), .B(\w3[0][59] ), .Z(out[59]) );
  XOR U726 ( .A(key[5]), .B(\w3[0][5] ), .Z(out[5]) );
  XOR U727 ( .A(key[60]), .B(\w3[0][60] ), .Z(out[60]) );
  XOR U728 ( .A(key[61]), .B(\w3[0][61] ), .Z(out[61]) );
  XOR U729 ( .A(key[62]), .B(\w3[0][62] ), .Z(out[62]) );
  XOR U730 ( .A(key[63]), .B(\w3[0][63] ), .Z(out[63]) );
  XOR U731 ( .A(key[64]), .B(\w3[0][64] ), .Z(out[64]) );
  XOR U732 ( .A(key[65]), .B(\w3[0][65] ), .Z(out[65]) );
  XOR U733 ( .A(key[66]), .B(\w3[0][66] ), .Z(out[66]) );
  XOR U734 ( .A(key[67]), .B(\w3[0][67] ), .Z(out[67]) );
  XOR U735 ( .A(key[68]), .B(\w3[0][68] ), .Z(out[68]) );
  XOR U736 ( .A(key[69]), .B(\w3[0][69] ), .Z(out[69]) );
  XOR U737 ( .A(key[6]), .B(\w3[0][6] ), .Z(out[6]) );
  XOR U738 ( .A(key[70]), .B(\w3[0][70] ), .Z(out[70]) );
  XOR U739 ( .A(key[71]), .B(\w3[0][71] ), .Z(out[71]) );
  XOR U740 ( .A(key[72]), .B(\w3[0][72] ), .Z(out[72]) );
  XOR U741 ( .A(key[73]), .B(\w3[0][73] ), .Z(out[73]) );
  XOR U742 ( .A(key[74]), .B(\w3[0][74] ), .Z(out[74]) );
  XOR U743 ( .A(key[75]), .B(\w3[0][75] ), .Z(out[75]) );
  XOR U744 ( .A(key[76]), .B(\w3[0][76] ), .Z(out[76]) );
  XOR U745 ( .A(key[77]), .B(\w3[0][77] ), .Z(out[77]) );
  XOR U746 ( .A(key[78]), .B(\w3[0][78] ), .Z(out[78]) );
  XOR U747 ( .A(key[79]), .B(\w3[0][79] ), .Z(out[79]) );
  XOR U748 ( .A(key[7]), .B(\w3[0][7] ), .Z(out[7]) );
  XOR U749 ( .A(key[80]), .B(\w3[0][80] ), .Z(out[80]) );
  XOR U750 ( .A(key[81]), .B(\w3[0][81] ), .Z(out[81]) );
  XOR U751 ( .A(key[82]), .B(\w3[0][82] ), .Z(out[82]) );
  XOR U752 ( .A(key[83]), .B(\w3[0][83] ), .Z(out[83]) );
  XOR U753 ( .A(key[84]), .B(\w3[0][84] ), .Z(out[84]) );
  XOR U754 ( .A(key[85]), .B(\w3[0][85] ), .Z(out[85]) );
  XOR U755 ( .A(key[86]), .B(\w3[0][86] ), .Z(out[86]) );
  XOR U756 ( .A(key[87]), .B(\w3[0][87] ), .Z(out[87]) );
  XOR U757 ( .A(key[88]), .B(\w3[0][88] ), .Z(out[88]) );
  XOR U758 ( .A(key[89]), .B(\w3[0][89] ), .Z(out[89]) );
  XOR U759 ( .A(key[8]), .B(\w3[0][8] ), .Z(out[8]) );
  XOR U760 ( .A(key[90]), .B(\w3[0][90] ), .Z(out[90]) );
  XOR U761 ( .A(key[91]), .B(\w3[0][91] ), .Z(out[91]) );
  XOR U762 ( .A(key[92]), .B(\w3[0][92] ), .Z(out[92]) );
  XOR U763 ( .A(key[93]), .B(\w3[0][93] ), .Z(out[93]) );
  XOR U764 ( .A(key[94]), .B(\w3[0][94] ), .Z(out[94]) );
  XOR U765 ( .A(key[95]), .B(\w3[0][95] ), .Z(out[95]) );
  XOR U766 ( .A(key[96]), .B(\w3[0][96] ), .Z(out[96]) );
  XOR U767 ( .A(key[97]), .B(\w3[0][97] ), .Z(out[97]) );
  XOR U768 ( .A(key[98]), .B(\w3[0][98] ), .Z(out[98]) );
  XOR U769 ( .A(key[99]), .B(\w3[0][99] ), .Z(out[99]) );
  XOR U770 ( .A(key[9]), .B(\w3[0][9] ), .Z(out[9]) );
  NAND U771 ( .A(state[0]), .B(init), .Z(n258) );
  NANDN U772 ( .A(init), .B(msg[0]), .Z(n257) );
  NAND U773 ( .A(n258), .B(n257), .Z(\w0[0][0] ) );
  NAND U774 ( .A(state[100]), .B(init), .Z(n260) );
  NANDN U775 ( .A(init), .B(msg[100]), .Z(n259) );
  NAND U776 ( .A(n260), .B(n259), .Z(\w0[0][100] ) );
  NAND U777 ( .A(state[101]), .B(init), .Z(n262) );
  NANDN U778 ( .A(init), .B(msg[101]), .Z(n261) );
  NAND U779 ( .A(n262), .B(n261), .Z(\w0[0][101] ) );
  NAND U780 ( .A(state[102]), .B(init), .Z(n264) );
  NANDN U781 ( .A(init), .B(msg[102]), .Z(n263) );
  NAND U782 ( .A(n264), .B(n263), .Z(\w0[0][102] ) );
  NAND U783 ( .A(state[103]), .B(init), .Z(n266) );
  NANDN U784 ( .A(init), .B(msg[103]), .Z(n265) );
  NAND U785 ( .A(n266), .B(n265), .Z(\w0[0][103] ) );
  NAND U786 ( .A(state[104]), .B(init), .Z(n268) );
  NANDN U787 ( .A(init), .B(msg[104]), .Z(n267) );
  NAND U788 ( .A(n268), .B(n267), .Z(\w0[0][104] ) );
  NAND U789 ( .A(state[105]), .B(init), .Z(n270) );
  NANDN U790 ( .A(init), .B(msg[105]), .Z(n269) );
  NAND U791 ( .A(n270), .B(n269), .Z(\w0[0][105] ) );
  NAND U792 ( .A(state[106]), .B(init), .Z(n272) );
  NANDN U793 ( .A(init), .B(msg[106]), .Z(n271) );
  NAND U794 ( .A(n272), .B(n271), .Z(\w0[0][106] ) );
  NAND U795 ( .A(state[107]), .B(init), .Z(n274) );
  NANDN U796 ( .A(init), .B(msg[107]), .Z(n273) );
  NAND U797 ( .A(n274), .B(n273), .Z(\w0[0][107] ) );
  NAND U798 ( .A(state[108]), .B(init), .Z(n276) );
  NANDN U799 ( .A(init), .B(msg[108]), .Z(n275) );
  NAND U800 ( .A(n276), .B(n275), .Z(\w0[0][108] ) );
  NAND U801 ( .A(state[109]), .B(init), .Z(n278) );
  NANDN U802 ( .A(init), .B(msg[109]), .Z(n277) );
  NAND U803 ( .A(n278), .B(n277), .Z(\w0[0][109] ) );
  NAND U804 ( .A(state[10]), .B(init), .Z(n280) );
  NANDN U805 ( .A(init), .B(msg[10]), .Z(n279) );
  NAND U806 ( .A(n280), .B(n279), .Z(\w0[0][10] ) );
  NAND U807 ( .A(state[110]), .B(init), .Z(n282) );
  NANDN U808 ( .A(init), .B(msg[110]), .Z(n281) );
  NAND U809 ( .A(n282), .B(n281), .Z(\w0[0][110] ) );
  NAND U810 ( .A(state[111]), .B(init), .Z(n284) );
  NANDN U811 ( .A(init), .B(msg[111]), .Z(n283) );
  NAND U812 ( .A(n284), .B(n283), .Z(\w0[0][111] ) );
  NAND U813 ( .A(state[112]), .B(init), .Z(n286) );
  NANDN U814 ( .A(init), .B(msg[112]), .Z(n285) );
  NAND U815 ( .A(n286), .B(n285), .Z(\w0[0][112] ) );
  NAND U816 ( .A(state[113]), .B(init), .Z(n288) );
  NANDN U817 ( .A(init), .B(msg[113]), .Z(n287) );
  NAND U818 ( .A(n288), .B(n287), .Z(\w0[0][113] ) );
  NAND U819 ( .A(state[114]), .B(init), .Z(n290) );
  NANDN U820 ( .A(init), .B(msg[114]), .Z(n289) );
  NAND U821 ( .A(n290), .B(n289), .Z(\w0[0][114] ) );
  NAND U822 ( .A(state[115]), .B(init), .Z(n292) );
  NANDN U823 ( .A(init), .B(msg[115]), .Z(n291) );
  NAND U824 ( .A(n292), .B(n291), .Z(\w0[0][115] ) );
  NAND U825 ( .A(state[116]), .B(init), .Z(n294) );
  NANDN U826 ( .A(init), .B(msg[116]), .Z(n293) );
  NAND U827 ( .A(n294), .B(n293), .Z(\w0[0][116] ) );
  NAND U828 ( .A(state[117]), .B(init), .Z(n296) );
  NANDN U829 ( .A(init), .B(msg[117]), .Z(n295) );
  NAND U830 ( .A(n296), .B(n295), .Z(\w0[0][117] ) );
  NAND U831 ( .A(state[118]), .B(init), .Z(n298) );
  NANDN U832 ( .A(init), .B(msg[118]), .Z(n297) );
  NAND U833 ( .A(n298), .B(n297), .Z(\w0[0][118] ) );
  NAND U834 ( .A(state[119]), .B(init), .Z(n300) );
  NANDN U835 ( .A(init), .B(msg[119]), .Z(n299) );
  NAND U836 ( .A(n300), .B(n299), .Z(\w0[0][119] ) );
  NAND U837 ( .A(state[11]), .B(init), .Z(n302) );
  NANDN U838 ( .A(init), .B(msg[11]), .Z(n301) );
  NAND U839 ( .A(n302), .B(n301), .Z(\w0[0][11] ) );
  NAND U840 ( .A(state[120]), .B(init), .Z(n304) );
  NANDN U841 ( .A(init), .B(msg[120]), .Z(n303) );
  NAND U842 ( .A(n304), .B(n303), .Z(\w0[0][120] ) );
  NAND U843 ( .A(state[121]), .B(init), .Z(n306) );
  NANDN U844 ( .A(init), .B(msg[121]), .Z(n305) );
  NAND U845 ( .A(n306), .B(n305), .Z(\w0[0][121] ) );
  NAND U846 ( .A(state[122]), .B(init), .Z(n308) );
  NANDN U847 ( .A(init), .B(msg[122]), .Z(n307) );
  NAND U848 ( .A(n308), .B(n307), .Z(\w0[0][122] ) );
  NAND U849 ( .A(state[123]), .B(init), .Z(n310) );
  NANDN U850 ( .A(init), .B(msg[123]), .Z(n309) );
  NAND U851 ( .A(n310), .B(n309), .Z(\w0[0][123] ) );
  NAND U852 ( .A(state[124]), .B(init), .Z(n312) );
  NANDN U853 ( .A(init), .B(msg[124]), .Z(n311) );
  NAND U854 ( .A(n312), .B(n311), .Z(\w0[0][124] ) );
  NAND U855 ( .A(state[125]), .B(init), .Z(n314) );
  NANDN U856 ( .A(init), .B(msg[125]), .Z(n313) );
  NAND U857 ( .A(n314), .B(n313), .Z(\w0[0][125] ) );
  NAND U858 ( .A(state[126]), .B(init), .Z(n316) );
  NANDN U859 ( .A(init), .B(msg[126]), .Z(n315) );
  NAND U860 ( .A(n316), .B(n315), .Z(\w0[0][126] ) );
  NAND U861 ( .A(state[127]), .B(init), .Z(n318) );
  NANDN U862 ( .A(init), .B(msg[127]), .Z(n317) );
  NAND U863 ( .A(n318), .B(n317), .Z(\w0[0][127] ) );
  NAND U864 ( .A(state[12]), .B(init), .Z(n320) );
  NANDN U865 ( .A(init), .B(msg[12]), .Z(n319) );
  NAND U866 ( .A(n320), .B(n319), .Z(\w0[0][12] ) );
  NAND U867 ( .A(state[13]), .B(init), .Z(n322) );
  NANDN U868 ( .A(init), .B(msg[13]), .Z(n321) );
  NAND U869 ( .A(n322), .B(n321), .Z(\w0[0][13] ) );
  NAND U870 ( .A(state[14]), .B(init), .Z(n324) );
  NANDN U871 ( .A(init), .B(msg[14]), .Z(n323) );
  NAND U872 ( .A(n324), .B(n323), .Z(\w0[0][14] ) );
  NAND U873 ( .A(state[15]), .B(init), .Z(n326) );
  NANDN U874 ( .A(init), .B(msg[15]), .Z(n325) );
  NAND U875 ( .A(n326), .B(n325), .Z(\w0[0][15] ) );
  NAND U876 ( .A(state[16]), .B(init), .Z(n328) );
  NANDN U877 ( .A(init), .B(msg[16]), .Z(n327) );
  NAND U878 ( .A(n328), .B(n327), .Z(\w0[0][16] ) );
  NAND U879 ( .A(state[17]), .B(init), .Z(n330) );
  NANDN U880 ( .A(init), .B(msg[17]), .Z(n329) );
  NAND U881 ( .A(n330), .B(n329), .Z(\w0[0][17] ) );
  NAND U882 ( .A(state[18]), .B(init), .Z(n332) );
  NANDN U883 ( .A(init), .B(msg[18]), .Z(n331) );
  NAND U884 ( .A(n332), .B(n331), .Z(\w0[0][18] ) );
  NAND U885 ( .A(state[19]), .B(init), .Z(n334) );
  NANDN U886 ( .A(init), .B(msg[19]), .Z(n333) );
  NAND U887 ( .A(n334), .B(n333), .Z(\w0[0][19] ) );
  NAND U888 ( .A(state[1]), .B(init), .Z(n336) );
  NANDN U889 ( .A(init), .B(msg[1]), .Z(n335) );
  NAND U890 ( .A(n336), .B(n335), .Z(\w0[0][1] ) );
  NAND U891 ( .A(state[20]), .B(init), .Z(n338) );
  NANDN U892 ( .A(init), .B(msg[20]), .Z(n337) );
  NAND U893 ( .A(n338), .B(n337), .Z(\w0[0][20] ) );
  NAND U894 ( .A(state[21]), .B(init), .Z(n340) );
  NANDN U895 ( .A(init), .B(msg[21]), .Z(n339) );
  NAND U896 ( .A(n340), .B(n339), .Z(\w0[0][21] ) );
  NAND U897 ( .A(state[22]), .B(init), .Z(n342) );
  NANDN U898 ( .A(init), .B(msg[22]), .Z(n341) );
  NAND U899 ( .A(n342), .B(n341), .Z(\w0[0][22] ) );
  NAND U900 ( .A(state[23]), .B(init), .Z(n344) );
  NANDN U901 ( .A(init), .B(msg[23]), .Z(n343) );
  NAND U902 ( .A(n344), .B(n343), .Z(\w0[0][23] ) );
  NAND U903 ( .A(state[24]), .B(init), .Z(n346) );
  NANDN U904 ( .A(init), .B(msg[24]), .Z(n345) );
  NAND U905 ( .A(n346), .B(n345), .Z(\w0[0][24] ) );
  NAND U906 ( .A(state[25]), .B(init), .Z(n348) );
  NANDN U907 ( .A(init), .B(msg[25]), .Z(n347) );
  NAND U908 ( .A(n348), .B(n347), .Z(\w0[0][25] ) );
  NAND U909 ( .A(state[26]), .B(init), .Z(n350) );
  NANDN U910 ( .A(init), .B(msg[26]), .Z(n349) );
  NAND U911 ( .A(n350), .B(n349), .Z(\w0[0][26] ) );
  NAND U912 ( .A(state[27]), .B(init), .Z(n352) );
  NANDN U913 ( .A(init), .B(msg[27]), .Z(n351) );
  NAND U914 ( .A(n352), .B(n351), .Z(\w0[0][27] ) );
  NAND U915 ( .A(state[28]), .B(init), .Z(n354) );
  NANDN U916 ( .A(init), .B(msg[28]), .Z(n353) );
  NAND U917 ( .A(n354), .B(n353), .Z(\w0[0][28] ) );
  NAND U918 ( .A(state[29]), .B(init), .Z(n356) );
  NANDN U919 ( .A(init), .B(msg[29]), .Z(n355) );
  NAND U920 ( .A(n356), .B(n355), .Z(\w0[0][29] ) );
  NAND U921 ( .A(state[2]), .B(init), .Z(n358) );
  NANDN U922 ( .A(init), .B(msg[2]), .Z(n357) );
  NAND U923 ( .A(n358), .B(n357), .Z(\w0[0][2] ) );
  NAND U924 ( .A(state[30]), .B(init), .Z(n360) );
  NANDN U925 ( .A(init), .B(msg[30]), .Z(n359) );
  NAND U926 ( .A(n360), .B(n359), .Z(\w0[0][30] ) );
  NAND U927 ( .A(state[31]), .B(init), .Z(n362) );
  NANDN U928 ( .A(init), .B(msg[31]), .Z(n361) );
  NAND U929 ( .A(n362), .B(n361), .Z(\w0[0][31] ) );
  NAND U930 ( .A(state[32]), .B(init), .Z(n364) );
  NANDN U931 ( .A(init), .B(msg[32]), .Z(n363) );
  NAND U932 ( .A(n364), .B(n363), .Z(\w0[0][32] ) );
  NAND U933 ( .A(state[33]), .B(init), .Z(n366) );
  NANDN U934 ( .A(init), .B(msg[33]), .Z(n365) );
  NAND U935 ( .A(n366), .B(n365), .Z(\w0[0][33] ) );
  NAND U936 ( .A(state[34]), .B(init), .Z(n368) );
  NANDN U937 ( .A(init), .B(msg[34]), .Z(n367) );
  NAND U938 ( .A(n368), .B(n367), .Z(\w0[0][34] ) );
  NAND U939 ( .A(state[35]), .B(init), .Z(n370) );
  NANDN U940 ( .A(init), .B(msg[35]), .Z(n369) );
  NAND U941 ( .A(n370), .B(n369), .Z(\w0[0][35] ) );
  NAND U942 ( .A(state[36]), .B(init), .Z(n372) );
  NANDN U943 ( .A(init), .B(msg[36]), .Z(n371) );
  NAND U944 ( .A(n372), .B(n371), .Z(\w0[0][36] ) );
  NAND U945 ( .A(state[37]), .B(init), .Z(n374) );
  NANDN U946 ( .A(init), .B(msg[37]), .Z(n373) );
  NAND U947 ( .A(n374), .B(n373), .Z(\w0[0][37] ) );
  NAND U948 ( .A(state[38]), .B(init), .Z(n376) );
  NANDN U949 ( .A(init), .B(msg[38]), .Z(n375) );
  NAND U950 ( .A(n376), .B(n375), .Z(\w0[0][38] ) );
  NAND U951 ( .A(state[39]), .B(init), .Z(n378) );
  NANDN U952 ( .A(init), .B(msg[39]), .Z(n377) );
  NAND U953 ( .A(n378), .B(n377), .Z(\w0[0][39] ) );
  NAND U954 ( .A(state[3]), .B(init), .Z(n380) );
  NANDN U955 ( .A(init), .B(msg[3]), .Z(n379) );
  NAND U956 ( .A(n380), .B(n379), .Z(\w0[0][3] ) );
  NAND U957 ( .A(state[40]), .B(init), .Z(n382) );
  NANDN U958 ( .A(init), .B(msg[40]), .Z(n381) );
  NAND U959 ( .A(n382), .B(n381), .Z(\w0[0][40] ) );
  NAND U960 ( .A(state[41]), .B(init), .Z(n384) );
  NANDN U961 ( .A(init), .B(msg[41]), .Z(n383) );
  NAND U962 ( .A(n384), .B(n383), .Z(\w0[0][41] ) );
  NAND U963 ( .A(state[42]), .B(init), .Z(n386) );
  NANDN U964 ( .A(init), .B(msg[42]), .Z(n385) );
  NAND U965 ( .A(n386), .B(n385), .Z(\w0[0][42] ) );
  NAND U966 ( .A(state[43]), .B(init), .Z(n388) );
  NANDN U967 ( .A(init), .B(msg[43]), .Z(n387) );
  NAND U968 ( .A(n388), .B(n387), .Z(\w0[0][43] ) );
  NAND U969 ( .A(state[44]), .B(init), .Z(n390) );
  NANDN U970 ( .A(init), .B(msg[44]), .Z(n389) );
  NAND U971 ( .A(n390), .B(n389), .Z(\w0[0][44] ) );
  NAND U972 ( .A(state[45]), .B(init), .Z(n392) );
  NANDN U973 ( .A(init), .B(msg[45]), .Z(n391) );
  NAND U974 ( .A(n392), .B(n391), .Z(\w0[0][45] ) );
  NAND U975 ( .A(state[46]), .B(init), .Z(n394) );
  NANDN U976 ( .A(init), .B(msg[46]), .Z(n393) );
  NAND U977 ( .A(n394), .B(n393), .Z(\w0[0][46] ) );
  NAND U978 ( .A(state[47]), .B(init), .Z(n396) );
  NANDN U979 ( .A(init), .B(msg[47]), .Z(n395) );
  NAND U980 ( .A(n396), .B(n395), .Z(\w0[0][47] ) );
  NAND U981 ( .A(state[48]), .B(init), .Z(n398) );
  NANDN U982 ( .A(init), .B(msg[48]), .Z(n397) );
  NAND U983 ( .A(n398), .B(n397), .Z(\w0[0][48] ) );
  NAND U984 ( .A(state[49]), .B(init), .Z(n400) );
  NANDN U985 ( .A(init), .B(msg[49]), .Z(n399) );
  NAND U986 ( .A(n400), .B(n399), .Z(\w0[0][49] ) );
  NAND U987 ( .A(state[4]), .B(init), .Z(n402) );
  NANDN U988 ( .A(init), .B(msg[4]), .Z(n401) );
  NAND U989 ( .A(n402), .B(n401), .Z(\w0[0][4] ) );
  NAND U990 ( .A(state[50]), .B(init), .Z(n404) );
  NANDN U991 ( .A(init), .B(msg[50]), .Z(n403) );
  NAND U992 ( .A(n404), .B(n403), .Z(\w0[0][50] ) );
  NAND U993 ( .A(state[51]), .B(init), .Z(n406) );
  NANDN U994 ( .A(init), .B(msg[51]), .Z(n405) );
  NAND U995 ( .A(n406), .B(n405), .Z(\w0[0][51] ) );
  NAND U996 ( .A(state[52]), .B(init), .Z(n408) );
  NANDN U997 ( .A(init), .B(msg[52]), .Z(n407) );
  NAND U998 ( .A(n408), .B(n407), .Z(\w0[0][52] ) );
  NAND U999 ( .A(state[53]), .B(init), .Z(n410) );
  NANDN U1000 ( .A(init), .B(msg[53]), .Z(n409) );
  NAND U1001 ( .A(n410), .B(n409), .Z(\w0[0][53] ) );
  NAND U1002 ( .A(state[54]), .B(init), .Z(n412) );
  NANDN U1003 ( .A(init), .B(msg[54]), .Z(n411) );
  NAND U1004 ( .A(n412), .B(n411), .Z(\w0[0][54] ) );
  NAND U1005 ( .A(state[55]), .B(init), .Z(n414) );
  NANDN U1006 ( .A(init), .B(msg[55]), .Z(n413) );
  NAND U1007 ( .A(n414), .B(n413), .Z(\w0[0][55] ) );
  NAND U1008 ( .A(state[56]), .B(init), .Z(n416) );
  NANDN U1009 ( .A(init), .B(msg[56]), .Z(n415) );
  NAND U1010 ( .A(n416), .B(n415), .Z(\w0[0][56] ) );
  NAND U1011 ( .A(state[57]), .B(init), .Z(n418) );
  NANDN U1012 ( .A(init), .B(msg[57]), .Z(n417) );
  NAND U1013 ( .A(n418), .B(n417), .Z(\w0[0][57] ) );
  NAND U1014 ( .A(state[58]), .B(init), .Z(n420) );
  NANDN U1015 ( .A(init), .B(msg[58]), .Z(n419) );
  NAND U1016 ( .A(n420), .B(n419), .Z(\w0[0][58] ) );
  NAND U1017 ( .A(state[59]), .B(init), .Z(n422) );
  NANDN U1018 ( .A(init), .B(msg[59]), .Z(n421) );
  NAND U1019 ( .A(n422), .B(n421), .Z(\w0[0][59] ) );
  NAND U1020 ( .A(state[5]), .B(init), .Z(n424) );
  NANDN U1021 ( .A(init), .B(msg[5]), .Z(n423) );
  NAND U1022 ( .A(n424), .B(n423), .Z(\w0[0][5] ) );
  NAND U1023 ( .A(state[60]), .B(init), .Z(n426) );
  NANDN U1024 ( .A(init), .B(msg[60]), .Z(n425) );
  NAND U1025 ( .A(n426), .B(n425), .Z(\w0[0][60] ) );
  NAND U1026 ( .A(state[61]), .B(init), .Z(n428) );
  NANDN U1027 ( .A(init), .B(msg[61]), .Z(n427) );
  NAND U1028 ( .A(n428), .B(n427), .Z(\w0[0][61] ) );
  NAND U1029 ( .A(state[62]), .B(init), .Z(n430) );
  NANDN U1030 ( .A(init), .B(msg[62]), .Z(n429) );
  NAND U1031 ( .A(n430), .B(n429), .Z(\w0[0][62] ) );
  NAND U1032 ( .A(state[63]), .B(init), .Z(n432) );
  NANDN U1033 ( .A(init), .B(msg[63]), .Z(n431) );
  NAND U1034 ( .A(n432), .B(n431), .Z(\w0[0][63] ) );
  NAND U1035 ( .A(state[64]), .B(init), .Z(n434) );
  NANDN U1036 ( .A(init), .B(msg[64]), .Z(n433) );
  NAND U1037 ( .A(n434), .B(n433), .Z(\w0[0][64] ) );
  NAND U1038 ( .A(state[65]), .B(init), .Z(n436) );
  NANDN U1039 ( .A(init), .B(msg[65]), .Z(n435) );
  NAND U1040 ( .A(n436), .B(n435), .Z(\w0[0][65] ) );
  NAND U1041 ( .A(state[66]), .B(init), .Z(n438) );
  NANDN U1042 ( .A(init), .B(msg[66]), .Z(n437) );
  NAND U1043 ( .A(n438), .B(n437), .Z(\w0[0][66] ) );
  NAND U1044 ( .A(state[67]), .B(init), .Z(n440) );
  NANDN U1045 ( .A(init), .B(msg[67]), .Z(n439) );
  NAND U1046 ( .A(n440), .B(n439), .Z(\w0[0][67] ) );
  NAND U1047 ( .A(state[68]), .B(init), .Z(n442) );
  NANDN U1048 ( .A(init), .B(msg[68]), .Z(n441) );
  NAND U1049 ( .A(n442), .B(n441), .Z(\w0[0][68] ) );
  NAND U1050 ( .A(state[69]), .B(init), .Z(n444) );
  NANDN U1051 ( .A(init), .B(msg[69]), .Z(n443) );
  NAND U1052 ( .A(n444), .B(n443), .Z(\w0[0][69] ) );
  NAND U1053 ( .A(state[6]), .B(init), .Z(n446) );
  NANDN U1054 ( .A(init), .B(msg[6]), .Z(n445) );
  NAND U1055 ( .A(n446), .B(n445), .Z(\w0[0][6] ) );
  NAND U1056 ( .A(state[70]), .B(init), .Z(n448) );
  NANDN U1057 ( .A(init), .B(msg[70]), .Z(n447) );
  NAND U1058 ( .A(n448), .B(n447), .Z(\w0[0][70] ) );
  NAND U1059 ( .A(state[71]), .B(init), .Z(n450) );
  NANDN U1060 ( .A(init), .B(msg[71]), .Z(n449) );
  NAND U1061 ( .A(n450), .B(n449), .Z(\w0[0][71] ) );
  NAND U1062 ( .A(state[72]), .B(init), .Z(n452) );
  NANDN U1063 ( .A(init), .B(msg[72]), .Z(n451) );
  NAND U1064 ( .A(n452), .B(n451), .Z(\w0[0][72] ) );
  NAND U1065 ( .A(state[73]), .B(init), .Z(n454) );
  NANDN U1066 ( .A(init), .B(msg[73]), .Z(n453) );
  NAND U1067 ( .A(n454), .B(n453), .Z(\w0[0][73] ) );
  NAND U1068 ( .A(state[74]), .B(init), .Z(n456) );
  NANDN U1069 ( .A(init), .B(msg[74]), .Z(n455) );
  NAND U1070 ( .A(n456), .B(n455), .Z(\w0[0][74] ) );
  NAND U1071 ( .A(state[75]), .B(init), .Z(n458) );
  NANDN U1072 ( .A(init), .B(msg[75]), .Z(n457) );
  NAND U1073 ( .A(n458), .B(n457), .Z(\w0[0][75] ) );
  NAND U1074 ( .A(state[76]), .B(init), .Z(n460) );
  NANDN U1075 ( .A(init), .B(msg[76]), .Z(n459) );
  NAND U1076 ( .A(n460), .B(n459), .Z(\w0[0][76] ) );
  NAND U1077 ( .A(state[77]), .B(init), .Z(n462) );
  NANDN U1078 ( .A(init), .B(msg[77]), .Z(n461) );
  NAND U1079 ( .A(n462), .B(n461), .Z(\w0[0][77] ) );
  NAND U1080 ( .A(state[78]), .B(init), .Z(n464) );
  NANDN U1081 ( .A(init), .B(msg[78]), .Z(n463) );
  NAND U1082 ( .A(n464), .B(n463), .Z(\w0[0][78] ) );
  NAND U1083 ( .A(state[79]), .B(init), .Z(n466) );
  NANDN U1084 ( .A(init), .B(msg[79]), .Z(n465) );
  NAND U1085 ( .A(n466), .B(n465), .Z(\w0[0][79] ) );
  NAND U1086 ( .A(state[7]), .B(init), .Z(n468) );
  NANDN U1087 ( .A(init), .B(msg[7]), .Z(n467) );
  NAND U1088 ( .A(n468), .B(n467), .Z(\w0[0][7] ) );
  NAND U1089 ( .A(state[80]), .B(init), .Z(n470) );
  NANDN U1090 ( .A(init), .B(msg[80]), .Z(n469) );
  NAND U1091 ( .A(n470), .B(n469), .Z(\w0[0][80] ) );
  NAND U1092 ( .A(state[81]), .B(init), .Z(n472) );
  NANDN U1093 ( .A(init), .B(msg[81]), .Z(n471) );
  NAND U1094 ( .A(n472), .B(n471), .Z(\w0[0][81] ) );
  NAND U1095 ( .A(state[82]), .B(init), .Z(n474) );
  NANDN U1096 ( .A(init), .B(msg[82]), .Z(n473) );
  NAND U1097 ( .A(n474), .B(n473), .Z(\w0[0][82] ) );
  NAND U1098 ( .A(state[83]), .B(init), .Z(n476) );
  NANDN U1099 ( .A(init), .B(msg[83]), .Z(n475) );
  NAND U1100 ( .A(n476), .B(n475), .Z(\w0[0][83] ) );
  NAND U1101 ( .A(state[84]), .B(init), .Z(n478) );
  NANDN U1102 ( .A(init), .B(msg[84]), .Z(n477) );
  NAND U1103 ( .A(n478), .B(n477), .Z(\w0[0][84] ) );
  NAND U1104 ( .A(state[85]), .B(init), .Z(n480) );
  NANDN U1105 ( .A(init), .B(msg[85]), .Z(n479) );
  NAND U1106 ( .A(n480), .B(n479), .Z(\w0[0][85] ) );
  NAND U1107 ( .A(state[86]), .B(init), .Z(n482) );
  NANDN U1108 ( .A(init), .B(msg[86]), .Z(n481) );
  NAND U1109 ( .A(n482), .B(n481), .Z(\w0[0][86] ) );
  NAND U1110 ( .A(state[87]), .B(init), .Z(n484) );
  NANDN U1111 ( .A(init), .B(msg[87]), .Z(n483) );
  NAND U1112 ( .A(n484), .B(n483), .Z(\w0[0][87] ) );
  NAND U1113 ( .A(state[88]), .B(init), .Z(n486) );
  NANDN U1114 ( .A(init), .B(msg[88]), .Z(n485) );
  NAND U1115 ( .A(n486), .B(n485), .Z(\w0[0][88] ) );
  NAND U1116 ( .A(state[89]), .B(init), .Z(n488) );
  NANDN U1117 ( .A(init), .B(msg[89]), .Z(n487) );
  NAND U1118 ( .A(n488), .B(n487), .Z(\w0[0][89] ) );
  NAND U1119 ( .A(state[8]), .B(init), .Z(n490) );
  NANDN U1120 ( .A(init), .B(msg[8]), .Z(n489) );
  NAND U1121 ( .A(n490), .B(n489), .Z(\w0[0][8] ) );
  NAND U1122 ( .A(state[90]), .B(init), .Z(n492) );
  NANDN U1123 ( .A(init), .B(msg[90]), .Z(n491) );
  NAND U1124 ( .A(n492), .B(n491), .Z(\w0[0][90] ) );
  NAND U1125 ( .A(state[91]), .B(init), .Z(n494) );
  NANDN U1126 ( .A(init), .B(msg[91]), .Z(n493) );
  NAND U1127 ( .A(n494), .B(n493), .Z(\w0[0][91] ) );
  NAND U1128 ( .A(state[92]), .B(init), .Z(n496) );
  NANDN U1129 ( .A(init), .B(msg[92]), .Z(n495) );
  NAND U1130 ( .A(n496), .B(n495), .Z(\w0[0][92] ) );
  NAND U1131 ( .A(state[93]), .B(init), .Z(n498) );
  NANDN U1132 ( .A(init), .B(msg[93]), .Z(n497) );
  NAND U1133 ( .A(n498), .B(n497), .Z(\w0[0][93] ) );
  NAND U1134 ( .A(state[94]), .B(init), .Z(n500) );
  NANDN U1135 ( .A(init), .B(msg[94]), .Z(n499) );
  NAND U1136 ( .A(n500), .B(n499), .Z(\w0[0][94] ) );
  NAND U1137 ( .A(state[95]), .B(init), .Z(n502) );
  NANDN U1138 ( .A(init), .B(msg[95]), .Z(n501) );
  NAND U1139 ( .A(n502), .B(n501), .Z(\w0[0][95] ) );
  NAND U1140 ( .A(state[96]), .B(init), .Z(n504) );
  NANDN U1141 ( .A(init), .B(msg[96]), .Z(n503) );
  NAND U1142 ( .A(n504), .B(n503), .Z(\w0[0][96] ) );
  NAND U1143 ( .A(state[97]), .B(init), .Z(n506) );
  NANDN U1144 ( .A(init), .B(msg[97]), .Z(n505) );
  NAND U1145 ( .A(n506), .B(n505), .Z(\w0[0][97] ) );
  NAND U1146 ( .A(state[98]), .B(init), .Z(n508) );
  NANDN U1147 ( .A(init), .B(msg[98]), .Z(n507) );
  NAND U1148 ( .A(n508), .B(n507), .Z(\w0[0][98] ) );
  NAND U1149 ( .A(state[99]), .B(init), .Z(n510) );
  NANDN U1150 ( .A(init), .B(msg[99]), .Z(n509) );
  NAND U1151 ( .A(n510), .B(n509), .Z(\w0[0][99] ) );
  NAND U1152 ( .A(state[9]), .B(init), .Z(n512) );
  NANDN U1153 ( .A(init), .B(msg[9]), .Z(n511) );
  NAND U1154 ( .A(n512), .B(n511), .Z(\w0[0][9] ) );
  XOR U1155 ( .A(key[0]), .B(\w0[0][0] ), .Z(\w1[0][0] ) );
  XOR U1156 ( .A(key[100]), .B(\w0[0][100] ), .Z(\w1[0][100] ) );
  XOR U1157 ( .A(key[101]), .B(\w0[0][101] ), .Z(\w1[0][101] ) );
  XOR U1158 ( .A(key[102]), .B(\w0[0][102] ), .Z(\w1[0][102] ) );
  XOR U1159 ( .A(key[103]), .B(\w0[0][103] ), .Z(\w1[0][103] ) );
  XOR U1160 ( .A(key[104]), .B(\w0[0][104] ), .Z(\w1[0][104] ) );
  XOR U1161 ( .A(key[105]), .B(\w0[0][105] ), .Z(\w1[0][105] ) );
  XOR U1162 ( .A(key[106]), .B(\w0[0][106] ), .Z(\w1[0][106] ) );
  XOR U1163 ( .A(key[107]), .B(\w0[0][107] ), .Z(\w1[0][107] ) );
  XOR U1164 ( .A(key[108]), .B(\w0[0][108] ), .Z(\w1[0][108] ) );
  XOR U1165 ( .A(key[109]), .B(\w0[0][109] ), .Z(\w1[0][109] ) );
  XOR U1166 ( .A(key[10]), .B(\w0[0][10] ), .Z(\w1[0][10] ) );
  XOR U1167 ( .A(key[110]), .B(\w0[0][110] ), .Z(\w1[0][110] ) );
  XOR U1168 ( .A(key[111]), .B(\w0[0][111] ), .Z(\w1[0][111] ) );
  XOR U1169 ( .A(key[112]), .B(\w0[0][112] ), .Z(\w1[0][112] ) );
  XOR U1170 ( .A(key[113]), .B(\w0[0][113] ), .Z(\w1[0][113] ) );
  XOR U1171 ( .A(key[114]), .B(\w0[0][114] ), .Z(\w1[0][114] ) );
  XOR U1172 ( .A(key[115]), .B(\w0[0][115] ), .Z(\w1[0][115] ) );
  XOR U1173 ( .A(key[116]), .B(\w0[0][116] ), .Z(\w1[0][116] ) );
  XOR U1174 ( .A(key[117]), .B(\w0[0][117] ), .Z(\w1[0][117] ) );
  XOR U1175 ( .A(key[118]), .B(\w0[0][118] ), .Z(\w1[0][118] ) );
  XOR U1176 ( .A(key[119]), .B(\w0[0][119] ), .Z(\w1[0][119] ) );
  XOR U1177 ( .A(key[11]), .B(\w0[0][11] ), .Z(\w1[0][11] ) );
  XOR U1178 ( .A(key[120]), .B(\w0[0][120] ), .Z(\w1[0][120] ) );
  XOR U1179 ( .A(key[121]), .B(\w0[0][121] ), .Z(\w1[0][121] ) );
  XOR U1180 ( .A(key[122]), .B(\w0[0][122] ), .Z(\w1[0][122] ) );
  XOR U1181 ( .A(key[123]), .B(\w0[0][123] ), .Z(\w1[0][123] ) );
  XOR U1182 ( .A(key[124]), .B(\w0[0][124] ), .Z(\w1[0][124] ) );
  XOR U1183 ( .A(key[125]), .B(\w0[0][125] ), .Z(\w1[0][125] ) );
  XOR U1184 ( .A(key[126]), .B(\w0[0][126] ), .Z(\w1[0][126] ) );
  XOR U1185 ( .A(key[127]), .B(\w0[0][127] ), .Z(\w1[0][127] ) );
  XOR U1186 ( .A(key[12]), .B(\w0[0][12] ), .Z(\w1[0][12] ) );
  XOR U1187 ( .A(key[13]), .B(\w0[0][13] ), .Z(\w1[0][13] ) );
  XOR U1188 ( .A(key[14]), .B(\w0[0][14] ), .Z(\w1[0][14] ) );
  XOR U1189 ( .A(key[15]), .B(\w0[0][15] ), .Z(\w1[0][15] ) );
  XOR U1190 ( .A(key[16]), .B(\w0[0][16] ), .Z(\w1[0][16] ) );
  XOR U1191 ( .A(key[17]), .B(\w0[0][17] ), .Z(\w1[0][17] ) );
  XOR U1192 ( .A(key[18]), .B(\w0[0][18] ), .Z(\w1[0][18] ) );
  XOR U1193 ( .A(key[19]), .B(\w0[0][19] ), .Z(\w1[0][19] ) );
  XOR U1194 ( .A(key[1]), .B(\w0[0][1] ), .Z(\w1[0][1] ) );
  XOR U1195 ( .A(key[20]), .B(\w0[0][20] ), .Z(\w1[0][20] ) );
  XOR U1196 ( .A(key[21]), .B(\w0[0][21] ), .Z(\w1[0][21] ) );
  XOR U1197 ( .A(key[22]), .B(\w0[0][22] ), .Z(\w1[0][22] ) );
  XOR U1198 ( .A(key[23]), .B(\w0[0][23] ), .Z(\w1[0][23] ) );
  XOR U1199 ( .A(key[24]), .B(\w0[0][24] ), .Z(\w1[0][24] ) );
  XOR U1200 ( .A(key[25]), .B(\w0[0][25] ), .Z(\w1[0][25] ) );
  XOR U1201 ( .A(key[26]), .B(\w0[0][26] ), .Z(\w1[0][26] ) );
  XOR U1202 ( .A(key[27]), .B(\w0[0][27] ), .Z(\w1[0][27] ) );
  XOR U1203 ( .A(key[28]), .B(\w0[0][28] ), .Z(\w1[0][28] ) );
  XOR U1204 ( .A(key[29]), .B(\w0[0][29] ), .Z(\w1[0][29] ) );
  XOR U1205 ( .A(key[2]), .B(\w0[0][2] ), .Z(\w1[0][2] ) );
  XOR U1206 ( .A(key[30]), .B(\w0[0][30] ), .Z(\w1[0][30] ) );
  XOR U1207 ( .A(key[31]), .B(\w0[0][31] ), .Z(\w1[0][31] ) );
  XOR U1208 ( .A(key[32]), .B(\w0[0][32] ), .Z(\w1[0][32] ) );
  XOR U1209 ( .A(key[33]), .B(\w0[0][33] ), .Z(\w1[0][33] ) );
  XOR U1210 ( .A(key[34]), .B(\w0[0][34] ), .Z(\w1[0][34] ) );
  XOR U1211 ( .A(key[35]), .B(\w0[0][35] ), .Z(\w1[0][35] ) );
  XOR U1212 ( .A(key[36]), .B(\w0[0][36] ), .Z(\w1[0][36] ) );
  XOR U1213 ( .A(key[37]), .B(\w0[0][37] ), .Z(\w1[0][37] ) );
  XOR U1214 ( .A(key[38]), .B(\w0[0][38] ), .Z(\w1[0][38] ) );
  XOR U1215 ( .A(key[39]), .B(\w0[0][39] ), .Z(\w1[0][39] ) );
  XOR U1216 ( .A(key[3]), .B(\w0[0][3] ), .Z(\w1[0][3] ) );
  XOR U1217 ( .A(key[40]), .B(\w0[0][40] ), .Z(\w1[0][40] ) );
  XOR U1218 ( .A(key[41]), .B(\w0[0][41] ), .Z(\w1[0][41] ) );
  XOR U1219 ( .A(key[42]), .B(\w0[0][42] ), .Z(\w1[0][42] ) );
  XOR U1220 ( .A(key[43]), .B(\w0[0][43] ), .Z(\w1[0][43] ) );
  XOR U1221 ( .A(key[44]), .B(\w0[0][44] ), .Z(\w1[0][44] ) );
  XOR U1222 ( .A(key[45]), .B(\w0[0][45] ), .Z(\w1[0][45] ) );
  XOR U1223 ( .A(key[46]), .B(\w0[0][46] ), .Z(\w1[0][46] ) );
  XOR U1224 ( .A(key[47]), .B(\w0[0][47] ), .Z(\w1[0][47] ) );
  XOR U1225 ( .A(key[48]), .B(\w0[0][48] ), .Z(\w1[0][48] ) );
  XOR U1226 ( .A(key[49]), .B(\w0[0][49] ), .Z(\w1[0][49] ) );
  XOR U1227 ( .A(key[4]), .B(\w0[0][4] ), .Z(\w1[0][4] ) );
  XOR U1228 ( .A(key[50]), .B(\w0[0][50] ), .Z(\w1[0][50] ) );
  XOR U1229 ( .A(key[51]), .B(\w0[0][51] ), .Z(\w1[0][51] ) );
  XOR U1230 ( .A(key[52]), .B(\w0[0][52] ), .Z(\w1[0][52] ) );
  XOR U1231 ( .A(key[53]), .B(\w0[0][53] ), .Z(\w1[0][53] ) );
  XOR U1232 ( .A(key[54]), .B(\w0[0][54] ), .Z(\w1[0][54] ) );
  XOR U1233 ( .A(key[55]), .B(\w0[0][55] ), .Z(\w1[0][55] ) );
  XOR U1234 ( .A(key[56]), .B(\w0[0][56] ), .Z(\w1[0][56] ) );
  XOR U1235 ( .A(key[57]), .B(\w0[0][57] ), .Z(\w1[0][57] ) );
  XOR U1236 ( .A(key[58]), .B(\w0[0][58] ), .Z(\w1[0][58] ) );
  XOR U1237 ( .A(key[59]), .B(\w0[0][59] ), .Z(\w1[0][59] ) );
  XOR U1238 ( .A(key[5]), .B(\w0[0][5] ), .Z(\w1[0][5] ) );
  XOR U1239 ( .A(key[60]), .B(\w0[0][60] ), .Z(\w1[0][60] ) );
  XOR U1240 ( .A(key[61]), .B(\w0[0][61] ), .Z(\w1[0][61] ) );
  XOR U1241 ( .A(key[62]), .B(\w0[0][62] ), .Z(\w1[0][62] ) );
  XOR U1242 ( .A(key[63]), .B(\w0[0][63] ), .Z(\w1[0][63] ) );
  XOR U1243 ( .A(key[64]), .B(\w0[0][64] ), .Z(\w1[0][64] ) );
  XOR U1244 ( .A(key[65]), .B(\w0[0][65] ), .Z(\w1[0][65] ) );
  XOR U1245 ( .A(key[66]), .B(\w0[0][66] ), .Z(\w1[0][66] ) );
  XOR U1246 ( .A(key[67]), .B(\w0[0][67] ), .Z(\w1[0][67] ) );
  XOR U1247 ( .A(key[68]), .B(\w0[0][68] ), .Z(\w1[0][68] ) );
  XOR U1248 ( .A(key[69]), .B(\w0[0][69] ), .Z(\w1[0][69] ) );
  XOR U1249 ( .A(key[6]), .B(\w0[0][6] ), .Z(\w1[0][6] ) );
  XOR U1250 ( .A(key[70]), .B(\w0[0][70] ), .Z(\w1[0][70] ) );
  XOR U1251 ( .A(key[71]), .B(\w0[0][71] ), .Z(\w1[0][71] ) );
  XOR U1252 ( .A(key[72]), .B(\w0[0][72] ), .Z(\w1[0][72] ) );
  XOR U1253 ( .A(key[73]), .B(\w0[0][73] ), .Z(\w1[0][73] ) );
  XOR U1254 ( .A(key[74]), .B(\w0[0][74] ), .Z(\w1[0][74] ) );
  XOR U1255 ( .A(key[75]), .B(\w0[0][75] ), .Z(\w1[0][75] ) );
  XOR U1256 ( .A(key[76]), .B(\w0[0][76] ), .Z(\w1[0][76] ) );
  XOR U1257 ( .A(key[77]), .B(\w0[0][77] ), .Z(\w1[0][77] ) );
  XOR U1258 ( .A(key[78]), .B(\w0[0][78] ), .Z(\w1[0][78] ) );
  XOR U1259 ( .A(key[79]), .B(\w0[0][79] ), .Z(\w1[0][79] ) );
  XOR U1260 ( .A(key[7]), .B(\w0[0][7] ), .Z(\w1[0][7] ) );
  XOR U1261 ( .A(key[80]), .B(\w0[0][80] ), .Z(\w1[0][80] ) );
  XOR U1262 ( .A(key[81]), .B(\w0[0][81] ), .Z(\w1[0][81] ) );
  XOR U1263 ( .A(key[82]), .B(\w0[0][82] ), .Z(\w1[0][82] ) );
  XOR U1264 ( .A(key[83]), .B(\w0[0][83] ), .Z(\w1[0][83] ) );
  XOR U1265 ( .A(key[84]), .B(\w0[0][84] ), .Z(\w1[0][84] ) );
  XOR U1266 ( .A(key[85]), .B(\w0[0][85] ), .Z(\w1[0][85] ) );
  XOR U1267 ( .A(key[86]), .B(\w0[0][86] ), .Z(\w1[0][86] ) );
  XOR U1268 ( .A(key[87]), .B(\w0[0][87] ), .Z(\w1[0][87] ) );
  XOR U1269 ( .A(key[88]), .B(\w0[0][88] ), .Z(\w1[0][88] ) );
  XOR U1270 ( .A(key[89]), .B(\w0[0][89] ), .Z(\w1[0][89] ) );
  XOR U1271 ( .A(key[8]), .B(\w0[0][8] ), .Z(\w1[0][8] ) );
  XOR U1272 ( .A(key[90]), .B(\w0[0][90] ), .Z(\w1[0][90] ) );
  XOR U1273 ( .A(key[91]), .B(\w0[0][91] ), .Z(\w1[0][91] ) );
  XOR U1274 ( .A(key[92]), .B(\w0[0][92] ), .Z(\w1[0][92] ) );
  XOR U1275 ( .A(key[93]), .B(\w0[0][93] ), .Z(\w1[0][93] ) );
  XOR U1276 ( .A(key[94]), .B(\w0[0][94] ), .Z(\w1[0][94] ) );
  XOR U1277 ( .A(key[95]), .B(\w0[0][95] ), .Z(\w1[0][95] ) );
  XOR U1278 ( .A(key[96]), .B(\w0[0][96] ), .Z(\w1[0][96] ) );
  XOR U1279 ( .A(key[97]), .B(\w0[0][97] ), .Z(\w1[0][97] ) );
  XOR U1280 ( .A(key[98]), .B(\w0[0][98] ), .Z(\w1[0][98] ) );
  XOR U1281 ( .A(key[99]), .B(\w0[0][99] ), .Z(\w1[0][99] ) );
  XOR U1282 ( .A(key[9]), .B(\w0[0][9] ), .Z(\w1[0][9] ) );
endmodule

