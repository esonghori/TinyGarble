
module hamming_N16000_CC32 ( clk, rst, x, y, o );
  input [499:0] x;
  input [499:0] y;
  output [13:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015;
  wire   [13:0] oglobal;

  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  XNOR U503 ( .A(n2717), .B(n2716), .Z(n2718) );
  XOR U504 ( .A(n2731), .B(n2730), .Z(n2700) );
  XNOR U505 ( .A(n1566), .B(n1565), .Z(n1567) );
  XNOR U506 ( .A(n2882), .B(n2881), .Z(n2870) );
  XNOR U507 ( .A(n2970), .B(n2969), .Z(n2971) );
  NAND U508 ( .A(n2278), .B(n2279), .Z(n1) );
  XOR U509 ( .A(n2278), .B(n2279), .Z(n2) );
  NANDN U510 ( .A(n2277), .B(n2), .Z(n3) );
  NAND U511 ( .A(n1), .B(n3), .Z(n2547) );
  XNOR U512 ( .A(n2656), .B(n2655), .Z(n2671) );
  XNOR U513 ( .A(n2847), .B(n2846), .Z(n2921) );
  XNOR U514 ( .A(n2129), .B(n2128), .Z(n2131) );
  XNOR U515 ( .A(n2063), .B(oglobal[1]), .Z(n2064) );
  XNOR U516 ( .A(n1668), .B(n1667), .Z(n1670) );
  XNOR U517 ( .A(n1674), .B(n1673), .Z(n1676) );
  XNOR U518 ( .A(n2475), .B(n2474), .Z(n2476) );
  XNOR U519 ( .A(n2469), .B(n2468), .Z(n2470) );
  XNOR U520 ( .A(n2348), .B(n2347), .Z(n2350) );
  XNOR U521 ( .A(n2863), .B(n2862), .Z(n2865) );
  XNOR U522 ( .A(n2875), .B(n2874), .Z(n2876) );
  XNOR U523 ( .A(n2529), .B(n2528), .Z(n2531) );
  XOR U524 ( .A(n1790), .B(n1789), .Z(n2266) );
  XNOR U525 ( .A(n2888), .B(n2887), .Z(n2918) );
  XNOR U526 ( .A(n2972), .B(n2971), .Z(n2952) );
  XOR U527 ( .A(n1562), .B(n1561), .Z(n2260) );
  XNOR U528 ( .A(n2983), .B(n2982), .Z(n2984) );
  NAND U529 ( .A(n2671), .B(n2673), .Z(n4) );
  XOR U530 ( .A(n2671), .B(n2673), .Z(n5) );
  NAND U531 ( .A(n5), .B(n2672), .Z(n6) );
  NAND U532 ( .A(n4), .B(n6), .Z(n2922) );
  XNOR U533 ( .A(n148), .B(n147), .Z(n149) );
  XNOR U534 ( .A(n385), .B(n384), .Z(n386) );
  XNOR U535 ( .A(n1608), .B(n1607), .Z(n1610) );
  XNOR U536 ( .A(n2117), .B(n2116), .Z(n2119) );
  XNOR U537 ( .A(n2189), .B(n2188), .Z(n2191) );
  XNOR U538 ( .A(n2195), .B(n2194), .Z(n2197) );
  XNOR U539 ( .A(n1656), .B(n1655), .Z(n1658) );
  XNOR U540 ( .A(n1746), .B(n1745), .Z(n1748) );
  XNOR U541 ( .A(n2147), .B(n2146), .Z(n2149) );
  XNOR U542 ( .A(n1910), .B(n1909), .Z(n1983) );
  XNOR U543 ( .A(n2396), .B(n2395), .Z(n2397) );
  XNOR U544 ( .A(n2390), .B(n2389), .Z(n2391) );
  XNOR U545 ( .A(n2451), .B(n2450), .Z(n2452) );
  XNOR U546 ( .A(n2457), .B(n2456), .Z(n2458) );
  XNOR U547 ( .A(n2483), .B(n2482), .Z(n2446) );
  XNOR U548 ( .A(n2402), .B(n2401), .Z(n2403) );
  XNOR U549 ( .A(n2336), .B(n2335), .Z(n2337) );
  XNOR U550 ( .A(n2324), .B(n2323), .Z(n2325) );
  XOR U551 ( .A(n2471), .B(n2470), .Z(n2464) );
  NAND U552 ( .A(n2019), .B(n2020), .Z(n7) );
  XOR U553 ( .A(n2019), .B(n2020), .Z(n8) );
  NANDN U554 ( .A(n2018), .B(n8), .Z(n9) );
  NAND U555 ( .A(n7), .B(n9), .Z(n2510) );
  NAND U556 ( .A(n1971), .B(n1972), .Z(n10) );
  XOR U557 ( .A(n1971), .B(n1972), .Z(n11) );
  NANDN U558 ( .A(n1970), .B(n11), .Z(n12) );
  NAND U559 ( .A(n10), .B(n12), .Z(n2499) );
  NAND U560 ( .A(n1953), .B(n1954), .Z(n13) );
  XOR U561 ( .A(n1953), .B(n1954), .Z(n14) );
  NANDN U562 ( .A(n1952), .B(n14), .Z(n15) );
  NAND U563 ( .A(n13), .B(n15), .Z(n2493) );
  XNOR U564 ( .A(n2417), .B(n2416), .Z(n2486) );
  XNOR U565 ( .A(n2735), .B(n2734), .Z(n2736) );
  XNOR U566 ( .A(n2705), .B(n2704), .Z(n2707) );
  XNOR U567 ( .A(n2772), .B(n2771), .Z(n2773) );
  XNOR U568 ( .A(n2778), .B(n2777), .Z(n2779) );
  XNOR U569 ( .A(n2687), .B(n2686), .Z(n2689) );
  XNOR U570 ( .A(n2681), .B(n2680), .Z(n2682) );
  XNOR U571 ( .A(n2869), .B(n2868), .Z(n2871) );
  XNOR U572 ( .A(n2886), .B(n2885), .Z(n2887) );
  XNOR U573 ( .A(n2808), .B(n2807), .Z(n2810) );
  XNOR U574 ( .A(n2916), .B(n2915), .Z(n2917) );
  XNOR U575 ( .A(n2953), .B(n2952), .Z(n2954) );
  XNOR U576 ( .A(n2557), .B(n2556), .Z(n2558) );
  XNOR U577 ( .A(n2666), .B(n2665), .Z(n2667) );
  NANDN U578 ( .A(n2254), .B(n2257), .Z(n16) );
  OR U579 ( .A(n2257), .B(n2256), .Z(n17) );
  NANDN U580 ( .A(n2255), .B(n17), .Z(n18) );
  NAND U581 ( .A(n16), .B(n18), .Z(n2542) );
  XNOR U582 ( .A(n2553), .B(n2552), .Z(n2548) );
  NAND U583 ( .A(n2921), .B(n2923), .Z(n19) );
  XOR U584 ( .A(n2921), .B(n2923), .Z(n20) );
  NAND U585 ( .A(n20), .B(n2922), .Z(n21) );
  NAND U586 ( .A(n19), .B(n21), .Z(n2938) );
  NAND U587 ( .A(n3007), .B(n3008), .Z(n22) );
  XOR U588 ( .A(n3007), .B(n3008), .Z(n23) );
  NAND U589 ( .A(n23), .B(n3006), .Z(n24) );
  NAND U590 ( .A(n22), .B(n24), .Z(n3010) );
  XNOR U591 ( .A(n715), .B(n714), .Z(n716) );
  XNOR U592 ( .A(n721), .B(n720), .Z(n722) );
  XNOR U593 ( .A(n703), .B(n702), .Z(n704) );
  XNOR U594 ( .A(n619), .B(n618), .Z(n620) );
  XNOR U595 ( .A(n1510), .B(n1509), .Z(n1511) );
  XNOR U596 ( .A(n1516), .B(n1515), .Z(n1517) );
  XNOR U597 ( .A(n1124), .B(n1123), .Z(n1125) );
  XNOR U598 ( .A(n1130), .B(n1129), .Z(n1131) );
  XNOR U599 ( .A(n583), .B(n582), .Z(n584) );
  XNOR U600 ( .A(n595), .B(n594), .Z(n596) );
  XNOR U601 ( .A(n1444), .B(n1443), .Z(n1445) );
  XNOR U602 ( .A(n1456), .B(n1455), .Z(n1457) );
  XNOR U603 ( .A(n99), .B(n98), .Z(n100) );
  XNOR U604 ( .A(n649), .B(n648), .Z(n650) );
  XNOR U605 ( .A(n655), .B(n654), .Z(n656) );
  XNOR U606 ( .A(n914), .B(n913), .Z(n915) );
  XNOR U607 ( .A(n124), .B(n123), .Z(n125) );
  XNOR U608 ( .A(n361), .B(n360), .Z(n362) );
  XNOR U609 ( .A(n697), .B(n696), .Z(n698) );
  XNOR U610 ( .A(n691), .B(n690), .Z(n692) );
  XNOR U611 ( .A(n1534), .B(n1533), .Z(n1535) );
  XNOR U612 ( .A(n1528), .B(n1527), .Z(n1529) );
  XNOR U613 ( .A(n631), .B(n630), .Z(n632) );
  XNOR U614 ( .A(n637), .B(n636), .Z(n638) );
  XNOR U615 ( .A(n475), .B(n474), .Z(n476) );
  XNOR U616 ( .A(n1142), .B(n1141), .Z(n1143) );
  XNOR U617 ( .A(n613), .B(n612), .Z(n614) );
  XNOR U618 ( .A(n1450), .B(n1449), .Z(n1451) );
  XNOR U619 ( .A(n1522), .B(n1521), .Z(n1523) );
  XNOR U620 ( .A(n1614), .B(n1613), .Z(n1616) );
  XNOR U621 ( .A(n2123), .B(n2122), .Z(n2125) );
  XNOR U622 ( .A(n2183), .B(n2182), .Z(n2185) );
  XNOR U623 ( .A(n2040), .B(n2039), .Z(n2042) );
  XNOR U624 ( .A(n1782), .B(n1781), .Z(n1784) );
  XNOR U625 ( .A(n1734), .B(n1733), .Z(n1736) );
  XNOR U626 ( .A(n2165), .B(n2164), .Z(n2167) );
  XNOR U627 ( .A(n2159), .B(n2158), .Z(n2161) );
  XNOR U628 ( .A(n2171), .B(n2170), .Z(n2173) );
  XNOR U629 ( .A(n2075), .B(n2074), .Z(n2077) );
  XNOR U630 ( .A(n2213), .B(n2212), .Z(n2215) );
  XNOR U631 ( .A(n2141), .B(n2140), .Z(n2143) );
  XNOR U632 ( .A(n1908), .B(n1907), .Z(n1909) );
  XNOR U633 ( .A(n1540), .B(n1539), .Z(n1541) );
  XNOR U634 ( .A(n93), .B(n92), .Z(n94) );
  XNOR U635 ( .A(n215), .B(n214), .Z(n216) );
  XNOR U636 ( .A(n130), .B(n129), .Z(n131) );
  XNOR U637 ( .A(n511), .B(n510), .Z(n512) );
  XNOR U638 ( .A(n908), .B(n907), .Z(n909) );
  XNOR U639 ( .A(n920), .B(n919), .Z(n921) );
  XNOR U640 ( .A(n2065), .B(n2064), .Z(n1939) );
  XNOR U641 ( .A(n2384), .B(n2383), .Z(n2385) );
  XNOR U642 ( .A(n2445), .B(n2444), .Z(n2447) );
  XNOR U643 ( .A(n2481), .B(n2480), .Z(n2482) );
  XNOR U644 ( .A(n2408), .B(n2407), .Z(n2409) );
  XNOR U645 ( .A(n2372), .B(n2371), .Z(n2373) );
  XNOR U646 ( .A(n2378), .B(n2377), .Z(n2379) );
  XOR U647 ( .A(n2404), .B(n2403), .Z(n2575) );
  XOR U648 ( .A(n2392), .B(n2391), .Z(n2422) );
  XOR U649 ( .A(n2477), .B(n2476), .Z(n2636) );
  XOR U650 ( .A(n2398), .B(n2397), .Z(n2642) );
  XNOR U651 ( .A(n2415), .B(n2414), .Z(n2416) );
  XNOR U652 ( .A(n2330), .B(n2329), .Z(n2332) );
  NAND U653 ( .A(n2016), .B(n2017), .Z(n25) );
  XOR U654 ( .A(n2016), .B(n2017), .Z(n26) );
  NANDN U655 ( .A(n2015), .B(n26), .Z(n27) );
  NAND U656 ( .A(n25), .B(n27), .Z(n2511) );
  NAND U657 ( .A(n1974), .B(n1975), .Z(n28) );
  XOR U658 ( .A(n1974), .B(n1975), .Z(n29) );
  NANDN U659 ( .A(n1973), .B(n29), .Z(n30) );
  NAND U660 ( .A(n28), .B(n30), .Z(n2498) );
  NAND U661 ( .A(n1956), .B(n1957), .Z(n31) );
  XOR U662 ( .A(n1956), .B(n1957), .Z(n32) );
  NANDN U663 ( .A(n1955), .B(n32), .Z(n33) );
  NAND U664 ( .A(n31), .B(n33), .Z(n2492) );
  XNOR U665 ( .A(n2326), .B(n2325), .Z(n2288) );
  NAND U666 ( .A(n1950), .B(n1951), .Z(n34) );
  XOR U667 ( .A(n1950), .B(n1951), .Z(n35) );
  NANDN U668 ( .A(n1949), .B(n35), .Z(n36) );
  NAND U669 ( .A(n34), .B(n36), .Z(n2342) );
  XNOR U670 ( .A(n2338), .B(n2337), .Z(n2488) );
  XNOR U671 ( .A(n2729), .B(n2728), .Z(n2730) );
  XNOR U672 ( .A(n2742), .B(n2741), .Z(n2743) );
  XNOR U673 ( .A(n2699), .B(n2698), .Z(n2701) );
  XOR U674 ( .A(n2006), .B(n2007), .Z(n37) );
  NANDN U675 ( .A(n2008), .B(n37), .Z(n38) );
  NAND U676 ( .A(n2006), .B(n2007), .Z(n39) );
  AND U677 ( .A(n38), .B(n39), .Z(n2360) );
  XOR U678 ( .A(n2354), .B(n2353), .Z(n2356) );
  XNOR U679 ( .A(n2683), .B(n2682), .Z(n2759) );
  XNOR U680 ( .A(n2780), .B(n2779), .Z(n2756) );
  XOR U681 ( .A(n2877), .B(n2876), .Z(n2864) );
  XNOR U682 ( .A(n2880), .B(oglobal[4]), .Z(n2881) );
  XNOR U683 ( .A(n2892), .B(n2891), .Z(n2893) );
  XNOR U684 ( .A(n2898), .B(n2897), .Z(n2899) );
  XNOR U685 ( .A(n1902), .B(n1901), .Z(n1903) );
  XNOR U686 ( .A(n1560), .B(n1559), .Z(n1561) );
  XOR U687 ( .A(n1568), .B(n1567), .Z(n2268) );
  XNOR U688 ( .A(n2959), .B(n2958), .Z(n2960) );
  XNOR U689 ( .A(n2918), .B(n2917), .Z(n2853) );
  XNOR U690 ( .A(n2841), .B(n2840), .Z(n2844) );
  XNOR U691 ( .A(n2668), .B(n2667), .Z(n2656) );
  XOR U692 ( .A(n2985), .B(n2984), .Z(n2977) );
  NAND U693 ( .A(n2548), .B(n2549), .Z(n40) );
  XOR U694 ( .A(n2548), .B(n2549), .Z(n41) );
  NANDN U695 ( .A(n2547), .B(n41), .Z(n42) );
  NAND U696 ( .A(n40), .B(n42), .Z(n2672) );
  NAND U697 ( .A(n2937), .B(n2939), .Z(n43) );
  XOR U698 ( .A(n2937), .B(n2939), .Z(n44) );
  NAND U699 ( .A(n44), .B(n2938), .Z(n45) );
  NAND U700 ( .A(n43), .B(n45), .Z(n2994) );
  XOR U701 ( .A(oglobal[8]), .B(n3010), .Z(n46) );
  NANDN U702 ( .A(n3011), .B(n46), .Z(n47) );
  NAND U703 ( .A(oglobal[8]), .B(n3010), .Z(n48) );
  AND U704 ( .A(n47), .B(n48), .Z(n3012) );
  NAND U705 ( .A(n3015), .B(oglobal[12]), .Z(n49) );
  XNOR U706 ( .A(oglobal[13]), .B(n49), .Z(o[13]) );
  XOR U707 ( .A(x[190]), .B(y[190]), .Z(n1042) );
  XOR U708 ( .A(x[163]), .B(y[163]), .Z(n1039) );
  XOR U709 ( .A(x[192]), .B(y[192]), .Z(n1040) );
  XOR U710 ( .A(n1039), .B(n1040), .Z(n1041) );
  XNOR U711 ( .A(n1042), .B(n1041), .Z(n1247) );
  XOR U712 ( .A(x[186]), .B(y[186]), .Z(n693) );
  XOR U713 ( .A(x[188]), .B(y[188]), .Z(n690) );
  XNOR U714 ( .A(x[469]), .B(y[469]), .Z(n691) );
  XNOR U715 ( .A(n693), .B(n692), .Z(n1245) );
  XOR U716 ( .A(x[178]), .B(y[178]), .Z(n699) );
  XOR U717 ( .A(x[167]), .B(y[167]), .Z(n696) );
  XNOR U718 ( .A(x[182]), .B(y[182]), .Z(n697) );
  XNOR U719 ( .A(n699), .B(n698), .Z(n1244) );
  XOR U720 ( .A(n1245), .B(n1244), .Z(n1246) );
  XOR U721 ( .A(n1247), .B(n1246), .Z(n263) );
  XOR U722 ( .A(x[174]), .B(y[174]), .Z(n687) );
  XOR U723 ( .A(x[176]), .B(y[176]), .Z(n684) );
  XOR U724 ( .A(x[467]), .B(y[467]), .Z(n685) );
  XOR U725 ( .A(n684), .B(n685), .Z(n686) );
  XNOR U726 ( .A(n687), .B(n686), .Z(n1314) );
  XOR U727 ( .A(x[170]), .B(y[170]), .Z(n675) );
  XOR U728 ( .A(x[171]), .B(y[171]), .Z(n672) );
  XOR U729 ( .A(x[172]), .B(y[172]), .Z(n673) );
  XOR U730 ( .A(n672), .B(n673), .Z(n674) );
  XNOR U731 ( .A(n675), .B(n674), .Z(n1312) );
  XOR U732 ( .A(x[164]), .B(y[164]), .Z(n681) );
  XOR U733 ( .A(x[168]), .B(y[168]), .Z(n678) );
  XOR U734 ( .A(x[465]), .B(y[465]), .Z(n679) );
  XOR U735 ( .A(n678), .B(n679), .Z(n680) );
  XNOR U736 ( .A(n681), .B(n680), .Z(n1311) );
  XOR U737 ( .A(n1312), .B(n1311), .Z(n1313) );
  XOR U738 ( .A(n1314), .B(n1313), .Z(n262) );
  XOR U739 ( .A(n263), .B(n262), .Z(n265) );
  XOR U740 ( .A(x[158]), .B(y[158]), .Z(n946) );
  XOR U741 ( .A(x[160]), .B(y[160]), .Z(n943) );
  XOR U742 ( .A(x[175]), .B(y[175]), .Z(n944) );
  XOR U743 ( .A(n943), .B(n944), .Z(n945) );
  XNOR U744 ( .A(n946), .B(n945), .Z(n1198) );
  XOR U745 ( .A(x[154]), .B(y[154]), .Z(n934) );
  XOR U746 ( .A(x[156]), .B(y[156]), .Z(n931) );
  XOR U747 ( .A(x[463]), .B(y[463]), .Z(n932) );
  XOR U748 ( .A(n931), .B(n932), .Z(n933) );
  XNOR U749 ( .A(n934), .B(n933), .Z(n1196) );
  XOR U750 ( .A(x[150]), .B(y[150]), .Z(n940) );
  XOR U751 ( .A(x[152]), .B(y[152]), .Z(n937) );
  XOR U752 ( .A(x[179]), .B(y[179]), .Z(n938) );
  XOR U753 ( .A(n937), .B(n938), .Z(n939) );
  XNOR U754 ( .A(n940), .B(n939), .Z(n1195) );
  XOR U755 ( .A(n1196), .B(n1195), .Z(n1197) );
  XOR U756 ( .A(n1198), .B(n1197), .Z(n264) );
  XNOR U757 ( .A(n265), .B(n264), .Z(n1174) );
  XOR U758 ( .A(x[142]), .B(y[142]), .Z(n1500) );
  XOR U759 ( .A(x[146]), .B(y[146]), .Z(n1497) );
  XOR U760 ( .A(x[461]), .B(y[461]), .Z(n1498) );
  XOR U761 ( .A(n1497), .B(n1498), .Z(n1499) );
  XNOR U762 ( .A(n1500), .B(n1499), .Z(n1271) );
  XOR U763 ( .A(x[138]), .B(y[138]), .Z(n1488) );
  XOR U764 ( .A(x[140]), .B(y[140]), .Z(n1485) );
  XOR U765 ( .A(x[183]), .B(y[183]), .Z(n1486) );
  XOR U766 ( .A(n1485), .B(n1486), .Z(n1487) );
  XNOR U767 ( .A(n1488), .B(n1487), .Z(n1269) );
  XOR U768 ( .A(x[134]), .B(y[134]), .Z(n1494) );
  XOR U769 ( .A(x[136]), .B(y[136]), .Z(n1491) );
  XOR U770 ( .A(x[459]), .B(y[459]), .Z(n1492) );
  XOR U771 ( .A(n1491), .B(n1492), .Z(n1493) );
  XNOR U772 ( .A(n1494), .B(n1493), .Z(n1268) );
  XOR U773 ( .A(n1269), .B(n1268), .Z(n1270) );
  XOR U774 ( .A(n1271), .B(n1270), .Z(n57) );
  XOR U775 ( .A(x[128]), .B(y[128]), .Z(n1440) );
  XOR U776 ( .A(x[132]), .B(y[132]), .Z(n1437) );
  XOR U777 ( .A(x[187]), .B(y[187]), .Z(n1438) );
  XOR U778 ( .A(n1437), .B(n1438), .Z(n1439) );
  XNOR U779 ( .A(n1440), .B(n1439), .Z(n1385) );
  XOR U780 ( .A(x[122]), .B(y[122]), .Z(n1428) );
  XOR U781 ( .A(x[124]), .B(y[124]), .Z(n1425) );
  XOR U782 ( .A(x[457]), .B(y[457]), .Z(n1426) );
  XOR U783 ( .A(n1425), .B(n1426), .Z(n1427) );
  XNOR U784 ( .A(n1428), .B(n1427), .Z(n1383) );
  XOR U785 ( .A(x[118]), .B(y[118]), .Z(n1434) );
  XOR U786 ( .A(x[120]), .B(y[120]), .Z(n1431) );
  XOR U787 ( .A(x[191]), .B(y[191]), .Z(n1432) );
  XOR U788 ( .A(n1431), .B(n1432), .Z(n1433) );
  XNOR U789 ( .A(n1434), .B(n1433), .Z(n1382) );
  XOR U790 ( .A(n1383), .B(n1382), .Z(n1384) );
  XOR U791 ( .A(n1385), .B(n1384), .Z(n56) );
  XOR U792 ( .A(n57), .B(n56), .Z(n59) );
  XOR U793 ( .A(x[114]), .B(y[114]), .Z(n826) );
  XOR U794 ( .A(x[116]), .B(y[116]), .Z(n823) );
  XOR U795 ( .A(x[455]), .B(y[455]), .Z(n824) );
  XOR U796 ( .A(n823), .B(n824), .Z(n825) );
  XNOR U797 ( .A(n826), .B(n825), .Z(n1421) );
  XOR U798 ( .A(x[106]), .B(y[106]), .Z(n814) );
  XOR U799 ( .A(x[110]), .B(y[110]), .Z(n811) );
  XOR U800 ( .A(x[195]), .B(y[195]), .Z(n812) );
  XOR U801 ( .A(n811), .B(n812), .Z(n813) );
  XNOR U802 ( .A(n814), .B(n813), .Z(n1419) );
  XOR U803 ( .A(x[102]), .B(y[102]), .Z(n820) );
  XOR U804 ( .A(x[104]), .B(y[104]), .Z(n817) );
  XOR U805 ( .A(x[453]), .B(y[453]), .Z(n818) );
  XOR U806 ( .A(n817), .B(n818), .Z(n819) );
  XNOR U807 ( .A(n820), .B(n819), .Z(n1418) );
  XOR U808 ( .A(n1419), .B(n1418), .Z(n1420) );
  XOR U809 ( .A(n1421), .B(n1420), .Z(n58) );
  XNOR U810 ( .A(n59), .B(n58), .Z(n1172) );
  XOR U811 ( .A(x[98]), .B(y[98]), .Z(n1415) );
  XOR U812 ( .A(x[100]), .B(y[100]), .Z(n1412) );
  XOR U813 ( .A(x[199]), .B(y[199]), .Z(n1413) );
  XOR U814 ( .A(n1412), .B(n1413), .Z(n1414) );
  XNOR U815 ( .A(n1415), .B(n1414), .Z(n1373) );
  XOR U816 ( .A(x[92]), .B(y[92]), .Z(n1403) );
  XOR U817 ( .A(x[96]), .B(y[96]), .Z(n1400) );
  XOR U818 ( .A(x[451]), .B(y[451]), .Z(n1401) );
  XOR U819 ( .A(n1400), .B(n1401), .Z(n1402) );
  XNOR U820 ( .A(n1403), .B(n1402), .Z(n1371) );
  XOR U821 ( .A(x[88]), .B(y[88]), .Z(n1409) );
  XOR U822 ( .A(x[90]), .B(y[90]), .Z(n1406) );
  XOR U823 ( .A(x[203]), .B(y[203]), .Z(n1407) );
  XOR U824 ( .A(n1406), .B(n1407), .Z(n1408) );
  XNOR U825 ( .A(n1409), .B(n1408), .Z(n1370) );
  XOR U826 ( .A(n1371), .B(n1370), .Z(n1372) );
  XOR U827 ( .A(n1373), .B(n1372), .Z(n337) );
  XOR U828 ( .A(x[84]), .B(y[84]), .Z(n964) );
  XOR U829 ( .A(x[86]), .B(y[86]), .Z(n961) );
  XOR U830 ( .A(x[449]), .B(y[449]), .Z(n962) );
  XOR U831 ( .A(n961), .B(n962), .Z(n963) );
  XNOR U832 ( .A(n964), .B(n963), .Z(n1548) );
  XOR U833 ( .A(x[80]), .B(y[80]), .Z(n952) );
  XOR U834 ( .A(x[82]), .B(y[82]), .Z(n949) );
  XOR U835 ( .A(x[207]), .B(y[207]), .Z(n950) );
  XOR U836 ( .A(n949), .B(n950), .Z(n951) );
  XNOR U837 ( .A(n952), .B(n951), .Z(n1546) );
  XOR U838 ( .A(x[76]), .B(y[76]), .Z(n958) );
  XOR U839 ( .A(x[78]), .B(y[78]), .Z(n955) );
  XOR U840 ( .A(x[447]), .B(y[447]), .Z(n956) );
  XOR U841 ( .A(n955), .B(n956), .Z(n957) );
  XNOR U842 ( .A(n958), .B(n957), .Z(n1545) );
  XOR U843 ( .A(n1546), .B(n1545), .Z(n1547) );
  XOR U844 ( .A(n1548), .B(n1547), .Z(n336) );
  XOR U845 ( .A(n337), .B(n336), .Z(n339) );
  XOR U846 ( .A(x[72]), .B(y[72]), .Z(n982) );
  XOR U847 ( .A(x[74]), .B(y[74]), .Z(n979) );
  XOR U848 ( .A(x[211]), .B(y[211]), .Z(n980) );
  XOR U849 ( .A(n979), .B(n980), .Z(n981) );
  XNOR U850 ( .A(n982), .B(n981), .Z(n1506) );
  XOR U851 ( .A(x[68]), .B(y[68]), .Z(n970) );
  XOR U852 ( .A(x[70]), .B(y[70]), .Z(n967) );
  XOR U853 ( .A(x[445]), .B(y[445]), .Z(n968) );
  XOR U854 ( .A(n967), .B(n968), .Z(n969) );
  XNOR U855 ( .A(n970), .B(n969), .Z(n1504) );
  XOR U856 ( .A(x[64]), .B(y[64]), .Z(n976) );
  XOR U857 ( .A(x[66]), .B(y[66]), .Z(n973) );
  XOR U858 ( .A(x[215]), .B(y[215]), .Z(n974) );
  XOR U859 ( .A(n973), .B(n974), .Z(n975) );
  XNOR U860 ( .A(n976), .B(n975), .Z(n1503) );
  XOR U861 ( .A(n1504), .B(n1503), .Z(n1505) );
  XOR U862 ( .A(n1506), .B(n1505), .Z(n338) );
  XNOR U863 ( .A(n339), .B(n338), .Z(n1171) );
  XOR U864 ( .A(n1172), .B(n1171), .Z(n1173) );
  XNOR U865 ( .A(n1174), .B(n1173), .Z(n1553) );
  XOR U866 ( .A(x[440]), .B(y[440]), .Z(n477) );
  XOR U867 ( .A(x[442]), .B(y[442]), .Z(n474) );
  XNOR U868 ( .A(x[444]), .B(y[444]), .Z(n475) );
  XOR U869 ( .A(n477), .B(n476), .Z(n986) );
  XOR U870 ( .A(x[446]), .B(y[446]), .Z(n387) );
  XOR U871 ( .A(x[198]), .B(y[198]), .Z(n384) );
  XNOR U872 ( .A(x[448]), .B(y[448]), .Z(n385) );
  XOR U873 ( .A(n387), .B(n386), .Z(n985) );
  XOR U874 ( .A(n986), .B(n985), .Z(n988) );
  XOR U875 ( .A(x[410]), .B(y[410]), .Z(n513) );
  XOR U876 ( .A(x[166]), .B(y[166]), .Z(n510) );
  XNOR U877 ( .A(x[412]), .B(y[412]), .Z(n511) );
  XOR U878 ( .A(n513), .B(n512), .Z(n987) );
  XNOR U879 ( .A(n988), .B(n987), .Z(n501) );
  XOR U880 ( .A(x[426]), .B(y[426]), .Z(n132) );
  XOR U881 ( .A(x[180]), .B(y[180]), .Z(n129) );
  XNOR U882 ( .A(x[428]), .B(y[428]), .Z(n130) );
  XNOR U883 ( .A(n132), .B(n131), .Z(n499) );
  XOR U884 ( .A(x[420]), .B(y[420]), .Z(n217) );
  XOR U885 ( .A(x[422]), .B(y[422]), .Z(n214) );
  XNOR U886 ( .A(x[424]), .B(y[424]), .Z(n215) );
  XNOR U887 ( .A(n217), .B(n216), .Z(n498) );
  XOR U888 ( .A(n499), .B(n498), .Z(n500) );
  XNOR U889 ( .A(n501), .B(n500), .Z(n1185) );
  XOR U890 ( .A(x[374]), .B(y[374]), .Z(n162) );
  XOR U891 ( .A(x[376]), .B(y[376]), .Z(n159) );
  XOR U892 ( .A(x[378]), .B(y[378]), .Z(n160) );
  XOR U893 ( .A(n159), .B(n160), .Z(n161) );
  XNOR U894 ( .A(n162), .B(n161), .Z(n1379) );
  XOR U895 ( .A(x[466]), .B(y[466]), .Z(n241) );
  XOR U896 ( .A(x[216]), .B(y[216]), .Z(n238) );
  XOR U897 ( .A(x[468]), .B(y[468]), .Z(n239) );
  XOR U898 ( .A(n238), .B(n239), .Z(n240) );
  XNOR U899 ( .A(n241), .B(n240), .Z(n1377) );
  XOR U900 ( .A(x[370]), .B(y[370]), .Z(n156) );
  XOR U901 ( .A(x[130]), .B(y[130]), .Z(n153) );
  XOR U902 ( .A(x[372]), .B(y[372]), .Z(n154) );
  XOR U903 ( .A(n153), .B(n154), .Z(n155) );
  XNOR U904 ( .A(n156), .B(n155), .Z(n1376) );
  XOR U905 ( .A(n1377), .B(n1376), .Z(n1378) );
  XNOR U906 ( .A(n1379), .B(n1378), .Z(n1184) );
  XOR U907 ( .A(x[394]), .B(y[394]), .Z(n211) );
  XOR U908 ( .A(x[396]), .B(y[396]), .Z(n208) );
  XOR U909 ( .A(x[398]), .B(y[398]), .Z(n209) );
  XOR U910 ( .A(n208), .B(n209), .Z(n210) );
  XOR U911 ( .A(n211), .B(n210), .Z(n1397) );
  XOR U912 ( .A(x[454]), .B(y[454]), .Z(n314) );
  XOR U913 ( .A(x[456]), .B(y[456]), .Z(n311) );
  XOR U914 ( .A(x[458]), .B(y[458]), .Z(n312) );
  XOR U915 ( .A(n311), .B(n312), .Z(n313) );
  XNOR U916 ( .A(n314), .B(n313), .Z(n1395) );
  XOR U917 ( .A(x[390]), .B(y[390]), .Z(n71) );
  XOR U918 ( .A(x[148]), .B(y[148]), .Z(n68) );
  XOR U919 ( .A(x[392]), .B(y[392]), .Z(n69) );
  XOR U920 ( .A(n68), .B(n69), .Z(n70) );
  XNOR U921 ( .A(n71), .B(n70), .Z(n1394) );
  XOR U922 ( .A(n1395), .B(n1394), .Z(n1396) );
  XOR U923 ( .A(n1397), .B(n1396), .Z(n1183) );
  XOR U924 ( .A(n1184), .B(n1183), .Z(n1186) );
  XNOR U925 ( .A(n1185), .B(n1186), .Z(n1551) );
  XOR U926 ( .A(x[310]), .B(y[310]), .Z(n192) );
  XOR U927 ( .A(x[111]), .B(y[111]), .Z(n189) );
  XOR U928 ( .A(x[312]), .B(y[312]), .Z(n190) );
  XOR U929 ( .A(n189), .B(n190), .Z(n191) );
  XNOR U930 ( .A(n192), .B(n191), .Z(n1253) );
  XOR U931 ( .A(x[244]), .B(y[244]), .Z(n1344) );
  XOR U932 ( .A(x[246]), .B(y[246]), .Z(n1341) );
  XOR U933 ( .A(x[498]), .B(y[498]), .Z(n1342) );
  XOR U934 ( .A(n1341), .B(n1342), .Z(n1343) );
  XNOR U935 ( .A(n1344), .B(n1343), .Z(n1251) );
  XOR U936 ( .A(x[306]), .B(y[306]), .Z(n186) );
  XOR U937 ( .A(x[308]), .B(y[308]), .Z(n183) );
  XOR U938 ( .A(x[495]), .B(y[495]), .Z(n184) );
  XOR U939 ( .A(n183), .B(n184), .Z(n185) );
  XNOR U940 ( .A(n186), .B(n185), .Z(n1250) );
  XOR U941 ( .A(n1251), .B(n1250), .Z(n1252) );
  XOR U942 ( .A(n1253), .B(n1252), .Z(n1300) );
  XOR U943 ( .A(x[302]), .B(y[302]), .Z(n253) );
  XOR U944 ( .A(x[115]), .B(y[115]), .Z(n250) );
  XOR U945 ( .A(x[304]), .B(y[304]), .Z(n251) );
  XOR U946 ( .A(n250), .B(n251), .Z(n252) );
  XNOR U947 ( .A(n253), .B(n252), .Z(n1241) );
  XOR U948 ( .A(x[298]), .B(y[298]), .Z(n247) );
  XOR U949 ( .A(x[300]), .B(y[300]), .Z(n244) );
  XOR U950 ( .A(x[493]), .B(y[493]), .Z(n245) );
  XOR U951 ( .A(n244), .B(n245), .Z(n246) );
  XNOR U952 ( .A(n247), .B(n246), .Z(n1239) );
  XOR U953 ( .A(x[294]), .B(y[294]), .Z(n101) );
  XOR U954 ( .A(x[119]), .B(y[119]), .Z(n98) );
  XNOR U955 ( .A(x[296]), .B(y[296]), .Z(n99) );
  XNOR U956 ( .A(n101), .B(n100), .Z(n1238) );
  XOR U957 ( .A(n1239), .B(n1238), .Z(n1240) );
  XOR U958 ( .A(n1241), .B(n1240), .Z(n1299) );
  XOR U959 ( .A(n1300), .B(n1299), .Z(n1302) );
  XOR U960 ( .A(x[290]), .B(y[290]), .Z(n95) );
  XOR U961 ( .A(x[292]), .B(y[292]), .Z(n92) );
  XNOR U962 ( .A(x[491]), .B(y[491]), .Z(n93) );
  XNOR U963 ( .A(n95), .B(n94), .Z(n1235) );
  XOR U964 ( .A(x[286]), .B(y[286]), .Z(n639) );
  XOR U965 ( .A(x[123]), .B(y[123]), .Z(n636) );
  XNOR U966 ( .A(x[288]), .B(y[288]), .Z(n637) );
  XNOR U967 ( .A(n639), .B(n638), .Z(n1233) );
  XOR U968 ( .A(x[282]), .B(y[282]), .Z(n633) );
  XOR U969 ( .A(x[284]), .B(y[284]), .Z(n630) );
  XNOR U970 ( .A(x[489]), .B(y[489]), .Z(n631) );
  XNOR U971 ( .A(n633), .B(n632), .Z(n1232) );
  XOR U972 ( .A(n1233), .B(n1232), .Z(n1234) );
  XOR U973 ( .A(n1235), .B(n1234), .Z(n1301) );
  XOR U974 ( .A(n1302), .B(n1301), .Z(n1156) );
  XOR U975 ( .A(x[236]), .B(y[236]), .Z(n1078) );
  XOR U976 ( .A(x[240]), .B(y[240]), .Z(n1075) );
  XOR U977 ( .A(x[479]), .B(y[479]), .Z(n1076) );
  XOR U978 ( .A(n1075), .B(n1076), .Z(n1077) );
  XNOR U979 ( .A(n1078), .B(n1077), .Z(n1295) );
  XOR U980 ( .A(x[230]), .B(y[230]), .Z(n1024) );
  XOR U981 ( .A(x[147]), .B(y[147]), .Z(n1021) );
  XOR U982 ( .A(x[232]), .B(y[232]), .Z(n1022) );
  XOR U983 ( .A(n1021), .B(n1022), .Z(n1023) );
  XNOR U984 ( .A(n1024), .B(n1023), .Z(n1293) );
  XOR U985 ( .A(x[226]), .B(y[226]), .Z(n1126) );
  XOR U986 ( .A(x[228]), .B(y[228]), .Z(n1123) );
  XNOR U987 ( .A(x[477]), .B(y[477]), .Z(n1124) );
  XNOR U988 ( .A(n1126), .B(n1125), .Z(n1292) );
  XOR U989 ( .A(n1293), .B(n1292), .Z(n1294) );
  XOR U990 ( .A(n1295), .B(n1294), .Z(n409) );
  XOR U991 ( .A(x[222]), .B(y[222]), .Z(n579) );
  XOR U992 ( .A(x[151]), .B(y[151]), .Z(n576) );
  XOR U993 ( .A(x[224]), .B(y[224]), .Z(n577) );
  XOR U994 ( .A(n576), .B(n577), .Z(n578) );
  XNOR U995 ( .A(n579), .B(n578), .Z(n1223) );
  XOR U996 ( .A(x[214]), .B(y[214]), .Z(n573) );
  XOR U997 ( .A(x[218]), .B(y[218]), .Z(n570) );
  XOR U998 ( .A(x[475]), .B(y[475]), .Z(n571) );
  XOR U999 ( .A(n570), .B(n571), .Z(n572) );
  XNOR U1000 ( .A(n573), .B(n572), .Z(n1221) );
  XOR U1001 ( .A(x[210]), .B(y[210]), .Z(n1132) );
  XOR U1002 ( .A(x[155]), .B(y[155]), .Z(n1129) );
  XNOR U1003 ( .A(x[212]), .B(y[212]), .Z(n1130) );
  XNOR U1004 ( .A(n1132), .B(n1131), .Z(n1220) );
  XOR U1005 ( .A(n1221), .B(n1220), .Z(n1222) );
  XOR U1006 ( .A(n1223), .B(n1222), .Z(n408) );
  XOR U1007 ( .A(n409), .B(n408), .Z(n411) );
  XOR U1008 ( .A(x[206]), .B(y[206]), .Z(n784) );
  XOR U1009 ( .A(x[208]), .B(y[208]), .Z(n781) );
  XOR U1010 ( .A(x[473]), .B(y[473]), .Z(n782) );
  XOR U1011 ( .A(n781), .B(n782), .Z(n783) );
  XNOR U1012 ( .A(n784), .B(n783), .Z(n1229) );
  XOR U1013 ( .A(x[200]), .B(y[200]), .Z(n705) );
  XOR U1014 ( .A(x[159]), .B(y[159]), .Z(n702) );
  XNOR U1015 ( .A(x[204]), .B(y[204]), .Z(n703) );
  XNOR U1016 ( .A(n705), .B(n704), .Z(n1227) );
  XOR U1017 ( .A(x[194]), .B(y[194]), .Z(n1036) );
  XOR U1018 ( .A(x[196]), .B(y[196]), .Z(n1033) );
  XOR U1019 ( .A(x[471]), .B(y[471]), .Z(n1034) );
  XOR U1020 ( .A(n1033), .B(n1034), .Z(n1035) );
  XNOR U1021 ( .A(n1036), .B(n1035), .Z(n1226) );
  XOR U1022 ( .A(n1227), .B(n1226), .Z(n1228) );
  XOR U1023 ( .A(n1229), .B(n1228), .Z(n410) );
  XOR U1024 ( .A(n411), .B(n410), .Z(n1154) );
  XOR U1025 ( .A(x[242]), .B(y[242]), .Z(n1018) );
  XOR U1026 ( .A(x[143]), .B(y[143]), .Z(n1015) );
  XOR U1027 ( .A(x[248]), .B(y[248]), .Z(n1016) );
  XOR U1028 ( .A(n1015), .B(n1016), .Z(n1017) );
  XOR U1029 ( .A(n1018), .B(n1017), .Z(n1215) );
  XOR U1030 ( .A(x[250]), .B(y[250]), .Z(n892) );
  XOR U1031 ( .A(x[252]), .B(y[252]), .Z(n889) );
  XOR U1032 ( .A(x[481]), .B(y[481]), .Z(n890) );
  XOR U1033 ( .A(n889), .B(n890), .Z(n891) );
  XOR U1034 ( .A(n892), .B(n891), .Z(n1214) );
  XOR U1035 ( .A(n1215), .B(n1214), .Z(n1217) );
  XOR U1036 ( .A(x[254]), .B(y[254]), .Z(n898) );
  XOR U1037 ( .A(x[139]), .B(y[139]), .Z(n895) );
  XOR U1038 ( .A(x[256]), .B(y[256]), .Z(n896) );
  XOR U1039 ( .A(n895), .B(n896), .Z(n897) );
  XOR U1040 ( .A(n898), .B(n897), .Z(n1216) );
  XNOR U1041 ( .A(n1217), .B(n1216), .Z(n1257) );
  XOR U1042 ( .A(x[278]), .B(y[278]), .Z(n657) );
  XOR U1043 ( .A(x[127]), .B(y[127]), .Z(n654) );
  XNOR U1044 ( .A(x[280]), .B(y[280]), .Z(n655) );
  XNOR U1045 ( .A(n657), .B(n656), .Z(n1283) );
  XOR U1046 ( .A(x[274]), .B(y[274]), .Z(n651) );
  XOR U1047 ( .A(x[276]), .B(y[276]), .Z(n648) );
  XNOR U1048 ( .A(x[487]), .B(y[487]), .Z(n649) );
  XNOR U1049 ( .A(n651), .B(n650), .Z(n1281) );
  XOR U1050 ( .A(x[270]), .B(y[270]), .Z(n621) );
  XOR U1051 ( .A(x[131]), .B(y[131]), .Z(n618) );
  XNOR U1052 ( .A(x[272]), .B(y[272]), .Z(n619) );
  XNOR U1053 ( .A(n621), .B(n620), .Z(n1280) );
  XOR U1054 ( .A(n1281), .B(n1280), .Z(n1282) );
  XOR U1055 ( .A(n1283), .B(n1282), .Z(n1256) );
  XOR U1056 ( .A(n1257), .B(n1256), .Z(n1259) );
  XOR U1057 ( .A(x[266]), .B(y[266]), .Z(n615) );
  XOR U1058 ( .A(x[268]), .B(y[268]), .Z(n612) );
  XNOR U1059 ( .A(x[485]), .B(y[485]), .Z(n613) );
  XNOR U1060 ( .A(n615), .B(n614), .Z(n1289) );
  XOR U1061 ( .A(x[262]), .B(y[262]), .Z(n723) );
  XOR U1062 ( .A(x[135]), .B(y[135]), .Z(n720) );
  XNOR U1063 ( .A(x[264]), .B(y[264]), .Z(n721) );
  XNOR U1064 ( .A(n723), .B(n722), .Z(n1287) );
  XOR U1065 ( .A(x[258]), .B(y[258]), .Z(n717) );
  XOR U1066 ( .A(x[260]), .B(y[260]), .Z(n714) );
  XNOR U1067 ( .A(x[483]), .B(y[483]), .Z(n715) );
  XNOR U1068 ( .A(n717), .B(n716), .Z(n1286) );
  XOR U1069 ( .A(n1287), .B(n1286), .Z(n1288) );
  XOR U1070 ( .A(n1289), .B(n1288), .Z(n1258) );
  XOR U1071 ( .A(n1259), .B(n1258), .Z(n1153) );
  XOR U1072 ( .A(n1154), .B(n1153), .Z(n1155) );
  XOR U1073 ( .A(n1156), .B(n1155), .Z(n1552) );
  XOR U1074 ( .A(n1551), .B(n1552), .Z(n1554) );
  XOR U1075 ( .A(n1553), .B(n1554), .Z(n531) );
  XOR U1076 ( .A(x[85]), .B(y[85]), .Z(n886) );
  XOR U1077 ( .A(x[81]), .B(y[81]), .Z(n883) );
  XOR U1078 ( .A(x[83]), .B(y[83]), .Z(n884) );
  XOR U1079 ( .A(n883), .B(n884), .Z(n885) );
  XNOR U1080 ( .A(n886), .B(n885), .Z(n332) );
  XOR U1081 ( .A(x[91]), .B(y[91]), .Z(n1012) );
  XOR U1082 ( .A(x[87]), .B(y[87]), .Z(n1009) );
  XOR U1083 ( .A(x[89]), .B(y[89]), .Z(n1010) );
  XOR U1084 ( .A(n1009), .B(n1010), .Z(n1011) );
  XNOR U1085 ( .A(n1012), .B(n1011), .Z(n330) );
  XOR U1086 ( .A(x[97]), .B(y[97]), .Z(n856) );
  XOR U1087 ( .A(x[93]), .B(y[93]), .Z(n853) );
  XOR U1088 ( .A(x[95]), .B(y[95]), .Z(n854) );
  XOR U1089 ( .A(n853), .B(n854), .Z(n855) );
  XNOR U1090 ( .A(n856), .B(n855), .Z(n329) );
  XOR U1091 ( .A(n330), .B(n329), .Z(n331) );
  XOR U1092 ( .A(n332), .B(n331), .Z(n541) );
  XOR U1093 ( .A(x[105]), .B(y[105]), .Z(n1066) );
  XOR U1094 ( .A(x[99]), .B(y[99]), .Z(n1063) );
  XOR U1095 ( .A(x[101]), .B(y[101]), .Z(n1064) );
  XOR U1096 ( .A(n1063), .B(n1064), .Z(n1065) );
  XNOR U1097 ( .A(n1066), .B(n1065), .Z(n495) );
  XOR U1098 ( .A(x[117]), .B(y[117]), .Z(n1120) );
  XOR U1099 ( .A(x[109]), .B(y[109]), .Z(n1117) );
  XOR U1100 ( .A(x[113]), .B(y[113]), .Z(n1118) );
  XOR U1101 ( .A(n1117), .B(n1118), .Z(n1119) );
  XNOR U1102 ( .A(n1120), .B(n1119), .Z(n493) );
  XOR U1103 ( .A(x[129]), .B(y[129]), .Z(n567) );
  XOR U1104 ( .A(x[121]), .B(y[121]), .Z(n564) );
  XOR U1105 ( .A(x[125]), .B(y[125]), .Z(n565) );
  XOR U1106 ( .A(n564), .B(n565), .Z(n566) );
  XNOR U1107 ( .A(n567), .B(n566), .Z(n492) );
  XOR U1108 ( .A(n493), .B(n492), .Z(n494) );
  XOR U1109 ( .A(n495), .B(n494), .Z(n540) );
  XOR U1110 ( .A(n541), .B(n540), .Z(n543) );
  XOR U1111 ( .A(x[141]), .B(y[141]), .Z(n1072) );
  XOR U1112 ( .A(x[133]), .B(y[133]), .Z(n1069) );
  XOR U1113 ( .A(x[137]), .B(y[137]), .Z(n1070) );
  XOR U1114 ( .A(n1069), .B(n1070), .Z(n1071) );
  XNOR U1115 ( .A(n1072), .B(n1071), .Z(n205) );
  XOR U1116 ( .A(x[153]), .B(y[153]), .Z(n465) );
  XOR U1117 ( .A(x[145]), .B(y[145]), .Z(n462) );
  XOR U1118 ( .A(x[149]), .B(y[149]), .Z(n463) );
  XOR U1119 ( .A(n462), .B(n463), .Z(n464) );
  XNOR U1120 ( .A(n465), .B(n464), .Z(n203) );
  XOR U1121 ( .A(x[165]), .B(y[165]), .Z(n453) );
  XOR U1122 ( .A(x[157]), .B(y[157]), .Z(n450) );
  XOR U1123 ( .A(x[161]), .B(y[161]), .Z(n451) );
  XOR U1124 ( .A(n450), .B(n451), .Z(n452) );
  XNOR U1125 ( .A(n453), .B(n452), .Z(n202) );
  XOR U1126 ( .A(n203), .B(n202), .Z(n204) );
  XOR U1127 ( .A(n205), .B(n204), .Z(n542) );
  XNOR U1128 ( .A(n543), .B(n542), .Z(n1211) );
  XOR U1129 ( .A(x[177]), .B(y[177]), .Z(n459) );
  XOR U1130 ( .A(x[169]), .B(y[169]), .Z(n456) );
  XOR U1131 ( .A(x[173]), .B(y[173]), .Z(n457) );
  XOR U1132 ( .A(n456), .B(n457), .Z(n458) );
  XNOR U1133 ( .A(n459), .B(n458), .Z(n138) );
  XOR U1134 ( .A(x[189]), .B(y[189]), .Z(n772) );
  XOR U1135 ( .A(x[181]), .B(y[181]), .Z(n769) );
  XOR U1136 ( .A(x[185]), .B(y[185]), .Z(n770) );
  XOR U1137 ( .A(n769), .B(n770), .Z(n771) );
  XNOR U1138 ( .A(n772), .B(n771), .Z(n136) );
  XOR U1139 ( .A(x[201]), .B(y[201]), .Z(n1030) );
  XOR U1140 ( .A(x[193]), .B(y[193]), .Z(n1027) );
  XOR U1141 ( .A(x[197]), .B(y[197]), .Z(n1028) );
  XOR U1142 ( .A(n1027), .B(n1028), .Z(n1029) );
  XNOR U1143 ( .A(n1030), .B(n1029), .Z(n135) );
  XOR U1144 ( .A(n136), .B(n135), .Z(n137) );
  XOR U1145 ( .A(n138), .B(n137), .Z(n535) );
  XOR U1146 ( .A(x[381]), .B(y[381]), .Z(n832) );
  XOR U1147 ( .A(x[379]), .B(y[379]), .Z(n829) );
  XOR U1148 ( .A(x[405]), .B(y[405]), .Z(n830) );
  XOR U1149 ( .A(n829), .B(n830), .Z(n831) );
  XNOR U1150 ( .A(n832), .B(n831), .Z(n808) );
  XOR U1151 ( .A(x[401]), .B(y[401]), .Z(n766) );
  XOR U1152 ( .A(x[397]), .B(y[397]), .Z(n763) );
  XOR U1153 ( .A(x[403]), .B(y[403]), .Z(n764) );
  XOR U1154 ( .A(n763), .B(n764), .Z(n765) );
  XNOR U1155 ( .A(n766), .B(n765), .Z(n806) );
  XOR U1156 ( .A(x[391]), .B(y[391]), .Z(n760) );
  XOR U1157 ( .A(x[385]), .B(y[385]), .Z(n757) );
  XOR U1158 ( .A(x[387]), .B(y[387]), .Z(n758) );
  XOR U1159 ( .A(n757), .B(n758), .Z(n759) );
  XNOR U1160 ( .A(n760), .B(n759), .Z(n805) );
  XOR U1161 ( .A(n806), .B(n805), .Z(n807) );
  XOR U1162 ( .A(n808), .B(n807), .Z(n534) );
  XOR U1163 ( .A(n535), .B(n534), .Z(n537) );
  XOR U1164 ( .A(x[213]), .B(y[213]), .Z(n778) );
  XOR U1165 ( .A(x[205]), .B(y[205]), .Z(n775) );
  XOR U1166 ( .A(x[209]), .B(y[209]), .Z(n776) );
  XOR U1167 ( .A(n775), .B(n776), .Z(n777) );
  XNOR U1168 ( .A(n778), .B(n777), .Z(n168) );
  XOR U1169 ( .A(x[225]), .B(y[225]), .Z(n1096) );
  XOR U1170 ( .A(x[217]), .B(y[217]), .Z(n1093) );
  XOR U1171 ( .A(x[221]), .B(y[221]), .Z(n1094) );
  XOR U1172 ( .A(n1093), .B(n1094), .Z(n1095) );
  XNOR U1173 ( .A(n1096), .B(n1095), .Z(n166) );
  XOR U1174 ( .A(x[235]), .B(y[235]), .Z(n1084) );
  XOR U1175 ( .A(x[229]), .B(y[229]), .Z(n1081) );
  XOR U1176 ( .A(x[233]), .B(y[233]), .Z(n1082) );
  XOR U1177 ( .A(n1081), .B(n1082), .Z(n1083) );
  XNOR U1178 ( .A(n1084), .B(n1083), .Z(n165) );
  XOR U1179 ( .A(n166), .B(n165), .Z(n167) );
  XOR U1180 ( .A(n168), .B(n167), .Z(n536) );
  XNOR U1181 ( .A(n537), .B(n536), .Z(n1209) );
  XOR U1182 ( .A(x[313]), .B(y[313]), .Z(n1108) );
  XOR U1183 ( .A(x[309]), .B(y[309]), .Z(n1105) );
  XOR U1184 ( .A(x[311]), .B(y[311]), .Z(n1106) );
  XOR U1185 ( .A(n1105), .B(n1106), .Z(n1107) );
  XNOR U1186 ( .A(n1108), .B(n1107), .Z(n375) );
  XOR U1187 ( .A(x[317]), .B(y[317]), .Z(n1060) );
  XOR U1188 ( .A(x[315]), .B(y[315]), .Z(n1057) );
  XOR U1189 ( .A(x[433]), .B(y[433]), .Z(n1058) );
  XOR U1190 ( .A(n1057), .B(n1058), .Z(n1059) );
  XNOR U1191 ( .A(n1060), .B(n1059), .Z(n373) );
  XOR U1192 ( .A(x[321]), .B(y[321]), .Z(n1048) );
  XOR U1193 ( .A(x[319]), .B(y[319]), .Z(n1045) );
  XOR U1194 ( .A(x[431]), .B(y[431]), .Z(n1046) );
  XOR U1195 ( .A(n1045), .B(n1046), .Z(n1047) );
  XNOR U1196 ( .A(n1048), .B(n1047), .Z(n372) );
  XOR U1197 ( .A(n373), .B(n372), .Z(n374) );
  XOR U1198 ( .A(n375), .B(n374), .Z(n661) );
  XOR U1199 ( .A(x[349]), .B(y[349]), .Z(n916) );
  XOR U1200 ( .A(x[347]), .B(y[347]), .Z(n913) );
  XNOR U1201 ( .A(x[417]), .B(y[417]), .Z(n914) );
  XNOR U1202 ( .A(n916), .B(n915), .Z(n381) );
  XOR U1203 ( .A(x[353]), .B(y[353]), .Z(n1150) );
  XOR U1204 ( .A(x[351]), .B(y[351]), .Z(n1147) );
  XOR U1205 ( .A(x[415]), .B(y[415]), .Z(n1148) );
  XOR U1206 ( .A(n1147), .B(n1148), .Z(n1149) );
  XNOR U1207 ( .A(n1150), .B(n1149), .Z(n379) );
  XOR U1208 ( .A(x[357]), .B(y[357]), .Z(n1138) );
  XOR U1209 ( .A(x[355]), .B(y[355]), .Z(n1135) );
  XOR U1210 ( .A(x[413]), .B(y[413]), .Z(n1136) );
  XOR U1211 ( .A(n1135), .B(n1136), .Z(n1137) );
  XNOR U1212 ( .A(n1138), .B(n1137), .Z(n378) );
  XOR U1213 ( .A(n379), .B(n378), .Z(n380) );
  XOR U1214 ( .A(n381), .B(n380), .Z(n660) );
  XOR U1215 ( .A(n661), .B(n660), .Z(n663) );
  XOR U1216 ( .A(x[325]), .B(y[325]), .Z(n1054) );
  XOR U1217 ( .A(x[323]), .B(y[323]), .Z(n1051) );
  XOR U1218 ( .A(x[429]), .B(y[429]), .Z(n1052) );
  XOR U1219 ( .A(n1051), .B(n1052), .Z(n1053) );
  XNOR U1220 ( .A(n1054), .B(n1053), .Z(n114) );
  XOR U1221 ( .A(x[329]), .B(y[329]), .Z(n1006) );
  XOR U1222 ( .A(x[327]), .B(y[327]), .Z(n1003) );
  XOR U1223 ( .A(x[427]), .B(y[427]), .Z(n1004) );
  XOR U1224 ( .A(n1003), .B(n1004), .Z(n1005) );
  XNOR U1225 ( .A(n1006), .B(n1005), .Z(n112) );
  XOR U1226 ( .A(x[333]), .B(y[333]), .Z(n994) );
  XOR U1227 ( .A(x[331]), .B(y[331]), .Z(n991) );
  XOR U1228 ( .A(x[425]), .B(y[425]), .Z(n992) );
  XOR U1229 ( .A(n991), .B(n992), .Z(n993) );
  XNOR U1230 ( .A(n994), .B(n993), .Z(n111) );
  XOR U1231 ( .A(n112), .B(n111), .Z(n113) );
  XOR U1232 ( .A(n114), .B(n113), .Z(n662) );
  XNOR U1233 ( .A(n663), .B(n662), .Z(n1208) );
  XOR U1234 ( .A(n1209), .B(n1208), .Z(n1210) );
  XOR U1235 ( .A(n1211), .B(n1210), .Z(n53) );
  XOR U1236 ( .A(x[60]), .B(y[60]), .Z(n880) );
  XOR U1237 ( .A(x[62]), .B(y[62]), .Z(n877) );
  XOR U1238 ( .A(x[443]), .B(y[443]), .Z(n878) );
  XOR U1239 ( .A(n877), .B(n878), .Z(n879) );
  XNOR U1240 ( .A(n880), .B(n879), .Z(n1464) );
  XOR U1241 ( .A(x[56]), .B(y[56]), .Z(n868) );
  XOR U1242 ( .A(x[58]), .B(y[58]), .Z(n865) );
  XOR U1243 ( .A(x[219]), .B(y[219]), .Z(n866) );
  XOR U1244 ( .A(n865), .B(n866), .Z(n867) );
  XNOR U1245 ( .A(n868), .B(n867), .Z(n1462) );
  XOR U1246 ( .A(x[52]), .B(y[52]), .Z(n874) );
  XOR U1247 ( .A(x[54]), .B(y[54]), .Z(n871) );
  XOR U1248 ( .A(x[441]), .B(y[441]), .Z(n872) );
  XOR U1249 ( .A(n871), .B(n872), .Z(n873) );
  XNOR U1250 ( .A(n874), .B(n873), .Z(n1461) );
  XOR U1251 ( .A(n1462), .B(n1461), .Z(n1463) );
  XOR U1252 ( .A(n1464), .B(n1463), .Z(n343) );
  XOR U1253 ( .A(x[48]), .B(y[48]), .Z(n1482) );
  XOR U1254 ( .A(x[50]), .B(y[50]), .Z(n1479) );
  XOR U1255 ( .A(x[223]), .B(y[223]), .Z(n1480) );
  XOR U1256 ( .A(n1479), .B(n1480), .Z(n1481) );
  XNOR U1257 ( .A(n1482), .B(n1481), .Z(n107) );
  XOR U1258 ( .A(x[44]), .B(y[44]), .Z(n1470) );
  XOR U1259 ( .A(x[46]), .B(y[46]), .Z(n1467) );
  XOR U1260 ( .A(x[439]), .B(y[439]), .Z(n1468) );
  XOR U1261 ( .A(n1467), .B(n1468), .Z(n1469) );
  XNOR U1262 ( .A(n1470), .B(n1469), .Z(n105) );
  XOR U1263 ( .A(x[40]), .B(y[40]), .Z(n1476) );
  XOR U1264 ( .A(x[42]), .B(y[42]), .Z(n1473) );
  XOR U1265 ( .A(x[227]), .B(y[227]), .Z(n1474) );
  XOR U1266 ( .A(n1473), .B(n1474), .Z(n1475) );
  XNOR U1267 ( .A(n1476), .B(n1475), .Z(n104) );
  XOR U1268 ( .A(n105), .B(n104), .Z(n106) );
  XOR U1269 ( .A(n107), .B(n106), .Z(n342) );
  XOR U1270 ( .A(n343), .B(n342), .Z(n345) );
  XOR U1271 ( .A(x[36]), .B(y[36]), .Z(n1542) );
  XOR U1272 ( .A(x[38]), .B(y[38]), .Z(n1539) );
  XNOR U1273 ( .A(x[437]), .B(y[437]), .Z(n1540) );
  XNOR U1274 ( .A(n1542), .B(n1541), .Z(n174) );
  XOR U1275 ( .A(x[32]), .B(y[32]), .Z(n1530) );
  XOR U1276 ( .A(x[34]), .B(y[34]), .Z(n1527) );
  XNOR U1277 ( .A(x[231]), .B(y[231]), .Z(n1528) );
  XNOR U1278 ( .A(n1530), .B(n1529), .Z(n172) );
  XOR U1279 ( .A(x[28]), .B(y[28]), .Z(n1536) );
  XOR U1280 ( .A(x[30]), .B(y[30]), .Z(n1533) );
  XNOR U1281 ( .A(x[435]), .B(y[435]), .Z(n1534) );
  XNOR U1282 ( .A(n1536), .B(n1535), .Z(n171) );
  XOR U1283 ( .A(n172), .B(n171), .Z(n173) );
  XOR U1284 ( .A(n174), .B(n173), .Z(n344) );
  XOR U1285 ( .A(n345), .B(n344), .Z(n1332) );
  XOR U1286 ( .A(x[31]), .B(y[31]), .Z(n1452) );
  XOR U1287 ( .A(x[27]), .B(y[27]), .Z(n1449) );
  XNOR U1288 ( .A(x[29]), .B(y[29]), .Z(n1450) );
  XNOR U1289 ( .A(n1452), .B(n1451), .Z(n296) );
  XOR U1290 ( .A(x[37]), .B(y[37]), .Z(n597) );
  XOR U1291 ( .A(x[33]), .B(y[33]), .Z(n594) );
  XNOR U1292 ( .A(x[35]), .B(y[35]), .Z(n595) );
  XNOR U1293 ( .A(n597), .B(n596), .Z(n294) );
  XOR U1294 ( .A(x[43]), .B(y[43]), .Z(n585) );
  XOR U1295 ( .A(x[39]), .B(y[39]), .Z(n582) );
  XNOR U1296 ( .A(x[41]), .B(y[41]), .Z(n583) );
  XNOR U1297 ( .A(n585), .B(n584), .Z(n293) );
  XOR U1298 ( .A(n294), .B(n293), .Z(n295) );
  XOR U1299 ( .A(n296), .B(n295), .Z(n667) );
  XOR U1300 ( .A(x[49]), .B(y[49]), .Z(n591) );
  XOR U1301 ( .A(x[45]), .B(y[45]), .Z(n588) );
  XOR U1302 ( .A(x[47]), .B(y[47]), .Z(n589) );
  XOR U1303 ( .A(n588), .B(n589), .Z(n590) );
  XNOR U1304 ( .A(n591), .B(n590), .Z(n235) );
  XOR U1305 ( .A(x[55]), .B(y[55]), .Z(n748) );
  XOR U1306 ( .A(x[51]), .B(y[51]), .Z(n745) );
  XOR U1307 ( .A(x[53]), .B(y[53]), .Z(n746) );
  XOR U1308 ( .A(n745), .B(n746), .Z(n747) );
  XNOR U1309 ( .A(n748), .B(n747), .Z(n233) );
  XOR U1310 ( .A(x[61]), .B(y[61]), .Z(n736) );
  XOR U1311 ( .A(x[57]), .B(y[57]), .Z(n733) );
  XOR U1312 ( .A(x[59]), .B(y[59]), .Z(n734) );
  XOR U1313 ( .A(n733), .B(n734), .Z(n735) );
  XNOR U1314 ( .A(n736), .B(n735), .Z(n232) );
  XOR U1315 ( .A(n233), .B(n232), .Z(n234) );
  XOR U1316 ( .A(n235), .B(n234), .Z(n666) );
  XOR U1317 ( .A(n667), .B(n666), .Z(n669) );
  XOR U1318 ( .A(x[67]), .B(y[67]), .Z(n742) );
  XOR U1319 ( .A(x[63]), .B(y[63]), .Z(n739) );
  XOR U1320 ( .A(x[65]), .B(y[65]), .Z(n740) );
  XOR U1321 ( .A(n739), .B(n740), .Z(n741) );
  XNOR U1322 ( .A(n742), .B(n741), .Z(n405) );
  XOR U1323 ( .A(x[73]), .B(y[73]), .Z(n862) );
  XOR U1324 ( .A(x[69]), .B(y[69]), .Z(n859) );
  XOR U1325 ( .A(x[71]), .B(y[71]), .Z(n860) );
  XOR U1326 ( .A(n859), .B(n860), .Z(n861) );
  XNOR U1327 ( .A(n862), .B(n861), .Z(n403) );
  XOR U1328 ( .A(x[79]), .B(y[79]), .Z(n850) );
  XOR U1329 ( .A(x[75]), .B(y[75]), .Z(n847) );
  XOR U1330 ( .A(x[77]), .B(y[77]), .Z(n848) );
  XOR U1331 ( .A(n847), .B(n848), .Z(n849) );
  XNOR U1332 ( .A(n850), .B(n849), .Z(n402) );
  XOR U1333 ( .A(n403), .B(n402), .Z(n404) );
  XOR U1334 ( .A(n405), .B(n404), .Z(n668) );
  XOR U1335 ( .A(n669), .B(n668), .Z(n1330) );
  XOR U1336 ( .A(x[22]), .B(y[22]), .Z(n1524) );
  XOR U1337 ( .A(x[24]), .B(y[24]), .Z(n1521) );
  XNOR U1338 ( .A(x[26]), .B(y[26]), .Z(n1522) );
  XNOR U1339 ( .A(n1524), .B(n1523), .Z(n198) );
  XOR U1340 ( .A(x[16]), .B(y[16]), .Z(n1512) );
  XOR U1341 ( .A(x[18]), .B(y[18]), .Z(n1509) );
  XNOR U1342 ( .A(x[20]), .B(y[20]), .Z(n1510) );
  XNOR U1343 ( .A(n1512), .B(n1511), .Z(n196) );
  XOR U1344 ( .A(x[10]), .B(y[10]), .Z(n1518) );
  XOR U1345 ( .A(x[12]), .B(y[12]), .Z(n1515) );
  XNOR U1346 ( .A(x[14]), .B(y[14]), .Z(n1516) );
  XNOR U1347 ( .A(n1518), .B(n1517), .Z(n195) );
  XOR U1348 ( .A(n196), .B(n195), .Z(n197) );
  XOR U1349 ( .A(n198), .B(n197), .Z(n601) );
  XOR U1350 ( .A(x[4]), .B(y[4]), .Z(n1367) );
  XOR U1351 ( .A(x[6]), .B(y[6]), .Z(n1364) );
  XOR U1352 ( .A(x[8]), .B(y[8]), .Z(n1365) );
  XOR U1353 ( .A(n1364), .B(n1365), .Z(n1366) );
  XNOR U1354 ( .A(n1367), .B(n1366), .Z(n308) );
  XOR U1355 ( .A(x[1]), .B(y[1]), .Z(n1361) );
  XOR U1356 ( .A(x[0]), .B(y[0]), .Z(n1358) );
  XOR U1357 ( .A(x[2]), .B(y[2]), .Z(n1359) );
  XOR U1358 ( .A(n1358), .B(n1359), .Z(n1360) );
  XNOR U1359 ( .A(n1361), .B(n1360), .Z(n306) );
  XOR U1360 ( .A(x[7]), .B(y[7]), .Z(n1355) );
  XOR U1361 ( .A(x[3]), .B(y[3]), .Z(n1352) );
  XOR U1362 ( .A(x[5]), .B(y[5]), .Z(n1353) );
  XOR U1363 ( .A(n1352), .B(n1353), .Z(n1354) );
  XNOR U1364 ( .A(n1355), .B(n1354), .Z(n305) );
  XOR U1365 ( .A(n306), .B(n305), .Z(n307) );
  XOR U1366 ( .A(n308), .B(n307), .Z(n600) );
  XOR U1367 ( .A(n601), .B(n600), .Z(n603) );
  XOR U1368 ( .A(x[13]), .B(y[13]), .Z(n1338) );
  XOR U1369 ( .A(x[9]), .B(y[9]), .Z(n1335) );
  XOR U1370 ( .A(x[11]), .B(y[11]), .Z(n1336) );
  XOR U1371 ( .A(n1335), .B(n1336), .Z(n1337) );
  XNOR U1372 ( .A(n1338), .B(n1337), .Z(n272) );
  XOR U1373 ( .A(x[19]), .B(y[19]), .Z(n1458) );
  XOR U1374 ( .A(x[15]), .B(y[15]), .Z(n1455) );
  XNOR U1375 ( .A(x[17]), .B(y[17]), .Z(n1456) );
  XNOR U1376 ( .A(n1458), .B(n1457), .Z(n270) );
  XOR U1377 ( .A(x[25]), .B(y[25]), .Z(n1446) );
  XOR U1378 ( .A(x[21]), .B(y[21]), .Z(n1443) );
  XNOR U1379 ( .A(x[23]), .B(y[23]), .Z(n1444) );
  XNOR U1380 ( .A(n1446), .B(n1445), .Z(n269) );
  XOR U1381 ( .A(n270), .B(n269), .Z(n271) );
  XOR U1382 ( .A(n272), .B(n271), .Z(n602) );
  XOR U1383 ( .A(n603), .B(n602), .Z(n1329) );
  XOR U1384 ( .A(n1330), .B(n1329), .Z(n1331) );
  XNOR U1385 ( .A(n1332), .B(n1331), .Z(n51) );
  XOR U1386 ( .A(x[366]), .B(y[366]), .Z(n357) );
  XOR U1387 ( .A(x[126]), .B(y[126]), .Z(n354) );
  XOR U1388 ( .A(x[368]), .B(y[368]), .Z(n355) );
  XOR U1389 ( .A(n354), .B(n355), .Z(n356) );
  XNOR U1390 ( .A(n357), .B(n356), .Z(n1277) );
  XOR U1391 ( .A(x[470]), .B(y[470]), .Z(n89) );
  XOR U1392 ( .A(x[220]), .B(y[220]), .Z(n86) );
  XOR U1393 ( .A(x[472]), .B(y[472]), .Z(n87) );
  XOR U1394 ( .A(n86), .B(n87), .Z(n88) );
  XNOR U1395 ( .A(n89), .B(n88), .Z(n1275) );
  XOR U1396 ( .A(x[360]), .B(y[360]), .Z(n120) );
  XOR U1397 ( .A(x[362]), .B(y[362]), .Z(n117) );
  XOR U1398 ( .A(x[364]), .B(y[364]), .Z(n118) );
  XOR U1399 ( .A(n117), .B(n118), .Z(n119) );
  XNOR U1400 ( .A(n120), .B(n119), .Z(n1274) );
  XOR U1401 ( .A(n1275), .B(n1274), .Z(n1276) );
  XOR U1402 ( .A(n1277), .B(n1276), .Z(n1178) );
  XOR U1403 ( .A(x[354]), .B(y[354]), .Z(n223) );
  XOR U1404 ( .A(x[356]), .B(y[356]), .Z(n220) );
  XOR U1405 ( .A(x[358]), .B(y[358]), .Z(n221) );
  XOR U1406 ( .A(n220), .B(n221), .Z(n222) );
  XNOR U1407 ( .A(n223), .B(n222), .Z(n1265) );
  XOR U1408 ( .A(x[474]), .B(y[474]), .Z(n627) );
  XOR U1409 ( .A(x[476]), .B(y[476]), .Z(n624) );
  XOR U1410 ( .A(x[478]), .B(y[478]), .Z(n625) );
  XOR U1411 ( .A(n624), .B(n625), .Z(n626) );
  XNOR U1412 ( .A(n627), .B(n626), .Z(n1263) );
  XOR U1413 ( .A(x[350]), .B(y[350]), .Z(n369) );
  XOR U1414 ( .A(x[112]), .B(y[112]), .Z(n366) );
  XOR U1415 ( .A(x[352]), .B(y[352]), .Z(n367) );
  XOR U1416 ( .A(n366), .B(n367), .Z(n368) );
  XNOR U1417 ( .A(n369), .B(n368), .Z(n1262) );
  XOR U1418 ( .A(n1263), .B(n1262), .Z(n1264) );
  XOR U1419 ( .A(n1265), .B(n1264), .Z(n1177) );
  XOR U1420 ( .A(n1178), .B(n1177), .Z(n1180) );
  XOR U1421 ( .A(x[346]), .B(y[346]), .Z(n489) );
  XOR U1422 ( .A(x[108]), .B(y[108]), .Z(n486) );
  XOR U1423 ( .A(x[348]), .B(y[348]), .Z(n487) );
  XOR U1424 ( .A(n486), .B(n487), .Z(n488) );
  XNOR U1425 ( .A(n489), .B(n488), .Z(n1204) );
  XOR U1426 ( .A(x[480]), .B(y[480]), .Z(n645) );
  XOR U1427 ( .A(x[482]), .B(y[482]), .Z(n642) );
  XOR U1428 ( .A(x[484]), .B(y[484]), .Z(n643) );
  XOR U1429 ( .A(n642), .B(n643), .Z(n644) );
  XNOR U1430 ( .A(n645), .B(n644), .Z(n1202) );
  XOR U1431 ( .A(x[340]), .B(y[340]), .Z(n483) );
  XOR U1432 ( .A(x[342]), .B(y[342]), .Z(n480) );
  XOR U1433 ( .A(x[344]), .B(y[344]), .Z(n481) );
  XOR U1434 ( .A(n480), .B(n481), .Z(n482) );
  XNOR U1435 ( .A(n483), .B(n482), .Z(n1201) );
  XOR U1436 ( .A(n1202), .B(n1201), .Z(n1203) );
  XOR U1437 ( .A(n1204), .B(n1203), .Z(n1179) );
  XNOR U1438 ( .A(n1180), .B(n1179), .Z(n1162) );
  XOR U1439 ( .A(x[400]), .B(y[400]), .Z(n77) );
  XOR U1440 ( .A(x[402]), .B(y[402]), .Z(n74) );
  XOR U1441 ( .A(x[404]), .B(y[404]), .Z(n75) );
  XOR U1442 ( .A(n74), .B(n75), .Z(n76) );
  XOR U1443 ( .A(n77), .B(n76), .Z(n926) );
  XOR U1444 ( .A(x[450]), .B(y[450]), .Z(n278) );
  XOR U1445 ( .A(x[202]), .B(y[202]), .Z(n275) );
  XOR U1446 ( .A(x[452]), .B(y[452]), .Z(n276) );
  XOR U1447 ( .A(n275), .B(n276), .Z(n277) );
  XOR U1448 ( .A(n278), .B(n277), .Z(n925) );
  XOR U1449 ( .A(n926), .B(n925), .Z(n928) );
  XOR U1450 ( .A(x[406]), .B(y[406]), .Z(n83) );
  XOR U1451 ( .A(x[162]), .B(y[162]), .Z(n80) );
  XOR U1452 ( .A(x[408]), .B(y[408]), .Z(n81) );
  XOR U1453 ( .A(n80), .B(n81), .Z(n82) );
  XOR U1454 ( .A(n83), .B(n82), .Z(n927) );
  XNOR U1455 ( .A(n928), .B(n927), .Z(n300) );
  XOR U1456 ( .A(x[430]), .B(y[430]), .Z(n126) );
  XOR U1457 ( .A(x[184]), .B(y[184]), .Z(n123) );
  XNOR U1458 ( .A(x[432]), .B(y[432]), .Z(n124) );
  XNOR U1459 ( .A(n126), .B(n125), .Z(n904) );
  XOR U1460 ( .A(x[434]), .B(y[434]), .Z(n363) );
  XOR U1461 ( .A(x[436]), .B(y[436]), .Z(n360) );
  XNOR U1462 ( .A(x[438]), .B(y[438]), .Z(n361) );
  XNOR U1463 ( .A(n363), .B(n362), .Z(n902) );
  XOR U1464 ( .A(x[414]), .B(y[414]), .Z(n150) );
  XOR U1465 ( .A(x[416]), .B(y[416]), .Z(n147) );
  XNOR U1466 ( .A(x[418]), .B(y[418]), .Z(n148) );
  XNOR U1467 ( .A(n150), .B(n149), .Z(n901) );
  XOR U1468 ( .A(n902), .B(n901), .Z(n903) );
  XOR U1469 ( .A(n904), .B(n903), .Z(n299) );
  XOR U1470 ( .A(n300), .B(n299), .Z(n302) );
  XOR U1471 ( .A(x[386]), .B(y[386]), .Z(n519) );
  XOR U1472 ( .A(x[144]), .B(y[144]), .Z(n516) );
  XOR U1473 ( .A(x[388]), .B(y[388]), .Z(n517) );
  XOR U1474 ( .A(n516), .B(n517), .Z(n518) );
  XNOR U1475 ( .A(n519), .B(n518), .Z(n1391) );
  XOR U1476 ( .A(x[460]), .B(y[460]), .Z(n180) );
  XOR U1477 ( .A(x[462]), .B(y[462]), .Z(n177) );
  XOR U1478 ( .A(x[464]), .B(y[464]), .Z(n178) );
  XOR U1479 ( .A(n177), .B(n178), .Z(n179) );
  XNOR U1480 ( .A(n180), .B(n179), .Z(n1389) );
  XOR U1481 ( .A(x[380]), .B(y[380]), .Z(n507) );
  XOR U1482 ( .A(x[382]), .B(y[382]), .Z(n504) );
  XOR U1483 ( .A(x[384]), .B(y[384]), .Z(n505) );
  XOR U1484 ( .A(n504), .B(n505), .Z(n506) );
  XNOR U1485 ( .A(n507), .B(n506), .Z(n1388) );
  XOR U1486 ( .A(n1389), .B(n1388), .Z(n1390) );
  XOR U1487 ( .A(n1391), .B(n1390), .Z(n301) );
  XNOR U1488 ( .A(n302), .B(n301), .Z(n1160) );
  XOR U1489 ( .A(x[334]), .B(y[334]), .Z(n399) );
  XOR U1490 ( .A(x[336]), .B(y[336]), .Z(n396) );
  XOR U1491 ( .A(x[338]), .B(y[338]), .Z(n397) );
  XOR U1492 ( .A(n396), .B(n397), .Z(n398) );
  XNOR U1493 ( .A(n399), .B(n398), .Z(n1192) );
  XOR U1494 ( .A(x[486]), .B(y[486]), .Z(n609) );
  XOR U1495 ( .A(x[234]), .B(y[234]), .Z(n606) );
  XOR U1496 ( .A(x[488]), .B(y[488]), .Z(n607) );
  XOR U1497 ( .A(n606), .B(n607), .Z(n608) );
  XNOR U1498 ( .A(n609), .B(n608), .Z(n1190) );
  XOR U1499 ( .A(x[330]), .B(y[330]), .Z(n393) );
  XOR U1500 ( .A(x[94]), .B(y[94]), .Z(n390) );
  XOR U1501 ( .A(x[332]), .B(y[332]), .Z(n391) );
  XOR U1502 ( .A(n390), .B(n391), .Z(n392) );
  XNOR U1503 ( .A(n393), .B(n392), .Z(n1189) );
  XOR U1504 ( .A(n1190), .B(n1189), .Z(n1191) );
  XOR U1505 ( .A(n1192), .B(n1191), .Z(n1324) );
  XOR U1506 ( .A(x[326]), .B(y[326]), .Z(n290) );
  XOR U1507 ( .A(x[103]), .B(y[103]), .Z(n287) );
  XOR U1508 ( .A(x[328]), .B(y[328]), .Z(n288) );
  XOR U1509 ( .A(n287), .B(n288), .Z(n289) );
  XNOR U1510 ( .A(n290), .B(n289), .Z(n1320) );
  XOR U1511 ( .A(x[490]), .B(y[490]), .Z(n711) );
  XOR U1512 ( .A(x[238]), .B(y[238]), .Z(n708) );
  XOR U1513 ( .A(x[492]), .B(y[492]), .Z(n709) );
  XOR U1514 ( .A(n708), .B(n709), .Z(n710) );
  XNOR U1515 ( .A(n711), .B(n710), .Z(n1318) );
  XOR U1516 ( .A(x[322]), .B(y[322]), .Z(n284) );
  XOR U1517 ( .A(x[324]), .B(y[324]), .Z(n281) );
  XOR U1518 ( .A(x[499]), .B(y[499]), .Z(n282) );
  XOR U1519 ( .A(n281), .B(n282), .Z(n283) );
  XNOR U1520 ( .A(n284), .B(n283), .Z(n1317) );
  XOR U1521 ( .A(n1318), .B(n1317), .Z(n1319) );
  XOR U1522 ( .A(n1320), .B(n1319), .Z(n1323) );
  XOR U1523 ( .A(n1324), .B(n1323), .Z(n1326) );
  XOR U1524 ( .A(x[318]), .B(y[318]), .Z(n326) );
  XOR U1525 ( .A(x[107]), .B(y[107]), .Z(n323) );
  XOR U1526 ( .A(x[320]), .B(y[320]), .Z(n324) );
  XOR U1527 ( .A(n323), .B(n324), .Z(n325) );
  XNOR U1528 ( .A(n326), .B(n325), .Z(n1308) );
  XOR U1529 ( .A(x[494]), .B(y[494]), .Z(n1349) );
  XOR U1530 ( .A(x[496]), .B(y[496]), .Z(n1347) );
  XOR U1531 ( .A(oglobal[0]), .B(n1347), .Z(n1348) );
  XNOR U1532 ( .A(n1349), .B(n1348), .Z(n1306) );
  XOR U1533 ( .A(x[314]), .B(y[314]), .Z(n320) );
  XOR U1534 ( .A(x[316]), .B(y[316]), .Z(n317) );
  XOR U1535 ( .A(x[497]), .B(y[497]), .Z(n318) );
  XOR U1536 ( .A(n317), .B(n318), .Z(n319) );
  XNOR U1537 ( .A(n320), .B(n319), .Z(n1305) );
  XOR U1538 ( .A(n1306), .B(n1305), .Z(n1307) );
  XOR U1539 ( .A(n1308), .B(n1307), .Z(n1325) );
  XNOR U1540 ( .A(n1326), .B(n1325), .Z(n1159) );
  XOR U1541 ( .A(n1160), .B(n1159), .Z(n1161) );
  XOR U1542 ( .A(n1162), .B(n1161), .Z(n50) );
  XOR U1543 ( .A(n51), .B(n50), .Z(n52) );
  XOR U1544 ( .A(n53), .B(n52), .Z(n529) );
  XOR U1545 ( .A(x[241]), .B(y[241]), .Z(n1090) );
  XOR U1546 ( .A(x[237]), .B(y[237]), .Z(n1087) );
  XOR U1547 ( .A(x[239]), .B(y[239]), .Z(n1088) );
  XOR U1548 ( .A(n1087), .B(n1088), .Z(n1089) );
  XNOR U1549 ( .A(n1090), .B(n1089), .Z(n525) );
  XOR U1550 ( .A(x[247]), .B(y[247]), .Z(n429) );
  XOR U1551 ( .A(x[243]), .B(y[243]), .Z(n426) );
  XOR U1552 ( .A(x[245]), .B(y[245]), .Z(n427) );
  XOR U1553 ( .A(n426), .B(n427), .Z(n428) );
  XNOR U1554 ( .A(n429), .B(n428), .Z(n523) );
  XOR U1555 ( .A(x[253]), .B(y[253]), .Z(n417) );
  XOR U1556 ( .A(x[249]), .B(y[249]), .Z(n414) );
  XOR U1557 ( .A(x[251]), .B(y[251]), .Z(n415) );
  XOR U1558 ( .A(n414), .B(n415), .Z(n416) );
  XNOR U1559 ( .A(n417), .B(n416), .Z(n522) );
  XOR U1560 ( .A(n523), .B(n522), .Z(n524) );
  XOR U1561 ( .A(n525), .B(n524), .Z(n727) );
  XOR U1562 ( .A(x[373]), .B(y[373]), .Z(n796) );
  XOR U1563 ( .A(x[371]), .B(y[371]), .Z(n793) );
  XOR U1564 ( .A(x[407]), .B(y[407]), .Z(n794) );
  XOR U1565 ( .A(n793), .B(n794), .Z(n795) );
  XNOR U1566 ( .A(n796), .B(n795), .Z(n754) );
  XOR U1567 ( .A(x[377]), .B(y[377]), .Z(n844) );
  XOR U1568 ( .A(x[375]), .B(y[375]), .Z(n841) );
  XOR U1569 ( .A(x[389]), .B(y[389]), .Z(n842) );
  XOR U1570 ( .A(n841), .B(n842), .Z(n843) );
  XNOR U1571 ( .A(n844), .B(n843), .Z(n752) );
  XOR U1572 ( .A(x[393]), .B(y[393]), .Z(n838) );
  XOR U1573 ( .A(x[395]), .B(y[395]), .Z(n835) );
  XOR U1574 ( .A(x[399]), .B(y[399]), .Z(n836) );
  XOR U1575 ( .A(n835), .B(n836), .Z(n837) );
  XNOR U1576 ( .A(n838), .B(n837), .Z(n751) );
  XOR U1577 ( .A(n752), .B(n751), .Z(n753) );
  XOR U1578 ( .A(n754), .B(n753), .Z(n726) );
  XOR U1579 ( .A(n727), .B(n726), .Z(n729) );
  XOR U1580 ( .A(x[259]), .B(y[259]), .Z(n423) );
  XOR U1581 ( .A(x[255]), .B(y[255]), .Z(n420) );
  XOR U1582 ( .A(x[257]), .B(y[257]), .Z(n421) );
  XOR U1583 ( .A(n420), .B(n421), .Z(n422) );
  XNOR U1584 ( .A(n423), .B(n422), .Z(n144) );
  XOR U1585 ( .A(x[265]), .B(y[265]), .Z(n447) );
  XOR U1586 ( .A(x[261]), .B(y[261]), .Z(n444) );
  XOR U1587 ( .A(x[263]), .B(y[263]), .Z(n445) );
  XOR U1588 ( .A(n444), .B(n445), .Z(n446) );
  XNOR U1589 ( .A(n447), .B(n446), .Z(n142) );
  XOR U1590 ( .A(x[271]), .B(y[271]), .Z(n435) );
  XOR U1591 ( .A(x[267]), .B(y[267]), .Z(n432) );
  XOR U1592 ( .A(x[269]), .B(y[269]), .Z(n433) );
  XOR U1593 ( .A(n432), .B(n433), .Z(n434) );
  XNOR U1594 ( .A(n435), .B(n434), .Z(n141) );
  XOR U1595 ( .A(n142), .B(n141), .Z(n143) );
  XOR U1596 ( .A(n144), .B(n143), .Z(n728) );
  XOR U1597 ( .A(n729), .B(n728), .Z(n1168) );
  XOR U1598 ( .A(x[277]), .B(y[277]), .Z(n441) );
  XOR U1599 ( .A(x[273]), .B(y[273]), .Z(n438) );
  XOR U1600 ( .A(x[275]), .B(y[275]), .Z(n439) );
  XOR U1601 ( .A(n438), .B(n439), .Z(n440) );
  XNOR U1602 ( .A(n441), .B(n440), .Z(n229) );
  XOR U1603 ( .A(x[283]), .B(y[283]), .Z(n561) );
  XOR U1604 ( .A(x[279]), .B(y[279]), .Z(n558) );
  XOR U1605 ( .A(x[281]), .B(y[281]), .Z(n559) );
  XOR U1606 ( .A(n558), .B(n559), .Z(n560) );
  XNOR U1607 ( .A(n561), .B(n560), .Z(n227) );
  XOR U1608 ( .A(x[289]), .B(y[289]), .Z(n549) );
  XOR U1609 ( .A(x[285]), .B(y[285]), .Z(n546) );
  XOR U1610 ( .A(x[287]), .B(y[287]), .Z(n547) );
  XOR U1611 ( .A(n546), .B(n547), .Z(n548) );
  XNOR U1612 ( .A(n549), .B(n548), .Z(n226) );
  XOR U1613 ( .A(n227), .B(n226), .Z(n228) );
  XOR U1614 ( .A(n229), .B(n228), .Z(n63) );
  XOR U1615 ( .A(x[361]), .B(y[361]), .Z(n1144) );
  XOR U1616 ( .A(x[359]), .B(y[359]), .Z(n1141) );
  XNOR U1617 ( .A(x[411]), .B(y[411]), .Z(n1142) );
  XNOR U1618 ( .A(n1144), .B(n1143), .Z(n259) );
  XOR U1619 ( .A(x[365]), .B(y[365]), .Z(n802) );
  XOR U1620 ( .A(x[363]), .B(y[363]), .Z(n799) );
  XOR U1621 ( .A(x[409]), .B(y[409]), .Z(n800) );
  XOR U1622 ( .A(n799), .B(n800), .Z(n801) );
  XNOR U1623 ( .A(n802), .B(n801), .Z(n257) );
  XOR U1624 ( .A(x[369]), .B(y[369]), .Z(n790) );
  XOR U1625 ( .A(x[367]), .B(y[367]), .Z(n787) );
  XOR U1626 ( .A(x[383]), .B(y[383]), .Z(n788) );
  XOR U1627 ( .A(n787), .B(n788), .Z(n789) );
  XNOR U1628 ( .A(n790), .B(n789), .Z(n256) );
  XOR U1629 ( .A(n257), .B(n256), .Z(n258) );
  XOR U1630 ( .A(n259), .B(n258), .Z(n62) );
  XOR U1631 ( .A(n63), .B(n62), .Z(n65) );
  XOR U1632 ( .A(x[295]), .B(y[295]), .Z(n555) );
  XOR U1633 ( .A(x[291]), .B(y[291]), .Z(n552) );
  XOR U1634 ( .A(x[293]), .B(y[293]), .Z(n553) );
  XOR U1635 ( .A(n552), .B(n553), .Z(n554) );
  XNOR U1636 ( .A(n555), .B(n554), .Z(n351) );
  XOR U1637 ( .A(x[301]), .B(y[301]), .Z(n1114) );
  XOR U1638 ( .A(x[297]), .B(y[297]), .Z(n1111) );
  XOR U1639 ( .A(x[299]), .B(y[299]), .Z(n1112) );
  XOR U1640 ( .A(n1111), .B(n1112), .Z(n1113) );
  XNOR U1641 ( .A(n1114), .B(n1113), .Z(n349) );
  XOR U1642 ( .A(x[307]), .B(y[307]), .Z(n1102) );
  XOR U1643 ( .A(x[303]), .B(y[303]), .Z(n1099) );
  XOR U1644 ( .A(x[305]), .B(y[305]), .Z(n1100) );
  XOR U1645 ( .A(n1099), .B(n1100), .Z(n1101) );
  XNOR U1646 ( .A(n1102), .B(n1101), .Z(n348) );
  XOR U1647 ( .A(n349), .B(n348), .Z(n350) );
  XOR U1648 ( .A(n351), .B(n350), .Z(n64) );
  XOR U1649 ( .A(n65), .B(n64), .Z(n1166) );
  XOR U1650 ( .A(x[337]), .B(y[337]), .Z(n1000) );
  XOR U1651 ( .A(x[335]), .B(y[335]), .Z(n997) );
  XOR U1652 ( .A(x[423]), .B(y[423]), .Z(n998) );
  XOR U1653 ( .A(n997), .B(n998), .Z(n999) );
  XNOR U1654 ( .A(n1000), .B(n999), .Z(n471) );
  XOR U1655 ( .A(x[341]), .B(y[341]), .Z(n922) );
  XOR U1656 ( .A(x[339]), .B(y[339]), .Z(n919) );
  XNOR U1657 ( .A(x[421]), .B(y[421]), .Z(n920) );
  XNOR U1658 ( .A(n922), .B(n921), .Z(n469) );
  XOR U1659 ( .A(x[345]), .B(y[345]), .Z(n910) );
  XOR U1660 ( .A(x[343]), .B(y[343]), .Z(n907) );
  XNOR U1661 ( .A(x[419]), .B(y[419]), .Z(n908) );
  XNOR U1662 ( .A(n910), .B(n909), .Z(n468) );
  XOR U1663 ( .A(n469), .B(n468), .Z(n470) );
  XOR U1664 ( .A(n471), .B(n470), .Z(n1165) );
  XOR U1665 ( .A(n1166), .B(n1165), .Z(n1167) );
  XOR U1666 ( .A(n1168), .B(n1167), .Z(n528) );
  XNOR U1667 ( .A(n529), .B(n528), .Z(n530) );
  XNOR U1668 ( .A(n531), .B(n530), .Z(o[0]) );
  NAND U1669 ( .A(n51), .B(n50), .Z(n55) );
  NAND U1670 ( .A(n53), .B(n52), .Z(n54) );
  AND U1671 ( .A(n55), .B(n54), .Z(n2274) );
  NAND U1672 ( .A(n57), .B(n56), .Z(n61) );
  NAND U1673 ( .A(n59), .B(n58), .Z(n60) );
  NAND U1674 ( .A(n61), .B(n60), .Z(n1972) );
  NAND U1675 ( .A(n63), .B(n62), .Z(n67) );
  NAND U1676 ( .A(n65), .B(n64), .Z(n66) );
  NAND U1677 ( .A(n67), .B(n66), .Z(n1971) );
  NAND U1678 ( .A(n69), .B(n68), .Z(n73) );
  NAND U1679 ( .A(n71), .B(n70), .Z(n72) );
  AND U1680 ( .A(n73), .B(n72), .Z(n1685) );
  NAND U1681 ( .A(n75), .B(n74), .Z(n79) );
  NAND U1682 ( .A(n77), .B(n76), .Z(n78) );
  AND U1683 ( .A(n79), .B(n78), .Z(n1686) );
  XOR U1684 ( .A(n1685), .B(n1686), .Z(n1688) );
  NAND U1685 ( .A(n81), .B(n80), .Z(n85) );
  NAND U1686 ( .A(n83), .B(n82), .Z(n84) );
  AND U1687 ( .A(n85), .B(n84), .Z(n1687) );
  XNOR U1688 ( .A(n1688), .B(n1687), .Z(n1850) );
  NAND U1689 ( .A(n87), .B(n86), .Z(n91) );
  NAND U1690 ( .A(n89), .B(n88), .Z(n90) );
  AND U1691 ( .A(n91), .B(n90), .Z(n2242) );
  NANDN U1692 ( .A(n93), .B(n92), .Z(n97) );
  NAND U1693 ( .A(n95), .B(n94), .Z(n96) );
  AND U1694 ( .A(n97), .B(n96), .Z(n2243) );
  XOR U1695 ( .A(n2242), .B(n2243), .Z(n2245) );
  NANDN U1696 ( .A(n99), .B(n98), .Z(n103) );
  NAND U1697 ( .A(n101), .B(n100), .Z(n102) );
  AND U1698 ( .A(n103), .B(n102), .Z(n2244) );
  XNOR U1699 ( .A(n2245), .B(n2244), .Z(n1848) );
  NAND U1700 ( .A(n105), .B(n104), .Z(n109) );
  NAND U1701 ( .A(n107), .B(n106), .Z(n108) );
  AND U1702 ( .A(n109), .B(n108), .Z(n1847) );
  XOR U1703 ( .A(n1848), .B(n1847), .Z(n1849) );
  XOR U1704 ( .A(n1850), .B(n1849), .Z(n1970) );
  XOR U1705 ( .A(n1971), .B(n1970), .Z(n110) );
  XOR U1706 ( .A(n1972), .B(n110), .Z(n2008) );
  NAND U1707 ( .A(n112), .B(n111), .Z(n116) );
  NAND U1708 ( .A(n114), .B(n113), .Z(n115) );
  AND U1709 ( .A(n116), .B(n115), .Z(n2137) );
  NAND U1710 ( .A(n118), .B(n117), .Z(n122) );
  NAND U1711 ( .A(n120), .B(n119), .Z(n121) );
  AND U1712 ( .A(n122), .B(n121), .Z(n2104) );
  NANDN U1713 ( .A(n124), .B(n123), .Z(n128) );
  NAND U1714 ( .A(n126), .B(n125), .Z(n127) );
  AND U1715 ( .A(n128), .B(n127), .Z(n2105) );
  XOR U1716 ( .A(n2104), .B(n2105), .Z(n2107) );
  NANDN U1717 ( .A(n130), .B(n129), .Z(n134) );
  NAND U1718 ( .A(n132), .B(n131), .Z(n133) );
  AND U1719 ( .A(n134), .B(n133), .Z(n2106) );
  XNOR U1720 ( .A(n2107), .B(n2106), .Z(n2135) );
  NAND U1721 ( .A(n136), .B(n135), .Z(n140) );
  NAND U1722 ( .A(n138), .B(n137), .Z(n139) );
  AND U1723 ( .A(n140), .B(n139), .Z(n2134) );
  XOR U1724 ( .A(n2135), .B(n2134), .Z(n2136) );
  XNOR U1725 ( .A(n2137), .B(n2136), .Z(n1954) );
  NAND U1726 ( .A(n142), .B(n141), .Z(n146) );
  NAND U1727 ( .A(n144), .B(n143), .Z(n145) );
  AND U1728 ( .A(n146), .B(n145), .Z(n2048) );
  NANDN U1729 ( .A(n148), .B(n147), .Z(n152) );
  NAND U1730 ( .A(n150), .B(n149), .Z(n151) );
  AND U1731 ( .A(n152), .B(n151), .Z(n2074) );
  NAND U1732 ( .A(n154), .B(n153), .Z(n158) );
  NAND U1733 ( .A(n156), .B(n155), .Z(n157) );
  NAND U1734 ( .A(n158), .B(n157), .Z(n2075) );
  NAND U1735 ( .A(n160), .B(n159), .Z(n164) );
  NAND U1736 ( .A(n162), .B(n161), .Z(n163) );
  AND U1737 ( .A(n164), .B(n163), .Z(n2076) );
  XNOR U1738 ( .A(n2077), .B(n2076), .Z(n2046) );
  NAND U1739 ( .A(n166), .B(n165), .Z(n170) );
  NAND U1740 ( .A(n168), .B(n167), .Z(n169) );
  AND U1741 ( .A(n170), .B(n169), .Z(n2045) );
  XOR U1742 ( .A(n2046), .B(n2045), .Z(n2047) );
  XNOR U1743 ( .A(n2048), .B(n2047), .Z(n1953) );
  NAND U1744 ( .A(n172), .B(n171), .Z(n176) );
  NAND U1745 ( .A(n174), .B(n173), .Z(n175) );
  AND U1746 ( .A(n176), .B(n175), .Z(n1604) );
  NAND U1747 ( .A(n178), .B(n177), .Z(n182) );
  NAND U1748 ( .A(n180), .B(n179), .Z(n181) );
  AND U1749 ( .A(n182), .B(n181), .Z(n2212) );
  NAND U1750 ( .A(n184), .B(n183), .Z(n188) );
  NAND U1751 ( .A(n186), .B(n185), .Z(n187) );
  NAND U1752 ( .A(n188), .B(n187), .Z(n2213) );
  NAND U1753 ( .A(n190), .B(n189), .Z(n194) );
  NAND U1754 ( .A(n192), .B(n191), .Z(n193) );
  AND U1755 ( .A(n194), .B(n193), .Z(n2214) );
  XNOR U1756 ( .A(n2215), .B(n2214), .Z(n1602) );
  NAND U1757 ( .A(n196), .B(n195), .Z(n200) );
  NAND U1758 ( .A(n198), .B(n197), .Z(n199) );
  AND U1759 ( .A(n200), .B(n199), .Z(n1601) );
  XOR U1760 ( .A(n1602), .B(n1601), .Z(n1603) );
  XOR U1761 ( .A(n1604), .B(n1603), .Z(n1952) );
  XOR U1762 ( .A(n1953), .B(n1952), .Z(n201) );
  XNOR U1763 ( .A(n1954), .B(n201), .Z(n2006) );
  NAND U1764 ( .A(n203), .B(n202), .Z(n207) );
  NAND U1765 ( .A(n205), .B(n204), .Z(n206) );
  AND U1766 ( .A(n207), .B(n206), .Z(n2089) );
  NAND U1767 ( .A(n209), .B(n208), .Z(n213) );
  NAND U1768 ( .A(n211), .B(n210), .Z(n212) );
  AND U1769 ( .A(n213), .B(n212), .Z(n2068) );
  NANDN U1770 ( .A(n215), .B(n214), .Z(n219) );
  NAND U1771 ( .A(n217), .B(n216), .Z(n218) );
  AND U1772 ( .A(n219), .B(n218), .Z(n2069) );
  XOR U1773 ( .A(n2068), .B(n2069), .Z(n2071) );
  NAND U1774 ( .A(n221), .B(n220), .Z(n225) );
  NAND U1775 ( .A(n223), .B(n222), .Z(n224) );
  AND U1776 ( .A(n225), .B(n224), .Z(n2070) );
  XNOR U1777 ( .A(n2071), .B(n2070), .Z(n2087) );
  NAND U1778 ( .A(n227), .B(n226), .Z(n231) );
  NAND U1779 ( .A(n229), .B(n228), .Z(n230) );
  AND U1780 ( .A(n231), .B(n230), .Z(n2086) );
  XOR U1781 ( .A(n2087), .B(n2086), .Z(n2088) );
  XNOR U1782 ( .A(n2089), .B(n2088), .Z(n1961) );
  NAND U1783 ( .A(n233), .B(n232), .Z(n237) );
  NAND U1784 ( .A(n235), .B(n234), .Z(n236) );
  AND U1785 ( .A(n237), .B(n236), .Z(n1586) );
  NAND U1786 ( .A(n239), .B(n238), .Z(n243) );
  NAND U1787 ( .A(n241), .B(n240), .Z(n242) );
  AND U1788 ( .A(n243), .B(n242), .Z(n2206) );
  NAND U1789 ( .A(n245), .B(n244), .Z(n249) );
  NAND U1790 ( .A(n247), .B(n246), .Z(n248) );
  AND U1791 ( .A(n249), .B(n248), .Z(n2207) );
  XOR U1792 ( .A(n2206), .B(n2207), .Z(n2209) );
  NAND U1793 ( .A(n251), .B(n250), .Z(n255) );
  NAND U1794 ( .A(n253), .B(n252), .Z(n254) );
  AND U1795 ( .A(n255), .B(n254), .Z(n2208) );
  XNOR U1796 ( .A(n2209), .B(n2208), .Z(n1584) );
  NAND U1797 ( .A(n257), .B(n256), .Z(n261) );
  NAND U1798 ( .A(n259), .B(n258), .Z(n260) );
  AND U1799 ( .A(n261), .B(n260), .Z(n1583) );
  XOR U1800 ( .A(n1584), .B(n1583), .Z(n1585) );
  XNOR U1801 ( .A(n1586), .B(n1585), .Z(n1959) );
  NAND U1802 ( .A(n263), .B(n262), .Z(n267) );
  NAND U1803 ( .A(n265), .B(n264), .Z(n266) );
  NAND U1804 ( .A(n267), .B(n266), .Z(n1958) );
  XOR U1805 ( .A(n1959), .B(n1958), .Z(n1960) );
  XOR U1806 ( .A(n1961), .B(n1960), .Z(n2007) );
  XOR U1807 ( .A(n2006), .B(n2007), .Z(n268) );
  XNOR U1808 ( .A(n2008), .B(n268), .Z(n2272) );
  NAND U1809 ( .A(n270), .B(n269), .Z(n274) );
  NAND U1810 ( .A(n272), .B(n271), .Z(n273) );
  AND U1811 ( .A(n274), .B(n273), .Z(n1766) );
  NAND U1812 ( .A(n276), .B(n275), .Z(n280) );
  NAND U1813 ( .A(n278), .B(n277), .Z(n279) );
  AND U1814 ( .A(n280), .B(n279), .Z(n1613) );
  NAND U1815 ( .A(n282), .B(n281), .Z(n286) );
  NAND U1816 ( .A(n284), .B(n283), .Z(n285) );
  NAND U1817 ( .A(n286), .B(n285), .Z(n1614) );
  NAND U1818 ( .A(n288), .B(n287), .Z(n292) );
  NAND U1819 ( .A(n290), .B(n289), .Z(n291) );
  AND U1820 ( .A(n292), .B(n291), .Z(n1615) );
  XNOR U1821 ( .A(n1616), .B(n1615), .Z(n1764) );
  NAND U1822 ( .A(n294), .B(n293), .Z(n298) );
  NAND U1823 ( .A(n296), .B(n295), .Z(n297) );
  AND U1824 ( .A(n298), .B(n297), .Z(n1763) );
  XOR U1825 ( .A(n1764), .B(n1763), .Z(n1765) );
  XOR U1826 ( .A(n1766), .B(n1765), .Z(n2020) );
  NAND U1827 ( .A(n300), .B(n299), .Z(n304) );
  NAND U1828 ( .A(n302), .B(n301), .Z(n303) );
  NAND U1829 ( .A(n304), .B(n303), .Z(n2018) );
  NAND U1830 ( .A(n306), .B(n305), .Z(n310) );
  NAND U1831 ( .A(n308), .B(n307), .Z(n309) );
  AND U1832 ( .A(n310), .B(n309), .Z(n1628) );
  NAND U1833 ( .A(n312), .B(n311), .Z(n316) );
  NAND U1834 ( .A(n314), .B(n313), .Z(n315) );
  AND U1835 ( .A(n316), .B(n315), .Z(n1607) );
  NAND U1836 ( .A(n318), .B(n317), .Z(n322) );
  NAND U1837 ( .A(n320), .B(n319), .Z(n321) );
  NAND U1838 ( .A(n322), .B(n321), .Z(n1608) );
  NAND U1839 ( .A(n324), .B(n323), .Z(n328) );
  NAND U1840 ( .A(n326), .B(n325), .Z(n327) );
  AND U1841 ( .A(n328), .B(n327), .Z(n1609) );
  XNOR U1842 ( .A(n1610), .B(n1609), .Z(n1626) );
  NAND U1843 ( .A(n330), .B(n329), .Z(n334) );
  NAND U1844 ( .A(n332), .B(n331), .Z(n333) );
  AND U1845 ( .A(n334), .B(n333), .Z(n1625) );
  XOR U1846 ( .A(n1626), .B(n1625), .Z(n1627) );
  XOR U1847 ( .A(n1628), .B(n1627), .Z(n2019) );
  XOR U1848 ( .A(n2018), .B(n2019), .Z(n335) );
  XOR U1849 ( .A(n2020), .B(n335), .Z(n1861) );
  NAND U1850 ( .A(n337), .B(n336), .Z(n341) );
  NAND U1851 ( .A(n339), .B(n338), .Z(n340) );
  NAND U1852 ( .A(n341), .B(n340), .Z(n1860) );
  NAND U1853 ( .A(n343), .B(n342), .Z(n347) );
  NAND U1854 ( .A(n345), .B(n344), .Z(n346) );
  NAND U1855 ( .A(n347), .B(n346), .Z(n1859) );
  XOR U1856 ( .A(n1860), .B(n1859), .Z(n1862) );
  XNOR U1857 ( .A(n1861), .B(n1862), .Z(n1795) );
  NAND U1858 ( .A(n349), .B(n348), .Z(n353) );
  NAND U1859 ( .A(n351), .B(n350), .Z(n352) );
  AND U1860 ( .A(n353), .B(n352), .Z(n2179) );
  NAND U1861 ( .A(n355), .B(n354), .Z(n359) );
  NAND U1862 ( .A(n357), .B(n356), .Z(n358) );
  AND U1863 ( .A(n359), .B(n358), .Z(n2092) );
  NANDN U1864 ( .A(n361), .B(n360), .Z(n365) );
  NAND U1865 ( .A(n363), .B(n362), .Z(n364) );
  AND U1866 ( .A(n365), .B(n364), .Z(n2093) );
  XOR U1867 ( .A(n2092), .B(n2093), .Z(n2095) );
  NAND U1868 ( .A(n367), .B(n366), .Z(n371) );
  NAND U1869 ( .A(n369), .B(n368), .Z(n370) );
  AND U1870 ( .A(n371), .B(n370), .Z(n2094) );
  XNOR U1871 ( .A(n2095), .B(n2094), .Z(n2177) );
  NAND U1872 ( .A(n373), .B(n372), .Z(n377) );
  NAND U1873 ( .A(n375), .B(n374), .Z(n376) );
  AND U1874 ( .A(n377), .B(n376), .Z(n2176) );
  XOR U1875 ( .A(n2177), .B(n2176), .Z(n2178) );
  XNOR U1876 ( .A(n2179), .B(n2178), .Z(n2251) );
  NAND U1877 ( .A(n379), .B(n378), .Z(n383) );
  NAND U1878 ( .A(n381), .B(n380), .Z(n382) );
  AND U1879 ( .A(n383), .B(n382), .Z(n1724) );
  NANDN U1880 ( .A(n385), .B(n384), .Z(n389) );
  NAND U1881 ( .A(n387), .B(n386), .Z(n388) );
  AND U1882 ( .A(n389), .B(n388), .Z(n2182) );
  NAND U1883 ( .A(n391), .B(n390), .Z(n395) );
  NAND U1884 ( .A(n393), .B(n392), .Z(n394) );
  NAND U1885 ( .A(n395), .B(n394), .Z(n2183) );
  NAND U1886 ( .A(n397), .B(n396), .Z(n401) );
  NAND U1887 ( .A(n399), .B(n398), .Z(n400) );
  AND U1888 ( .A(n401), .B(n400), .Z(n2184) );
  XNOR U1889 ( .A(n2185), .B(n2184), .Z(n1722) );
  NAND U1890 ( .A(n403), .B(n402), .Z(n407) );
  NAND U1891 ( .A(n405), .B(n404), .Z(n406) );
  AND U1892 ( .A(n407), .B(n406), .Z(n1721) );
  XOR U1893 ( .A(n1722), .B(n1721), .Z(n1723) );
  XNOR U1894 ( .A(n1724), .B(n1723), .Z(n2249) );
  NAND U1895 ( .A(n409), .B(n408), .Z(n413) );
  NAND U1896 ( .A(n411), .B(n410), .Z(n412) );
  NAND U1897 ( .A(n413), .B(n412), .Z(n2248) );
  XOR U1898 ( .A(n2249), .B(n2248), .Z(n2250) );
  XNOR U1899 ( .A(n2251), .B(n2250), .Z(n1793) );
  NAND U1900 ( .A(n415), .B(n414), .Z(n419) );
  NAND U1901 ( .A(n417), .B(n416), .Z(n418) );
  AND U1902 ( .A(n419), .B(n418), .Z(n2158) );
  NAND U1903 ( .A(n421), .B(n420), .Z(n425) );
  NAND U1904 ( .A(n423), .B(n422), .Z(n424) );
  NAND U1905 ( .A(n425), .B(n424), .Z(n2159) );
  NAND U1906 ( .A(n427), .B(n426), .Z(n431) );
  NAND U1907 ( .A(n429), .B(n428), .Z(n430) );
  AND U1908 ( .A(n431), .B(n430), .Z(n2160) );
  XNOR U1909 ( .A(n2161), .B(n2160), .Z(n1946) );
  NAND U1910 ( .A(n433), .B(n432), .Z(n437) );
  NAND U1911 ( .A(n435), .B(n434), .Z(n436) );
  AND U1912 ( .A(n437), .B(n436), .Z(n2164) );
  NAND U1913 ( .A(n439), .B(n438), .Z(n443) );
  NAND U1914 ( .A(n441), .B(n440), .Z(n442) );
  NAND U1915 ( .A(n443), .B(n442), .Z(n2165) );
  NAND U1916 ( .A(n445), .B(n444), .Z(n449) );
  NAND U1917 ( .A(n447), .B(n446), .Z(n448) );
  AND U1918 ( .A(n449), .B(n448), .Z(n2166) );
  XNOR U1919 ( .A(n2167), .B(n2166), .Z(n1944) );
  NAND U1920 ( .A(n451), .B(n450), .Z(n455) );
  NAND U1921 ( .A(n453), .B(n452), .Z(n454) );
  AND U1922 ( .A(n455), .B(n454), .Z(n1667) );
  NAND U1923 ( .A(n457), .B(n456), .Z(n461) );
  NAND U1924 ( .A(n459), .B(n458), .Z(n460) );
  NAND U1925 ( .A(n461), .B(n460), .Z(n1668) );
  NAND U1926 ( .A(n463), .B(n462), .Z(n467) );
  NAND U1927 ( .A(n465), .B(n464), .Z(n466) );
  AND U1928 ( .A(n467), .B(n466), .Z(n1669) );
  XNOR U1929 ( .A(n1670), .B(n1669), .Z(n1943) );
  XOR U1930 ( .A(n1944), .B(n1943), .Z(n1945) );
  XOR U1931 ( .A(n1946), .B(n1945), .Z(n2010) );
  NAND U1932 ( .A(n469), .B(n468), .Z(n473) );
  NAND U1933 ( .A(n471), .B(n470), .Z(n472) );
  AND U1934 ( .A(n473), .B(n472), .Z(n2227) );
  NANDN U1935 ( .A(n475), .B(n474), .Z(n479) );
  NAND U1936 ( .A(n477), .B(n476), .Z(n478) );
  AND U1937 ( .A(n479), .B(n478), .Z(n2188) );
  NAND U1938 ( .A(n481), .B(n480), .Z(n485) );
  NAND U1939 ( .A(n483), .B(n482), .Z(n484) );
  NAND U1940 ( .A(n485), .B(n484), .Z(n2189) );
  NAND U1941 ( .A(n487), .B(n486), .Z(n491) );
  NAND U1942 ( .A(n489), .B(n488), .Z(n490) );
  AND U1943 ( .A(n491), .B(n490), .Z(n2190) );
  XNOR U1944 ( .A(n2191), .B(n2190), .Z(n2225) );
  NAND U1945 ( .A(n493), .B(n492), .Z(n497) );
  NAND U1946 ( .A(n495), .B(n494), .Z(n496) );
  AND U1947 ( .A(n497), .B(n496), .Z(n2224) );
  XOR U1948 ( .A(n2225), .B(n2224), .Z(n2226) );
  XOR U1949 ( .A(n2227), .B(n2226), .Z(n2009) );
  XOR U1950 ( .A(n2010), .B(n2009), .Z(n2012) );
  NAND U1951 ( .A(n499), .B(n498), .Z(n503) );
  NAND U1952 ( .A(n501), .B(n500), .Z(n502) );
  AND U1953 ( .A(n503), .B(n502), .Z(n1700) );
  NAND U1954 ( .A(n505), .B(n504), .Z(n509) );
  NAND U1955 ( .A(n507), .B(n506), .Z(n508) );
  AND U1956 ( .A(n509), .B(n508), .Z(n2051) );
  NANDN U1957 ( .A(n511), .B(n510), .Z(n515) );
  NAND U1958 ( .A(n513), .B(n512), .Z(n514) );
  AND U1959 ( .A(n515), .B(n514), .Z(n2052) );
  XOR U1960 ( .A(n2051), .B(n2052), .Z(n2054) );
  NAND U1961 ( .A(n517), .B(n516), .Z(n521) );
  NAND U1962 ( .A(n519), .B(n518), .Z(n520) );
  AND U1963 ( .A(n521), .B(n520), .Z(n2053) );
  XNOR U1964 ( .A(n2054), .B(n2053), .Z(n1698) );
  NAND U1965 ( .A(n523), .B(n522), .Z(n527) );
  NAND U1966 ( .A(n525), .B(n524), .Z(n526) );
  AND U1967 ( .A(n527), .B(n526), .Z(n1697) );
  XOR U1968 ( .A(n1698), .B(n1697), .Z(n1699) );
  XOR U1969 ( .A(n1700), .B(n1699), .Z(n2011) );
  XOR U1970 ( .A(n2012), .B(n2011), .Z(n1794) );
  XOR U1971 ( .A(n1793), .B(n1794), .Z(n1796) );
  XNOR U1972 ( .A(n1795), .B(n1796), .Z(n2271) );
  XOR U1973 ( .A(n2272), .B(n2271), .Z(n2273) );
  XNOR U1974 ( .A(n2274), .B(n2273), .Z(n2279) );
  NANDN U1975 ( .A(n529), .B(n528), .Z(n533) );
  NAND U1976 ( .A(n531), .B(n530), .Z(n532) );
  AND U1977 ( .A(n533), .B(n532), .Z(n2278) );
  NAND U1978 ( .A(n535), .B(n534), .Z(n539) );
  NAND U1979 ( .A(n537), .B(n536), .Z(n538) );
  NAND U1980 ( .A(n539), .B(n538), .Z(n1997) );
  NAND U1981 ( .A(n541), .B(n540), .Z(n545) );
  NAND U1982 ( .A(n543), .B(n542), .Z(n544) );
  NAND U1983 ( .A(n545), .B(n544), .Z(n1995) );
  NAND U1984 ( .A(n547), .B(n546), .Z(n551) );
  NAND U1985 ( .A(n549), .B(n548), .Z(n550) );
  AND U1986 ( .A(n551), .B(n550), .Z(n1703) );
  NAND U1987 ( .A(n553), .B(n552), .Z(n557) );
  NAND U1988 ( .A(n555), .B(n554), .Z(n556) );
  AND U1989 ( .A(n557), .B(n556), .Z(n1704) );
  XOR U1990 ( .A(n1703), .B(n1704), .Z(n1706) );
  NAND U1991 ( .A(n559), .B(n558), .Z(n563) );
  NAND U1992 ( .A(n561), .B(n560), .Z(n562) );
  AND U1993 ( .A(n563), .B(n562), .Z(n1705) );
  XOR U1994 ( .A(n1706), .B(n1705), .Z(n1880) );
  NAND U1995 ( .A(n565), .B(n564), .Z(n569) );
  NAND U1996 ( .A(n567), .B(n566), .Z(n568) );
  AND U1997 ( .A(n569), .B(n568), .Z(n1727) );
  NAND U1998 ( .A(n571), .B(n570), .Z(n575) );
  NAND U1999 ( .A(n573), .B(n572), .Z(n574) );
  AND U2000 ( .A(n575), .B(n574), .Z(n1728) );
  XOR U2001 ( .A(n1727), .B(n1728), .Z(n1730) );
  NAND U2002 ( .A(n577), .B(n576), .Z(n581) );
  NAND U2003 ( .A(n579), .B(n578), .Z(n580) );
  AND U2004 ( .A(n581), .B(n580), .Z(n1729) );
  XNOR U2005 ( .A(n1730), .B(n1729), .Z(n1878) );
  NANDN U2006 ( .A(n583), .B(n582), .Z(n587) );
  NAND U2007 ( .A(n585), .B(n584), .Z(n586) );
  AND U2008 ( .A(n587), .B(n586), .Z(n1661) );
  NAND U2009 ( .A(n589), .B(n588), .Z(n593) );
  NAND U2010 ( .A(n591), .B(n590), .Z(n592) );
  AND U2011 ( .A(n593), .B(n592), .Z(n1662) );
  XOR U2012 ( .A(n1661), .B(n1662), .Z(n1664) );
  NANDN U2013 ( .A(n595), .B(n594), .Z(n599) );
  NAND U2014 ( .A(n597), .B(n596), .Z(n598) );
  AND U2015 ( .A(n599), .B(n598), .Z(n1663) );
  XNOR U2016 ( .A(n1664), .B(n1663), .Z(n1877) );
  XOR U2017 ( .A(n1878), .B(n1877), .Z(n1879) );
  XOR U2018 ( .A(n1880), .B(n1879), .Z(n1994) );
  XOR U2019 ( .A(n1995), .B(n1994), .Z(n1996) );
  XNOR U2020 ( .A(n1997), .B(n1996), .Z(n1951) );
  NAND U2021 ( .A(n601), .B(n600), .Z(n605) );
  NAND U2022 ( .A(n603), .B(n602), .Z(n604) );
  NAND U2023 ( .A(n605), .B(n604), .Z(n2113) );
  NAND U2024 ( .A(n607), .B(n606), .Z(n611) );
  NAND U2025 ( .A(n609), .B(n608), .Z(n610) );
  AND U2026 ( .A(n611), .B(n610), .Z(n2194) );
  NANDN U2027 ( .A(n613), .B(n612), .Z(n617) );
  NAND U2028 ( .A(n615), .B(n614), .Z(n616) );
  NAND U2029 ( .A(n617), .B(n616), .Z(n2195) );
  NANDN U2030 ( .A(n619), .B(n618), .Z(n623) );
  NAND U2031 ( .A(n621), .B(n620), .Z(n622) );
  AND U2032 ( .A(n623), .B(n622), .Z(n2196) );
  XNOR U2033 ( .A(n2197), .B(n2196), .Z(n1832) );
  NAND U2034 ( .A(n625), .B(n624), .Z(n629) );
  NAND U2035 ( .A(n627), .B(n626), .Z(n628) );
  AND U2036 ( .A(n629), .B(n628), .Z(n2236) );
  NANDN U2037 ( .A(n631), .B(n630), .Z(n635) );
  NAND U2038 ( .A(n633), .B(n632), .Z(n634) );
  AND U2039 ( .A(n635), .B(n634), .Z(n2237) );
  XOR U2040 ( .A(n2236), .B(n2237), .Z(n2239) );
  NANDN U2041 ( .A(n637), .B(n636), .Z(n641) );
  NAND U2042 ( .A(n639), .B(n638), .Z(n640) );
  AND U2043 ( .A(n641), .B(n640), .Z(n2238) );
  XNOR U2044 ( .A(n2239), .B(n2238), .Z(n1830) );
  NAND U2045 ( .A(n643), .B(n642), .Z(n647) );
  NAND U2046 ( .A(n645), .B(n644), .Z(n646) );
  AND U2047 ( .A(n647), .B(n646), .Z(n2218) );
  NANDN U2048 ( .A(n649), .B(n648), .Z(n653) );
  NAND U2049 ( .A(n651), .B(n650), .Z(n652) );
  AND U2050 ( .A(n653), .B(n652), .Z(n2219) );
  XOR U2051 ( .A(n2218), .B(n2219), .Z(n2221) );
  NANDN U2052 ( .A(n655), .B(n654), .Z(n659) );
  NAND U2053 ( .A(n657), .B(n656), .Z(n658) );
  AND U2054 ( .A(n659), .B(n658), .Z(n2220) );
  XNOR U2055 ( .A(n2221), .B(n2220), .Z(n1829) );
  XOR U2056 ( .A(n1830), .B(n1829), .Z(n1831) );
  XNOR U2057 ( .A(n1832), .B(n1831), .Z(n2111) );
  NAND U2058 ( .A(n661), .B(n660), .Z(n665) );
  NAND U2059 ( .A(n663), .B(n662), .Z(n664) );
  NAND U2060 ( .A(n665), .B(n664), .Z(n2110) );
  XOR U2061 ( .A(n2111), .B(n2110), .Z(n2112) );
  XNOR U2062 ( .A(n2113), .B(n2112), .Z(n1950) );
  NAND U2063 ( .A(n667), .B(n666), .Z(n671) );
  NAND U2064 ( .A(n669), .B(n668), .Z(n670) );
  NAND U2065 ( .A(n671), .B(n670), .Z(n1967) );
  NAND U2066 ( .A(n673), .B(n672), .Z(n677) );
  NAND U2067 ( .A(n675), .B(n674), .Z(n676) );
  AND U2068 ( .A(n677), .B(n676), .Z(n2080) );
  NAND U2069 ( .A(n679), .B(n678), .Z(n683) );
  NAND U2070 ( .A(n681), .B(n680), .Z(n682) );
  AND U2071 ( .A(n683), .B(n682), .Z(n2081) );
  XOR U2072 ( .A(n2080), .B(n2081), .Z(n2083) );
  NAND U2073 ( .A(n685), .B(n684), .Z(n689) );
  NAND U2074 ( .A(n687), .B(n686), .Z(n688) );
  AND U2075 ( .A(n689), .B(n688), .Z(n2082) );
  XNOR U2076 ( .A(n2083), .B(n2082), .Z(n1814) );
  NANDN U2077 ( .A(n691), .B(n690), .Z(n695) );
  NAND U2078 ( .A(n693), .B(n692), .Z(n694) );
  AND U2079 ( .A(n695), .B(n694), .Z(n2128) );
  NANDN U2080 ( .A(n697), .B(n696), .Z(n701) );
  NAND U2081 ( .A(n699), .B(n698), .Z(n700) );
  NAND U2082 ( .A(n701), .B(n700), .Z(n2129) );
  NANDN U2083 ( .A(n703), .B(n702), .Z(n707) );
  NAND U2084 ( .A(n705), .B(n704), .Z(n706) );
  AND U2085 ( .A(n707), .B(n706), .Z(n2130) );
  XNOR U2086 ( .A(n2131), .B(n2130), .Z(n1812) );
  NAND U2087 ( .A(n709), .B(n708), .Z(n713) );
  NAND U2088 ( .A(n711), .B(n710), .Z(n712) );
  AND U2089 ( .A(n713), .B(n712), .Z(n1619) );
  NANDN U2090 ( .A(n715), .B(n714), .Z(n719) );
  NAND U2091 ( .A(n717), .B(n716), .Z(n718) );
  AND U2092 ( .A(n719), .B(n718), .Z(n1620) );
  XOR U2093 ( .A(n1619), .B(n1620), .Z(n1622) );
  NANDN U2094 ( .A(n721), .B(n720), .Z(n725) );
  NAND U2095 ( .A(n723), .B(n722), .Z(n724) );
  AND U2096 ( .A(n725), .B(n724), .Z(n1621) );
  XNOR U2097 ( .A(n1622), .B(n1621), .Z(n1811) );
  XOR U2098 ( .A(n1812), .B(n1811), .Z(n1813) );
  XNOR U2099 ( .A(n1814), .B(n1813), .Z(n1965) );
  NAND U2100 ( .A(n727), .B(n726), .Z(n731) );
  NAND U2101 ( .A(n729), .B(n728), .Z(n730) );
  NAND U2102 ( .A(n731), .B(n730), .Z(n1964) );
  XOR U2103 ( .A(n1965), .B(n1964), .Z(n1966) );
  XOR U2104 ( .A(n1967), .B(n1966), .Z(n1949) );
  XOR U2105 ( .A(n1950), .B(n1949), .Z(n732) );
  XNOR U2106 ( .A(n1951), .B(n732), .Z(n2261) );
  NAND U2107 ( .A(n734), .B(n733), .Z(n738) );
  NAND U2108 ( .A(n736), .B(n735), .Z(n737) );
  AND U2109 ( .A(n738), .B(n737), .Z(n1673) );
  NAND U2110 ( .A(n740), .B(n739), .Z(n744) );
  NAND U2111 ( .A(n742), .B(n741), .Z(n743) );
  NAND U2112 ( .A(n744), .B(n743), .Z(n1674) );
  NAND U2113 ( .A(n746), .B(n745), .Z(n750) );
  NAND U2114 ( .A(n748), .B(n747), .Z(n749) );
  AND U2115 ( .A(n750), .B(n749), .Z(n1675) );
  XNOR U2116 ( .A(n1676), .B(n1675), .Z(n1938) );
  NAND U2117 ( .A(n752), .B(n751), .Z(n756) );
  NAND U2118 ( .A(n754), .B(n753), .Z(n755) );
  AND U2119 ( .A(n756), .B(n755), .Z(n1937) );
  XOR U2120 ( .A(n1938), .B(n1937), .Z(n1940) );
  NAND U2121 ( .A(n758), .B(n757), .Z(n762) );
  NAND U2122 ( .A(n760), .B(n759), .Z(n761) );
  AND U2123 ( .A(n762), .B(n761), .Z(n2065) );
  NAND U2124 ( .A(n764), .B(n763), .Z(n768) );
  NAND U2125 ( .A(n766), .B(n765), .Z(n767) );
  AND U2126 ( .A(n768), .B(n767), .Z(n2063) );
  XOR U2127 ( .A(n1940), .B(n1939), .Z(n1989) );
  NAND U2128 ( .A(n770), .B(n769), .Z(n774) );
  NAND U2129 ( .A(n772), .B(n771), .Z(n773) );
  AND U2130 ( .A(n774), .B(n773), .Z(n1745) );
  NAND U2131 ( .A(n776), .B(n775), .Z(n780) );
  NAND U2132 ( .A(n778), .B(n777), .Z(n779) );
  NAND U2133 ( .A(n780), .B(n779), .Z(n1746) );
  NAND U2134 ( .A(n782), .B(n781), .Z(n786) );
  NAND U2135 ( .A(n784), .B(n783), .Z(n785) );
  AND U2136 ( .A(n786), .B(n785), .Z(n1747) );
  XNOR U2137 ( .A(n1748), .B(n1747), .Z(n1934) );
  NAND U2138 ( .A(n788), .B(n787), .Z(n792) );
  NAND U2139 ( .A(n790), .B(n789), .Z(n791) );
  AND U2140 ( .A(n792), .B(n791), .Z(n2027) );
  NAND U2141 ( .A(n794), .B(n793), .Z(n798) );
  NAND U2142 ( .A(n796), .B(n795), .Z(n797) );
  AND U2143 ( .A(n798), .B(n797), .Z(n2028) );
  XOR U2144 ( .A(n2027), .B(n2028), .Z(n2030) );
  NAND U2145 ( .A(n800), .B(n799), .Z(n804) );
  NAND U2146 ( .A(n802), .B(n801), .Z(n803) );
  AND U2147 ( .A(n804), .B(n803), .Z(n2029) );
  XNOR U2148 ( .A(n2030), .B(n2029), .Z(n1932) );
  NAND U2149 ( .A(n806), .B(n805), .Z(n810) );
  NAND U2150 ( .A(n808), .B(n807), .Z(n809) );
  AND U2151 ( .A(n810), .B(n809), .Z(n1931) );
  XOR U2152 ( .A(n1932), .B(n1931), .Z(n1933) );
  XOR U2153 ( .A(n1934), .B(n1933), .Z(n1988) );
  XOR U2154 ( .A(n1989), .B(n1988), .Z(n1991) );
  NAND U2155 ( .A(n812), .B(n811), .Z(n816) );
  NAND U2156 ( .A(n814), .B(n813), .Z(n815) );
  AND U2157 ( .A(n816), .B(n815), .Z(n1679) );
  NAND U2158 ( .A(n818), .B(n817), .Z(n822) );
  NAND U2159 ( .A(n820), .B(n819), .Z(n821) );
  AND U2160 ( .A(n822), .B(n821), .Z(n1680) );
  XOR U2161 ( .A(n1679), .B(n1680), .Z(n1682) );
  NAND U2162 ( .A(n824), .B(n823), .Z(n828) );
  NAND U2163 ( .A(n826), .B(n825), .Z(n827) );
  AND U2164 ( .A(n828), .B(n827), .Z(n1681) );
  XNOR U2165 ( .A(n1682), .B(n1681), .Z(n1922) );
  NAND U2166 ( .A(n830), .B(n829), .Z(n834) );
  NAND U2167 ( .A(n832), .B(n831), .Z(n833) );
  AND U2168 ( .A(n834), .B(n833), .Z(n2033) );
  NAND U2169 ( .A(n836), .B(n835), .Z(n840) );
  NAND U2170 ( .A(n838), .B(n837), .Z(n839) );
  AND U2171 ( .A(n840), .B(n839), .Z(n2034) );
  XOR U2172 ( .A(n2033), .B(n2034), .Z(n2036) );
  NAND U2173 ( .A(n842), .B(n841), .Z(n846) );
  NAND U2174 ( .A(n844), .B(n843), .Z(n845) );
  AND U2175 ( .A(n846), .B(n845), .Z(n2035) );
  XNOR U2176 ( .A(n2036), .B(n2035), .Z(n1920) );
  NAND U2177 ( .A(n848), .B(n847), .Z(n852) );
  NAND U2178 ( .A(n850), .B(n849), .Z(n851) );
  AND U2179 ( .A(n852), .B(n851), .Z(n1751) );
  NAND U2180 ( .A(n854), .B(n853), .Z(n858) );
  NAND U2181 ( .A(n856), .B(n855), .Z(n857) );
  AND U2182 ( .A(n858), .B(n857), .Z(n1752) );
  XOR U2183 ( .A(n1751), .B(n1752), .Z(n1754) );
  NAND U2184 ( .A(n860), .B(n859), .Z(n864) );
  NAND U2185 ( .A(n862), .B(n861), .Z(n863) );
  AND U2186 ( .A(n864), .B(n863), .Z(n1753) );
  XNOR U2187 ( .A(n1754), .B(n1753), .Z(n1919) );
  XOR U2188 ( .A(n1920), .B(n1919), .Z(n1921) );
  XOR U2189 ( .A(n1922), .B(n1921), .Z(n1990) );
  XOR U2190 ( .A(n1991), .B(n1990), .Z(n1562) );
  NAND U2191 ( .A(n866), .B(n865), .Z(n870) );
  NAND U2192 ( .A(n868), .B(n867), .Z(n869) );
  AND U2193 ( .A(n870), .B(n869), .Z(n2170) );
  NAND U2194 ( .A(n872), .B(n871), .Z(n876) );
  NAND U2195 ( .A(n874), .B(n873), .Z(n875) );
  NAND U2196 ( .A(n876), .B(n875), .Z(n2171) );
  NAND U2197 ( .A(n878), .B(n877), .Z(n882) );
  NAND U2198 ( .A(n880), .B(n879), .Z(n881) );
  AND U2199 ( .A(n882), .B(n881), .Z(n2172) );
  XNOR U2200 ( .A(n2173), .B(n2172), .Z(n1898) );
  NAND U2201 ( .A(n884), .B(n883), .Z(n888) );
  NAND U2202 ( .A(n886), .B(n885), .Z(n887) );
  AND U2203 ( .A(n888), .B(n887), .Z(n1733) );
  NAND U2204 ( .A(n890), .B(n889), .Z(n894) );
  NAND U2205 ( .A(n892), .B(n891), .Z(n893) );
  NAND U2206 ( .A(n894), .B(n893), .Z(n1734) );
  NAND U2207 ( .A(n896), .B(n895), .Z(n900) );
  NAND U2208 ( .A(n898), .B(n897), .Z(n899) );
  AND U2209 ( .A(n900), .B(n899), .Z(n1735) );
  XNOR U2210 ( .A(n1736), .B(n1735), .Z(n1896) );
  NAND U2211 ( .A(n902), .B(n901), .Z(n906) );
  NAND U2212 ( .A(n904), .B(n903), .Z(n905) );
  AND U2213 ( .A(n906), .B(n905), .Z(n1895) );
  XOR U2214 ( .A(n1896), .B(n1895), .Z(n1897) );
  XOR U2215 ( .A(n1898), .B(n1897), .Z(n1985) );
  NANDN U2216 ( .A(n908), .B(n907), .Z(n912) );
  NAND U2217 ( .A(n910), .B(n909), .Z(n911) );
  AND U2218 ( .A(n912), .B(n911), .Z(n2152) );
  NANDN U2219 ( .A(n914), .B(n913), .Z(n918) );
  NAND U2220 ( .A(n916), .B(n915), .Z(n917) );
  AND U2221 ( .A(n918), .B(n917), .Z(n2153) );
  XOR U2222 ( .A(n2152), .B(n2153), .Z(n2155) );
  NANDN U2223 ( .A(n920), .B(n919), .Z(n924) );
  NAND U2224 ( .A(n922), .B(n921), .Z(n923) );
  AND U2225 ( .A(n924), .B(n923), .Z(n2154) );
  XOR U2226 ( .A(n2155), .B(n2154), .Z(n1910) );
  NAND U2227 ( .A(n926), .B(n925), .Z(n930) );
  NAND U2228 ( .A(n928), .B(n927), .Z(n929) );
  AND U2229 ( .A(n930), .B(n929), .Z(n1908) );
  NAND U2230 ( .A(n932), .B(n931), .Z(n936) );
  NAND U2231 ( .A(n934), .B(n933), .Z(n935) );
  AND U2232 ( .A(n936), .B(n935), .Z(n2098) );
  NAND U2233 ( .A(n938), .B(n937), .Z(n942) );
  NAND U2234 ( .A(n940), .B(n939), .Z(n941) );
  AND U2235 ( .A(n942), .B(n941), .Z(n2099) );
  XOR U2236 ( .A(n2098), .B(n2099), .Z(n2101) );
  NAND U2237 ( .A(n944), .B(n943), .Z(n948) );
  NAND U2238 ( .A(n946), .B(n945), .Z(n947) );
  AND U2239 ( .A(n948), .B(n947), .Z(n2100) );
  XNOR U2240 ( .A(n2101), .B(n2100), .Z(n1907) );
  NAND U2241 ( .A(n950), .B(n949), .Z(n954) );
  NAND U2242 ( .A(n952), .B(n951), .Z(n953) );
  AND U2243 ( .A(n954), .B(n953), .Z(n2039) );
  NAND U2244 ( .A(n956), .B(n955), .Z(n960) );
  NAND U2245 ( .A(n958), .B(n957), .Z(n959) );
  NAND U2246 ( .A(n960), .B(n959), .Z(n2040) );
  NAND U2247 ( .A(n962), .B(n961), .Z(n966) );
  NAND U2248 ( .A(n964), .B(n963), .Z(n965) );
  AND U2249 ( .A(n966), .B(n965), .Z(n2041) );
  XNOR U2250 ( .A(n2042), .B(n2041), .Z(n1886) );
  NAND U2251 ( .A(n968), .B(n967), .Z(n972) );
  NAND U2252 ( .A(n970), .B(n969), .Z(n971) );
  AND U2253 ( .A(n972), .B(n971), .Z(n2140) );
  NAND U2254 ( .A(n974), .B(n973), .Z(n978) );
  NAND U2255 ( .A(n976), .B(n975), .Z(n977) );
  NAND U2256 ( .A(n978), .B(n977), .Z(n2141) );
  NAND U2257 ( .A(n980), .B(n979), .Z(n984) );
  NAND U2258 ( .A(n982), .B(n981), .Z(n983) );
  AND U2259 ( .A(n984), .B(n983), .Z(n2142) );
  XNOR U2260 ( .A(n2143), .B(n2142), .Z(n1884) );
  NAND U2261 ( .A(n986), .B(n985), .Z(n990) );
  NAND U2262 ( .A(n988), .B(n987), .Z(n989) );
  NAND U2263 ( .A(n990), .B(n989), .Z(n1883) );
  XOR U2264 ( .A(n1884), .B(n1883), .Z(n1885) );
  XOR U2265 ( .A(n1886), .B(n1885), .Z(n1982) );
  XOR U2266 ( .A(n1983), .B(n1982), .Z(n1984) );
  XOR U2267 ( .A(n1985), .B(n1984), .Z(n1560) );
  NAND U2268 ( .A(n992), .B(n991), .Z(n996) );
  NAND U2269 ( .A(n994), .B(n993), .Z(n995) );
  AND U2270 ( .A(n996), .B(n995), .Z(n2122) );
  NAND U2271 ( .A(n998), .B(n997), .Z(n1002) );
  NAND U2272 ( .A(n1000), .B(n999), .Z(n1001) );
  NAND U2273 ( .A(n1002), .B(n1001), .Z(n2123) );
  NAND U2274 ( .A(n1004), .B(n1003), .Z(n1008) );
  NAND U2275 ( .A(n1006), .B(n1005), .Z(n1007) );
  AND U2276 ( .A(n1008), .B(n1007), .Z(n2124) );
  XNOR U2277 ( .A(n2125), .B(n2124), .Z(n1892) );
  NAND U2278 ( .A(n1010), .B(n1009), .Z(n1014) );
  NAND U2279 ( .A(n1012), .B(n1011), .Z(n1013) );
  AND U2280 ( .A(n1014), .B(n1013), .Z(n1655) );
  NAND U2281 ( .A(n1016), .B(n1015), .Z(n1020) );
  NAND U2282 ( .A(n1018), .B(n1017), .Z(n1019) );
  NAND U2283 ( .A(n1020), .B(n1019), .Z(n1656) );
  NAND U2284 ( .A(n1022), .B(n1021), .Z(n1026) );
  NAND U2285 ( .A(n1024), .B(n1023), .Z(n1025) );
  AND U2286 ( .A(n1026), .B(n1025), .Z(n1657) );
  XNOR U2287 ( .A(n1658), .B(n1657), .Z(n1890) );
  NAND U2288 ( .A(n1028), .B(n1027), .Z(n1032) );
  NAND U2289 ( .A(n1030), .B(n1029), .Z(n1031) );
  AND U2290 ( .A(n1032), .B(n1031), .Z(n1781) );
  NAND U2291 ( .A(n1034), .B(n1033), .Z(n1038) );
  NAND U2292 ( .A(n1036), .B(n1035), .Z(n1037) );
  NAND U2293 ( .A(n1038), .B(n1037), .Z(n1782) );
  NAND U2294 ( .A(n1040), .B(n1039), .Z(n1044) );
  NAND U2295 ( .A(n1042), .B(n1041), .Z(n1043) );
  AND U2296 ( .A(n1044), .B(n1043), .Z(n1783) );
  XNOR U2297 ( .A(n1784), .B(n1783), .Z(n1889) );
  XOR U2298 ( .A(n1890), .B(n1889), .Z(n1891) );
  XOR U2299 ( .A(n1892), .B(n1891), .Z(n1977) );
  NAND U2300 ( .A(n1046), .B(n1045), .Z(n1050) );
  NAND U2301 ( .A(n1048), .B(n1047), .Z(n1049) );
  AND U2302 ( .A(n1050), .B(n1049), .Z(n2116) );
  NAND U2303 ( .A(n1052), .B(n1051), .Z(n1056) );
  NAND U2304 ( .A(n1054), .B(n1053), .Z(n1055) );
  NAND U2305 ( .A(n1056), .B(n1055), .Z(n2117) );
  NAND U2306 ( .A(n1058), .B(n1057), .Z(n1062) );
  NAND U2307 ( .A(n1060), .B(n1059), .Z(n1061) );
  AND U2308 ( .A(n1062), .B(n1061), .Z(n2118) );
  XNOR U2309 ( .A(n2119), .B(n2118), .Z(n1916) );
  NAND U2310 ( .A(n1064), .B(n1063), .Z(n1068) );
  NAND U2311 ( .A(n1066), .B(n1065), .Z(n1067) );
  AND U2312 ( .A(n1068), .B(n1067), .Z(n1739) );
  NAND U2313 ( .A(n1070), .B(n1069), .Z(n1074) );
  NAND U2314 ( .A(n1072), .B(n1071), .Z(n1073) );
  AND U2315 ( .A(n1074), .B(n1073), .Z(n1740) );
  XOR U2316 ( .A(n1739), .B(n1740), .Z(n1742) );
  NAND U2317 ( .A(n1076), .B(n1075), .Z(n1080) );
  NAND U2318 ( .A(n1078), .B(n1077), .Z(n1079) );
  AND U2319 ( .A(n1080), .B(n1079), .Z(n1741) );
  XNOR U2320 ( .A(n1742), .B(n1741), .Z(n1914) );
  NAND U2321 ( .A(n1082), .B(n1081), .Z(n1086) );
  NAND U2322 ( .A(n1084), .B(n1083), .Z(n1085) );
  AND U2323 ( .A(n1086), .B(n1085), .Z(n1643) );
  NAND U2324 ( .A(n1088), .B(n1087), .Z(n1092) );
  NAND U2325 ( .A(n1090), .B(n1089), .Z(n1091) );
  AND U2326 ( .A(n1092), .B(n1091), .Z(n1644) );
  XOR U2327 ( .A(n1643), .B(n1644), .Z(n1646) );
  NAND U2328 ( .A(n1094), .B(n1093), .Z(n1098) );
  NAND U2329 ( .A(n1096), .B(n1095), .Z(n1097) );
  AND U2330 ( .A(n1098), .B(n1097), .Z(n1645) );
  XNOR U2331 ( .A(n1646), .B(n1645), .Z(n1913) );
  XOR U2332 ( .A(n1914), .B(n1913), .Z(n1915) );
  XOR U2333 ( .A(n1916), .B(n1915), .Z(n1976) );
  XOR U2334 ( .A(n1977), .B(n1976), .Z(n1979) );
  NAND U2335 ( .A(n1100), .B(n1099), .Z(n1104) );
  NAND U2336 ( .A(n1102), .B(n1101), .Z(n1103) );
  AND U2337 ( .A(n1104), .B(n1103), .Z(n1709) );
  NAND U2338 ( .A(n1106), .B(n1105), .Z(n1110) );
  NAND U2339 ( .A(n1108), .B(n1107), .Z(n1109) );
  AND U2340 ( .A(n1110), .B(n1109), .Z(n1710) );
  XOR U2341 ( .A(n1709), .B(n1710), .Z(n1712) );
  NAND U2342 ( .A(n1112), .B(n1111), .Z(n1116) );
  NAND U2343 ( .A(n1114), .B(n1113), .Z(n1115) );
  AND U2344 ( .A(n1116), .B(n1115), .Z(n1711) );
  XNOR U2345 ( .A(n1712), .B(n1711), .Z(n1928) );
  NAND U2346 ( .A(n1118), .B(n1117), .Z(n1122) );
  NAND U2347 ( .A(n1120), .B(n1119), .Z(n1121) );
  AND U2348 ( .A(n1122), .B(n1121), .Z(n1649) );
  NANDN U2349 ( .A(n1124), .B(n1123), .Z(n1128) );
  NAND U2350 ( .A(n1126), .B(n1125), .Z(n1127) );
  AND U2351 ( .A(n1128), .B(n1127), .Z(n1650) );
  XOR U2352 ( .A(n1649), .B(n1650), .Z(n1652) );
  NANDN U2353 ( .A(n1130), .B(n1129), .Z(n1134) );
  NAND U2354 ( .A(n1132), .B(n1131), .Z(n1133) );
  AND U2355 ( .A(n1134), .B(n1133), .Z(n1651) );
  XNOR U2356 ( .A(n1652), .B(n1651), .Z(n1926) );
  NAND U2357 ( .A(n1136), .B(n1135), .Z(n1140) );
  NAND U2358 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U2359 ( .A(n1140), .B(n1139), .Z(n2146) );
  NANDN U2360 ( .A(n1142), .B(n1141), .Z(n1146) );
  NAND U2361 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U2362 ( .A(n1146), .B(n1145), .Z(n2147) );
  NAND U2363 ( .A(n1148), .B(n1147), .Z(n1152) );
  NAND U2364 ( .A(n1150), .B(n1149), .Z(n1151) );
  AND U2365 ( .A(n1152), .B(n1151), .Z(n2148) );
  XNOR U2366 ( .A(n2149), .B(n2148), .Z(n1925) );
  XOR U2367 ( .A(n1926), .B(n1925), .Z(n1927) );
  XOR U2368 ( .A(n1928), .B(n1927), .Z(n1978) );
  XNOR U2369 ( .A(n1979), .B(n1978), .Z(n1559) );
  NAND U2370 ( .A(n1154), .B(n1153), .Z(n1158) );
  NAND U2371 ( .A(n1156), .B(n1155), .Z(n1157) );
  AND U2372 ( .A(n1158), .B(n1157), .Z(n1904) );
  NAND U2373 ( .A(n1160), .B(n1159), .Z(n1164) );
  NAND U2374 ( .A(n1162), .B(n1161), .Z(n1163) );
  AND U2375 ( .A(n1164), .B(n1163), .Z(n1902) );
  NAND U2376 ( .A(n1166), .B(n1165), .Z(n1170) );
  NAND U2377 ( .A(n1168), .B(n1167), .Z(n1169) );
  AND U2378 ( .A(n1170), .B(n1169), .Z(n1901) );
  XOR U2379 ( .A(n1904), .B(n1903), .Z(n2259) );
  XNOR U2380 ( .A(n2260), .B(n2259), .Z(n2262) );
  XOR U2381 ( .A(n2261), .B(n2262), .Z(n2257) );
  NAND U2382 ( .A(n1172), .B(n1171), .Z(n1176) );
  NAND U2383 ( .A(n1174), .B(n1173), .Z(n1175) );
  AND U2384 ( .A(n1176), .B(n1175), .Z(n1856) );
  NAND U2385 ( .A(n1178), .B(n1177), .Z(n1182) );
  NAND U2386 ( .A(n1180), .B(n1179), .Z(n1181) );
  NAND U2387 ( .A(n1182), .B(n1181), .Z(n2017) );
  NAND U2388 ( .A(n1184), .B(n1183), .Z(n1188) );
  NAND U2389 ( .A(n1186), .B(n1185), .Z(n1187) );
  NAND U2390 ( .A(n1188), .B(n1187), .Z(n2015) );
  NAND U2391 ( .A(n1190), .B(n1189), .Z(n1194) );
  NAND U2392 ( .A(n1192), .B(n1191), .Z(n1193) );
  AND U2393 ( .A(n1194), .B(n1193), .Z(n1844) );
  NAND U2394 ( .A(n1196), .B(n1195), .Z(n1200) );
  NAND U2395 ( .A(n1198), .B(n1197), .Z(n1199) );
  AND U2396 ( .A(n1200), .B(n1199), .Z(n1841) );
  NAND U2397 ( .A(n1202), .B(n1201), .Z(n1206) );
  NAND U2398 ( .A(n1204), .B(n1203), .Z(n1205) );
  AND U2399 ( .A(n1206), .B(n1205), .Z(n1842) );
  XOR U2400 ( .A(n1841), .B(n1842), .Z(n1843) );
  XNOR U2401 ( .A(n1844), .B(n1843), .Z(n2016) );
  XNOR U2402 ( .A(n2015), .B(n2016), .Z(n1207) );
  XOR U2403 ( .A(n2017), .B(n1207), .Z(n1853) );
  NAND U2404 ( .A(n1209), .B(n1208), .Z(n1213) );
  NAND U2405 ( .A(n1211), .B(n1210), .Z(n1212) );
  AND U2406 ( .A(n1213), .B(n1212), .Z(n1854) );
  XOR U2407 ( .A(n1853), .B(n1854), .Z(n1855) );
  XOR U2408 ( .A(n1856), .B(n1855), .Z(n2265) );
  NAND U2409 ( .A(n1215), .B(n1214), .Z(n1219) );
  NAND U2410 ( .A(n1217), .B(n1216), .Z(n1218) );
  NAND U2411 ( .A(n1219), .B(n1218), .Z(n2022) );
  NAND U2412 ( .A(n1221), .B(n1220), .Z(n1225) );
  NAND U2413 ( .A(n1223), .B(n1222), .Z(n1224) );
  AND U2414 ( .A(n1225), .B(n1224), .Z(n1592) );
  NAND U2415 ( .A(n1227), .B(n1226), .Z(n1231) );
  NAND U2416 ( .A(n1229), .B(n1228), .Z(n1230) );
  AND U2417 ( .A(n1231), .B(n1230), .Z(n1589) );
  NAND U2418 ( .A(n1233), .B(n1232), .Z(n1237) );
  NAND U2419 ( .A(n1235), .B(n1234), .Z(n1236) );
  AND U2420 ( .A(n1237), .B(n1236), .Z(n1590) );
  XOR U2421 ( .A(n1589), .B(n1590), .Z(n1591) );
  XOR U2422 ( .A(n1592), .B(n1591), .Z(n2021) );
  XOR U2423 ( .A(n2022), .B(n2021), .Z(n2024) );
  NAND U2424 ( .A(n1239), .B(n1238), .Z(n1243) );
  NAND U2425 ( .A(n1241), .B(n1240), .Z(n1242) );
  AND U2426 ( .A(n1243), .B(n1242), .Z(n1580) );
  NAND U2427 ( .A(n1245), .B(n1244), .Z(n1249) );
  NAND U2428 ( .A(n1247), .B(n1246), .Z(n1248) );
  AND U2429 ( .A(n1249), .B(n1248), .Z(n1577) );
  NAND U2430 ( .A(n1251), .B(n1250), .Z(n1255) );
  NAND U2431 ( .A(n1253), .B(n1252), .Z(n1254) );
  AND U2432 ( .A(n1255), .B(n1254), .Z(n1578) );
  XOR U2433 ( .A(n1577), .B(n1578), .Z(n1579) );
  XOR U2434 ( .A(n1580), .B(n1579), .Z(n2023) );
  XOR U2435 ( .A(n2024), .B(n2023), .Z(n1790) );
  NAND U2436 ( .A(n1257), .B(n1256), .Z(n1261) );
  NAND U2437 ( .A(n1259), .B(n1258), .Z(n1260) );
  AND U2438 ( .A(n1261), .B(n1260), .Z(n1957) );
  NAND U2439 ( .A(n1263), .B(n1262), .Z(n1267) );
  NAND U2440 ( .A(n1265), .B(n1264), .Z(n1266) );
  AND U2441 ( .A(n1267), .B(n1266), .Z(n1838) );
  NAND U2442 ( .A(n1269), .B(n1268), .Z(n1273) );
  NAND U2443 ( .A(n1271), .B(n1270), .Z(n1272) );
  AND U2444 ( .A(n1273), .B(n1272), .Z(n1835) );
  NAND U2445 ( .A(n1275), .B(n1274), .Z(n1279) );
  NAND U2446 ( .A(n1277), .B(n1276), .Z(n1278) );
  AND U2447 ( .A(n1279), .B(n1278), .Z(n1836) );
  XOR U2448 ( .A(n1835), .B(n1836), .Z(n1837) );
  XNOR U2449 ( .A(n1838), .B(n1837), .Z(n1955) );
  NAND U2450 ( .A(n1281), .B(n1280), .Z(n1285) );
  NAND U2451 ( .A(n1283), .B(n1282), .Z(n1284) );
  AND U2452 ( .A(n1285), .B(n1284), .Z(n1598) );
  NAND U2453 ( .A(n1287), .B(n1286), .Z(n1291) );
  NAND U2454 ( .A(n1289), .B(n1288), .Z(n1290) );
  AND U2455 ( .A(n1291), .B(n1290), .Z(n1595) );
  NAND U2456 ( .A(n1293), .B(n1292), .Z(n1297) );
  NAND U2457 ( .A(n1295), .B(n1294), .Z(n1296) );
  AND U2458 ( .A(n1297), .B(n1296), .Z(n1596) );
  XOR U2459 ( .A(n1595), .B(n1596), .Z(n1597) );
  XOR U2460 ( .A(n1598), .B(n1597), .Z(n1956) );
  XOR U2461 ( .A(n1955), .B(n1956), .Z(n1298) );
  XOR U2462 ( .A(n1957), .B(n1298), .Z(n1787) );
  NAND U2463 ( .A(n1300), .B(n1299), .Z(n1304) );
  NAND U2464 ( .A(n1302), .B(n1301), .Z(n1303) );
  NAND U2465 ( .A(n1304), .B(n1303), .Z(n2203) );
  NAND U2466 ( .A(n1306), .B(n1305), .Z(n1310) );
  NAND U2467 ( .A(n1308), .B(n1307), .Z(n1309) );
  AND U2468 ( .A(n1310), .B(n1309), .Z(n1574) );
  NAND U2469 ( .A(n1312), .B(n1311), .Z(n1316) );
  NAND U2470 ( .A(n1314), .B(n1313), .Z(n1315) );
  AND U2471 ( .A(n1316), .B(n1315), .Z(n1571) );
  NAND U2472 ( .A(n1318), .B(n1317), .Z(n1322) );
  NAND U2473 ( .A(n1320), .B(n1319), .Z(n1321) );
  AND U2474 ( .A(n1322), .B(n1321), .Z(n1572) );
  XOR U2475 ( .A(n1571), .B(n1572), .Z(n1573) );
  XNOR U2476 ( .A(n1574), .B(n1573), .Z(n2201) );
  NAND U2477 ( .A(n1324), .B(n1323), .Z(n1328) );
  NAND U2478 ( .A(n1326), .B(n1325), .Z(n1327) );
  NAND U2479 ( .A(n1328), .B(n1327), .Z(n2200) );
  XOR U2480 ( .A(n2201), .B(n2200), .Z(n2202) );
  XOR U2481 ( .A(n2203), .B(n2202), .Z(n1788) );
  XOR U2482 ( .A(n1787), .B(n1788), .Z(n1789) );
  XNOR U2483 ( .A(n2265), .B(n2266), .Z(n2267) );
  NAND U2484 ( .A(n1330), .B(n1329), .Z(n1334) );
  NAND U2485 ( .A(n1332), .B(n1331), .Z(n1333) );
  AND U2486 ( .A(n1334), .B(n1333), .Z(n1568) );
  NAND U2487 ( .A(n1336), .B(n1335), .Z(n1340) );
  NAND U2488 ( .A(n1338), .B(n1337), .Z(n1339) );
  AND U2489 ( .A(n1340), .B(n1339), .Z(n1769) );
  NAND U2490 ( .A(n1342), .B(n1341), .Z(n1346) );
  NAND U2491 ( .A(n1344), .B(n1343), .Z(n1345) );
  AND U2492 ( .A(n1346), .B(n1345), .Z(n1770) );
  XOR U2493 ( .A(n1769), .B(n1770), .Z(n1772) );
  NAND U2494 ( .A(n1347), .B(oglobal[0]), .Z(n1351) );
  NAND U2495 ( .A(n1349), .B(n1348), .Z(n1350) );
  AND U2496 ( .A(n1351), .B(n1350), .Z(n1771) );
  XOR U2497 ( .A(n1772), .B(n1771), .Z(n1808) );
  NAND U2498 ( .A(n1353), .B(n1352), .Z(n1357) );
  NAND U2499 ( .A(n1355), .B(n1354), .Z(n1356) );
  AND U2500 ( .A(n1357), .B(n1356), .Z(n1775) );
  NAND U2501 ( .A(n1359), .B(n1358), .Z(n1363) );
  NAND U2502 ( .A(n1361), .B(n1360), .Z(n1362) );
  AND U2503 ( .A(n1363), .B(n1362), .Z(n1776) );
  XOR U2504 ( .A(n1775), .B(n1776), .Z(n1778) );
  NAND U2505 ( .A(n1365), .B(n1364), .Z(n1369) );
  NAND U2506 ( .A(n1367), .B(n1366), .Z(n1368) );
  AND U2507 ( .A(n1369), .B(n1368), .Z(n1777) );
  XNOR U2508 ( .A(n1778), .B(n1777), .Z(n1806) );
  NAND U2509 ( .A(n1371), .B(n1370), .Z(n1375) );
  NAND U2510 ( .A(n1373), .B(n1372), .Z(n1374) );
  AND U2511 ( .A(n1375), .B(n1374), .Z(n1805) );
  XOR U2512 ( .A(n1806), .B(n1805), .Z(n1807) );
  XOR U2513 ( .A(n1808), .B(n1807), .Z(n1975) );
  NAND U2514 ( .A(n1377), .B(n1376), .Z(n1381) );
  NAND U2515 ( .A(n1379), .B(n1378), .Z(n1380) );
  AND U2516 ( .A(n1381), .B(n1380), .Z(n1826) );
  NAND U2517 ( .A(n1383), .B(n1382), .Z(n1387) );
  NAND U2518 ( .A(n1385), .B(n1384), .Z(n1386) );
  AND U2519 ( .A(n1387), .B(n1386), .Z(n1823) );
  NAND U2520 ( .A(n1389), .B(n1388), .Z(n1393) );
  NAND U2521 ( .A(n1391), .B(n1390), .Z(n1392) );
  AND U2522 ( .A(n1393), .B(n1392), .Z(n1824) );
  XOR U2523 ( .A(n1823), .B(n1824), .Z(n1825) );
  XNOR U2524 ( .A(n1826), .B(n1825), .Z(n1974) );
  NAND U2525 ( .A(n1395), .B(n1394), .Z(n1399) );
  NANDN U2526 ( .A(n1397), .B(n1396), .Z(n1398) );
  AND U2527 ( .A(n1399), .B(n1398), .Z(n1820) );
  NAND U2528 ( .A(n1401), .B(n1400), .Z(n1405) );
  NAND U2529 ( .A(n1403), .B(n1402), .Z(n1404) );
  AND U2530 ( .A(n1405), .B(n1404), .Z(n2057) );
  NAND U2531 ( .A(n1407), .B(n1406), .Z(n1411) );
  NAND U2532 ( .A(n1409), .B(n1408), .Z(n1410) );
  AND U2533 ( .A(n1411), .B(n1410), .Z(n2058) );
  XOR U2534 ( .A(n2057), .B(n2058), .Z(n2060) );
  NAND U2535 ( .A(n1413), .B(n1412), .Z(n1417) );
  NAND U2536 ( .A(n1415), .B(n1414), .Z(n1416) );
  AND U2537 ( .A(n1417), .B(n1416), .Z(n2059) );
  XNOR U2538 ( .A(n2060), .B(n2059), .Z(n1818) );
  NAND U2539 ( .A(n1419), .B(n1418), .Z(n1423) );
  NAND U2540 ( .A(n1421), .B(n1420), .Z(n1422) );
  AND U2541 ( .A(n1423), .B(n1422), .Z(n1817) );
  XOR U2542 ( .A(n1818), .B(n1817), .Z(n1819) );
  XOR U2543 ( .A(n1820), .B(n1819), .Z(n1973) );
  XOR U2544 ( .A(n1974), .B(n1973), .Z(n1424) );
  XOR U2545 ( .A(n1975), .B(n1424), .Z(n1566) );
  NAND U2546 ( .A(n1426), .B(n1425), .Z(n1430) );
  NAND U2547 ( .A(n1428), .B(n1427), .Z(n1429) );
  AND U2548 ( .A(n1430), .B(n1429), .Z(n1691) );
  NAND U2549 ( .A(n1432), .B(n1431), .Z(n1436) );
  NAND U2550 ( .A(n1434), .B(n1433), .Z(n1435) );
  AND U2551 ( .A(n1436), .B(n1435), .Z(n1692) );
  XOR U2552 ( .A(n1691), .B(n1692), .Z(n1694) );
  NAND U2553 ( .A(n1438), .B(n1437), .Z(n1442) );
  NAND U2554 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U2555 ( .A(n1442), .B(n1441), .Z(n1693) );
  XNOR U2556 ( .A(n1694), .B(n1693), .Z(n1868) );
  NANDN U2557 ( .A(n1444), .B(n1443), .Z(n1448) );
  NAND U2558 ( .A(n1446), .B(n1445), .Z(n1447) );
  AND U2559 ( .A(n1448), .B(n1447), .Z(n1757) );
  NANDN U2560 ( .A(n1450), .B(n1449), .Z(n1454) );
  NAND U2561 ( .A(n1452), .B(n1451), .Z(n1453) );
  AND U2562 ( .A(n1454), .B(n1453), .Z(n1758) );
  XOR U2563 ( .A(n1757), .B(n1758), .Z(n1760) );
  NANDN U2564 ( .A(n1456), .B(n1455), .Z(n1460) );
  NAND U2565 ( .A(n1458), .B(n1457), .Z(n1459) );
  AND U2566 ( .A(n1460), .B(n1459), .Z(n1759) );
  XNOR U2567 ( .A(n1760), .B(n1759), .Z(n1866) );
  NAND U2568 ( .A(n1462), .B(n1461), .Z(n1466) );
  NAND U2569 ( .A(n1464), .B(n1463), .Z(n1465) );
  AND U2570 ( .A(n1466), .B(n1465), .Z(n1865) );
  XOR U2571 ( .A(n1866), .B(n1865), .Z(n1867) );
  XNOR U2572 ( .A(n1868), .B(n1867), .Z(n2002) );
  NAND U2573 ( .A(n1468), .B(n1467), .Z(n1472) );
  NAND U2574 ( .A(n1470), .B(n1469), .Z(n1471) );
  AND U2575 ( .A(n1472), .B(n1471), .Z(n2230) );
  NAND U2576 ( .A(n1474), .B(n1473), .Z(n1478) );
  NAND U2577 ( .A(n1476), .B(n1475), .Z(n1477) );
  AND U2578 ( .A(n1478), .B(n1477), .Z(n2231) );
  XOR U2579 ( .A(n2230), .B(n2231), .Z(n2233) );
  NAND U2580 ( .A(n1480), .B(n1479), .Z(n1484) );
  NAND U2581 ( .A(n1482), .B(n1481), .Z(n1483) );
  AND U2582 ( .A(n1484), .B(n1483), .Z(n2232) );
  XNOR U2583 ( .A(n2233), .B(n2232), .Z(n1874) );
  NAND U2584 ( .A(n1486), .B(n1485), .Z(n1490) );
  NAND U2585 ( .A(n1488), .B(n1487), .Z(n1489) );
  AND U2586 ( .A(n1490), .B(n1489), .Z(n1715) );
  NAND U2587 ( .A(n1492), .B(n1491), .Z(n1496) );
  NAND U2588 ( .A(n1494), .B(n1493), .Z(n1495) );
  AND U2589 ( .A(n1496), .B(n1495), .Z(n1716) );
  XOR U2590 ( .A(n1715), .B(n1716), .Z(n1718) );
  NAND U2591 ( .A(n1498), .B(n1497), .Z(n1502) );
  NAND U2592 ( .A(n1500), .B(n1499), .Z(n1501) );
  AND U2593 ( .A(n1502), .B(n1501), .Z(n1717) );
  XNOR U2594 ( .A(n1718), .B(n1717), .Z(n1872) );
  NAND U2595 ( .A(n1504), .B(n1503), .Z(n1508) );
  NAND U2596 ( .A(n1506), .B(n1505), .Z(n1507) );
  AND U2597 ( .A(n1508), .B(n1507), .Z(n1871) );
  XOR U2598 ( .A(n1872), .B(n1871), .Z(n1873) );
  XNOR U2599 ( .A(n1874), .B(n1873), .Z(n2001) );
  NANDN U2600 ( .A(n1510), .B(n1509), .Z(n1514) );
  NAND U2601 ( .A(n1512), .B(n1511), .Z(n1513) );
  AND U2602 ( .A(n1514), .B(n1513), .Z(n1631) );
  NANDN U2603 ( .A(n1516), .B(n1515), .Z(n1520) );
  NAND U2604 ( .A(n1518), .B(n1517), .Z(n1519) );
  AND U2605 ( .A(n1520), .B(n1519), .Z(n1632) );
  XOR U2606 ( .A(n1631), .B(n1632), .Z(n1634) );
  NANDN U2607 ( .A(n1522), .B(n1521), .Z(n1526) );
  NAND U2608 ( .A(n1524), .B(n1523), .Z(n1525) );
  AND U2609 ( .A(n1526), .B(n1525), .Z(n1633) );
  XOR U2610 ( .A(n1634), .B(n1633), .Z(n1802) );
  NANDN U2611 ( .A(n1528), .B(n1527), .Z(n1532) );
  NAND U2612 ( .A(n1530), .B(n1529), .Z(n1531) );
  AND U2613 ( .A(n1532), .B(n1531), .Z(n1637) );
  NANDN U2614 ( .A(n1534), .B(n1533), .Z(n1538) );
  NAND U2615 ( .A(n1536), .B(n1535), .Z(n1537) );
  AND U2616 ( .A(n1538), .B(n1537), .Z(n1638) );
  XOR U2617 ( .A(n1637), .B(n1638), .Z(n1640) );
  NANDN U2618 ( .A(n1540), .B(n1539), .Z(n1544) );
  NAND U2619 ( .A(n1542), .B(n1541), .Z(n1543) );
  AND U2620 ( .A(n1544), .B(n1543), .Z(n1639) );
  XNOR U2621 ( .A(n1640), .B(n1639), .Z(n1800) );
  NAND U2622 ( .A(n1546), .B(n1545), .Z(n1550) );
  NAND U2623 ( .A(n1548), .B(n1547), .Z(n1549) );
  AND U2624 ( .A(n1550), .B(n1549), .Z(n1799) );
  XOR U2625 ( .A(n1800), .B(n1799), .Z(n1801) );
  XOR U2626 ( .A(n1802), .B(n1801), .Z(n2000) );
  XOR U2627 ( .A(n2001), .B(n2000), .Z(n2003) );
  XOR U2628 ( .A(n2002), .B(n2003), .Z(n1565) );
  XNOR U2629 ( .A(n2267), .B(n2268), .Z(n2256) );
  IV U2630 ( .A(n2256), .Z(n2254) );
  NAND U2631 ( .A(n1552), .B(n1551), .Z(n1556) );
  NAND U2632 ( .A(n1554), .B(n1553), .Z(n1555) );
  AND U2633 ( .A(n1556), .B(n1555), .Z(n2255) );
  XOR U2634 ( .A(n2254), .B(n2255), .Z(n1557) );
  XOR U2635 ( .A(n2257), .B(n1557), .Z(n2277) );
  XOR U2636 ( .A(n2278), .B(n2277), .Z(n1558) );
  XNOR U2637 ( .A(n2279), .B(n1558), .Z(o[1]) );
  NANDN U2638 ( .A(n1560), .B(n1559), .Z(n1564) );
  NANDN U2639 ( .A(n1562), .B(n1561), .Z(n1563) );
  AND U2640 ( .A(n1564), .B(n1563), .Z(n2528) );
  NANDN U2641 ( .A(n1566), .B(n1565), .Z(n1570) );
  NANDN U2642 ( .A(n1568), .B(n1567), .Z(n1569) );
  NAND U2643 ( .A(n1570), .B(n1569), .Z(n2529) );
  NAND U2644 ( .A(n1572), .B(n1571), .Z(n1576) );
  NAND U2645 ( .A(n1574), .B(n1573), .Z(n1575) );
  AND U2646 ( .A(n1576), .B(n1575), .Z(n2326) );
  NAND U2647 ( .A(n1578), .B(n1577), .Z(n1582) );
  NAND U2648 ( .A(n1580), .B(n1579), .Z(n1581) );
  AND U2649 ( .A(n1582), .B(n1581), .Z(n2324) );
  NAND U2650 ( .A(n1584), .B(n1583), .Z(n1588) );
  NAND U2651 ( .A(n1586), .B(n1585), .Z(n1587) );
  NAND U2652 ( .A(n1588), .B(n1587), .Z(n2323) );
  NAND U2653 ( .A(n1590), .B(n1589), .Z(n1594) );
  NAND U2654 ( .A(n1592), .B(n1591), .Z(n1593) );
  NAND U2655 ( .A(n1594), .B(n1593), .Z(n2631) );
  NAND U2656 ( .A(n1596), .B(n1595), .Z(n1600) );
  NAND U2657 ( .A(n1598), .B(n1597), .Z(n1599) );
  NAND U2658 ( .A(n1600), .B(n1599), .Z(n2629) );
  NAND U2659 ( .A(n1602), .B(n1601), .Z(n1606) );
  NAND U2660 ( .A(n1604), .B(n1603), .Z(n1605) );
  NAND U2661 ( .A(n1606), .B(n1605), .Z(n2628) );
  XOR U2662 ( .A(n2629), .B(n2628), .Z(n2630) );
  XOR U2663 ( .A(n2631), .B(n2630), .Z(n2287) );
  XOR U2664 ( .A(n2288), .B(n2287), .Z(n2290) );
  NANDN U2665 ( .A(n1608), .B(n1607), .Z(n1612) );
  NAND U2666 ( .A(n1610), .B(n1609), .Z(n1611) );
  AND U2667 ( .A(n1612), .B(n1611), .Z(n2398) );
  NANDN U2668 ( .A(n1614), .B(n1613), .Z(n1618) );
  NAND U2669 ( .A(n1616), .B(n1615), .Z(n1617) );
  AND U2670 ( .A(n1618), .B(n1617), .Z(n2396) );
  NAND U2671 ( .A(n1620), .B(n1619), .Z(n1624) );
  NAND U2672 ( .A(n1622), .B(n1621), .Z(n1623) );
  NAND U2673 ( .A(n1624), .B(n1623), .Z(n2395) );
  NAND U2674 ( .A(n1626), .B(n1625), .Z(n1630) );
  NAND U2675 ( .A(n1628), .B(n1627), .Z(n1629) );
  NAND U2676 ( .A(n1630), .B(n1629), .Z(n2641) );
  NAND U2677 ( .A(n1632), .B(n1631), .Z(n1636) );
  NAND U2678 ( .A(n1634), .B(n1633), .Z(n1635) );
  AND U2679 ( .A(n1636), .B(n1635), .Z(n2459) );
  NAND U2680 ( .A(n1638), .B(n1637), .Z(n1642) );
  NAND U2681 ( .A(n1640), .B(n1639), .Z(n1641) );
  AND U2682 ( .A(n1642), .B(n1641), .Z(n2457) );
  NAND U2683 ( .A(n1644), .B(n1643), .Z(n1648) );
  NAND U2684 ( .A(n1646), .B(n1645), .Z(n1647) );
  NAND U2685 ( .A(n1648), .B(n1647), .Z(n2456) );
  XOR U2686 ( .A(n2459), .B(n2458), .Z(n2640) );
  XOR U2687 ( .A(n2641), .B(n2640), .Z(n2643) );
  XOR U2688 ( .A(n2642), .B(n2643), .Z(n2289) );
  XOR U2689 ( .A(n2290), .B(n2289), .Z(n2355) );
  NAND U2690 ( .A(n1650), .B(n1649), .Z(n1654) );
  NAND U2691 ( .A(n1652), .B(n1651), .Z(n1653) );
  AND U2692 ( .A(n1654), .B(n1653), .Z(n2445) );
  NANDN U2693 ( .A(n1656), .B(n1655), .Z(n1660) );
  NAND U2694 ( .A(n1658), .B(n1657), .Z(n1659) );
  NAND U2695 ( .A(n1660), .B(n1659), .Z(n2444) );
  NAND U2696 ( .A(n1662), .B(n1661), .Z(n1666) );
  NAND U2697 ( .A(n1664), .B(n1663), .Z(n1665) );
  AND U2698 ( .A(n1666), .B(n1665), .Z(n2483) );
  NANDN U2699 ( .A(n1668), .B(n1667), .Z(n1672) );
  NAND U2700 ( .A(n1670), .B(n1669), .Z(n1671) );
  AND U2701 ( .A(n1672), .B(n1671), .Z(n2481) );
  NANDN U2702 ( .A(n1674), .B(n1673), .Z(n1678) );
  NAND U2703 ( .A(n1676), .B(n1675), .Z(n1677) );
  NAND U2704 ( .A(n1678), .B(n1677), .Z(n2480) );
  XNOR U2705 ( .A(n2447), .B(n2446), .Z(n2577) );
  NAND U2706 ( .A(n1680), .B(n1679), .Z(n1684) );
  NAND U2707 ( .A(n1682), .B(n1681), .Z(n1683) );
  AND U2708 ( .A(n1684), .B(n1683), .Z(n2413) );
  XOR U2709 ( .A(n2413), .B(oglobal[2]), .Z(n2404) );
  NAND U2710 ( .A(n1686), .B(n1685), .Z(n1690) );
  NAND U2711 ( .A(n1688), .B(n1687), .Z(n1689) );
  AND U2712 ( .A(n1690), .B(n1689), .Z(n2402) );
  NAND U2713 ( .A(n1692), .B(n1691), .Z(n1696) );
  NAND U2714 ( .A(n1694), .B(n1693), .Z(n1695) );
  NAND U2715 ( .A(n1696), .B(n1695), .Z(n2401) );
  NAND U2716 ( .A(n1698), .B(n1697), .Z(n1702) );
  NAND U2717 ( .A(n1700), .B(n1699), .Z(n1701) );
  NAND U2718 ( .A(n1702), .B(n1701), .Z(n2574) );
  XOR U2719 ( .A(n2575), .B(n2574), .Z(n2576) );
  XNOR U2720 ( .A(n2577), .B(n2576), .Z(n2283) );
  NAND U2721 ( .A(n1704), .B(n1703), .Z(n1708) );
  NAND U2722 ( .A(n1706), .B(n1705), .Z(n1707) );
  NAND U2723 ( .A(n1708), .B(n1707), .Z(n2595) );
  NAND U2724 ( .A(n1710), .B(n1709), .Z(n1714) );
  NAND U2725 ( .A(n1712), .B(n1711), .Z(n1713) );
  NAND U2726 ( .A(n1714), .B(n1713), .Z(n2593) );
  NAND U2727 ( .A(n1716), .B(n1715), .Z(n1720) );
  NAND U2728 ( .A(n1718), .B(n1717), .Z(n1719) );
  NAND U2729 ( .A(n1720), .B(n1719), .Z(n2592) );
  XOR U2730 ( .A(n2593), .B(n2592), .Z(n2594) );
  XNOR U2731 ( .A(n2595), .B(n2594), .Z(n2331) );
  NAND U2732 ( .A(n1722), .B(n1721), .Z(n1726) );
  NAND U2733 ( .A(n1724), .B(n1723), .Z(n1725) );
  AND U2734 ( .A(n1726), .B(n1725), .Z(n2330) );
  NAND U2735 ( .A(n1728), .B(n1727), .Z(n1732) );
  NAND U2736 ( .A(n1730), .B(n1729), .Z(n1731) );
  AND U2737 ( .A(n1732), .B(n1731), .Z(n2607) );
  NANDN U2738 ( .A(n1734), .B(n1733), .Z(n1738) );
  NAND U2739 ( .A(n1736), .B(n1735), .Z(n1737) );
  NAND U2740 ( .A(n1738), .B(n1737), .Z(n2605) );
  NAND U2741 ( .A(n1740), .B(n1739), .Z(n1744) );
  NAND U2742 ( .A(n1742), .B(n1741), .Z(n1743) );
  NAND U2743 ( .A(n1744), .B(n1743), .Z(n2604) );
  XOR U2744 ( .A(n2605), .B(n2604), .Z(n2606) );
  XOR U2745 ( .A(n2607), .B(n2606), .Z(n2329) );
  XNOR U2746 ( .A(n2331), .B(n2332), .Z(n2282) );
  NANDN U2747 ( .A(n1746), .B(n1745), .Z(n1750) );
  NAND U2748 ( .A(n1748), .B(n1747), .Z(n1749) );
  AND U2749 ( .A(n1750), .B(n1749), .Z(n2477) );
  NAND U2750 ( .A(n1752), .B(n1751), .Z(n1756) );
  NAND U2751 ( .A(n1754), .B(n1753), .Z(n1755) );
  AND U2752 ( .A(n1756), .B(n1755), .Z(n2475) );
  NAND U2753 ( .A(n1758), .B(n1757), .Z(n1762) );
  NAND U2754 ( .A(n1760), .B(n1759), .Z(n1761) );
  NAND U2755 ( .A(n1762), .B(n1761), .Z(n2474) );
  NAND U2756 ( .A(n1764), .B(n1763), .Z(n1768) );
  NAND U2757 ( .A(n1766), .B(n1765), .Z(n1767) );
  NAND U2758 ( .A(n1768), .B(n1767), .Z(n2635) );
  NAND U2759 ( .A(n1770), .B(n1769), .Z(n1774) );
  NAND U2760 ( .A(n1772), .B(n1771), .Z(n1773) );
  AND U2761 ( .A(n1774), .B(n1773), .Z(n2613) );
  NAND U2762 ( .A(n1776), .B(n1775), .Z(n1780) );
  NAND U2763 ( .A(n1778), .B(n1777), .Z(n1779) );
  NAND U2764 ( .A(n1780), .B(n1779), .Z(n2611) );
  NANDN U2765 ( .A(n1782), .B(n1781), .Z(n1786) );
  NAND U2766 ( .A(n1784), .B(n1783), .Z(n1785) );
  NAND U2767 ( .A(n1786), .B(n1785), .Z(n2610) );
  XOR U2768 ( .A(n2611), .B(n2610), .Z(n2612) );
  XOR U2769 ( .A(n2613), .B(n2612), .Z(n2634) );
  XOR U2770 ( .A(n2635), .B(n2634), .Z(n2637) );
  XNOR U2771 ( .A(n2636), .B(n2637), .Z(n2281) );
  XOR U2772 ( .A(n2282), .B(n2281), .Z(n2284) );
  XOR U2773 ( .A(n2283), .B(n2284), .Z(n2354) );
  NAND U2774 ( .A(n1788), .B(n1787), .Z(n1792) );
  NANDN U2775 ( .A(n1790), .B(n1789), .Z(n1791) );
  AND U2776 ( .A(n1792), .B(n1791), .Z(n2353) );
  XNOR U2777 ( .A(n2355), .B(n2356), .Z(n2530) );
  XOR U2778 ( .A(n2531), .B(n2530), .Z(n2559) );
  NAND U2779 ( .A(n1794), .B(n1793), .Z(n1798) );
  NAND U2780 ( .A(n1796), .B(n1795), .Z(n1797) );
  NAND U2781 ( .A(n1798), .B(n1797), .Z(n2563) );
  NAND U2782 ( .A(n1800), .B(n1799), .Z(n1804) );
  NANDN U2783 ( .A(n1802), .B(n1801), .Z(n1803) );
  NAND U2784 ( .A(n1804), .B(n1803), .Z(n2435) );
  NAND U2785 ( .A(n1806), .B(n1805), .Z(n1810) );
  NANDN U2786 ( .A(n1808), .B(n1807), .Z(n1809) );
  NAND U2787 ( .A(n1810), .B(n1809), .Z(n2433) );
  NAND U2788 ( .A(n1812), .B(n1811), .Z(n1816) );
  NAND U2789 ( .A(n1814), .B(n1813), .Z(n1815) );
  NAND U2790 ( .A(n1816), .B(n1815), .Z(n2432) );
  XOR U2791 ( .A(n2433), .B(n2432), .Z(n2434) );
  XOR U2792 ( .A(n2435), .B(n2434), .Z(n2487) );
  NAND U2793 ( .A(n1818), .B(n1817), .Z(n1822) );
  NAND U2794 ( .A(n1820), .B(n1819), .Z(n1821) );
  AND U2795 ( .A(n1822), .B(n1821), .Z(n2417) );
  NAND U2796 ( .A(n1824), .B(n1823), .Z(n1828) );
  NAND U2797 ( .A(n1826), .B(n1825), .Z(n1827) );
  AND U2798 ( .A(n1828), .B(n1827), .Z(n2415) );
  NAND U2799 ( .A(n1830), .B(n1829), .Z(n1834) );
  NAND U2800 ( .A(n1832), .B(n1831), .Z(n1833) );
  NAND U2801 ( .A(n1834), .B(n1833), .Z(n2414) );
  XOR U2802 ( .A(n2487), .B(n2486), .Z(n2489) );
  NAND U2803 ( .A(n1836), .B(n1835), .Z(n1840) );
  NAND U2804 ( .A(n1838), .B(n1837), .Z(n1839) );
  AND U2805 ( .A(n1840), .B(n1839), .Z(n2338) );
  NAND U2806 ( .A(n1842), .B(n1841), .Z(n1846) );
  NAND U2807 ( .A(n1844), .B(n1843), .Z(n1845) );
  AND U2808 ( .A(n1846), .B(n1845), .Z(n2336) );
  NAND U2809 ( .A(n1848), .B(n1847), .Z(n1852) );
  NAND U2810 ( .A(n1850), .B(n1849), .Z(n1851) );
  NAND U2811 ( .A(n1852), .B(n1851), .Z(n2335) );
  XOR U2812 ( .A(n2489), .B(n2488), .Z(n2562) );
  XOR U2813 ( .A(n2563), .B(n2562), .Z(n2564) );
  NAND U2814 ( .A(n1854), .B(n1853), .Z(n1858) );
  NAND U2815 ( .A(n1856), .B(n1855), .Z(n1857) );
  AND U2816 ( .A(n1858), .B(n1857), .Z(n2565) );
  XOR U2817 ( .A(n2564), .B(n2565), .Z(n2556) );
  NAND U2818 ( .A(n1860), .B(n1859), .Z(n1864) );
  NAND U2819 ( .A(n1862), .B(n1861), .Z(n1863) );
  NAND U2820 ( .A(n1864), .B(n1863), .Z(n2320) );
  NAND U2821 ( .A(n1866), .B(n1865), .Z(n1870) );
  NAND U2822 ( .A(n1868), .B(n1867), .Z(n1869) );
  NAND U2823 ( .A(n1870), .B(n1869), .Z(n2308) );
  NAND U2824 ( .A(n1872), .B(n1871), .Z(n1876) );
  NAND U2825 ( .A(n1874), .B(n1873), .Z(n1875) );
  NAND U2826 ( .A(n1876), .B(n1875), .Z(n2306) );
  NAND U2827 ( .A(n1878), .B(n1877), .Z(n1882) );
  NANDN U2828 ( .A(n1880), .B(n1879), .Z(n1881) );
  NAND U2829 ( .A(n1882), .B(n1881), .Z(n2305) );
  XOR U2830 ( .A(n2306), .B(n2305), .Z(n2307) );
  XNOR U2831 ( .A(n2308), .B(n2307), .Z(n2318) );
  NAND U2832 ( .A(n1884), .B(n1883), .Z(n1888) );
  NAND U2833 ( .A(n1886), .B(n1885), .Z(n1887) );
  AND U2834 ( .A(n1888), .B(n1887), .Z(n2601) );
  NAND U2835 ( .A(n1890), .B(n1889), .Z(n1894) );
  NAND U2836 ( .A(n1892), .B(n1891), .Z(n1893) );
  NAND U2837 ( .A(n1894), .B(n1893), .Z(n2599) );
  NAND U2838 ( .A(n1896), .B(n1895), .Z(n1900) );
  NAND U2839 ( .A(n1898), .B(n1897), .Z(n1899) );
  NAND U2840 ( .A(n1900), .B(n1899), .Z(n2598) );
  XOR U2841 ( .A(n2599), .B(n2598), .Z(n2600) );
  XOR U2842 ( .A(n2601), .B(n2600), .Z(n2317) );
  XOR U2843 ( .A(n2318), .B(n2317), .Z(n2319) );
  XNOR U2844 ( .A(n2320), .B(n2319), .Z(n2349) );
  NANDN U2845 ( .A(n1902), .B(n1901), .Z(n1906) );
  NAND U2846 ( .A(n1904), .B(n1903), .Z(n1905) );
  AND U2847 ( .A(n1906), .B(n1905), .Z(n2348) );
  NANDN U2848 ( .A(n1908), .B(n1907), .Z(n1912) );
  NANDN U2849 ( .A(n1910), .B(n1909), .Z(n1911) );
  NAND U2850 ( .A(n1912), .B(n1911), .Z(n2366) );
  NAND U2851 ( .A(n1914), .B(n1913), .Z(n1918) );
  NAND U2852 ( .A(n1916), .B(n1915), .Z(n1917) );
  NAND U2853 ( .A(n1918), .B(n1917), .Z(n2302) );
  NAND U2854 ( .A(n1920), .B(n1919), .Z(n1924) );
  NAND U2855 ( .A(n1922), .B(n1921), .Z(n1923) );
  NAND U2856 ( .A(n1924), .B(n1923), .Z(n2300) );
  NAND U2857 ( .A(n1926), .B(n1925), .Z(n1930) );
  NAND U2858 ( .A(n1928), .B(n1927), .Z(n1929) );
  NAND U2859 ( .A(n1930), .B(n1929), .Z(n2299) );
  XOR U2860 ( .A(n2300), .B(n2299), .Z(n2301) );
  XOR U2861 ( .A(n2302), .B(n2301), .Z(n2365) );
  XOR U2862 ( .A(n2366), .B(n2365), .Z(n2368) );
  NAND U2863 ( .A(n1932), .B(n1931), .Z(n1936) );
  NAND U2864 ( .A(n1934), .B(n1933), .Z(n1935) );
  NAND U2865 ( .A(n1936), .B(n1935), .Z(n2625) );
  NAND U2866 ( .A(n1938), .B(n1937), .Z(n1942) );
  NAND U2867 ( .A(n1940), .B(n1939), .Z(n1941) );
  NAND U2868 ( .A(n1942), .B(n1941), .Z(n2623) );
  NAND U2869 ( .A(n1944), .B(n1943), .Z(n1948) );
  NAND U2870 ( .A(n1946), .B(n1945), .Z(n1947) );
  NAND U2871 ( .A(n1948), .B(n1947), .Z(n2622) );
  XOR U2872 ( .A(n2623), .B(n2622), .Z(n2624) );
  XOR U2873 ( .A(n2625), .B(n2624), .Z(n2367) );
  XOR U2874 ( .A(n2368), .B(n2367), .Z(n2347) );
  XNOR U2875 ( .A(n2349), .B(n2350), .Z(n2557) );
  XNOR U2876 ( .A(n2559), .B(n2558), .Z(n2543) );
  XNOR U2877 ( .A(n2493), .B(n2492), .Z(n2495) );
  NAND U2878 ( .A(n1959), .B(n1958), .Z(n1963) );
  NAND U2879 ( .A(n1961), .B(n1960), .Z(n1962) );
  AND U2880 ( .A(n1963), .B(n1962), .Z(n2494) );
  XNOR U2881 ( .A(n2495), .B(n2494), .Z(n2341) );
  XNOR U2882 ( .A(n2342), .B(n2341), .Z(n2344) );
  NAND U2883 ( .A(n1965), .B(n1964), .Z(n1969) );
  NAND U2884 ( .A(n1967), .B(n1966), .Z(n1968) );
  AND U2885 ( .A(n1969), .B(n1968), .Z(n2501) );
  XOR U2886 ( .A(n2499), .B(n2498), .Z(n2500) );
  XNOR U2887 ( .A(n2501), .B(n2500), .Z(n2314) );
  NAND U2888 ( .A(n1977), .B(n1976), .Z(n1981) );
  NAND U2889 ( .A(n1979), .B(n1978), .Z(n1980) );
  AND U2890 ( .A(n1981), .B(n1980), .Z(n2311) );
  NAND U2891 ( .A(n1983), .B(n1982), .Z(n1987) );
  NAND U2892 ( .A(n1985), .B(n1984), .Z(n1986) );
  AND U2893 ( .A(n1987), .B(n1986), .Z(n2312) );
  XOR U2894 ( .A(n2311), .B(n2312), .Z(n2313) );
  XOR U2895 ( .A(n2314), .B(n2313), .Z(n2343) );
  XOR U2896 ( .A(n2344), .B(n2343), .Z(n2535) );
  NAND U2897 ( .A(n1989), .B(n1988), .Z(n1993) );
  NAND U2898 ( .A(n1991), .B(n1990), .Z(n1992) );
  NAND U2899 ( .A(n1993), .B(n1992), .Z(n2439) );
  NAND U2900 ( .A(n1995), .B(n1994), .Z(n1999) );
  NAND U2901 ( .A(n1997), .B(n1996), .Z(n1998) );
  AND U2902 ( .A(n1999), .B(n1998), .Z(n2438) );
  XOR U2903 ( .A(n2439), .B(n2438), .Z(n2441) );
  NAND U2904 ( .A(n2001), .B(n2000), .Z(n2005) );
  NAND U2905 ( .A(n2003), .B(n2002), .Z(n2004) );
  AND U2906 ( .A(n2005), .B(n2004), .Z(n2440) );
  XNOR U2907 ( .A(n2441), .B(n2440), .Z(n2362) );
  NAND U2908 ( .A(n2010), .B(n2009), .Z(n2014) );
  NAND U2909 ( .A(n2012), .B(n2011), .Z(n2013) );
  NAND U2910 ( .A(n2014), .B(n2013), .Z(n2512) );
  XOR U2911 ( .A(n2511), .B(n2510), .Z(n2513) );
  XOR U2912 ( .A(n2512), .B(n2513), .Z(n2359) );
  XNOR U2913 ( .A(n2360), .B(n2359), .Z(n2361) );
  XOR U2914 ( .A(n2362), .B(n2361), .Z(n2534) );
  XOR U2915 ( .A(n2535), .B(n2534), .Z(n2537) );
  NAND U2916 ( .A(n2022), .B(n2021), .Z(n2026) );
  NAND U2917 ( .A(n2024), .B(n2023), .Z(n2025) );
  NAND U2918 ( .A(n2026), .B(n2025), .Z(n2505) );
  NAND U2919 ( .A(n2028), .B(n2027), .Z(n2032) );
  NAND U2920 ( .A(n2030), .B(n2029), .Z(n2031) );
  NAND U2921 ( .A(n2032), .B(n2031), .Z(n2619) );
  NAND U2922 ( .A(n2034), .B(n2033), .Z(n2038) );
  NAND U2923 ( .A(n2036), .B(n2035), .Z(n2037) );
  NAND U2924 ( .A(n2038), .B(n2037), .Z(n2617) );
  NANDN U2925 ( .A(n2040), .B(n2039), .Z(n2044) );
  NAND U2926 ( .A(n2042), .B(n2041), .Z(n2043) );
  NAND U2927 ( .A(n2044), .B(n2043), .Z(n2616) );
  XOR U2928 ( .A(n2617), .B(n2616), .Z(n2618) );
  XNOR U2929 ( .A(n2619), .B(n2618), .Z(n2570) );
  NAND U2930 ( .A(n2046), .B(n2045), .Z(n2050) );
  NAND U2931 ( .A(n2048), .B(n2047), .Z(n2049) );
  NAND U2932 ( .A(n2050), .B(n2049), .Z(n2569) );
  NAND U2933 ( .A(n2052), .B(n2051), .Z(n2056) );
  NAND U2934 ( .A(n2054), .B(n2053), .Z(n2055) );
  AND U2935 ( .A(n2056), .B(n2055), .Z(n2453) );
  NAND U2936 ( .A(n2058), .B(n2057), .Z(n2062) );
  NAND U2937 ( .A(n2060), .B(n2059), .Z(n2061) );
  AND U2938 ( .A(n2062), .B(n2061), .Z(n2451) );
  NANDN U2939 ( .A(n2063), .B(oglobal[1]), .Z(n2067) );
  NANDN U2940 ( .A(n2065), .B(n2064), .Z(n2066) );
  AND U2941 ( .A(n2067), .B(n2066), .Z(n2450) );
  XOR U2942 ( .A(n2453), .B(n2452), .Z(n2568) );
  XOR U2943 ( .A(n2569), .B(n2568), .Z(n2571) );
  XOR U2944 ( .A(n2570), .B(n2571), .Z(n2504) );
  XOR U2945 ( .A(n2505), .B(n2504), .Z(n2507) );
  NAND U2946 ( .A(n2069), .B(n2068), .Z(n2073) );
  NAND U2947 ( .A(n2071), .B(n2070), .Z(n2072) );
  NAND U2948 ( .A(n2073), .B(n2072), .Z(n2589) );
  NANDN U2949 ( .A(n2075), .B(n2074), .Z(n2079) );
  NAND U2950 ( .A(n2077), .B(n2076), .Z(n2078) );
  NAND U2951 ( .A(n2079), .B(n2078), .Z(n2587) );
  NAND U2952 ( .A(n2081), .B(n2080), .Z(n2085) );
  NAND U2953 ( .A(n2083), .B(n2082), .Z(n2084) );
  NAND U2954 ( .A(n2085), .B(n2084), .Z(n2586) );
  XOR U2955 ( .A(n2587), .B(n2586), .Z(n2588) );
  XNOR U2956 ( .A(n2589), .B(n2588), .Z(n2428) );
  NAND U2957 ( .A(n2087), .B(n2086), .Z(n2091) );
  NAND U2958 ( .A(n2089), .B(n2088), .Z(n2090) );
  NAND U2959 ( .A(n2091), .B(n2090), .Z(n2427) );
  NAND U2960 ( .A(n2093), .B(n2092), .Z(n2097) );
  NAND U2961 ( .A(n2095), .B(n2094), .Z(n2096) );
  AND U2962 ( .A(n2097), .B(n2096), .Z(n2380) );
  NAND U2963 ( .A(n2099), .B(n2098), .Z(n2103) );
  NAND U2964 ( .A(n2101), .B(n2100), .Z(n2102) );
  AND U2965 ( .A(n2103), .B(n2102), .Z(n2378) );
  NAND U2966 ( .A(n2105), .B(n2104), .Z(n2109) );
  NAND U2967 ( .A(n2107), .B(n2106), .Z(n2108) );
  NAND U2968 ( .A(n2109), .B(n2108), .Z(n2377) );
  XOR U2969 ( .A(n2380), .B(n2379), .Z(n2426) );
  XOR U2970 ( .A(n2427), .B(n2426), .Z(n2429) );
  XOR U2971 ( .A(n2428), .B(n2429), .Z(n2506) );
  XNOR U2972 ( .A(n2507), .B(n2506), .Z(n2649) );
  NAND U2973 ( .A(n2111), .B(n2110), .Z(n2115) );
  NAND U2974 ( .A(n2113), .B(n2112), .Z(n2114) );
  AND U2975 ( .A(n2115), .B(n2114), .Z(n2517) );
  NANDN U2976 ( .A(n2117), .B(n2116), .Z(n2121) );
  NAND U2977 ( .A(n2119), .B(n2118), .Z(n2120) );
  AND U2978 ( .A(n2121), .B(n2120), .Z(n2392) );
  NANDN U2979 ( .A(n2123), .B(n2122), .Z(n2127) );
  NAND U2980 ( .A(n2125), .B(n2124), .Z(n2126) );
  AND U2981 ( .A(n2127), .B(n2126), .Z(n2390) );
  NANDN U2982 ( .A(n2129), .B(n2128), .Z(n2133) );
  NAND U2983 ( .A(n2131), .B(n2130), .Z(n2132) );
  NAND U2984 ( .A(n2133), .B(n2132), .Z(n2389) );
  NAND U2985 ( .A(n2135), .B(n2134), .Z(n2139) );
  NAND U2986 ( .A(n2137), .B(n2136), .Z(n2138) );
  NAND U2987 ( .A(n2139), .B(n2138), .Z(n2421) );
  NANDN U2988 ( .A(n2141), .B(n2140), .Z(n2145) );
  NAND U2989 ( .A(n2143), .B(n2142), .Z(n2144) );
  AND U2990 ( .A(n2145), .B(n2144), .Z(n2374) );
  NANDN U2991 ( .A(n2147), .B(n2146), .Z(n2151) );
  NAND U2992 ( .A(n2149), .B(n2148), .Z(n2150) );
  AND U2993 ( .A(n2151), .B(n2150), .Z(n2371) );
  NAND U2994 ( .A(n2153), .B(n2152), .Z(n2157) );
  NAND U2995 ( .A(n2155), .B(n2154), .Z(n2156) );
  NAND U2996 ( .A(n2157), .B(n2156), .Z(n2372) );
  XOR U2997 ( .A(n2374), .B(n2373), .Z(n2420) );
  XOR U2998 ( .A(n2421), .B(n2420), .Z(n2423) );
  XOR U2999 ( .A(n2422), .B(n2423), .Z(n2516) );
  XOR U3000 ( .A(n2517), .B(n2516), .Z(n2519) );
  NANDN U3001 ( .A(n2159), .B(n2158), .Z(n2163) );
  NAND U3002 ( .A(n2161), .B(n2160), .Z(n2162) );
  AND U3003 ( .A(n2163), .B(n2162), .Z(n2471) );
  NANDN U3004 ( .A(n2165), .B(n2164), .Z(n2169) );
  NAND U3005 ( .A(n2167), .B(n2166), .Z(n2168) );
  AND U3006 ( .A(n2169), .B(n2168), .Z(n2469) );
  NANDN U3007 ( .A(n2171), .B(n2170), .Z(n2175) );
  NAND U3008 ( .A(n2173), .B(n2172), .Z(n2174) );
  NAND U3009 ( .A(n2175), .B(n2174), .Z(n2468) );
  NAND U3010 ( .A(n2177), .B(n2176), .Z(n2181) );
  NAND U3011 ( .A(n2179), .B(n2178), .Z(n2180) );
  NAND U3012 ( .A(n2181), .B(n2180), .Z(n2463) );
  NANDN U3013 ( .A(n2183), .B(n2182), .Z(n2187) );
  NAND U3014 ( .A(n2185), .B(n2184), .Z(n2186) );
  AND U3015 ( .A(n2187), .B(n2186), .Z(n2386) );
  NANDN U3016 ( .A(n2189), .B(n2188), .Z(n2193) );
  NAND U3017 ( .A(n2191), .B(n2190), .Z(n2192) );
  AND U3018 ( .A(n2193), .B(n2192), .Z(n2384) );
  NANDN U3019 ( .A(n2195), .B(n2194), .Z(n2199) );
  NAND U3020 ( .A(n2197), .B(n2196), .Z(n2198) );
  NAND U3021 ( .A(n2199), .B(n2198), .Z(n2383) );
  XOR U3022 ( .A(n2386), .B(n2385), .Z(n2462) );
  XOR U3023 ( .A(n2463), .B(n2462), .Z(n2465) );
  XOR U3024 ( .A(n2464), .B(n2465), .Z(n2518) );
  XNOR U3025 ( .A(n2519), .B(n2518), .Z(n2647) );
  NAND U3026 ( .A(n2201), .B(n2200), .Z(n2205) );
  NAND U3027 ( .A(n2203), .B(n2202), .Z(n2204) );
  AND U3028 ( .A(n2205), .B(n2204), .Z(n2523) );
  NAND U3029 ( .A(n2207), .B(n2206), .Z(n2211) );
  NAND U3030 ( .A(n2209), .B(n2208), .Z(n2210) );
  NAND U3031 ( .A(n2211), .B(n2210), .Z(n2583) );
  NANDN U3032 ( .A(n2213), .B(n2212), .Z(n2217) );
  NAND U3033 ( .A(n2215), .B(n2214), .Z(n2216) );
  NAND U3034 ( .A(n2217), .B(n2216), .Z(n2581) );
  NAND U3035 ( .A(n2219), .B(n2218), .Z(n2223) );
  NAND U3036 ( .A(n2221), .B(n2220), .Z(n2222) );
  NAND U3037 ( .A(n2223), .B(n2222), .Z(n2580) );
  XOR U3038 ( .A(n2581), .B(n2580), .Z(n2582) );
  XNOR U3039 ( .A(n2583), .B(n2582), .Z(n2295) );
  NAND U3040 ( .A(n2225), .B(n2224), .Z(n2229) );
  NAND U3041 ( .A(n2227), .B(n2226), .Z(n2228) );
  NAND U3042 ( .A(n2229), .B(n2228), .Z(n2294) );
  NAND U3043 ( .A(n2231), .B(n2230), .Z(n2235) );
  NAND U3044 ( .A(n2233), .B(n2232), .Z(n2234) );
  AND U3045 ( .A(n2235), .B(n2234), .Z(n2410) );
  NAND U3046 ( .A(n2237), .B(n2236), .Z(n2241) );
  NAND U3047 ( .A(n2239), .B(n2238), .Z(n2240) );
  AND U3048 ( .A(n2241), .B(n2240), .Z(n2408) );
  NAND U3049 ( .A(n2243), .B(n2242), .Z(n2247) );
  NAND U3050 ( .A(n2245), .B(n2244), .Z(n2246) );
  NAND U3051 ( .A(n2247), .B(n2246), .Z(n2407) );
  XOR U3052 ( .A(n2410), .B(n2409), .Z(n2293) );
  XOR U3053 ( .A(n2294), .B(n2293), .Z(n2296) );
  XOR U3054 ( .A(n2295), .B(n2296), .Z(n2522) );
  XOR U3055 ( .A(n2523), .B(n2522), .Z(n2525) );
  NAND U3056 ( .A(n2249), .B(n2248), .Z(n2253) );
  NAND U3057 ( .A(n2251), .B(n2250), .Z(n2252) );
  AND U3058 ( .A(n2253), .B(n2252), .Z(n2524) );
  XNOR U3059 ( .A(n2525), .B(n2524), .Z(n2646) );
  XOR U3060 ( .A(n2647), .B(n2646), .Z(n2648) );
  XOR U3061 ( .A(n2649), .B(n2648), .Z(n2536) );
  XOR U3062 ( .A(n2537), .B(n2536), .Z(n2540) );
  IV U3063 ( .A(n2540), .Z(n2541) );
  XOR U3064 ( .A(n2541), .B(n2542), .Z(n2258) );
  XNOR U3065 ( .A(n2543), .B(n2258), .Z(n2549) );
  NAND U3066 ( .A(n2260), .B(n2259), .Z(n2264) );
  NANDN U3067 ( .A(n2262), .B(n2261), .Z(n2263) );
  AND U3068 ( .A(n2264), .B(n2263), .Z(n2552) );
  NANDN U3069 ( .A(n2266), .B(n2265), .Z(n2270) );
  NANDN U3070 ( .A(n2268), .B(n2267), .Z(n2269) );
  NAND U3071 ( .A(n2270), .B(n2269), .Z(n2551) );
  NAND U3072 ( .A(n2272), .B(n2271), .Z(n2276) );
  NAND U3073 ( .A(n2274), .B(n2273), .Z(n2275) );
  NAND U3074 ( .A(n2276), .B(n2275), .Z(n2550) );
  XNOR U3075 ( .A(n2551), .B(n2550), .Z(n2553) );
  XNOR U3076 ( .A(n2548), .B(n2547), .Z(n2280) );
  XNOR U3077 ( .A(n2549), .B(n2280), .Z(o[2]) );
  NAND U3078 ( .A(n2282), .B(n2281), .Z(n2286) );
  NAND U3079 ( .A(n2284), .B(n2283), .Z(n2285) );
  NAND U3080 ( .A(n2286), .B(n2285), .Z(n2762) );
  NAND U3081 ( .A(n2288), .B(n2287), .Z(n2292) );
  NAND U3082 ( .A(n2290), .B(n2289), .Z(n2291) );
  AND U3083 ( .A(n2292), .B(n2291), .Z(n2760) );
  NAND U3084 ( .A(n2294), .B(n2293), .Z(n2298) );
  NAND U3085 ( .A(n2296), .B(n2295), .Z(n2297) );
  AND U3086 ( .A(n2298), .B(n2297), .Z(n2680) );
  NAND U3087 ( .A(n2300), .B(n2299), .Z(n2304) );
  NAND U3088 ( .A(n2302), .B(n2301), .Z(n2303) );
  NAND U3089 ( .A(n2304), .B(n2303), .Z(n2681) );
  NAND U3090 ( .A(n2306), .B(n2305), .Z(n2310) );
  NAND U3091 ( .A(n2308), .B(n2307), .Z(n2309) );
  NAND U3092 ( .A(n2310), .B(n2309), .Z(n2683) );
  XOR U3093 ( .A(n2760), .B(n2759), .Z(n2761) );
  XNOR U3094 ( .A(n2762), .B(n2761), .Z(n2791) );
  NAND U3095 ( .A(n2312), .B(n2311), .Z(n2316) );
  NAND U3096 ( .A(n2314), .B(n2313), .Z(n2315) );
  NAND U3097 ( .A(n2316), .B(n2315), .Z(n2750) );
  NAND U3098 ( .A(n2318), .B(n2317), .Z(n2322) );
  NAND U3099 ( .A(n2320), .B(n2319), .Z(n2321) );
  NAND U3100 ( .A(n2322), .B(n2321), .Z(n2748) );
  NANDN U3101 ( .A(n2324), .B(n2323), .Z(n2328) );
  NANDN U3102 ( .A(n2326), .B(n2325), .Z(n2327) );
  AND U3103 ( .A(n2328), .B(n2327), .Z(n2695) );
  NANDN U3104 ( .A(n2330), .B(n2329), .Z(n2334) );
  NAND U3105 ( .A(n2332), .B(n2331), .Z(n2333) );
  AND U3106 ( .A(n2334), .B(n2333), .Z(n2692) );
  NANDN U3107 ( .A(n2336), .B(n2335), .Z(n2340) );
  NANDN U3108 ( .A(n2338), .B(n2337), .Z(n2339) );
  AND U3109 ( .A(n2340), .B(n2339), .Z(n2693) );
  XOR U3110 ( .A(n2692), .B(n2693), .Z(n2694) );
  XOR U3111 ( .A(n2695), .B(n2694), .Z(n2747) );
  XOR U3112 ( .A(n2748), .B(n2747), .Z(n2749) );
  XNOR U3113 ( .A(n2750), .B(n2749), .Z(n2789) );
  NANDN U3114 ( .A(n2342), .B(n2341), .Z(n2346) );
  NAND U3115 ( .A(n2344), .B(n2343), .Z(n2345) );
  AND U3116 ( .A(n2346), .B(n2345), .Z(n2790) );
  XOR U3117 ( .A(n2789), .B(n2790), .Z(n2792) );
  XNOR U3118 ( .A(n2791), .B(n2792), .Z(n2809) );
  NANDN U3119 ( .A(n2348), .B(n2347), .Z(n2352) );
  NAND U3120 ( .A(n2350), .B(n2349), .Z(n2351) );
  AND U3121 ( .A(n2352), .B(n2351), .Z(n2807) );
  NANDN U3122 ( .A(n2354), .B(n2353), .Z(n2358) );
  NANDN U3123 ( .A(n2356), .B(n2355), .Z(n2357) );
  NAND U3124 ( .A(n2358), .B(n2357), .Z(n2808) );
  XOR U3125 ( .A(n2809), .B(n2810), .Z(n2668) );
  NANDN U3126 ( .A(n2360), .B(n2359), .Z(n2364) );
  NAND U3127 ( .A(n2362), .B(n2361), .Z(n2363) );
  NAND U3128 ( .A(n2364), .B(n2363), .Z(n2804) );
  NAND U3129 ( .A(n2366), .B(n2365), .Z(n2370) );
  NAND U3130 ( .A(n2368), .B(n2367), .Z(n2369) );
  NAND U3131 ( .A(n2370), .B(n2369), .Z(n2826) );
  NANDN U3132 ( .A(n2372), .B(n2371), .Z(n2376) );
  NAND U3133 ( .A(n2374), .B(n2373), .Z(n2375) );
  AND U3134 ( .A(n2376), .B(n2375), .Z(n2705) );
  NANDN U3135 ( .A(n2378), .B(n2377), .Z(n2382) );
  NANDN U3136 ( .A(n2380), .B(n2379), .Z(n2381) );
  AND U3137 ( .A(n2382), .B(n2381), .Z(n2704) );
  NANDN U3138 ( .A(n2384), .B(n2383), .Z(n2388) );
  NANDN U3139 ( .A(n2386), .B(n2385), .Z(n2387) );
  AND U3140 ( .A(n2388), .B(n2387), .Z(n2725) );
  NANDN U3141 ( .A(n2390), .B(n2389), .Z(n2394) );
  NANDN U3142 ( .A(n2392), .B(n2391), .Z(n2393) );
  AND U3143 ( .A(n2394), .B(n2393), .Z(n2723) );
  NANDN U3144 ( .A(n2396), .B(n2395), .Z(n2400) );
  NANDN U3145 ( .A(n2398), .B(n2397), .Z(n2399) );
  AND U3146 ( .A(n2400), .B(n2399), .Z(n2722) );
  XOR U3147 ( .A(n2723), .B(n2722), .Z(n2724) );
  XOR U3148 ( .A(n2725), .B(n2724), .Z(n2706) );
  XOR U3149 ( .A(n2707), .B(n2706), .Z(n2677) );
  NANDN U3150 ( .A(n2402), .B(n2401), .Z(n2406) );
  NANDN U3151 ( .A(n2404), .B(n2403), .Z(n2405) );
  AND U3152 ( .A(n2406), .B(n2405), .Z(n2713) );
  NANDN U3153 ( .A(n2408), .B(n2407), .Z(n2412) );
  NANDN U3154 ( .A(n2410), .B(n2409), .Z(n2411) );
  AND U3155 ( .A(n2412), .B(n2411), .Z(n2711) );
  AND U3156 ( .A(n2413), .B(oglobal[2]), .Z(n2740) );
  XOR U3157 ( .A(oglobal[3]), .B(n2740), .Z(n2710) );
  XOR U3158 ( .A(n2711), .B(n2710), .Z(n2712) );
  XNOR U3159 ( .A(n2713), .B(n2712), .Z(n2675) );
  NANDN U3160 ( .A(n2415), .B(n2414), .Z(n2419) );
  NANDN U3161 ( .A(n2417), .B(n2416), .Z(n2418) );
  AND U3162 ( .A(n2419), .B(n2418), .Z(n2674) );
  XOR U3163 ( .A(n2675), .B(n2674), .Z(n2676) );
  XOR U3164 ( .A(n2677), .B(n2676), .Z(n2825) );
  XOR U3165 ( .A(n2826), .B(n2825), .Z(n2828) );
  NAND U3166 ( .A(n2421), .B(n2420), .Z(n2425) );
  NAND U3167 ( .A(n2423), .B(n2422), .Z(n2424) );
  NAND U3168 ( .A(n2425), .B(n2424), .Z(n2768) );
  NAND U3169 ( .A(n2427), .B(n2426), .Z(n2431) );
  NAND U3170 ( .A(n2429), .B(n2428), .Z(n2430) );
  NAND U3171 ( .A(n2431), .B(n2430), .Z(n2766) );
  NAND U3172 ( .A(n2433), .B(n2432), .Z(n2437) );
  NAND U3173 ( .A(n2435), .B(n2434), .Z(n2436) );
  NAND U3174 ( .A(n2437), .B(n2436), .Z(n2765) );
  XOR U3175 ( .A(n2766), .B(n2765), .Z(n2767) );
  XOR U3176 ( .A(n2768), .B(n2767), .Z(n2827) );
  XNOR U3177 ( .A(n2828), .B(n2827), .Z(n2802) );
  NAND U3178 ( .A(n2439), .B(n2438), .Z(n2443) );
  NAND U3179 ( .A(n2441), .B(n2440), .Z(n2442) );
  AND U3180 ( .A(n2443), .B(n2442), .Z(n2786) );
  NANDN U3181 ( .A(n2445), .B(n2444), .Z(n2449) );
  NAND U3182 ( .A(n2447), .B(n2446), .Z(n2448) );
  AND U3183 ( .A(n2449), .B(n2448), .Z(n2731) );
  NANDN U3184 ( .A(n2451), .B(n2450), .Z(n2455) );
  NANDN U3185 ( .A(n2453), .B(n2452), .Z(n2454) );
  AND U3186 ( .A(n2455), .B(n2454), .Z(n2729) );
  NANDN U3187 ( .A(n2457), .B(n2456), .Z(n2461) );
  NANDN U3188 ( .A(n2459), .B(n2458), .Z(n2460) );
  NAND U3189 ( .A(n2461), .B(n2460), .Z(n2728) );
  NAND U3190 ( .A(n2463), .B(n2462), .Z(n2467) );
  NAND U3191 ( .A(n2465), .B(n2464), .Z(n2466) );
  AND U3192 ( .A(n2467), .B(n2466), .Z(n2699) );
  NANDN U3193 ( .A(n2469), .B(n2468), .Z(n2473) );
  NANDN U3194 ( .A(n2471), .B(n2470), .Z(n2472) );
  AND U3195 ( .A(n2473), .B(n2472), .Z(n2737) );
  NANDN U3196 ( .A(n2475), .B(n2474), .Z(n2479) );
  NANDN U3197 ( .A(n2477), .B(n2476), .Z(n2478) );
  AND U3198 ( .A(n2479), .B(n2478), .Z(n2734) );
  NANDN U3199 ( .A(n2481), .B(n2480), .Z(n2485) );
  NANDN U3200 ( .A(n2483), .B(n2482), .Z(n2484) );
  NAND U3201 ( .A(n2485), .B(n2484), .Z(n2735) );
  XOR U3202 ( .A(n2737), .B(n2736), .Z(n2698) );
  XNOR U3203 ( .A(n2700), .B(n2701), .Z(n2783) );
  NAND U3204 ( .A(n2487), .B(n2486), .Z(n2491) );
  NAND U3205 ( .A(n2489), .B(n2488), .Z(n2490) );
  AND U3206 ( .A(n2491), .B(n2490), .Z(n2784) );
  XOR U3207 ( .A(n2783), .B(n2784), .Z(n2785) );
  XOR U3208 ( .A(n2786), .B(n2785), .Z(n2801) );
  XOR U3209 ( .A(n2802), .B(n2801), .Z(n2803) );
  XOR U3210 ( .A(n2804), .B(n2803), .Z(n2666) );
  NANDN U3211 ( .A(n2493), .B(n2492), .Z(n2497) );
  NAND U3212 ( .A(n2495), .B(n2494), .Z(n2496) );
  NAND U3213 ( .A(n2497), .B(n2496), .Z(n2816) );
  OR U3214 ( .A(n2499), .B(n2498), .Z(n2503) );
  NAND U3215 ( .A(n2501), .B(n2500), .Z(n2502) );
  NAND U3216 ( .A(n2503), .B(n2502), .Z(n2814) );
  NAND U3217 ( .A(n2505), .B(n2504), .Z(n2509) );
  NAND U3218 ( .A(n2507), .B(n2506), .Z(n2508) );
  NAND U3219 ( .A(n2509), .B(n2508), .Z(n2813) );
  XOR U3220 ( .A(n2814), .B(n2813), .Z(n2815) );
  XNOR U3221 ( .A(n2816), .B(n2815), .Z(n2832) );
  NANDN U3222 ( .A(n2511), .B(n2510), .Z(n2515) );
  NANDN U3223 ( .A(n2513), .B(n2512), .Z(n2514) );
  AND U3224 ( .A(n2515), .B(n2514), .Z(n2822) );
  NAND U3225 ( .A(n2517), .B(n2516), .Z(n2521) );
  NAND U3226 ( .A(n2519), .B(n2518), .Z(n2520) );
  NAND U3227 ( .A(n2521), .B(n2520), .Z(n2820) );
  NAND U3228 ( .A(n2523), .B(n2522), .Z(n2527) );
  NAND U3229 ( .A(n2525), .B(n2524), .Z(n2526) );
  NAND U3230 ( .A(n2527), .B(n2526), .Z(n2819) );
  XOR U3231 ( .A(n2820), .B(n2819), .Z(n2821) );
  XOR U3232 ( .A(n2822), .B(n2821), .Z(n2831) );
  XOR U3233 ( .A(n2832), .B(n2831), .Z(n2834) );
  NANDN U3234 ( .A(n2529), .B(n2528), .Z(n2533) );
  NAND U3235 ( .A(n2531), .B(n2530), .Z(n2532) );
  AND U3236 ( .A(n2533), .B(n2532), .Z(n2833) );
  XNOR U3237 ( .A(n2834), .B(n2833), .Z(n2665) );
  NAND U3238 ( .A(n2535), .B(n2534), .Z(n2539) );
  NAND U3239 ( .A(n2537), .B(n2536), .Z(n2538) );
  NAND U3240 ( .A(n2539), .B(n2538), .Z(n2653) );
  OR U3241 ( .A(n2542), .B(n2540), .Z(n2546) );
  ANDN U3242 ( .B(n2542), .A(n2541), .Z(n2544) );
  OR U3243 ( .A(n2544), .B(n2543), .Z(n2545) );
  AND U3244 ( .A(n2546), .B(n2545), .Z(n2654) );
  XOR U3245 ( .A(n2653), .B(n2654), .Z(n2655) );
  NAND U3246 ( .A(n2551), .B(n2550), .Z(n2555) );
  NANDN U3247 ( .A(n2553), .B(n2552), .Z(n2554) );
  NAND U3248 ( .A(n2555), .B(n2554), .Z(n2661) );
  NANDN U3249 ( .A(n2557), .B(n2556), .Z(n2561) );
  NAND U3250 ( .A(n2559), .B(n2558), .Z(n2560) );
  AND U3251 ( .A(n2561), .B(n2560), .Z(n2660) );
  NAND U3252 ( .A(n2563), .B(n2562), .Z(n2567) );
  NAND U3253 ( .A(n2565), .B(n2564), .Z(n2566) );
  AND U3254 ( .A(n2567), .B(n2566), .Z(n2798) );
  NAND U3255 ( .A(n2569), .B(n2568), .Z(n2573) );
  NAND U3256 ( .A(n2571), .B(n2570), .Z(n2572) );
  AND U3257 ( .A(n2573), .B(n2572), .Z(n2780) );
  NAND U3258 ( .A(n2575), .B(n2574), .Z(n2579) );
  NAND U3259 ( .A(n2577), .B(n2576), .Z(n2578) );
  AND U3260 ( .A(n2579), .B(n2578), .Z(n2778) );
  NAND U3261 ( .A(n2581), .B(n2580), .Z(n2585) );
  NAND U3262 ( .A(n2583), .B(n2582), .Z(n2584) );
  AND U3263 ( .A(n2585), .B(n2584), .Z(n2719) );
  NAND U3264 ( .A(n2587), .B(n2586), .Z(n2591) );
  NAND U3265 ( .A(n2589), .B(n2588), .Z(n2590) );
  AND U3266 ( .A(n2591), .B(n2590), .Z(n2716) );
  NAND U3267 ( .A(n2593), .B(n2592), .Z(n2597) );
  NAND U3268 ( .A(n2595), .B(n2594), .Z(n2596) );
  NAND U3269 ( .A(n2597), .B(n2596), .Z(n2717) );
  XOR U3270 ( .A(n2719), .B(n2718), .Z(n2777) );
  NAND U3271 ( .A(n2599), .B(n2598), .Z(n2603) );
  NANDN U3272 ( .A(n2601), .B(n2600), .Z(n2602) );
  AND U3273 ( .A(n2603), .B(n2602), .Z(n2774) );
  NAND U3274 ( .A(n2605), .B(n2604), .Z(n2609) );
  NANDN U3275 ( .A(n2607), .B(n2606), .Z(n2608) );
  AND U3276 ( .A(n2609), .B(n2608), .Z(n2744) );
  NAND U3277 ( .A(n2611), .B(n2610), .Z(n2615) );
  NANDN U3278 ( .A(n2613), .B(n2612), .Z(n2614) );
  AND U3279 ( .A(n2615), .B(n2614), .Z(n2741) );
  NAND U3280 ( .A(n2617), .B(n2616), .Z(n2621) );
  NAND U3281 ( .A(n2619), .B(n2618), .Z(n2620) );
  NAND U3282 ( .A(n2621), .B(n2620), .Z(n2742) );
  XOR U3283 ( .A(n2744), .B(n2743), .Z(n2772) );
  NAND U3284 ( .A(n2623), .B(n2622), .Z(n2627) );
  NAND U3285 ( .A(n2625), .B(n2624), .Z(n2626) );
  AND U3286 ( .A(n2627), .B(n2626), .Z(n2771) );
  XNOR U3287 ( .A(n2774), .B(n2773), .Z(n2754) );
  NAND U3288 ( .A(n2629), .B(n2628), .Z(n2633) );
  NAND U3289 ( .A(n2631), .B(n2630), .Z(n2632) );
  AND U3290 ( .A(n2633), .B(n2632), .Z(n2686) );
  NAND U3291 ( .A(n2635), .B(n2634), .Z(n2639) );
  NAND U3292 ( .A(n2637), .B(n2636), .Z(n2638) );
  NAND U3293 ( .A(n2639), .B(n2638), .Z(n2687) );
  NAND U3294 ( .A(n2641), .B(n2640), .Z(n2645) );
  NAND U3295 ( .A(n2643), .B(n2642), .Z(n2644) );
  AND U3296 ( .A(n2645), .B(n2644), .Z(n2688) );
  XNOR U3297 ( .A(n2689), .B(n2688), .Z(n2753) );
  XOR U3298 ( .A(n2754), .B(n2753), .Z(n2755) );
  XNOR U3299 ( .A(n2756), .B(n2755), .Z(n2796) );
  NAND U3300 ( .A(n2647), .B(n2646), .Z(n2651) );
  NAND U3301 ( .A(n2649), .B(n2648), .Z(n2650) );
  NAND U3302 ( .A(n2651), .B(n2650), .Z(n2795) );
  XOR U3303 ( .A(n2796), .B(n2795), .Z(n2797) );
  XOR U3304 ( .A(n2798), .B(n2797), .Z(n2659) );
  XOR U3305 ( .A(n2660), .B(n2659), .Z(n2662) );
  XOR U3306 ( .A(n2661), .B(n2662), .Z(n2673) );
  XNOR U3307 ( .A(n2672), .B(n2673), .Z(n2652) );
  XOR U3308 ( .A(n2671), .B(n2652), .Z(o[3]) );
  NAND U3309 ( .A(n2654), .B(n2653), .Z(n2658) );
  NANDN U3310 ( .A(n2656), .B(n2655), .Z(n2657) );
  AND U3311 ( .A(n2658), .B(n2657), .Z(n2927) );
  NAND U3312 ( .A(n2660), .B(n2659), .Z(n2664) );
  NAND U3313 ( .A(n2662), .B(n2661), .Z(n2663) );
  AND U3314 ( .A(n2664), .B(n2663), .Z(n2925) );
  NANDN U3315 ( .A(n2666), .B(n2665), .Z(n2670) );
  NANDN U3316 ( .A(n2668), .B(n2667), .Z(n2669) );
  NAND U3317 ( .A(n2670), .B(n2669), .Z(n2924) );
  XOR U3318 ( .A(n2925), .B(n2924), .Z(n2926) );
  XNOR U3319 ( .A(n2927), .B(n2926), .Z(n2923) );
  NAND U3320 ( .A(n2675), .B(n2674), .Z(n2679) );
  NANDN U3321 ( .A(n2677), .B(n2676), .Z(n2678) );
  AND U3322 ( .A(n2679), .B(n2678), .Z(n2900) );
  NANDN U3323 ( .A(n2681), .B(n2680), .Z(n2685) );
  NANDN U3324 ( .A(n2683), .B(n2682), .Z(n2684) );
  AND U3325 ( .A(n2685), .B(n2684), .Z(n2897) );
  NANDN U3326 ( .A(n2687), .B(n2686), .Z(n2691) );
  NAND U3327 ( .A(n2689), .B(n2688), .Z(n2690) );
  NAND U3328 ( .A(n2691), .B(n2690), .Z(n2898) );
  XOR U3329 ( .A(n2900), .B(n2899), .Z(n2888) );
  NAND U3330 ( .A(n2693), .B(n2692), .Z(n2697) );
  NAND U3331 ( .A(n2695), .B(n2694), .Z(n2696) );
  AND U3332 ( .A(n2697), .B(n2696), .Z(n2886) );
  NANDN U3333 ( .A(n2699), .B(n2698), .Z(n2703) );
  NAND U3334 ( .A(n2701), .B(n2700), .Z(n2702) );
  AND U3335 ( .A(n2703), .B(n2702), .Z(n2885) );
  NANDN U3336 ( .A(n2705), .B(n2704), .Z(n2709) );
  NAND U3337 ( .A(n2707), .B(n2706), .Z(n2708) );
  AND U3338 ( .A(n2709), .B(n2708), .Z(n2877) );
  NAND U3339 ( .A(n2711), .B(n2710), .Z(n2715) );
  NAND U3340 ( .A(n2713), .B(n2712), .Z(n2714) );
  AND U3341 ( .A(n2715), .B(n2714), .Z(n2875) );
  NANDN U3342 ( .A(n2717), .B(n2716), .Z(n2721) );
  NAND U3343 ( .A(n2719), .B(n2718), .Z(n2720) );
  NAND U3344 ( .A(n2721), .B(n2720), .Z(n2874) );
  NAND U3345 ( .A(n2723), .B(n2722), .Z(n2727) );
  NAND U3346 ( .A(n2725), .B(n2724), .Z(n2726) );
  AND U3347 ( .A(n2727), .B(n2726), .Z(n2869) );
  NANDN U3348 ( .A(n2729), .B(n2728), .Z(n2733) );
  NANDN U3349 ( .A(n2731), .B(n2730), .Z(n2732) );
  AND U3350 ( .A(n2733), .B(n2732), .Z(n2868) );
  NANDN U3351 ( .A(n2735), .B(n2734), .Z(n2739) );
  NAND U3352 ( .A(n2737), .B(n2736), .Z(n2738) );
  AND U3353 ( .A(n2739), .B(n2738), .Z(n2882) );
  NAND U3354 ( .A(n2740), .B(oglobal[3]), .Z(n2880) );
  XOR U3355 ( .A(n2871), .B(n2870), .Z(n2863) );
  NANDN U3356 ( .A(n2742), .B(n2741), .Z(n2746) );
  NAND U3357 ( .A(n2744), .B(n2743), .Z(n2745) );
  AND U3358 ( .A(n2746), .B(n2745), .Z(n2862) );
  XOR U3359 ( .A(n2864), .B(n2865), .Z(n2916) );
  NAND U3360 ( .A(n2748), .B(n2747), .Z(n2752) );
  NAND U3361 ( .A(n2750), .B(n2749), .Z(n2751) );
  AND U3362 ( .A(n2752), .B(n2751), .Z(n2915) );
  NAND U3363 ( .A(n2754), .B(n2753), .Z(n2758) );
  NAND U3364 ( .A(n2756), .B(n2755), .Z(n2757) );
  AND U3365 ( .A(n2758), .B(n2757), .Z(n2912) );
  NAND U3366 ( .A(n2760), .B(n2759), .Z(n2764) );
  NAND U3367 ( .A(n2762), .B(n2761), .Z(n2763) );
  NAND U3368 ( .A(n2764), .B(n2763), .Z(n2909) );
  NAND U3369 ( .A(n2766), .B(n2765), .Z(n2770) );
  NAND U3370 ( .A(n2768), .B(n2767), .Z(n2769) );
  AND U3371 ( .A(n2770), .B(n2769), .Z(n2894) );
  NANDN U3372 ( .A(n2772), .B(n2771), .Z(n2776) );
  NAND U3373 ( .A(n2774), .B(n2773), .Z(n2775) );
  AND U3374 ( .A(n2776), .B(n2775), .Z(n2892) );
  NANDN U3375 ( .A(n2778), .B(n2777), .Z(n2782) );
  NANDN U3376 ( .A(n2780), .B(n2779), .Z(n2781) );
  AND U3377 ( .A(n2782), .B(n2781), .Z(n2891) );
  XOR U3378 ( .A(n2894), .B(n2893), .Z(n2910) );
  XOR U3379 ( .A(n2909), .B(n2910), .Z(n2911) );
  XNOR U3380 ( .A(n2912), .B(n2911), .Z(n2851) );
  NAND U3381 ( .A(n2784), .B(n2783), .Z(n2788) );
  NAND U3382 ( .A(n2786), .B(n2785), .Z(n2787) );
  AND U3383 ( .A(n2788), .B(n2787), .Z(n2850) );
  XOR U3384 ( .A(n2851), .B(n2850), .Z(n2852) );
  XOR U3385 ( .A(n2853), .B(n2852), .Z(n2847) );
  NAND U3386 ( .A(n2790), .B(n2789), .Z(n2794) );
  NAND U3387 ( .A(n2792), .B(n2791), .Z(n2793) );
  AND U3388 ( .A(n2794), .B(n2793), .Z(n2906) );
  NAND U3389 ( .A(n2796), .B(n2795), .Z(n2800) );
  NAND U3390 ( .A(n2798), .B(n2797), .Z(n2799) );
  NAND U3391 ( .A(n2800), .B(n2799), .Z(n2904) );
  NAND U3392 ( .A(n2802), .B(n2801), .Z(n2806) );
  NAND U3393 ( .A(n2804), .B(n2803), .Z(n2805) );
  NAND U3394 ( .A(n2806), .B(n2805), .Z(n2903) );
  XOR U3395 ( .A(n2904), .B(n2903), .Z(n2905) );
  XOR U3396 ( .A(n2906), .B(n2905), .Z(n2845) );
  NANDN U3397 ( .A(n2808), .B(n2807), .Z(n2812) );
  NAND U3398 ( .A(n2810), .B(n2809), .Z(n2811) );
  AND U3399 ( .A(n2812), .B(n2811), .Z(n2841) );
  NAND U3400 ( .A(n2814), .B(n2813), .Z(n2818) );
  NAND U3401 ( .A(n2816), .B(n2815), .Z(n2817) );
  NAND U3402 ( .A(n2818), .B(n2817), .Z(n2859) );
  NAND U3403 ( .A(n2820), .B(n2819), .Z(n2824) );
  NANDN U3404 ( .A(n2822), .B(n2821), .Z(n2823) );
  NAND U3405 ( .A(n2824), .B(n2823), .Z(n2857) );
  NAND U3406 ( .A(n2826), .B(n2825), .Z(n2830) );
  NAND U3407 ( .A(n2828), .B(n2827), .Z(n2829) );
  NAND U3408 ( .A(n2830), .B(n2829), .Z(n2856) );
  XOR U3409 ( .A(n2857), .B(n2856), .Z(n2858) );
  XNOR U3410 ( .A(n2859), .B(n2858), .Z(n2839) );
  NAND U3411 ( .A(n2832), .B(n2831), .Z(n2836) );
  NAND U3412 ( .A(n2834), .B(n2833), .Z(n2835) );
  NAND U3413 ( .A(n2836), .B(n2835), .Z(n2838) );
  XOR U3414 ( .A(n2839), .B(n2838), .Z(n2840) );
  XOR U3415 ( .A(n2845), .B(n2844), .Z(n2846) );
  XOR U3416 ( .A(n2922), .B(n2921), .Z(n2837) );
  XNOR U3417 ( .A(n2923), .B(n2837), .Z(o[4]) );
  NAND U3418 ( .A(n2839), .B(n2838), .Z(n2843) );
  NANDN U3419 ( .A(n2841), .B(n2840), .Z(n2842) );
  NAND U3420 ( .A(n2843), .B(n2842), .Z(n2932) );
  NAND U3421 ( .A(n2845), .B(n2844), .Z(n2849) );
  NANDN U3422 ( .A(n2847), .B(n2846), .Z(n2848) );
  NAND U3423 ( .A(n2849), .B(n2848), .Z(n2931) );
  XOR U3424 ( .A(n2932), .B(n2931), .Z(n2934) );
  NAND U3425 ( .A(n2851), .B(n2850), .Z(n2855) );
  NAND U3426 ( .A(n2853), .B(n2852), .Z(n2854) );
  AND U3427 ( .A(n2855), .B(n2854), .Z(n2941) );
  NAND U3428 ( .A(n2857), .B(n2856), .Z(n2861) );
  NAND U3429 ( .A(n2859), .B(n2858), .Z(n2860) );
  AND U3430 ( .A(n2861), .B(n2860), .Z(n2955) );
  NANDN U3431 ( .A(n2863), .B(n2862), .Z(n2867) );
  NAND U3432 ( .A(n2865), .B(n2864), .Z(n2866) );
  AND U3433 ( .A(n2867), .B(n2866), .Z(n2961) );
  NANDN U3434 ( .A(n2869), .B(n2868), .Z(n2873) );
  NAND U3435 ( .A(n2871), .B(n2870), .Z(n2872) );
  AND U3436 ( .A(n2873), .B(n2872), .Z(n2959) );
  NANDN U3437 ( .A(n2875), .B(n2874), .Z(n2879) );
  NANDN U3438 ( .A(n2877), .B(n2876), .Z(n2878) );
  NAND U3439 ( .A(n2879), .B(n2878), .Z(n2965) );
  NANDN U3440 ( .A(n2880), .B(oglobal[4]), .Z(n2884) );
  NANDN U3441 ( .A(n2882), .B(n2881), .Z(n2883) );
  NAND U3442 ( .A(n2884), .B(n2883), .Z(n2964) );
  XOR U3443 ( .A(n2964), .B(oglobal[5]), .Z(n2966) );
  XOR U3444 ( .A(n2965), .B(n2966), .Z(n2958) );
  XOR U3445 ( .A(n2961), .B(n2960), .Z(n2953) );
  NANDN U3446 ( .A(n2886), .B(n2885), .Z(n2890) );
  NANDN U3447 ( .A(n2888), .B(n2887), .Z(n2889) );
  AND U3448 ( .A(n2890), .B(n2889), .Z(n2972) );
  NANDN U3449 ( .A(n2892), .B(n2891), .Z(n2896) );
  NAND U3450 ( .A(n2894), .B(n2893), .Z(n2895) );
  AND U3451 ( .A(n2896), .B(n2895), .Z(n2970) );
  NANDN U3452 ( .A(n2898), .B(n2897), .Z(n2902) );
  NAND U3453 ( .A(n2900), .B(n2899), .Z(n2901) );
  AND U3454 ( .A(n2902), .B(n2901), .Z(n2969) );
  XOR U3455 ( .A(n2955), .B(n2954), .Z(n2940) );
  XOR U3456 ( .A(n2941), .B(n2940), .Z(n2943) );
  NAND U3457 ( .A(n2904), .B(n2903), .Z(n2908) );
  NAND U3458 ( .A(n2906), .B(n2905), .Z(n2907) );
  NAND U3459 ( .A(n2908), .B(n2907), .Z(n2948) );
  NAND U3460 ( .A(n2910), .B(n2909), .Z(n2914) );
  NAND U3461 ( .A(n2912), .B(n2911), .Z(n2913) );
  NAND U3462 ( .A(n2914), .B(n2913), .Z(n2946) );
  NANDN U3463 ( .A(n2916), .B(n2915), .Z(n2920) );
  NANDN U3464 ( .A(n2918), .B(n2917), .Z(n2919) );
  AND U3465 ( .A(n2920), .B(n2919), .Z(n2947) );
  XOR U3466 ( .A(n2946), .B(n2947), .Z(n2949) );
  XOR U3467 ( .A(n2948), .B(n2949), .Z(n2942) );
  XOR U3468 ( .A(n2943), .B(n2942), .Z(n2933) );
  XOR U3469 ( .A(n2934), .B(n2933), .Z(n2937) );
  NAND U3470 ( .A(n2925), .B(n2924), .Z(n2929) );
  NAND U3471 ( .A(n2927), .B(n2926), .Z(n2928) );
  AND U3472 ( .A(n2929), .B(n2928), .Z(n2939) );
  XNOR U3473 ( .A(n2938), .B(n2939), .Z(n2930) );
  XOR U3474 ( .A(n2937), .B(n2930), .Z(o[5]) );
  NAND U3475 ( .A(n2932), .B(n2931), .Z(n2936) );
  NAND U3476 ( .A(n2934), .B(n2933), .Z(n2935) );
  AND U3477 ( .A(n2936), .B(n2935), .Z(n2996) );
  NAND U3478 ( .A(n2941), .B(n2940), .Z(n2945) );
  NAND U3479 ( .A(n2943), .B(n2942), .Z(n2944) );
  NAND U3480 ( .A(n2945), .B(n2944), .Z(n2978) );
  NAND U3481 ( .A(n2947), .B(n2946), .Z(n2951) );
  NAND U3482 ( .A(n2949), .B(n2948), .Z(n2950) );
  NAND U3483 ( .A(n2951), .B(n2950), .Z(n2976) );
  NANDN U3484 ( .A(n2953), .B(n2952), .Z(n2957) );
  NAND U3485 ( .A(n2955), .B(n2954), .Z(n2956) );
  AND U3486 ( .A(n2957), .B(n2956), .Z(n2985) );
  NANDN U3487 ( .A(n2959), .B(n2958), .Z(n2963) );
  NAND U3488 ( .A(n2961), .B(n2960), .Z(n2962) );
  NAND U3489 ( .A(n2963), .B(n2962), .Z(n2988) );
  XOR U3490 ( .A(n2988), .B(oglobal[6]), .Z(n2990) );
  NAND U3491 ( .A(oglobal[5]), .B(n2964), .Z(n2968) );
  NAND U3492 ( .A(n2966), .B(n2965), .Z(n2967) );
  NAND U3493 ( .A(n2968), .B(n2967), .Z(n2989) );
  XOR U3494 ( .A(n2990), .B(n2989), .Z(n2983) );
  NANDN U3495 ( .A(n2970), .B(n2969), .Z(n2974) );
  NANDN U3496 ( .A(n2972), .B(n2971), .Z(n2973) );
  NAND U3497 ( .A(n2974), .B(n2973), .Z(n2982) );
  XOR U3498 ( .A(n2976), .B(n2977), .Z(n2979) );
  XNOR U3499 ( .A(n2978), .B(n2979), .Z(n2995) );
  IV U3500 ( .A(n2995), .Z(n2993) );
  XOR U3501 ( .A(n2994), .B(n2993), .Z(n2975) );
  XNOR U3502 ( .A(n2996), .B(n2975), .Z(o[6]) );
  NANDN U3503 ( .A(n2977), .B(n2976), .Z(n2981) );
  NANDN U3504 ( .A(n2979), .B(n2978), .Z(n2980) );
  AND U3505 ( .A(n2981), .B(n2980), .Z(n3008) );
  NANDN U3506 ( .A(n2983), .B(n2982), .Z(n2987) );
  NANDN U3507 ( .A(n2985), .B(n2984), .Z(n2986) );
  AND U3508 ( .A(n2987), .B(n2986), .Z(n3003) );
  NAND U3509 ( .A(oglobal[6]), .B(n2988), .Z(n2992) );
  NAND U3510 ( .A(n2990), .B(n2989), .Z(n2991) );
  NAND U3511 ( .A(n2992), .B(n2991), .Z(n3001) );
  XOR U3512 ( .A(oglobal[7]), .B(n3001), .Z(n3002) );
  XOR U3513 ( .A(n3003), .B(n3002), .Z(n3007) );
  NANDN U3514 ( .A(n2993), .B(n2994), .Z(n2999) );
  NOR U3515 ( .A(n2995), .B(n2994), .Z(n2997) );
  OR U3516 ( .A(n2997), .B(n2996), .Z(n2998) );
  AND U3517 ( .A(n2999), .B(n2998), .Z(n3006) );
  XNOR U3518 ( .A(n3007), .B(n3006), .Z(n3000) );
  XNOR U3519 ( .A(n3008), .B(n3000), .Z(o[7]) );
  NAND U3520 ( .A(oglobal[7]), .B(n3001), .Z(n3005) );
  NAND U3521 ( .A(n3003), .B(n3002), .Z(n3004) );
  AND U3522 ( .A(n3005), .B(n3004), .Z(n3011) );
  XOR U3523 ( .A(n3010), .B(oglobal[8]), .Z(n3009) );
  XNOR U3524 ( .A(n3011), .B(n3009), .Z(o[8]) );
  XNOR U3525 ( .A(n3012), .B(oglobal[9]), .Z(o[9]) );
  ANDN U3526 ( .B(oglobal[9]), .A(n3012), .Z(n3013) );
  XOR U3527 ( .A(n3013), .B(oglobal[10]), .Z(o[10]) );
  AND U3528 ( .A(n3013), .B(oglobal[10]), .Z(n3014) );
  XOR U3529 ( .A(n3014), .B(oglobal[11]), .Z(o[11]) );
  AND U3530 ( .A(n3014), .B(oglobal[11]), .Z(n3015) );
  XOR U3531 ( .A(oglobal[12]), .B(n3015), .Z(o[12]) );
endmodule

