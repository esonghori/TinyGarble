
module hamming_N1600_CC16 ( clk, rst, x, y, o );
  input [99:0] x;
  input [99:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U103 ( .A(n93), .B(n92), .Z(n1) );
  NANDN U104 ( .A(n91), .B(n90), .Z(n2) );
  AND U105 ( .A(n1), .B(n2), .Z(n414) );
  NAND U106 ( .A(n393), .B(n392), .Z(n3) );
  NANDN U107 ( .A(n391), .B(n390), .Z(n4) );
  NAND U108 ( .A(n3), .B(n4), .Z(n531) );
  XOR U109 ( .A(n476), .B(n475), .Z(n5) );
  NANDN U110 ( .A(n474), .B(n5), .Z(n6) );
  NAND U111 ( .A(n476), .B(n475), .Z(n7) );
  AND U112 ( .A(n6), .B(n7), .Z(n525) );
  XOR U113 ( .A(n89), .B(n88), .Z(n8) );
  NANDN U114 ( .A(n87), .B(n8), .Z(n9) );
  NAND U115 ( .A(n89), .B(n88), .Z(n10) );
  AND U116 ( .A(n9), .B(n10), .Z(n413) );
  OR U117 ( .A(n245), .B(n246), .Z(n11) );
  NANDN U118 ( .A(n248), .B(n247), .Z(n12) );
  AND U119 ( .A(n11), .B(n12), .Z(n424) );
  XOR U120 ( .A(n302), .B(n301), .Z(n13) );
  NANDN U121 ( .A(n300), .B(n13), .Z(n14) );
  NAND U122 ( .A(n302), .B(n301), .Z(n15) );
  AND U123 ( .A(n14), .B(n15), .Z(n483) );
  XOR U124 ( .A(n210), .B(n209), .Z(n16) );
  NANDN U125 ( .A(n208), .B(n16), .Z(n17) );
  NAND U126 ( .A(n210), .B(n209), .Z(n18) );
  AND U127 ( .A(n17), .B(n18), .Z(n474) );
  NAND U128 ( .A(n534), .B(n533), .Z(n19) );
  NANDN U129 ( .A(n532), .B(n531), .Z(n20) );
  NAND U130 ( .A(n19), .B(n20), .Z(n565) );
  XOR U131 ( .A(n369), .B(n368), .Z(n21) );
  NANDN U132 ( .A(n367), .B(n21), .Z(n22) );
  NAND U133 ( .A(n369), .B(n368), .Z(n23) );
  AND U134 ( .A(n22), .B(n23), .Z(n543) );
  OR U135 ( .A(n241), .B(n242), .Z(n24) );
  NANDN U136 ( .A(n244), .B(n243), .Z(n25) );
  AND U137 ( .A(n24), .B(n25), .Z(n423) );
  OR U138 ( .A(n296), .B(n295), .Z(n26) );
  NANDN U139 ( .A(n298), .B(n297), .Z(n27) );
  NAND U140 ( .A(n26), .B(n27), .Z(n444) );
  NAND U141 ( .A(n305), .B(n306), .Z(n28) );
  NANDN U142 ( .A(n304), .B(n303), .Z(n29) );
  NAND U143 ( .A(n28), .B(n29), .Z(n455) );
  XOR U144 ( .A(n249), .B(n250), .Z(n30) );
  NANDN U145 ( .A(n251), .B(n30), .Z(n31) );
  NAND U146 ( .A(n249), .B(n250), .Z(n32) );
  AND U147 ( .A(n31), .B(n32), .Z(n388) );
  NANDN U148 ( .A(n416), .B(n415), .Z(n33) );
  NANDN U149 ( .A(n414), .B(n413), .Z(n34) );
  AND U150 ( .A(n33), .B(n34), .Z(n535) );
  NAND U151 ( .A(n524), .B(n523), .Z(n35) );
  XOR U152 ( .A(n523), .B(n524), .Z(n36) );
  NAND U153 ( .A(n36), .B(n522), .Z(n37) );
  NAND U154 ( .A(n35), .B(n37), .Z(n556) );
  XOR U155 ( .A(n578), .B(n579), .Z(n572) );
  XOR U156 ( .A(n545), .B(n544), .Z(n38) );
  NANDN U157 ( .A(n543), .B(n38), .Z(n39) );
  NAND U158 ( .A(n545), .B(n544), .Z(n40) );
  AND U159 ( .A(n39), .B(n40), .Z(n553) );
  OR U160 ( .A(n383), .B(n384), .Z(n41) );
  NANDN U161 ( .A(n386), .B(n385), .Z(n42) );
  AND U162 ( .A(n41), .B(n42), .Z(n492) );
  OR U163 ( .A(n177), .B(n176), .Z(n43) );
  NANDN U164 ( .A(n179), .B(n178), .Z(n44) );
  NAND U165 ( .A(n43), .B(n44), .Z(n439) );
  OR U166 ( .A(n111), .B(n110), .Z(n45) );
  NANDN U167 ( .A(n113), .B(n112), .Z(n46) );
  NAND U168 ( .A(n45), .B(n46), .Z(n470) );
  NAND U169 ( .A(n182), .B(n183), .Z(n47) );
  NANDN U170 ( .A(n181), .B(n180), .Z(n48) );
  NAND U171 ( .A(n47), .B(n48), .Z(n477) );
  NAND U172 ( .A(n86), .B(n85), .Z(n49) );
  NANDN U173 ( .A(n84), .B(n83), .Z(n50) );
  AND U174 ( .A(n49), .B(n50), .Z(n416) );
  XOR U175 ( .A(n511), .B(n512), .Z(n536) );
  XOR U176 ( .A(n388), .B(n387), .Z(n51) );
  NANDN U177 ( .A(n389), .B(n51), .Z(n52) );
  NAND U178 ( .A(n388), .B(n387), .Z(n53) );
  AND U179 ( .A(n52), .B(n53), .Z(n532) );
  XOR U180 ( .A(n445), .B(n444), .Z(n54) );
  NANDN U181 ( .A(n443), .B(n54), .Z(n55) );
  NAND U182 ( .A(n445), .B(n444), .Z(n56) );
  AND U183 ( .A(n55), .B(n56), .Z(n503) );
  NAND U184 ( .A(n460), .B(n459), .Z(n57) );
  XOR U185 ( .A(n459), .B(n460), .Z(n58) );
  NANDN U186 ( .A(n461), .B(n58), .Z(n59) );
  NAND U187 ( .A(n57), .B(n59), .Z(n495) );
  NAND U188 ( .A(n97), .B(n96), .Z(n60) );
  NANDN U189 ( .A(n95), .B(n94), .Z(n61) );
  NAND U190 ( .A(n60), .B(n61), .Z(n361) );
  NAND U191 ( .A(n502), .B(n500), .Z(n62) );
  XOR U192 ( .A(n500), .B(n502), .Z(n63) );
  NANDN U193 ( .A(n501), .B(n63), .Z(n64) );
  NAND U194 ( .A(n62), .B(n64), .Z(n570) );
  NAND U195 ( .A(n339), .B(n340), .Z(n65) );
  XOR U196 ( .A(n340), .B(n339), .Z(n66) );
  NANDN U197 ( .A(n341), .B(n66), .Z(n67) );
  NAND U198 ( .A(n65), .B(n67), .Z(n367) );
  NAND U199 ( .A(n493), .B(n491), .Z(n68) );
  XOR U200 ( .A(n491), .B(n493), .Z(n69) );
  NANDN U201 ( .A(n492), .B(n69), .Z(n70) );
  NAND U202 ( .A(n68), .B(n70), .Z(n583) );
  NAND U203 ( .A(n555), .B(n554), .Z(n71) );
  XOR U204 ( .A(n554), .B(n555), .Z(n72) );
  NAND U205 ( .A(n72), .B(n553), .Z(n73) );
  NAND U206 ( .A(n71), .B(n73), .Z(n596) );
  NAND U207 ( .A(n603), .B(n602), .Z(n74) );
  NANDN U208 ( .A(n603), .B(n604), .Z(n75) );
  NANDN U209 ( .A(n605), .B(n75), .Z(n76) );
  NAND U210 ( .A(n74), .B(n76), .Z(n608) );
  XNOR U211 ( .A(x[78]), .B(y[78]), .Z(n256) );
  XNOR U212 ( .A(x[82]), .B(y[82]), .Z(n254) );
  XNOR U213 ( .A(x[80]), .B(y[80]), .Z(n253) );
  XNOR U214 ( .A(n254), .B(n253), .Z(n255) );
  XNOR U215 ( .A(n256), .B(n255), .Z(n182) );
  XNOR U216 ( .A(x[84]), .B(y[84]), .Z(n322) );
  XNOR U217 ( .A(x[88]), .B(y[88]), .Z(n320) );
  XNOR U218 ( .A(x[86]), .B(y[86]), .Z(n319) );
  XNOR U219 ( .A(n320), .B(n319), .Z(n321) );
  XNOR U220 ( .A(n322), .B(n321), .Z(n180) );
  XNOR U221 ( .A(x[90]), .B(y[90]), .Z(n238) );
  XNOR U222 ( .A(x[92]), .B(y[92]), .Z(n236) );
  XOR U223 ( .A(oglobal[0]), .B(n236), .Z(n237) );
  XOR U224 ( .A(n238), .B(n237), .Z(n181) );
  XNOR U225 ( .A(n180), .B(n181), .Z(n183) );
  XNOR U226 ( .A(n182), .B(n183), .Z(n335) );
  XNOR U227 ( .A(x[6]), .B(y[6]), .Z(n316) );
  XNOR U228 ( .A(x[10]), .B(y[10]), .Z(n314) );
  XNOR U229 ( .A(x[8]), .B(y[8]), .Z(n313) );
  XNOR U230 ( .A(n314), .B(n313), .Z(n315) );
  XOR U231 ( .A(n316), .B(n315), .Z(n231) );
  XNOR U232 ( .A(x[0]), .B(y[0]), .Z(n248) );
  XNOR U233 ( .A(x[4]), .B(y[4]), .Z(n246) );
  XNOR U234 ( .A(x[2]), .B(y[2]), .Z(n245) );
  XOR U235 ( .A(n246), .B(n245), .Z(n247) );
  XNOR U236 ( .A(n248), .B(n247), .Z(n230) );
  XOR U237 ( .A(n231), .B(n230), .Z(n233) );
  XNOR U238 ( .A(x[5]), .B(y[5]), .Z(n244) );
  XNOR U239 ( .A(x[3]), .B(y[3]), .Z(n242) );
  XNOR U240 ( .A(x[1]), .B(y[1]), .Z(n241) );
  XOR U241 ( .A(n242), .B(n241), .Z(n243) );
  XNOR U242 ( .A(n244), .B(n243), .Z(n232) );
  XOR U243 ( .A(n233), .B(n232), .Z(n333) );
  XNOR U244 ( .A(x[12]), .B(y[12]), .Z(n310) );
  XNOR U245 ( .A(x[16]), .B(y[16]), .Z(n308) );
  XNOR U246 ( .A(x[14]), .B(y[14]), .Z(n307) );
  XNOR U247 ( .A(n308), .B(n307), .Z(n309) );
  XNOR U248 ( .A(n310), .B(n309), .Z(n85) );
  XNOR U249 ( .A(x[18]), .B(y[18]), .Z(n268) );
  XNOR U250 ( .A(x[20]), .B(y[20]), .Z(n266) );
  XNOR U251 ( .A(x[22]), .B(y[22]), .Z(n265) );
  XNOR U252 ( .A(n266), .B(n265), .Z(n267) );
  XNOR U253 ( .A(n268), .B(n267), .Z(n83) );
  XNOR U254 ( .A(x[24]), .B(y[24]), .Z(n262) );
  XNOR U255 ( .A(x[28]), .B(y[28]), .Z(n260) );
  XNOR U256 ( .A(x[26]), .B(y[26]), .Z(n259) );
  XNOR U257 ( .A(n260), .B(n259), .Z(n261) );
  XOR U258 ( .A(n262), .B(n261), .Z(n84) );
  XNOR U259 ( .A(n83), .B(n84), .Z(n86) );
  XNOR U260 ( .A(n85), .B(n86), .Z(n334) );
  XNOR U261 ( .A(n333), .B(n334), .Z(n336) );
  XNOR U262 ( .A(n335), .B(n336), .Z(n349) );
  XNOR U263 ( .A(x[61]), .B(y[61]), .Z(n129) );
  XNOR U264 ( .A(x[97]), .B(y[97]), .Z(n127) );
  XNOR U265 ( .A(x[59]), .B(y[59]), .Z(n126) );
  XNOR U266 ( .A(n127), .B(n126), .Z(n128) );
  XNOR U267 ( .A(n129), .B(n128), .Z(n251) );
  XNOR U268 ( .A(x[77]), .B(y[77]), .Z(n160) );
  XNOR U269 ( .A(x[89]), .B(y[89]), .Z(n158) );
  XNOR U270 ( .A(x[75]), .B(y[75]), .Z(n157) );
  XNOR U271 ( .A(n158), .B(n157), .Z(n159) );
  XNOR U272 ( .A(n160), .B(n159), .Z(n141) );
  XNOR U273 ( .A(x[85]), .B(y[85]), .Z(n139) );
  XNOR U274 ( .A(x[83]), .B(y[83]), .Z(n138) );
  XNOR U275 ( .A(n139), .B(n138), .Z(n140) );
  XOR U276 ( .A(n141), .B(n140), .Z(n250) );
  XNOR U277 ( .A(x[69]), .B(y[69]), .Z(n147) );
  XNOR U278 ( .A(x[93]), .B(y[93]), .Z(n145) );
  XNOR U279 ( .A(x[67]), .B(y[67]), .Z(n144) );
  XNOR U280 ( .A(n145), .B(n144), .Z(n146) );
  XOR U281 ( .A(n147), .B(n146), .Z(n249) );
  XNOR U282 ( .A(n250), .B(n249), .Z(n77) );
  XNOR U283 ( .A(n251), .B(n77), .Z(n95) );
  XNOR U284 ( .A(x[81]), .B(y[81]), .Z(n135) );
  XNOR U285 ( .A(x[87]), .B(y[87]), .Z(n133) );
  XNOR U286 ( .A(x[79]), .B(y[79]), .Z(n132) );
  XNOR U287 ( .A(n133), .B(n132), .Z(n134) );
  XOR U288 ( .A(n135), .B(n134), .Z(n210) );
  XNOR U289 ( .A(x[73]), .B(y[73]), .Z(n154) );
  XNOR U290 ( .A(x[91]), .B(y[91]), .Z(n152) );
  XNOR U291 ( .A(x[71]), .B(y[71]), .Z(n151) );
  XNOR U292 ( .A(n152), .B(n151), .Z(n153) );
  XOR U293 ( .A(n154), .B(n153), .Z(n209) );
  XNOR U294 ( .A(x[65]), .B(y[65]), .Z(n117) );
  XNOR U295 ( .A(x[95]), .B(y[95]), .Z(n115) );
  XNOR U296 ( .A(x[63]), .B(y[63]), .Z(n114) );
  XNOR U297 ( .A(n115), .B(n114), .Z(n116) );
  XNOR U298 ( .A(n117), .B(n116), .Z(n208) );
  XOR U299 ( .A(n209), .B(n208), .Z(n78) );
  XNOR U300 ( .A(n210), .B(n78), .Z(n94) );
  XNOR U301 ( .A(n95), .B(n94), .Z(n96) );
  XNOR U302 ( .A(x[30]), .B(y[30]), .Z(n286) );
  XNOR U303 ( .A(x[34]), .B(y[34]), .Z(n284) );
  XNOR U304 ( .A(x[32]), .B(y[32]), .Z(n283) );
  XOR U305 ( .A(n284), .B(n283), .Z(n285) );
  XNOR U306 ( .A(n286), .B(n285), .Z(n186) );
  XNOR U307 ( .A(x[42]), .B(y[42]), .Z(n220) );
  XNOR U308 ( .A(x[46]), .B(y[46]), .Z(n218) );
  XNOR U309 ( .A(x[44]), .B(y[44]), .Z(n217) );
  XOR U310 ( .A(n218), .B(n217), .Z(n219) );
  XNOR U311 ( .A(n220), .B(n219), .Z(n184) );
  XNOR U312 ( .A(x[36]), .B(y[36]), .Z(n292) );
  XNOR U313 ( .A(x[40]), .B(y[40]), .Z(n290) );
  XNOR U314 ( .A(x[38]), .B(y[38]), .Z(n289) );
  XNOR U315 ( .A(n290), .B(n289), .Z(n291) );
  XOR U316 ( .A(n292), .B(n291), .Z(n185) );
  XNOR U317 ( .A(n184), .B(n185), .Z(n187) );
  XNOR U318 ( .A(n186), .B(n187), .Z(n343) );
  XNOR U319 ( .A(x[72]), .B(y[72]), .Z(n298) );
  XNOR U320 ( .A(x[76]), .B(y[76]), .Z(n296) );
  XNOR U321 ( .A(x[74]), .B(y[74]), .Z(n295) );
  XOR U322 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U323 ( .A(n298), .B(n297), .Z(n89) );
  XNOR U324 ( .A(x[66]), .B(y[66]), .Z(n226) );
  XNOR U325 ( .A(x[68]), .B(y[68]), .Z(n224) );
  XNOR U326 ( .A(x[70]), .B(y[70]), .Z(n223) );
  XOR U327 ( .A(n224), .B(n223), .Z(n225) );
  XNOR U328 ( .A(n226), .B(n225), .Z(n88) );
  XNOR U329 ( .A(x[94]), .B(y[94]), .Z(n113) );
  XNOR U330 ( .A(x[98]), .B(y[98]), .Z(n111) );
  XNOR U331 ( .A(x[96]), .B(y[96]), .Z(n110) );
  XOR U332 ( .A(n111), .B(n110), .Z(n112) );
  XOR U333 ( .A(n113), .B(n112), .Z(n87) );
  XOR U334 ( .A(n88), .B(n87), .Z(n79) );
  XNOR U335 ( .A(n89), .B(n79), .Z(n342) );
  XNOR U336 ( .A(n343), .B(n342), .Z(n345) );
  XNOR U337 ( .A(x[48]), .B(y[48]), .Z(n274) );
  XNOR U338 ( .A(x[50]), .B(y[50]), .Z(n272) );
  XNOR U339 ( .A(x[52]), .B(y[52]), .Z(n271) );
  XNOR U340 ( .A(n272), .B(n271), .Z(n273) );
  XNOR U341 ( .A(n274), .B(n273), .Z(n92) );
  XNOR U342 ( .A(x[60]), .B(y[60]), .Z(n214) );
  XNOR U343 ( .A(x[62]), .B(y[62]), .Z(n212) );
  XNOR U344 ( .A(x[64]), .B(y[64]), .Z(n211) );
  XNOR U345 ( .A(n212), .B(n211), .Z(n213) );
  XNOR U346 ( .A(n214), .B(n213), .Z(n90) );
  XNOR U347 ( .A(x[54]), .B(y[54]), .Z(n280) );
  XNOR U348 ( .A(x[58]), .B(y[58]), .Z(n278) );
  XNOR U349 ( .A(x[56]), .B(y[56]), .Z(n277) );
  XNOR U350 ( .A(n278), .B(n277), .Z(n279) );
  XOR U351 ( .A(n280), .B(n279), .Z(n91) );
  XNOR U352 ( .A(n90), .B(n91), .Z(n93) );
  XNOR U353 ( .A(n92), .B(n93), .Z(n344) );
  XNOR U354 ( .A(n345), .B(n344), .Z(n97) );
  XOR U355 ( .A(n96), .B(n97), .Z(n350) );
  XOR U356 ( .A(n349), .B(n350), .Z(n351) );
  XNOR U357 ( .A(x[35]), .B(y[35]), .Z(n193) );
  XNOR U358 ( .A(x[33]), .B(y[33]), .Z(n191) );
  XNOR U359 ( .A(x[31]), .B(y[31]), .Z(n190) );
  XNOR U360 ( .A(n191), .B(n190), .Z(n192) );
  XOR U361 ( .A(n193), .B(n192), .Z(n326) );
  IV U362 ( .A(n326), .Z(n325) );
  XNOR U363 ( .A(x[41]), .B(y[41]), .Z(n173) );
  XNOR U364 ( .A(x[39]), .B(y[39]), .Z(n171) );
  XNOR U365 ( .A(x[37]), .B(y[37]), .Z(n170) );
  XNOR U366 ( .A(n171), .B(n170), .Z(n172) );
  XNOR U367 ( .A(n173), .B(n172), .Z(n329) );
  XNOR U368 ( .A(x[29]), .B(y[29]), .Z(n205) );
  XNOR U369 ( .A(x[25]), .B(y[25]), .Z(n203) );
  XNOR U370 ( .A(x[27]), .B(y[27]), .Z(n202) );
  XNOR U371 ( .A(n203), .B(n202), .Z(n204) );
  XNOR U372 ( .A(n205), .B(n204), .Z(n327) );
  XNOR U373 ( .A(n329), .B(n327), .Z(n80) );
  XNOR U374 ( .A(n325), .B(n80), .Z(n341) );
  XNOR U375 ( .A(x[23]), .B(y[23]), .Z(n199) );
  XNOR U376 ( .A(x[21]), .B(y[21]), .Z(n197) );
  XNOR U377 ( .A(x[19]), .B(y[19]), .Z(n196) );
  XNOR U378 ( .A(n197), .B(n196), .Z(n198) );
  XNOR U379 ( .A(n199), .B(n198), .Z(n305) );
  XNOR U380 ( .A(x[17]), .B(y[17]), .Z(n101) );
  XNOR U381 ( .A(x[15]), .B(y[15]), .Z(n99) );
  XNOR U382 ( .A(x[13]), .B(y[13]), .Z(n98) );
  XNOR U383 ( .A(n99), .B(n98), .Z(n100) );
  XNOR U384 ( .A(n101), .B(n100), .Z(n303) );
  XNOR U385 ( .A(x[11]), .B(y[11]), .Z(n107) );
  XNOR U386 ( .A(x[9]), .B(y[9]), .Z(n105) );
  XNOR U387 ( .A(x[7]), .B(y[7]), .Z(n104) );
  XNOR U388 ( .A(n105), .B(n104), .Z(n106) );
  XOR U389 ( .A(n107), .B(n106), .Z(n304) );
  XNOR U390 ( .A(n303), .B(n304), .Z(n306) );
  XNOR U391 ( .A(n305), .B(n306), .Z(n340) );
  XNOR U392 ( .A(x[57]), .B(y[57]), .Z(n123) );
  XNOR U393 ( .A(x[99]), .B(y[99]), .Z(n121) );
  XNOR U394 ( .A(x[55]), .B(y[55]), .Z(n120) );
  XNOR U395 ( .A(n121), .B(n120), .Z(n122) );
  XOR U396 ( .A(n123), .B(n122), .Z(n302) );
  XNOR U397 ( .A(x[53]), .B(y[53]), .Z(n167) );
  XNOR U398 ( .A(x[51]), .B(y[51]), .Z(n165) );
  XNOR U399 ( .A(x[49]), .B(y[49]), .Z(n164) );
  XOR U400 ( .A(n165), .B(n164), .Z(n166) );
  XNOR U401 ( .A(n167), .B(n166), .Z(n301) );
  XNOR U402 ( .A(x[47]), .B(y[47]), .Z(n179) );
  XNOR U403 ( .A(x[45]), .B(y[45]), .Z(n177) );
  XNOR U404 ( .A(x[43]), .B(y[43]), .Z(n176) );
  XOR U405 ( .A(n177), .B(n176), .Z(n178) );
  XOR U406 ( .A(n179), .B(n178), .Z(n300) );
  XOR U407 ( .A(n301), .B(n300), .Z(n81) );
  XNOR U408 ( .A(n302), .B(n81), .Z(n339) );
  XOR U409 ( .A(n340), .B(n339), .Z(n82) );
  XNOR U410 ( .A(n341), .B(n82), .Z(n352) );
  XOR U411 ( .A(n351), .B(n352), .Z(o[0]) );
  XNOR U412 ( .A(n413), .B(n414), .Z(n415) );
  XNOR U413 ( .A(n416), .B(n415), .Z(n364) );
  OR U414 ( .A(n99), .B(n98), .Z(n103) );
  OR U415 ( .A(n101), .B(n100), .Z(n102) );
  NAND U416 ( .A(n103), .B(n102), .Z(n469) );
  OR U417 ( .A(n105), .B(n104), .Z(n109) );
  OR U418 ( .A(n107), .B(n106), .Z(n108) );
  NAND U419 ( .A(n109), .B(n108), .Z(n468) );
  XNOR U420 ( .A(n469), .B(n468), .Z(n471) );
  XNOR U421 ( .A(n471), .B(n470), .Z(n391) );
  OR U422 ( .A(n115), .B(n114), .Z(n119) );
  OR U423 ( .A(n117), .B(n116), .Z(n118) );
  NAND U424 ( .A(n119), .B(n118), .Z(n463) );
  OR U425 ( .A(n121), .B(n120), .Z(n125) );
  OR U426 ( .A(n123), .B(n122), .Z(n124) );
  NAND U427 ( .A(n125), .B(n124), .Z(n462) );
  XNOR U428 ( .A(n463), .B(n462), .Z(n465) );
  OR U429 ( .A(n127), .B(n126), .Z(n131) );
  OR U430 ( .A(n129), .B(n128), .Z(n130) );
  NAND U431 ( .A(n131), .B(n130), .Z(n464) );
  XOR U432 ( .A(n465), .B(n464), .Z(n390) );
  XNOR U433 ( .A(n391), .B(n390), .Z(n393) );
  OR U434 ( .A(n133), .B(n132), .Z(n137) );
  OR U435 ( .A(n135), .B(n134), .Z(n136) );
  AND U436 ( .A(n137), .B(n136), .Z(n460) );
  OR U437 ( .A(n139), .B(n138), .Z(n143) );
  OR U438 ( .A(n141), .B(n140), .Z(n142) );
  NAND U439 ( .A(n143), .B(n142), .Z(n461) );
  OR U440 ( .A(n145), .B(n144), .Z(n149) );
  OR U441 ( .A(n147), .B(n146), .Z(n148) );
  AND U442 ( .A(n149), .B(n148), .Z(n459) );
  XOR U443 ( .A(n461), .B(n459), .Z(n150) );
  XNOR U444 ( .A(n460), .B(n150), .Z(n392) );
  XOR U445 ( .A(n393), .B(n392), .Z(n362) );
  XNOR U446 ( .A(n361), .B(n362), .Z(n363) );
  XNOR U447 ( .A(n364), .B(n363), .Z(n379) );
  OR U448 ( .A(n152), .B(n151), .Z(n156) );
  OR U449 ( .A(n154), .B(n153), .Z(n155) );
  AND U450 ( .A(n156), .B(n155), .Z(n430) );
  IV U451 ( .A(n430), .Z(n431) );
  OR U452 ( .A(n158), .B(n157), .Z(n162) );
  OR U453 ( .A(n160), .B(n159), .Z(n161) );
  AND U454 ( .A(n162), .B(n161), .Z(n432) );
  IV U455 ( .A(n432), .Z(n429) );
  XOR U456 ( .A(n429), .B(oglobal[1]), .Z(n163) );
  XNOR U457 ( .A(n431), .B(n163), .Z(n480) );
  OR U458 ( .A(n165), .B(n164), .Z(n169) );
  NANDN U459 ( .A(n167), .B(n166), .Z(n168) );
  NAND U460 ( .A(n169), .B(n168), .Z(n438) );
  OR U461 ( .A(n171), .B(n170), .Z(n175) );
  OR U462 ( .A(n173), .B(n172), .Z(n174) );
  NAND U463 ( .A(n175), .B(n174), .Z(n437) );
  XNOR U464 ( .A(n438), .B(n437), .Z(n440) );
  XNOR U465 ( .A(n440), .B(n439), .Z(n478) );
  XNOR U466 ( .A(n478), .B(n477), .Z(n479) );
  XOR U467 ( .A(n480), .B(n479), .Z(n383) );
  OR U468 ( .A(n185), .B(n184), .Z(n189) );
  OR U469 ( .A(n187), .B(n186), .Z(n188) );
  NAND U470 ( .A(n189), .B(n188), .Z(n384) );
  XNOR U471 ( .A(n383), .B(n384), .Z(n386) );
  OR U472 ( .A(n191), .B(n190), .Z(n195) );
  OR U473 ( .A(n193), .B(n192), .Z(n194) );
  NAND U474 ( .A(n195), .B(n194), .Z(n447) );
  OR U475 ( .A(n197), .B(n196), .Z(n201) );
  OR U476 ( .A(n199), .B(n198), .Z(n200) );
  NAND U477 ( .A(n201), .B(n200), .Z(n446) );
  XNOR U478 ( .A(n447), .B(n446), .Z(n449) );
  OR U479 ( .A(n203), .B(n202), .Z(n207) );
  OR U480 ( .A(n205), .B(n204), .Z(n206) );
  NAND U481 ( .A(n207), .B(n206), .Z(n448) );
  XNOR U482 ( .A(n449), .B(n448), .Z(n476) );
  OR U483 ( .A(n212), .B(n211), .Z(n216) );
  OR U484 ( .A(n214), .B(n213), .Z(n215) );
  NAND U485 ( .A(n216), .B(n215), .Z(n395) );
  OR U486 ( .A(n218), .B(n217), .Z(n222) );
  NANDN U487 ( .A(n220), .B(n219), .Z(n221) );
  NAND U488 ( .A(n222), .B(n221), .Z(n394) );
  XNOR U489 ( .A(n395), .B(n394), .Z(n397) );
  OR U490 ( .A(n224), .B(n223), .Z(n228) );
  NANDN U491 ( .A(n226), .B(n225), .Z(n227) );
  NAND U492 ( .A(n228), .B(n227), .Z(n396) );
  XNOR U493 ( .A(n397), .B(n396), .Z(n475) );
  XOR U494 ( .A(n474), .B(n475), .Z(n229) );
  XNOR U495 ( .A(n476), .B(n229), .Z(n385) );
  XNOR U496 ( .A(n386), .B(n385), .Z(n377) );
  NAND U497 ( .A(n231), .B(n230), .Z(n235) );
  NAND U498 ( .A(n233), .B(n232), .Z(n234) );
  NAND U499 ( .A(n235), .B(n234), .Z(n389) );
  NANDN U500 ( .A(n236), .B(oglobal[0]), .Z(n240) );
  OR U501 ( .A(n238), .B(n237), .Z(n239) );
  AND U502 ( .A(n240), .B(n239), .Z(n426) );
  XNOR U503 ( .A(n423), .B(n424), .Z(n425) );
  XNOR U504 ( .A(n426), .B(n425), .Z(n387) );
  XOR U505 ( .A(n387), .B(n388), .Z(n252) );
  XOR U506 ( .A(n389), .B(n252), .Z(n373) );
  OR U507 ( .A(n254), .B(n253), .Z(n258) );
  OR U508 ( .A(n256), .B(n255), .Z(n257) );
  NAND U509 ( .A(n258), .B(n257), .Z(n408) );
  OR U510 ( .A(n260), .B(n259), .Z(n264) );
  OR U511 ( .A(n262), .B(n261), .Z(n263) );
  AND U512 ( .A(n264), .B(n263), .Z(n406) );
  OR U513 ( .A(n266), .B(n265), .Z(n270) );
  OR U514 ( .A(n268), .B(n267), .Z(n269) );
  AND U515 ( .A(n270), .B(n269), .Z(n407) );
  XNOR U516 ( .A(n406), .B(n407), .Z(n409) );
  XOR U517 ( .A(n408), .B(n409), .Z(n485) );
  OR U518 ( .A(n272), .B(n271), .Z(n276) );
  OR U519 ( .A(n274), .B(n273), .Z(n275) );
  NAND U520 ( .A(n276), .B(n275), .Z(n401) );
  OR U521 ( .A(n278), .B(n277), .Z(n282) );
  OR U522 ( .A(n280), .B(n279), .Z(n281) );
  NAND U523 ( .A(n282), .B(n281), .Z(n400) );
  XNOR U524 ( .A(n401), .B(n400), .Z(n403) );
  OR U525 ( .A(n284), .B(n283), .Z(n288) );
  NANDN U526 ( .A(n286), .B(n285), .Z(n287) );
  AND U527 ( .A(n288), .B(n287), .Z(n443) );
  OR U528 ( .A(n290), .B(n289), .Z(n294) );
  OR U529 ( .A(n292), .B(n291), .Z(n293) );
  NAND U530 ( .A(n294), .B(n293), .Z(n445) );
  XNOR U531 ( .A(n445), .B(n444), .Z(n299) );
  XOR U532 ( .A(n443), .B(n299), .Z(n402) );
  XNOR U533 ( .A(n403), .B(n402), .Z(n484) );
  XOR U534 ( .A(n484), .B(n483), .Z(n486) );
  XOR U535 ( .A(n485), .B(n486), .Z(n370) );
  OR U536 ( .A(n308), .B(n307), .Z(n312) );
  OR U537 ( .A(n310), .B(n309), .Z(n311) );
  NAND U538 ( .A(n312), .B(n311), .Z(n418) );
  OR U539 ( .A(n314), .B(n313), .Z(n318) );
  OR U540 ( .A(n316), .B(n315), .Z(n317) );
  NAND U541 ( .A(n318), .B(n317), .Z(n417) );
  XNOR U542 ( .A(n418), .B(n417), .Z(n420) );
  OR U543 ( .A(n320), .B(n319), .Z(n324) );
  OR U544 ( .A(n322), .B(n321), .Z(n323) );
  NAND U545 ( .A(n324), .B(n323), .Z(n419) );
  XNOR U546 ( .A(n420), .B(n419), .Z(n454) );
  OR U547 ( .A(n327), .B(n325), .Z(n331) );
  ANDN U548 ( .B(n327), .A(n326), .Z(n328) );
  OR U549 ( .A(n329), .B(n328), .Z(n330) );
  AND U550 ( .A(n331), .B(n330), .Z(n453) );
  IV U551 ( .A(n453), .Z(n452) );
  XNOR U552 ( .A(n454), .B(n452), .Z(n332) );
  XNOR U553 ( .A(n455), .B(n332), .Z(n371) );
  XNOR U554 ( .A(n370), .B(n371), .Z(n372) );
  XOR U555 ( .A(n373), .B(n372), .Z(n378) );
  XOR U556 ( .A(n377), .B(n378), .Z(n380) );
  XOR U557 ( .A(n379), .B(n380), .Z(n355) );
  NAND U558 ( .A(n334), .B(n333), .Z(n338) );
  NANDN U559 ( .A(n336), .B(n335), .Z(n337) );
  AND U560 ( .A(n338), .B(n337), .Z(n369) );
  NAND U561 ( .A(n343), .B(n342), .Z(n347) );
  NANDN U562 ( .A(n345), .B(n344), .Z(n346) );
  AND U563 ( .A(n347), .B(n346), .Z(n368) );
  XOR U564 ( .A(n367), .B(n368), .Z(n348) );
  XOR U565 ( .A(n369), .B(n348), .Z(n356) );
  XOR U566 ( .A(n355), .B(n356), .Z(n357) );
  NAND U567 ( .A(n350), .B(n349), .Z(n354) );
  NAND U568 ( .A(n352), .B(n351), .Z(n353) );
  AND U569 ( .A(n354), .B(n353), .Z(n358) );
  XNOR U570 ( .A(n357), .B(n358), .Z(o[1]) );
  NAND U571 ( .A(n356), .B(n355), .Z(n360) );
  NANDN U572 ( .A(n358), .B(n357), .Z(n359) );
  NAND U573 ( .A(n360), .B(n359), .Z(n547) );
  NANDN U574 ( .A(n362), .B(n361), .Z(n366) );
  NANDN U575 ( .A(n364), .B(n363), .Z(n365) );
  AND U576 ( .A(n366), .B(n365), .Z(n545) );
  NANDN U577 ( .A(n371), .B(n370), .Z(n375) );
  NAND U578 ( .A(n373), .B(n372), .Z(n374) );
  AND U579 ( .A(n375), .B(n374), .Z(n544) );
  XOR U580 ( .A(n543), .B(n544), .Z(n376) );
  XNOR U581 ( .A(n545), .B(n376), .Z(n548) );
  XNOR U582 ( .A(n547), .B(n548), .Z(n549) );
  NAND U583 ( .A(n378), .B(n377), .Z(n382) );
  NAND U584 ( .A(n380), .B(n379), .Z(n381) );
  NAND U585 ( .A(n382), .B(n381), .Z(n491) );
  XNOR U586 ( .A(n532), .B(n531), .Z(n533) );
  OR U587 ( .A(n395), .B(n394), .Z(n399) );
  OR U588 ( .A(n397), .B(n396), .Z(n398) );
  AND U589 ( .A(n399), .B(n398), .Z(n501) );
  OR U590 ( .A(n401), .B(n400), .Z(n405) );
  OR U591 ( .A(n403), .B(n402), .Z(n404) );
  NAND U592 ( .A(n405), .B(n404), .Z(n502) );
  OR U593 ( .A(n407), .B(n406), .Z(n411) );
  NANDN U594 ( .A(n409), .B(n408), .Z(n410) );
  AND U595 ( .A(n411), .B(n410), .Z(n500) );
  XOR U596 ( .A(n502), .B(n500), .Z(n412) );
  XNOR U597 ( .A(n501), .B(n412), .Z(n538) );
  IV U598 ( .A(n535), .Z(n537) );
  OR U599 ( .A(n418), .B(n417), .Z(n422) );
  OR U600 ( .A(n420), .B(n419), .Z(n421) );
  AND U601 ( .A(n422), .B(n421), .Z(n512) );
  OR U602 ( .A(n424), .B(n423), .Z(n428) );
  OR U603 ( .A(n426), .B(n425), .Z(n427) );
  AND U604 ( .A(n428), .B(n427), .Z(n515) );
  XNOR U605 ( .A(oglobal[2]), .B(n515), .Z(n509) );
  NANDN U606 ( .A(n430), .B(n429), .Z(n435) );
  ANDN U607 ( .B(n432), .A(n431), .Z(n433) );
  NANDN U608 ( .A(n433), .B(oglobal[1]), .Z(n434) );
  NAND U609 ( .A(n435), .B(n434), .Z(n510) );
  XNOR U610 ( .A(n509), .B(n510), .Z(n511) );
  XOR U611 ( .A(n537), .B(n536), .Z(n436) );
  XOR U612 ( .A(n538), .B(n436), .Z(n534) );
  XOR U613 ( .A(n533), .B(n534), .Z(n524) );
  OR U614 ( .A(n438), .B(n437), .Z(n442) );
  OR U615 ( .A(n440), .B(n439), .Z(n441) );
  NAND U616 ( .A(n442), .B(n441), .Z(n506) );
  OR U617 ( .A(n447), .B(n446), .Z(n451) );
  OR U618 ( .A(n449), .B(n448), .Z(n450) );
  AND U619 ( .A(n451), .B(n450), .Z(n504) );
  XNOR U620 ( .A(n503), .B(n504), .Z(n505) );
  XNOR U621 ( .A(n506), .B(n505), .Z(n518) );
  OR U622 ( .A(n454), .B(n452), .Z(n458) );
  ANDN U623 ( .B(n454), .A(n453), .Z(n456) );
  NANDN U624 ( .A(n456), .B(n455), .Z(n457) );
  NAND U625 ( .A(n458), .B(n457), .Z(n516) );
  OR U626 ( .A(n463), .B(n462), .Z(n467) );
  OR U627 ( .A(n465), .B(n464), .Z(n466) );
  AND U628 ( .A(n467), .B(n466), .Z(n494) );
  XNOR U629 ( .A(n495), .B(n494), .Z(n496) );
  OR U630 ( .A(n469), .B(n468), .Z(n473) );
  OR U631 ( .A(n471), .B(n470), .Z(n472) );
  NAND U632 ( .A(n473), .B(n472), .Z(n497) );
  XNOR U633 ( .A(n496), .B(n497), .Z(n517) );
  XOR U634 ( .A(n516), .B(n517), .Z(n519) );
  XOR U635 ( .A(n518), .B(n519), .Z(n523) );
  NANDN U636 ( .A(n478), .B(n477), .Z(n482) );
  NAND U637 ( .A(n480), .B(n479), .Z(n481) );
  AND U638 ( .A(n482), .B(n481), .Z(n526) );
  XOR U639 ( .A(n525), .B(n526), .Z(n528) );
  NANDN U640 ( .A(n484), .B(n483), .Z(n488) );
  NANDN U641 ( .A(n486), .B(n485), .Z(n487) );
  AND U642 ( .A(n488), .B(n487), .Z(n527) );
  XOR U643 ( .A(n528), .B(n527), .Z(n522) );
  XNOR U644 ( .A(n523), .B(n522), .Z(n489) );
  XOR U645 ( .A(n524), .B(n489), .Z(n493) );
  XOR U646 ( .A(n492), .B(n493), .Z(n490) );
  XNOR U647 ( .A(n491), .B(n490), .Z(n550) );
  XOR U648 ( .A(n549), .B(n550), .Z(o[2]) );
  NANDN U649 ( .A(n495), .B(n494), .Z(n499) );
  NANDN U650 ( .A(n497), .B(n496), .Z(n498) );
  NAND U651 ( .A(n499), .B(n498), .Z(n571) );
  XOR U652 ( .A(n571), .B(n570), .Z(n573) );
  NANDN U653 ( .A(n504), .B(n503), .Z(n508) );
  NAND U654 ( .A(n506), .B(n505), .Z(n507) );
  AND U655 ( .A(n508), .B(n507), .Z(n576) );
  OR U656 ( .A(n510), .B(n509), .Z(n514) );
  OR U657 ( .A(n512), .B(n511), .Z(n513) );
  AND U658 ( .A(n514), .B(n513), .Z(n577) );
  XNOR U659 ( .A(n576), .B(n577), .Z(n578) );
  NANDN U660 ( .A(n515), .B(oglobal[2]), .Z(n569) );
  XNOR U661 ( .A(n569), .B(oglobal[3]), .Z(n579) );
  XOR U662 ( .A(n573), .B(n572), .Z(n559) );
  NANDN U663 ( .A(n517), .B(n516), .Z(n521) );
  OR U664 ( .A(n519), .B(n518), .Z(n520) );
  AND U665 ( .A(n521), .B(n520), .Z(n557) );
  XOR U666 ( .A(n557), .B(n556), .Z(n558) );
  XNOR U667 ( .A(n559), .B(n558), .Z(n555) );
  NANDN U668 ( .A(n526), .B(n525), .Z(n530) );
  OR U669 ( .A(n528), .B(n527), .Z(n529) );
  AND U670 ( .A(n530), .B(n529), .Z(n564) );
  NANDN U671 ( .A(n535), .B(n536), .Z(n541) );
  NOR U672 ( .A(n537), .B(n536), .Z(n539) );
  NANDN U673 ( .A(n539), .B(n538), .Z(n540) );
  AND U674 ( .A(n541), .B(n540), .Z(n562) );
  IV U675 ( .A(n562), .Z(n563) );
  XNOR U676 ( .A(n565), .B(n563), .Z(n542) );
  XNOR U677 ( .A(n564), .B(n542), .Z(n554) );
  XOR U678 ( .A(n554), .B(n553), .Z(n546) );
  XOR U679 ( .A(n555), .B(n546), .Z(n584) );
  XOR U680 ( .A(n583), .B(n584), .Z(n585) );
  NANDN U681 ( .A(n548), .B(n547), .Z(n552) );
  NAND U682 ( .A(n550), .B(n549), .Z(n551) );
  AND U683 ( .A(n552), .B(n551), .Z(n586) );
  XNOR U684 ( .A(n585), .B(n586), .Z(o[3]) );
  NANDN U685 ( .A(n557), .B(n556), .Z(n561) );
  OR U686 ( .A(n559), .B(n558), .Z(n560) );
  NAND U687 ( .A(n561), .B(n560), .Z(n605) );
  OR U688 ( .A(n564), .B(n562), .Z(n568) );
  ANDN U689 ( .B(n564), .A(n563), .Z(n566) );
  NANDN U690 ( .A(n566), .B(n565), .Z(n567) );
  AND U691 ( .A(n568), .B(n567), .Z(n602) );
  IV U692 ( .A(n602), .Z(n604) );
  NANDN U693 ( .A(n569), .B(oglobal[3]), .Z(n589) );
  XOR U694 ( .A(oglobal[4]), .B(n589), .Z(n592) );
  NANDN U695 ( .A(n571), .B(n570), .Z(n575) );
  NANDN U696 ( .A(n573), .B(n572), .Z(n574) );
  AND U697 ( .A(n575), .B(n574), .Z(n591) );
  OR U698 ( .A(n577), .B(n576), .Z(n581) );
  OR U699 ( .A(n579), .B(n578), .Z(n580) );
  AND U700 ( .A(n581), .B(n580), .Z(n590) );
  XNOR U701 ( .A(n591), .B(n590), .Z(n593) );
  XOR U702 ( .A(n592), .B(n593), .Z(n603) );
  XOR U703 ( .A(n604), .B(n603), .Z(n582) );
  XNOR U704 ( .A(n605), .B(n582), .Z(n597) );
  XOR U705 ( .A(n596), .B(n597), .Z(n599) );
  NAND U706 ( .A(n584), .B(n583), .Z(n588) );
  NANDN U707 ( .A(n586), .B(n585), .Z(n587) );
  AND U708 ( .A(n588), .B(n587), .Z(n598) );
  XOR U709 ( .A(n599), .B(n598), .Z(o[4]) );
  NANDN U710 ( .A(n589), .B(oglobal[4]), .Z(n612) );
  XOR U711 ( .A(oglobal[5]), .B(n612), .Z(n614) );
  OR U712 ( .A(n591), .B(n590), .Z(n595) );
  NANDN U713 ( .A(n593), .B(n592), .Z(n594) );
  NAND U714 ( .A(n595), .B(n594), .Z(n613) );
  XOR U715 ( .A(n614), .B(n613), .Z(n607) );
  NANDN U716 ( .A(n597), .B(n596), .Z(n601) );
  OR U717 ( .A(n599), .B(n598), .Z(n600) );
  NAND U718 ( .A(n601), .B(n600), .Z(n609) );
  XOR U719 ( .A(n609), .B(n608), .Z(n606) );
  XOR U720 ( .A(n607), .B(n606), .Z(o[5]) );
  NANDN U721 ( .A(n607), .B(n606), .Z(n611) );
  OR U722 ( .A(n609), .B(n608), .Z(n610) );
  AND U723 ( .A(n611), .B(n610), .Z(n617) );
  XNOR U724 ( .A(n617), .B(oglobal[6]), .Z(n619) );
  NANDN U725 ( .A(n612), .B(oglobal[5]), .Z(n616) );
  OR U726 ( .A(n614), .B(n613), .Z(n615) );
  AND U727 ( .A(n616), .B(n615), .Z(n618) );
  XOR U728 ( .A(n619), .B(n618), .Z(o[6]) );
  NAND U729 ( .A(n617), .B(oglobal[6]), .Z(n621) );
  OR U730 ( .A(n619), .B(n618), .Z(n620) );
  AND U731 ( .A(n621), .B(n620), .Z(n622) );
  XNOR U732 ( .A(oglobal[7]), .B(n622), .Z(o[7]) );
  NANDN U733 ( .A(n622), .B(oglobal[7]), .Z(n623) );
  XNOR U734 ( .A(n623), .B(oglobal[8]), .Z(o[8]) );
  NANDN U735 ( .A(n623), .B(oglobal[8]), .Z(n624) );
  XNOR U736 ( .A(oglobal[9]), .B(n624), .Z(o[9]) );
  NANDN U737 ( .A(n624), .B(oglobal[9]), .Z(n625) );
  XNOR U738 ( .A(oglobal[10]), .B(n625), .Z(o[10]) );
endmodule

