
module hamming_N16000_CC4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;

  XNOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U18 ( .A(B[1]), .B(A[1]), .Z(n18) );
  XOR U19 ( .A(A[13]), .B(n19), .Z(SUM[13]) );
  AND U20 ( .A(A[12]), .B(n20), .Z(n19) );
  XOR U21 ( .A(A[12]), .B(n20), .Z(SUM[12]) );
  NAND U22 ( .A(n21), .B(n22), .Z(n20) );
  NAND U23 ( .A(B[11]), .B(n23), .Z(n22) );
  NANDN U24 ( .A(A[11]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(n24), .B(A[11]), .Z(n21) );
  XOR U26 ( .A(n24), .B(n25), .Z(SUM[11]) );
  XNOR U27 ( .A(B[11]), .B(A[11]), .Z(n25) );
  AND U28 ( .A(n26), .B(n27), .Z(n24) );
  NAND U29 ( .A(B[10]), .B(n28), .Z(n27) );
  NANDN U30 ( .A(A[10]), .B(n29), .Z(n28) );
  NANDN U31 ( .A(n29), .B(A[10]), .Z(n26) );
  XOR U32 ( .A(n29), .B(n30), .Z(SUM[10]) );
  XNOR U33 ( .A(B[10]), .B(A[10]), .Z(n30) );
  AND U34 ( .A(n31), .B(n32), .Z(n29) );
  NAND U35 ( .A(B[9]), .B(n33), .Z(n32) );
  OR U36 ( .A(n1), .B(A[9]), .Z(n33) );
  NAND U37 ( .A(A[9]), .B(n1), .Z(n31) );
  NAND U38 ( .A(n34), .B(n35), .Z(n1) );
  NAND U39 ( .A(B[8]), .B(n36), .Z(n35) );
  NANDN U40 ( .A(A[8]), .B(n3), .Z(n36) );
  NANDN U41 ( .A(n3), .B(A[8]), .Z(n34) );
  AND U42 ( .A(n37), .B(n38), .Z(n3) );
  NAND U43 ( .A(B[7]), .B(n39), .Z(n38) );
  NANDN U44 ( .A(A[7]), .B(n5), .Z(n39) );
  NANDN U45 ( .A(n5), .B(A[7]), .Z(n37) );
  AND U46 ( .A(n40), .B(n41), .Z(n5) );
  NAND U47 ( .A(B[6]), .B(n42), .Z(n41) );
  NANDN U48 ( .A(A[6]), .B(n7), .Z(n42) );
  NANDN U49 ( .A(n7), .B(A[6]), .Z(n40) );
  AND U50 ( .A(n43), .B(n44), .Z(n7) );
  NAND U51 ( .A(B[5]), .B(n45), .Z(n44) );
  NANDN U52 ( .A(A[5]), .B(n9), .Z(n45) );
  NANDN U53 ( .A(n9), .B(A[5]), .Z(n43) );
  AND U54 ( .A(n46), .B(n47), .Z(n9) );
  NAND U55 ( .A(B[4]), .B(n48), .Z(n47) );
  NANDN U56 ( .A(A[4]), .B(n11), .Z(n48) );
  NANDN U57 ( .A(n11), .B(A[4]), .Z(n46) );
  AND U58 ( .A(n49), .B(n50), .Z(n11) );
  NAND U59 ( .A(B[3]), .B(n51), .Z(n50) );
  NANDN U60 ( .A(A[3]), .B(n13), .Z(n51) );
  NANDN U61 ( .A(n13), .B(A[3]), .Z(n49) );
  AND U62 ( .A(n52), .B(n53), .Z(n13) );
  NAND U63 ( .A(B[2]), .B(n54), .Z(n53) );
  NANDN U64 ( .A(A[2]), .B(n15), .Z(n54) );
  NANDN U65 ( .A(n15), .B(A[2]), .Z(n52) );
  AND U66 ( .A(n55), .B(n56), .Z(n15) );
  NAND U67 ( .A(B[1]), .B(n57), .Z(n56) );
  OR U68 ( .A(n17), .B(A[1]), .Z(n57) );
  NAND U69 ( .A(A[1]), .B(n17), .Z(n55) );
  AND U70 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U71 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52;

  IV U1 ( .A(B[11]), .Z(n1) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  XOR U20 ( .A(n20), .B(n1), .Z(SUM[11]) );
  AND U21 ( .A(n21), .B(n22), .Z(n20) );
  NAND U22 ( .A(B[10]), .B(n23), .Z(n22) );
  NANDN U23 ( .A(A[10]), .B(n24), .Z(n23) );
  NANDN U24 ( .A(n24), .B(A[10]), .Z(n21) );
  XOR U25 ( .A(n24), .B(n25), .Z(SUM[10]) );
  XNOR U26 ( .A(B[10]), .B(A[10]), .Z(n25) );
  AND U27 ( .A(n26), .B(n27), .Z(n24) );
  NAND U28 ( .A(B[9]), .B(n28), .Z(n27) );
  OR U29 ( .A(n2), .B(A[9]), .Z(n28) );
  NAND U30 ( .A(A[9]), .B(n2), .Z(n26) );
  NAND U31 ( .A(n29), .B(n30), .Z(n2) );
  NAND U32 ( .A(B[8]), .B(n31), .Z(n30) );
  NANDN U33 ( .A(A[8]), .B(n4), .Z(n31) );
  NANDN U34 ( .A(n4), .B(A[8]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n4) );
  NAND U36 ( .A(B[7]), .B(n34), .Z(n33) );
  NANDN U37 ( .A(A[7]), .B(n6), .Z(n34) );
  NANDN U38 ( .A(n6), .B(A[7]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n6) );
  NAND U40 ( .A(B[6]), .B(n37), .Z(n36) );
  NANDN U41 ( .A(A[6]), .B(n8), .Z(n37) );
  NANDN U42 ( .A(n8), .B(A[6]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n8) );
  NAND U44 ( .A(B[5]), .B(n40), .Z(n39) );
  NANDN U45 ( .A(A[5]), .B(n10), .Z(n40) );
  NANDN U46 ( .A(n10), .B(A[5]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n10) );
  NAND U48 ( .A(B[4]), .B(n43), .Z(n42) );
  NANDN U49 ( .A(A[4]), .B(n12), .Z(n43) );
  NANDN U50 ( .A(n12), .B(A[4]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n12) );
  NAND U52 ( .A(B[3]), .B(n46), .Z(n45) );
  NANDN U53 ( .A(A[3]), .B(n14), .Z(n46) );
  NANDN U54 ( .A(n14), .B(A[3]), .Z(n44) );
  AND U55 ( .A(n47), .B(n48), .Z(n14) );
  NAND U56 ( .A(B[2]), .B(n49), .Z(n48) );
  NANDN U57 ( .A(A[2]), .B(n16), .Z(n49) );
  NANDN U58 ( .A(n16), .B(A[2]), .Z(n47) );
  AND U59 ( .A(n50), .B(n51), .Z(n16) );
  NAND U60 ( .A(B[1]), .B(n52), .Z(n51) );
  OR U61 ( .A(n18), .B(A[1]), .Z(n52) );
  NAND U62 ( .A(A[1]), .B(n18), .Z(n50) );
  AND U63 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U64 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_2 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[11]) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(B[10]), .B(n22), .Z(n21) );
  NANDN U21 ( .A(A[10]), .B(n23), .Z(n22) );
  NANDN U22 ( .A(n23), .B(A[10]), .Z(n20) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[10]) );
  XNOR U24 ( .A(B[10]), .B(A[10]), .Z(n24) );
  AND U25 ( .A(n25), .B(n26), .Z(n23) );
  NAND U26 ( .A(B[9]), .B(n27), .Z(n26) );
  OR U27 ( .A(n2), .B(A[9]), .Z(n27) );
  NAND U28 ( .A(A[9]), .B(n2), .Z(n25) );
  NAND U29 ( .A(n28), .B(n29), .Z(n2) );
  NAND U30 ( .A(B[8]), .B(n30), .Z(n29) );
  NANDN U31 ( .A(A[8]), .B(n4), .Z(n30) );
  NANDN U32 ( .A(n4), .B(A[8]), .Z(n28) );
  AND U33 ( .A(n31), .B(n32), .Z(n4) );
  NAND U34 ( .A(B[7]), .B(n33), .Z(n32) );
  NANDN U35 ( .A(A[7]), .B(n6), .Z(n33) );
  NANDN U36 ( .A(n6), .B(A[7]), .Z(n31) );
  AND U37 ( .A(n34), .B(n35), .Z(n6) );
  NAND U38 ( .A(B[6]), .B(n36), .Z(n35) );
  NANDN U39 ( .A(A[6]), .B(n8), .Z(n36) );
  NANDN U40 ( .A(n8), .B(A[6]), .Z(n34) );
  AND U41 ( .A(n37), .B(n38), .Z(n8) );
  NAND U42 ( .A(B[5]), .B(n39), .Z(n38) );
  NANDN U43 ( .A(A[5]), .B(n10), .Z(n39) );
  NANDN U44 ( .A(n10), .B(A[5]), .Z(n37) );
  AND U45 ( .A(n40), .B(n41), .Z(n10) );
  NAND U46 ( .A(B[4]), .B(n42), .Z(n41) );
  NANDN U47 ( .A(A[4]), .B(n12), .Z(n42) );
  NANDN U48 ( .A(n12), .B(A[4]), .Z(n40) );
  AND U49 ( .A(n43), .B(n44), .Z(n12) );
  NAND U50 ( .A(B[3]), .B(n45), .Z(n44) );
  NANDN U51 ( .A(A[3]), .B(n14), .Z(n45) );
  NANDN U52 ( .A(n14), .B(A[3]), .Z(n43) );
  AND U53 ( .A(n46), .B(n47), .Z(n14) );
  NAND U54 ( .A(B[2]), .B(n48), .Z(n47) );
  NANDN U55 ( .A(A[2]), .B(n16), .Z(n48) );
  NANDN U56 ( .A(n16), .B(A[2]), .Z(n46) );
  AND U57 ( .A(n49), .B(n50), .Z(n16) );
  NAND U58 ( .A(B[1]), .B(n51), .Z(n50) );
  OR U59 ( .A(n18), .B(A[1]), .Z(n51) );
  NAND U60 ( .A(A[1]), .B(n18), .Z(n49) );
  AND U61 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U62 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_3 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(B[9]), .B(n22), .Z(n21) );
  OR U21 ( .A(n2), .B(A[9]), .Z(n22) );
  NAND U22 ( .A(A[9]), .B(n2), .Z(n20) );
  NAND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(B[8]), .B(n25), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(B[7]), .B(n28), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(B[6]), .B(n31), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(B[5]), .B(n34), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(B[4]), .B(n37), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(B[3]), .B(n40), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(B[2]), .B(n43), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(B[1]), .B(n46), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(A[1]), .B(n18), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_4 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(B[9]), .B(n22), .Z(n21) );
  OR U21 ( .A(n2), .B(A[9]), .Z(n22) );
  NAND U22 ( .A(A[9]), .B(n2), .Z(n20) );
  NAND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(B[8]), .B(n25), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(B[7]), .B(n28), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(B[6]), .B(n31), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(B[5]), .B(n34), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(B[4]), .B(n37), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(B[3]), .B(n40), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(B[2]), .B(n43), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(B[1]), .B(n46), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(A[1]), .B(n18), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_5 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AND U1 ( .A(B[9]), .B(n19), .Z(SUM[10]) );
  IV U2 ( .A(B[9]), .Z(n2) );
  XNOR U3 ( .A(n19), .B(n2), .Z(SUM[9]) );
  XOR U4 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U6 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U8 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U10 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U12 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U14 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U16 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U18 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n18) );
  NAND U20 ( .A(n20), .B(n21), .Z(n19) );
  NAND U21 ( .A(B[8]), .B(n22), .Z(n21) );
  NANDN U22 ( .A(A[8]), .B(n3), .Z(n22) );
  NANDN U23 ( .A(n3), .B(A[8]), .Z(n20) );
  AND U24 ( .A(n23), .B(n24), .Z(n3) );
  NAND U25 ( .A(B[7]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(A[7]), .B(n5), .Z(n25) );
  NANDN U27 ( .A(n5), .B(A[7]), .Z(n23) );
  AND U28 ( .A(n26), .B(n27), .Z(n5) );
  NAND U29 ( .A(B[6]), .B(n28), .Z(n27) );
  NANDN U30 ( .A(A[6]), .B(n7), .Z(n28) );
  NANDN U31 ( .A(n7), .B(A[6]), .Z(n26) );
  AND U32 ( .A(n29), .B(n30), .Z(n7) );
  NAND U33 ( .A(B[5]), .B(n31), .Z(n30) );
  NANDN U34 ( .A(A[5]), .B(n9), .Z(n31) );
  NANDN U35 ( .A(n9), .B(A[5]), .Z(n29) );
  AND U36 ( .A(n32), .B(n33), .Z(n9) );
  NAND U37 ( .A(B[4]), .B(n34), .Z(n33) );
  NANDN U38 ( .A(A[4]), .B(n11), .Z(n34) );
  NANDN U39 ( .A(n11), .B(A[4]), .Z(n32) );
  AND U40 ( .A(n35), .B(n36), .Z(n11) );
  NAND U41 ( .A(B[3]), .B(n37), .Z(n36) );
  NANDN U42 ( .A(A[3]), .B(n13), .Z(n37) );
  NANDN U43 ( .A(n13), .B(A[3]), .Z(n35) );
  AND U44 ( .A(n38), .B(n39), .Z(n13) );
  NAND U45 ( .A(B[2]), .B(n40), .Z(n39) );
  NANDN U46 ( .A(A[2]), .B(n15), .Z(n40) );
  NANDN U47 ( .A(n15), .B(A[2]), .Z(n38) );
  AND U48 ( .A(n41), .B(n42), .Z(n15) );
  NAND U49 ( .A(B[1]), .B(n43), .Z(n42) );
  OR U50 ( .A(n17), .B(A[1]), .Z(n43) );
  NAND U51 ( .A(A[1]), .B(n17), .Z(n41) );
  AND U52 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U53 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_6 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_7 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_8 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_9 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_10 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39;

  AND U1 ( .A(B[8]), .B(n2), .Z(SUM[9]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[8]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U18 ( .A(B[1]), .B(A[1]), .Z(n18) );
  AND U19 ( .A(n19), .B(n20), .Z(n4) );
  NAND U20 ( .A(B[7]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[7]), .B(n5), .Z(n21) );
  NANDN U22 ( .A(n5), .B(A[7]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n5) );
  NAND U24 ( .A(B[6]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[6]), .B(n7), .Z(n24) );
  NANDN U26 ( .A(n7), .B(A[6]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n7) );
  NAND U28 ( .A(B[5]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[5]), .B(n9), .Z(n27) );
  NANDN U30 ( .A(n9), .B(A[5]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n9) );
  NAND U32 ( .A(B[4]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[4]), .B(n11), .Z(n30) );
  NANDN U34 ( .A(n11), .B(A[4]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n11) );
  NAND U36 ( .A(B[3]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[3]), .B(n13), .Z(n33) );
  NANDN U38 ( .A(n13), .B(A[3]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n13) );
  NAND U40 ( .A(B[2]), .B(n36), .Z(n35) );
  NANDN U41 ( .A(A[2]), .B(n15), .Z(n36) );
  NANDN U42 ( .A(n15), .B(A[2]), .Z(n34) );
  AND U43 ( .A(n37), .B(n38), .Z(n15) );
  NAND U44 ( .A(B[1]), .B(n39), .Z(n38) );
  OR U45 ( .A(n17), .B(A[1]), .Z(n39) );
  NAND U46 ( .A(A[1]), .B(n17), .Z(n37) );
  AND U47 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U48 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_11 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_12 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_13 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_14 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_15 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_16 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_17 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_18 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_19 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_20 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_21 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_22 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_23 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_24 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_25 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_26 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_27 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_28 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_29 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_30 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_31 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_32 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_33 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_34 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_35 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_36 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_37 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_38 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_39 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_40 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_41 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_42 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_43 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_44 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_45 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_46 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_47 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_48 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_49 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_50 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_51 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_52 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_53 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_54 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_55 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_56 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_57 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_58 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_59 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_60 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_61 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_62 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_63 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_64 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_65 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_66 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_67 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_68 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_69 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_70 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_71 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_72 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_73 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_74 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_75 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_76 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_77 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_78 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_79 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_80 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_81 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_82 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_83 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;

  AND U1 ( .A(B[5]), .B(n2), .Z(SUM[6]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[5]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[3]) );
  XNOR U8 ( .A(B[3]), .B(A[3]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[2]) );
  XNOR U10 ( .A(B[2]), .B(A[2]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[1]) );
  XOR U12 ( .A(B[1]), .B(A[1]), .Z(n12) );
  AND U13 ( .A(n13), .B(n14), .Z(n4) );
  NAND U14 ( .A(B[4]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[4]), .B(n5), .Z(n15) );
  NANDN U16 ( .A(n5), .B(A[4]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n5) );
  NAND U18 ( .A(B[3]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[3]), .B(n7), .Z(n18) );
  NANDN U20 ( .A(n7), .B(A[3]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n7) );
  NAND U22 ( .A(B[2]), .B(n21), .Z(n20) );
  NANDN U23 ( .A(A[2]), .B(n9), .Z(n21) );
  NANDN U24 ( .A(n9), .B(A[2]), .Z(n19) );
  AND U25 ( .A(n22), .B(n23), .Z(n9) );
  NAND U26 ( .A(B[1]), .B(n24), .Z(n23) );
  OR U27 ( .A(n11), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(A[1]), .B(n11), .Z(n22) );
  AND U29 ( .A(B[0]), .B(A[0]), .Z(n11) );
  XOR U30 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_84 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_85 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_86 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_87 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_88 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_89 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_90 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_91 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_92 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_93 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_94 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_95 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_96 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_97 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_98 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_99 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_100 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_101 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_102 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_103 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_104 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_105 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_106 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_107 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_108 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_109 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_110 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_111 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_112 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_113 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_114 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_115 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_116 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_117 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_118 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_119 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_120 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_121 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_122 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_123 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_124 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_125 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_126 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_127 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_128 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_129 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_130 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_131 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_132 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_133 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_134 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_135 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_136 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_137 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_138 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_139 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_140 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_141 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_142 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_143 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_144 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_145 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_146 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_147 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_148 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_149 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_150 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_151 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_152 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_153 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_154 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_155 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_156 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_157 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_158 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_159 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_160 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_161 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_162 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_163 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_164 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_165 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4_DW01_add_166 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC4 ( clk, rst, x, y, o );
  input [3999:0] x;
  input [3999:0] y;
  output [13:0] o;
  input clk, rst;
  wire   N27929, N27930, N27931, N27932, N27933, N27941, N27942, N27943,
         N27944, N27945, N27953, N27954, N27955, N27956, N27957, N27965,
         N27966, N27967, N27968, N27969, N27977, N27978, N27979, N27980,
         N27981, N27989, N27990, N27991, N27992, N27993, N28001, N28002,
         N28003, N28004, N28005, N28013, N28014, N28015, N28016, N28017,
         N28025, N28026, N28027, N28028, N28029, N28037, N28038, N28039,
         N28040, N28041, N28049, N28050, N28051, N28052, N28053, N28061,
         N28062, N28063, N28064, N28065, N28073, N28074, N28075, N28076,
         N28077, N28085, N28086, N28087, N28088, N28089, N28097, N28098,
         N28099, N28100, N28101, N28109, N28110, N28111, N28112, N28113,
         N28121, N28122, N28123, N28124, N28125, N28133, N28134, N28135,
         N28136, N28137, N28145, N28146, N28147, N28148, N28149, N28157,
         N28158, N28159, N28160, N28161, N28169, N28170, N28171, N28172,
         N28173, N28181, N28182, N28183, N28184, N28185, N28193, N28194,
         N28195, N28196, N28197, N28205, N28206, N28207, N28208, N28209,
         N28217, N28218, N28219, N28220, N28221, N28229, N28230, N28231,
         N28232, N28233, N28241, N28242, N28243, N28244, N28245, N28253,
         N28254, N28255, N28256, N28257, N28265, N28266, N28267, N28268,
         N28269, N28277, N28278, N28279, N28280, N28281, N28289, N28290,
         N28291, N28292, N28293, N28301, N28302, N28303, N28304, N28305,
         N28313, N28314, N28315, N28316, N28317, N28325, N28326, N28327,
         N28328, N28329, N28337, N28338, N28339, N28340, N28341, N28349,
         N28350, N28351, N28352, N28353, N28361, N28362, N28363, N28364,
         N28365, N28373, N28374, N28375, N28376, N28377, N28385, N28386,
         N28387, N28388, N28389, N28397, N28398, N28399, N28400, N28401,
         N28409, N28410, N28411, N28412, N28413, N28421, N28422, N28423,
         N28424, N28425, N28433, N28434, N28435, N28436, N28437, N28445,
         N28446, N28447, N28448, N28449, N28457, N28458, N28459, N28460,
         N28461, N28469, N28470, N28471, N28472, N28473, N28481, N28482,
         N28483, N28484, N28485, N28493, N28494, N28495, N28496, N28497,
         N28505, N28506, N28507, N28508, N28509, N28517, N28518, N28519,
         N28520, N28521, N28529, N28530, N28531, N28532, N28533, N28541,
         N28542, N28543, N28544, N28545, N28553, N28554, N28555, N28556,
         N28557, N28565, N28566, N28567, N28568, N28569, N28577, N28578,
         N28579, N28580, N28581, N28589, N28590, N28591, N28592, N28593,
         N28601, N28602, N28603, N28604, N28605, N28613, N28614, N28615,
         N28616, N28617, N28625, N28626, N28627, N28628, N28629, N28637,
         N28638, N28639, N28640, N28641, N28649, N28650, N28651, N28652,
         N28653, N28661, N28662, N28663, N28664, N28665, N28673, N28674,
         N28675, N28676, N28677, N28685, N28686, N28687, N28688, N28689,
         N28697, N28698, N28699, N28700, N28701, N28709, N28710, N28711,
         N28712, N28713, N28721, N28722, N28723, N28724, N28725, N28733,
         N28734, N28735, N28736, N28737, N28745, N28746, N28747, N28748,
         N28749, N28757, N28758, N28759, N28760, N28761, N28769, N28770,
         N28771, N28772, N28773, N28781, N28782, N28783, N28784, N28785,
         N28793, N28794, N28795, N28796, N28797, N28805, N28806, N28807,
         N28808, N28809, N28817, N28818, N28819, N28820, N28821, N28829,
         N28830, N28831, N28832, N28833, N28841, N28842, N28843, N28844,
         N28845, N28853, N28854, N28855, N28856, N28857, N28865, N28866,
         N28867, N28868, N28869, N28877, N28878, N28879, N28880, N28881,
         N28889, N28890, N28891, N28892, N28893, N28901, N28902, N28903,
         N28904, N28905, N28913, N28914, N28915, N28916, N28917, N28925,
         N28926, N28927, N28928, N28929, N28937, N28938, N28939, N28940,
         N28941, N28949, N28950, N28951, N28952, N28953, N28961, N28962,
         N28963, N28964, N28965, N28973, N28974, N28975, N28976, N28977,
         N28985, N28986, N28987, N28988, N28989, N28997, N28998, N28999,
         N29000, N29001, N29009, N29010, N29011, N29012, N29013, N29021,
         N29022, N29023, N29024, N29025, N29033, N29034, N29035, N29036,
         N29037, N29045, N29046, N29047, N29048, N29049, N29057, N29058,
         N29059, N29060, N29061, N29069, N29070, N29071, N29072, N29073,
         N29081, N29082, N29083, N29084, N29085, N29093, N29094, N29095,
         N29096, N29097, N29105, N29106, N29107, N29108, N29109, N29117,
         N29118, N29119, N29120, N29121, N29129, N29130, N29131, N29132,
         N29133, N29141, N29142, N29143, N29144, N29145, N29153, N29154,
         N29155, N29156, N29157, N29165, N29166, N29167, N29168, N29169,
         N29177, N29178, N29179, N29180, N29181, N29189, N29190, N29191,
         N29192, N29193, N29201, N29202, N29203, N29204, N29205, N29213,
         N29214, N29215, N29216, N29217, N29225, N29226, N29227, N29228,
         N29229, N29237, N29238, N29239, N29240, N29241, N29249, N29250,
         N29251, N29252, N29253, N29261, N29262, N29263, N29264, N29265,
         N29273, N29274, N29275, N29276, N29277, N29285, N29286, N29287,
         N29288, N29289, N29297, N29298, N29299, N29300, N29301, N29309,
         N29310, N29311, N29312, N29313, N29321, N29322, N29323, N29324,
         N29325, N29333, N29334, N29335, N29336, N29337, N29345, N29346,
         N29347, N29348, N29349, N29357, N29358, N29359, N29360, N29361,
         N29369, N29370, N29371, N29372, N29373, N29381, N29382, N29383,
         N29384, N29385, N29393, N29394, N29395, N29396, N29397, N29405,
         N29406, N29407, N29408, N29409, N29417, N29418, N29419, N29420,
         N29421, N29429, N29430, N29431, N29432, N29433, N29441, N29442,
         N29443, N29444, N29445, N29453, N29454, N29455, N29456, N29457,
         N29465, N29466, N29467, N29468, N29469, N29477, N29478, N29479,
         N29480, N29481, N29489, N29490, N29491, N29492, N29493, N29501,
         N29502, N29503, N29504, N29505, N29513, N29514, N29515, N29516,
         N29517, N29525, N29526, N29527, N29528, N29529, N29537, N29538,
         N29539, N29540, N29541, N29549, N29550, N29551, N29552, N29553,
         N29561, N29562, N29563, N29564, N29565, N29573, N29574, N29575,
         N29576, N29577, N29585, N29586, N29587, N29588, N29589, N29597,
         N29598, N29599, N29600, N29601, N29609, N29610, N29611, N29612,
         N29613, N29621, N29622, N29623, N29624, N29625, N29633, N29634,
         N29635, N29636, N29637, N29645, N29646, N29647, N29648, N29649,
         N29657, N29658, N29659, N29660, N29661, N29669, N29670, N29671,
         N29672, N29673, N29681, N29682, N29683, N29684, N29685, N29693,
         N29694, N29695, N29696, N29697, N29705, N29706, N29707, N29708,
         N29709, N29717, N29718, N29719, N29720, N29721, N29729, N29730,
         N29731, N29732, N29733, N29741, N29742, N29743, N29744, N29745,
         N29753, N29754, N29755, N29756, N29757, N29765, N29766, N29767,
         N29768, N29769, N29777, N29778, N29779, N29780, N29781, N29789,
         N29790, N29791, N29792, N29793, N29801, N29802, N29803, N29804,
         N29805, N29813, N29814, N29815, N29816, N29817, N29825, N29826,
         N29827, N29828, N29829, N29837, N29838, N29839, N29840, N29841,
         N29849, N29850, N29851, N29852, N29853, N29861, N29862, N29863,
         N29864, N29865, N29873, N29874, N29875, N29876, N29877, N29885,
         N29886, N29887, N29888, N29889, N29897, N29898, N29899, N29900,
         N29901, N29909, N29910, N29911, N29912, N29913, N29921, N29922,
         N29923, N29924, N29925, N29933, N29934, N29935, N29936, N29937,
         N29938, N29945, N29946, N29947, N29948, N29949, N29950, N29957,
         N29958, N29959, N29960, N29961, N29962, N29969, N29970, N29971,
         N29972, N29973, N29974, N29981, N29982, N29983, N29984, N29985,
         N29986, N29993, N29994, N29995, N29996, N29997, N29998, N30005,
         N30006, N30007, N30008, N30009, N30010, N30017, N30018, N30019,
         N30020, N30021, N30022, N30029, N30030, N30031, N30032, N30033,
         N30034, N30041, N30042, N30043, N30044, N30045, N30046, N30053,
         N30054, N30055, N30056, N30057, N30058, N30065, N30066, N30067,
         N30068, N30069, N30070, N30077, N30078, N30079, N30080, N30081,
         N30082, N30089, N30090, N30091, N30092, N30093, N30094, N30101,
         N30102, N30103, N30104, N30105, N30106, N30113, N30114, N30115,
         N30116, N30117, N30118, N30125, N30126, N30127, N30128, N30129,
         N30130, N30137, N30138, N30139, N30140, N30141, N30142, N30149,
         N30150, N30151, N30152, N30153, N30154, N30161, N30162, N30163,
         N30164, N30165, N30166, N30173, N30174, N30175, N30176, N30177,
         N30178, N30185, N30186, N30187, N30188, N30189, N30190, N30197,
         N30198, N30199, N30200, N30201, N30202, N30209, N30210, N30211,
         N30212, N30213, N30214, N30221, N30222, N30223, N30224, N30225,
         N30226, N30233, N30234, N30235, N30236, N30237, N30238, N30245,
         N30246, N30247, N30248, N30249, N30250, N30257, N30258, N30259,
         N30260, N30261, N30262, N30269, N30270, N30271, N30272, N30273,
         N30274, N30281, N30282, N30283, N30284, N30285, N30286, N30293,
         N30294, N30295, N30296, N30297, N30298, N30305, N30306, N30307,
         N30308, N30309, N30310, N30317, N30318, N30319, N30320, N30321,
         N30322, N30329, N30330, N30331, N30332, N30333, N30334, N30341,
         N30342, N30343, N30344, N30345, N30346, N30353, N30354, N30355,
         N30356, N30357, N30358, N30365, N30366, N30367, N30368, N30369,
         N30370, N30377, N30378, N30379, N30380, N30381, N30382, N30389,
         N30390, N30391, N30392, N30393, N30394, N30401, N30402, N30403,
         N30404, N30405, N30406, N30413, N30414, N30415, N30416, N30417,
         N30418, N30425, N30426, N30427, N30428, N30429, N30430, N30437,
         N30438, N30439, N30440, N30441, N30442, N30449, N30450, N30451,
         N30452, N30453, N30454, N30461, N30462, N30463, N30464, N30465,
         N30466, N30473, N30474, N30475, N30476, N30477, N30478, N30485,
         N30486, N30487, N30488, N30489, N30490, N30497, N30498, N30499,
         N30500, N30501, N30502, N30509, N30510, N30511, N30512, N30513,
         N30514, N30521, N30522, N30523, N30524, N30525, N30526, N30533,
         N30534, N30535, N30536, N30537, N30538, N30545, N30546, N30547,
         N30548, N30549, N30550, N30557, N30558, N30559, N30560, N30561,
         N30562, N30569, N30570, N30571, N30572, N30573, N30574, N30581,
         N30582, N30583, N30584, N30585, N30586, N30593, N30594, N30595,
         N30596, N30597, N30598, N30605, N30606, N30607, N30608, N30609,
         N30610, N30617, N30618, N30619, N30620, N30621, N30622, N30629,
         N30630, N30631, N30632, N30633, N30634, N30641, N30642, N30643,
         N30644, N30645, N30646, N30653, N30654, N30655, N30656, N30657,
         N30658, N30665, N30666, N30667, N30668, N30669, N30670, N30677,
         N30678, N30679, N30680, N30681, N30682, N30689, N30690, N30691,
         N30692, N30693, N30694, N30701, N30702, N30703, N30704, N30705,
         N30706, N30713, N30714, N30715, N30716, N30717, N30718, N30725,
         N30726, N30727, N30728, N30729, N30730, N30737, N30738, N30739,
         N30740, N30741, N30742, N30749, N30750, N30751, N30752, N30753,
         N30754, N30761, N30762, N30763, N30764, N30765, N30766, N30773,
         N30774, N30775, N30776, N30777, N30778, N30785, N30786, N30787,
         N30788, N30789, N30790, N30797, N30798, N30799, N30800, N30801,
         N30802, N30809, N30810, N30811, N30812, N30813, N30814, N30821,
         N30822, N30823, N30824, N30825, N30826, N30833, N30834, N30835,
         N30836, N30837, N30838, N30845, N30846, N30847, N30848, N30849,
         N30850, N30857, N30858, N30859, N30860, N30861, N30862, N30869,
         N30870, N30871, N30872, N30873, N30874, N30881, N30882, N30883,
         N30884, N30885, N30886, N30893, N30894, N30895, N30896, N30897,
         N30898, N30905, N30906, N30907, N30908, N30909, N30910, N30917,
         N30918, N30919, N30920, N30921, N30922, N30929, N30930, N30931,
         N30932, N30933, N30934, N30935, N30941, N30942, N30943, N30944,
         N30945, N30946, N30947, N30953, N30954, N30955, N30956, N30957,
         N30958, N30959, N30965, N30966, N30967, N30968, N30969, N30970,
         N30971, N30977, N30978, N30979, N30980, N30981, N30982, N30983,
         N30989, N30990, N30991, N30992, N30993, N30994, N30995, N31001,
         N31002, N31003, N31004, N31005, N31006, N31007, N31013, N31014,
         N31015, N31016, N31017, N31018, N31019, N31025, N31026, N31027,
         N31028, N31029, N31030, N31031, N31037, N31038, N31039, N31040,
         N31041, N31042, N31043, N31049, N31050, N31051, N31052, N31053,
         N31054, N31055, N31061, N31062, N31063, N31064, N31065, N31066,
         N31067, N31073, N31074, N31075, N31076, N31077, N31078, N31079,
         N31085, N31086, N31087, N31088, N31089, N31090, N31091, N31097,
         N31098, N31099, N31100, N31101, N31102, N31103, N31109, N31110,
         N31111, N31112, N31113, N31114, N31115, N31121, N31122, N31123,
         N31124, N31125, N31126, N31127, N31133, N31134, N31135, N31136,
         N31137, N31138, N31139, N31145, N31146, N31147, N31148, N31149,
         N31150, N31151, N31157, N31158, N31159, N31160, N31161, N31162,
         N31163, N31169, N31170, N31171, N31172, N31173, N31174, N31175,
         N31181, N31182, N31183, N31184, N31185, N31186, N31187, N31193,
         N31194, N31195, N31196, N31197, N31198, N31199, N31205, N31206,
         N31207, N31208, N31209, N31210, N31211, N31217, N31218, N31219,
         N31220, N31221, N31222, N31223, N31229, N31230, N31231, N31232,
         N31233, N31234, N31235, N31241, N31242, N31243, N31244, N31245,
         N31246, N31247, N31253, N31254, N31255, N31256, N31257, N31258,
         N31259, N31265, N31266, N31267, N31268, N31269, N31270, N31271,
         N31277, N31278, N31279, N31280, N31281, N31282, N31283, N31289,
         N31290, N31291, N31292, N31293, N31294, N31295, N31301, N31302,
         N31303, N31304, N31305, N31306, N31307, N31313, N31314, N31315,
         N31316, N31317, N31318, N31319, N31325, N31326, N31327, N31328,
         N31329, N31330, N31331, N31337, N31338, N31339, N31340, N31341,
         N31342, N31343, N31349, N31350, N31351, N31352, N31353, N31354,
         N31355, N31361, N31362, N31363, N31364, N31365, N31366, N31367,
         N31373, N31374, N31375, N31376, N31377, N31378, N31379, N31385,
         N31386, N31387, N31388, N31389, N31390, N31391, N31397, N31398,
         N31399, N31400, N31401, N31402, N31403, N31409, N31410, N31411,
         N31412, N31413, N31414, N31415, N31421, N31422, N31423, N31424,
         N31425, N31426, N31427, N31433, N31434, N31435, N31436, N31437,
         N31438, N31439, N31440, N31445, N31446, N31447, N31448, N31449,
         N31450, N31451, N31452, N31457, N31458, N31459, N31460, N31461,
         N31462, N31463, N31464, N31469, N31470, N31471, N31472, N31473,
         N31474, N31475, N31476, N31481, N31482, N31483, N31484, N31485,
         N31486, N31487, N31488, N31493, N31494, N31495, N31496, N31497,
         N31498, N31499, N31500, N31505, N31506, N31507, N31508, N31509,
         N31510, N31511, N31512, N31517, N31518, N31519, N31520, N31521,
         N31522, N31523, N31524, N31529, N31530, N31531, N31532, N31533,
         N31534, N31535, N31536, N31541, N31542, N31543, N31544, N31545,
         N31546, N31547, N31548, N31553, N31554, N31555, N31556, N31557,
         N31558, N31559, N31560, N31565, N31566, N31567, N31568, N31569,
         N31570, N31571, N31572, N31577, N31578, N31579, N31580, N31581,
         N31582, N31583, N31584, N31589, N31590, N31591, N31592, N31593,
         N31594, N31595, N31596, N31601, N31602, N31603, N31604, N31605,
         N31606, N31607, N31608, N31613, N31614, N31615, N31616, N31617,
         N31618, N31619, N31620, N31625, N31626, N31627, N31628, N31629,
         N31630, N31631, N31632, N31637, N31638, N31639, N31640, N31641,
         N31642, N31643, N31644, N31649, N31650, N31651, N31652, N31653,
         N31654, N31655, N31656, N31661, N31662, N31663, N31664, N31665,
         N31666, N31667, N31668, N31673, N31674, N31675, N31676, N31677,
         N31678, N31679, N31680, N31685, N31686, N31687, N31688, N31689,
         N31690, N31691, N31692, N31693, N31697, N31698, N31699, N31700,
         N31701, N31702, N31703, N31704, N31705, N31709, N31710, N31711,
         N31712, N31713, N31714, N31715, N31716, N31717, N31721, N31722,
         N31723, N31724, N31725, N31726, N31727, N31728, N31729, N31733,
         N31734, N31735, N31736, N31737, N31738, N31739, N31740, N31741,
         N31745, N31746, N31747, N31748, N31749, N31750, N31751, N31752,
         N31753, N31757, N31758, N31759, N31760, N31761, N31762, N31763,
         N31764, N31765, N31769, N31770, N31771, N31772, N31773, N31774,
         N31775, N31776, N31777, N31781, N31782, N31783, N31784, N31785,
         N31786, N31787, N31788, N31789, N31793, N31794, N31795, N31796,
         N31797, N31798, N31799, N31800, N31801, N31805, N31806, N31807,
         N31808, N31809, N31810, N31811, N31812, N31813, N31814, N31817,
         N31818, N31819, N31820, N31821, N31822, N31823, N31824, N31825,
         N31826, N31829, N31830, N31831, N31832, N31833, N31834, N31835,
         N31836, N31837, N31838, N31841, N31842, N31843, N31844, N31845,
         N31846, N31847, N31848, N31849, N31850, N31853, N31854, N31855,
         N31856, N31857, N31858, N31859, N31860, N31861, N31862, N31865,
         N31866, N31867, N31868, N31869, N31870, N31871, N31872, N31873,
         N31874, N31875, N31877, N31878, N31879, N31880, N31881, N31882,
         N31883, N31884, N31885, N31886, N31887, N31889, N31890, N31891,
         N31892, N31893, N31894, N31895, N31896, N31897, N31898, N31899,
         N31901, N31902, N31903, N31904, N31905, N31906, N31907, N31908,
         N31909, N31910, N31911, N31912, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
         n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
         n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
         n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
         n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
         n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695,
         n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719,
         n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
         n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
         n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
         n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
         n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
         n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791,
         n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
         n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
         n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
         n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
         n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
         n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847,
         n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
         n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863,
         n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
         n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879,
         n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887,
         n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
         n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903,
         n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911,
         n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919,
         n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927,
         n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935,
         n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943,
         n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
         n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959,
         n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967,
         n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975,
         n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983,
         n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
         n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999,
         n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007,
         n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
         n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
         n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031,
         n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039,
         n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
         n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055,
         n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063,
         n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
         n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079,
         n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087,
         n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095,
         n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103,
         n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111,
         n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119,
         n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127,
         n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
         n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
         n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151,
         n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
         n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167,
         n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175,
         n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183,
         n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191,
         n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199,
         n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207,
         n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
         n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223,
         n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
         n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239,
         n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247,
         n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
         n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263,
         n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
         n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279,
         n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
         n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295,
         n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303,
         n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
         n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319,
         n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327,
         n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335,
         n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343,
         n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351,
         n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
         n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
         n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375,
         n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
         n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391,
         n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399,
         n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407,
         n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415,
         n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423,
         n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
         n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439,
         n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447,
         n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455,
         n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463,
         n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471,
         n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479,
         n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487,
         n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495,
         n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503,
         n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511,
         n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519,
         n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
         n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535,
         n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543,
         n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551,
         n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559,
         n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567,
         n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575,
         n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583,
         n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591,
         n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599,
         n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607,
         n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615,
         n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623,
         n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
         n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
         n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
         n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
         n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663,
         n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
         n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679,
         n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
         n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
         n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703,
         n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
         n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719,
         n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727,
         n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735,
         n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743,
         n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751,
         n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
         n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
         n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
         n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
         n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
         n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799,
         n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807,
         n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815,
         n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823,
         n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
         n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847,
         n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855,
         n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
         n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871,
         n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879,
         n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887,
         n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895,
         n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903,
         n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
         n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919,
         n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927,
         n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
         n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943,
         n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951,
         n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959,
         n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967,
         n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
         n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
         n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991,
         n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999,
         n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
         n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015,
         n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023,
         n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031,
         n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039,
         n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047,
         n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
         n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063,
         n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071,
         n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
         n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087,
         n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095,
         n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103,
         n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111,
         n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119,
         n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
         n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135,
         n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143,
         n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
         n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159,
         n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167,
         n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175,
         n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183,
         n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191,
         n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199,
         n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207,
         n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215,
         n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
         n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231,
         n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239,
         n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247,
         n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255,
         n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
         n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271,
         n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279,
         n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287,
         n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
         n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303,
         n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311,
         n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319,
         n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327,
         n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
         n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343,
         n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351,
         n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359,
         n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367,
         n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375,
         n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383,
         n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391,
         n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399,
         n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
         n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
         n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423,
         n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431,
         n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
         n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447,
         n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455,
         n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463,
         n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471,
         n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
         n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487,
         n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495,
         n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503,
         n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511,
         n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519,
         n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527,
         n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535,
         n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543,
         n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
         n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559,
         n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567,
         n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
         n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
         n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591,
         n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599,
         n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607,
         n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615,
         n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
         n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631,
         n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639,
         n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647,
         n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
         n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663,
         n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671,
         n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679,
         n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687,
         n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695,
         n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703,
         n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711,
         n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719,
         n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727,
         n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735,
         n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743,
         n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751,
         n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759,
         n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767,
         n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775,
         n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783,
         n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791,
         n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799,
         n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807,
         n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815,
         n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823,
         n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831,
         n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839,
         n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847,
         n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855,
         n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863,
         n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871,
         n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879,
         n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887,
         n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895,
         n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903,
         n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911,
         n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
         n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927,
         n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
         n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943,
         n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951,
         n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959,
         n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967,
         n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975,
         n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983,
         n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991,
         n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999,
         n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
         n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015,
         n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023,
         n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031,
         n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
         n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047,
         n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055,
         n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063,
         n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071,
         n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079,
         n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087,
         n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095,
         n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103,
         n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111,
         n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119,
         n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127,
         n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135,
         n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143,
         n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151,
         n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159,
         n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167,
         n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175,
         n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183,
         n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191,
         n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199,
         n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207,
         n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215,
         n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223,
         n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231,
         n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239,
         n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247,
         n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255,
         n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263,
         n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271,
         n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279,
         n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287,
         n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295,
         n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303,
         n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311,
         n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319,
         n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327,
         n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335,
         n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343,
         n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351,
         n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359,
         n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367,
         n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375,
         n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383,
         n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391,
         n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399,
         n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407,
         n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
         n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423,
         n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431,
         n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439,
         n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
         n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455,
         n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463,
         n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471,
         n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479,
         n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487,
         n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495,
         n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503,
         n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511,
         n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519,
         n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527,
         n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535,
         n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543,
         n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551,
         n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559,
         n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567,
         n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575,
         n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583,
         n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591,
         n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599,
         n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607,
         n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615,
         n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623,
         n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631,
         n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639,
         n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647,
         n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655,
         n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663,
         n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671,
         n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679,
         n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687,
         n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695,
         n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703,
         n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711,
         n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719,
         n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727,
         n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735,
         n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743,
         n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751,
         n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759,
         n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767,
         n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775,
         n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783,
         n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791,
         n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799,
         n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807,
         n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815,
         n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823,
         n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831,
         n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839,
         n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847,
         n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855,
         n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863,
         n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871,
         n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879,
         n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887,
         n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895,
         n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903,
         n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911,
         n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919,
         n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927,
         n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935,
         n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943,
         n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951,
         n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959,
         n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967,
         n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975,
         n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983,
         n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991,
         n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999,
         n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007,
         n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015,
         n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023,
         n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031,
         n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039,
         n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047,
         n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055,
         n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063,
         n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
         n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079,
         n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087,
         n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095,
         n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103,
         n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111,
         n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119,
         n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127,
         n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
         n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143,
         n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151,
         n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159,
         n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167,
         n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175,
         n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183,
         n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191,
         n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199,
         n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207,
         n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215,
         n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223,
         n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231,
         n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239,
         n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247,
         n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255,
         n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263,
         n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271,
         n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
         n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287,
         n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295,
         n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303,
         n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311,
         n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319,
         n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327,
         n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335,
         n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343,
         n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351,
         n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359,
         n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367,
         n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375,
         n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383,
         n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391,
         n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399,
         n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
         n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415,
         n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
         n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431,
         n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439,
         n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447,
         n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455,
         n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463,
         n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471,
         n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479,
         n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487,
         n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
         n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503,
         n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511,
         n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519,
         n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
         n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535,
         n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543,
         n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551,
         n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559,
         n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567,
         n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575,
         n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583,
         n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591,
         n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599,
         n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607,
         n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615,
         n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623,
         n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631,
         n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639,
         n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647,
         n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655,
         n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663,
         n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671,
         n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679,
         n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687,
         n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695,
         n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703,
         n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711,
         n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719,
         n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727,
         n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735,
         n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743,
         n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751,
         n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759,
         n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767,
         n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775,
         n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
         n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791,
         n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799,
         n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807,
         n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
         n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823,
         n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831,
         n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839,
         n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847,
         n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855,
         n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863,
         n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871,
         n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879,
         n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887,
         n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895,
         n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903,
         n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911,
         n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919,
         n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927,
         n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935,
         n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943,
         n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951,
         n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
         n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967,
         n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975,
         n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
         n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991,
         n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999,
         n27000, n27001, n27002, n27003;
  wire   [11:0] olocal;
  wire   [13:0] oglobal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, 
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, 
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, 
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        SYNOPSYS_UNCONNECTED__352, SYNOPSYS_UNCONNECTED__353, 
        SYNOPSYS_UNCONNECTED__354, SYNOPSYS_UNCONNECTED__355, 
        SYNOPSYS_UNCONNECTED__356, SYNOPSYS_UNCONNECTED__357, 
        SYNOPSYS_UNCONNECTED__358, SYNOPSYS_UNCONNECTED__359, 
        SYNOPSYS_UNCONNECTED__360, SYNOPSYS_UNCONNECTED__361, 
        SYNOPSYS_UNCONNECTED__362, SYNOPSYS_UNCONNECTED__363, 
        SYNOPSYS_UNCONNECTED__364, SYNOPSYS_UNCONNECTED__365, 
        SYNOPSYS_UNCONNECTED__366, SYNOPSYS_UNCONNECTED__367, 
        SYNOPSYS_UNCONNECTED__368, SYNOPSYS_UNCONNECTED__369, 
        SYNOPSYS_UNCONNECTED__370, SYNOPSYS_UNCONNECTED__371, 
        SYNOPSYS_UNCONNECTED__372, SYNOPSYS_UNCONNECTED__373, 
        SYNOPSYS_UNCONNECTED__374, SYNOPSYS_UNCONNECTED__375, 
        SYNOPSYS_UNCONNECTED__376, SYNOPSYS_UNCONNECTED__377, 
        SYNOPSYS_UNCONNECTED__378, SYNOPSYS_UNCONNECTED__379, 
        SYNOPSYS_UNCONNECTED__380, SYNOPSYS_UNCONNECTED__381, 
        SYNOPSYS_UNCONNECTED__382, SYNOPSYS_UNCONNECTED__383, 
        SYNOPSYS_UNCONNECTED__384, SYNOPSYS_UNCONNECTED__385, 
        SYNOPSYS_UNCONNECTED__386, SYNOPSYS_UNCONNECTED__387, 
        SYNOPSYS_UNCONNECTED__388, SYNOPSYS_UNCONNECTED__389, 
        SYNOPSYS_UNCONNECTED__390, SYNOPSYS_UNCONNECTED__391, 
        SYNOPSYS_UNCONNECTED__392, SYNOPSYS_UNCONNECTED__393, 
        SYNOPSYS_UNCONNECTED__394, SYNOPSYS_UNCONNECTED__395, 
        SYNOPSYS_UNCONNECTED__396, SYNOPSYS_UNCONNECTED__397, 
        SYNOPSYS_UNCONNECTED__398, SYNOPSYS_UNCONNECTED__399, 
        SYNOPSYS_UNCONNECTED__400, SYNOPSYS_UNCONNECTED__401, 
        SYNOPSYS_UNCONNECTED__402, SYNOPSYS_UNCONNECTED__403, 
        SYNOPSYS_UNCONNECTED__404, SYNOPSYS_UNCONNECTED__405, 
        SYNOPSYS_UNCONNECTED__406, SYNOPSYS_UNCONNECTED__407, 
        SYNOPSYS_UNCONNECTED__408, SYNOPSYS_UNCONNECTED__409, 
        SYNOPSYS_UNCONNECTED__410, SYNOPSYS_UNCONNECTED__411, 
        SYNOPSYS_UNCONNECTED__412, SYNOPSYS_UNCONNECTED__413, 
        SYNOPSYS_UNCONNECTED__414, SYNOPSYS_UNCONNECTED__415, 
        SYNOPSYS_UNCONNECTED__416, SYNOPSYS_UNCONNECTED__417, 
        SYNOPSYS_UNCONNECTED__418, SYNOPSYS_UNCONNECTED__419, 
        SYNOPSYS_UNCONNECTED__420, SYNOPSYS_UNCONNECTED__421, 
        SYNOPSYS_UNCONNECTED__422, SYNOPSYS_UNCONNECTED__423, 
        SYNOPSYS_UNCONNECTED__424, SYNOPSYS_UNCONNECTED__425, 
        SYNOPSYS_UNCONNECTED__426, SYNOPSYS_UNCONNECTED__427, 
        SYNOPSYS_UNCONNECTED__428, SYNOPSYS_UNCONNECTED__429, 
        SYNOPSYS_UNCONNECTED__430, SYNOPSYS_UNCONNECTED__431, 
        SYNOPSYS_UNCONNECTED__432, SYNOPSYS_UNCONNECTED__433, 
        SYNOPSYS_UNCONNECTED__434, SYNOPSYS_UNCONNECTED__435, 
        SYNOPSYS_UNCONNECTED__436, SYNOPSYS_UNCONNECTED__437, 
        SYNOPSYS_UNCONNECTED__438, SYNOPSYS_UNCONNECTED__439, 
        SYNOPSYS_UNCONNECTED__440, SYNOPSYS_UNCONNECTED__441, 
        SYNOPSYS_UNCONNECTED__442, SYNOPSYS_UNCONNECTED__443, 
        SYNOPSYS_UNCONNECTED__444, SYNOPSYS_UNCONNECTED__445, 
        SYNOPSYS_UNCONNECTED__446, SYNOPSYS_UNCONNECTED__447, 
        SYNOPSYS_UNCONNECTED__448, SYNOPSYS_UNCONNECTED__449, 
        SYNOPSYS_UNCONNECTED__450, SYNOPSYS_UNCONNECTED__451, 
        SYNOPSYS_UNCONNECTED__452, SYNOPSYS_UNCONNECTED__453, 
        SYNOPSYS_UNCONNECTED__454, SYNOPSYS_UNCONNECTED__455, 
        SYNOPSYS_UNCONNECTED__456, SYNOPSYS_UNCONNECTED__457, 
        SYNOPSYS_UNCONNECTED__458, SYNOPSYS_UNCONNECTED__459, 
        SYNOPSYS_UNCONNECTED__460, SYNOPSYS_UNCONNECTED__461, 
        SYNOPSYS_UNCONNECTED__462, SYNOPSYS_UNCONNECTED__463, 
        SYNOPSYS_UNCONNECTED__464, SYNOPSYS_UNCONNECTED__465, 
        SYNOPSYS_UNCONNECTED__466, SYNOPSYS_UNCONNECTED__467, 
        SYNOPSYS_UNCONNECTED__468, SYNOPSYS_UNCONNECTED__469, 
        SYNOPSYS_UNCONNECTED__470, SYNOPSYS_UNCONNECTED__471, 
        SYNOPSYS_UNCONNECTED__472, SYNOPSYS_UNCONNECTED__473, 
        SYNOPSYS_UNCONNECTED__474, SYNOPSYS_UNCONNECTED__475, 
        SYNOPSYS_UNCONNECTED__476, SYNOPSYS_UNCONNECTED__477, 
        SYNOPSYS_UNCONNECTED__478, SYNOPSYS_UNCONNECTED__479, 
        SYNOPSYS_UNCONNECTED__480, SYNOPSYS_UNCONNECTED__481, 
        SYNOPSYS_UNCONNECTED__482, SYNOPSYS_UNCONNECTED__483, 
        SYNOPSYS_UNCONNECTED__484, SYNOPSYS_UNCONNECTED__485, 
        SYNOPSYS_UNCONNECTED__486, SYNOPSYS_UNCONNECTED__487, 
        SYNOPSYS_UNCONNECTED__488, SYNOPSYS_UNCONNECTED__489, 
        SYNOPSYS_UNCONNECTED__490, SYNOPSYS_UNCONNECTED__491, 
        SYNOPSYS_UNCONNECTED__492, SYNOPSYS_UNCONNECTED__493, 
        SYNOPSYS_UNCONNECTED__494, SYNOPSYS_UNCONNECTED__495, 
        SYNOPSYS_UNCONNECTED__496, SYNOPSYS_UNCONNECTED__497, 
        SYNOPSYS_UNCONNECTED__498, SYNOPSYS_UNCONNECTED__499, 
        SYNOPSYS_UNCONNECTED__500, SYNOPSYS_UNCONNECTED__501, 
        SYNOPSYS_UNCONNECTED__502, SYNOPSYS_UNCONNECTED__503, 
        SYNOPSYS_UNCONNECTED__504, SYNOPSYS_UNCONNECTED__505, 
        SYNOPSYS_UNCONNECTED__506, SYNOPSYS_UNCONNECTED__507, 
        SYNOPSYS_UNCONNECTED__508, SYNOPSYS_UNCONNECTED__509, 
        SYNOPSYS_UNCONNECTED__510, SYNOPSYS_UNCONNECTED__511, 
        SYNOPSYS_UNCONNECTED__512, SYNOPSYS_UNCONNECTED__513, 
        SYNOPSYS_UNCONNECTED__514, SYNOPSYS_UNCONNECTED__515, 
        SYNOPSYS_UNCONNECTED__516, SYNOPSYS_UNCONNECTED__517, 
        SYNOPSYS_UNCONNECTED__518, SYNOPSYS_UNCONNECTED__519, 
        SYNOPSYS_UNCONNECTED__520, SYNOPSYS_UNCONNECTED__521, 
        SYNOPSYS_UNCONNECTED__522, SYNOPSYS_UNCONNECTED__523, 
        SYNOPSYS_UNCONNECTED__524, SYNOPSYS_UNCONNECTED__525, 
        SYNOPSYS_UNCONNECTED__526, SYNOPSYS_UNCONNECTED__527, 
        SYNOPSYS_UNCONNECTED__528, SYNOPSYS_UNCONNECTED__529, 
        SYNOPSYS_UNCONNECTED__530, SYNOPSYS_UNCONNECTED__531, 
        SYNOPSYS_UNCONNECTED__532, SYNOPSYS_UNCONNECTED__533, 
        SYNOPSYS_UNCONNECTED__534, SYNOPSYS_UNCONNECTED__535, 
        SYNOPSYS_UNCONNECTED__536, SYNOPSYS_UNCONNECTED__537, 
        SYNOPSYS_UNCONNECTED__538, SYNOPSYS_UNCONNECTED__539, 
        SYNOPSYS_UNCONNECTED__540, SYNOPSYS_UNCONNECTED__541, 
        SYNOPSYS_UNCONNECTED__542, SYNOPSYS_UNCONNECTED__543, 
        SYNOPSYS_UNCONNECTED__544, SYNOPSYS_UNCONNECTED__545, 
        SYNOPSYS_UNCONNECTED__546, SYNOPSYS_UNCONNECTED__547, 
        SYNOPSYS_UNCONNECTED__548, SYNOPSYS_UNCONNECTED__549, 
        SYNOPSYS_UNCONNECTED__550, SYNOPSYS_UNCONNECTED__551, 
        SYNOPSYS_UNCONNECTED__552, SYNOPSYS_UNCONNECTED__553, 
        SYNOPSYS_UNCONNECTED__554, SYNOPSYS_UNCONNECTED__555, 
        SYNOPSYS_UNCONNECTED__556, SYNOPSYS_UNCONNECTED__557, 
        SYNOPSYS_UNCONNECTED__558, SYNOPSYS_UNCONNECTED__559, 
        SYNOPSYS_UNCONNECTED__560, SYNOPSYS_UNCONNECTED__561, 
        SYNOPSYS_UNCONNECTED__562, SYNOPSYS_UNCONNECTED__563, 
        SYNOPSYS_UNCONNECTED__564, SYNOPSYS_UNCONNECTED__565, 
        SYNOPSYS_UNCONNECTED__566, SYNOPSYS_UNCONNECTED__567, 
        SYNOPSYS_UNCONNECTED__568, SYNOPSYS_UNCONNECTED__569, 
        SYNOPSYS_UNCONNECTED__570, SYNOPSYS_UNCONNECTED__571, 
        SYNOPSYS_UNCONNECTED__572, SYNOPSYS_UNCONNECTED__573, 
        SYNOPSYS_UNCONNECTED__574, SYNOPSYS_UNCONNECTED__575, 
        SYNOPSYS_UNCONNECTED__576, SYNOPSYS_UNCONNECTED__577, 
        SYNOPSYS_UNCONNECTED__578, SYNOPSYS_UNCONNECTED__579, 
        SYNOPSYS_UNCONNECTED__580, SYNOPSYS_UNCONNECTED__581, 
        SYNOPSYS_UNCONNECTED__582, SYNOPSYS_UNCONNECTED__583, 
        SYNOPSYS_UNCONNECTED__584, SYNOPSYS_UNCONNECTED__585, 
        SYNOPSYS_UNCONNECTED__586, SYNOPSYS_UNCONNECTED__587, 
        SYNOPSYS_UNCONNECTED__588, SYNOPSYS_UNCONNECTED__589, 
        SYNOPSYS_UNCONNECTED__590, SYNOPSYS_UNCONNECTED__591, 
        SYNOPSYS_UNCONNECTED__592, SYNOPSYS_UNCONNECTED__593, 
        SYNOPSYS_UNCONNECTED__594, SYNOPSYS_UNCONNECTED__595, 
        SYNOPSYS_UNCONNECTED__596, SYNOPSYS_UNCONNECTED__597, 
        SYNOPSYS_UNCONNECTED__598, SYNOPSYS_UNCONNECTED__599, 
        SYNOPSYS_UNCONNECTED__600, SYNOPSYS_UNCONNECTED__601, 
        SYNOPSYS_UNCONNECTED__602, SYNOPSYS_UNCONNECTED__603, 
        SYNOPSYS_UNCONNECTED__604, SYNOPSYS_UNCONNECTED__605, 
        SYNOPSYS_UNCONNECTED__606, SYNOPSYS_UNCONNECTED__607, 
        SYNOPSYS_UNCONNECTED__608, SYNOPSYS_UNCONNECTED__609, 
        SYNOPSYS_UNCONNECTED__610, SYNOPSYS_UNCONNECTED__611, 
        SYNOPSYS_UNCONNECTED__612, SYNOPSYS_UNCONNECTED__613, 
        SYNOPSYS_UNCONNECTED__614, SYNOPSYS_UNCONNECTED__615, 
        SYNOPSYS_UNCONNECTED__616, SYNOPSYS_UNCONNECTED__617, 
        SYNOPSYS_UNCONNECTED__618, SYNOPSYS_UNCONNECTED__619, 
        SYNOPSYS_UNCONNECTED__620, SYNOPSYS_UNCONNECTED__621, 
        SYNOPSYS_UNCONNECTED__622, SYNOPSYS_UNCONNECTED__623, 
        SYNOPSYS_UNCONNECTED__624, SYNOPSYS_UNCONNECTED__625, 
        SYNOPSYS_UNCONNECTED__626, SYNOPSYS_UNCONNECTED__627, 
        SYNOPSYS_UNCONNECTED__628, SYNOPSYS_UNCONNECTED__629, 
        SYNOPSYS_UNCONNECTED__630, SYNOPSYS_UNCONNECTED__631, 
        SYNOPSYS_UNCONNECTED__632, SYNOPSYS_UNCONNECTED__633, 
        SYNOPSYS_UNCONNECTED__634, SYNOPSYS_UNCONNECTED__635, 
        SYNOPSYS_UNCONNECTED__636, SYNOPSYS_UNCONNECTED__637, 
        SYNOPSYS_UNCONNECTED__638, SYNOPSYS_UNCONNECTED__639, 
        SYNOPSYS_UNCONNECTED__640, SYNOPSYS_UNCONNECTED__641, 
        SYNOPSYS_UNCONNECTED__642, SYNOPSYS_UNCONNECTED__643, 
        SYNOPSYS_UNCONNECTED__644, SYNOPSYS_UNCONNECTED__645, 
        SYNOPSYS_UNCONNECTED__646, SYNOPSYS_UNCONNECTED__647, 
        SYNOPSYS_UNCONNECTED__648, SYNOPSYS_UNCONNECTED__649, 
        SYNOPSYS_UNCONNECTED__650, SYNOPSYS_UNCONNECTED__651, 
        SYNOPSYS_UNCONNECTED__652, SYNOPSYS_UNCONNECTED__653, 
        SYNOPSYS_UNCONNECTED__654, SYNOPSYS_UNCONNECTED__655, 
        SYNOPSYS_UNCONNECTED__656, SYNOPSYS_UNCONNECTED__657, 
        SYNOPSYS_UNCONNECTED__658, SYNOPSYS_UNCONNECTED__659, 
        SYNOPSYS_UNCONNECTED__660, SYNOPSYS_UNCONNECTED__661, 
        SYNOPSYS_UNCONNECTED__662, SYNOPSYS_UNCONNECTED__663, 
        SYNOPSYS_UNCONNECTED__664, SYNOPSYS_UNCONNECTED__665, 
        SYNOPSYS_UNCONNECTED__666, SYNOPSYS_UNCONNECTED__667, 
        SYNOPSYS_UNCONNECTED__668, SYNOPSYS_UNCONNECTED__669, 
        SYNOPSYS_UNCONNECTED__670, SYNOPSYS_UNCONNECTED__671, 
        SYNOPSYS_UNCONNECTED__672, SYNOPSYS_UNCONNECTED__673, 
        SYNOPSYS_UNCONNECTED__674, SYNOPSYS_UNCONNECTED__675, 
        SYNOPSYS_UNCONNECTED__676, SYNOPSYS_UNCONNECTED__677, 
        SYNOPSYS_UNCONNECTED__678, SYNOPSYS_UNCONNECTED__679, 
        SYNOPSYS_UNCONNECTED__680, SYNOPSYS_UNCONNECTED__681, 
        SYNOPSYS_UNCONNECTED__682, SYNOPSYS_UNCONNECTED__683, 
        SYNOPSYS_UNCONNECTED__684, SYNOPSYS_UNCONNECTED__685, 
        SYNOPSYS_UNCONNECTED__686, SYNOPSYS_UNCONNECTED__687, 
        SYNOPSYS_UNCONNECTED__688, SYNOPSYS_UNCONNECTED__689, 
        SYNOPSYS_UNCONNECTED__690, SYNOPSYS_UNCONNECTED__691, 
        SYNOPSYS_UNCONNECTED__692, SYNOPSYS_UNCONNECTED__693, 
        SYNOPSYS_UNCONNECTED__694, SYNOPSYS_UNCONNECTED__695, 
        SYNOPSYS_UNCONNECTED__696, SYNOPSYS_UNCONNECTED__697, 
        SYNOPSYS_UNCONNECTED__698, SYNOPSYS_UNCONNECTED__699, 
        SYNOPSYS_UNCONNECTED__700, SYNOPSYS_UNCONNECTED__701, 
        SYNOPSYS_UNCONNECTED__702, SYNOPSYS_UNCONNECTED__703, 
        SYNOPSYS_UNCONNECTED__704, SYNOPSYS_UNCONNECTED__705, 
        SYNOPSYS_UNCONNECTED__706, SYNOPSYS_UNCONNECTED__707, 
        SYNOPSYS_UNCONNECTED__708, SYNOPSYS_UNCONNECTED__709, 
        SYNOPSYS_UNCONNECTED__710, SYNOPSYS_UNCONNECTED__711, 
        SYNOPSYS_UNCONNECTED__712, SYNOPSYS_UNCONNECTED__713, 
        SYNOPSYS_UNCONNECTED__714, SYNOPSYS_UNCONNECTED__715, 
        SYNOPSYS_UNCONNECTED__716, SYNOPSYS_UNCONNECTED__717, 
        SYNOPSYS_UNCONNECTED__718, SYNOPSYS_UNCONNECTED__719, 
        SYNOPSYS_UNCONNECTED__720, SYNOPSYS_UNCONNECTED__721, 
        SYNOPSYS_UNCONNECTED__722, SYNOPSYS_UNCONNECTED__723, 
        SYNOPSYS_UNCONNECTED__724, SYNOPSYS_UNCONNECTED__725, 
        SYNOPSYS_UNCONNECTED__726, SYNOPSYS_UNCONNECTED__727, 
        SYNOPSYS_UNCONNECTED__728, SYNOPSYS_UNCONNECTED__729, 
        SYNOPSYS_UNCONNECTED__730, SYNOPSYS_UNCONNECTED__731, 
        SYNOPSYS_UNCONNECTED__732, SYNOPSYS_UNCONNECTED__733, 
        SYNOPSYS_UNCONNECTED__734, SYNOPSYS_UNCONNECTED__735, 
        SYNOPSYS_UNCONNECTED__736, SYNOPSYS_UNCONNECTED__737, 
        SYNOPSYS_UNCONNECTED__738, SYNOPSYS_UNCONNECTED__739, 
        SYNOPSYS_UNCONNECTED__740, SYNOPSYS_UNCONNECTED__741, 
        SYNOPSYS_UNCONNECTED__742, SYNOPSYS_UNCONNECTED__743, 
        SYNOPSYS_UNCONNECTED__744, SYNOPSYS_UNCONNECTED__745, 
        SYNOPSYS_UNCONNECTED__746, SYNOPSYS_UNCONNECTED__747, 
        SYNOPSYS_UNCONNECTED__748, SYNOPSYS_UNCONNECTED__749, 
        SYNOPSYS_UNCONNECTED__750, SYNOPSYS_UNCONNECTED__751, 
        SYNOPSYS_UNCONNECTED__752, SYNOPSYS_UNCONNECTED__753, 
        SYNOPSYS_UNCONNECTED__754, SYNOPSYS_UNCONNECTED__755, 
        SYNOPSYS_UNCONNECTED__756, SYNOPSYS_UNCONNECTED__757, 
        SYNOPSYS_UNCONNECTED__758, SYNOPSYS_UNCONNECTED__759, 
        SYNOPSYS_UNCONNECTED__760, SYNOPSYS_UNCONNECTED__761, 
        SYNOPSYS_UNCONNECTED__762, SYNOPSYS_UNCONNECTED__763, 
        SYNOPSYS_UNCONNECTED__764, SYNOPSYS_UNCONNECTED__765, 
        SYNOPSYS_UNCONNECTED__766, SYNOPSYS_UNCONNECTED__767, 
        SYNOPSYS_UNCONNECTED__768, SYNOPSYS_UNCONNECTED__769, 
        SYNOPSYS_UNCONNECTED__770, SYNOPSYS_UNCONNECTED__771, 
        SYNOPSYS_UNCONNECTED__772, SYNOPSYS_UNCONNECTED__773, 
        SYNOPSYS_UNCONNECTED__774, SYNOPSYS_UNCONNECTED__775, 
        SYNOPSYS_UNCONNECTED__776, SYNOPSYS_UNCONNECTED__777, 
        SYNOPSYS_UNCONNECTED__778, SYNOPSYS_UNCONNECTED__779, 
        SYNOPSYS_UNCONNECTED__780, SYNOPSYS_UNCONNECTED__781, 
        SYNOPSYS_UNCONNECTED__782, SYNOPSYS_UNCONNECTED__783, 
        SYNOPSYS_UNCONNECTED__784, SYNOPSYS_UNCONNECTED__785, 
        SYNOPSYS_UNCONNECTED__786, SYNOPSYS_UNCONNECTED__787, 
        SYNOPSYS_UNCONNECTED__788, SYNOPSYS_UNCONNECTED__789, 
        SYNOPSYS_UNCONNECTED__790, SYNOPSYS_UNCONNECTED__791, 
        SYNOPSYS_UNCONNECTED__792, SYNOPSYS_UNCONNECTED__793, 
        SYNOPSYS_UNCONNECTED__794, SYNOPSYS_UNCONNECTED__795, 
        SYNOPSYS_UNCONNECTED__796, SYNOPSYS_UNCONNECTED__797, 
        SYNOPSYS_UNCONNECTED__798, SYNOPSYS_UNCONNECTED__799, 
        SYNOPSYS_UNCONNECTED__800, SYNOPSYS_UNCONNECTED__801, 
        SYNOPSYS_UNCONNECTED__802, SYNOPSYS_UNCONNECTED__803, 
        SYNOPSYS_UNCONNECTED__804, SYNOPSYS_UNCONNECTED__805, 
        SYNOPSYS_UNCONNECTED__806, SYNOPSYS_UNCONNECTED__807, 
        SYNOPSYS_UNCONNECTED__808, SYNOPSYS_UNCONNECTED__809, 
        SYNOPSYS_UNCONNECTED__810, SYNOPSYS_UNCONNECTED__811, 
        SYNOPSYS_UNCONNECTED__812, SYNOPSYS_UNCONNECTED__813, 
        SYNOPSYS_UNCONNECTED__814, SYNOPSYS_UNCONNECTED__815, 
        SYNOPSYS_UNCONNECTED__816, SYNOPSYS_UNCONNECTED__817, 
        SYNOPSYS_UNCONNECTED__818, SYNOPSYS_UNCONNECTED__819, 
        SYNOPSYS_UNCONNECTED__820, SYNOPSYS_UNCONNECTED__821, 
        SYNOPSYS_UNCONNECTED__822, SYNOPSYS_UNCONNECTED__823, 
        SYNOPSYS_UNCONNECTED__824, SYNOPSYS_UNCONNECTED__825, 
        SYNOPSYS_UNCONNECTED__826, SYNOPSYS_UNCONNECTED__827, 
        SYNOPSYS_UNCONNECTED__828, SYNOPSYS_UNCONNECTED__829, 
        SYNOPSYS_UNCONNECTED__830, SYNOPSYS_UNCONNECTED__831, 
        SYNOPSYS_UNCONNECTED__832, SYNOPSYS_UNCONNECTED__833, 
        SYNOPSYS_UNCONNECTED__834;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  hamming_N16000_CC4_DW01_add_0 add_97 ( .A(oglobal), .B({1'b0, 1'b0, olocal}), 
        .CI(1'b0), .SUM(o) );
  hamming_N16000_CC4_DW01_add_1 add_1334_root_add_71_I928 ( .A({1'b0, N31899, 
        N31898, N31897, N31896, N31895, N31894, N31893, N31892, N31891, N31890, 
        N31889}), .B({N31912, N31911, N31910, N31909, N31908, N31907, N31906, 
        N31905, N31904, N31903, N31902, N31901}), .CI(1'b0), .SUM(olocal) );
  hamming_N16000_CC4_DW01_add_2 add_1335_root_add_71_I928 ( .A({1'b0, N31875, 
        N31874, N31873, N31872, N31871, N31870, N31869, N31868, N31867, N31866, 
        N31865}), .B({1'b0, N31887, N31886, N31885, N31884, N31883, N31882, 
        N31881, N31880, N31879, N31878, N31877}), .CI(1'b0), .SUM({N31912, 
        N31911, N31910, N31909, N31908, N31907, N31906, N31905, N31904, N31903, 
        N31902, N31901}) );
  hamming_N16000_CC4_DW01_add_3 add_1336_root_add_71_I928 ( .A({1'b0, 1'b0, 
        N31850, N31849, N31848, N31847, N31846, N31845, N31844, N31843, N31842, 
        N31841}), .B({1'b0, 1'b0, N31862, N31861, N31860, N31859, N31858, 
        N31857, N31856, N31855, N31854, N31853}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, N31899, N31898, N31897, N31896, N31895, 
        N31894, N31893, N31892, N31891, N31890, N31889}) );
  hamming_N16000_CC4_DW01_add_4 add_1337_root_add_71_I928 ( .A({1'b0, 1'b0, 
        N31826, N31825, N31824, N31823, N31822, N31821, N31820, N31819, N31818, 
        N31817}), .B({1'b0, 1'b0, N31838, N31837, N31836, N31835, N31834, 
        N31833, N31832, N31831, N31830, N31829}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1, N31887, N31886, N31885, N31884, N31883, 
        N31882, N31881, N31880, N31879, N31878, N31877}) );
  hamming_N16000_CC4_DW01_add_5 add_1338_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, N31801, N31800, N31799, N31798, N31797, N31796, N31795, N31794, 
        N31793}), .B({1'b0, 1'b0, N31814, N31813, N31812, N31811, N31810, 
        N31809, N31808, N31807, N31806, N31805}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__2, N31875, N31874, N31873, N31872, N31871, 
        N31870, N31869, N31868, N31867, N31866, N31865}) );
  hamming_N16000_CC4_DW01_add_6 add_1339_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, N31777, N31776, N31775, N31774, N31773, N31772, N31771, N31770, 
        N31769}), .B({1'b0, 1'b0, 1'b0, N31789, N31788, N31787, N31786, N31785, 
        N31784, N31783, N31782, N31781}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, N31862, N31861, 
        N31860, N31859, N31858, N31857, N31856, N31855, N31854, N31853}) );
  hamming_N16000_CC4_DW01_add_7 add_1340_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, N31753, N31752, N31751, N31750, N31749, N31748, N31747, N31746, 
        N31745}), .B({1'b0, 1'b0, 1'b0, N31765, N31764, N31763, N31762, N31761, 
        N31760, N31759, N31758, N31757}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, N31850, N31849, 
        N31848, N31847, N31846, N31845, N31844, N31843, N31842, N31841}) );
  hamming_N16000_CC4_DW01_add_8 add_1341_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, N31729, N31728, N31727, N31726, N31725, N31724, N31723, N31722, 
        N31721}), .B({1'b0, 1'b0, 1'b0, N31741, N31740, N31739, N31738, N31737, 
        N31736, N31735, N31734, N31733}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, N31838, N31837, 
        N31836, N31835, N31834, N31833, N31832, N31831, N31830, N31829}) );
  hamming_N16000_CC4_DW01_add_9 add_1342_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, N31705, N31704, N31703, N31702, N31701, N31700, N31699, N31698, 
        N31697}), .B({1'b0, 1'b0, 1'b0, N31717, N31716, N31715, N31714, N31713, 
        N31712, N31711, N31710, N31709}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, N31826, N31825, 
        N31824, N31823, N31822, N31821, N31820, N31819, N31818, N31817}) );
  hamming_N16000_CC4_DW01_add_10 add_1343_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31680, N31679, N31678, N31677, N31676, N31675, N31674, 
        N31673}), .B({1'b0, 1'b0, 1'b0, N31693, N31692, N31691, N31690, N31689, 
        N31688, N31687, N31686, N31685}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, N31814, N31813, 
        N31812, N31811, N31810, N31809, N31808, N31807, N31806, N31805}) );
  hamming_N16000_CC4_DW01_add_11 add_1344_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31656, N31655, N31654, N31653, N31652, N31651, N31650, 
        N31649}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31668, N31667, N31666, N31665, 
        N31664, N31663, N31662, N31661}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N31801, N31800, N31799, N31798, N31797, 
        N31796, N31795, N31794, N31793}) );
  hamming_N16000_CC4_DW01_add_12 add_1345_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31632, N31631, N31630, N31629, N31628, N31627, N31626, 
        N31625}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31644, N31643, N31642, N31641, 
        N31640, N31639, N31638, N31637}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, N31789, N31788, N31787, N31786, N31785, 
        N31784, N31783, N31782, N31781}) );
  hamming_N16000_CC4_DW01_add_13 add_1346_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31608, N31607, N31606, N31605, N31604, N31603, N31602, 
        N31601}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31620, N31619, N31618, N31617, 
        N31616, N31615, N31614, N31613}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, N31777, N31776, N31775, N31774, N31773, 
        N31772, N31771, N31770, N31769}) );
  hamming_N16000_CC4_DW01_add_14 add_1347_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31584, N31583, N31582, N31581, N31580, N31579, N31578, 
        N31577}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31596, N31595, N31594, N31593, 
        N31592, N31591, N31590, N31589}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, N31765, N31764, N31763, N31762, N31761, 
        N31760, N31759, N31758, N31757}) );
  hamming_N16000_CC4_DW01_add_15 add_1348_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31560, N31559, N31558, N31557, N31556, N31555, N31554, 
        N31553}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31572, N31571, N31570, N31569, 
        N31568, N31567, N31566, N31565}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, N31753, N31752, N31751, N31750, N31749, 
        N31748, N31747, N31746, N31745}) );
  hamming_N16000_CC4_DW01_add_16 add_1349_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31536, N31535, N31534, N31533, N31532, N31531, N31530, 
        N31529}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31548, N31547, N31546, N31545, 
        N31544, N31543, N31542, N31541}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, N31741, N31740, N31739, N31738, N31737, 
        N31736, N31735, N31734, N31733}) );
  hamming_N16000_CC4_DW01_add_17 add_1350_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31512, N31511, N31510, N31509, N31508, N31507, N31506, 
        N31505}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31524, N31523, N31522, N31521, 
        N31520, N31519, N31518, N31517}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, N31729, N31728, N31727, N31726, N31725, 
        N31724, N31723, N31722, N31721}) );
  hamming_N16000_CC4_DW01_add_18 add_1351_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31488, N31487, N31486, N31485, N31484, N31483, N31482, 
        N31481}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31500, N31499, N31498, N31497, 
        N31496, N31495, N31494, N31493}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, N31717, N31716, N31715, N31714, N31713, 
        N31712, N31711, N31710, N31709}) );
  hamming_N16000_CC4_DW01_add_19 add_1352_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31464, N31463, N31462, N31461, N31460, N31459, N31458, 
        N31457}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31476, N31475, N31474, N31473, 
        N31472, N31471, N31470, N31469}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, N31705, N31704, N31703, N31702, N31701, 
        N31700, N31699, N31698, N31697}) );
  hamming_N16000_CC4_DW01_add_20 add_1353_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N31440, N31439, N31438, N31437, N31436, N31435, N31434, 
        N31433}), .B({1'b0, 1'b0, 1'b0, 1'b0, N31452, N31451, N31450, N31449, 
        N31448, N31447, N31446, N31445}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, N31693, N31692, N31691, N31690, N31689, 
        N31688, N31687, N31686, N31685}) );
  hamming_N16000_CC4_DW01_add_21 add_1354_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31415, N31414, N31413, N31412, N31411, N31410, 
        N31409}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31427, N31426, N31425, 
        N31424, N31423, N31422, N31421}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, N31680, N31679, 
        N31678, N31677, N31676, N31675, N31674, N31673}) );
  hamming_N16000_CC4_DW01_add_22 add_1355_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31391, N31390, N31389, N31388, N31387, N31386, 
        N31385}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31403, N31402, N31401, 
        N31400, N31399, N31398, N31397}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, N31668, N31667, 
        N31666, N31665, N31664, N31663, N31662, N31661}) );
  hamming_N16000_CC4_DW01_add_23 add_1356_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31367, N31366, N31365, N31364, N31363, N31362, 
        N31361}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31379, N31378, N31377, 
        N31376, N31375, N31374, N31373}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, N31656, N31655, 
        N31654, N31653, N31652, N31651, N31650, N31649}) );
  hamming_N16000_CC4_DW01_add_24 add_1357_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31343, N31342, N31341, N31340, N31339, N31338, 
        N31337}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31355, N31354, N31353, 
        N31352, N31351, N31350, N31349}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, N31644, N31643, 
        N31642, N31641, N31640, N31639, N31638, N31637}) );
  hamming_N16000_CC4_DW01_add_25 add_1358_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31319, N31318, N31317, N31316, N31315, N31314, 
        N31313}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31331, N31330, N31329, 
        N31328, N31327, N31326, N31325}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, N31632, N31631, 
        N31630, N31629, N31628, N31627, N31626, N31625}) );
  hamming_N16000_CC4_DW01_add_26 add_1359_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31295, N31294, N31293, N31292, N31291, N31290, 
        N31289}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31307, N31306, N31305, 
        N31304, N31303, N31302, N31301}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, N31620, N31619, 
        N31618, N31617, N31616, N31615, N31614, N31613}) );
  hamming_N16000_CC4_DW01_add_27 add_1360_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31271, N31270, N31269, N31268, N31267, N31266, 
        N31265}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31283, N31282, N31281, 
        N31280, N31279, N31278, N31277}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, N31608, N31607, 
        N31606, N31605, N31604, N31603, N31602, N31601}) );
  hamming_N16000_CC4_DW01_add_28 add_1361_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31247, N31246, N31245, N31244, N31243, N31242, 
        N31241}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31259, N31258, N31257, 
        N31256, N31255, N31254, N31253}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, N31596, N31595, 
        N31594, N31593, N31592, N31591, N31590, N31589}) );
  hamming_N16000_CC4_DW01_add_29 add_1362_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31223, N31222, N31221, N31220, N31219, N31218, 
        N31217}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31235, N31234, N31233, 
        N31232, N31231, N31230, N31229}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, N31584, N31583, 
        N31582, N31581, N31580, N31579, N31578, N31577}) );
  hamming_N16000_CC4_DW01_add_30 add_1363_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31199, N31198, N31197, N31196, N31195, N31194, 
        N31193}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31211, N31210, N31209, 
        N31208, N31207, N31206, N31205}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, N31572, N31571, 
        N31570, N31569, N31568, N31567, N31566, N31565}) );
  hamming_N16000_CC4_DW01_add_31 add_1364_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31175, N31174, N31173, N31172, N31171, N31170, 
        N31169}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31187, N31186, N31185, 
        N31184, N31183, N31182, N31181}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, N31560, N31559, 
        N31558, N31557, N31556, N31555, N31554, N31553}) );
  hamming_N16000_CC4_DW01_add_32 add_1365_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31151, N31150, N31149, N31148, N31147, N31146, 
        N31145}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31163, N31162, N31161, 
        N31160, N31159, N31158, N31157}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, N31548, N31547, 
        N31546, N31545, N31544, N31543, N31542, N31541}) );
  hamming_N16000_CC4_DW01_add_33 add_1366_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31127, N31126, N31125, N31124, N31123, N31122, 
        N31121}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31139, N31138, N31137, 
        N31136, N31135, N31134, N31133}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, N31536, N31535, 
        N31534, N31533, N31532, N31531, N31530, N31529}) );
  hamming_N16000_CC4_DW01_add_34 add_1367_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31103, N31102, N31101, N31100, N31099, N31098, 
        N31097}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31115, N31114, N31113, 
        N31112, N31111, N31110, N31109}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, N31524, N31523, 
        N31522, N31521, N31520, N31519, N31518, N31517}) );
  hamming_N16000_CC4_DW01_add_35 add_1368_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31079, N31078, N31077, N31076, N31075, N31074, 
        N31073}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31091, N31090, N31089, 
        N31088, N31087, N31086, N31085}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, N31512, N31511, 
        N31510, N31509, N31508, N31507, N31506, N31505}) );
  hamming_N16000_CC4_DW01_add_36 add_1369_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31055, N31054, N31053, N31052, N31051, N31050, 
        N31049}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31067, N31066, N31065, 
        N31064, N31063, N31062, N31061}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, N31500, N31499, 
        N31498, N31497, N31496, N31495, N31494, N31493}) );
  hamming_N16000_CC4_DW01_add_37 add_1370_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31031, N31030, N31029, N31028, N31027, N31026, 
        N31025}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31043, N31042, N31041, 
        N31040, N31039, N31038, N31037}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, N31488, N31487, 
        N31486, N31485, N31484, N31483, N31482, N31481}) );
  hamming_N16000_CC4_DW01_add_38 add_1371_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N31007, N31006, N31005, N31004, N31003, N31002, 
        N31001}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N31019, N31018, N31017, 
        N31016, N31015, N31014, N31013}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, N31476, N31475, 
        N31474, N31473, N31472, N31471, N31470, N31469}) );
  hamming_N16000_CC4_DW01_add_39 add_1372_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N30983, N30982, N30981, N30980, N30979, N30978, 
        N30977}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30995, N30994, N30993, 
        N30992, N30991, N30990, N30989}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, N31464, N31463, 
        N31462, N31461, N31460, N31459, N31458, N31457}) );
  hamming_N16000_CC4_DW01_add_40 add_1373_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N30959, N30958, N30957, N30956, N30955, N30954, 
        N30953}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30971, N30970, N30969, 
        N30968, N30967, N30966, N30965}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, N31452, N31451, 
        N31450, N31449, N31448, N31447, N31446, N31445}) );
  hamming_N16000_CC4_DW01_add_41 add_1374_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N30935, N30934, N30933, N30932, N30931, N30930, 
        N30929}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30947, N30946, N30945, 
        N30944, N30943, N30942, N30941}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, N31440, N31439, 
        N31438, N31437, N31436, N31435, N31434, N31433}) );
  hamming_N16000_CC4_DW01_add_42 add_1375_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30910, N30909, N30908, N30907, N30906, N30905}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30922, N30921, N30920, N30919, 
        N30918, N30917}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, N31427, N31426, 
        N31425, N31424, N31423, N31422, N31421}) );
  hamming_N16000_CC4_DW01_add_43 add_1376_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30886, N30885, N30884, N30883, N30882, N30881}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30898, N30897, N30896, N30895, 
        N30894, N30893}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, N31415, N31414, 
        N31413, N31412, N31411, N31410, N31409}) );
  hamming_N16000_CC4_DW01_add_44 add_1377_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30862, N30861, N30860, N30859, N30858, N30857}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30874, N30873, N30872, N30871, 
        N30870, N30869}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, N31403, N31402, 
        N31401, N31400, N31399, N31398, N31397}) );
  hamming_N16000_CC4_DW01_add_45 add_1378_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30838, N30837, N30836, N30835, N30834, N30833}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30850, N30849, N30848, N30847, 
        N30846, N30845}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__142, 
        SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, N31391, N31390, 
        N31389, N31388, N31387, N31386, N31385}) );
  hamming_N16000_CC4_DW01_add_46 add_1379_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30814, N30813, N30812, N30811, N30810, N30809}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30826, N30825, N30824, N30823, 
        N30822, N30821}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, N31379, N31378, 
        N31377, N31376, N31375, N31374, N31373}) );
  hamming_N16000_CC4_DW01_add_47 add_1380_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30790, N30789, N30788, N30787, N30786, N30785}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30802, N30801, N30800, N30799, 
        N30798, N30797}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__152, 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, N31367, N31366, 
        N31365, N31364, N31363, N31362, N31361}) );
  hamming_N16000_CC4_DW01_add_48 add_1381_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30766, N30765, N30764, N30763, N30762, N30761}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30778, N30777, N30776, N30775, 
        N30774, N30773}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, N31355, N31354, 
        N31353, N31352, N31351, N31350, N31349}) );
  hamming_N16000_CC4_DW01_add_49 add_1382_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30742, N30741, N30740, N30739, N30738, N30737}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30754, N30753, N30752, N30751, 
        N30750, N30749}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, N31343, N31342, 
        N31341, N31340, N31339, N31338, N31337}) );
  hamming_N16000_CC4_DW01_add_50 add_1383_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30718, N30717, N30716, N30715, N30714, N30713}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30730, N30729, N30728, N30727, 
        N30726, N30725}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, N31331, N31330, 
        N31329, N31328, N31327, N31326, N31325}) );
  hamming_N16000_CC4_DW01_add_51 add_1384_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30694, N30693, N30692, N30691, N30690, N30689}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30706, N30705, N30704, N30703, 
        N30702, N30701}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__172, 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, N31319, N31318, 
        N31317, N31316, N31315, N31314, N31313}) );
  hamming_N16000_CC4_DW01_add_52 add_1385_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30670, N30669, N30668, N30667, N30666, N30665}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30682, N30681, N30680, N30679, 
        N30678, N30677}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, N31307, N31306, 
        N31305, N31304, N31303, N31302, N31301}) );
  hamming_N16000_CC4_DW01_add_53 add_1386_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30646, N30645, N30644, N30643, N30642, N30641}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30658, N30657, N30656, N30655, 
        N30654, N30653}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__182, 
        SYNOPSYS_UNCONNECTED__183, SYNOPSYS_UNCONNECTED__184, 
        SYNOPSYS_UNCONNECTED__185, SYNOPSYS_UNCONNECTED__186, N31295, N31294, 
        N31293, N31292, N31291, N31290, N31289}) );
  hamming_N16000_CC4_DW01_add_54 add_1387_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30622, N30621, N30620, N30619, N30618, N30617}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30634, N30633, N30632, N30631, 
        N30630, N30629}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, N31283, N31282, 
        N31281, N31280, N31279, N31278, N31277}) );
  hamming_N16000_CC4_DW01_add_55 add_1388_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30598, N30597, N30596, N30595, N30594, N30593}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30610, N30609, N30608, N30607, 
        N30606, N30605}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__192, 
        SYNOPSYS_UNCONNECTED__193, SYNOPSYS_UNCONNECTED__194, 
        SYNOPSYS_UNCONNECTED__195, SYNOPSYS_UNCONNECTED__196, N31271, N31270, 
        N31269, N31268, N31267, N31266, N31265}) );
  hamming_N16000_CC4_DW01_add_56 add_1389_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30574, N30573, N30572, N30571, N30570, N30569}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30586, N30585, N30584, N30583, 
        N30582, N30581}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, N31259, N31258, 
        N31257, N31256, N31255, N31254, N31253}) );
  hamming_N16000_CC4_DW01_add_57 add_1390_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30550, N30549, N30548, N30547, N30546, N30545}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30562, N30561, N30560, N30559, 
        N30558, N30557}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__202, 
        SYNOPSYS_UNCONNECTED__203, SYNOPSYS_UNCONNECTED__204, 
        SYNOPSYS_UNCONNECTED__205, SYNOPSYS_UNCONNECTED__206, N31247, N31246, 
        N31245, N31244, N31243, N31242, N31241}) );
  hamming_N16000_CC4_DW01_add_58 add_1391_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30526, N30525, N30524, N30523, N30522, N30521}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30538, N30537, N30536, N30535, 
        N30534, N30533}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, N31235, N31234, 
        N31233, N31232, N31231, N31230, N31229}) );
  hamming_N16000_CC4_DW01_add_59 add_1392_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30502, N30501, N30500, N30499, N30498, N30497}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30514, N30513, N30512, N30511, 
        N30510, N30509}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__212, 
        SYNOPSYS_UNCONNECTED__213, SYNOPSYS_UNCONNECTED__214, 
        SYNOPSYS_UNCONNECTED__215, SYNOPSYS_UNCONNECTED__216, N31223, N31222, 
        N31221, N31220, N31219, N31218, N31217}) );
  hamming_N16000_CC4_DW01_add_60 add_1393_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30478, N30477, N30476, N30475, N30474, N30473}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30490, N30489, N30488, N30487, 
        N30486, N30485}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, N31211, N31210, 
        N31209, N31208, N31207, N31206, N31205}) );
  hamming_N16000_CC4_DW01_add_61 add_1394_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30454, N30453, N30452, N30451, N30450, N30449}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30466, N30465, N30464, N30463, 
        N30462, N30461}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__222, 
        SYNOPSYS_UNCONNECTED__223, SYNOPSYS_UNCONNECTED__224, 
        SYNOPSYS_UNCONNECTED__225, SYNOPSYS_UNCONNECTED__226, N31199, N31198, 
        N31197, N31196, N31195, N31194, N31193}) );
  hamming_N16000_CC4_DW01_add_62 add_1395_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30430, N30429, N30428, N30427, N30426, N30425}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30442, N30441, N30440, N30439, 
        N30438, N30437}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, N31187, N31186, 
        N31185, N31184, N31183, N31182, N31181}) );
  hamming_N16000_CC4_DW01_add_63 add_1396_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30406, N30405, N30404, N30403, N30402, N30401}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30418, N30417, N30416, N30415, 
        N30414, N30413}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__232, 
        SYNOPSYS_UNCONNECTED__233, SYNOPSYS_UNCONNECTED__234, 
        SYNOPSYS_UNCONNECTED__235, SYNOPSYS_UNCONNECTED__236, N31175, N31174, 
        N31173, N31172, N31171, N31170, N31169}) );
  hamming_N16000_CC4_DW01_add_64 add_1397_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30382, N30381, N30380, N30379, N30378, N30377}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30394, N30393, N30392, N30391, 
        N30390, N30389}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, N31163, N31162, 
        N31161, N31160, N31159, N31158, N31157}) );
  hamming_N16000_CC4_DW01_add_65 add_1398_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30358, N30357, N30356, N30355, N30354, N30353}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30370, N30369, N30368, N30367, 
        N30366, N30365}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__242, 
        SYNOPSYS_UNCONNECTED__243, SYNOPSYS_UNCONNECTED__244, 
        SYNOPSYS_UNCONNECTED__245, SYNOPSYS_UNCONNECTED__246, N31151, N31150, 
        N31149, N31148, N31147, N31146, N31145}) );
  hamming_N16000_CC4_DW01_add_66 add_1399_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30334, N30333, N30332, N30331, N30330, N30329}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30346, N30345, N30344, N30343, 
        N30342, N30341}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, N31139, N31138, 
        N31137, N31136, N31135, N31134, N31133}) );
  hamming_N16000_CC4_DW01_add_67 add_1400_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30310, N30309, N30308, N30307, N30306, N30305}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30322, N30321, N30320, N30319, 
        N30318, N30317}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__252, 
        SYNOPSYS_UNCONNECTED__253, SYNOPSYS_UNCONNECTED__254, 
        SYNOPSYS_UNCONNECTED__255, SYNOPSYS_UNCONNECTED__256, N31127, N31126, 
        N31125, N31124, N31123, N31122, N31121}) );
  hamming_N16000_CC4_DW01_add_68 add_1401_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30286, N30285, N30284, N30283, N30282, N30281}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30298, N30297, N30296, N30295, 
        N30294, N30293}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, N31115, N31114, 
        N31113, N31112, N31111, N31110, N31109}) );
  hamming_N16000_CC4_DW01_add_69 add_1402_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30262, N30261, N30260, N30259, N30258, N30257}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30274, N30273, N30272, N30271, 
        N30270, N30269}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__262, 
        SYNOPSYS_UNCONNECTED__263, SYNOPSYS_UNCONNECTED__264, 
        SYNOPSYS_UNCONNECTED__265, SYNOPSYS_UNCONNECTED__266, N31103, N31102, 
        N31101, N31100, N31099, N31098, N31097}) );
  hamming_N16000_CC4_DW01_add_70 add_1403_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30238, N30237, N30236, N30235, N30234, N30233}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30250, N30249, N30248, N30247, 
        N30246, N30245}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, N31091, N31090, 
        N31089, N31088, N31087, N31086, N31085}) );
  hamming_N16000_CC4_DW01_add_71 add_1404_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30214, N30213, N30212, N30211, N30210, N30209}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30226, N30225, N30224, N30223, 
        N30222, N30221}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__272, 
        SYNOPSYS_UNCONNECTED__273, SYNOPSYS_UNCONNECTED__274, 
        SYNOPSYS_UNCONNECTED__275, SYNOPSYS_UNCONNECTED__276, N31079, N31078, 
        N31077, N31076, N31075, N31074, N31073}) );
  hamming_N16000_CC4_DW01_add_72 add_1405_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30190, N30189, N30188, N30187, N30186, N30185}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30202, N30201, N30200, N30199, 
        N30198, N30197}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, N31067, N31066, 
        N31065, N31064, N31063, N31062, N31061}) );
  hamming_N16000_CC4_DW01_add_73 add_1406_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30166, N30165, N30164, N30163, N30162, N30161}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30178, N30177, N30176, N30175, 
        N30174, N30173}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__282, 
        SYNOPSYS_UNCONNECTED__283, SYNOPSYS_UNCONNECTED__284, 
        SYNOPSYS_UNCONNECTED__285, SYNOPSYS_UNCONNECTED__286, N31055, N31054, 
        N31053, N31052, N31051, N31050, N31049}) );
  hamming_N16000_CC4_DW01_add_74 add_1407_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30142, N30141, N30140, N30139, N30138, N30137}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30154, N30153, N30152, N30151, 
        N30150, N30149}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, N31043, N31042, 
        N31041, N31040, N31039, N31038, N31037}) );
  hamming_N16000_CC4_DW01_add_75 add_1408_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30118, N30117, N30116, N30115, N30114, N30113}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30130, N30129, N30128, N30127, 
        N30126, N30125}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__292, 
        SYNOPSYS_UNCONNECTED__293, SYNOPSYS_UNCONNECTED__294, 
        SYNOPSYS_UNCONNECTED__295, SYNOPSYS_UNCONNECTED__296, N31031, N31030, 
        N31029, N31028, N31027, N31026, N31025}) );
  hamming_N16000_CC4_DW01_add_76 add_1409_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30094, N30093, N30092, N30091, N30090, N30089}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30106, N30105, N30104, N30103, 
        N30102, N30101}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, N31019, N31018, 
        N31017, N31016, N31015, N31014, N31013}) );
  hamming_N16000_CC4_DW01_add_77 add_1410_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30070, N30069, N30068, N30067, N30066, N30065}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30082, N30081, N30080, N30079, 
        N30078, N30077}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__302, 
        SYNOPSYS_UNCONNECTED__303, SYNOPSYS_UNCONNECTED__304, 
        SYNOPSYS_UNCONNECTED__305, SYNOPSYS_UNCONNECTED__306, N31007, N31006, 
        N31005, N31004, N31003, N31002, N31001}) );
  hamming_N16000_CC4_DW01_add_78 add_1411_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30046, N30045, N30044, N30043, N30042, N30041}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30058, N30057, N30056, N30055, 
        N30054, N30053}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, N30995, N30994, 
        N30993, N30992, N30991, N30990, N30989}) );
  hamming_N16000_CC4_DW01_add_79 add_1412_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N30022, N30021, N30020, N30019, N30018, N30017}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30034, N30033, N30032, N30031, 
        N30030, N30029}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__312, 
        SYNOPSYS_UNCONNECTED__313, SYNOPSYS_UNCONNECTED__314, 
        SYNOPSYS_UNCONNECTED__315, SYNOPSYS_UNCONNECTED__316, N30983, N30982, 
        N30981, N30980, N30979, N30978, N30977}) );
  hamming_N16000_CC4_DW01_add_80 add_1413_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N29998, N29997, N29996, N29995, N29994, N29993}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N30010, N30009, N30008, N30007, 
        N30006, N30005}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, N30971, N30970, 
        N30969, N30968, N30967, N30966, N30965}) );
  hamming_N16000_CC4_DW01_add_81 add_1414_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N29974, N29973, N29972, N29971, N29970, N29969}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29986, N29985, N29984, N29983, 
        N29982, N29981}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__322, 
        SYNOPSYS_UNCONNECTED__323, SYNOPSYS_UNCONNECTED__324, 
        SYNOPSYS_UNCONNECTED__325, SYNOPSYS_UNCONNECTED__326, N30959, N30958, 
        N30957, N30956, N30955, N30954, N30953}) );
  hamming_N16000_CC4_DW01_add_82 add_1415_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N29950, N29949, N29948, N29947, N29946, N29945}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29962, N29961, N29960, N29959, 
        N29958, N29957}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, N30947, N30946, 
        N30945, N30944, N30943, N30942, N30941}) );
  hamming_N16000_CC4_DW01_add_83 add_1416_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29925, N29924, N29923, N29922, N29921}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29938, N29937, N29936, N29935, 
        N29934, N29933}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__332, 
        SYNOPSYS_UNCONNECTED__333, SYNOPSYS_UNCONNECTED__334, 
        SYNOPSYS_UNCONNECTED__335, SYNOPSYS_UNCONNECTED__336, N30935, N30934, 
        N30933, N30932, N30931, N30930, N30929}) );
  hamming_N16000_CC4_DW01_add_84 add_1417_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29901, N29900, N29899, N29898, N29897}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29913, N29912, N29911, 
        N29910, N29909}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, N30922, N30921, N30920, N30919, N30918, 
        N30917}) );
  hamming_N16000_CC4_DW01_add_85 add_1418_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29877, N29876, N29875, N29874, N29873}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29889, N29888, N29887, 
        N29886, N29885}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, N30910, N30909, N30908, N30907, N30906, 
        N30905}) );
  hamming_N16000_CC4_DW01_add_86 add_1419_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29853, N29852, N29851, N29850, N29849}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29865, N29864, N29863, 
        N29862, N29861}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        SYNOPSYS_UNCONNECTED__352, SYNOPSYS_UNCONNECTED__353, 
        SYNOPSYS_UNCONNECTED__354, N30898, N30897, N30896, N30895, N30894, 
        N30893}) );
  hamming_N16000_CC4_DW01_add_87 add_1420_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29829, N29828, N29827, N29826, N29825}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29841, N29840, N29839, 
        N29838, N29837}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__355, 
        SYNOPSYS_UNCONNECTED__356, SYNOPSYS_UNCONNECTED__357, 
        SYNOPSYS_UNCONNECTED__358, SYNOPSYS_UNCONNECTED__359, 
        SYNOPSYS_UNCONNECTED__360, N30886, N30885, N30884, N30883, N30882, 
        N30881}) );
  hamming_N16000_CC4_DW01_add_88 add_1421_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29805, N29804, N29803, N29802, N29801}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29817, N29816, N29815, 
        N29814, N29813}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__361, 
        SYNOPSYS_UNCONNECTED__362, SYNOPSYS_UNCONNECTED__363, 
        SYNOPSYS_UNCONNECTED__364, SYNOPSYS_UNCONNECTED__365, 
        SYNOPSYS_UNCONNECTED__366, N30874, N30873, N30872, N30871, N30870, 
        N30869}) );
  hamming_N16000_CC4_DW01_add_89 add_1422_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29781, N29780, N29779, N29778, N29777}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29793, N29792, N29791, 
        N29790, N29789}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__367, 
        SYNOPSYS_UNCONNECTED__368, SYNOPSYS_UNCONNECTED__369, 
        SYNOPSYS_UNCONNECTED__370, SYNOPSYS_UNCONNECTED__371, 
        SYNOPSYS_UNCONNECTED__372, N30862, N30861, N30860, N30859, N30858, 
        N30857}) );
  hamming_N16000_CC4_DW01_add_90 add_1423_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29757, N29756, N29755, N29754, N29753}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29769, N29768, N29767, 
        N29766, N29765}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__373, 
        SYNOPSYS_UNCONNECTED__374, SYNOPSYS_UNCONNECTED__375, 
        SYNOPSYS_UNCONNECTED__376, SYNOPSYS_UNCONNECTED__377, 
        SYNOPSYS_UNCONNECTED__378, N30850, N30849, N30848, N30847, N30846, 
        N30845}) );
  hamming_N16000_CC4_DW01_add_91 add_1424_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29733, N29732, N29731, N29730, N29729}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29745, N29744, N29743, 
        N29742, N29741}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__379, 
        SYNOPSYS_UNCONNECTED__380, SYNOPSYS_UNCONNECTED__381, 
        SYNOPSYS_UNCONNECTED__382, SYNOPSYS_UNCONNECTED__383, 
        SYNOPSYS_UNCONNECTED__384, N30838, N30837, N30836, N30835, N30834, 
        N30833}) );
  hamming_N16000_CC4_DW01_add_92 add_1425_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29709, N29708, N29707, N29706, N29705}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29721, N29720, N29719, 
        N29718, N29717}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__385, 
        SYNOPSYS_UNCONNECTED__386, SYNOPSYS_UNCONNECTED__387, 
        SYNOPSYS_UNCONNECTED__388, SYNOPSYS_UNCONNECTED__389, 
        SYNOPSYS_UNCONNECTED__390, N30826, N30825, N30824, N30823, N30822, 
        N30821}) );
  hamming_N16000_CC4_DW01_add_93 add_1426_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29685, N29684, N29683, N29682, N29681}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29697, N29696, N29695, 
        N29694, N29693}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__391, 
        SYNOPSYS_UNCONNECTED__392, SYNOPSYS_UNCONNECTED__393, 
        SYNOPSYS_UNCONNECTED__394, SYNOPSYS_UNCONNECTED__395, 
        SYNOPSYS_UNCONNECTED__396, N30814, N30813, N30812, N30811, N30810, 
        N30809}) );
  hamming_N16000_CC4_DW01_add_94 add_1427_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29661, N29660, N29659, N29658, N29657}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29673, N29672, N29671, 
        N29670, N29669}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__397, 
        SYNOPSYS_UNCONNECTED__398, SYNOPSYS_UNCONNECTED__399, 
        SYNOPSYS_UNCONNECTED__400, SYNOPSYS_UNCONNECTED__401, 
        SYNOPSYS_UNCONNECTED__402, N30802, N30801, N30800, N30799, N30798, 
        N30797}) );
  hamming_N16000_CC4_DW01_add_95 add_1428_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29637, N29636, N29635, N29634, N29633}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29649, N29648, N29647, 
        N29646, N29645}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__403, 
        SYNOPSYS_UNCONNECTED__404, SYNOPSYS_UNCONNECTED__405, 
        SYNOPSYS_UNCONNECTED__406, SYNOPSYS_UNCONNECTED__407, 
        SYNOPSYS_UNCONNECTED__408, N30790, N30789, N30788, N30787, N30786, 
        N30785}) );
  hamming_N16000_CC4_DW01_add_96 add_1429_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29613, N29612, N29611, N29610, N29609}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29625, N29624, N29623, 
        N29622, N29621}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__409, 
        SYNOPSYS_UNCONNECTED__410, SYNOPSYS_UNCONNECTED__411, 
        SYNOPSYS_UNCONNECTED__412, SYNOPSYS_UNCONNECTED__413, 
        SYNOPSYS_UNCONNECTED__414, N30778, N30777, N30776, N30775, N30774, 
        N30773}) );
  hamming_N16000_CC4_DW01_add_97 add_1430_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29589, N29588, N29587, N29586, N29585}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29601, N29600, N29599, 
        N29598, N29597}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__415, 
        SYNOPSYS_UNCONNECTED__416, SYNOPSYS_UNCONNECTED__417, 
        SYNOPSYS_UNCONNECTED__418, SYNOPSYS_UNCONNECTED__419, 
        SYNOPSYS_UNCONNECTED__420, N30766, N30765, N30764, N30763, N30762, 
        N30761}) );
  hamming_N16000_CC4_DW01_add_98 add_1431_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29565, N29564, N29563, N29562, N29561}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29577, N29576, N29575, 
        N29574, N29573}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__421, 
        SYNOPSYS_UNCONNECTED__422, SYNOPSYS_UNCONNECTED__423, 
        SYNOPSYS_UNCONNECTED__424, SYNOPSYS_UNCONNECTED__425, 
        SYNOPSYS_UNCONNECTED__426, N30754, N30753, N30752, N30751, N30750, 
        N30749}) );
  hamming_N16000_CC4_DW01_add_99 add_1432_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29541, N29540, N29539, N29538, N29537}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29553, N29552, N29551, 
        N29550, N29549}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__427, 
        SYNOPSYS_UNCONNECTED__428, SYNOPSYS_UNCONNECTED__429, 
        SYNOPSYS_UNCONNECTED__430, SYNOPSYS_UNCONNECTED__431, 
        SYNOPSYS_UNCONNECTED__432, N30742, N30741, N30740, N30739, N30738, 
        N30737}) );
  hamming_N16000_CC4_DW01_add_100 add_1433_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29517, N29516, N29515, N29514, N29513}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29529, N29528, N29527, 
        N29526, N29525}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__433, 
        SYNOPSYS_UNCONNECTED__434, SYNOPSYS_UNCONNECTED__435, 
        SYNOPSYS_UNCONNECTED__436, SYNOPSYS_UNCONNECTED__437, 
        SYNOPSYS_UNCONNECTED__438, N30730, N30729, N30728, N30727, N30726, 
        N30725}) );
  hamming_N16000_CC4_DW01_add_101 add_1434_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29493, N29492, N29491, N29490, N29489}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29505, N29504, N29503, 
        N29502, N29501}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__439, 
        SYNOPSYS_UNCONNECTED__440, SYNOPSYS_UNCONNECTED__441, 
        SYNOPSYS_UNCONNECTED__442, SYNOPSYS_UNCONNECTED__443, 
        SYNOPSYS_UNCONNECTED__444, N30718, N30717, N30716, N30715, N30714, 
        N30713}) );
  hamming_N16000_CC4_DW01_add_102 add_1435_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29469, N29468, N29467, N29466, N29465}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29481, N29480, N29479, 
        N29478, N29477}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__445, 
        SYNOPSYS_UNCONNECTED__446, SYNOPSYS_UNCONNECTED__447, 
        SYNOPSYS_UNCONNECTED__448, SYNOPSYS_UNCONNECTED__449, 
        SYNOPSYS_UNCONNECTED__450, N30706, N30705, N30704, N30703, N30702, 
        N30701}) );
  hamming_N16000_CC4_DW01_add_103 add_1436_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29445, N29444, N29443, N29442, N29441}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29457, N29456, N29455, 
        N29454, N29453}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__451, 
        SYNOPSYS_UNCONNECTED__452, SYNOPSYS_UNCONNECTED__453, 
        SYNOPSYS_UNCONNECTED__454, SYNOPSYS_UNCONNECTED__455, 
        SYNOPSYS_UNCONNECTED__456, N30694, N30693, N30692, N30691, N30690, 
        N30689}) );
  hamming_N16000_CC4_DW01_add_104 add_1437_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29421, N29420, N29419, N29418, N29417}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29433, N29432, N29431, 
        N29430, N29429}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__457, 
        SYNOPSYS_UNCONNECTED__458, SYNOPSYS_UNCONNECTED__459, 
        SYNOPSYS_UNCONNECTED__460, SYNOPSYS_UNCONNECTED__461, 
        SYNOPSYS_UNCONNECTED__462, N30682, N30681, N30680, N30679, N30678, 
        N30677}) );
  hamming_N16000_CC4_DW01_add_105 add_1438_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29397, N29396, N29395, N29394, N29393}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29409, N29408, N29407, 
        N29406, N29405}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__463, 
        SYNOPSYS_UNCONNECTED__464, SYNOPSYS_UNCONNECTED__465, 
        SYNOPSYS_UNCONNECTED__466, SYNOPSYS_UNCONNECTED__467, 
        SYNOPSYS_UNCONNECTED__468, N30670, N30669, N30668, N30667, N30666, 
        N30665}) );
  hamming_N16000_CC4_DW01_add_106 add_1439_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29373, N29372, N29371, N29370, N29369}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29385, N29384, N29383, 
        N29382, N29381}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__469, 
        SYNOPSYS_UNCONNECTED__470, SYNOPSYS_UNCONNECTED__471, 
        SYNOPSYS_UNCONNECTED__472, SYNOPSYS_UNCONNECTED__473, 
        SYNOPSYS_UNCONNECTED__474, N30658, N30657, N30656, N30655, N30654, 
        N30653}) );
  hamming_N16000_CC4_DW01_add_107 add_1440_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29349, N29348, N29347, N29346, N29345}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29361, N29360, N29359, 
        N29358, N29357}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__475, 
        SYNOPSYS_UNCONNECTED__476, SYNOPSYS_UNCONNECTED__477, 
        SYNOPSYS_UNCONNECTED__478, SYNOPSYS_UNCONNECTED__479, 
        SYNOPSYS_UNCONNECTED__480, N30646, N30645, N30644, N30643, N30642, 
        N30641}) );
  hamming_N16000_CC4_DW01_add_108 add_1441_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29325, N29324, N29323, N29322, N29321}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29337, N29336, N29335, 
        N29334, N29333}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__481, 
        SYNOPSYS_UNCONNECTED__482, SYNOPSYS_UNCONNECTED__483, 
        SYNOPSYS_UNCONNECTED__484, SYNOPSYS_UNCONNECTED__485, 
        SYNOPSYS_UNCONNECTED__486, N30634, N30633, N30632, N30631, N30630, 
        N30629}) );
  hamming_N16000_CC4_DW01_add_109 add_1442_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29301, N29300, N29299, N29298, N29297}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29313, N29312, N29311, 
        N29310, N29309}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__487, 
        SYNOPSYS_UNCONNECTED__488, SYNOPSYS_UNCONNECTED__489, 
        SYNOPSYS_UNCONNECTED__490, SYNOPSYS_UNCONNECTED__491, 
        SYNOPSYS_UNCONNECTED__492, N30622, N30621, N30620, N30619, N30618, 
        N30617}) );
  hamming_N16000_CC4_DW01_add_110 add_1443_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29277, N29276, N29275, N29274, N29273}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29289, N29288, N29287, 
        N29286, N29285}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__493, 
        SYNOPSYS_UNCONNECTED__494, SYNOPSYS_UNCONNECTED__495, 
        SYNOPSYS_UNCONNECTED__496, SYNOPSYS_UNCONNECTED__497, 
        SYNOPSYS_UNCONNECTED__498, N30610, N30609, N30608, N30607, N30606, 
        N30605}) );
  hamming_N16000_CC4_DW01_add_111 add_1444_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29253, N29252, N29251, N29250, N29249}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29265, N29264, N29263, 
        N29262, N29261}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__499, 
        SYNOPSYS_UNCONNECTED__500, SYNOPSYS_UNCONNECTED__501, 
        SYNOPSYS_UNCONNECTED__502, SYNOPSYS_UNCONNECTED__503, 
        SYNOPSYS_UNCONNECTED__504, N30598, N30597, N30596, N30595, N30594, 
        N30593}) );
  hamming_N16000_CC4_DW01_add_112 add_1445_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29229, N29228, N29227, N29226, N29225}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29241, N29240, N29239, 
        N29238, N29237}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__505, 
        SYNOPSYS_UNCONNECTED__506, SYNOPSYS_UNCONNECTED__507, 
        SYNOPSYS_UNCONNECTED__508, SYNOPSYS_UNCONNECTED__509, 
        SYNOPSYS_UNCONNECTED__510, N30586, N30585, N30584, N30583, N30582, 
        N30581}) );
  hamming_N16000_CC4_DW01_add_113 add_1446_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29205, N29204, N29203, N29202, N29201}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29217, N29216, N29215, 
        N29214, N29213}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__511, 
        SYNOPSYS_UNCONNECTED__512, SYNOPSYS_UNCONNECTED__513, 
        SYNOPSYS_UNCONNECTED__514, SYNOPSYS_UNCONNECTED__515, 
        SYNOPSYS_UNCONNECTED__516, N30574, N30573, N30572, N30571, N30570, 
        N30569}) );
  hamming_N16000_CC4_DW01_add_114 add_1447_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29181, N29180, N29179, N29178, N29177}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29193, N29192, N29191, 
        N29190, N29189}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__517, 
        SYNOPSYS_UNCONNECTED__518, SYNOPSYS_UNCONNECTED__519, 
        SYNOPSYS_UNCONNECTED__520, SYNOPSYS_UNCONNECTED__521, 
        SYNOPSYS_UNCONNECTED__522, N30562, N30561, N30560, N30559, N30558, 
        N30557}) );
  hamming_N16000_CC4_DW01_add_115 add_1448_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29157, N29156, N29155, N29154, N29153}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29169, N29168, N29167, 
        N29166, N29165}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__523, 
        SYNOPSYS_UNCONNECTED__524, SYNOPSYS_UNCONNECTED__525, 
        SYNOPSYS_UNCONNECTED__526, SYNOPSYS_UNCONNECTED__527, 
        SYNOPSYS_UNCONNECTED__528, N30550, N30549, N30548, N30547, N30546, 
        N30545}) );
  hamming_N16000_CC4_DW01_add_116 add_1449_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29133, N29132, N29131, N29130, N29129}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29145, N29144, N29143, 
        N29142, N29141}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__529, 
        SYNOPSYS_UNCONNECTED__530, SYNOPSYS_UNCONNECTED__531, 
        SYNOPSYS_UNCONNECTED__532, SYNOPSYS_UNCONNECTED__533, 
        SYNOPSYS_UNCONNECTED__534, N30538, N30537, N30536, N30535, N30534, 
        N30533}) );
  hamming_N16000_CC4_DW01_add_117 add_1450_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29109, N29108, N29107, N29106, N29105}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29121, N29120, N29119, 
        N29118, N29117}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__535, 
        SYNOPSYS_UNCONNECTED__536, SYNOPSYS_UNCONNECTED__537, 
        SYNOPSYS_UNCONNECTED__538, SYNOPSYS_UNCONNECTED__539, 
        SYNOPSYS_UNCONNECTED__540, N30526, N30525, N30524, N30523, N30522, 
        N30521}) );
  hamming_N16000_CC4_DW01_add_118 add_1451_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29085, N29084, N29083, N29082, N29081}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29097, N29096, N29095, 
        N29094, N29093}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__541, 
        SYNOPSYS_UNCONNECTED__542, SYNOPSYS_UNCONNECTED__543, 
        SYNOPSYS_UNCONNECTED__544, SYNOPSYS_UNCONNECTED__545, 
        SYNOPSYS_UNCONNECTED__546, N30514, N30513, N30512, N30511, N30510, 
        N30509}) );
  hamming_N16000_CC4_DW01_add_119 add_1452_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29061, N29060, N29059, N29058, N29057}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29073, N29072, N29071, 
        N29070, N29069}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__547, 
        SYNOPSYS_UNCONNECTED__548, SYNOPSYS_UNCONNECTED__549, 
        SYNOPSYS_UNCONNECTED__550, SYNOPSYS_UNCONNECTED__551, 
        SYNOPSYS_UNCONNECTED__552, N30502, N30501, N30500, N30499, N30498, 
        N30497}) );
  hamming_N16000_CC4_DW01_add_120 add_1453_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29037, N29036, N29035, N29034, N29033}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29049, N29048, N29047, 
        N29046, N29045}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__553, 
        SYNOPSYS_UNCONNECTED__554, SYNOPSYS_UNCONNECTED__555, 
        SYNOPSYS_UNCONNECTED__556, SYNOPSYS_UNCONNECTED__557, 
        SYNOPSYS_UNCONNECTED__558, N30490, N30489, N30488, N30487, N30486, 
        N30485}) );
  hamming_N16000_CC4_DW01_add_121 add_1454_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29013, N29012, N29011, N29010, N29009}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29025, N29024, N29023, 
        N29022, N29021}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__559, 
        SYNOPSYS_UNCONNECTED__560, SYNOPSYS_UNCONNECTED__561, 
        SYNOPSYS_UNCONNECTED__562, SYNOPSYS_UNCONNECTED__563, 
        SYNOPSYS_UNCONNECTED__564, N30478, N30477, N30476, N30475, N30474, 
        N30473}) );
  hamming_N16000_CC4_DW01_add_122 add_1455_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28989, N28988, N28987, N28986, N28985}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N29001, N29000, N28999, 
        N28998, N28997}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__565, 
        SYNOPSYS_UNCONNECTED__566, SYNOPSYS_UNCONNECTED__567, 
        SYNOPSYS_UNCONNECTED__568, SYNOPSYS_UNCONNECTED__569, 
        SYNOPSYS_UNCONNECTED__570, N30466, N30465, N30464, N30463, N30462, 
        N30461}) );
  hamming_N16000_CC4_DW01_add_123 add_1456_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28965, N28964, N28963, N28962, N28961}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28977, N28976, N28975, 
        N28974, N28973}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__571, 
        SYNOPSYS_UNCONNECTED__572, SYNOPSYS_UNCONNECTED__573, 
        SYNOPSYS_UNCONNECTED__574, SYNOPSYS_UNCONNECTED__575, 
        SYNOPSYS_UNCONNECTED__576, N30454, N30453, N30452, N30451, N30450, 
        N30449}) );
  hamming_N16000_CC4_DW01_add_124 add_1457_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28941, N28940, N28939, N28938, N28937}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28953, N28952, N28951, 
        N28950, N28949}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__577, 
        SYNOPSYS_UNCONNECTED__578, SYNOPSYS_UNCONNECTED__579, 
        SYNOPSYS_UNCONNECTED__580, SYNOPSYS_UNCONNECTED__581, 
        SYNOPSYS_UNCONNECTED__582, N30442, N30441, N30440, N30439, N30438, 
        N30437}) );
  hamming_N16000_CC4_DW01_add_125 add_1458_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28917, N28916, N28915, N28914, N28913}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28929, N28928, N28927, 
        N28926, N28925}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__583, 
        SYNOPSYS_UNCONNECTED__584, SYNOPSYS_UNCONNECTED__585, 
        SYNOPSYS_UNCONNECTED__586, SYNOPSYS_UNCONNECTED__587, 
        SYNOPSYS_UNCONNECTED__588, N30430, N30429, N30428, N30427, N30426, 
        N30425}) );
  hamming_N16000_CC4_DW01_add_126 add_1459_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28893, N28892, N28891, N28890, N28889}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28905, N28904, N28903, 
        N28902, N28901}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__589, 
        SYNOPSYS_UNCONNECTED__590, SYNOPSYS_UNCONNECTED__591, 
        SYNOPSYS_UNCONNECTED__592, SYNOPSYS_UNCONNECTED__593, 
        SYNOPSYS_UNCONNECTED__594, N30418, N30417, N30416, N30415, N30414, 
        N30413}) );
  hamming_N16000_CC4_DW01_add_127 add_1460_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28869, N28868, N28867, N28866, N28865}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28881, N28880, N28879, 
        N28878, N28877}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__595, 
        SYNOPSYS_UNCONNECTED__596, SYNOPSYS_UNCONNECTED__597, 
        SYNOPSYS_UNCONNECTED__598, SYNOPSYS_UNCONNECTED__599, 
        SYNOPSYS_UNCONNECTED__600, N30406, N30405, N30404, N30403, N30402, 
        N30401}) );
  hamming_N16000_CC4_DW01_add_128 add_1461_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28845, N28844, N28843, N28842, N28841}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28857, N28856, N28855, 
        N28854, N28853}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__601, 
        SYNOPSYS_UNCONNECTED__602, SYNOPSYS_UNCONNECTED__603, 
        SYNOPSYS_UNCONNECTED__604, SYNOPSYS_UNCONNECTED__605, 
        SYNOPSYS_UNCONNECTED__606, N30394, N30393, N30392, N30391, N30390, 
        N30389}) );
  hamming_N16000_CC4_DW01_add_129 add_1462_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28821, N28820, N28819, N28818, N28817}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28833, N28832, N28831, 
        N28830, N28829}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__607, 
        SYNOPSYS_UNCONNECTED__608, SYNOPSYS_UNCONNECTED__609, 
        SYNOPSYS_UNCONNECTED__610, SYNOPSYS_UNCONNECTED__611, 
        SYNOPSYS_UNCONNECTED__612, N30382, N30381, N30380, N30379, N30378, 
        N30377}) );
  hamming_N16000_CC4_DW01_add_130 add_1463_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28797, N28796, N28795, N28794, N28793}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28809, N28808, N28807, 
        N28806, N28805}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__613, 
        SYNOPSYS_UNCONNECTED__614, SYNOPSYS_UNCONNECTED__615, 
        SYNOPSYS_UNCONNECTED__616, SYNOPSYS_UNCONNECTED__617, 
        SYNOPSYS_UNCONNECTED__618, N30370, N30369, N30368, N30367, N30366, 
        N30365}) );
  hamming_N16000_CC4_DW01_add_131 add_1464_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28773, N28772, N28771, N28770, N28769}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28785, N28784, N28783, 
        N28782, N28781}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__619, 
        SYNOPSYS_UNCONNECTED__620, SYNOPSYS_UNCONNECTED__621, 
        SYNOPSYS_UNCONNECTED__622, SYNOPSYS_UNCONNECTED__623, 
        SYNOPSYS_UNCONNECTED__624, N30358, N30357, N30356, N30355, N30354, 
        N30353}) );
  hamming_N16000_CC4_DW01_add_132 add_1465_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28749, N28748, N28747, N28746, N28745}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28761, N28760, N28759, 
        N28758, N28757}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__625, 
        SYNOPSYS_UNCONNECTED__626, SYNOPSYS_UNCONNECTED__627, 
        SYNOPSYS_UNCONNECTED__628, SYNOPSYS_UNCONNECTED__629, 
        SYNOPSYS_UNCONNECTED__630, N30346, N30345, N30344, N30343, N30342, 
        N30341}) );
  hamming_N16000_CC4_DW01_add_133 add_1466_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28725, N28724, N28723, N28722, N28721}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28737, N28736, N28735, 
        N28734, N28733}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__631, 
        SYNOPSYS_UNCONNECTED__632, SYNOPSYS_UNCONNECTED__633, 
        SYNOPSYS_UNCONNECTED__634, SYNOPSYS_UNCONNECTED__635, 
        SYNOPSYS_UNCONNECTED__636, N30334, N30333, N30332, N30331, N30330, 
        N30329}) );
  hamming_N16000_CC4_DW01_add_134 add_1467_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28701, N28700, N28699, N28698, N28697}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28713, N28712, N28711, 
        N28710, N28709}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__637, 
        SYNOPSYS_UNCONNECTED__638, SYNOPSYS_UNCONNECTED__639, 
        SYNOPSYS_UNCONNECTED__640, SYNOPSYS_UNCONNECTED__641, 
        SYNOPSYS_UNCONNECTED__642, N30322, N30321, N30320, N30319, N30318, 
        N30317}) );
  hamming_N16000_CC4_DW01_add_135 add_1468_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28677, N28676, N28675, N28674, N28673}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28689, N28688, N28687, 
        N28686, N28685}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__643, 
        SYNOPSYS_UNCONNECTED__644, SYNOPSYS_UNCONNECTED__645, 
        SYNOPSYS_UNCONNECTED__646, SYNOPSYS_UNCONNECTED__647, 
        SYNOPSYS_UNCONNECTED__648, N30310, N30309, N30308, N30307, N30306, 
        N30305}) );
  hamming_N16000_CC4_DW01_add_136 add_1469_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28653, N28652, N28651, N28650, N28649}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28665, N28664, N28663, 
        N28662, N28661}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__649, 
        SYNOPSYS_UNCONNECTED__650, SYNOPSYS_UNCONNECTED__651, 
        SYNOPSYS_UNCONNECTED__652, SYNOPSYS_UNCONNECTED__653, 
        SYNOPSYS_UNCONNECTED__654, N30298, N30297, N30296, N30295, N30294, 
        N30293}) );
  hamming_N16000_CC4_DW01_add_137 add_1470_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28629, N28628, N28627, N28626, N28625}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28641, N28640, N28639, 
        N28638, N28637}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__655, 
        SYNOPSYS_UNCONNECTED__656, SYNOPSYS_UNCONNECTED__657, 
        SYNOPSYS_UNCONNECTED__658, SYNOPSYS_UNCONNECTED__659, 
        SYNOPSYS_UNCONNECTED__660, N30286, N30285, N30284, N30283, N30282, 
        N30281}) );
  hamming_N16000_CC4_DW01_add_138 add_1471_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28605, N28604, N28603, N28602, N28601}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28617, N28616, N28615, 
        N28614, N28613}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__661, 
        SYNOPSYS_UNCONNECTED__662, SYNOPSYS_UNCONNECTED__663, 
        SYNOPSYS_UNCONNECTED__664, SYNOPSYS_UNCONNECTED__665, 
        SYNOPSYS_UNCONNECTED__666, N30274, N30273, N30272, N30271, N30270, 
        N30269}) );
  hamming_N16000_CC4_DW01_add_139 add_1472_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28581, N28580, N28579, N28578, N28577}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28593, N28592, N28591, 
        N28590, N28589}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__667, 
        SYNOPSYS_UNCONNECTED__668, SYNOPSYS_UNCONNECTED__669, 
        SYNOPSYS_UNCONNECTED__670, SYNOPSYS_UNCONNECTED__671, 
        SYNOPSYS_UNCONNECTED__672, N30262, N30261, N30260, N30259, N30258, 
        N30257}) );
  hamming_N16000_CC4_DW01_add_140 add_1473_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28557, N28556, N28555, N28554, N28553}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28569, N28568, N28567, 
        N28566, N28565}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__673, 
        SYNOPSYS_UNCONNECTED__674, SYNOPSYS_UNCONNECTED__675, 
        SYNOPSYS_UNCONNECTED__676, SYNOPSYS_UNCONNECTED__677, 
        SYNOPSYS_UNCONNECTED__678, N30250, N30249, N30248, N30247, N30246, 
        N30245}) );
  hamming_N16000_CC4_DW01_add_141 add_1474_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28533, N28532, N28531, N28530, N28529}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28545, N28544, N28543, 
        N28542, N28541}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__679, 
        SYNOPSYS_UNCONNECTED__680, SYNOPSYS_UNCONNECTED__681, 
        SYNOPSYS_UNCONNECTED__682, SYNOPSYS_UNCONNECTED__683, 
        SYNOPSYS_UNCONNECTED__684, N30238, N30237, N30236, N30235, N30234, 
        N30233}) );
  hamming_N16000_CC4_DW01_add_142 add_1475_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28509, N28508, N28507, N28506, N28505}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28521, N28520, N28519, 
        N28518, N28517}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__685, 
        SYNOPSYS_UNCONNECTED__686, SYNOPSYS_UNCONNECTED__687, 
        SYNOPSYS_UNCONNECTED__688, SYNOPSYS_UNCONNECTED__689, 
        SYNOPSYS_UNCONNECTED__690, N30226, N30225, N30224, N30223, N30222, 
        N30221}) );
  hamming_N16000_CC4_DW01_add_143 add_1476_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28485, N28484, N28483, N28482, N28481}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28497, N28496, N28495, 
        N28494, N28493}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__691, 
        SYNOPSYS_UNCONNECTED__692, SYNOPSYS_UNCONNECTED__693, 
        SYNOPSYS_UNCONNECTED__694, SYNOPSYS_UNCONNECTED__695, 
        SYNOPSYS_UNCONNECTED__696, N30214, N30213, N30212, N30211, N30210, 
        N30209}) );
  hamming_N16000_CC4_DW01_add_144 add_1477_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28461, N28460, N28459, N28458, N28457}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28473, N28472, N28471, 
        N28470, N28469}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__697, 
        SYNOPSYS_UNCONNECTED__698, SYNOPSYS_UNCONNECTED__699, 
        SYNOPSYS_UNCONNECTED__700, SYNOPSYS_UNCONNECTED__701, 
        SYNOPSYS_UNCONNECTED__702, N30202, N30201, N30200, N30199, N30198, 
        N30197}) );
  hamming_N16000_CC4_DW01_add_145 add_1478_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28437, N28436, N28435, N28434, N28433}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28449, N28448, N28447, 
        N28446, N28445}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__703, 
        SYNOPSYS_UNCONNECTED__704, SYNOPSYS_UNCONNECTED__705, 
        SYNOPSYS_UNCONNECTED__706, SYNOPSYS_UNCONNECTED__707, 
        SYNOPSYS_UNCONNECTED__708, N30190, N30189, N30188, N30187, N30186, 
        N30185}) );
  hamming_N16000_CC4_DW01_add_146 add_1479_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28413, N28412, N28411, N28410, N28409}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28425, N28424, N28423, 
        N28422, N28421}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__709, 
        SYNOPSYS_UNCONNECTED__710, SYNOPSYS_UNCONNECTED__711, 
        SYNOPSYS_UNCONNECTED__712, SYNOPSYS_UNCONNECTED__713, 
        SYNOPSYS_UNCONNECTED__714, N30178, N30177, N30176, N30175, N30174, 
        N30173}) );
  hamming_N16000_CC4_DW01_add_147 add_1480_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28389, N28388, N28387, N28386, N28385}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28401, N28400, N28399, 
        N28398, N28397}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__715, 
        SYNOPSYS_UNCONNECTED__716, SYNOPSYS_UNCONNECTED__717, 
        SYNOPSYS_UNCONNECTED__718, SYNOPSYS_UNCONNECTED__719, 
        SYNOPSYS_UNCONNECTED__720, N30166, N30165, N30164, N30163, N30162, 
        N30161}) );
  hamming_N16000_CC4_DW01_add_148 add_1481_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28365, N28364, N28363, N28362, N28361}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28377, N28376, N28375, 
        N28374, N28373}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__721, 
        SYNOPSYS_UNCONNECTED__722, SYNOPSYS_UNCONNECTED__723, 
        SYNOPSYS_UNCONNECTED__724, SYNOPSYS_UNCONNECTED__725, 
        SYNOPSYS_UNCONNECTED__726, N30154, N30153, N30152, N30151, N30150, 
        N30149}) );
  hamming_N16000_CC4_DW01_add_149 add_1482_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28341, N28340, N28339, N28338, N28337}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28353, N28352, N28351, 
        N28350, N28349}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__727, 
        SYNOPSYS_UNCONNECTED__728, SYNOPSYS_UNCONNECTED__729, 
        SYNOPSYS_UNCONNECTED__730, SYNOPSYS_UNCONNECTED__731, 
        SYNOPSYS_UNCONNECTED__732, N30142, N30141, N30140, N30139, N30138, 
        N30137}) );
  hamming_N16000_CC4_DW01_add_150 add_1483_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28317, N28316, N28315, N28314, N28313}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28329, N28328, N28327, 
        N28326, N28325}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__733, 
        SYNOPSYS_UNCONNECTED__734, SYNOPSYS_UNCONNECTED__735, 
        SYNOPSYS_UNCONNECTED__736, SYNOPSYS_UNCONNECTED__737, 
        SYNOPSYS_UNCONNECTED__738, N30130, N30129, N30128, N30127, N30126, 
        N30125}) );
  hamming_N16000_CC4_DW01_add_151 add_1484_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28293, N28292, N28291, N28290, N28289}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28305, N28304, N28303, 
        N28302, N28301}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__739, 
        SYNOPSYS_UNCONNECTED__740, SYNOPSYS_UNCONNECTED__741, 
        SYNOPSYS_UNCONNECTED__742, SYNOPSYS_UNCONNECTED__743, 
        SYNOPSYS_UNCONNECTED__744, N30118, N30117, N30116, N30115, N30114, 
        N30113}) );
  hamming_N16000_CC4_DW01_add_152 add_1485_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28269, N28268, N28267, N28266, N28265}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28281, N28280, N28279, 
        N28278, N28277}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__745, 
        SYNOPSYS_UNCONNECTED__746, SYNOPSYS_UNCONNECTED__747, 
        SYNOPSYS_UNCONNECTED__748, SYNOPSYS_UNCONNECTED__749, 
        SYNOPSYS_UNCONNECTED__750, N30106, N30105, N30104, N30103, N30102, 
        N30101}) );
  hamming_N16000_CC4_DW01_add_153 add_1486_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28245, N28244, N28243, N28242, N28241}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28257, N28256, N28255, 
        N28254, N28253}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__751, 
        SYNOPSYS_UNCONNECTED__752, SYNOPSYS_UNCONNECTED__753, 
        SYNOPSYS_UNCONNECTED__754, SYNOPSYS_UNCONNECTED__755, 
        SYNOPSYS_UNCONNECTED__756, N30094, N30093, N30092, N30091, N30090, 
        N30089}) );
  hamming_N16000_CC4_DW01_add_154 add_1487_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28221, N28220, N28219, N28218, N28217}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28233, N28232, N28231, 
        N28230, N28229}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__757, 
        SYNOPSYS_UNCONNECTED__758, SYNOPSYS_UNCONNECTED__759, 
        SYNOPSYS_UNCONNECTED__760, SYNOPSYS_UNCONNECTED__761, 
        SYNOPSYS_UNCONNECTED__762, N30082, N30081, N30080, N30079, N30078, 
        N30077}) );
  hamming_N16000_CC4_DW01_add_155 add_1488_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28197, N28196, N28195, N28194, N28193}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28209, N28208, N28207, 
        N28206, N28205}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__763, 
        SYNOPSYS_UNCONNECTED__764, SYNOPSYS_UNCONNECTED__765, 
        SYNOPSYS_UNCONNECTED__766, SYNOPSYS_UNCONNECTED__767, 
        SYNOPSYS_UNCONNECTED__768, N30070, N30069, N30068, N30067, N30066, 
        N30065}) );
  hamming_N16000_CC4_DW01_add_156 add_1489_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28173, N28172, N28171, N28170, N28169}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28185, N28184, N28183, 
        N28182, N28181}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__769, 
        SYNOPSYS_UNCONNECTED__770, SYNOPSYS_UNCONNECTED__771, 
        SYNOPSYS_UNCONNECTED__772, SYNOPSYS_UNCONNECTED__773, 
        SYNOPSYS_UNCONNECTED__774, N30058, N30057, N30056, N30055, N30054, 
        N30053}) );
  hamming_N16000_CC4_DW01_add_157 add_1490_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28149, N28148, N28147, N28146, N28145}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28161, N28160, N28159, 
        N28158, N28157}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__775, 
        SYNOPSYS_UNCONNECTED__776, SYNOPSYS_UNCONNECTED__777, 
        SYNOPSYS_UNCONNECTED__778, SYNOPSYS_UNCONNECTED__779, 
        SYNOPSYS_UNCONNECTED__780, N30046, N30045, N30044, N30043, N30042, 
        N30041}) );
  hamming_N16000_CC4_DW01_add_158 add_1491_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28125, N28124, N28123, N28122, N28121}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28137, N28136, N28135, 
        N28134, N28133}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__781, 
        SYNOPSYS_UNCONNECTED__782, SYNOPSYS_UNCONNECTED__783, 
        SYNOPSYS_UNCONNECTED__784, SYNOPSYS_UNCONNECTED__785, 
        SYNOPSYS_UNCONNECTED__786, N30034, N30033, N30032, N30031, N30030, 
        N30029}) );
  hamming_N16000_CC4_DW01_add_159 add_1492_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28101, N28100, N28099, N28098, N28097}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28113, N28112, N28111, 
        N28110, N28109}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__787, 
        SYNOPSYS_UNCONNECTED__788, SYNOPSYS_UNCONNECTED__789, 
        SYNOPSYS_UNCONNECTED__790, SYNOPSYS_UNCONNECTED__791, 
        SYNOPSYS_UNCONNECTED__792, N30022, N30021, N30020, N30019, N30018, 
        N30017}) );
  hamming_N16000_CC4_DW01_add_160 add_1493_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28077, N28076, N28075, N28074, N28073}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28089, N28088, N28087, 
        N28086, N28085}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__793, 
        SYNOPSYS_UNCONNECTED__794, SYNOPSYS_UNCONNECTED__795, 
        SYNOPSYS_UNCONNECTED__796, SYNOPSYS_UNCONNECTED__797, 
        SYNOPSYS_UNCONNECTED__798, N30010, N30009, N30008, N30007, N30006, 
        N30005}) );
  hamming_N16000_CC4_DW01_add_161 add_1494_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28053, N28052, N28051, N28050, N28049}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28065, N28064, N28063, 
        N28062, N28061}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__799, 
        SYNOPSYS_UNCONNECTED__800, SYNOPSYS_UNCONNECTED__801, 
        SYNOPSYS_UNCONNECTED__802, SYNOPSYS_UNCONNECTED__803, 
        SYNOPSYS_UNCONNECTED__804, N29998, N29997, N29996, N29995, N29994, 
        N29993}) );
  hamming_N16000_CC4_DW01_add_162 add_1495_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28029, N28028, N28027, N28026, N28025}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28041, N28040, N28039, 
        N28038, N28037}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__805, 
        SYNOPSYS_UNCONNECTED__806, SYNOPSYS_UNCONNECTED__807, 
        SYNOPSYS_UNCONNECTED__808, SYNOPSYS_UNCONNECTED__809, 
        SYNOPSYS_UNCONNECTED__810, N29986, N29985, N29984, N29983, N29982, 
        N29981}) );
  hamming_N16000_CC4_DW01_add_163 add_1496_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28005, N28004, N28003, N28002, N28001}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N28017, N28016, N28015, 
        N28014, N28013}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__811, 
        SYNOPSYS_UNCONNECTED__812, SYNOPSYS_UNCONNECTED__813, 
        SYNOPSYS_UNCONNECTED__814, SYNOPSYS_UNCONNECTED__815, 
        SYNOPSYS_UNCONNECTED__816, N29974, N29973, N29972, N29971, N29970, 
        N29969}) );
  hamming_N16000_CC4_DW01_add_164 add_1497_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27981, N27980, N27979, N27978, N27977}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27993, N27992, N27991, 
        N27990, N27989}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__817, 
        SYNOPSYS_UNCONNECTED__818, SYNOPSYS_UNCONNECTED__819, 
        SYNOPSYS_UNCONNECTED__820, SYNOPSYS_UNCONNECTED__821, 
        SYNOPSYS_UNCONNECTED__822, N29962, N29961, N29960, N29959, N29958, 
        N29957}) );
  hamming_N16000_CC4_DW01_add_165 add_1498_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27957, N27956, N27955, N27954, N27953}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27969, N27968, N27967, 
        N27966, N27965}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__823, 
        SYNOPSYS_UNCONNECTED__824, SYNOPSYS_UNCONNECTED__825, 
        SYNOPSYS_UNCONNECTED__826, SYNOPSYS_UNCONNECTED__827, 
        SYNOPSYS_UNCONNECTED__828, N29950, N29949, N29948, N29947, N29946, 
        N29945}) );
  hamming_N16000_CC4_DW01_add_166 add_1499_root_add_71_I928 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27933, N27932, N27931, N27930, N27929}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N27945, N27944, N27943, 
        N27942, N27941}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__829, 
        SYNOPSYS_UNCONNECTED__830, SYNOPSYS_UNCONNECTED__831, 
        SYNOPSYS_UNCONNECTED__832, SYNOPSYS_UNCONNECTED__833, 
        SYNOPSYS_UNCONNECTED__834, N29938, N29937, N29936, N29935, N29934, 
        N29933}) );
  NAND U6683 ( .A(n2684), .B(n2685), .Z(N29925) );
  NAND U6684 ( .A(n2686), .B(n2687), .Z(n2685) );
  NANDN U6685 ( .A(n2688), .B(n2689), .Z(n2687) );
  NANDN U6686 ( .A(n2689), .B(n2688), .Z(n2684) );
  XOR U6687 ( .A(n2688), .B(n2690), .Z(N29924) );
  XNOR U6688 ( .A(n2686), .B(n2689), .Z(n2690) );
  NAND U6689 ( .A(n2691), .B(n2692), .Z(n2689) );
  NAND U6690 ( .A(n2693), .B(n2694), .Z(n2692) );
  NANDN U6691 ( .A(n2695), .B(n2696), .Z(n2694) );
  NANDN U6692 ( .A(n2696), .B(n2695), .Z(n2691) );
  AND U6693 ( .A(n2697), .B(n2698), .Z(n2686) );
  NAND U6694 ( .A(n2699), .B(n2700), .Z(n2698) );
  OR U6695 ( .A(n2701), .B(n2702), .Z(n2700) );
  NAND U6696 ( .A(n2702), .B(n2701), .Z(n2697) );
  IV U6697 ( .A(n2703), .Z(n2702) );
  AND U6698 ( .A(n2704), .B(n2705), .Z(n2688) );
  NAND U6699 ( .A(n2706), .B(n2707), .Z(n2705) );
  NANDN U6700 ( .A(n2708), .B(n2709), .Z(n2707) );
  NANDN U6701 ( .A(n2709), .B(n2708), .Z(n2704) );
  XOR U6702 ( .A(n2701), .B(n2710), .Z(N29923) );
  XOR U6703 ( .A(n2699), .B(n2703), .Z(n2710) );
  XNOR U6704 ( .A(n2696), .B(n2711), .Z(n2703) );
  XNOR U6705 ( .A(n2693), .B(n2695), .Z(n2711) );
  AND U6706 ( .A(n2712), .B(n2713), .Z(n2695) );
  NANDN U6707 ( .A(n2714), .B(n2715), .Z(n2713) );
  NANDN U6708 ( .A(n2716), .B(n2717), .Z(n2715) );
  IV U6709 ( .A(n2718), .Z(n2717) );
  NAND U6710 ( .A(n2718), .B(n2716), .Z(n2712) );
  AND U6711 ( .A(n2719), .B(n2720), .Z(n2693) );
  NAND U6712 ( .A(n2721), .B(n2722), .Z(n2720) );
  OR U6713 ( .A(n2723), .B(n2724), .Z(n2722) );
  NAND U6714 ( .A(n2724), .B(n2723), .Z(n2719) );
  IV U6715 ( .A(n2725), .Z(n2724) );
  NAND U6716 ( .A(n2726), .B(n2727), .Z(n2696) );
  NANDN U6717 ( .A(n2728), .B(n2729), .Z(n2727) );
  NAND U6718 ( .A(n2730), .B(n2731), .Z(n2729) );
  OR U6719 ( .A(n2731), .B(n2730), .Z(n2726) );
  IV U6720 ( .A(n2732), .Z(n2730) );
  AND U6721 ( .A(n2733), .B(n2734), .Z(n2699) );
  NAND U6722 ( .A(n2735), .B(n2736), .Z(n2734) );
  NANDN U6723 ( .A(n2737), .B(n2738), .Z(n2736) );
  NANDN U6724 ( .A(n2738), .B(n2737), .Z(n2733) );
  XOR U6725 ( .A(n2709), .B(n2739), .Z(n2701) );
  XNOR U6726 ( .A(n2706), .B(n2708), .Z(n2739) );
  AND U6727 ( .A(n2740), .B(n2741), .Z(n2708) );
  NANDN U6728 ( .A(n2742), .B(n2743), .Z(n2741) );
  NANDN U6729 ( .A(n2744), .B(n2745), .Z(n2743) );
  IV U6730 ( .A(n2746), .Z(n2745) );
  NAND U6731 ( .A(n2746), .B(n2744), .Z(n2740) );
  AND U6732 ( .A(n2747), .B(n2748), .Z(n2706) );
  NAND U6733 ( .A(n2749), .B(n2750), .Z(n2748) );
  OR U6734 ( .A(n2751), .B(n2752), .Z(n2750) );
  NAND U6735 ( .A(n2752), .B(n2751), .Z(n2747) );
  IV U6736 ( .A(n2753), .Z(n2752) );
  NAND U6737 ( .A(n2754), .B(n2755), .Z(n2709) );
  NANDN U6738 ( .A(n2756), .B(n2757), .Z(n2755) );
  NAND U6739 ( .A(n2758), .B(n2759), .Z(n2757) );
  OR U6740 ( .A(n2759), .B(n2758), .Z(n2754) );
  IV U6741 ( .A(n2760), .Z(n2758) );
  XOR U6742 ( .A(n2735), .B(n2761), .Z(N29922) );
  XNOR U6743 ( .A(n2738), .B(n2737), .Z(n2761) );
  XNOR U6744 ( .A(n2749), .B(n2762), .Z(n2737) );
  XOR U6745 ( .A(n2753), .B(n2751), .Z(n2762) );
  XOR U6746 ( .A(n2759), .B(n2763), .Z(n2751) );
  XOR U6747 ( .A(n2756), .B(n2760), .Z(n2763) );
  NAND U6748 ( .A(n2764), .B(n2765), .Z(n2760) );
  NAND U6749 ( .A(n2766), .B(n2767), .Z(n2765) );
  NAND U6750 ( .A(n2768), .B(n2769), .Z(n2764) );
  AND U6751 ( .A(n2770), .B(n2771), .Z(n2756) );
  NAND U6752 ( .A(n2772), .B(n2773), .Z(n2771) );
  NAND U6753 ( .A(n2774), .B(n2775), .Z(n2770) );
  NANDN U6754 ( .A(n2776), .B(n2777), .Z(n2759) );
  NANDN U6755 ( .A(n2778), .B(n2779), .Z(n2753) );
  XNOR U6756 ( .A(n2744), .B(n2780), .Z(n2749) );
  XOR U6757 ( .A(n2742), .B(n2746), .Z(n2780) );
  NAND U6758 ( .A(n2781), .B(n2782), .Z(n2746) );
  NAND U6759 ( .A(n2783), .B(n2784), .Z(n2782) );
  NAND U6760 ( .A(n2785), .B(n2786), .Z(n2781) );
  AND U6761 ( .A(n2787), .B(n2788), .Z(n2742) );
  NAND U6762 ( .A(n2789), .B(n2790), .Z(n2788) );
  NAND U6763 ( .A(n2791), .B(n2792), .Z(n2787) );
  AND U6764 ( .A(n2793), .B(n2794), .Z(n2744) );
  NAND U6765 ( .A(n2795), .B(n2796), .Z(n2738) );
  XNOR U6766 ( .A(n2721), .B(n2797), .Z(n2735) );
  XOR U6767 ( .A(n2725), .B(n2723), .Z(n2797) );
  XOR U6768 ( .A(n2731), .B(n2798), .Z(n2723) );
  XOR U6769 ( .A(n2728), .B(n2732), .Z(n2798) );
  NAND U6770 ( .A(n2799), .B(n2800), .Z(n2732) );
  NAND U6771 ( .A(n2801), .B(n2802), .Z(n2800) );
  NAND U6772 ( .A(n2803), .B(n2804), .Z(n2799) );
  AND U6773 ( .A(n2805), .B(n2806), .Z(n2728) );
  NAND U6774 ( .A(n2807), .B(n2808), .Z(n2806) );
  NAND U6775 ( .A(n2809), .B(n2810), .Z(n2805) );
  NANDN U6776 ( .A(n2811), .B(n2812), .Z(n2731) );
  NANDN U6777 ( .A(n2813), .B(n2814), .Z(n2725) );
  XNOR U6778 ( .A(n2716), .B(n2815), .Z(n2721) );
  XOR U6779 ( .A(n2714), .B(n2718), .Z(n2815) );
  NAND U6780 ( .A(n2816), .B(n2817), .Z(n2718) );
  NAND U6781 ( .A(n2818), .B(n2819), .Z(n2817) );
  NAND U6782 ( .A(n2820), .B(n2821), .Z(n2816) );
  AND U6783 ( .A(n2822), .B(n2823), .Z(n2714) );
  NAND U6784 ( .A(n2824), .B(n2825), .Z(n2823) );
  NAND U6785 ( .A(n2826), .B(n2827), .Z(n2822) );
  AND U6786 ( .A(n2828), .B(n2829), .Z(n2716) );
  XOR U6787 ( .A(n2796), .B(n2795), .Z(N29921) );
  XNOR U6788 ( .A(n2814), .B(n2813), .Z(n2795) );
  XNOR U6789 ( .A(n2828), .B(n2829), .Z(n2813) );
  XOR U6790 ( .A(n2825), .B(n2824), .Z(n2829) );
  XOR U6791 ( .A(y[3987]), .B(x[3987]), .Z(n2824) );
  XOR U6792 ( .A(n2827), .B(n2826), .Z(n2825) );
  XOR U6793 ( .A(y[3989]), .B(x[3989]), .Z(n2826) );
  XOR U6794 ( .A(y[3988]), .B(x[3988]), .Z(n2827) );
  XOR U6795 ( .A(n2819), .B(n2818), .Z(n2828) );
  XOR U6796 ( .A(n2821), .B(n2820), .Z(n2818) );
  XOR U6797 ( .A(y[3986]), .B(x[3986]), .Z(n2820) );
  XOR U6798 ( .A(y[3985]), .B(x[3985]), .Z(n2821) );
  XOR U6799 ( .A(y[3984]), .B(x[3984]), .Z(n2819) );
  XNOR U6800 ( .A(n2812), .B(n2811), .Z(n2814) );
  XNOR U6801 ( .A(n2808), .B(n2807), .Z(n2811) );
  XOR U6802 ( .A(n2810), .B(n2809), .Z(n2807) );
  XOR U6803 ( .A(y[3983]), .B(x[3983]), .Z(n2809) );
  XOR U6804 ( .A(y[3982]), .B(x[3982]), .Z(n2810) );
  XOR U6805 ( .A(y[3981]), .B(x[3981]), .Z(n2808) );
  XOR U6806 ( .A(n2802), .B(n2801), .Z(n2812) );
  XOR U6807 ( .A(n2804), .B(n2803), .Z(n2801) );
  XOR U6808 ( .A(y[3980]), .B(x[3980]), .Z(n2803) );
  XOR U6809 ( .A(y[3979]), .B(x[3979]), .Z(n2804) );
  XOR U6810 ( .A(y[3978]), .B(x[3978]), .Z(n2802) );
  XNOR U6811 ( .A(n2779), .B(n2778), .Z(n2796) );
  XNOR U6812 ( .A(n2793), .B(n2794), .Z(n2778) );
  XOR U6813 ( .A(n2790), .B(n2789), .Z(n2794) );
  XOR U6814 ( .A(y[3975]), .B(x[3975]), .Z(n2789) );
  XOR U6815 ( .A(n2792), .B(n2791), .Z(n2790) );
  XOR U6816 ( .A(y[3977]), .B(x[3977]), .Z(n2791) );
  XOR U6817 ( .A(y[3976]), .B(x[3976]), .Z(n2792) );
  XOR U6818 ( .A(n2784), .B(n2783), .Z(n2793) );
  XOR U6819 ( .A(n2786), .B(n2785), .Z(n2783) );
  XOR U6820 ( .A(y[3974]), .B(x[3974]), .Z(n2785) );
  XOR U6821 ( .A(y[3973]), .B(x[3973]), .Z(n2786) );
  XOR U6822 ( .A(y[3972]), .B(x[3972]), .Z(n2784) );
  XNOR U6823 ( .A(n2777), .B(n2776), .Z(n2779) );
  XNOR U6824 ( .A(n2773), .B(n2772), .Z(n2776) );
  XOR U6825 ( .A(n2775), .B(n2774), .Z(n2772) );
  XOR U6826 ( .A(y[3971]), .B(x[3971]), .Z(n2774) );
  XOR U6827 ( .A(y[3970]), .B(x[3970]), .Z(n2775) );
  XOR U6828 ( .A(y[3969]), .B(x[3969]), .Z(n2773) );
  XOR U6829 ( .A(n2767), .B(n2766), .Z(n2777) );
  XOR U6830 ( .A(n2769), .B(n2768), .Z(n2766) );
  XOR U6831 ( .A(y[3968]), .B(x[3968]), .Z(n2768) );
  XOR U6832 ( .A(y[3967]), .B(x[3967]), .Z(n2769) );
  XOR U6833 ( .A(y[3966]), .B(x[3966]), .Z(n2767) );
  NAND U6834 ( .A(n2830), .B(n2831), .Z(N29913) );
  NAND U6835 ( .A(n2832), .B(n2833), .Z(n2831) );
  NANDN U6836 ( .A(n2834), .B(n2835), .Z(n2833) );
  NANDN U6837 ( .A(n2835), .B(n2834), .Z(n2830) );
  XOR U6838 ( .A(n2834), .B(n2836), .Z(N29912) );
  XNOR U6839 ( .A(n2832), .B(n2835), .Z(n2836) );
  NAND U6840 ( .A(n2837), .B(n2838), .Z(n2835) );
  NAND U6841 ( .A(n2839), .B(n2840), .Z(n2838) );
  NANDN U6842 ( .A(n2841), .B(n2842), .Z(n2840) );
  NANDN U6843 ( .A(n2842), .B(n2841), .Z(n2837) );
  AND U6844 ( .A(n2843), .B(n2844), .Z(n2832) );
  NAND U6845 ( .A(n2845), .B(n2846), .Z(n2844) );
  OR U6846 ( .A(n2847), .B(n2848), .Z(n2846) );
  NAND U6847 ( .A(n2848), .B(n2847), .Z(n2843) );
  IV U6848 ( .A(n2849), .Z(n2848) );
  AND U6849 ( .A(n2850), .B(n2851), .Z(n2834) );
  NAND U6850 ( .A(n2852), .B(n2853), .Z(n2851) );
  NANDN U6851 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U6852 ( .A(n2855), .B(n2854), .Z(n2850) );
  XOR U6853 ( .A(n2847), .B(n2856), .Z(N29911) );
  XOR U6854 ( .A(n2845), .B(n2849), .Z(n2856) );
  XNOR U6855 ( .A(n2842), .B(n2857), .Z(n2849) );
  XNOR U6856 ( .A(n2839), .B(n2841), .Z(n2857) );
  AND U6857 ( .A(n2858), .B(n2859), .Z(n2841) );
  NANDN U6858 ( .A(n2860), .B(n2861), .Z(n2859) );
  NANDN U6859 ( .A(n2862), .B(n2863), .Z(n2861) );
  IV U6860 ( .A(n2864), .Z(n2863) );
  NAND U6861 ( .A(n2864), .B(n2862), .Z(n2858) );
  AND U6862 ( .A(n2865), .B(n2866), .Z(n2839) );
  NAND U6863 ( .A(n2867), .B(n2868), .Z(n2866) );
  OR U6864 ( .A(n2869), .B(n2870), .Z(n2868) );
  NAND U6865 ( .A(n2870), .B(n2869), .Z(n2865) );
  IV U6866 ( .A(n2871), .Z(n2870) );
  NAND U6867 ( .A(n2872), .B(n2873), .Z(n2842) );
  NANDN U6868 ( .A(n2874), .B(n2875), .Z(n2873) );
  NAND U6869 ( .A(n2876), .B(n2877), .Z(n2875) );
  OR U6870 ( .A(n2877), .B(n2876), .Z(n2872) );
  IV U6871 ( .A(n2878), .Z(n2876) );
  AND U6872 ( .A(n2879), .B(n2880), .Z(n2845) );
  NAND U6873 ( .A(n2881), .B(n2882), .Z(n2880) );
  NANDN U6874 ( .A(n2883), .B(n2884), .Z(n2882) );
  NANDN U6875 ( .A(n2884), .B(n2883), .Z(n2879) );
  XOR U6876 ( .A(n2855), .B(n2885), .Z(n2847) );
  XNOR U6877 ( .A(n2852), .B(n2854), .Z(n2885) );
  AND U6878 ( .A(n2886), .B(n2887), .Z(n2854) );
  NANDN U6879 ( .A(n2888), .B(n2889), .Z(n2887) );
  NANDN U6880 ( .A(n2890), .B(n2891), .Z(n2889) );
  IV U6881 ( .A(n2892), .Z(n2891) );
  NAND U6882 ( .A(n2892), .B(n2890), .Z(n2886) );
  AND U6883 ( .A(n2893), .B(n2894), .Z(n2852) );
  NAND U6884 ( .A(n2895), .B(n2896), .Z(n2894) );
  OR U6885 ( .A(n2897), .B(n2898), .Z(n2896) );
  NAND U6886 ( .A(n2898), .B(n2897), .Z(n2893) );
  IV U6887 ( .A(n2899), .Z(n2898) );
  NAND U6888 ( .A(n2900), .B(n2901), .Z(n2855) );
  NANDN U6889 ( .A(n2902), .B(n2903), .Z(n2901) );
  NAND U6890 ( .A(n2904), .B(n2905), .Z(n2903) );
  OR U6891 ( .A(n2905), .B(n2904), .Z(n2900) );
  IV U6892 ( .A(n2906), .Z(n2904) );
  XOR U6893 ( .A(n2881), .B(n2907), .Z(N29910) );
  XNOR U6894 ( .A(n2884), .B(n2883), .Z(n2907) );
  XNOR U6895 ( .A(n2895), .B(n2908), .Z(n2883) );
  XOR U6896 ( .A(n2899), .B(n2897), .Z(n2908) );
  XOR U6897 ( .A(n2905), .B(n2909), .Z(n2897) );
  XOR U6898 ( .A(n2902), .B(n2906), .Z(n2909) );
  NAND U6899 ( .A(n2910), .B(n2911), .Z(n2906) );
  NAND U6900 ( .A(n2912), .B(n2913), .Z(n2911) );
  NAND U6901 ( .A(n2914), .B(n2915), .Z(n2910) );
  AND U6902 ( .A(n2916), .B(n2917), .Z(n2902) );
  NAND U6903 ( .A(n2918), .B(n2919), .Z(n2917) );
  NAND U6904 ( .A(n2920), .B(n2921), .Z(n2916) );
  NANDN U6905 ( .A(n2922), .B(n2923), .Z(n2905) );
  NANDN U6906 ( .A(n2924), .B(n2925), .Z(n2899) );
  XNOR U6907 ( .A(n2890), .B(n2926), .Z(n2895) );
  XOR U6908 ( .A(n2888), .B(n2892), .Z(n2926) );
  NAND U6909 ( .A(n2927), .B(n2928), .Z(n2892) );
  NAND U6910 ( .A(n2929), .B(n2930), .Z(n2928) );
  NAND U6911 ( .A(n2931), .B(n2932), .Z(n2927) );
  AND U6912 ( .A(n2933), .B(n2934), .Z(n2888) );
  NAND U6913 ( .A(n2935), .B(n2936), .Z(n2934) );
  NAND U6914 ( .A(n2937), .B(n2938), .Z(n2933) );
  AND U6915 ( .A(n2939), .B(n2940), .Z(n2890) );
  NAND U6916 ( .A(n2941), .B(n2942), .Z(n2884) );
  XNOR U6917 ( .A(n2867), .B(n2943), .Z(n2881) );
  XOR U6918 ( .A(n2871), .B(n2869), .Z(n2943) );
  XOR U6919 ( .A(n2877), .B(n2944), .Z(n2869) );
  XOR U6920 ( .A(n2874), .B(n2878), .Z(n2944) );
  NAND U6921 ( .A(n2945), .B(n2946), .Z(n2878) );
  NAND U6922 ( .A(n2947), .B(n2948), .Z(n2946) );
  NAND U6923 ( .A(n2949), .B(n2950), .Z(n2945) );
  AND U6924 ( .A(n2951), .B(n2952), .Z(n2874) );
  NAND U6925 ( .A(n2953), .B(n2954), .Z(n2952) );
  NAND U6926 ( .A(n2955), .B(n2956), .Z(n2951) );
  NANDN U6927 ( .A(n2957), .B(n2958), .Z(n2877) );
  NANDN U6928 ( .A(n2959), .B(n2960), .Z(n2871) );
  XNOR U6929 ( .A(n2862), .B(n2961), .Z(n2867) );
  XOR U6930 ( .A(n2860), .B(n2864), .Z(n2961) );
  NAND U6931 ( .A(n2962), .B(n2963), .Z(n2864) );
  NAND U6932 ( .A(n2964), .B(n2965), .Z(n2963) );
  NAND U6933 ( .A(n2966), .B(n2967), .Z(n2962) );
  AND U6934 ( .A(n2968), .B(n2969), .Z(n2860) );
  NAND U6935 ( .A(n2970), .B(n2971), .Z(n2969) );
  NAND U6936 ( .A(n2972), .B(n2973), .Z(n2968) );
  AND U6937 ( .A(n2974), .B(n2975), .Z(n2862) );
  XOR U6938 ( .A(n2942), .B(n2941), .Z(N29909) );
  XNOR U6939 ( .A(n2960), .B(n2959), .Z(n2941) );
  XNOR U6940 ( .A(n2974), .B(n2975), .Z(n2959) );
  XOR U6941 ( .A(n2971), .B(n2970), .Z(n2975) );
  XOR U6942 ( .A(y[3963]), .B(x[3963]), .Z(n2970) );
  XOR U6943 ( .A(n2973), .B(n2972), .Z(n2971) );
  XOR U6944 ( .A(y[3965]), .B(x[3965]), .Z(n2972) );
  XOR U6945 ( .A(y[3964]), .B(x[3964]), .Z(n2973) );
  XOR U6946 ( .A(n2965), .B(n2964), .Z(n2974) );
  XOR U6947 ( .A(n2967), .B(n2966), .Z(n2964) );
  XOR U6948 ( .A(y[3962]), .B(x[3962]), .Z(n2966) );
  XOR U6949 ( .A(y[3961]), .B(x[3961]), .Z(n2967) );
  XOR U6950 ( .A(y[3960]), .B(x[3960]), .Z(n2965) );
  XNOR U6951 ( .A(n2958), .B(n2957), .Z(n2960) );
  XNOR U6952 ( .A(n2954), .B(n2953), .Z(n2957) );
  XOR U6953 ( .A(n2956), .B(n2955), .Z(n2953) );
  XOR U6954 ( .A(y[3959]), .B(x[3959]), .Z(n2955) );
  XOR U6955 ( .A(y[3958]), .B(x[3958]), .Z(n2956) );
  XOR U6956 ( .A(y[3957]), .B(x[3957]), .Z(n2954) );
  XOR U6957 ( .A(n2948), .B(n2947), .Z(n2958) );
  XOR U6958 ( .A(n2950), .B(n2949), .Z(n2947) );
  XOR U6959 ( .A(y[3956]), .B(x[3956]), .Z(n2949) );
  XOR U6960 ( .A(y[3955]), .B(x[3955]), .Z(n2950) );
  XOR U6961 ( .A(y[3954]), .B(x[3954]), .Z(n2948) );
  XNOR U6962 ( .A(n2925), .B(n2924), .Z(n2942) );
  XNOR U6963 ( .A(n2939), .B(n2940), .Z(n2924) );
  XOR U6964 ( .A(n2936), .B(n2935), .Z(n2940) );
  XOR U6965 ( .A(y[3951]), .B(x[3951]), .Z(n2935) );
  XOR U6966 ( .A(n2938), .B(n2937), .Z(n2936) );
  XOR U6967 ( .A(y[3953]), .B(x[3953]), .Z(n2937) );
  XOR U6968 ( .A(y[3952]), .B(x[3952]), .Z(n2938) );
  XOR U6969 ( .A(n2930), .B(n2929), .Z(n2939) );
  XOR U6970 ( .A(n2932), .B(n2931), .Z(n2929) );
  XOR U6971 ( .A(y[3950]), .B(x[3950]), .Z(n2931) );
  XOR U6972 ( .A(y[3949]), .B(x[3949]), .Z(n2932) );
  XOR U6973 ( .A(y[3948]), .B(x[3948]), .Z(n2930) );
  XNOR U6974 ( .A(n2923), .B(n2922), .Z(n2925) );
  XNOR U6975 ( .A(n2919), .B(n2918), .Z(n2922) );
  XOR U6976 ( .A(n2921), .B(n2920), .Z(n2918) );
  XOR U6977 ( .A(y[3947]), .B(x[3947]), .Z(n2920) );
  XOR U6978 ( .A(y[3946]), .B(x[3946]), .Z(n2921) );
  XOR U6979 ( .A(y[3945]), .B(x[3945]), .Z(n2919) );
  XOR U6980 ( .A(n2913), .B(n2912), .Z(n2923) );
  XOR U6981 ( .A(n2915), .B(n2914), .Z(n2912) );
  XOR U6982 ( .A(y[3944]), .B(x[3944]), .Z(n2914) );
  XOR U6983 ( .A(y[3943]), .B(x[3943]), .Z(n2915) );
  XOR U6984 ( .A(y[3942]), .B(x[3942]), .Z(n2913) );
  NAND U6985 ( .A(n2976), .B(n2977), .Z(N29901) );
  NAND U6986 ( .A(n2978), .B(n2979), .Z(n2977) );
  NANDN U6987 ( .A(n2980), .B(n2981), .Z(n2979) );
  NANDN U6988 ( .A(n2981), .B(n2980), .Z(n2976) );
  XOR U6989 ( .A(n2980), .B(n2982), .Z(N29900) );
  XNOR U6990 ( .A(n2978), .B(n2981), .Z(n2982) );
  NAND U6991 ( .A(n2983), .B(n2984), .Z(n2981) );
  NAND U6992 ( .A(n2985), .B(n2986), .Z(n2984) );
  NANDN U6993 ( .A(n2987), .B(n2988), .Z(n2986) );
  NANDN U6994 ( .A(n2988), .B(n2987), .Z(n2983) );
  AND U6995 ( .A(n2989), .B(n2990), .Z(n2978) );
  NAND U6996 ( .A(n2991), .B(n2992), .Z(n2990) );
  OR U6997 ( .A(n2993), .B(n2994), .Z(n2992) );
  NAND U6998 ( .A(n2994), .B(n2993), .Z(n2989) );
  IV U6999 ( .A(n2995), .Z(n2994) );
  AND U7000 ( .A(n2996), .B(n2997), .Z(n2980) );
  NAND U7001 ( .A(n2998), .B(n2999), .Z(n2997) );
  NANDN U7002 ( .A(n3000), .B(n3001), .Z(n2999) );
  NANDN U7003 ( .A(n3001), .B(n3000), .Z(n2996) );
  XOR U7004 ( .A(n2993), .B(n3002), .Z(N29899) );
  XOR U7005 ( .A(n2991), .B(n2995), .Z(n3002) );
  XNOR U7006 ( .A(n2988), .B(n3003), .Z(n2995) );
  XNOR U7007 ( .A(n2985), .B(n2987), .Z(n3003) );
  AND U7008 ( .A(n3004), .B(n3005), .Z(n2987) );
  NANDN U7009 ( .A(n3006), .B(n3007), .Z(n3005) );
  NANDN U7010 ( .A(n3008), .B(n3009), .Z(n3007) );
  IV U7011 ( .A(n3010), .Z(n3009) );
  NAND U7012 ( .A(n3010), .B(n3008), .Z(n3004) );
  AND U7013 ( .A(n3011), .B(n3012), .Z(n2985) );
  NAND U7014 ( .A(n3013), .B(n3014), .Z(n3012) );
  OR U7015 ( .A(n3015), .B(n3016), .Z(n3014) );
  NAND U7016 ( .A(n3016), .B(n3015), .Z(n3011) );
  IV U7017 ( .A(n3017), .Z(n3016) );
  NAND U7018 ( .A(n3018), .B(n3019), .Z(n2988) );
  NANDN U7019 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U7020 ( .A(n3022), .B(n3023), .Z(n3021) );
  OR U7021 ( .A(n3023), .B(n3022), .Z(n3018) );
  IV U7022 ( .A(n3024), .Z(n3022) );
  AND U7023 ( .A(n3025), .B(n3026), .Z(n2991) );
  NAND U7024 ( .A(n3027), .B(n3028), .Z(n3026) );
  NANDN U7025 ( .A(n3029), .B(n3030), .Z(n3028) );
  NANDN U7026 ( .A(n3030), .B(n3029), .Z(n3025) );
  XOR U7027 ( .A(n3001), .B(n3031), .Z(n2993) );
  XNOR U7028 ( .A(n2998), .B(n3000), .Z(n3031) );
  AND U7029 ( .A(n3032), .B(n3033), .Z(n3000) );
  NANDN U7030 ( .A(n3034), .B(n3035), .Z(n3033) );
  NANDN U7031 ( .A(n3036), .B(n3037), .Z(n3035) );
  IV U7032 ( .A(n3038), .Z(n3037) );
  NAND U7033 ( .A(n3038), .B(n3036), .Z(n3032) );
  AND U7034 ( .A(n3039), .B(n3040), .Z(n2998) );
  NAND U7035 ( .A(n3041), .B(n3042), .Z(n3040) );
  OR U7036 ( .A(n3043), .B(n3044), .Z(n3042) );
  NAND U7037 ( .A(n3044), .B(n3043), .Z(n3039) );
  IV U7038 ( .A(n3045), .Z(n3044) );
  NAND U7039 ( .A(n3046), .B(n3047), .Z(n3001) );
  NANDN U7040 ( .A(n3048), .B(n3049), .Z(n3047) );
  NAND U7041 ( .A(n3050), .B(n3051), .Z(n3049) );
  OR U7042 ( .A(n3051), .B(n3050), .Z(n3046) );
  IV U7043 ( .A(n3052), .Z(n3050) );
  XOR U7044 ( .A(n3027), .B(n3053), .Z(N29898) );
  XNOR U7045 ( .A(n3030), .B(n3029), .Z(n3053) );
  XNOR U7046 ( .A(n3041), .B(n3054), .Z(n3029) );
  XOR U7047 ( .A(n3045), .B(n3043), .Z(n3054) );
  XOR U7048 ( .A(n3051), .B(n3055), .Z(n3043) );
  XOR U7049 ( .A(n3048), .B(n3052), .Z(n3055) );
  NAND U7050 ( .A(n3056), .B(n3057), .Z(n3052) );
  NAND U7051 ( .A(n3058), .B(n3059), .Z(n3057) );
  NAND U7052 ( .A(n3060), .B(n3061), .Z(n3056) );
  AND U7053 ( .A(n3062), .B(n3063), .Z(n3048) );
  NAND U7054 ( .A(n3064), .B(n3065), .Z(n3063) );
  NAND U7055 ( .A(n3066), .B(n3067), .Z(n3062) );
  NANDN U7056 ( .A(n3068), .B(n3069), .Z(n3051) );
  NANDN U7057 ( .A(n3070), .B(n3071), .Z(n3045) );
  XNOR U7058 ( .A(n3036), .B(n3072), .Z(n3041) );
  XOR U7059 ( .A(n3034), .B(n3038), .Z(n3072) );
  NAND U7060 ( .A(n3073), .B(n3074), .Z(n3038) );
  NAND U7061 ( .A(n3075), .B(n3076), .Z(n3074) );
  NAND U7062 ( .A(n3077), .B(n3078), .Z(n3073) );
  AND U7063 ( .A(n3079), .B(n3080), .Z(n3034) );
  NAND U7064 ( .A(n3081), .B(n3082), .Z(n3080) );
  NAND U7065 ( .A(n3083), .B(n3084), .Z(n3079) );
  AND U7066 ( .A(n3085), .B(n3086), .Z(n3036) );
  NAND U7067 ( .A(n3087), .B(n3088), .Z(n3030) );
  XNOR U7068 ( .A(n3013), .B(n3089), .Z(n3027) );
  XOR U7069 ( .A(n3017), .B(n3015), .Z(n3089) );
  XOR U7070 ( .A(n3023), .B(n3090), .Z(n3015) );
  XOR U7071 ( .A(n3020), .B(n3024), .Z(n3090) );
  NAND U7072 ( .A(n3091), .B(n3092), .Z(n3024) );
  NAND U7073 ( .A(n3093), .B(n3094), .Z(n3092) );
  NAND U7074 ( .A(n3095), .B(n3096), .Z(n3091) );
  AND U7075 ( .A(n3097), .B(n3098), .Z(n3020) );
  NAND U7076 ( .A(n3099), .B(n3100), .Z(n3098) );
  NAND U7077 ( .A(n3101), .B(n3102), .Z(n3097) );
  NANDN U7078 ( .A(n3103), .B(n3104), .Z(n3023) );
  NANDN U7079 ( .A(n3105), .B(n3106), .Z(n3017) );
  XNOR U7080 ( .A(n3008), .B(n3107), .Z(n3013) );
  XOR U7081 ( .A(n3006), .B(n3010), .Z(n3107) );
  NAND U7082 ( .A(n3108), .B(n3109), .Z(n3010) );
  NAND U7083 ( .A(n3110), .B(n3111), .Z(n3109) );
  NAND U7084 ( .A(n3112), .B(n3113), .Z(n3108) );
  AND U7085 ( .A(n3114), .B(n3115), .Z(n3006) );
  NAND U7086 ( .A(n3116), .B(n3117), .Z(n3115) );
  NAND U7087 ( .A(n3118), .B(n3119), .Z(n3114) );
  AND U7088 ( .A(n3120), .B(n3121), .Z(n3008) );
  XOR U7089 ( .A(n3088), .B(n3087), .Z(N29897) );
  XNOR U7090 ( .A(n3106), .B(n3105), .Z(n3087) );
  XNOR U7091 ( .A(n3120), .B(n3121), .Z(n3105) );
  XOR U7092 ( .A(n3117), .B(n3116), .Z(n3121) );
  XOR U7093 ( .A(y[3939]), .B(x[3939]), .Z(n3116) );
  XOR U7094 ( .A(n3119), .B(n3118), .Z(n3117) );
  XOR U7095 ( .A(y[3941]), .B(x[3941]), .Z(n3118) );
  XOR U7096 ( .A(y[3940]), .B(x[3940]), .Z(n3119) );
  XOR U7097 ( .A(n3111), .B(n3110), .Z(n3120) );
  XOR U7098 ( .A(n3113), .B(n3112), .Z(n3110) );
  XOR U7099 ( .A(y[3938]), .B(x[3938]), .Z(n3112) );
  XOR U7100 ( .A(y[3937]), .B(x[3937]), .Z(n3113) );
  XOR U7101 ( .A(y[3936]), .B(x[3936]), .Z(n3111) );
  XNOR U7102 ( .A(n3104), .B(n3103), .Z(n3106) );
  XNOR U7103 ( .A(n3100), .B(n3099), .Z(n3103) );
  XOR U7104 ( .A(n3102), .B(n3101), .Z(n3099) );
  XOR U7105 ( .A(y[3935]), .B(x[3935]), .Z(n3101) );
  XOR U7106 ( .A(y[3934]), .B(x[3934]), .Z(n3102) );
  XOR U7107 ( .A(y[3933]), .B(x[3933]), .Z(n3100) );
  XOR U7108 ( .A(n3094), .B(n3093), .Z(n3104) );
  XOR U7109 ( .A(n3096), .B(n3095), .Z(n3093) );
  XOR U7110 ( .A(y[3932]), .B(x[3932]), .Z(n3095) );
  XOR U7111 ( .A(y[3931]), .B(x[3931]), .Z(n3096) );
  XOR U7112 ( .A(y[3930]), .B(x[3930]), .Z(n3094) );
  XNOR U7113 ( .A(n3071), .B(n3070), .Z(n3088) );
  XNOR U7114 ( .A(n3085), .B(n3086), .Z(n3070) );
  XOR U7115 ( .A(n3082), .B(n3081), .Z(n3086) );
  XOR U7116 ( .A(y[3927]), .B(x[3927]), .Z(n3081) );
  XOR U7117 ( .A(n3084), .B(n3083), .Z(n3082) );
  XOR U7118 ( .A(y[3929]), .B(x[3929]), .Z(n3083) );
  XOR U7119 ( .A(y[3928]), .B(x[3928]), .Z(n3084) );
  XOR U7120 ( .A(n3076), .B(n3075), .Z(n3085) );
  XOR U7121 ( .A(n3078), .B(n3077), .Z(n3075) );
  XOR U7122 ( .A(y[3926]), .B(x[3926]), .Z(n3077) );
  XOR U7123 ( .A(y[3925]), .B(x[3925]), .Z(n3078) );
  XOR U7124 ( .A(y[3924]), .B(x[3924]), .Z(n3076) );
  XNOR U7125 ( .A(n3069), .B(n3068), .Z(n3071) );
  XNOR U7126 ( .A(n3065), .B(n3064), .Z(n3068) );
  XOR U7127 ( .A(n3067), .B(n3066), .Z(n3064) );
  XOR U7128 ( .A(y[3923]), .B(x[3923]), .Z(n3066) );
  XOR U7129 ( .A(y[3922]), .B(x[3922]), .Z(n3067) );
  XOR U7130 ( .A(y[3921]), .B(x[3921]), .Z(n3065) );
  XOR U7131 ( .A(n3059), .B(n3058), .Z(n3069) );
  XOR U7132 ( .A(n3061), .B(n3060), .Z(n3058) );
  XOR U7133 ( .A(y[3920]), .B(x[3920]), .Z(n3060) );
  XOR U7134 ( .A(y[3919]), .B(x[3919]), .Z(n3061) );
  XOR U7135 ( .A(y[3918]), .B(x[3918]), .Z(n3059) );
  NAND U7136 ( .A(n3122), .B(n3123), .Z(N29889) );
  NAND U7137 ( .A(n3124), .B(n3125), .Z(n3123) );
  NANDN U7138 ( .A(n3126), .B(n3127), .Z(n3125) );
  NANDN U7139 ( .A(n3127), .B(n3126), .Z(n3122) );
  XOR U7140 ( .A(n3126), .B(n3128), .Z(N29888) );
  XNOR U7141 ( .A(n3124), .B(n3127), .Z(n3128) );
  NAND U7142 ( .A(n3129), .B(n3130), .Z(n3127) );
  NAND U7143 ( .A(n3131), .B(n3132), .Z(n3130) );
  NANDN U7144 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U7145 ( .A(n3134), .B(n3133), .Z(n3129) );
  AND U7146 ( .A(n3135), .B(n3136), .Z(n3124) );
  NAND U7147 ( .A(n3137), .B(n3138), .Z(n3136) );
  OR U7148 ( .A(n3139), .B(n3140), .Z(n3138) );
  NAND U7149 ( .A(n3140), .B(n3139), .Z(n3135) );
  IV U7150 ( .A(n3141), .Z(n3140) );
  AND U7151 ( .A(n3142), .B(n3143), .Z(n3126) );
  NAND U7152 ( .A(n3144), .B(n3145), .Z(n3143) );
  NANDN U7153 ( .A(n3146), .B(n3147), .Z(n3145) );
  NANDN U7154 ( .A(n3147), .B(n3146), .Z(n3142) );
  XOR U7155 ( .A(n3139), .B(n3148), .Z(N29887) );
  XOR U7156 ( .A(n3137), .B(n3141), .Z(n3148) );
  XNOR U7157 ( .A(n3134), .B(n3149), .Z(n3141) );
  XNOR U7158 ( .A(n3131), .B(n3133), .Z(n3149) );
  AND U7159 ( .A(n3150), .B(n3151), .Z(n3133) );
  NANDN U7160 ( .A(n3152), .B(n3153), .Z(n3151) );
  NANDN U7161 ( .A(n3154), .B(n3155), .Z(n3153) );
  IV U7162 ( .A(n3156), .Z(n3155) );
  NAND U7163 ( .A(n3156), .B(n3154), .Z(n3150) );
  AND U7164 ( .A(n3157), .B(n3158), .Z(n3131) );
  NAND U7165 ( .A(n3159), .B(n3160), .Z(n3158) );
  OR U7166 ( .A(n3161), .B(n3162), .Z(n3160) );
  NAND U7167 ( .A(n3162), .B(n3161), .Z(n3157) );
  IV U7168 ( .A(n3163), .Z(n3162) );
  NAND U7169 ( .A(n3164), .B(n3165), .Z(n3134) );
  NANDN U7170 ( .A(n3166), .B(n3167), .Z(n3165) );
  NAND U7171 ( .A(n3168), .B(n3169), .Z(n3167) );
  OR U7172 ( .A(n3169), .B(n3168), .Z(n3164) );
  IV U7173 ( .A(n3170), .Z(n3168) );
  AND U7174 ( .A(n3171), .B(n3172), .Z(n3137) );
  NAND U7175 ( .A(n3173), .B(n3174), .Z(n3172) );
  NANDN U7176 ( .A(n3175), .B(n3176), .Z(n3174) );
  NANDN U7177 ( .A(n3176), .B(n3175), .Z(n3171) );
  XOR U7178 ( .A(n3147), .B(n3177), .Z(n3139) );
  XNOR U7179 ( .A(n3144), .B(n3146), .Z(n3177) );
  AND U7180 ( .A(n3178), .B(n3179), .Z(n3146) );
  NANDN U7181 ( .A(n3180), .B(n3181), .Z(n3179) );
  NANDN U7182 ( .A(n3182), .B(n3183), .Z(n3181) );
  IV U7183 ( .A(n3184), .Z(n3183) );
  NAND U7184 ( .A(n3184), .B(n3182), .Z(n3178) );
  AND U7185 ( .A(n3185), .B(n3186), .Z(n3144) );
  NAND U7186 ( .A(n3187), .B(n3188), .Z(n3186) );
  OR U7187 ( .A(n3189), .B(n3190), .Z(n3188) );
  NAND U7188 ( .A(n3190), .B(n3189), .Z(n3185) );
  IV U7189 ( .A(n3191), .Z(n3190) );
  NAND U7190 ( .A(n3192), .B(n3193), .Z(n3147) );
  NANDN U7191 ( .A(n3194), .B(n3195), .Z(n3193) );
  NAND U7192 ( .A(n3196), .B(n3197), .Z(n3195) );
  OR U7193 ( .A(n3197), .B(n3196), .Z(n3192) );
  IV U7194 ( .A(n3198), .Z(n3196) );
  XOR U7195 ( .A(n3173), .B(n3199), .Z(N29886) );
  XNOR U7196 ( .A(n3176), .B(n3175), .Z(n3199) );
  XNOR U7197 ( .A(n3187), .B(n3200), .Z(n3175) );
  XOR U7198 ( .A(n3191), .B(n3189), .Z(n3200) );
  XOR U7199 ( .A(n3197), .B(n3201), .Z(n3189) );
  XOR U7200 ( .A(n3194), .B(n3198), .Z(n3201) );
  NAND U7201 ( .A(n3202), .B(n3203), .Z(n3198) );
  NAND U7202 ( .A(n3204), .B(n3205), .Z(n3203) );
  NAND U7203 ( .A(n3206), .B(n3207), .Z(n3202) );
  AND U7204 ( .A(n3208), .B(n3209), .Z(n3194) );
  NAND U7205 ( .A(n3210), .B(n3211), .Z(n3209) );
  NAND U7206 ( .A(n3212), .B(n3213), .Z(n3208) );
  NANDN U7207 ( .A(n3214), .B(n3215), .Z(n3197) );
  NANDN U7208 ( .A(n3216), .B(n3217), .Z(n3191) );
  XNOR U7209 ( .A(n3182), .B(n3218), .Z(n3187) );
  XOR U7210 ( .A(n3180), .B(n3184), .Z(n3218) );
  NAND U7211 ( .A(n3219), .B(n3220), .Z(n3184) );
  NAND U7212 ( .A(n3221), .B(n3222), .Z(n3220) );
  NAND U7213 ( .A(n3223), .B(n3224), .Z(n3219) );
  AND U7214 ( .A(n3225), .B(n3226), .Z(n3180) );
  NAND U7215 ( .A(n3227), .B(n3228), .Z(n3226) );
  NAND U7216 ( .A(n3229), .B(n3230), .Z(n3225) );
  AND U7217 ( .A(n3231), .B(n3232), .Z(n3182) );
  NAND U7218 ( .A(n3233), .B(n3234), .Z(n3176) );
  XNOR U7219 ( .A(n3159), .B(n3235), .Z(n3173) );
  XOR U7220 ( .A(n3163), .B(n3161), .Z(n3235) );
  XOR U7221 ( .A(n3169), .B(n3236), .Z(n3161) );
  XOR U7222 ( .A(n3166), .B(n3170), .Z(n3236) );
  NAND U7223 ( .A(n3237), .B(n3238), .Z(n3170) );
  NAND U7224 ( .A(n3239), .B(n3240), .Z(n3238) );
  NAND U7225 ( .A(n3241), .B(n3242), .Z(n3237) );
  AND U7226 ( .A(n3243), .B(n3244), .Z(n3166) );
  NAND U7227 ( .A(n3245), .B(n3246), .Z(n3244) );
  NAND U7228 ( .A(n3247), .B(n3248), .Z(n3243) );
  NANDN U7229 ( .A(n3249), .B(n3250), .Z(n3169) );
  NANDN U7230 ( .A(n3251), .B(n3252), .Z(n3163) );
  XNOR U7231 ( .A(n3154), .B(n3253), .Z(n3159) );
  XOR U7232 ( .A(n3152), .B(n3156), .Z(n3253) );
  NAND U7233 ( .A(n3254), .B(n3255), .Z(n3156) );
  NAND U7234 ( .A(n3256), .B(n3257), .Z(n3255) );
  NAND U7235 ( .A(n3258), .B(n3259), .Z(n3254) );
  AND U7236 ( .A(n3260), .B(n3261), .Z(n3152) );
  NAND U7237 ( .A(n3262), .B(n3263), .Z(n3261) );
  NAND U7238 ( .A(n3264), .B(n3265), .Z(n3260) );
  AND U7239 ( .A(n3266), .B(n3267), .Z(n3154) );
  XOR U7240 ( .A(n3234), .B(n3233), .Z(N29885) );
  XNOR U7241 ( .A(n3252), .B(n3251), .Z(n3233) );
  XNOR U7242 ( .A(n3266), .B(n3267), .Z(n3251) );
  XOR U7243 ( .A(n3263), .B(n3262), .Z(n3267) );
  XOR U7244 ( .A(y[3915]), .B(x[3915]), .Z(n3262) );
  XOR U7245 ( .A(n3265), .B(n3264), .Z(n3263) );
  XOR U7246 ( .A(y[3917]), .B(x[3917]), .Z(n3264) );
  XOR U7247 ( .A(y[3916]), .B(x[3916]), .Z(n3265) );
  XOR U7248 ( .A(n3257), .B(n3256), .Z(n3266) );
  XOR U7249 ( .A(n3259), .B(n3258), .Z(n3256) );
  XOR U7250 ( .A(y[3914]), .B(x[3914]), .Z(n3258) );
  XOR U7251 ( .A(y[3913]), .B(x[3913]), .Z(n3259) );
  XOR U7252 ( .A(y[3912]), .B(x[3912]), .Z(n3257) );
  XNOR U7253 ( .A(n3250), .B(n3249), .Z(n3252) );
  XNOR U7254 ( .A(n3246), .B(n3245), .Z(n3249) );
  XOR U7255 ( .A(n3248), .B(n3247), .Z(n3245) );
  XOR U7256 ( .A(y[3911]), .B(x[3911]), .Z(n3247) );
  XOR U7257 ( .A(y[3910]), .B(x[3910]), .Z(n3248) );
  XOR U7258 ( .A(y[3909]), .B(x[3909]), .Z(n3246) );
  XOR U7259 ( .A(n3240), .B(n3239), .Z(n3250) );
  XOR U7260 ( .A(n3242), .B(n3241), .Z(n3239) );
  XOR U7261 ( .A(y[3908]), .B(x[3908]), .Z(n3241) );
  XOR U7262 ( .A(y[3907]), .B(x[3907]), .Z(n3242) );
  XOR U7263 ( .A(y[3906]), .B(x[3906]), .Z(n3240) );
  XNOR U7264 ( .A(n3217), .B(n3216), .Z(n3234) );
  XNOR U7265 ( .A(n3231), .B(n3232), .Z(n3216) );
  XOR U7266 ( .A(n3228), .B(n3227), .Z(n3232) );
  XOR U7267 ( .A(y[3903]), .B(x[3903]), .Z(n3227) );
  XOR U7268 ( .A(n3230), .B(n3229), .Z(n3228) );
  XOR U7269 ( .A(y[3905]), .B(x[3905]), .Z(n3229) );
  XOR U7270 ( .A(y[3904]), .B(x[3904]), .Z(n3230) );
  XOR U7271 ( .A(n3222), .B(n3221), .Z(n3231) );
  XOR U7272 ( .A(n3224), .B(n3223), .Z(n3221) );
  XOR U7273 ( .A(y[3902]), .B(x[3902]), .Z(n3223) );
  XOR U7274 ( .A(y[3901]), .B(x[3901]), .Z(n3224) );
  XOR U7275 ( .A(y[3900]), .B(x[3900]), .Z(n3222) );
  XNOR U7276 ( .A(n3215), .B(n3214), .Z(n3217) );
  XNOR U7277 ( .A(n3211), .B(n3210), .Z(n3214) );
  XOR U7278 ( .A(n3213), .B(n3212), .Z(n3210) );
  XOR U7279 ( .A(y[3899]), .B(x[3899]), .Z(n3212) );
  XOR U7280 ( .A(y[3898]), .B(x[3898]), .Z(n3213) );
  XOR U7281 ( .A(y[3897]), .B(x[3897]), .Z(n3211) );
  XOR U7282 ( .A(n3205), .B(n3204), .Z(n3215) );
  XOR U7283 ( .A(n3207), .B(n3206), .Z(n3204) );
  XOR U7284 ( .A(y[3896]), .B(x[3896]), .Z(n3206) );
  XOR U7285 ( .A(y[3895]), .B(x[3895]), .Z(n3207) );
  XOR U7286 ( .A(y[3894]), .B(x[3894]), .Z(n3205) );
  NAND U7287 ( .A(n3268), .B(n3269), .Z(N29877) );
  NAND U7288 ( .A(n3270), .B(n3271), .Z(n3269) );
  NANDN U7289 ( .A(n3272), .B(n3273), .Z(n3271) );
  NANDN U7290 ( .A(n3273), .B(n3272), .Z(n3268) );
  XOR U7291 ( .A(n3272), .B(n3274), .Z(N29876) );
  XNOR U7292 ( .A(n3270), .B(n3273), .Z(n3274) );
  NAND U7293 ( .A(n3275), .B(n3276), .Z(n3273) );
  NAND U7294 ( .A(n3277), .B(n3278), .Z(n3276) );
  NANDN U7295 ( .A(n3279), .B(n3280), .Z(n3278) );
  NANDN U7296 ( .A(n3280), .B(n3279), .Z(n3275) );
  AND U7297 ( .A(n3281), .B(n3282), .Z(n3270) );
  NAND U7298 ( .A(n3283), .B(n3284), .Z(n3282) );
  OR U7299 ( .A(n3285), .B(n3286), .Z(n3284) );
  NAND U7300 ( .A(n3286), .B(n3285), .Z(n3281) );
  IV U7301 ( .A(n3287), .Z(n3286) );
  AND U7302 ( .A(n3288), .B(n3289), .Z(n3272) );
  NAND U7303 ( .A(n3290), .B(n3291), .Z(n3289) );
  NANDN U7304 ( .A(n3292), .B(n3293), .Z(n3291) );
  NANDN U7305 ( .A(n3293), .B(n3292), .Z(n3288) );
  XOR U7306 ( .A(n3285), .B(n3294), .Z(N29875) );
  XOR U7307 ( .A(n3283), .B(n3287), .Z(n3294) );
  XNOR U7308 ( .A(n3280), .B(n3295), .Z(n3287) );
  XNOR U7309 ( .A(n3277), .B(n3279), .Z(n3295) );
  AND U7310 ( .A(n3296), .B(n3297), .Z(n3279) );
  NANDN U7311 ( .A(n3298), .B(n3299), .Z(n3297) );
  NANDN U7312 ( .A(n3300), .B(n3301), .Z(n3299) );
  IV U7313 ( .A(n3302), .Z(n3301) );
  NAND U7314 ( .A(n3302), .B(n3300), .Z(n3296) );
  AND U7315 ( .A(n3303), .B(n3304), .Z(n3277) );
  NAND U7316 ( .A(n3305), .B(n3306), .Z(n3304) );
  OR U7317 ( .A(n3307), .B(n3308), .Z(n3306) );
  NAND U7318 ( .A(n3308), .B(n3307), .Z(n3303) );
  IV U7319 ( .A(n3309), .Z(n3308) );
  NAND U7320 ( .A(n3310), .B(n3311), .Z(n3280) );
  NANDN U7321 ( .A(n3312), .B(n3313), .Z(n3311) );
  NAND U7322 ( .A(n3314), .B(n3315), .Z(n3313) );
  OR U7323 ( .A(n3315), .B(n3314), .Z(n3310) );
  IV U7324 ( .A(n3316), .Z(n3314) );
  AND U7325 ( .A(n3317), .B(n3318), .Z(n3283) );
  NAND U7326 ( .A(n3319), .B(n3320), .Z(n3318) );
  NANDN U7327 ( .A(n3321), .B(n3322), .Z(n3320) );
  NANDN U7328 ( .A(n3322), .B(n3321), .Z(n3317) );
  XOR U7329 ( .A(n3293), .B(n3323), .Z(n3285) );
  XNOR U7330 ( .A(n3290), .B(n3292), .Z(n3323) );
  AND U7331 ( .A(n3324), .B(n3325), .Z(n3292) );
  NANDN U7332 ( .A(n3326), .B(n3327), .Z(n3325) );
  NANDN U7333 ( .A(n3328), .B(n3329), .Z(n3327) );
  IV U7334 ( .A(n3330), .Z(n3329) );
  NAND U7335 ( .A(n3330), .B(n3328), .Z(n3324) );
  AND U7336 ( .A(n3331), .B(n3332), .Z(n3290) );
  NAND U7337 ( .A(n3333), .B(n3334), .Z(n3332) );
  OR U7338 ( .A(n3335), .B(n3336), .Z(n3334) );
  NAND U7339 ( .A(n3336), .B(n3335), .Z(n3331) );
  IV U7340 ( .A(n3337), .Z(n3336) );
  NAND U7341 ( .A(n3338), .B(n3339), .Z(n3293) );
  NANDN U7342 ( .A(n3340), .B(n3341), .Z(n3339) );
  NAND U7343 ( .A(n3342), .B(n3343), .Z(n3341) );
  OR U7344 ( .A(n3343), .B(n3342), .Z(n3338) );
  IV U7345 ( .A(n3344), .Z(n3342) );
  XOR U7346 ( .A(n3319), .B(n3345), .Z(N29874) );
  XNOR U7347 ( .A(n3322), .B(n3321), .Z(n3345) );
  XNOR U7348 ( .A(n3333), .B(n3346), .Z(n3321) );
  XOR U7349 ( .A(n3337), .B(n3335), .Z(n3346) );
  XOR U7350 ( .A(n3343), .B(n3347), .Z(n3335) );
  XOR U7351 ( .A(n3340), .B(n3344), .Z(n3347) );
  NAND U7352 ( .A(n3348), .B(n3349), .Z(n3344) );
  NAND U7353 ( .A(n3350), .B(n3351), .Z(n3349) );
  NAND U7354 ( .A(n3352), .B(n3353), .Z(n3348) );
  AND U7355 ( .A(n3354), .B(n3355), .Z(n3340) );
  NAND U7356 ( .A(n3356), .B(n3357), .Z(n3355) );
  NAND U7357 ( .A(n3358), .B(n3359), .Z(n3354) );
  NANDN U7358 ( .A(n3360), .B(n3361), .Z(n3343) );
  NANDN U7359 ( .A(n3362), .B(n3363), .Z(n3337) );
  XNOR U7360 ( .A(n3328), .B(n3364), .Z(n3333) );
  XOR U7361 ( .A(n3326), .B(n3330), .Z(n3364) );
  NAND U7362 ( .A(n3365), .B(n3366), .Z(n3330) );
  NAND U7363 ( .A(n3367), .B(n3368), .Z(n3366) );
  NAND U7364 ( .A(n3369), .B(n3370), .Z(n3365) );
  AND U7365 ( .A(n3371), .B(n3372), .Z(n3326) );
  NAND U7366 ( .A(n3373), .B(n3374), .Z(n3372) );
  NAND U7367 ( .A(n3375), .B(n3376), .Z(n3371) );
  AND U7368 ( .A(n3377), .B(n3378), .Z(n3328) );
  NAND U7369 ( .A(n3379), .B(n3380), .Z(n3322) );
  XNOR U7370 ( .A(n3305), .B(n3381), .Z(n3319) );
  XOR U7371 ( .A(n3309), .B(n3307), .Z(n3381) );
  XOR U7372 ( .A(n3315), .B(n3382), .Z(n3307) );
  XOR U7373 ( .A(n3312), .B(n3316), .Z(n3382) );
  NAND U7374 ( .A(n3383), .B(n3384), .Z(n3316) );
  NAND U7375 ( .A(n3385), .B(n3386), .Z(n3384) );
  NAND U7376 ( .A(n3387), .B(n3388), .Z(n3383) );
  AND U7377 ( .A(n3389), .B(n3390), .Z(n3312) );
  NAND U7378 ( .A(n3391), .B(n3392), .Z(n3390) );
  NAND U7379 ( .A(n3393), .B(n3394), .Z(n3389) );
  NANDN U7380 ( .A(n3395), .B(n3396), .Z(n3315) );
  NANDN U7381 ( .A(n3397), .B(n3398), .Z(n3309) );
  XNOR U7382 ( .A(n3300), .B(n3399), .Z(n3305) );
  XOR U7383 ( .A(n3298), .B(n3302), .Z(n3399) );
  NAND U7384 ( .A(n3400), .B(n3401), .Z(n3302) );
  NAND U7385 ( .A(n3402), .B(n3403), .Z(n3401) );
  NAND U7386 ( .A(n3404), .B(n3405), .Z(n3400) );
  AND U7387 ( .A(n3406), .B(n3407), .Z(n3298) );
  NAND U7388 ( .A(n3408), .B(n3409), .Z(n3407) );
  NAND U7389 ( .A(n3410), .B(n3411), .Z(n3406) );
  AND U7390 ( .A(n3412), .B(n3413), .Z(n3300) );
  XOR U7391 ( .A(n3380), .B(n3379), .Z(N29873) );
  XNOR U7392 ( .A(n3398), .B(n3397), .Z(n3379) );
  XNOR U7393 ( .A(n3412), .B(n3413), .Z(n3397) );
  XOR U7394 ( .A(n3409), .B(n3408), .Z(n3413) );
  XOR U7395 ( .A(y[3891]), .B(x[3891]), .Z(n3408) );
  XOR U7396 ( .A(n3411), .B(n3410), .Z(n3409) );
  XOR U7397 ( .A(y[3893]), .B(x[3893]), .Z(n3410) );
  XOR U7398 ( .A(y[3892]), .B(x[3892]), .Z(n3411) );
  XOR U7399 ( .A(n3403), .B(n3402), .Z(n3412) );
  XOR U7400 ( .A(n3405), .B(n3404), .Z(n3402) );
  XOR U7401 ( .A(y[3890]), .B(x[3890]), .Z(n3404) );
  XOR U7402 ( .A(y[3889]), .B(x[3889]), .Z(n3405) );
  XOR U7403 ( .A(y[3888]), .B(x[3888]), .Z(n3403) );
  XNOR U7404 ( .A(n3396), .B(n3395), .Z(n3398) );
  XNOR U7405 ( .A(n3392), .B(n3391), .Z(n3395) );
  XOR U7406 ( .A(n3394), .B(n3393), .Z(n3391) );
  XOR U7407 ( .A(y[3887]), .B(x[3887]), .Z(n3393) );
  XOR U7408 ( .A(y[3886]), .B(x[3886]), .Z(n3394) );
  XOR U7409 ( .A(y[3885]), .B(x[3885]), .Z(n3392) );
  XOR U7410 ( .A(n3386), .B(n3385), .Z(n3396) );
  XOR U7411 ( .A(n3388), .B(n3387), .Z(n3385) );
  XOR U7412 ( .A(y[3884]), .B(x[3884]), .Z(n3387) );
  XOR U7413 ( .A(y[3883]), .B(x[3883]), .Z(n3388) );
  XOR U7414 ( .A(y[3882]), .B(x[3882]), .Z(n3386) );
  XNOR U7415 ( .A(n3363), .B(n3362), .Z(n3380) );
  XNOR U7416 ( .A(n3377), .B(n3378), .Z(n3362) );
  XOR U7417 ( .A(n3374), .B(n3373), .Z(n3378) );
  XOR U7418 ( .A(y[3879]), .B(x[3879]), .Z(n3373) );
  XOR U7419 ( .A(n3376), .B(n3375), .Z(n3374) );
  XOR U7420 ( .A(y[3881]), .B(x[3881]), .Z(n3375) );
  XOR U7421 ( .A(y[3880]), .B(x[3880]), .Z(n3376) );
  XOR U7422 ( .A(n3368), .B(n3367), .Z(n3377) );
  XOR U7423 ( .A(n3370), .B(n3369), .Z(n3367) );
  XOR U7424 ( .A(y[3878]), .B(x[3878]), .Z(n3369) );
  XOR U7425 ( .A(y[3877]), .B(x[3877]), .Z(n3370) );
  XOR U7426 ( .A(y[3876]), .B(x[3876]), .Z(n3368) );
  XNOR U7427 ( .A(n3361), .B(n3360), .Z(n3363) );
  XNOR U7428 ( .A(n3357), .B(n3356), .Z(n3360) );
  XOR U7429 ( .A(n3359), .B(n3358), .Z(n3356) );
  XOR U7430 ( .A(y[3875]), .B(x[3875]), .Z(n3358) );
  XOR U7431 ( .A(y[3874]), .B(x[3874]), .Z(n3359) );
  XOR U7432 ( .A(y[3873]), .B(x[3873]), .Z(n3357) );
  XOR U7433 ( .A(n3351), .B(n3350), .Z(n3361) );
  XOR U7434 ( .A(n3353), .B(n3352), .Z(n3350) );
  XOR U7435 ( .A(y[3872]), .B(x[3872]), .Z(n3352) );
  XOR U7436 ( .A(y[3871]), .B(x[3871]), .Z(n3353) );
  XOR U7437 ( .A(y[3870]), .B(x[3870]), .Z(n3351) );
  NAND U7438 ( .A(n3414), .B(n3415), .Z(N29865) );
  NAND U7439 ( .A(n3416), .B(n3417), .Z(n3415) );
  NANDN U7440 ( .A(n3418), .B(n3419), .Z(n3417) );
  NANDN U7441 ( .A(n3419), .B(n3418), .Z(n3414) );
  XOR U7442 ( .A(n3418), .B(n3420), .Z(N29864) );
  XNOR U7443 ( .A(n3416), .B(n3419), .Z(n3420) );
  NAND U7444 ( .A(n3421), .B(n3422), .Z(n3419) );
  NAND U7445 ( .A(n3423), .B(n3424), .Z(n3422) );
  NANDN U7446 ( .A(n3425), .B(n3426), .Z(n3424) );
  NANDN U7447 ( .A(n3426), .B(n3425), .Z(n3421) );
  AND U7448 ( .A(n3427), .B(n3428), .Z(n3416) );
  NAND U7449 ( .A(n3429), .B(n3430), .Z(n3428) );
  OR U7450 ( .A(n3431), .B(n3432), .Z(n3430) );
  NAND U7451 ( .A(n3432), .B(n3431), .Z(n3427) );
  IV U7452 ( .A(n3433), .Z(n3432) );
  AND U7453 ( .A(n3434), .B(n3435), .Z(n3418) );
  NAND U7454 ( .A(n3436), .B(n3437), .Z(n3435) );
  NANDN U7455 ( .A(n3438), .B(n3439), .Z(n3437) );
  NANDN U7456 ( .A(n3439), .B(n3438), .Z(n3434) );
  XOR U7457 ( .A(n3431), .B(n3440), .Z(N29863) );
  XOR U7458 ( .A(n3429), .B(n3433), .Z(n3440) );
  XNOR U7459 ( .A(n3426), .B(n3441), .Z(n3433) );
  XNOR U7460 ( .A(n3423), .B(n3425), .Z(n3441) );
  AND U7461 ( .A(n3442), .B(n3443), .Z(n3425) );
  NANDN U7462 ( .A(n3444), .B(n3445), .Z(n3443) );
  NANDN U7463 ( .A(n3446), .B(n3447), .Z(n3445) );
  IV U7464 ( .A(n3448), .Z(n3447) );
  NAND U7465 ( .A(n3448), .B(n3446), .Z(n3442) );
  AND U7466 ( .A(n3449), .B(n3450), .Z(n3423) );
  NAND U7467 ( .A(n3451), .B(n3452), .Z(n3450) );
  OR U7468 ( .A(n3453), .B(n3454), .Z(n3452) );
  NAND U7469 ( .A(n3454), .B(n3453), .Z(n3449) );
  IV U7470 ( .A(n3455), .Z(n3454) );
  NAND U7471 ( .A(n3456), .B(n3457), .Z(n3426) );
  NANDN U7472 ( .A(n3458), .B(n3459), .Z(n3457) );
  NAND U7473 ( .A(n3460), .B(n3461), .Z(n3459) );
  OR U7474 ( .A(n3461), .B(n3460), .Z(n3456) );
  IV U7475 ( .A(n3462), .Z(n3460) );
  AND U7476 ( .A(n3463), .B(n3464), .Z(n3429) );
  NAND U7477 ( .A(n3465), .B(n3466), .Z(n3464) );
  NANDN U7478 ( .A(n3467), .B(n3468), .Z(n3466) );
  NANDN U7479 ( .A(n3468), .B(n3467), .Z(n3463) );
  XOR U7480 ( .A(n3439), .B(n3469), .Z(n3431) );
  XNOR U7481 ( .A(n3436), .B(n3438), .Z(n3469) );
  AND U7482 ( .A(n3470), .B(n3471), .Z(n3438) );
  NANDN U7483 ( .A(n3472), .B(n3473), .Z(n3471) );
  NANDN U7484 ( .A(n3474), .B(n3475), .Z(n3473) );
  IV U7485 ( .A(n3476), .Z(n3475) );
  NAND U7486 ( .A(n3476), .B(n3474), .Z(n3470) );
  AND U7487 ( .A(n3477), .B(n3478), .Z(n3436) );
  NAND U7488 ( .A(n3479), .B(n3480), .Z(n3478) );
  OR U7489 ( .A(n3481), .B(n3482), .Z(n3480) );
  NAND U7490 ( .A(n3482), .B(n3481), .Z(n3477) );
  IV U7491 ( .A(n3483), .Z(n3482) );
  NAND U7492 ( .A(n3484), .B(n3485), .Z(n3439) );
  NANDN U7493 ( .A(n3486), .B(n3487), .Z(n3485) );
  NAND U7494 ( .A(n3488), .B(n3489), .Z(n3487) );
  OR U7495 ( .A(n3489), .B(n3488), .Z(n3484) );
  IV U7496 ( .A(n3490), .Z(n3488) );
  XOR U7497 ( .A(n3465), .B(n3491), .Z(N29862) );
  XNOR U7498 ( .A(n3468), .B(n3467), .Z(n3491) );
  XNOR U7499 ( .A(n3479), .B(n3492), .Z(n3467) );
  XOR U7500 ( .A(n3483), .B(n3481), .Z(n3492) );
  XOR U7501 ( .A(n3489), .B(n3493), .Z(n3481) );
  XOR U7502 ( .A(n3486), .B(n3490), .Z(n3493) );
  NAND U7503 ( .A(n3494), .B(n3495), .Z(n3490) );
  NAND U7504 ( .A(n3496), .B(n3497), .Z(n3495) );
  NAND U7505 ( .A(n3498), .B(n3499), .Z(n3494) );
  AND U7506 ( .A(n3500), .B(n3501), .Z(n3486) );
  NAND U7507 ( .A(n3502), .B(n3503), .Z(n3501) );
  NAND U7508 ( .A(n3504), .B(n3505), .Z(n3500) );
  NANDN U7509 ( .A(n3506), .B(n3507), .Z(n3489) );
  NANDN U7510 ( .A(n3508), .B(n3509), .Z(n3483) );
  XNOR U7511 ( .A(n3474), .B(n3510), .Z(n3479) );
  XOR U7512 ( .A(n3472), .B(n3476), .Z(n3510) );
  NAND U7513 ( .A(n3511), .B(n3512), .Z(n3476) );
  NAND U7514 ( .A(n3513), .B(n3514), .Z(n3512) );
  NAND U7515 ( .A(n3515), .B(n3516), .Z(n3511) );
  AND U7516 ( .A(n3517), .B(n3518), .Z(n3472) );
  NAND U7517 ( .A(n3519), .B(n3520), .Z(n3518) );
  NAND U7518 ( .A(n3521), .B(n3522), .Z(n3517) );
  AND U7519 ( .A(n3523), .B(n3524), .Z(n3474) );
  NAND U7520 ( .A(n3525), .B(n3526), .Z(n3468) );
  XNOR U7521 ( .A(n3451), .B(n3527), .Z(n3465) );
  XOR U7522 ( .A(n3455), .B(n3453), .Z(n3527) );
  XOR U7523 ( .A(n3461), .B(n3528), .Z(n3453) );
  XOR U7524 ( .A(n3458), .B(n3462), .Z(n3528) );
  NAND U7525 ( .A(n3529), .B(n3530), .Z(n3462) );
  NAND U7526 ( .A(n3531), .B(n3532), .Z(n3530) );
  NAND U7527 ( .A(n3533), .B(n3534), .Z(n3529) );
  AND U7528 ( .A(n3535), .B(n3536), .Z(n3458) );
  NAND U7529 ( .A(n3537), .B(n3538), .Z(n3536) );
  NAND U7530 ( .A(n3539), .B(n3540), .Z(n3535) );
  NANDN U7531 ( .A(n3541), .B(n3542), .Z(n3461) );
  NANDN U7532 ( .A(n3543), .B(n3544), .Z(n3455) );
  XNOR U7533 ( .A(n3446), .B(n3545), .Z(n3451) );
  XOR U7534 ( .A(n3444), .B(n3448), .Z(n3545) );
  NAND U7535 ( .A(n3546), .B(n3547), .Z(n3448) );
  NAND U7536 ( .A(n3548), .B(n3549), .Z(n3547) );
  NAND U7537 ( .A(n3550), .B(n3551), .Z(n3546) );
  AND U7538 ( .A(n3552), .B(n3553), .Z(n3444) );
  NAND U7539 ( .A(n3554), .B(n3555), .Z(n3553) );
  NAND U7540 ( .A(n3556), .B(n3557), .Z(n3552) );
  AND U7541 ( .A(n3558), .B(n3559), .Z(n3446) );
  XOR U7542 ( .A(n3526), .B(n3525), .Z(N29861) );
  XNOR U7543 ( .A(n3544), .B(n3543), .Z(n3525) );
  XNOR U7544 ( .A(n3558), .B(n3559), .Z(n3543) );
  XOR U7545 ( .A(n3555), .B(n3554), .Z(n3559) );
  XOR U7546 ( .A(y[3867]), .B(x[3867]), .Z(n3554) );
  XOR U7547 ( .A(n3557), .B(n3556), .Z(n3555) );
  XOR U7548 ( .A(y[3869]), .B(x[3869]), .Z(n3556) );
  XOR U7549 ( .A(y[3868]), .B(x[3868]), .Z(n3557) );
  XOR U7550 ( .A(n3549), .B(n3548), .Z(n3558) );
  XOR U7551 ( .A(n3551), .B(n3550), .Z(n3548) );
  XOR U7552 ( .A(y[3866]), .B(x[3866]), .Z(n3550) );
  XOR U7553 ( .A(y[3865]), .B(x[3865]), .Z(n3551) );
  XOR U7554 ( .A(y[3864]), .B(x[3864]), .Z(n3549) );
  XNOR U7555 ( .A(n3542), .B(n3541), .Z(n3544) );
  XNOR U7556 ( .A(n3538), .B(n3537), .Z(n3541) );
  XOR U7557 ( .A(n3540), .B(n3539), .Z(n3537) );
  XOR U7558 ( .A(y[3863]), .B(x[3863]), .Z(n3539) );
  XOR U7559 ( .A(y[3862]), .B(x[3862]), .Z(n3540) );
  XOR U7560 ( .A(y[3861]), .B(x[3861]), .Z(n3538) );
  XOR U7561 ( .A(n3532), .B(n3531), .Z(n3542) );
  XOR U7562 ( .A(n3534), .B(n3533), .Z(n3531) );
  XOR U7563 ( .A(y[3860]), .B(x[3860]), .Z(n3533) );
  XOR U7564 ( .A(y[3859]), .B(x[3859]), .Z(n3534) );
  XOR U7565 ( .A(y[3858]), .B(x[3858]), .Z(n3532) );
  XNOR U7566 ( .A(n3509), .B(n3508), .Z(n3526) );
  XNOR U7567 ( .A(n3523), .B(n3524), .Z(n3508) );
  XOR U7568 ( .A(n3520), .B(n3519), .Z(n3524) );
  XOR U7569 ( .A(y[3855]), .B(x[3855]), .Z(n3519) );
  XOR U7570 ( .A(n3522), .B(n3521), .Z(n3520) );
  XOR U7571 ( .A(y[3857]), .B(x[3857]), .Z(n3521) );
  XOR U7572 ( .A(y[3856]), .B(x[3856]), .Z(n3522) );
  XOR U7573 ( .A(n3514), .B(n3513), .Z(n3523) );
  XOR U7574 ( .A(n3516), .B(n3515), .Z(n3513) );
  XOR U7575 ( .A(y[3854]), .B(x[3854]), .Z(n3515) );
  XOR U7576 ( .A(y[3853]), .B(x[3853]), .Z(n3516) );
  XOR U7577 ( .A(y[3852]), .B(x[3852]), .Z(n3514) );
  XNOR U7578 ( .A(n3507), .B(n3506), .Z(n3509) );
  XNOR U7579 ( .A(n3503), .B(n3502), .Z(n3506) );
  XOR U7580 ( .A(n3505), .B(n3504), .Z(n3502) );
  XOR U7581 ( .A(y[3851]), .B(x[3851]), .Z(n3504) );
  XOR U7582 ( .A(y[3850]), .B(x[3850]), .Z(n3505) );
  XOR U7583 ( .A(y[3849]), .B(x[3849]), .Z(n3503) );
  XOR U7584 ( .A(n3497), .B(n3496), .Z(n3507) );
  XOR U7585 ( .A(n3499), .B(n3498), .Z(n3496) );
  XOR U7586 ( .A(y[3848]), .B(x[3848]), .Z(n3498) );
  XOR U7587 ( .A(y[3847]), .B(x[3847]), .Z(n3499) );
  XOR U7588 ( .A(y[3846]), .B(x[3846]), .Z(n3497) );
  NAND U7589 ( .A(n3560), .B(n3561), .Z(N29853) );
  NAND U7590 ( .A(n3562), .B(n3563), .Z(n3561) );
  NANDN U7591 ( .A(n3564), .B(n3565), .Z(n3563) );
  NANDN U7592 ( .A(n3565), .B(n3564), .Z(n3560) );
  XOR U7593 ( .A(n3564), .B(n3566), .Z(N29852) );
  XNOR U7594 ( .A(n3562), .B(n3565), .Z(n3566) );
  NAND U7595 ( .A(n3567), .B(n3568), .Z(n3565) );
  NAND U7596 ( .A(n3569), .B(n3570), .Z(n3568) );
  NANDN U7597 ( .A(n3571), .B(n3572), .Z(n3570) );
  NANDN U7598 ( .A(n3572), .B(n3571), .Z(n3567) );
  AND U7599 ( .A(n3573), .B(n3574), .Z(n3562) );
  NAND U7600 ( .A(n3575), .B(n3576), .Z(n3574) );
  OR U7601 ( .A(n3577), .B(n3578), .Z(n3576) );
  NAND U7602 ( .A(n3578), .B(n3577), .Z(n3573) );
  IV U7603 ( .A(n3579), .Z(n3578) );
  AND U7604 ( .A(n3580), .B(n3581), .Z(n3564) );
  NAND U7605 ( .A(n3582), .B(n3583), .Z(n3581) );
  NANDN U7606 ( .A(n3584), .B(n3585), .Z(n3583) );
  NANDN U7607 ( .A(n3585), .B(n3584), .Z(n3580) );
  XOR U7608 ( .A(n3577), .B(n3586), .Z(N29851) );
  XOR U7609 ( .A(n3575), .B(n3579), .Z(n3586) );
  XNOR U7610 ( .A(n3572), .B(n3587), .Z(n3579) );
  XNOR U7611 ( .A(n3569), .B(n3571), .Z(n3587) );
  AND U7612 ( .A(n3588), .B(n3589), .Z(n3571) );
  NANDN U7613 ( .A(n3590), .B(n3591), .Z(n3589) );
  NANDN U7614 ( .A(n3592), .B(n3593), .Z(n3591) );
  IV U7615 ( .A(n3594), .Z(n3593) );
  NAND U7616 ( .A(n3594), .B(n3592), .Z(n3588) );
  AND U7617 ( .A(n3595), .B(n3596), .Z(n3569) );
  NAND U7618 ( .A(n3597), .B(n3598), .Z(n3596) );
  OR U7619 ( .A(n3599), .B(n3600), .Z(n3598) );
  NAND U7620 ( .A(n3600), .B(n3599), .Z(n3595) );
  IV U7621 ( .A(n3601), .Z(n3600) );
  NAND U7622 ( .A(n3602), .B(n3603), .Z(n3572) );
  NANDN U7623 ( .A(n3604), .B(n3605), .Z(n3603) );
  NAND U7624 ( .A(n3606), .B(n3607), .Z(n3605) );
  OR U7625 ( .A(n3607), .B(n3606), .Z(n3602) );
  IV U7626 ( .A(n3608), .Z(n3606) );
  AND U7627 ( .A(n3609), .B(n3610), .Z(n3575) );
  NAND U7628 ( .A(n3611), .B(n3612), .Z(n3610) );
  NANDN U7629 ( .A(n3613), .B(n3614), .Z(n3612) );
  NANDN U7630 ( .A(n3614), .B(n3613), .Z(n3609) );
  XOR U7631 ( .A(n3585), .B(n3615), .Z(n3577) );
  XNOR U7632 ( .A(n3582), .B(n3584), .Z(n3615) );
  AND U7633 ( .A(n3616), .B(n3617), .Z(n3584) );
  NANDN U7634 ( .A(n3618), .B(n3619), .Z(n3617) );
  NANDN U7635 ( .A(n3620), .B(n3621), .Z(n3619) );
  IV U7636 ( .A(n3622), .Z(n3621) );
  NAND U7637 ( .A(n3622), .B(n3620), .Z(n3616) );
  AND U7638 ( .A(n3623), .B(n3624), .Z(n3582) );
  NAND U7639 ( .A(n3625), .B(n3626), .Z(n3624) );
  OR U7640 ( .A(n3627), .B(n3628), .Z(n3626) );
  NAND U7641 ( .A(n3628), .B(n3627), .Z(n3623) );
  IV U7642 ( .A(n3629), .Z(n3628) );
  NAND U7643 ( .A(n3630), .B(n3631), .Z(n3585) );
  NANDN U7644 ( .A(n3632), .B(n3633), .Z(n3631) );
  NAND U7645 ( .A(n3634), .B(n3635), .Z(n3633) );
  OR U7646 ( .A(n3635), .B(n3634), .Z(n3630) );
  IV U7647 ( .A(n3636), .Z(n3634) );
  XOR U7648 ( .A(n3611), .B(n3637), .Z(N29850) );
  XNOR U7649 ( .A(n3614), .B(n3613), .Z(n3637) );
  XNOR U7650 ( .A(n3625), .B(n3638), .Z(n3613) );
  XOR U7651 ( .A(n3629), .B(n3627), .Z(n3638) );
  XOR U7652 ( .A(n3635), .B(n3639), .Z(n3627) );
  XOR U7653 ( .A(n3632), .B(n3636), .Z(n3639) );
  NAND U7654 ( .A(n3640), .B(n3641), .Z(n3636) );
  NAND U7655 ( .A(n3642), .B(n3643), .Z(n3641) );
  NAND U7656 ( .A(n3644), .B(n3645), .Z(n3640) );
  AND U7657 ( .A(n3646), .B(n3647), .Z(n3632) );
  NAND U7658 ( .A(n3648), .B(n3649), .Z(n3647) );
  NAND U7659 ( .A(n3650), .B(n3651), .Z(n3646) );
  NANDN U7660 ( .A(n3652), .B(n3653), .Z(n3635) );
  NANDN U7661 ( .A(n3654), .B(n3655), .Z(n3629) );
  XNOR U7662 ( .A(n3620), .B(n3656), .Z(n3625) );
  XOR U7663 ( .A(n3618), .B(n3622), .Z(n3656) );
  NAND U7664 ( .A(n3657), .B(n3658), .Z(n3622) );
  NAND U7665 ( .A(n3659), .B(n3660), .Z(n3658) );
  NAND U7666 ( .A(n3661), .B(n3662), .Z(n3657) );
  AND U7667 ( .A(n3663), .B(n3664), .Z(n3618) );
  NAND U7668 ( .A(n3665), .B(n3666), .Z(n3664) );
  NAND U7669 ( .A(n3667), .B(n3668), .Z(n3663) );
  AND U7670 ( .A(n3669), .B(n3670), .Z(n3620) );
  NAND U7671 ( .A(n3671), .B(n3672), .Z(n3614) );
  XNOR U7672 ( .A(n3597), .B(n3673), .Z(n3611) );
  XOR U7673 ( .A(n3601), .B(n3599), .Z(n3673) );
  XOR U7674 ( .A(n3607), .B(n3674), .Z(n3599) );
  XOR U7675 ( .A(n3604), .B(n3608), .Z(n3674) );
  NAND U7676 ( .A(n3675), .B(n3676), .Z(n3608) );
  NAND U7677 ( .A(n3677), .B(n3678), .Z(n3676) );
  NAND U7678 ( .A(n3679), .B(n3680), .Z(n3675) );
  AND U7679 ( .A(n3681), .B(n3682), .Z(n3604) );
  NAND U7680 ( .A(n3683), .B(n3684), .Z(n3682) );
  NAND U7681 ( .A(n3685), .B(n3686), .Z(n3681) );
  NANDN U7682 ( .A(n3687), .B(n3688), .Z(n3607) );
  NANDN U7683 ( .A(n3689), .B(n3690), .Z(n3601) );
  XNOR U7684 ( .A(n3592), .B(n3691), .Z(n3597) );
  XOR U7685 ( .A(n3590), .B(n3594), .Z(n3691) );
  NAND U7686 ( .A(n3692), .B(n3693), .Z(n3594) );
  NAND U7687 ( .A(n3694), .B(n3695), .Z(n3693) );
  NAND U7688 ( .A(n3696), .B(n3697), .Z(n3692) );
  AND U7689 ( .A(n3698), .B(n3699), .Z(n3590) );
  NAND U7690 ( .A(n3700), .B(n3701), .Z(n3699) );
  NAND U7691 ( .A(n3702), .B(n3703), .Z(n3698) );
  AND U7692 ( .A(n3704), .B(n3705), .Z(n3592) );
  XOR U7693 ( .A(n3672), .B(n3671), .Z(N29849) );
  XNOR U7694 ( .A(n3690), .B(n3689), .Z(n3671) );
  XNOR U7695 ( .A(n3704), .B(n3705), .Z(n3689) );
  XOR U7696 ( .A(n3701), .B(n3700), .Z(n3705) );
  XOR U7697 ( .A(y[3843]), .B(x[3843]), .Z(n3700) );
  XOR U7698 ( .A(n3703), .B(n3702), .Z(n3701) );
  XOR U7699 ( .A(y[3845]), .B(x[3845]), .Z(n3702) );
  XOR U7700 ( .A(y[3844]), .B(x[3844]), .Z(n3703) );
  XOR U7701 ( .A(n3695), .B(n3694), .Z(n3704) );
  XOR U7702 ( .A(n3697), .B(n3696), .Z(n3694) );
  XOR U7703 ( .A(y[3842]), .B(x[3842]), .Z(n3696) );
  XOR U7704 ( .A(y[3841]), .B(x[3841]), .Z(n3697) );
  XOR U7705 ( .A(y[3840]), .B(x[3840]), .Z(n3695) );
  XNOR U7706 ( .A(n3688), .B(n3687), .Z(n3690) );
  XNOR U7707 ( .A(n3684), .B(n3683), .Z(n3687) );
  XOR U7708 ( .A(n3686), .B(n3685), .Z(n3683) );
  XOR U7709 ( .A(y[3839]), .B(x[3839]), .Z(n3685) );
  XOR U7710 ( .A(y[3838]), .B(x[3838]), .Z(n3686) );
  XOR U7711 ( .A(y[3837]), .B(x[3837]), .Z(n3684) );
  XOR U7712 ( .A(n3678), .B(n3677), .Z(n3688) );
  XOR U7713 ( .A(n3680), .B(n3679), .Z(n3677) );
  XOR U7714 ( .A(y[3836]), .B(x[3836]), .Z(n3679) );
  XOR U7715 ( .A(y[3835]), .B(x[3835]), .Z(n3680) );
  XOR U7716 ( .A(y[3834]), .B(x[3834]), .Z(n3678) );
  XNOR U7717 ( .A(n3655), .B(n3654), .Z(n3672) );
  XNOR U7718 ( .A(n3669), .B(n3670), .Z(n3654) );
  XOR U7719 ( .A(n3666), .B(n3665), .Z(n3670) );
  XOR U7720 ( .A(y[3831]), .B(x[3831]), .Z(n3665) );
  XOR U7721 ( .A(n3668), .B(n3667), .Z(n3666) );
  XOR U7722 ( .A(y[3833]), .B(x[3833]), .Z(n3667) );
  XOR U7723 ( .A(y[3832]), .B(x[3832]), .Z(n3668) );
  XOR U7724 ( .A(n3660), .B(n3659), .Z(n3669) );
  XOR U7725 ( .A(n3662), .B(n3661), .Z(n3659) );
  XOR U7726 ( .A(y[3830]), .B(x[3830]), .Z(n3661) );
  XOR U7727 ( .A(y[3829]), .B(x[3829]), .Z(n3662) );
  XOR U7728 ( .A(y[3828]), .B(x[3828]), .Z(n3660) );
  XNOR U7729 ( .A(n3653), .B(n3652), .Z(n3655) );
  XNOR U7730 ( .A(n3649), .B(n3648), .Z(n3652) );
  XOR U7731 ( .A(n3651), .B(n3650), .Z(n3648) );
  XOR U7732 ( .A(y[3827]), .B(x[3827]), .Z(n3650) );
  XOR U7733 ( .A(y[3826]), .B(x[3826]), .Z(n3651) );
  XOR U7734 ( .A(y[3825]), .B(x[3825]), .Z(n3649) );
  XOR U7735 ( .A(n3643), .B(n3642), .Z(n3653) );
  XOR U7736 ( .A(n3645), .B(n3644), .Z(n3642) );
  XOR U7737 ( .A(y[3824]), .B(x[3824]), .Z(n3644) );
  XOR U7738 ( .A(y[3823]), .B(x[3823]), .Z(n3645) );
  XOR U7739 ( .A(y[3822]), .B(x[3822]), .Z(n3643) );
  NAND U7740 ( .A(n3706), .B(n3707), .Z(N29841) );
  NAND U7741 ( .A(n3708), .B(n3709), .Z(n3707) );
  NANDN U7742 ( .A(n3710), .B(n3711), .Z(n3709) );
  NANDN U7743 ( .A(n3711), .B(n3710), .Z(n3706) );
  XOR U7744 ( .A(n3710), .B(n3712), .Z(N29840) );
  XNOR U7745 ( .A(n3708), .B(n3711), .Z(n3712) );
  NAND U7746 ( .A(n3713), .B(n3714), .Z(n3711) );
  NAND U7747 ( .A(n3715), .B(n3716), .Z(n3714) );
  NANDN U7748 ( .A(n3717), .B(n3718), .Z(n3716) );
  NANDN U7749 ( .A(n3718), .B(n3717), .Z(n3713) );
  AND U7750 ( .A(n3719), .B(n3720), .Z(n3708) );
  NAND U7751 ( .A(n3721), .B(n3722), .Z(n3720) );
  OR U7752 ( .A(n3723), .B(n3724), .Z(n3722) );
  NAND U7753 ( .A(n3724), .B(n3723), .Z(n3719) );
  IV U7754 ( .A(n3725), .Z(n3724) );
  AND U7755 ( .A(n3726), .B(n3727), .Z(n3710) );
  NAND U7756 ( .A(n3728), .B(n3729), .Z(n3727) );
  NANDN U7757 ( .A(n3730), .B(n3731), .Z(n3729) );
  NANDN U7758 ( .A(n3731), .B(n3730), .Z(n3726) );
  XOR U7759 ( .A(n3723), .B(n3732), .Z(N29839) );
  XOR U7760 ( .A(n3721), .B(n3725), .Z(n3732) );
  XNOR U7761 ( .A(n3718), .B(n3733), .Z(n3725) );
  XNOR U7762 ( .A(n3715), .B(n3717), .Z(n3733) );
  AND U7763 ( .A(n3734), .B(n3735), .Z(n3717) );
  NANDN U7764 ( .A(n3736), .B(n3737), .Z(n3735) );
  NANDN U7765 ( .A(n3738), .B(n3739), .Z(n3737) );
  IV U7766 ( .A(n3740), .Z(n3739) );
  NAND U7767 ( .A(n3740), .B(n3738), .Z(n3734) );
  AND U7768 ( .A(n3741), .B(n3742), .Z(n3715) );
  NAND U7769 ( .A(n3743), .B(n3744), .Z(n3742) );
  OR U7770 ( .A(n3745), .B(n3746), .Z(n3744) );
  NAND U7771 ( .A(n3746), .B(n3745), .Z(n3741) );
  IV U7772 ( .A(n3747), .Z(n3746) );
  NAND U7773 ( .A(n3748), .B(n3749), .Z(n3718) );
  NANDN U7774 ( .A(n3750), .B(n3751), .Z(n3749) );
  NAND U7775 ( .A(n3752), .B(n3753), .Z(n3751) );
  OR U7776 ( .A(n3753), .B(n3752), .Z(n3748) );
  IV U7777 ( .A(n3754), .Z(n3752) );
  AND U7778 ( .A(n3755), .B(n3756), .Z(n3721) );
  NAND U7779 ( .A(n3757), .B(n3758), .Z(n3756) );
  NANDN U7780 ( .A(n3759), .B(n3760), .Z(n3758) );
  NANDN U7781 ( .A(n3760), .B(n3759), .Z(n3755) );
  XOR U7782 ( .A(n3731), .B(n3761), .Z(n3723) );
  XNOR U7783 ( .A(n3728), .B(n3730), .Z(n3761) );
  AND U7784 ( .A(n3762), .B(n3763), .Z(n3730) );
  NANDN U7785 ( .A(n3764), .B(n3765), .Z(n3763) );
  NANDN U7786 ( .A(n3766), .B(n3767), .Z(n3765) );
  IV U7787 ( .A(n3768), .Z(n3767) );
  NAND U7788 ( .A(n3768), .B(n3766), .Z(n3762) );
  AND U7789 ( .A(n3769), .B(n3770), .Z(n3728) );
  NAND U7790 ( .A(n3771), .B(n3772), .Z(n3770) );
  OR U7791 ( .A(n3773), .B(n3774), .Z(n3772) );
  NAND U7792 ( .A(n3774), .B(n3773), .Z(n3769) );
  IV U7793 ( .A(n3775), .Z(n3774) );
  NAND U7794 ( .A(n3776), .B(n3777), .Z(n3731) );
  NANDN U7795 ( .A(n3778), .B(n3779), .Z(n3777) );
  NAND U7796 ( .A(n3780), .B(n3781), .Z(n3779) );
  OR U7797 ( .A(n3781), .B(n3780), .Z(n3776) );
  IV U7798 ( .A(n3782), .Z(n3780) );
  XOR U7799 ( .A(n3757), .B(n3783), .Z(N29838) );
  XNOR U7800 ( .A(n3760), .B(n3759), .Z(n3783) );
  XNOR U7801 ( .A(n3771), .B(n3784), .Z(n3759) );
  XOR U7802 ( .A(n3775), .B(n3773), .Z(n3784) );
  XOR U7803 ( .A(n3781), .B(n3785), .Z(n3773) );
  XOR U7804 ( .A(n3778), .B(n3782), .Z(n3785) );
  NAND U7805 ( .A(n3786), .B(n3787), .Z(n3782) );
  NAND U7806 ( .A(n3788), .B(n3789), .Z(n3787) );
  NAND U7807 ( .A(n3790), .B(n3791), .Z(n3786) );
  AND U7808 ( .A(n3792), .B(n3793), .Z(n3778) );
  NAND U7809 ( .A(n3794), .B(n3795), .Z(n3793) );
  NAND U7810 ( .A(n3796), .B(n3797), .Z(n3792) );
  NANDN U7811 ( .A(n3798), .B(n3799), .Z(n3781) );
  NANDN U7812 ( .A(n3800), .B(n3801), .Z(n3775) );
  XNOR U7813 ( .A(n3766), .B(n3802), .Z(n3771) );
  XOR U7814 ( .A(n3764), .B(n3768), .Z(n3802) );
  NAND U7815 ( .A(n3803), .B(n3804), .Z(n3768) );
  NAND U7816 ( .A(n3805), .B(n3806), .Z(n3804) );
  NAND U7817 ( .A(n3807), .B(n3808), .Z(n3803) );
  AND U7818 ( .A(n3809), .B(n3810), .Z(n3764) );
  NAND U7819 ( .A(n3811), .B(n3812), .Z(n3810) );
  NAND U7820 ( .A(n3813), .B(n3814), .Z(n3809) );
  AND U7821 ( .A(n3815), .B(n3816), .Z(n3766) );
  NAND U7822 ( .A(n3817), .B(n3818), .Z(n3760) );
  XNOR U7823 ( .A(n3743), .B(n3819), .Z(n3757) );
  XOR U7824 ( .A(n3747), .B(n3745), .Z(n3819) );
  XOR U7825 ( .A(n3753), .B(n3820), .Z(n3745) );
  XOR U7826 ( .A(n3750), .B(n3754), .Z(n3820) );
  NAND U7827 ( .A(n3821), .B(n3822), .Z(n3754) );
  NAND U7828 ( .A(n3823), .B(n3824), .Z(n3822) );
  NAND U7829 ( .A(n3825), .B(n3826), .Z(n3821) );
  AND U7830 ( .A(n3827), .B(n3828), .Z(n3750) );
  NAND U7831 ( .A(n3829), .B(n3830), .Z(n3828) );
  NAND U7832 ( .A(n3831), .B(n3832), .Z(n3827) );
  NANDN U7833 ( .A(n3833), .B(n3834), .Z(n3753) );
  NANDN U7834 ( .A(n3835), .B(n3836), .Z(n3747) );
  XNOR U7835 ( .A(n3738), .B(n3837), .Z(n3743) );
  XOR U7836 ( .A(n3736), .B(n3740), .Z(n3837) );
  NAND U7837 ( .A(n3838), .B(n3839), .Z(n3740) );
  NAND U7838 ( .A(n3840), .B(n3841), .Z(n3839) );
  NAND U7839 ( .A(n3842), .B(n3843), .Z(n3838) );
  AND U7840 ( .A(n3844), .B(n3845), .Z(n3736) );
  NAND U7841 ( .A(n3846), .B(n3847), .Z(n3845) );
  NAND U7842 ( .A(n3848), .B(n3849), .Z(n3844) );
  AND U7843 ( .A(n3850), .B(n3851), .Z(n3738) );
  XOR U7844 ( .A(n3818), .B(n3817), .Z(N29837) );
  XNOR U7845 ( .A(n3836), .B(n3835), .Z(n3817) );
  XNOR U7846 ( .A(n3850), .B(n3851), .Z(n3835) );
  XOR U7847 ( .A(n3847), .B(n3846), .Z(n3851) );
  XOR U7848 ( .A(y[3819]), .B(x[3819]), .Z(n3846) );
  XOR U7849 ( .A(n3849), .B(n3848), .Z(n3847) );
  XOR U7850 ( .A(y[3821]), .B(x[3821]), .Z(n3848) );
  XOR U7851 ( .A(y[3820]), .B(x[3820]), .Z(n3849) );
  XOR U7852 ( .A(n3841), .B(n3840), .Z(n3850) );
  XOR U7853 ( .A(n3843), .B(n3842), .Z(n3840) );
  XOR U7854 ( .A(y[3818]), .B(x[3818]), .Z(n3842) );
  XOR U7855 ( .A(y[3817]), .B(x[3817]), .Z(n3843) );
  XOR U7856 ( .A(y[3816]), .B(x[3816]), .Z(n3841) );
  XNOR U7857 ( .A(n3834), .B(n3833), .Z(n3836) );
  XNOR U7858 ( .A(n3830), .B(n3829), .Z(n3833) );
  XOR U7859 ( .A(n3832), .B(n3831), .Z(n3829) );
  XOR U7860 ( .A(y[3815]), .B(x[3815]), .Z(n3831) );
  XOR U7861 ( .A(y[3814]), .B(x[3814]), .Z(n3832) );
  XOR U7862 ( .A(y[3813]), .B(x[3813]), .Z(n3830) );
  XOR U7863 ( .A(n3824), .B(n3823), .Z(n3834) );
  XOR U7864 ( .A(n3826), .B(n3825), .Z(n3823) );
  XOR U7865 ( .A(y[3812]), .B(x[3812]), .Z(n3825) );
  XOR U7866 ( .A(y[3811]), .B(x[3811]), .Z(n3826) );
  XOR U7867 ( .A(y[3810]), .B(x[3810]), .Z(n3824) );
  XNOR U7868 ( .A(n3801), .B(n3800), .Z(n3818) );
  XNOR U7869 ( .A(n3815), .B(n3816), .Z(n3800) );
  XOR U7870 ( .A(n3812), .B(n3811), .Z(n3816) );
  XOR U7871 ( .A(y[3807]), .B(x[3807]), .Z(n3811) );
  XOR U7872 ( .A(n3814), .B(n3813), .Z(n3812) );
  XOR U7873 ( .A(y[3809]), .B(x[3809]), .Z(n3813) );
  XOR U7874 ( .A(y[3808]), .B(x[3808]), .Z(n3814) );
  XOR U7875 ( .A(n3806), .B(n3805), .Z(n3815) );
  XOR U7876 ( .A(n3808), .B(n3807), .Z(n3805) );
  XOR U7877 ( .A(y[3806]), .B(x[3806]), .Z(n3807) );
  XOR U7878 ( .A(y[3805]), .B(x[3805]), .Z(n3808) );
  XOR U7879 ( .A(y[3804]), .B(x[3804]), .Z(n3806) );
  XNOR U7880 ( .A(n3799), .B(n3798), .Z(n3801) );
  XNOR U7881 ( .A(n3795), .B(n3794), .Z(n3798) );
  XOR U7882 ( .A(n3797), .B(n3796), .Z(n3794) );
  XOR U7883 ( .A(y[3803]), .B(x[3803]), .Z(n3796) );
  XOR U7884 ( .A(y[3802]), .B(x[3802]), .Z(n3797) );
  XOR U7885 ( .A(y[3801]), .B(x[3801]), .Z(n3795) );
  XOR U7886 ( .A(n3789), .B(n3788), .Z(n3799) );
  XOR U7887 ( .A(n3791), .B(n3790), .Z(n3788) );
  XOR U7888 ( .A(y[3800]), .B(x[3800]), .Z(n3790) );
  XOR U7889 ( .A(y[3799]), .B(x[3799]), .Z(n3791) );
  XOR U7890 ( .A(y[3798]), .B(x[3798]), .Z(n3789) );
  NAND U7891 ( .A(n3852), .B(n3853), .Z(N29829) );
  NAND U7892 ( .A(n3854), .B(n3855), .Z(n3853) );
  NANDN U7893 ( .A(n3856), .B(n3857), .Z(n3855) );
  NANDN U7894 ( .A(n3857), .B(n3856), .Z(n3852) );
  XOR U7895 ( .A(n3856), .B(n3858), .Z(N29828) );
  XNOR U7896 ( .A(n3854), .B(n3857), .Z(n3858) );
  NAND U7897 ( .A(n3859), .B(n3860), .Z(n3857) );
  NAND U7898 ( .A(n3861), .B(n3862), .Z(n3860) );
  NANDN U7899 ( .A(n3863), .B(n3864), .Z(n3862) );
  NANDN U7900 ( .A(n3864), .B(n3863), .Z(n3859) );
  AND U7901 ( .A(n3865), .B(n3866), .Z(n3854) );
  NAND U7902 ( .A(n3867), .B(n3868), .Z(n3866) );
  OR U7903 ( .A(n3869), .B(n3870), .Z(n3868) );
  NAND U7904 ( .A(n3870), .B(n3869), .Z(n3865) );
  IV U7905 ( .A(n3871), .Z(n3870) );
  AND U7906 ( .A(n3872), .B(n3873), .Z(n3856) );
  NAND U7907 ( .A(n3874), .B(n3875), .Z(n3873) );
  NANDN U7908 ( .A(n3876), .B(n3877), .Z(n3875) );
  NANDN U7909 ( .A(n3877), .B(n3876), .Z(n3872) );
  XOR U7910 ( .A(n3869), .B(n3878), .Z(N29827) );
  XOR U7911 ( .A(n3867), .B(n3871), .Z(n3878) );
  XNOR U7912 ( .A(n3864), .B(n3879), .Z(n3871) );
  XNOR U7913 ( .A(n3861), .B(n3863), .Z(n3879) );
  AND U7914 ( .A(n3880), .B(n3881), .Z(n3863) );
  NANDN U7915 ( .A(n3882), .B(n3883), .Z(n3881) );
  NANDN U7916 ( .A(n3884), .B(n3885), .Z(n3883) );
  IV U7917 ( .A(n3886), .Z(n3885) );
  NAND U7918 ( .A(n3886), .B(n3884), .Z(n3880) );
  AND U7919 ( .A(n3887), .B(n3888), .Z(n3861) );
  NAND U7920 ( .A(n3889), .B(n3890), .Z(n3888) );
  OR U7921 ( .A(n3891), .B(n3892), .Z(n3890) );
  NAND U7922 ( .A(n3892), .B(n3891), .Z(n3887) );
  IV U7923 ( .A(n3893), .Z(n3892) );
  NAND U7924 ( .A(n3894), .B(n3895), .Z(n3864) );
  NANDN U7925 ( .A(n3896), .B(n3897), .Z(n3895) );
  NAND U7926 ( .A(n3898), .B(n3899), .Z(n3897) );
  OR U7927 ( .A(n3899), .B(n3898), .Z(n3894) );
  IV U7928 ( .A(n3900), .Z(n3898) );
  AND U7929 ( .A(n3901), .B(n3902), .Z(n3867) );
  NAND U7930 ( .A(n3903), .B(n3904), .Z(n3902) );
  NANDN U7931 ( .A(n3905), .B(n3906), .Z(n3904) );
  NANDN U7932 ( .A(n3906), .B(n3905), .Z(n3901) );
  XOR U7933 ( .A(n3877), .B(n3907), .Z(n3869) );
  XNOR U7934 ( .A(n3874), .B(n3876), .Z(n3907) );
  AND U7935 ( .A(n3908), .B(n3909), .Z(n3876) );
  NANDN U7936 ( .A(n3910), .B(n3911), .Z(n3909) );
  NANDN U7937 ( .A(n3912), .B(n3913), .Z(n3911) );
  IV U7938 ( .A(n3914), .Z(n3913) );
  NAND U7939 ( .A(n3914), .B(n3912), .Z(n3908) );
  AND U7940 ( .A(n3915), .B(n3916), .Z(n3874) );
  NAND U7941 ( .A(n3917), .B(n3918), .Z(n3916) );
  OR U7942 ( .A(n3919), .B(n3920), .Z(n3918) );
  NAND U7943 ( .A(n3920), .B(n3919), .Z(n3915) );
  IV U7944 ( .A(n3921), .Z(n3920) );
  NAND U7945 ( .A(n3922), .B(n3923), .Z(n3877) );
  NANDN U7946 ( .A(n3924), .B(n3925), .Z(n3923) );
  NAND U7947 ( .A(n3926), .B(n3927), .Z(n3925) );
  OR U7948 ( .A(n3927), .B(n3926), .Z(n3922) );
  IV U7949 ( .A(n3928), .Z(n3926) );
  XOR U7950 ( .A(n3903), .B(n3929), .Z(N29826) );
  XNOR U7951 ( .A(n3906), .B(n3905), .Z(n3929) );
  XNOR U7952 ( .A(n3917), .B(n3930), .Z(n3905) );
  XOR U7953 ( .A(n3921), .B(n3919), .Z(n3930) );
  XOR U7954 ( .A(n3927), .B(n3931), .Z(n3919) );
  XOR U7955 ( .A(n3924), .B(n3928), .Z(n3931) );
  NAND U7956 ( .A(n3932), .B(n3933), .Z(n3928) );
  NAND U7957 ( .A(n3934), .B(n3935), .Z(n3933) );
  NAND U7958 ( .A(n3936), .B(n3937), .Z(n3932) );
  AND U7959 ( .A(n3938), .B(n3939), .Z(n3924) );
  NAND U7960 ( .A(n3940), .B(n3941), .Z(n3939) );
  NAND U7961 ( .A(n3942), .B(n3943), .Z(n3938) );
  NANDN U7962 ( .A(n3944), .B(n3945), .Z(n3927) );
  NANDN U7963 ( .A(n3946), .B(n3947), .Z(n3921) );
  XNOR U7964 ( .A(n3912), .B(n3948), .Z(n3917) );
  XOR U7965 ( .A(n3910), .B(n3914), .Z(n3948) );
  NAND U7966 ( .A(n3949), .B(n3950), .Z(n3914) );
  NAND U7967 ( .A(n3951), .B(n3952), .Z(n3950) );
  NAND U7968 ( .A(n3953), .B(n3954), .Z(n3949) );
  AND U7969 ( .A(n3955), .B(n3956), .Z(n3910) );
  NAND U7970 ( .A(n3957), .B(n3958), .Z(n3956) );
  NAND U7971 ( .A(n3959), .B(n3960), .Z(n3955) );
  AND U7972 ( .A(n3961), .B(n3962), .Z(n3912) );
  NAND U7973 ( .A(n3963), .B(n3964), .Z(n3906) );
  XNOR U7974 ( .A(n3889), .B(n3965), .Z(n3903) );
  XOR U7975 ( .A(n3893), .B(n3891), .Z(n3965) );
  XOR U7976 ( .A(n3899), .B(n3966), .Z(n3891) );
  XOR U7977 ( .A(n3896), .B(n3900), .Z(n3966) );
  NAND U7978 ( .A(n3967), .B(n3968), .Z(n3900) );
  NAND U7979 ( .A(n3969), .B(n3970), .Z(n3968) );
  NAND U7980 ( .A(n3971), .B(n3972), .Z(n3967) );
  AND U7981 ( .A(n3973), .B(n3974), .Z(n3896) );
  NAND U7982 ( .A(n3975), .B(n3976), .Z(n3974) );
  NAND U7983 ( .A(n3977), .B(n3978), .Z(n3973) );
  NANDN U7984 ( .A(n3979), .B(n3980), .Z(n3899) );
  NANDN U7985 ( .A(n3981), .B(n3982), .Z(n3893) );
  XNOR U7986 ( .A(n3884), .B(n3983), .Z(n3889) );
  XOR U7987 ( .A(n3882), .B(n3886), .Z(n3983) );
  NAND U7988 ( .A(n3984), .B(n3985), .Z(n3886) );
  NAND U7989 ( .A(n3986), .B(n3987), .Z(n3985) );
  NAND U7990 ( .A(n3988), .B(n3989), .Z(n3984) );
  AND U7991 ( .A(n3990), .B(n3991), .Z(n3882) );
  NAND U7992 ( .A(n3992), .B(n3993), .Z(n3991) );
  NAND U7993 ( .A(n3994), .B(n3995), .Z(n3990) );
  AND U7994 ( .A(n3996), .B(n3997), .Z(n3884) );
  XOR U7995 ( .A(n3964), .B(n3963), .Z(N29825) );
  XNOR U7996 ( .A(n3982), .B(n3981), .Z(n3963) );
  XNOR U7997 ( .A(n3996), .B(n3997), .Z(n3981) );
  XOR U7998 ( .A(n3993), .B(n3992), .Z(n3997) );
  XOR U7999 ( .A(y[3795]), .B(x[3795]), .Z(n3992) );
  XOR U8000 ( .A(n3995), .B(n3994), .Z(n3993) );
  XOR U8001 ( .A(y[3797]), .B(x[3797]), .Z(n3994) );
  XOR U8002 ( .A(y[3796]), .B(x[3796]), .Z(n3995) );
  XOR U8003 ( .A(n3987), .B(n3986), .Z(n3996) );
  XOR U8004 ( .A(n3989), .B(n3988), .Z(n3986) );
  XOR U8005 ( .A(y[3794]), .B(x[3794]), .Z(n3988) );
  XOR U8006 ( .A(y[3793]), .B(x[3793]), .Z(n3989) );
  XOR U8007 ( .A(y[3792]), .B(x[3792]), .Z(n3987) );
  XNOR U8008 ( .A(n3980), .B(n3979), .Z(n3982) );
  XNOR U8009 ( .A(n3976), .B(n3975), .Z(n3979) );
  XOR U8010 ( .A(n3978), .B(n3977), .Z(n3975) );
  XOR U8011 ( .A(y[3791]), .B(x[3791]), .Z(n3977) );
  XOR U8012 ( .A(y[3790]), .B(x[3790]), .Z(n3978) );
  XOR U8013 ( .A(y[3789]), .B(x[3789]), .Z(n3976) );
  XOR U8014 ( .A(n3970), .B(n3969), .Z(n3980) );
  XOR U8015 ( .A(n3972), .B(n3971), .Z(n3969) );
  XOR U8016 ( .A(y[3788]), .B(x[3788]), .Z(n3971) );
  XOR U8017 ( .A(y[3787]), .B(x[3787]), .Z(n3972) );
  XOR U8018 ( .A(y[3786]), .B(x[3786]), .Z(n3970) );
  XNOR U8019 ( .A(n3947), .B(n3946), .Z(n3964) );
  XNOR U8020 ( .A(n3961), .B(n3962), .Z(n3946) );
  XOR U8021 ( .A(n3958), .B(n3957), .Z(n3962) );
  XOR U8022 ( .A(y[3783]), .B(x[3783]), .Z(n3957) );
  XOR U8023 ( .A(n3960), .B(n3959), .Z(n3958) );
  XOR U8024 ( .A(y[3785]), .B(x[3785]), .Z(n3959) );
  XOR U8025 ( .A(y[3784]), .B(x[3784]), .Z(n3960) );
  XOR U8026 ( .A(n3952), .B(n3951), .Z(n3961) );
  XOR U8027 ( .A(n3954), .B(n3953), .Z(n3951) );
  XOR U8028 ( .A(y[3782]), .B(x[3782]), .Z(n3953) );
  XOR U8029 ( .A(y[3781]), .B(x[3781]), .Z(n3954) );
  XOR U8030 ( .A(y[3780]), .B(x[3780]), .Z(n3952) );
  XNOR U8031 ( .A(n3945), .B(n3944), .Z(n3947) );
  XNOR U8032 ( .A(n3941), .B(n3940), .Z(n3944) );
  XOR U8033 ( .A(n3943), .B(n3942), .Z(n3940) );
  XOR U8034 ( .A(y[3779]), .B(x[3779]), .Z(n3942) );
  XOR U8035 ( .A(y[3778]), .B(x[3778]), .Z(n3943) );
  XOR U8036 ( .A(y[3777]), .B(x[3777]), .Z(n3941) );
  XOR U8037 ( .A(n3935), .B(n3934), .Z(n3945) );
  XOR U8038 ( .A(n3937), .B(n3936), .Z(n3934) );
  XOR U8039 ( .A(y[3776]), .B(x[3776]), .Z(n3936) );
  XOR U8040 ( .A(y[3775]), .B(x[3775]), .Z(n3937) );
  XOR U8041 ( .A(y[3774]), .B(x[3774]), .Z(n3935) );
  NAND U8042 ( .A(n3998), .B(n3999), .Z(N29817) );
  NAND U8043 ( .A(n4000), .B(n4001), .Z(n3999) );
  NANDN U8044 ( .A(n4002), .B(n4003), .Z(n4001) );
  NANDN U8045 ( .A(n4003), .B(n4002), .Z(n3998) );
  XOR U8046 ( .A(n4002), .B(n4004), .Z(N29816) );
  XNOR U8047 ( .A(n4000), .B(n4003), .Z(n4004) );
  NAND U8048 ( .A(n4005), .B(n4006), .Z(n4003) );
  NAND U8049 ( .A(n4007), .B(n4008), .Z(n4006) );
  NANDN U8050 ( .A(n4009), .B(n4010), .Z(n4008) );
  NANDN U8051 ( .A(n4010), .B(n4009), .Z(n4005) );
  AND U8052 ( .A(n4011), .B(n4012), .Z(n4000) );
  NAND U8053 ( .A(n4013), .B(n4014), .Z(n4012) );
  OR U8054 ( .A(n4015), .B(n4016), .Z(n4014) );
  NAND U8055 ( .A(n4016), .B(n4015), .Z(n4011) );
  IV U8056 ( .A(n4017), .Z(n4016) );
  AND U8057 ( .A(n4018), .B(n4019), .Z(n4002) );
  NAND U8058 ( .A(n4020), .B(n4021), .Z(n4019) );
  NANDN U8059 ( .A(n4022), .B(n4023), .Z(n4021) );
  NANDN U8060 ( .A(n4023), .B(n4022), .Z(n4018) );
  XOR U8061 ( .A(n4015), .B(n4024), .Z(N29815) );
  XOR U8062 ( .A(n4013), .B(n4017), .Z(n4024) );
  XNOR U8063 ( .A(n4010), .B(n4025), .Z(n4017) );
  XNOR U8064 ( .A(n4007), .B(n4009), .Z(n4025) );
  AND U8065 ( .A(n4026), .B(n4027), .Z(n4009) );
  NANDN U8066 ( .A(n4028), .B(n4029), .Z(n4027) );
  NANDN U8067 ( .A(n4030), .B(n4031), .Z(n4029) );
  IV U8068 ( .A(n4032), .Z(n4031) );
  NAND U8069 ( .A(n4032), .B(n4030), .Z(n4026) );
  AND U8070 ( .A(n4033), .B(n4034), .Z(n4007) );
  NAND U8071 ( .A(n4035), .B(n4036), .Z(n4034) );
  OR U8072 ( .A(n4037), .B(n4038), .Z(n4036) );
  NAND U8073 ( .A(n4038), .B(n4037), .Z(n4033) );
  IV U8074 ( .A(n4039), .Z(n4038) );
  NAND U8075 ( .A(n4040), .B(n4041), .Z(n4010) );
  NANDN U8076 ( .A(n4042), .B(n4043), .Z(n4041) );
  NAND U8077 ( .A(n4044), .B(n4045), .Z(n4043) );
  OR U8078 ( .A(n4045), .B(n4044), .Z(n4040) );
  IV U8079 ( .A(n4046), .Z(n4044) );
  AND U8080 ( .A(n4047), .B(n4048), .Z(n4013) );
  NAND U8081 ( .A(n4049), .B(n4050), .Z(n4048) );
  NANDN U8082 ( .A(n4051), .B(n4052), .Z(n4050) );
  NANDN U8083 ( .A(n4052), .B(n4051), .Z(n4047) );
  XOR U8084 ( .A(n4023), .B(n4053), .Z(n4015) );
  XNOR U8085 ( .A(n4020), .B(n4022), .Z(n4053) );
  AND U8086 ( .A(n4054), .B(n4055), .Z(n4022) );
  NANDN U8087 ( .A(n4056), .B(n4057), .Z(n4055) );
  NANDN U8088 ( .A(n4058), .B(n4059), .Z(n4057) );
  IV U8089 ( .A(n4060), .Z(n4059) );
  NAND U8090 ( .A(n4060), .B(n4058), .Z(n4054) );
  AND U8091 ( .A(n4061), .B(n4062), .Z(n4020) );
  NAND U8092 ( .A(n4063), .B(n4064), .Z(n4062) );
  OR U8093 ( .A(n4065), .B(n4066), .Z(n4064) );
  NAND U8094 ( .A(n4066), .B(n4065), .Z(n4061) );
  IV U8095 ( .A(n4067), .Z(n4066) );
  NAND U8096 ( .A(n4068), .B(n4069), .Z(n4023) );
  NANDN U8097 ( .A(n4070), .B(n4071), .Z(n4069) );
  NAND U8098 ( .A(n4072), .B(n4073), .Z(n4071) );
  OR U8099 ( .A(n4073), .B(n4072), .Z(n4068) );
  IV U8100 ( .A(n4074), .Z(n4072) );
  XOR U8101 ( .A(n4049), .B(n4075), .Z(N29814) );
  XNOR U8102 ( .A(n4052), .B(n4051), .Z(n4075) );
  XNOR U8103 ( .A(n4063), .B(n4076), .Z(n4051) );
  XOR U8104 ( .A(n4067), .B(n4065), .Z(n4076) );
  XOR U8105 ( .A(n4073), .B(n4077), .Z(n4065) );
  XOR U8106 ( .A(n4070), .B(n4074), .Z(n4077) );
  NAND U8107 ( .A(n4078), .B(n4079), .Z(n4074) );
  NAND U8108 ( .A(n4080), .B(n4081), .Z(n4079) );
  NAND U8109 ( .A(n4082), .B(n4083), .Z(n4078) );
  AND U8110 ( .A(n4084), .B(n4085), .Z(n4070) );
  NAND U8111 ( .A(n4086), .B(n4087), .Z(n4085) );
  NAND U8112 ( .A(n4088), .B(n4089), .Z(n4084) );
  NANDN U8113 ( .A(n4090), .B(n4091), .Z(n4073) );
  NANDN U8114 ( .A(n4092), .B(n4093), .Z(n4067) );
  XNOR U8115 ( .A(n4058), .B(n4094), .Z(n4063) );
  XOR U8116 ( .A(n4056), .B(n4060), .Z(n4094) );
  NAND U8117 ( .A(n4095), .B(n4096), .Z(n4060) );
  NAND U8118 ( .A(n4097), .B(n4098), .Z(n4096) );
  NAND U8119 ( .A(n4099), .B(n4100), .Z(n4095) );
  AND U8120 ( .A(n4101), .B(n4102), .Z(n4056) );
  NAND U8121 ( .A(n4103), .B(n4104), .Z(n4102) );
  NAND U8122 ( .A(n4105), .B(n4106), .Z(n4101) );
  AND U8123 ( .A(n4107), .B(n4108), .Z(n4058) );
  NAND U8124 ( .A(n4109), .B(n4110), .Z(n4052) );
  XNOR U8125 ( .A(n4035), .B(n4111), .Z(n4049) );
  XOR U8126 ( .A(n4039), .B(n4037), .Z(n4111) );
  XOR U8127 ( .A(n4045), .B(n4112), .Z(n4037) );
  XOR U8128 ( .A(n4042), .B(n4046), .Z(n4112) );
  NAND U8129 ( .A(n4113), .B(n4114), .Z(n4046) );
  NAND U8130 ( .A(n4115), .B(n4116), .Z(n4114) );
  NAND U8131 ( .A(n4117), .B(n4118), .Z(n4113) );
  AND U8132 ( .A(n4119), .B(n4120), .Z(n4042) );
  NAND U8133 ( .A(n4121), .B(n4122), .Z(n4120) );
  NAND U8134 ( .A(n4123), .B(n4124), .Z(n4119) );
  NANDN U8135 ( .A(n4125), .B(n4126), .Z(n4045) );
  NANDN U8136 ( .A(n4127), .B(n4128), .Z(n4039) );
  XNOR U8137 ( .A(n4030), .B(n4129), .Z(n4035) );
  XOR U8138 ( .A(n4028), .B(n4032), .Z(n4129) );
  NAND U8139 ( .A(n4130), .B(n4131), .Z(n4032) );
  NAND U8140 ( .A(n4132), .B(n4133), .Z(n4131) );
  NAND U8141 ( .A(n4134), .B(n4135), .Z(n4130) );
  AND U8142 ( .A(n4136), .B(n4137), .Z(n4028) );
  NAND U8143 ( .A(n4138), .B(n4139), .Z(n4137) );
  NAND U8144 ( .A(n4140), .B(n4141), .Z(n4136) );
  AND U8145 ( .A(n4142), .B(n4143), .Z(n4030) );
  XOR U8146 ( .A(n4110), .B(n4109), .Z(N29813) );
  XNOR U8147 ( .A(n4128), .B(n4127), .Z(n4109) );
  XNOR U8148 ( .A(n4142), .B(n4143), .Z(n4127) );
  XOR U8149 ( .A(n4139), .B(n4138), .Z(n4143) );
  XOR U8150 ( .A(y[3771]), .B(x[3771]), .Z(n4138) );
  XOR U8151 ( .A(n4141), .B(n4140), .Z(n4139) );
  XOR U8152 ( .A(y[3773]), .B(x[3773]), .Z(n4140) );
  XOR U8153 ( .A(y[3772]), .B(x[3772]), .Z(n4141) );
  XOR U8154 ( .A(n4133), .B(n4132), .Z(n4142) );
  XOR U8155 ( .A(n4135), .B(n4134), .Z(n4132) );
  XOR U8156 ( .A(y[3770]), .B(x[3770]), .Z(n4134) );
  XOR U8157 ( .A(y[3769]), .B(x[3769]), .Z(n4135) );
  XOR U8158 ( .A(y[3768]), .B(x[3768]), .Z(n4133) );
  XNOR U8159 ( .A(n4126), .B(n4125), .Z(n4128) );
  XNOR U8160 ( .A(n4122), .B(n4121), .Z(n4125) );
  XOR U8161 ( .A(n4124), .B(n4123), .Z(n4121) );
  XOR U8162 ( .A(y[3767]), .B(x[3767]), .Z(n4123) );
  XOR U8163 ( .A(y[3766]), .B(x[3766]), .Z(n4124) );
  XOR U8164 ( .A(y[3765]), .B(x[3765]), .Z(n4122) );
  XOR U8165 ( .A(n4116), .B(n4115), .Z(n4126) );
  XOR U8166 ( .A(n4118), .B(n4117), .Z(n4115) );
  XOR U8167 ( .A(y[3764]), .B(x[3764]), .Z(n4117) );
  XOR U8168 ( .A(y[3763]), .B(x[3763]), .Z(n4118) );
  XOR U8169 ( .A(y[3762]), .B(x[3762]), .Z(n4116) );
  XNOR U8170 ( .A(n4093), .B(n4092), .Z(n4110) );
  XNOR U8171 ( .A(n4107), .B(n4108), .Z(n4092) );
  XOR U8172 ( .A(n4104), .B(n4103), .Z(n4108) );
  XOR U8173 ( .A(y[3759]), .B(x[3759]), .Z(n4103) );
  XOR U8174 ( .A(n4106), .B(n4105), .Z(n4104) );
  XOR U8175 ( .A(y[3761]), .B(x[3761]), .Z(n4105) );
  XOR U8176 ( .A(y[3760]), .B(x[3760]), .Z(n4106) );
  XOR U8177 ( .A(n4098), .B(n4097), .Z(n4107) );
  XOR U8178 ( .A(n4100), .B(n4099), .Z(n4097) );
  XOR U8179 ( .A(y[3758]), .B(x[3758]), .Z(n4099) );
  XOR U8180 ( .A(y[3757]), .B(x[3757]), .Z(n4100) );
  XOR U8181 ( .A(y[3756]), .B(x[3756]), .Z(n4098) );
  XNOR U8182 ( .A(n4091), .B(n4090), .Z(n4093) );
  XNOR U8183 ( .A(n4087), .B(n4086), .Z(n4090) );
  XOR U8184 ( .A(n4089), .B(n4088), .Z(n4086) );
  XOR U8185 ( .A(y[3755]), .B(x[3755]), .Z(n4088) );
  XOR U8186 ( .A(y[3754]), .B(x[3754]), .Z(n4089) );
  XOR U8187 ( .A(y[3753]), .B(x[3753]), .Z(n4087) );
  XOR U8188 ( .A(n4081), .B(n4080), .Z(n4091) );
  XOR U8189 ( .A(n4083), .B(n4082), .Z(n4080) );
  XOR U8190 ( .A(y[3752]), .B(x[3752]), .Z(n4082) );
  XOR U8191 ( .A(y[3751]), .B(x[3751]), .Z(n4083) );
  XOR U8192 ( .A(y[3750]), .B(x[3750]), .Z(n4081) );
  NAND U8193 ( .A(n4144), .B(n4145), .Z(N29805) );
  NAND U8194 ( .A(n4146), .B(n4147), .Z(n4145) );
  NANDN U8195 ( .A(n4148), .B(n4149), .Z(n4147) );
  NANDN U8196 ( .A(n4149), .B(n4148), .Z(n4144) );
  XOR U8197 ( .A(n4148), .B(n4150), .Z(N29804) );
  XNOR U8198 ( .A(n4146), .B(n4149), .Z(n4150) );
  NAND U8199 ( .A(n4151), .B(n4152), .Z(n4149) );
  NAND U8200 ( .A(n4153), .B(n4154), .Z(n4152) );
  NANDN U8201 ( .A(n4155), .B(n4156), .Z(n4154) );
  NANDN U8202 ( .A(n4156), .B(n4155), .Z(n4151) );
  AND U8203 ( .A(n4157), .B(n4158), .Z(n4146) );
  NAND U8204 ( .A(n4159), .B(n4160), .Z(n4158) );
  OR U8205 ( .A(n4161), .B(n4162), .Z(n4160) );
  NAND U8206 ( .A(n4162), .B(n4161), .Z(n4157) );
  IV U8207 ( .A(n4163), .Z(n4162) );
  AND U8208 ( .A(n4164), .B(n4165), .Z(n4148) );
  NAND U8209 ( .A(n4166), .B(n4167), .Z(n4165) );
  NANDN U8210 ( .A(n4168), .B(n4169), .Z(n4167) );
  NANDN U8211 ( .A(n4169), .B(n4168), .Z(n4164) );
  XOR U8212 ( .A(n4161), .B(n4170), .Z(N29803) );
  XOR U8213 ( .A(n4159), .B(n4163), .Z(n4170) );
  XNOR U8214 ( .A(n4156), .B(n4171), .Z(n4163) );
  XNOR U8215 ( .A(n4153), .B(n4155), .Z(n4171) );
  AND U8216 ( .A(n4172), .B(n4173), .Z(n4155) );
  NANDN U8217 ( .A(n4174), .B(n4175), .Z(n4173) );
  NANDN U8218 ( .A(n4176), .B(n4177), .Z(n4175) );
  IV U8219 ( .A(n4178), .Z(n4177) );
  NAND U8220 ( .A(n4178), .B(n4176), .Z(n4172) );
  AND U8221 ( .A(n4179), .B(n4180), .Z(n4153) );
  NAND U8222 ( .A(n4181), .B(n4182), .Z(n4180) );
  OR U8223 ( .A(n4183), .B(n4184), .Z(n4182) );
  NAND U8224 ( .A(n4184), .B(n4183), .Z(n4179) );
  IV U8225 ( .A(n4185), .Z(n4184) );
  NAND U8226 ( .A(n4186), .B(n4187), .Z(n4156) );
  NANDN U8227 ( .A(n4188), .B(n4189), .Z(n4187) );
  NAND U8228 ( .A(n4190), .B(n4191), .Z(n4189) );
  OR U8229 ( .A(n4191), .B(n4190), .Z(n4186) );
  IV U8230 ( .A(n4192), .Z(n4190) );
  AND U8231 ( .A(n4193), .B(n4194), .Z(n4159) );
  NAND U8232 ( .A(n4195), .B(n4196), .Z(n4194) );
  NANDN U8233 ( .A(n4197), .B(n4198), .Z(n4196) );
  NANDN U8234 ( .A(n4198), .B(n4197), .Z(n4193) );
  XOR U8235 ( .A(n4169), .B(n4199), .Z(n4161) );
  XNOR U8236 ( .A(n4166), .B(n4168), .Z(n4199) );
  AND U8237 ( .A(n4200), .B(n4201), .Z(n4168) );
  NANDN U8238 ( .A(n4202), .B(n4203), .Z(n4201) );
  NANDN U8239 ( .A(n4204), .B(n4205), .Z(n4203) );
  IV U8240 ( .A(n4206), .Z(n4205) );
  NAND U8241 ( .A(n4206), .B(n4204), .Z(n4200) );
  AND U8242 ( .A(n4207), .B(n4208), .Z(n4166) );
  NAND U8243 ( .A(n4209), .B(n4210), .Z(n4208) );
  OR U8244 ( .A(n4211), .B(n4212), .Z(n4210) );
  NAND U8245 ( .A(n4212), .B(n4211), .Z(n4207) );
  IV U8246 ( .A(n4213), .Z(n4212) );
  NAND U8247 ( .A(n4214), .B(n4215), .Z(n4169) );
  NANDN U8248 ( .A(n4216), .B(n4217), .Z(n4215) );
  NAND U8249 ( .A(n4218), .B(n4219), .Z(n4217) );
  OR U8250 ( .A(n4219), .B(n4218), .Z(n4214) );
  IV U8251 ( .A(n4220), .Z(n4218) );
  XOR U8252 ( .A(n4195), .B(n4221), .Z(N29802) );
  XNOR U8253 ( .A(n4198), .B(n4197), .Z(n4221) );
  XNOR U8254 ( .A(n4209), .B(n4222), .Z(n4197) );
  XOR U8255 ( .A(n4213), .B(n4211), .Z(n4222) );
  XOR U8256 ( .A(n4219), .B(n4223), .Z(n4211) );
  XOR U8257 ( .A(n4216), .B(n4220), .Z(n4223) );
  NAND U8258 ( .A(n4224), .B(n4225), .Z(n4220) );
  NAND U8259 ( .A(n4226), .B(n4227), .Z(n4225) );
  NAND U8260 ( .A(n4228), .B(n4229), .Z(n4224) );
  AND U8261 ( .A(n4230), .B(n4231), .Z(n4216) );
  NAND U8262 ( .A(n4232), .B(n4233), .Z(n4231) );
  NAND U8263 ( .A(n4234), .B(n4235), .Z(n4230) );
  NANDN U8264 ( .A(n4236), .B(n4237), .Z(n4219) );
  NANDN U8265 ( .A(n4238), .B(n4239), .Z(n4213) );
  XNOR U8266 ( .A(n4204), .B(n4240), .Z(n4209) );
  XOR U8267 ( .A(n4202), .B(n4206), .Z(n4240) );
  NAND U8268 ( .A(n4241), .B(n4242), .Z(n4206) );
  NAND U8269 ( .A(n4243), .B(n4244), .Z(n4242) );
  NAND U8270 ( .A(n4245), .B(n4246), .Z(n4241) );
  AND U8271 ( .A(n4247), .B(n4248), .Z(n4202) );
  NAND U8272 ( .A(n4249), .B(n4250), .Z(n4248) );
  NAND U8273 ( .A(n4251), .B(n4252), .Z(n4247) );
  AND U8274 ( .A(n4253), .B(n4254), .Z(n4204) );
  NAND U8275 ( .A(n4255), .B(n4256), .Z(n4198) );
  XNOR U8276 ( .A(n4181), .B(n4257), .Z(n4195) );
  XOR U8277 ( .A(n4185), .B(n4183), .Z(n4257) );
  XOR U8278 ( .A(n4191), .B(n4258), .Z(n4183) );
  XOR U8279 ( .A(n4188), .B(n4192), .Z(n4258) );
  NAND U8280 ( .A(n4259), .B(n4260), .Z(n4192) );
  NAND U8281 ( .A(n4261), .B(n4262), .Z(n4260) );
  NAND U8282 ( .A(n4263), .B(n4264), .Z(n4259) );
  AND U8283 ( .A(n4265), .B(n4266), .Z(n4188) );
  NAND U8284 ( .A(n4267), .B(n4268), .Z(n4266) );
  NAND U8285 ( .A(n4269), .B(n4270), .Z(n4265) );
  NANDN U8286 ( .A(n4271), .B(n4272), .Z(n4191) );
  NANDN U8287 ( .A(n4273), .B(n4274), .Z(n4185) );
  XNOR U8288 ( .A(n4176), .B(n4275), .Z(n4181) );
  XOR U8289 ( .A(n4174), .B(n4178), .Z(n4275) );
  NAND U8290 ( .A(n4276), .B(n4277), .Z(n4178) );
  NAND U8291 ( .A(n4278), .B(n4279), .Z(n4277) );
  NAND U8292 ( .A(n4280), .B(n4281), .Z(n4276) );
  AND U8293 ( .A(n4282), .B(n4283), .Z(n4174) );
  NAND U8294 ( .A(n4284), .B(n4285), .Z(n4283) );
  NAND U8295 ( .A(n4286), .B(n4287), .Z(n4282) );
  AND U8296 ( .A(n4288), .B(n4289), .Z(n4176) );
  XOR U8297 ( .A(n4256), .B(n4255), .Z(N29801) );
  XNOR U8298 ( .A(n4274), .B(n4273), .Z(n4255) );
  XNOR U8299 ( .A(n4288), .B(n4289), .Z(n4273) );
  XOR U8300 ( .A(n4285), .B(n4284), .Z(n4289) );
  XOR U8301 ( .A(y[3747]), .B(x[3747]), .Z(n4284) );
  XOR U8302 ( .A(n4287), .B(n4286), .Z(n4285) );
  XOR U8303 ( .A(y[3749]), .B(x[3749]), .Z(n4286) );
  XOR U8304 ( .A(y[3748]), .B(x[3748]), .Z(n4287) );
  XOR U8305 ( .A(n4279), .B(n4278), .Z(n4288) );
  XOR U8306 ( .A(n4281), .B(n4280), .Z(n4278) );
  XOR U8307 ( .A(y[3746]), .B(x[3746]), .Z(n4280) );
  XOR U8308 ( .A(y[3745]), .B(x[3745]), .Z(n4281) );
  XOR U8309 ( .A(y[3744]), .B(x[3744]), .Z(n4279) );
  XNOR U8310 ( .A(n4272), .B(n4271), .Z(n4274) );
  XNOR U8311 ( .A(n4268), .B(n4267), .Z(n4271) );
  XOR U8312 ( .A(n4270), .B(n4269), .Z(n4267) );
  XOR U8313 ( .A(y[3743]), .B(x[3743]), .Z(n4269) );
  XOR U8314 ( .A(y[3742]), .B(x[3742]), .Z(n4270) );
  XOR U8315 ( .A(y[3741]), .B(x[3741]), .Z(n4268) );
  XOR U8316 ( .A(n4262), .B(n4261), .Z(n4272) );
  XOR U8317 ( .A(n4264), .B(n4263), .Z(n4261) );
  XOR U8318 ( .A(y[3740]), .B(x[3740]), .Z(n4263) );
  XOR U8319 ( .A(y[3739]), .B(x[3739]), .Z(n4264) );
  XOR U8320 ( .A(y[3738]), .B(x[3738]), .Z(n4262) );
  XNOR U8321 ( .A(n4239), .B(n4238), .Z(n4256) );
  XNOR U8322 ( .A(n4253), .B(n4254), .Z(n4238) );
  XOR U8323 ( .A(n4250), .B(n4249), .Z(n4254) );
  XOR U8324 ( .A(y[3735]), .B(x[3735]), .Z(n4249) );
  XOR U8325 ( .A(n4252), .B(n4251), .Z(n4250) );
  XOR U8326 ( .A(y[3737]), .B(x[3737]), .Z(n4251) );
  XOR U8327 ( .A(y[3736]), .B(x[3736]), .Z(n4252) );
  XOR U8328 ( .A(n4244), .B(n4243), .Z(n4253) );
  XOR U8329 ( .A(n4246), .B(n4245), .Z(n4243) );
  XOR U8330 ( .A(y[3734]), .B(x[3734]), .Z(n4245) );
  XOR U8331 ( .A(y[3733]), .B(x[3733]), .Z(n4246) );
  XOR U8332 ( .A(y[3732]), .B(x[3732]), .Z(n4244) );
  XNOR U8333 ( .A(n4237), .B(n4236), .Z(n4239) );
  XNOR U8334 ( .A(n4233), .B(n4232), .Z(n4236) );
  XOR U8335 ( .A(n4235), .B(n4234), .Z(n4232) );
  XOR U8336 ( .A(y[3731]), .B(x[3731]), .Z(n4234) );
  XOR U8337 ( .A(y[3730]), .B(x[3730]), .Z(n4235) );
  XOR U8338 ( .A(y[3729]), .B(x[3729]), .Z(n4233) );
  XOR U8339 ( .A(n4227), .B(n4226), .Z(n4237) );
  XOR U8340 ( .A(n4229), .B(n4228), .Z(n4226) );
  XOR U8341 ( .A(y[3728]), .B(x[3728]), .Z(n4228) );
  XOR U8342 ( .A(y[3727]), .B(x[3727]), .Z(n4229) );
  XOR U8343 ( .A(y[3726]), .B(x[3726]), .Z(n4227) );
  NAND U8344 ( .A(n4290), .B(n4291), .Z(N29793) );
  NAND U8345 ( .A(n4292), .B(n4293), .Z(n4291) );
  NANDN U8346 ( .A(n4294), .B(n4295), .Z(n4293) );
  NANDN U8347 ( .A(n4295), .B(n4294), .Z(n4290) );
  XOR U8348 ( .A(n4294), .B(n4296), .Z(N29792) );
  XNOR U8349 ( .A(n4292), .B(n4295), .Z(n4296) );
  NAND U8350 ( .A(n4297), .B(n4298), .Z(n4295) );
  NAND U8351 ( .A(n4299), .B(n4300), .Z(n4298) );
  NANDN U8352 ( .A(n4301), .B(n4302), .Z(n4300) );
  NANDN U8353 ( .A(n4302), .B(n4301), .Z(n4297) );
  AND U8354 ( .A(n4303), .B(n4304), .Z(n4292) );
  NAND U8355 ( .A(n4305), .B(n4306), .Z(n4304) );
  OR U8356 ( .A(n4307), .B(n4308), .Z(n4306) );
  NAND U8357 ( .A(n4308), .B(n4307), .Z(n4303) );
  IV U8358 ( .A(n4309), .Z(n4308) );
  AND U8359 ( .A(n4310), .B(n4311), .Z(n4294) );
  NAND U8360 ( .A(n4312), .B(n4313), .Z(n4311) );
  NANDN U8361 ( .A(n4314), .B(n4315), .Z(n4313) );
  NANDN U8362 ( .A(n4315), .B(n4314), .Z(n4310) );
  XOR U8363 ( .A(n4307), .B(n4316), .Z(N29791) );
  XOR U8364 ( .A(n4305), .B(n4309), .Z(n4316) );
  XNOR U8365 ( .A(n4302), .B(n4317), .Z(n4309) );
  XNOR U8366 ( .A(n4299), .B(n4301), .Z(n4317) );
  AND U8367 ( .A(n4318), .B(n4319), .Z(n4301) );
  NANDN U8368 ( .A(n4320), .B(n4321), .Z(n4319) );
  NANDN U8369 ( .A(n4322), .B(n4323), .Z(n4321) );
  IV U8370 ( .A(n4324), .Z(n4323) );
  NAND U8371 ( .A(n4324), .B(n4322), .Z(n4318) );
  AND U8372 ( .A(n4325), .B(n4326), .Z(n4299) );
  NAND U8373 ( .A(n4327), .B(n4328), .Z(n4326) );
  OR U8374 ( .A(n4329), .B(n4330), .Z(n4328) );
  NAND U8375 ( .A(n4330), .B(n4329), .Z(n4325) );
  IV U8376 ( .A(n4331), .Z(n4330) );
  NAND U8377 ( .A(n4332), .B(n4333), .Z(n4302) );
  NANDN U8378 ( .A(n4334), .B(n4335), .Z(n4333) );
  NAND U8379 ( .A(n4336), .B(n4337), .Z(n4335) );
  OR U8380 ( .A(n4337), .B(n4336), .Z(n4332) );
  IV U8381 ( .A(n4338), .Z(n4336) );
  AND U8382 ( .A(n4339), .B(n4340), .Z(n4305) );
  NAND U8383 ( .A(n4341), .B(n4342), .Z(n4340) );
  NANDN U8384 ( .A(n4343), .B(n4344), .Z(n4342) );
  NANDN U8385 ( .A(n4344), .B(n4343), .Z(n4339) );
  XOR U8386 ( .A(n4315), .B(n4345), .Z(n4307) );
  XNOR U8387 ( .A(n4312), .B(n4314), .Z(n4345) );
  AND U8388 ( .A(n4346), .B(n4347), .Z(n4314) );
  NANDN U8389 ( .A(n4348), .B(n4349), .Z(n4347) );
  NANDN U8390 ( .A(n4350), .B(n4351), .Z(n4349) );
  IV U8391 ( .A(n4352), .Z(n4351) );
  NAND U8392 ( .A(n4352), .B(n4350), .Z(n4346) );
  AND U8393 ( .A(n4353), .B(n4354), .Z(n4312) );
  NAND U8394 ( .A(n4355), .B(n4356), .Z(n4354) );
  OR U8395 ( .A(n4357), .B(n4358), .Z(n4356) );
  NAND U8396 ( .A(n4358), .B(n4357), .Z(n4353) );
  IV U8397 ( .A(n4359), .Z(n4358) );
  NAND U8398 ( .A(n4360), .B(n4361), .Z(n4315) );
  NANDN U8399 ( .A(n4362), .B(n4363), .Z(n4361) );
  NAND U8400 ( .A(n4364), .B(n4365), .Z(n4363) );
  OR U8401 ( .A(n4365), .B(n4364), .Z(n4360) );
  IV U8402 ( .A(n4366), .Z(n4364) );
  XOR U8403 ( .A(n4341), .B(n4367), .Z(N29790) );
  XNOR U8404 ( .A(n4344), .B(n4343), .Z(n4367) );
  XNOR U8405 ( .A(n4355), .B(n4368), .Z(n4343) );
  XOR U8406 ( .A(n4359), .B(n4357), .Z(n4368) );
  XOR U8407 ( .A(n4365), .B(n4369), .Z(n4357) );
  XOR U8408 ( .A(n4362), .B(n4366), .Z(n4369) );
  NAND U8409 ( .A(n4370), .B(n4371), .Z(n4366) );
  NAND U8410 ( .A(n4372), .B(n4373), .Z(n4371) );
  NAND U8411 ( .A(n4374), .B(n4375), .Z(n4370) );
  AND U8412 ( .A(n4376), .B(n4377), .Z(n4362) );
  NAND U8413 ( .A(n4378), .B(n4379), .Z(n4377) );
  NAND U8414 ( .A(n4380), .B(n4381), .Z(n4376) );
  NANDN U8415 ( .A(n4382), .B(n4383), .Z(n4365) );
  NANDN U8416 ( .A(n4384), .B(n4385), .Z(n4359) );
  XNOR U8417 ( .A(n4350), .B(n4386), .Z(n4355) );
  XOR U8418 ( .A(n4348), .B(n4352), .Z(n4386) );
  NAND U8419 ( .A(n4387), .B(n4388), .Z(n4352) );
  NAND U8420 ( .A(n4389), .B(n4390), .Z(n4388) );
  NAND U8421 ( .A(n4391), .B(n4392), .Z(n4387) );
  AND U8422 ( .A(n4393), .B(n4394), .Z(n4348) );
  NAND U8423 ( .A(n4395), .B(n4396), .Z(n4394) );
  NAND U8424 ( .A(n4397), .B(n4398), .Z(n4393) );
  AND U8425 ( .A(n4399), .B(n4400), .Z(n4350) );
  NAND U8426 ( .A(n4401), .B(n4402), .Z(n4344) );
  XNOR U8427 ( .A(n4327), .B(n4403), .Z(n4341) );
  XOR U8428 ( .A(n4331), .B(n4329), .Z(n4403) );
  XOR U8429 ( .A(n4337), .B(n4404), .Z(n4329) );
  XOR U8430 ( .A(n4334), .B(n4338), .Z(n4404) );
  NAND U8431 ( .A(n4405), .B(n4406), .Z(n4338) );
  NAND U8432 ( .A(n4407), .B(n4408), .Z(n4406) );
  NAND U8433 ( .A(n4409), .B(n4410), .Z(n4405) );
  AND U8434 ( .A(n4411), .B(n4412), .Z(n4334) );
  NAND U8435 ( .A(n4413), .B(n4414), .Z(n4412) );
  NAND U8436 ( .A(n4415), .B(n4416), .Z(n4411) );
  NANDN U8437 ( .A(n4417), .B(n4418), .Z(n4337) );
  NANDN U8438 ( .A(n4419), .B(n4420), .Z(n4331) );
  XNOR U8439 ( .A(n4322), .B(n4421), .Z(n4327) );
  XOR U8440 ( .A(n4320), .B(n4324), .Z(n4421) );
  NAND U8441 ( .A(n4422), .B(n4423), .Z(n4324) );
  NAND U8442 ( .A(n4424), .B(n4425), .Z(n4423) );
  NAND U8443 ( .A(n4426), .B(n4427), .Z(n4422) );
  AND U8444 ( .A(n4428), .B(n4429), .Z(n4320) );
  NAND U8445 ( .A(n4430), .B(n4431), .Z(n4429) );
  NAND U8446 ( .A(n4432), .B(n4433), .Z(n4428) );
  AND U8447 ( .A(n4434), .B(n4435), .Z(n4322) );
  XOR U8448 ( .A(n4402), .B(n4401), .Z(N29789) );
  XNOR U8449 ( .A(n4420), .B(n4419), .Z(n4401) );
  XNOR U8450 ( .A(n4434), .B(n4435), .Z(n4419) );
  XOR U8451 ( .A(n4431), .B(n4430), .Z(n4435) );
  XOR U8452 ( .A(y[3723]), .B(x[3723]), .Z(n4430) );
  XOR U8453 ( .A(n4433), .B(n4432), .Z(n4431) );
  XOR U8454 ( .A(y[3725]), .B(x[3725]), .Z(n4432) );
  XOR U8455 ( .A(y[3724]), .B(x[3724]), .Z(n4433) );
  XOR U8456 ( .A(n4425), .B(n4424), .Z(n4434) );
  XOR U8457 ( .A(n4427), .B(n4426), .Z(n4424) );
  XOR U8458 ( .A(y[3722]), .B(x[3722]), .Z(n4426) );
  XOR U8459 ( .A(y[3721]), .B(x[3721]), .Z(n4427) );
  XOR U8460 ( .A(y[3720]), .B(x[3720]), .Z(n4425) );
  XNOR U8461 ( .A(n4418), .B(n4417), .Z(n4420) );
  XNOR U8462 ( .A(n4414), .B(n4413), .Z(n4417) );
  XOR U8463 ( .A(n4416), .B(n4415), .Z(n4413) );
  XOR U8464 ( .A(y[3719]), .B(x[3719]), .Z(n4415) );
  XOR U8465 ( .A(y[3718]), .B(x[3718]), .Z(n4416) );
  XOR U8466 ( .A(y[3717]), .B(x[3717]), .Z(n4414) );
  XOR U8467 ( .A(n4408), .B(n4407), .Z(n4418) );
  XOR U8468 ( .A(n4410), .B(n4409), .Z(n4407) );
  XOR U8469 ( .A(y[3716]), .B(x[3716]), .Z(n4409) );
  XOR U8470 ( .A(y[3715]), .B(x[3715]), .Z(n4410) );
  XOR U8471 ( .A(y[3714]), .B(x[3714]), .Z(n4408) );
  XNOR U8472 ( .A(n4385), .B(n4384), .Z(n4402) );
  XNOR U8473 ( .A(n4399), .B(n4400), .Z(n4384) );
  XOR U8474 ( .A(n4396), .B(n4395), .Z(n4400) );
  XOR U8475 ( .A(y[3711]), .B(x[3711]), .Z(n4395) );
  XOR U8476 ( .A(n4398), .B(n4397), .Z(n4396) );
  XOR U8477 ( .A(y[3713]), .B(x[3713]), .Z(n4397) );
  XOR U8478 ( .A(y[3712]), .B(x[3712]), .Z(n4398) );
  XOR U8479 ( .A(n4390), .B(n4389), .Z(n4399) );
  XOR U8480 ( .A(n4392), .B(n4391), .Z(n4389) );
  XOR U8481 ( .A(y[3710]), .B(x[3710]), .Z(n4391) );
  XOR U8482 ( .A(y[3709]), .B(x[3709]), .Z(n4392) );
  XOR U8483 ( .A(y[3708]), .B(x[3708]), .Z(n4390) );
  XNOR U8484 ( .A(n4383), .B(n4382), .Z(n4385) );
  XNOR U8485 ( .A(n4379), .B(n4378), .Z(n4382) );
  XOR U8486 ( .A(n4381), .B(n4380), .Z(n4378) );
  XOR U8487 ( .A(y[3707]), .B(x[3707]), .Z(n4380) );
  XOR U8488 ( .A(y[3706]), .B(x[3706]), .Z(n4381) );
  XOR U8489 ( .A(y[3705]), .B(x[3705]), .Z(n4379) );
  XOR U8490 ( .A(n4373), .B(n4372), .Z(n4383) );
  XOR U8491 ( .A(n4375), .B(n4374), .Z(n4372) );
  XOR U8492 ( .A(y[3704]), .B(x[3704]), .Z(n4374) );
  XOR U8493 ( .A(y[3703]), .B(x[3703]), .Z(n4375) );
  XOR U8494 ( .A(y[3702]), .B(x[3702]), .Z(n4373) );
  NAND U8495 ( .A(n4436), .B(n4437), .Z(N29781) );
  NAND U8496 ( .A(n4438), .B(n4439), .Z(n4437) );
  NANDN U8497 ( .A(n4440), .B(n4441), .Z(n4439) );
  NANDN U8498 ( .A(n4441), .B(n4440), .Z(n4436) );
  XOR U8499 ( .A(n4440), .B(n4442), .Z(N29780) );
  XNOR U8500 ( .A(n4438), .B(n4441), .Z(n4442) );
  NAND U8501 ( .A(n4443), .B(n4444), .Z(n4441) );
  NAND U8502 ( .A(n4445), .B(n4446), .Z(n4444) );
  NANDN U8503 ( .A(n4447), .B(n4448), .Z(n4446) );
  NANDN U8504 ( .A(n4448), .B(n4447), .Z(n4443) );
  AND U8505 ( .A(n4449), .B(n4450), .Z(n4438) );
  NAND U8506 ( .A(n4451), .B(n4452), .Z(n4450) );
  OR U8507 ( .A(n4453), .B(n4454), .Z(n4452) );
  NAND U8508 ( .A(n4454), .B(n4453), .Z(n4449) );
  IV U8509 ( .A(n4455), .Z(n4454) );
  AND U8510 ( .A(n4456), .B(n4457), .Z(n4440) );
  NAND U8511 ( .A(n4458), .B(n4459), .Z(n4457) );
  NANDN U8512 ( .A(n4460), .B(n4461), .Z(n4459) );
  NANDN U8513 ( .A(n4461), .B(n4460), .Z(n4456) );
  XOR U8514 ( .A(n4453), .B(n4462), .Z(N29779) );
  XOR U8515 ( .A(n4451), .B(n4455), .Z(n4462) );
  XNOR U8516 ( .A(n4448), .B(n4463), .Z(n4455) );
  XNOR U8517 ( .A(n4445), .B(n4447), .Z(n4463) );
  AND U8518 ( .A(n4464), .B(n4465), .Z(n4447) );
  NANDN U8519 ( .A(n4466), .B(n4467), .Z(n4465) );
  NANDN U8520 ( .A(n4468), .B(n4469), .Z(n4467) );
  IV U8521 ( .A(n4470), .Z(n4469) );
  NAND U8522 ( .A(n4470), .B(n4468), .Z(n4464) );
  AND U8523 ( .A(n4471), .B(n4472), .Z(n4445) );
  NAND U8524 ( .A(n4473), .B(n4474), .Z(n4472) );
  OR U8525 ( .A(n4475), .B(n4476), .Z(n4474) );
  NAND U8526 ( .A(n4476), .B(n4475), .Z(n4471) );
  IV U8527 ( .A(n4477), .Z(n4476) );
  NAND U8528 ( .A(n4478), .B(n4479), .Z(n4448) );
  NANDN U8529 ( .A(n4480), .B(n4481), .Z(n4479) );
  NAND U8530 ( .A(n4482), .B(n4483), .Z(n4481) );
  OR U8531 ( .A(n4483), .B(n4482), .Z(n4478) );
  IV U8532 ( .A(n4484), .Z(n4482) );
  AND U8533 ( .A(n4485), .B(n4486), .Z(n4451) );
  NAND U8534 ( .A(n4487), .B(n4488), .Z(n4486) );
  NANDN U8535 ( .A(n4489), .B(n4490), .Z(n4488) );
  NANDN U8536 ( .A(n4490), .B(n4489), .Z(n4485) );
  XOR U8537 ( .A(n4461), .B(n4491), .Z(n4453) );
  XNOR U8538 ( .A(n4458), .B(n4460), .Z(n4491) );
  AND U8539 ( .A(n4492), .B(n4493), .Z(n4460) );
  NANDN U8540 ( .A(n4494), .B(n4495), .Z(n4493) );
  NANDN U8541 ( .A(n4496), .B(n4497), .Z(n4495) );
  IV U8542 ( .A(n4498), .Z(n4497) );
  NAND U8543 ( .A(n4498), .B(n4496), .Z(n4492) );
  AND U8544 ( .A(n4499), .B(n4500), .Z(n4458) );
  NAND U8545 ( .A(n4501), .B(n4502), .Z(n4500) );
  OR U8546 ( .A(n4503), .B(n4504), .Z(n4502) );
  NAND U8547 ( .A(n4504), .B(n4503), .Z(n4499) );
  IV U8548 ( .A(n4505), .Z(n4504) );
  NAND U8549 ( .A(n4506), .B(n4507), .Z(n4461) );
  NANDN U8550 ( .A(n4508), .B(n4509), .Z(n4507) );
  NAND U8551 ( .A(n4510), .B(n4511), .Z(n4509) );
  OR U8552 ( .A(n4511), .B(n4510), .Z(n4506) );
  IV U8553 ( .A(n4512), .Z(n4510) );
  XOR U8554 ( .A(n4487), .B(n4513), .Z(N29778) );
  XNOR U8555 ( .A(n4490), .B(n4489), .Z(n4513) );
  XNOR U8556 ( .A(n4501), .B(n4514), .Z(n4489) );
  XOR U8557 ( .A(n4505), .B(n4503), .Z(n4514) );
  XOR U8558 ( .A(n4511), .B(n4515), .Z(n4503) );
  XOR U8559 ( .A(n4508), .B(n4512), .Z(n4515) );
  NAND U8560 ( .A(n4516), .B(n4517), .Z(n4512) );
  NAND U8561 ( .A(n4518), .B(n4519), .Z(n4517) );
  NAND U8562 ( .A(n4520), .B(n4521), .Z(n4516) );
  AND U8563 ( .A(n4522), .B(n4523), .Z(n4508) );
  NAND U8564 ( .A(n4524), .B(n4525), .Z(n4523) );
  NAND U8565 ( .A(n4526), .B(n4527), .Z(n4522) );
  NANDN U8566 ( .A(n4528), .B(n4529), .Z(n4511) );
  NANDN U8567 ( .A(n4530), .B(n4531), .Z(n4505) );
  XNOR U8568 ( .A(n4496), .B(n4532), .Z(n4501) );
  XOR U8569 ( .A(n4494), .B(n4498), .Z(n4532) );
  NAND U8570 ( .A(n4533), .B(n4534), .Z(n4498) );
  NAND U8571 ( .A(n4535), .B(n4536), .Z(n4534) );
  NAND U8572 ( .A(n4537), .B(n4538), .Z(n4533) );
  AND U8573 ( .A(n4539), .B(n4540), .Z(n4494) );
  NAND U8574 ( .A(n4541), .B(n4542), .Z(n4540) );
  NAND U8575 ( .A(n4543), .B(n4544), .Z(n4539) );
  AND U8576 ( .A(n4545), .B(n4546), .Z(n4496) );
  NAND U8577 ( .A(n4547), .B(n4548), .Z(n4490) );
  XNOR U8578 ( .A(n4473), .B(n4549), .Z(n4487) );
  XOR U8579 ( .A(n4477), .B(n4475), .Z(n4549) );
  XOR U8580 ( .A(n4483), .B(n4550), .Z(n4475) );
  XOR U8581 ( .A(n4480), .B(n4484), .Z(n4550) );
  NAND U8582 ( .A(n4551), .B(n4552), .Z(n4484) );
  NAND U8583 ( .A(n4553), .B(n4554), .Z(n4552) );
  NAND U8584 ( .A(n4555), .B(n4556), .Z(n4551) );
  AND U8585 ( .A(n4557), .B(n4558), .Z(n4480) );
  NAND U8586 ( .A(n4559), .B(n4560), .Z(n4558) );
  NAND U8587 ( .A(n4561), .B(n4562), .Z(n4557) );
  NANDN U8588 ( .A(n4563), .B(n4564), .Z(n4483) );
  NANDN U8589 ( .A(n4565), .B(n4566), .Z(n4477) );
  XNOR U8590 ( .A(n4468), .B(n4567), .Z(n4473) );
  XOR U8591 ( .A(n4466), .B(n4470), .Z(n4567) );
  NAND U8592 ( .A(n4568), .B(n4569), .Z(n4470) );
  NAND U8593 ( .A(n4570), .B(n4571), .Z(n4569) );
  NAND U8594 ( .A(n4572), .B(n4573), .Z(n4568) );
  AND U8595 ( .A(n4574), .B(n4575), .Z(n4466) );
  NAND U8596 ( .A(n4576), .B(n4577), .Z(n4575) );
  NAND U8597 ( .A(n4578), .B(n4579), .Z(n4574) );
  AND U8598 ( .A(n4580), .B(n4581), .Z(n4468) );
  XOR U8599 ( .A(n4548), .B(n4547), .Z(N29777) );
  XNOR U8600 ( .A(n4566), .B(n4565), .Z(n4547) );
  XNOR U8601 ( .A(n4580), .B(n4581), .Z(n4565) );
  XOR U8602 ( .A(n4577), .B(n4576), .Z(n4581) );
  XOR U8603 ( .A(y[3699]), .B(x[3699]), .Z(n4576) );
  XOR U8604 ( .A(n4579), .B(n4578), .Z(n4577) );
  XOR U8605 ( .A(y[3701]), .B(x[3701]), .Z(n4578) );
  XOR U8606 ( .A(y[3700]), .B(x[3700]), .Z(n4579) );
  XOR U8607 ( .A(n4571), .B(n4570), .Z(n4580) );
  XOR U8608 ( .A(n4573), .B(n4572), .Z(n4570) );
  XOR U8609 ( .A(y[3698]), .B(x[3698]), .Z(n4572) );
  XOR U8610 ( .A(y[3697]), .B(x[3697]), .Z(n4573) );
  XOR U8611 ( .A(y[3696]), .B(x[3696]), .Z(n4571) );
  XNOR U8612 ( .A(n4564), .B(n4563), .Z(n4566) );
  XNOR U8613 ( .A(n4560), .B(n4559), .Z(n4563) );
  XOR U8614 ( .A(n4562), .B(n4561), .Z(n4559) );
  XOR U8615 ( .A(y[3695]), .B(x[3695]), .Z(n4561) );
  XOR U8616 ( .A(y[3694]), .B(x[3694]), .Z(n4562) );
  XOR U8617 ( .A(y[3693]), .B(x[3693]), .Z(n4560) );
  XOR U8618 ( .A(n4554), .B(n4553), .Z(n4564) );
  XOR U8619 ( .A(n4556), .B(n4555), .Z(n4553) );
  XOR U8620 ( .A(y[3692]), .B(x[3692]), .Z(n4555) );
  XOR U8621 ( .A(y[3691]), .B(x[3691]), .Z(n4556) );
  XOR U8622 ( .A(y[3690]), .B(x[3690]), .Z(n4554) );
  XNOR U8623 ( .A(n4531), .B(n4530), .Z(n4548) );
  XNOR U8624 ( .A(n4545), .B(n4546), .Z(n4530) );
  XOR U8625 ( .A(n4542), .B(n4541), .Z(n4546) );
  XOR U8626 ( .A(y[3687]), .B(x[3687]), .Z(n4541) );
  XOR U8627 ( .A(n4544), .B(n4543), .Z(n4542) );
  XOR U8628 ( .A(y[3689]), .B(x[3689]), .Z(n4543) );
  XOR U8629 ( .A(y[3688]), .B(x[3688]), .Z(n4544) );
  XOR U8630 ( .A(n4536), .B(n4535), .Z(n4545) );
  XOR U8631 ( .A(n4538), .B(n4537), .Z(n4535) );
  XOR U8632 ( .A(y[3686]), .B(x[3686]), .Z(n4537) );
  XOR U8633 ( .A(y[3685]), .B(x[3685]), .Z(n4538) );
  XOR U8634 ( .A(y[3684]), .B(x[3684]), .Z(n4536) );
  XNOR U8635 ( .A(n4529), .B(n4528), .Z(n4531) );
  XNOR U8636 ( .A(n4525), .B(n4524), .Z(n4528) );
  XOR U8637 ( .A(n4527), .B(n4526), .Z(n4524) );
  XOR U8638 ( .A(y[3683]), .B(x[3683]), .Z(n4526) );
  XOR U8639 ( .A(y[3682]), .B(x[3682]), .Z(n4527) );
  XOR U8640 ( .A(y[3681]), .B(x[3681]), .Z(n4525) );
  XOR U8641 ( .A(n4519), .B(n4518), .Z(n4529) );
  XOR U8642 ( .A(n4521), .B(n4520), .Z(n4518) );
  XOR U8643 ( .A(y[3680]), .B(x[3680]), .Z(n4520) );
  XOR U8644 ( .A(y[3679]), .B(x[3679]), .Z(n4521) );
  XOR U8645 ( .A(y[3678]), .B(x[3678]), .Z(n4519) );
  NAND U8646 ( .A(n4582), .B(n4583), .Z(N29769) );
  NAND U8647 ( .A(n4584), .B(n4585), .Z(n4583) );
  NANDN U8648 ( .A(n4586), .B(n4587), .Z(n4585) );
  NANDN U8649 ( .A(n4587), .B(n4586), .Z(n4582) );
  XOR U8650 ( .A(n4586), .B(n4588), .Z(N29768) );
  XNOR U8651 ( .A(n4584), .B(n4587), .Z(n4588) );
  NAND U8652 ( .A(n4589), .B(n4590), .Z(n4587) );
  NAND U8653 ( .A(n4591), .B(n4592), .Z(n4590) );
  NANDN U8654 ( .A(n4593), .B(n4594), .Z(n4592) );
  NANDN U8655 ( .A(n4594), .B(n4593), .Z(n4589) );
  AND U8656 ( .A(n4595), .B(n4596), .Z(n4584) );
  NAND U8657 ( .A(n4597), .B(n4598), .Z(n4596) );
  OR U8658 ( .A(n4599), .B(n4600), .Z(n4598) );
  NAND U8659 ( .A(n4600), .B(n4599), .Z(n4595) );
  IV U8660 ( .A(n4601), .Z(n4600) );
  AND U8661 ( .A(n4602), .B(n4603), .Z(n4586) );
  NAND U8662 ( .A(n4604), .B(n4605), .Z(n4603) );
  NANDN U8663 ( .A(n4606), .B(n4607), .Z(n4605) );
  NANDN U8664 ( .A(n4607), .B(n4606), .Z(n4602) );
  XOR U8665 ( .A(n4599), .B(n4608), .Z(N29767) );
  XOR U8666 ( .A(n4597), .B(n4601), .Z(n4608) );
  XNOR U8667 ( .A(n4594), .B(n4609), .Z(n4601) );
  XNOR U8668 ( .A(n4591), .B(n4593), .Z(n4609) );
  AND U8669 ( .A(n4610), .B(n4611), .Z(n4593) );
  NANDN U8670 ( .A(n4612), .B(n4613), .Z(n4611) );
  NANDN U8671 ( .A(n4614), .B(n4615), .Z(n4613) );
  IV U8672 ( .A(n4616), .Z(n4615) );
  NAND U8673 ( .A(n4616), .B(n4614), .Z(n4610) );
  AND U8674 ( .A(n4617), .B(n4618), .Z(n4591) );
  NAND U8675 ( .A(n4619), .B(n4620), .Z(n4618) );
  OR U8676 ( .A(n4621), .B(n4622), .Z(n4620) );
  NAND U8677 ( .A(n4622), .B(n4621), .Z(n4617) );
  IV U8678 ( .A(n4623), .Z(n4622) );
  NAND U8679 ( .A(n4624), .B(n4625), .Z(n4594) );
  NANDN U8680 ( .A(n4626), .B(n4627), .Z(n4625) );
  NAND U8681 ( .A(n4628), .B(n4629), .Z(n4627) );
  OR U8682 ( .A(n4629), .B(n4628), .Z(n4624) );
  IV U8683 ( .A(n4630), .Z(n4628) );
  AND U8684 ( .A(n4631), .B(n4632), .Z(n4597) );
  NAND U8685 ( .A(n4633), .B(n4634), .Z(n4632) );
  NANDN U8686 ( .A(n4635), .B(n4636), .Z(n4634) );
  NANDN U8687 ( .A(n4636), .B(n4635), .Z(n4631) );
  XOR U8688 ( .A(n4607), .B(n4637), .Z(n4599) );
  XNOR U8689 ( .A(n4604), .B(n4606), .Z(n4637) );
  AND U8690 ( .A(n4638), .B(n4639), .Z(n4606) );
  NANDN U8691 ( .A(n4640), .B(n4641), .Z(n4639) );
  NANDN U8692 ( .A(n4642), .B(n4643), .Z(n4641) );
  IV U8693 ( .A(n4644), .Z(n4643) );
  NAND U8694 ( .A(n4644), .B(n4642), .Z(n4638) );
  AND U8695 ( .A(n4645), .B(n4646), .Z(n4604) );
  NAND U8696 ( .A(n4647), .B(n4648), .Z(n4646) );
  OR U8697 ( .A(n4649), .B(n4650), .Z(n4648) );
  NAND U8698 ( .A(n4650), .B(n4649), .Z(n4645) );
  IV U8699 ( .A(n4651), .Z(n4650) );
  NAND U8700 ( .A(n4652), .B(n4653), .Z(n4607) );
  NANDN U8701 ( .A(n4654), .B(n4655), .Z(n4653) );
  NAND U8702 ( .A(n4656), .B(n4657), .Z(n4655) );
  OR U8703 ( .A(n4657), .B(n4656), .Z(n4652) );
  IV U8704 ( .A(n4658), .Z(n4656) );
  XOR U8705 ( .A(n4633), .B(n4659), .Z(N29766) );
  XNOR U8706 ( .A(n4636), .B(n4635), .Z(n4659) );
  XNOR U8707 ( .A(n4647), .B(n4660), .Z(n4635) );
  XOR U8708 ( .A(n4651), .B(n4649), .Z(n4660) );
  XOR U8709 ( .A(n4657), .B(n4661), .Z(n4649) );
  XOR U8710 ( .A(n4654), .B(n4658), .Z(n4661) );
  NAND U8711 ( .A(n4662), .B(n4663), .Z(n4658) );
  NAND U8712 ( .A(n4664), .B(n4665), .Z(n4663) );
  NAND U8713 ( .A(n4666), .B(n4667), .Z(n4662) );
  AND U8714 ( .A(n4668), .B(n4669), .Z(n4654) );
  NAND U8715 ( .A(n4670), .B(n4671), .Z(n4669) );
  NAND U8716 ( .A(n4672), .B(n4673), .Z(n4668) );
  NANDN U8717 ( .A(n4674), .B(n4675), .Z(n4657) );
  NANDN U8718 ( .A(n4676), .B(n4677), .Z(n4651) );
  XNOR U8719 ( .A(n4642), .B(n4678), .Z(n4647) );
  XOR U8720 ( .A(n4640), .B(n4644), .Z(n4678) );
  NAND U8721 ( .A(n4679), .B(n4680), .Z(n4644) );
  NAND U8722 ( .A(n4681), .B(n4682), .Z(n4680) );
  NAND U8723 ( .A(n4683), .B(n4684), .Z(n4679) );
  AND U8724 ( .A(n4685), .B(n4686), .Z(n4640) );
  NAND U8725 ( .A(n4687), .B(n4688), .Z(n4686) );
  NAND U8726 ( .A(n4689), .B(n4690), .Z(n4685) );
  AND U8727 ( .A(n4691), .B(n4692), .Z(n4642) );
  NAND U8728 ( .A(n4693), .B(n4694), .Z(n4636) );
  XNOR U8729 ( .A(n4619), .B(n4695), .Z(n4633) );
  XOR U8730 ( .A(n4623), .B(n4621), .Z(n4695) );
  XOR U8731 ( .A(n4629), .B(n4696), .Z(n4621) );
  XOR U8732 ( .A(n4626), .B(n4630), .Z(n4696) );
  NAND U8733 ( .A(n4697), .B(n4698), .Z(n4630) );
  NAND U8734 ( .A(n4699), .B(n4700), .Z(n4698) );
  NAND U8735 ( .A(n4701), .B(n4702), .Z(n4697) );
  AND U8736 ( .A(n4703), .B(n4704), .Z(n4626) );
  NAND U8737 ( .A(n4705), .B(n4706), .Z(n4704) );
  NAND U8738 ( .A(n4707), .B(n4708), .Z(n4703) );
  NANDN U8739 ( .A(n4709), .B(n4710), .Z(n4629) );
  NANDN U8740 ( .A(n4711), .B(n4712), .Z(n4623) );
  XNOR U8741 ( .A(n4614), .B(n4713), .Z(n4619) );
  XOR U8742 ( .A(n4612), .B(n4616), .Z(n4713) );
  NAND U8743 ( .A(n4714), .B(n4715), .Z(n4616) );
  NAND U8744 ( .A(n4716), .B(n4717), .Z(n4715) );
  NAND U8745 ( .A(n4718), .B(n4719), .Z(n4714) );
  AND U8746 ( .A(n4720), .B(n4721), .Z(n4612) );
  NAND U8747 ( .A(n4722), .B(n4723), .Z(n4721) );
  NAND U8748 ( .A(n4724), .B(n4725), .Z(n4720) );
  AND U8749 ( .A(n4726), .B(n4727), .Z(n4614) );
  XOR U8750 ( .A(n4694), .B(n4693), .Z(N29765) );
  XNOR U8751 ( .A(n4712), .B(n4711), .Z(n4693) );
  XNOR U8752 ( .A(n4726), .B(n4727), .Z(n4711) );
  XOR U8753 ( .A(n4723), .B(n4722), .Z(n4727) );
  XOR U8754 ( .A(y[3675]), .B(x[3675]), .Z(n4722) );
  XOR U8755 ( .A(n4725), .B(n4724), .Z(n4723) );
  XOR U8756 ( .A(y[3677]), .B(x[3677]), .Z(n4724) );
  XOR U8757 ( .A(y[3676]), .B(x[3676]), .Z(n4725) );
  XOR U8758 ( .A(n4717), .B(n4716), .Z(n4726) );
  XOR U8759 ( .A(n4719), .B(n4718), .Z(n4716) );
  XOR U8760 ( .A(y[3674]), .B(x[3674]), .Z(n4718) );
  XOR U8761 ( .A(y[3673]), .B(x[3673]), .Z(n4719) );
  XOR U8762 ( .A(y[3672]), .B(x[3672]), .Z(n4717) );
  XNOR U8763 ( .A(n4710), .B(n4709), .Z(n4712) );
  XNOR U8764 ( .A(n4706), .B(n4705), .Z(n4709) );
  XOR U8765 ( .A(n4708), .B(n4707), .Z(n4705) );
  XOR U8766 ( .A(y[3671]), .B(x[3671]), .Z(n4707) );
  XOR U8767 ( .A(y[3670]), .B(x[3670]), .Z(n4708) );
  XOR U8768 ( .A(y[3669]), .B(x[3669]), .Z(n4706) );
  XOR U8769 ( .A(n4700), .B(n4699), .Z(n4710) );
  XOR U8770 ( .A(n4702), .B(n4701), .Z(n4699) );
  XOR U8771 ( .A(y[3668]), .B(x[3668]), .Z(n4701) );
  XOR U8772 ( .A(y[3667]), .B(x[3667]), .Z(n4702) );
  XOR U8773 ( .A(y[3666]), .B(x[3666]), .Z(n4700) );
  XNOR U8774 ( .A(n4677), .B(n4676), .Z(n4694) );
  XNOR U8775 ( .A(n4691), .B(n4692), .Z(n4676) );
  XOR U8776 ( .A(n4688), .B(n4687), .Z(n4692) );
  XOR U8777 ( .A(y[3663]), .B(x[3663]), .Z(n4687) );
  XOR U8778 ( .A(n4690), .B(n4689), .Z(n4688) );
  XOR U8779 ( .A(y[3665]), .B(x[3665]), .Z(n4689) );
  XOR U8780 ( .A(y[3664]), .B(x[3664]), .Z(n4690) );
  XOR U8781 ( .A(n4682), .B(n4681), .Z(n4691) );
  XOR U8782 ( .A(n4684), .B(n4683), .Z(n4681) );
  XOR U8783 ( .A(y[3662]), .B(x[3662]), .Z(n4683) );
  XOR U8784 ( .A(y[3661]), .B(x[3661]), .Z(n4684) );
  XOR U8785 ( .A(y[3660]), .B(x[3660]), .Z(n4682) );
  XNOR U8786 ( .A(n4675), .B(n4674), .Z(n4677) );
  XNOR U8787 ( .A(n4671), .B(n4670), .Z(n4674) );
  XOR U8788 ( .A(n4673), .B(n4672), .Z(n4670) );
  XOR U8789 ( .A(y[3659]), .B(x[3659]), .Z(n4672) );
  XOR U8790 ( .A(y[3658]), .B(x[3658]), .Z(n4673) );
  XOR U8791 ( .A(y[3657]), .B(x[3657]), .Z(n4671) );
  XOR U8792 ( .A(n4665), .B(n4664), .Z(n4675) );
  XOR U8793 ( .A(n4667), .B(n4666), .Z(n4664) );
  XOR U8794 ( .A(y[3656]), .B(x[3656]), .Z(n4666) );
  XOR U8795 ( .A(y[3655]), .B(x[3655]), .Z(n4667) );
  XOR U8796 ( .A(y[3654]), .B(x[3654]), .Z(n4665) );
  NAND U8797 ( .A(n4728), .B(n4729), .Z(N29757) );
  NAND U8798 ( .A(n4730), .B(n4731), .Z(n4729) );
  NANDN U8799 ( .A(n4732), .B(n4733), .Z(n4731) );
  NANDN U8800 ( .A(n4733), .B(n4732), .Z(n4728) );
  XOR U8801 ( .A(n4732), .B(n4734), .Z(N29756) );
  XNOR U8802 ( .A(n4730), .B(n4733), .Z(n4734) );
  NAND U8803 ( .A(n4735), .B(n4736), .Z(n4733) );
  NAND U8804 ( .A(n4737), .B(n4738), .Z(n4736) );
  NANDN U8805 ( .A(n4739), .B(n4740), .Z(n4738) );
  NANDN U8806 ( .A(n4740), .B(n4739), .Z(n4735) );
  AND U8807 ( .A(n4741), .B(n4742), .Z(n4730) );
  NAND U8808 ( .A(n4743), .B(n4744), .Z(n4742) );
  OR U8809 ( .A(n4745), .B(n4746), .Z(n4744) );
  NAND U8810 ( .A(n4746), .B(n4745), .Z(n4741) );
  IV U8811 ( .A(n4747), .Z(n4746) );
  AND U8812 ( .A(n4748), .B(n4749), .Z(n4732) );
  NAND U8813 ( .A(n4750), .B(n4751), .Z(n4749) );
  NANDN U8814 ( .A(n4752), .B(n4753), .Z(n4751) );
  NANDN U8815 ( .A(n4753), .B(n4752), .Z(n4748) );
  XOR U8816 ( .A(n4745), .B(n4754), .Z(N29755) );
  XOR U8817 ( .A(n4743), .B(n4747), .Z(n4754) );
  XNOR U8818 ( .A(n4740), .B(n4755), .Z(n4747) );
  XNOR U8819 ( .A(n4737), .B(n4739), .Z(n4755) );
  AND U8820 ( .A(n4756), .B(n4757), .Z(n4739) );
  NANDN U8821 ( .A(n4758), .B(n4759), .Z(n4757) );
  NANDN U8822 ( .A(n4760), .B(n4761), .Z(n4759) );
  IV U8823 ( .A(n4762), .Z(n4761) );
  NAND U8824 ( .A(n4762), .B(n4760), .Z(n4756) );
  AND U8825 ( .A(n4763), .B(n4764), .Z(n4737) );
  NAND U8826 ( .A(n4765), .B(n4766), .Z(n4764) );
  OR U8827 ( .A(n4767), .B(n4768), .Z(n4766) );
  NAND U8828 ( .A(n4768), .B(n4767), .Z(n4763) );
  IV U8829 ( .A(n4769), .Z(n4768) );
  NAND U8830 ( .A(n4770), .B(n4771), .Z(n4740) );
  NANDN U8831 ( .A(n4772), .B(n4773), .Z(n4771) );
  NAND U8832 ( .A(n4774), .B(n4775), .Z(n4773) );
  OR U8833 ( .A(n4775), .B(n4774), .Z(n4770) );
  IV U8834 ( .A(n4776), .Z(n4774) );
  AND U8835 ( .A(n4777), .B(n4778), .Z(n4743) );
  NAND U8836 ( .A(n4779), .B(n4780), .Z(n4778) );
  NANDN U8837 ( .A(n4781), .B(n4782), .Z(n4780) );
  NANDN U8838 ( .A(n4782), .B(n4781), .Z(n4777) );
  XOR U8839 ( .A(n4753), .B(n4783), .Z(n4745) );
  XNOR U8840 ( .A(n4750), .B(n4752), .Z(n4783) );
  AND U8841 ( .A(n4784), .B(n4785), .Z(n4752) );
  NANDN U8842 ( .A(n4786), .B(n4787), .Z(n4785) );
  NANDN U8843 ( .A(n4788), .B(n4789), .Z(n4787) );
  IV U8844 ( .A(n4790), .Z(n4789) );
  NAND U8845 ( .A(n4790), .B(n4788), .Z(n4784) );
  AND U8846 ( .A(n4791), .B(n4792), .Z(n4750) );
  NAND U8847 ( .A(n4793), .B(n4794), .Z(n4792) );
  OR U8848 ( .A(n4795), .B(n4796), .Z(n4794) );
  NAND U8849 ( .A(n4796), .B(n4795), .Z(n4791) );
  IV U8850 ( .A(n4797), .Z(n4796) );
  NAND U8851 ( .A(n4798), .B(n4799), .Z(n4753) );
  NANDN U8852 ( .A(n4800), .B(n4801), .Z(n4799) );
  NAND U8853 ( .A(n4802), .B(n4803), .Z(n4801) );
  OR U8854 ( .A(n4803), .B(n4802), .Z(n4798) );
  IV U8855 ( .A(n4804), .Z(n4802) );
  XOR U8856 ( .A(n4779), .B(n4805), .Z(N29754) );
  XNOR U8857 ( .A(n4782), .B(n4781), .Z(n4805) );
  XNOR U8858 ( .A(n4793), .B(n4806), .Z(n4781) );
  XOR U8859 ( .A(n4797), .B(n4795), .Z(n4806) );
  XOR U8860 ( .A(n4803), .B(n4807), .Z(n4795) );
  XOR U8861 ( .A(n4800), .B(n4804), .Z(n4807) );
  NAND U8862 ( .A(n4808), .B(n4809), .Z(n4804) );
  NAND U8863 ( .A(n4810), .B(n4811), .Z(n4809) );
  NAND U8864 ( .A(n4812), .B(n4813), .Z(n4808) );
  AND U8865 ( .A(n4814), .B(n4815), .Z(n4800) );
  NAND U8866 ( .A(n4816), .B(n4817), .Z(n4815) );
  NAND U8867 ( .A(n4818), .B(n4819), .Z(n4814) );
  NANDN U8868 ( .A(n4820), .B(n4821), .Z(n4803) );
  NANDN U8869 ( .A(n4822), .B(n4823), .Z(n4797) );
  XNOR U8870 ( .A(n4788), .B(n4824), .Z(n4793) );
  XOR U8871 ( .A(n4786), .B(n4790), .Z(n4824) );
  NAND U8872 ( .A(n4825), .B(n4826), .Z(n4790) );
  NAND U8873 ( .A(n4827), .B(n4828), .Z(n4826) );
  NAND U8874 ( .A(n4829), .B(n4830), .Z(n4825) );
  AND U8875 ( .A(n4831), .B(n4832), .Z(n4786) );
  NAND U8876 ( .A(n4833), .B(n4834), .Z(n4832) );
  NAND U8877 ( .A(n4835), .B(n4836), .Z(n4831) );
  AND U8878 ( .A(n4837), .B(n4838), .Z(n4788) );
  NAND U8879 ( .A(n4839), .B(n4840), .Z(n4782) );
  XNOR U8880 ( .A(n4765), .B(n4841), .Z(n4779) );
  XOR U8881 ( .A(n4769), .B(n4767), .Z(n4841) );
  XOR U8882 ( .A(n4775), .B(n4842), .Z(n4767) );
  XOR U8883 ( .A(n4772), .B(n4776), .Z(n4842) );
  NAND U8884 ( .A(n4843), .B(n4844), .Z(n4776) );
  NAND U8885 ( .A(n4845), .B(n4846), .Z(n4844) );
  NAND U8886 ( .A(n4847), .B(n4848), .Z(n4843) );
  AND U8887 ( .A(n4849), .B(n4850), .Z(n4772) );
  NAND U8888 ( .A(n4851), .B(n4852), .Z(n4850) );
  NAND U8889 ( .A(n4853), .B(n4854), .Z(n4849) );
  NANDN U8890 ( .A(n4855), .B(n4856), .Z(n4775) );
  NANDN U8891 ( .A(n4857), .B(n4858), .Z(n4769) );
  XNOR U8892 ( .A(n4760), .B(n4859), .Z(n4765) );
  XOR U8893 ( .A(n4758), .B(n4762), .Z(n4859) );
  NAND U8894 ( .A(n4860), .B(n4861), .Z(n4762) );
  NAND U8895 ( .A(n4862), .B(n4863), .Z(n4861) );
  NAND U8896 ( .A(n4864), .B(n4865), .Z(n4860) );
  AND U8897 ( .A(n4866), .B(n4867), .Z(n4758) );
  NAND U8898 ( .A(n4868), .B(n4869), .Z(n4867) );
  NAND U8899 ( .A(n4870), .B(n4871), .Z(n4866) );
  AND U8900 ( .A(n4872), .B(n4873), .Z(n4760) );
  XOR U8901 ( .A(n4840), .B(n4839), .Z(N29753) );
  XNOR U8902 ( .A(n4858), .B(n4857), .Z(n4839) );
  XNOR U8903 ( .A(n4872), .B(n4873), .Z(n4857) );
  XOR U8904 ( .A(n4869), .B(n4868), .Z(n4873) );
  XOR U8905 ( .A(y[3651]), .B(x[3651]), .Z(n4868) );
  XOR U8906 ( .A(n4871), .B(n4870), .Z(n4869) );
  XOR U8907 ( .A(y[3653]), .B(x[3653]), .Z(n4870) );
  XOR U8908 ( .A(y[3652]), .B(x[3652]), .Z(n4871) );
  XOR U8909 ( .A(n4863), .B(n4862), .Z(n4872) );
  XOR U8910 ( .A(n4865), .B(n4864), .Z(n4862) );
  XOR U8911 ( .A(y[3650]), .B(x[3650]), .Z(n4864) );
  XOR U8912 ( .A(y[3649]), .B(x[3649]), .Z(n4865) );
  XOR U8913 ( .A(y[3648]), .B(x[3648]), .Z(n4863) );
  XNOR U8914 ( .A(n4856), .B(n4855), .Z(n4858) );
  XNOR U8915 ( .A(n4852), .B(n4851), .Z(n4855) );
  XOR U8916 ( .A(n4854), .B(n4853), .Z(n4851) );
  XOR U8917 ( .A(y[3647]), .B(x[3647]), .Z(n4853) );
  XOR U8918 ( .A(y[3646]), .B(x[3646]), .Z(n4854) );
  XOR U8919 ( .A(y[3645]), .B(x[3645]), .Z(n4852) );
  XOR U8920 ( .A(n4846), .B(n4845), .Z(n4856) );
  XOR U8921 ( .A(n4848), .B(n4847), .Z(n4845) );
  XOR U8922 ( .A(y[3644]), .B(x[3644]), .Z(n4847) );
  XOR U8923 ( .A(y[3643]), .B(x[3643]), .Z(n4848) );
  XOR U8924 ( .A(y[3642]), .B(x[3642]), .Z(n4846) );
  XNOR U8925 ( .A(n4823), .B(n4822), .Z(n4840) );
  XNOR U8926 ( .A(n4837), .B(n4838), .Z(n4822) );
  XOR U8927 ( .A(n4834), .B(n4833), .Z(n4838) );
  XOR U8928 ( .A(y[3639]), .B(x[3639]), .Z(n4833) );
  XOR U8929 ( .A(n4836), .B(n4835), .Z(n4834) );
  XOR U8930 ( .A(y[3641]), .B(x[3641]), .Z(n4835) );
  XOR U8931 ( .A(y[3640]), .B(x[3640]), .Z(n4836) );
  XOR U8932 ( .A(n4828), .B(n4827), .Z(n4837) );
  XOR U8933 ( .A(n4830), .B(n4829), .Z(n4827) );
  XOR U8934 ( .A(y[3638]), .B(x[3638]), .Z(n4829) );
  XOR U8935 ( .A(y[3637]), .B(x[3637]), .Z(n4830) );
  XOR U8936 ( .A(y[3636]), .B(x[3636]), .Z(n4828) );
  XNOR U8937 ( .A(n4821), .B(n4820), .Z(n4823) );
  XNOR U8938 ( .A(n4817), .B(n4816), .Z(n4820) );
  XOR U8939 ( .A(n4819), .B(n4818), .Z(n4816) );
  XOR U8940 ( .A(y[3635]), .B(x[3635]), .Z(n4818) );
  XOR U8941 ( .A(y[3634]), .B(x[3634]), .Z(n4819) );
  XOR U8942 ( .A(y[3633]), .B(x[3633]), .Z(n4817) );
  XOR U8943 ( .A(n4811), .B(n4810), .Z(n4821) );
  XOR U8944 ( .A(n4813), .B(n4812), .Z(n4810) );
  XOR U8945 ( .A(y[3632]), .B(x[3632]), .Z(n4812) );
  XOR U8946 ( .A(y[3631]), .B(x[3631]), .Z(n4813) );
  XOR U8947 ( .A(y[3630]), .B(x[3630]), .Z(n4811) );
  NAND U8948 ( .A(n4874), .B(n4875), .Z(N29745) );
  NAND U8949 ( .A(n4876), .B(n4877), .Z(n4875) );
  NANDN U8950 ( .A(n4878), .B(n4879), .Z(n4877) );
  NANDN U8951 ( .A(n4879), .B(n4878), .Z(n4874) );
  XOR U8952 ( .A(n4878), .B(n4880), .Z(N29744) );
  XNOR U8953 ( .A(n4876), .B(n4879), .Z(n4880) );
  NAND U8954 ( .A(n4881), .B(n4882), .Z(n4879) );
  NAND U8955 ( .A(n4883), .B(n4884), .Z(n4882) );
  NANDN U8956 ( .A(n4885), .B(n4886), .Z(n4884) );
  NANDN U8957 ( .A(n4886), .B(n4885), .Z(n4881) );
  AND U8958 ( .A(n4887), .B(n4888), .Z(n4876) );
  NAND U8959 ( .A(n4889), .B(n4890), .Z(n4888) );
  OR U8960 ( .A(n4891), .B(n4892), .Z(n4890) );
  NAND U8961 ( .A(n4892), .B(n4891), .Z(n4887) );
  IV U8962 ( .A(n4893), .Z(n4892) );
  AND U8963 ( .A(n4894), .B(n4895), .Z(n4878) );
  NAND U8964 ( .A(n4896), .B(n4897), .Z(n4895) );
  NANDN U8965 ( .A(n4898), .B(n4899), .Z(n4897) );
  NANDN U8966 ( .A(n4899), .B(n4898), .Z(n4894) );
  XOR U8967 ( .A(n4891), .B(n4900), .Z(N29743) );
  XOR U8968 ( .A(n4889), .B(n4893), .Z(n4900) );
  XNOR U8969 ( .A(n4886), .B(n4901), .Z(n4893) );
  XNOR U8970 ( .A(n4883), .B(n4885), .Z(n4901) );
  AND U8971 ( .A(n4902), .B(n4903), .Z(n4885) );
  NANDN U8972 ( .A(n4904), .B(n4905), .Z(n4903) );
  NANDN U8973 ( .A(n4906), .B(n4907), .Z(n4905) );
  IV U8974 ( .A(n4908), .Z(n4907) );
  NAND U8975 ( .A(n4908), .B(n4906), .Z(n4902) );
  AND U8976 ( .A(n4909), .B(n4910), .Z(n4883) );
  NAND U8977 ( .A(n4911), .B(n4912), .Z(n4910) );
  OR U8978 ( .A(n4913), .B(n4914), .Z(n4912) );
  NAND U8979 ( .A(n4914), .B(n4913), .Z(n4909) );
  IV U8980 ( .A(n4915), .Z(n4914) );
  NAND U8981 ( .A(n4916), .B(n4917), .Z(n4886) );
  NANDN U8982 ( .A(n4918), .B(n4919), .Z(n4917) );
  NAND U8983 ( .A(n4920), .B(n4921), .Z(n4919) );
  OR U8984 ( .A(n4921), .B(n4920), .Z(n4916) );
  IV U8985 ( .A(n4922), .Z(n4920) );
  AND U8986 ( .A(n4923), .B(n4924), .Z(n4889) );
  NAND U8987 ( .A(n4925), .B(n4926), .Z(n4924) );
  NANDN U8988 ( .A(n4927), .B(n4928), .Z(n4926) );
  NANDN U8989 ( .A(n4928), .B(n4927), .Z(n4923) );
  XOR U8990 ( .A(n4899), .B(n4929), .Z(n4891) );
  XNOR U8991 ( .A(n4896), .B(n4898), .Z(n4929) );
  AND U8992 ( .A(n4930), .B(n4931), .Z(n4898) );
  NANDN U8993 ( .A(n4932), .B(n4933), .Z(n4931) );
  NANDN U8994 ( .A(n4934), .B(n4935), .Z(n4933) );
  IV U8995 ( .A(n4936), .Z(n4935) );
  NAND U8996 ( .A(n4936), .B(n4934), .Z(n4930) );
  AND U8997 ( .A(n4937), .B(n4938), .Z(n4896) );
  NAND U8998 ( .A(n4939), .B(n4940), .Z(n4938) );
  OR U8999 ( .A(n4941), .B(n4942), .Z(n4940) );
  NAND U9000 ( .A(n4942), .B(n4941), .Z(n4937) );
  IV U9001 ( .A(n4943), .Z(n4942) );
  NAND U9002 ( .A(n4944), .B(n4945), .Z(n4899) );
  NANDN U9003 ( .A(n4946), .B(n4947), .Z(n4945) );
  NAND U9004 ( .A(n4948), .B(n4949), .Z(n4947) );
  OR U9005 ( .A(n4949), .B(n4948), .Z(n4944) );
  IV U9006 ( .A(n4950), .Z(n4948) );
  XOR U9007 ( .A(n4925), .B(n4951), .Z(N29742) );
  XNOR U9008 ( .A(n4928), .B(n4927), .Z(n4951) );
  XNOR U9009 ( .A(n4939), .B(n4952), .Z(n4927) );
  XOR U9010 ( .A(n4943), .B(n4941), .Z(n4952) );
  XOR U9011 ( .A(n4949), .B(n4953), .Z(n4941) );
  XOR U9012 ( .A(n4946), .B(n4950), .Z(n4953) );
  NAND U9013 ( .A(n4954), .B(n4955), .Z(n4950) );
  NAND U9014 ( .A(n4956), .B(n4957), .Z(n4955) );
  NAND U9015 ( .A(n4958), .B(n4959), .Z(n4954) );
  AND U9016 ( .A(n4960), .B(n4961), .Z(n4946) );
  NAND U9017 ( .A(n4962), .B(n4963), .Z(n4961) );
  NAND U9018 ( .A(n4964), .B(n4965), .Z(n4960) );
  NANDN U9019 ( .A(n4966), .B(n4967), .Z(n4949) );
  NANDN U9020 ( .A(n4968), .B(n4969), .Z(n4943) );
  XNOR U9021 ( .A(n4934), .B(n4970), .Z(n4939) );
  XOR U9022 ( .A(n4932), .B(n4936), .Z(n4970) );
  NAND U9023 ( .A(n4971), .B(n4972), .Z(n4936) );
  NAND U9024 ( .A(n4973), .B(n4974), .Z(n4972) );
  NAND U9025 ( .A(n4975), .B(n4976), .Z(n4971) );
  AND U9026 ( .A(n4977), .B(n4978), .Z(n4932) );
  NAND U9027 ( .A(n4979), .B(n4980), .Z(n4978) );
  NAND U9028 ( .A(n4981), .B(n4982), .Z(n4977) );
  AND U9029 ( .A(n4983), .B(n4984), .Z(n4934) );
  NAND U9030 ( .A(n4985), .B(n4986), .Z(n4928) );
  XNOR U9031 ( .A(n4911), .B(n4987), .Z(n4925) );
  XOR U9032 ( .A(n4915), .B(n4913), .Z(n4987) );
  XOR U9033 ( .A(n4921), .B(n4988), .Z(n4913) );
  XOR U9034 ( .A(n4918), .B(n4922), .Z(n4988) );
  NAND U9035 ( .A(n4989), .B(n4990), .Z(n4922) );
  NAND U9036 ( .A(n4991), .B(n4992), .Z(n4990) );
  NAND U9037 ( .A(n4993), .B(n4994), .Z(n4989) );
  AND U9038 ( .A(n4995), .B(n4996), .Z(n4918) );
  NAND U9039 ( .A(n4997), .B(n4998), .Z(n4996) );
  NAND U9040 ( .A(n4999), .B(n5000), .Z(n4995) );
  NANDN U9041 ( .A(n5001), .B(n5002), .Z(n4921) );
  NANDN U9042 ( .A(n5003), .B(n5004), .Z(n4915) );
  XNOR U9043 ( .A(n4906), .B(n5005), .Z(n4911) );
  XOR U9044 ( .A(n4904), .B(n4908), .Z(n5005) );
  NAND U9045 ( .A(n5006), .B(n5007), .Z(n4908) );
  NAND U9046 ( .A(n5008), .B(n5009), .Z(n5007) );
  NAND U9047 ( .A(n5010), .B(n5011), .Z(n5006) );
  AND U9048 ( .A(n5012), .B(n5013), .Z(n4904) );
  NAND U9049 ( .A(n5014), .B(n5015), .Z(n5013) );
  NAND U9050 ( .A(n5016), .B(n5017), .Z(n5012) );
  AND U9051 ( .A(n5018), .B(n5019), .Z(n4906) );
  XOR U9052 ( .A(n4986), .B(n4985), .Z(N29741) );
  XNOR U9053 ( .A(n5004), .B(n5003), .Z(n4985) );
  XNOR U9054 ( .A(n5018), .B(n5019), .Z(n5003) );
  XOR U9055 ( .A(n5015), .B(n5014), .Z(n5019) );
  XOR U9056 ( .A(y[3627]), .B(x[3627]), .Z(n5014) );
  XOR U9057 ( .A(n5017), .B(n5016), .Z(n5015) );
  XOR U9058 ( .A(y[3629]), .B(x[3629]), .Z(n5016) );
  XOR U9059 ( .A(y[3628]), .B(x[3628]), .Z(n5017) );
  XOR U9060 ( .A(n5009), .B(n5008), .Z(n5018) );
  XOR U9061 ( .A(n5011), .B(n5010), .Z(n5008) );
  XOR U9062 ( .A(y[3626]), .B(x[3626]), .Z(n5010) );
  XOR U9063 ( .A(y[3625]), .B(x[3625]), .Z(n5011) );
  XOR U9064 ( .A(y[3624]), .B(x[3624]), .Z(n5009) );
  XNOR U9065 ( .A(n5002), .B(n5001), .Z(n5004) );
  XNOR U9066 ( .A(n4998), .B(n4997), .Z(n5001) );
  XOR U9067 ( .A(n5000), .B(n4999), .Z(n4997) );
  XOR U9068 ( .A(y[3623]), .B(x[3623]), .Z(n4999) );
  XOR U9069 ( .A(y[3622]), .B(x[3622]), .Z(n5000) );
  XOR U9070 ( .A(y[3621]), .B(x[3621]), .Z(n4998) );
  XOR U9071 ( .A(n4992), .B(n4991), .Z(n5002) );
  XOR U9072 ( .A(n4994), .B(n4993), .Z(n4991) );
  XOR U9073 ( .A(y[3620]), .B(x[3620]), .Z(n4993) );
  XOR U9074 ( .A(y[3619]), .B(x[3619]), .Z(n4994) );
  XOR U9075 ( .A(y[3618]), .B(x[3618]), .Z(n4992) );
  XNOR U9076 ( .A(n4969), .B(n4968), .Z(n4986) );
  XNOR U9077 ( .A(n4983), .B(n4984), .Z(n4968) );
  XOR U9078 ( .A(n4980), .B(n4979), .Z(n4984) );
  XOR U9079 ( .A(y[3615]), .B(x[3615]), .Z(n4979) );
  XOR U9080 ( .A(n4982), .B(n4981), .Z(n4980) );
  XOR U9081 ( .A(y[3617]), .B(x[3617]), .Z(n4981) );
  XOR U9082 ( .A(y[3616]), .B(x[3616]), .Z(n4982) );
  XOR U9083 ( .A(n4974), .B(n4973), .Z(n4983) );
  XOR U9084 ( .A(n4976), .B(n4975), .Z(n4973) );
  XOR U9085 ( .A(y[3614]), .B(x[3614]), .Z(n4975) );
  XOR U9086 ( .A(y[3613]), .B(x[3613]), .Z(n4976) );
  XOR U9087 ( .A(y[3612]), .B(x[3612]), .Z(n4974) );
  XNOR U9088 ( .A(n4967), .B(n4966), .Z(n4969) );
  XNOR U9089 ( .A(n4963), .B(n4962), .Z(n4966) );
  XOR U9090 ( .A(n4965), .B(n4964), .Z(n4962) );
  XOR U9091 ( .A(y[3611]), .B(x[3611]), .Z(n4964) );
  XOR U9092 ( .A(y[3610]), .B(x[3610]), .Z(n4965) );
  XOR U9093 ( .A(y[3609]), .B(x[3609]), .Z(n4963) );
  XOR U9094 ( .A(n4957), .B(n4956), .Z(n4967) );
  XOR U9095 ( .A(n4959), .B(n4958), .Z(n4956) );
  XOR U9096 ( .A(y[3608]), .B(x[3608]), .Z(n4958) );
  XOR U9097 ( .A(y[3607]), .B(x[3607]), .Z(n4959) );
  XOR U9098 ( .A(y[3606]), .B(x[3606]), .Z(n4957) );
  NAND U9099 ( .A(n5020), .B(n5021), .Z(N29733) );
  NAND U9100 ( .A(n5022), .B(n5023), .Z(n5021) );
  NANDN U9101 ( .A(n5024), .B(n5025), .Z(n5023) );
  NANDN U9102 ( .A(n5025), .B(n5024), .Z(n5020) );
  XOR U9103 ( .A(n5024), .B(n5026), .Z(N29732) );
  XNOR U9104 ( .A(n5022), .B(n5025), .Z(n5026) );
  NAND U9105 ( .A(n5027), .B(n5028), .Z(n5025) );
  NAND U9106 ( .A(n5029), .B(n5030), .Z(n5028) );
  NANDN U9107 ( .A(n5031), .B(n5032), .Z(n5030) );
  NANDN U9108 ( .A(n5032), .B(n5031), .Z(n5027) );
  AND U9109 ( .A(n5033), .B(n5034), .Z(n5022) );
  NAND U9110 ( .A(n5035), .B(n5036), .Z(n5034) );
  OR U9111 ( .A(n5037), .B(n5038), .Z(n5036) );
  NAND U9112 ( .A(n5038), .B(n5037), .Z(n5033) );
  IV U9113 ( .A(n5039), .Z(n5038) );
  AND U9114 ( .A(n5040), .B(n5041), .Z(n5024) );
  NAND U9115 ( .A(n5042), .B(n5043), .Z(n5041) );
  NANDN U9116 ( .A(n5044), .B(n5045), .Z(n5043) );
  NANDN U9117 ( .A(n5045), .B(n5044), .Z(n5040) );
  XOR U9118 ( .A(n5037), .B(n5046), .Z(N29731) );
  XOR U9119 ( .A(n5035), .B(n5039), .Z(n5046) );
  XNOR U9120 ( .A(n5032), .B(n5047), .Z(n5039) );
  XNOR U9121 ( .A(n5029), .B(n5031), .Z(n5047) );
  AND U9122 ( .A(n5048), .B(n5049), .Z(n5031) );
  NANDN U9123 ( .A(n5050), .B(n5051), .Z(n5049) );
  NANDN U9124 ( .A(n5052), .B(n5053), .Z(n5051) );
  IV U9125 ( .A(n5054), .Z(n5053) );
  NAND U9126 ( .A(n5054), .B(n5052), .Z(n5048) );
  AND U9127 ( .A(n5055), .B(n5056), .Z(n5029) );
  NAND U9128 ( .A(n5057), .B(n5058), .Z(n5056) );
  OR U9129 ( .A(n5059), .B(n5060), .Z(n5058) );
  NAND U9130 ( .A(n5060), .B(n5059), .Z(n5055) );
  IV U9131 ( .A(n5061), .Z(n5060) );
  NAND U9132 ( .A(n5062), .B(n5063), .Z(n5032) );
  NANDN U9133 ( .A(n5064), .B(n5065), .Z(n5063) );
  NAND U9134 ( .A(n5066), .B(n5067), .Z(n5065) );
  OR U9135 ( .A(n5067), .B(n5066), .Z(n5062) );
  IV U9136 ( .A(n5068), .Z(n5066) );
  AND U9137 ( .A(n5069), .B(n5070), .Z(n5035) );
  NAND U9138 ( .A(n5071), .B(n5072), .Z(n5070) );
  NANDN U9139 ( .A(n5073), .B(n5074), .Z(n5072) );
  NANDN U9140 ( .A(n5074), .B(n5073), .Z(n5069) );
  XOR U9141 ( .A(n5045), .B(n5075), .Z(n5037) );
  XNOR U9142 ( .A(n5042), .B(n5044), .Z(n5075) );
  AND U9143 ( .A(n5076), .B(n5077), .Z(n5044) );
  NANDN U9144 ( .A(n5078), .B(n5079), .Z(n5077) );
  NANDN U9145 ( .A(n5080), .B(n5081), .Z(n5079) );
  IV U9146 ( .A(n5082), .Z(n5081) );
  NAND U9147 ( .A(n5082), .B(n5080), .Z(n5076) );
  AND U9148 ( .A(n5083), .B(n5084), .Z(n5042) );
  NAND U9149 ( .A(n5085), .B(n5086), .Z(n5084) );
  OR U9150 ( .A(n5087), .B(n5088), .Z(n5086) );
  NAND U9151 ( .A(n5088), .B(n5087), .Z(n5083) );
  IV U9152 ( .A(n5089), .Z(n5088) );
  NAND U9153 ( .A(n5090), .B(n5091), .Z(n5045) );
  NANDN U9154 ( .A(n5092), .B(n5093), .Z(n5091) );
  NAND U9155 ( .A(n5094), .B(n5095), .Z(n5093) );
  OR U9156 ( .A(n5095), .B(n5094), .Z(n5090) );
  IV U9157 ( .A(n5096), .Z(n5094) );
  XOR U9158 ( .A(n5071), .B(n5097), .Z(N29730) );
  XNOR U9159 ( .A(n5074), .B(n5073), .Z(n5097) );
  XNOR U9160 ( .A(n5085), .B(n5098), .Z(n5073) );
  XOR U9161 ( .A(n5089), .B(n5087), .Z(n5098) );
  XOR U9162 ( .A(n5095), .B(n5099), .Z(n5087) );
  XOR U9163 ( .A(n5092), .B(n5096), .Z(n5099) );
  NAND U9164 ( .A(n5100), .B(n5101), .Z(n5096) );
  NAND U9165 ( .A(n5102), .B(n5103), .Z(n5101) );
  NAND U9166 ( .A(n5104), .B(n5105), .Z(n5100) );
  AND U9167 ( .A(n5106), .B(n5107), .Z(n5092) );
  NAND U9168 ( .A(n5108), .B(n5109), .Z(n5107) );
  NAND U9169 ( .A(n5110), .B(n5111), .Z(n5106) );
  NANDN U9170 ( .A(n5112), .B(n5113), .Z(n5095) );
  NANDN U9171 ( .A(n5114), .B(n5115), .Z(n5089) );
  XNOR U9172 ( .A(n5080), .B(n5116), .Z(n5085) );
  XOR U9173 ( .A(n5078), .B(n5082), .Z(n5116) );
  NAND U9174 ( .A(n5117), .B(n5118), .Z(n5082) );
  NAND U9175 ( .A(n5119), .B(n5120), .Z(n5118) );
  NAND U9176 ( .A(n5121), .B(n5122), .Z(n5117) );
  AND U9177 ( .A(n5123), .B(n5124), .Z(n5078) );
  NAND U9178 ( .A(n5125), .B(n5126), .Z(n5124) );
  NAND U9179 ( .A(n5127), .B(n5128), .Z(n5123) );
  AND U9180 ( .A(n5129), .B(n5130), .Z(n5080) );
  NAND U9181 ( .A(n5131), .B(n5132), .Z(n5074) );
  XNOR U9182 ( .A(n5057), .B(n5133), .Z(n5071) );
  XOR U9183 ( .A(n5061), .B(n5059), .Z(n5133) );
  XOR U9184 ( .A(n5067), .B(n5134), .Z(n5059) );
  XOR U9185 ( .A(n5064), .B(n5068), .Z(n5134) );
  NAND U9186 ( .A(n5135), .B(n5136), .Z(n5068) );
  NAND U9187 ( .A(n5137), .B(n5138), .Z(n5136) );
  NAND U9188 ( .A(n5139), .B(n5140), .Z(n5135) );
  AND U9189 ( .A(n5141), .B(n5142), .Z(n5064) );
  NAND U9190 ( .A(n5143), .B(n5144), .Z(n5142) );
  NAND U9191 ( .A(n5145), .B(n5146), .Z(n5141) );
  NANDN U9192 ( .A(n5147), .B(n5148), .Z(n5067) );
  NANDN U9193 ( .A(n5149), .B(n5150), .Z(n5061) );
  XNOR U9194 ( .A(n5052), .B(n5151), .Z(n5057) );
  XOR U9195 ( .A(n5050), .B(n5054), .Z(n5151) );
  NAND U9196 ( .A(n5152), .B(n5153), .Z(n5054) );
  NAND U9197 ( .A(n5154), .B(n5155), .Z(n5153) );
  NAND U9198 ( .A(n5156), .B(n5157), .Z(n5152) );
  AND U9199 ( .A(n5158), .B(n5159), .Z(n5050) );
  NAND U9200 ( .A(n5160), .B(n5161), .Z(n5159) );
  NAND U9201 ( .A(n5162), .B(n5163), .Z(n5158) );
  AND U9202 ( .A(n5164), .B(n5165), .Z(n5052) );
  XOR U9203 ( .A(n5132), .B(n5131), .Z(N29729) );
  XNOR U9204 ( .A(n5150), .B(n5149), .Z(n5131) );
  XNOR U9205 ( .A(n5164), .B(n5165), .Z(n5149) );
  XOR U9206 ( .A(n5161), .B(n5160), .Z(n5165) );
  XOR U9207 ( .A(y[3603]), .B(x[3603]), .Z(n5160) );
  XOR U9208 ( .A(n5163), .B(n5162), .Z(n5161) );
  XOR U9209 ( .A(y[3605]), .B(x[3605]), .Z(n5162) );
  XOR U9210 ( .A(y[3604]), .B(x[3604]), .Z(n5163) );
  XOR U9211 ( .A(n5155), .B(n5154), .Z(n5164) );
  XOR U9212 ( .A(n5157), .B(n5156), .Z(n5154) );
  XOR U9213 ( .A(y[3602]), .B(x[3602]), .Z(n5156) );
  XOR U9214 ( .A(y[3601]), .B(x[3601]), .Z(n5157) );
  XOR U9215 ( .A(y[3600]), .B(x[3600]), .Z(n5155) );
  XNOR U9216 ( .A(n5148), .B(n5147), .Z(n5150) );
  XNOR U9217 ( .A(n5144), .B(n5143), .Z(n5147) );
  XOR U9218 ( .A(n5146), .B(n5145), .Z(n5143) );
  XOR U9219 ( .A(y[3599]), .B(x[3599]), .Z(n5145) );
  XOR U9220 ( .A(y[3598]), .B(x[3598]), .Z(n5146) );
  XOR U9221 ( .A(y[3597]), .B(x[3597]), .Z(n5144) );
  XOR U9222 ( .A(n5138), .B(n5137), .Z(n5148) );
  XOR U9223 ( .A(n5140), .B(n5139), .Z(n5137) );
  XOR U9224 ( .A(y[3596]), .B(x[3596]), .Z(n5139) );
  XOR U9225 ( .A(y[3595]), .B(x[3595]), .Z(n5140) );
  XOR U9226 ( .A(y[3594]), .B(x[3594]), .Z(n5138) );
  XNOR U9227 ( .A(n5115), .B(n5114), .Z(n5132) );
  XNOR U9228 ( .A(n5129), .B(n5130), .Z(n5114) );
  XOR U9229 ( .A(n5126), .B(n5125), .Z(n5130) );
  XOR U9230 ( .A(y[3591]), .B(x[3591]), .Z(n5125) );
  XOR U9231 ( .A(n5128), .B(n5127), .Z(n5126) );
  XOR U9232 ( .A(y[3593]), .B(x[3593]), .Z(n5127) );
  XOR U9233 ( .A(y[3592]), .B(x[3592]), .Z(n5128) );
  XOR U9234 ( .A(n5120), .B(n5119), .Z(n5129) );
  XOR U9235 ( .A(n5122), .B(n5121), .Z(n5119) );
  XOR U9236 ( .A(y[3590]), .B(x[3590]), .Z(n5121) );
  XOR U9237 ( .A(y[3589]), .B(x[3589]), .Z(n5122) );
  XOR U9238 ( .A(y[3588]), .B(x[3588]), .Z(n5120) );
  XNOR U9239 ( .A(n5113), .B(n5112), .Z(n5115) );
  XNOR U9240 ( .A(n5109), .B(n5108), .Z(n5112) );
  XOR U9241 ( .A(n5111), .B(n5110), .Z(n5108) );
  XOR U9242 ( .A(y[3587]), .B(x[3587]), .Z(n5110) );
  XOR U9243 ( .A(y[3586]), .B(x[3586]), .Z(n5111) );
  XOR U9244 ( .A(y[3585]), .B(x[3585]), .Z(n5109) );
  XOR U9245 ( .A(n5103), .B(n5102), .Z(n5113) );
  XOR U9246 ( .A(n5105), .B(n5104), .Z(n5102) );
  XOR U9247 ( .A(y[3584]), .B(x[3584]), .Z(n5104) );
  XOR U9248 ( .A(y[3583]), .B(x[3583]), .Z(n5105) );
  XOR U9249 ( .A(y[3582]), .B(x[3582]), .Z(n5103) );
  NAND U9250 ( .A(n5166), .B(n5167), .Z(N29721) );
  NAND U9251 ( .A(n5168), .B(n5169), .Z(n5167) );
  NANDN U9252 ( .A(n5170), .B(n5171), .Z(n5169) );
  NANDN U9253 ( .A(n5171), .B(n5170), .Z(n5166) );
  XOR U9254 ( .A(n5170), .B(n5172), .Z(N29720) );
  XNOR U9255 ( .A(n5168), .B(n5171), .Z(n5172) );
  NAND U9256 ( .A(n5173), .B(n5174), .Z(n5171) );
  NAND U9257 ( .A(n5175), .B(n5176), .Z(n5174) );
  NANDN U9258 ( .A(n5177), .B(n5178), .Z(n5176) );
  NANDN U9259 ( .A(n5178), .B(n5177), .Z(n5173) );
  AND U9260 ( .A(n5179), .B(n5180), .Z(n5168) );
  NAND U9261 ( .A(n5181), .B(n5182), .Z(n5180) );
  OR U9262 ( .A(n5183), .B(n5184), .Z(n5182) );
  NAND U9263 ( .A(n5184), .B(n5183), .Z(n5179) );
  IV U9264 ( .A(n5185), .Z(n5184) );
  AND U9265 ( .A(n5186), .B(n5187), .Z(n5170) );
  NAND U9266 ( .A(n5188), .B(n5189), .Z(n5187) );
  NANDN U9267 ( .A(n5190), .B(n5191), .Z(n5189) );
  NANDN U9268 ( .A(n5191), .B(n5190), .Z(n5186) );
  XOR U9269 ( .A(n5183), .B(n5192), .Z(N29719) );
  XOR U9270 ( .A(n5181), .B(n5185), .Z(n5192) );
  XNOR U9271 ( .A(n5178), .B(n5193), .Z(n5185) );
  XNOR U9272 ( .A(n5175), .B(n5177), .Z(n5193) );
  AND U9273 ( .A(n5194), .B(n5195), .Z(n5177) );
  NANDN U9274 ( .A(n5196), .B(n5197), .Z(n5195) );
  NANDN U9275 ( .A(n5198), .B(n5199), .Z(n5197) );
  IV U9276 ( .A(n5200), .Z(n5199) );
  NAND U9277 ( .A(n5200), .B(n5198), .Z(n5194) );
  AND U9278 ( .A(n5201), .B(n5202), .Z(n5175) );
  NAND U9279 ( .A(n5203), .B(n5204), .Z(n5202) );
  OR U9280 ( .A(n5205), .B(n5206), .Z(n5204) );
  NAND U9281 ( .A(n5206), .B(n5205), .Z(n5201) );
  IV U9282 ( .A(n5207), .Z(n5206) );
  NAND U9283 ( .A(n5208), .B(n5209), .Z(n5178) );
  NANDN U9284 ( .A(n5210), .B(n5211), .Z(n5209) );
  NAND U9285 ( .A(n5212), .B(n5213), .Z(n5211) );
  OR U9286 ( .A(n5213), .B(n5212), .Z(n5208) );
  IV U9287 ( .A(n5214), .Z(n5212) );
  AND U9288 ( .A(n5215), .B(n5216), .Z(n5181) );
  NAND U9289 ( .A(n5217), .B(n5218), .Z(n5216) );
  NANDN U9290 ( .A(n5219), .B(n5220), .Z(n5218) );
  NANDN U9291 ( .A(n5220), .B(n5219), .Z(n5215) );
  XOR U9292 ( .A(n5191), .B(n5221), .Z(n5183) );
  XNOR U9293 ( .A(n5188), .B(n5190), .Z(n5221) );
  AND U9294 ( .A(n5222), .B(n5223), .Z(n5190) );
  NANDN U9295 ( .A(n5224), .B(n5225), .Z(n5223) );
  NANDN U9296 ( .A(n5226), .B(n5227), .Z(n5225) );
  IV U9297 ( .A(n5228), .Z(n5227) );
  NAND U9298 ( .A(n5228), .B(n5226), .Z(n5222) );
  AND U9299 ( .A(n5229), .B(n5230), .Z(n5188) );
  NAND U9300 ( .A(n5231), .B(n5232), .Z(n5230) );
  OR U9301 ( .A(n5233), .B(n5234), .Z(n5232) );
  NAND U9302 ( .A(n5234), .B(n5233), .Z(n5229) );
  IV U9303 ( .A(n5235), .Z(n5234) );
  NAND U9304 ( .A(n5236), .B(n5237), .Z(n5191) );
  NANDN U9305 ( .A(n5238), .B(n5239), .Z(n5237) );
  NAND U9306 ( .A(n5240), .B(n5241), .Z(n5239) );
  OR U9307 ( .A(n5241), .B(n5240), .Z(n5236) );
  IV U9308 ( .A(n5242), .Z(n5240) );
  XOR U9309 ( .A(n5217), .B(n5243), .Z(N29718) );
  XNOR U9310 ( .A(n5220), .B(n5219), .Z(n5243) );
  XNOR U9311 ( .A(n5231), .B(n5244), .Z(n5219) );
  XOR U9312 ( .A(n5235), .B(n5233), .Z(n5244) );
  XOR U9313 ( .A(n5241), .B(n5245), .Z(n5233) );
  XOR U9314 ( .A(n5238), .B(n5242), .Z(n5245) );
  NAND U9315 ( .A(n5246), .B(n5247), .Z(n5242) );
  NAND U9316 ( .A(n5248), .B(n5249), .Z(n5247) );
  NAND U9317 ( .A(n5250), .B(n5251), .Z(n5246) );
  AND U9318 ( .A(n5252), .B(n5253), .Z(n5238) );
  NAND U9319 ( .A(n5254), .B(n5255), .Z(n5253) );
  NAND U9320 ( .A(n5256), .B(n5257), .Z(n5252) );
  NANDN U9321 ( .A(n5258), .B(n5259), .Z(n5241) );
  NANDN U9322 ( .A(n5260), .B(n5261), .Z(n5235) );
  XNOR U9323 ( .A(n5226), .B(n5262), .Z(n5231) );
  XOR U9324 ( .A(n5224), .B(n5228), .Z(n5262) );
  NAND U9325 ( .A(n5263), .B(n5264), .Z(n5228) );
  NAND U9326 ( .A(n5265), .B(n5266), .Z(n5264) );
  NAND U9327 ( .A(n5267), .B(n5268), .Z(n5263) );
  AND U9328 ( .A(n5269), .B(n5270), .Z(n5224) );
  NAND U9329 ( .A(n5271), .B(n5272), .Z(n5270) );
  NAND U9330 ( .A(n5273), .B(n5274), .Z(n5269) );
  AND U9331 ( .A(n5275), .B(n5276), .Z(n5226) );
  NAND U9332 ( .A(n5277), .B(n5278), .Z(n5220) );
  XNOR U9333 ( .A(n5203), .B(n5279), .Z(n5217) );
  XOR U9334 ( .A(n5207), .B(n5205), .Z(n5279) );
  XOR U9335 ( .A(n5213), .B(n5280), .Z(n5205) );
  XOR U9336 ( .A(n5210), .B(n5214), .Z(n5280) );
  NAND U9337 ( .A(n5281), .B(n5282), .Z(n5214) );
  NAND U9338 ( .A(n5283), .B(n5284), .Z(n5282) );
  NAND U9339 ( .A(n5285), .B(n5286), .Z(n5281) );
  AND U9340 ( .A(n5287), .B(n5288), .Z(n5210) );
  NAND U9341 ( .A(n5289), .B(n5290), .Z(n5288) );
  NAND U9342 ( .A(n5291), .B(n5292), .Z(n5287) );
  NANDN U9343 ( .A(n5293), .B(n5294), .Z(n5213) );
  NANDN U9344 ( .A(n5295), .B(n5296), .Z(n5207) );
  XNOR U9345 ( .A(n5198), .B(n5297), .Z(n5203) );
  XOR U9346 ( .A(n5196), .B(n5200), .Z(n5297) );
  NAND U9347 ( .A(n5298), .B(n5299), .Z(n5200) );
  NAND U9348 ( .A(n5300), .B(n5301), .Z(n5299) );
  NAND U9349 ( .A(n5302), .B(n5303), .Z(n5298) );
  AND U9350 ( .A(n5304), .B(n5305), .Z(n5196) );
  NAND U9351 ( .A(n5306), .B(n5307), .Z(n5305) );
  NAND U9352 ( .A(n5308), .B(n5309), .Z(n5304) );
  AND U9353 ( .A(n5310), .B(n5311), .Z(n5198) );
  XOR U9354 ( .A(n5278), .B(n5277), .Z(N29717) );
  XNOR U9355 ( .A(n5296), .B(n5295), .Z(n5277) );
  XNOR U9356 ( .A(n5310), .B(n5311), .Z(n5295) );
  XOR U9357 ( .A(n5307), .B(n5306), .Z(n5311) );
  XOR U9358 ( .A(y[3579]), .B(x[3579]), .Z(n5306) );
  XOR U9359 ( .A(n5309), .B(n5308), .Z(n5307) );
  XOR U9360 ( .A(y[3581]), .B(x[3581]), .Z(n5308) );
  XOR U9361 ( .A(y[3580]), .B(x[3580]), .Z(n5309) );
  XOR U9362 ( .A(n5301), .B(n5300), .Z(n5310) );
  XOR U9363 ( .A(n5303), .B(n5302), .Z(n5300) );
  XOR U9364 ( .A(y[3578]), .B(x[3578]), .Z(n5302) );
  XOR U9365 ( .A(y[3577]), .B(x[3577]), .Z(n5303) );
  XOR U9366 ( .A(y[3576]), .B(x[3576]), .Z(n5301) );
  XNOR U9367 ( .A(n5294), .B(n5293), .Z(n5296) );
  XNOR U9368 ( .A(n5290), .B(n5289), .Z(n5293) );
  XOR U9369 ( .A(n5292), .B(n5291), .Z(n5289) );
  XOR U9370 ( .A(y[3575]), .B(x[3575]), .Z(n5291) );
  XOR U9371 ( .A(y[3574]), .B(x[3574]), .Z(n5292) );
  XOR U9372 ( .A(y[3573]), .B(x[3573]), .Z(n5290) );
  XOR U9373 ( .A(n5284), .B(n5283), .Z(n5294) );
  XOR U9374 ( .A(n5286), .B(n5285), .Z(n5283) );
  XOR U9375 ( .A(y[3572]), .B(x[3572]), .Z(n5285) );
  XOR U9376 ( .A(y[3571]), .B(x[3571]), .Z(n5286) );
  XOR U9377 ( .A(y[3570]), .B(x[3570]), .Z(n5284) );
  XNOR U9378 ( .A(n5261), .B(n5260), .Z(n5278) );
  XNOR U9379 ( .A(n5275), .B(n5276), .Z(n5260) );
  XOR U9380 ( .A(n5272), .B(n5271), .Z(n5276) );
  XOR U9381 ( .A(y[3567]), .B(x[3567]), .Z(n5271) );
  XOR U9382 ( .A(n5274), .B(n5273), .Z(n5272) );
  XOR U9383 ( .A(y[3569]), .B(x[3569]), .Z(n5273) );
  XOR U9384 ( .A(y[3568]), .B(x[3568]), .Z(n5274) );
  XOR U9385 ( .A(n5266), .B(n5265), .Z(n5275) );
  XOR U9386 ( .A(n5268), .B(n5267), .Z(n5265) );
  XOR U9387 ( .A(y[3566]), .B(x[3566]), .Z(n5267) );
  XOR U9388 ( .A(y[3565]), .B(x[3565]), .Z(n5268) );
  XOR U9389 ( .A(y[3564]), .B(x[3564]), .Z(n5266) );
  XNOR U9390 ( .A(n5259), .B(n5258), .Z(n5261) );
  XNOR U9391 ( .A(n5255), .B(n5254), .Z(n5258) );
  XOR U9392 ( .A(n5257), .B(n5256), .Z(n5254) );
  XOR U9393 ( .A(y[3563]), .B(x[3563]), .Z(n5256) );
  XOR U9394 ( .A(y[3562]), .B(x[3562]), .Z(n5257) );
  XOR U9395 ( .A(y[3561]), .B(x[3561]), .Z(n5255) );
  XOR U9396 ( .A(n5249), .B(n5248), .Z(n5259) );
  XOR U9397 ( .A(n5251), .B(n5250), .Z(n5248) );
  XOR U9398 ( .A(y[3560]), .B(x[3560]), .Z(n5250) );
  XOR U9399 ( .A(y[3559]), .B(x[3559]), .Z(n5251) );
  XOR U9400 ( .A(y[3558]), .B(x[3558]), .Z(n5249) );
  NAND U9401 ( .A(n5312), .B(n5313), .Z(N29709) );
  NAND U9402 ( .A(n5314), .B(n5315), .Z(n5313) );
  NANDN U9403 ( .A(n5316), .B(n5317), .Z(n5315) );
  NANDN U9404 ( .A(n5317), .B(n5316), .Z(n5312) );
  XOR U9405 ( .A(n5316), .B(n5318), .Z(N29708) );
  XNOR U9406 ( .A(n5314), .B(n5317), .Z(n5318) );
  NAND U9407 ( .A(n5319), .B(n5320), .Z(n5317) );
  NAND U9408 ( .A(n5321), .B(n5322), .Z(n5320) );
  NANDN U9409 ( .A(n5323), .B(n5324), .Z(n5322) );
  NANDN U9410 ( .A(n5324), .B(n5323), .Z(n5319) );
  AND U9411 ( .A(n5325), .B(n5326), .Z(n5314) );
  NAND U9412 ( .A(n5327), .B(n5328), .Z(n5326) );
  OR U9413 ( .A(n5329), .B(n5330), .Z(n5328) );
  NAND U9414 ( .A(n5330), .B(n5329), .Z(n5325) );
  IV U9415 ( .A(n5331), .Z(n5330) );
  AND U9416 ( .A(n5332), .B(n5333), .Z(n5316) );
  NAND U9417 ( .A(n5334), .B(n5335), .Z(n5333) );
  NANDN U9418 ( .A(n5336), .B(n5337), .Z(n5335) );
  NANDN U9419 ( .A(n5337), .B(n5336), .Z(n5332) );
  XOR U9420 ( .A(n5329), .B(n5338), .Z(N29707) );
  XOR U9421 ( .A(n5327), .B(n5331), .Z(n5338) );
  XNOR U9422 ( .A(n5324), .B(n5339), .Z(n5331) );
  XNOR U9423 ( .A(n5321), .B(n5323), .Z(n5339) );
  AND U9424 ( .A(n5340), .B(n5341), .Z(n5323) );
  NANDN U9425 ( .A(n5342), .B(n5343), .Z(n5341) );
  NANDN U9426 ( .A(n5344), .B(n5345), .Z(n5343) );
  IV U9427 ( .A(n5346), .Z(n5345) );
  NAND U9428 ( .A(n5346), .B(n5344), .Z(n5340) );
  AND U9429 ( .A(n5347), .B(n5348), .Z(n5321) );
  NAND U9430 ( .A(n5349), .B(n5350), .Z(n5348) );
  OR U9431 ( .A(n5351), .B(n5352), .Z(n5350) );
  NAND U9432 ( .A(n5352), .B(n5351), .Z(n5347) );
  IV U9433 ( .A(n5353), .Z(n5352) );
  NAND U9434 ( .A(n5354), .B(n5355), .Z(n5324) );
  NANDN U9435 ( .A(n5356), .B(n5357), .Z(n5355) );
  NAND U9436 ( .A(n5358), .B(n5359), .Z(n5357) );
  OR U9437 ( .A(n5359), .B(n5358), .Z(n5354) );
  IV U9438 ( .A(n5360), .Z(n5358) );
  AND U9439 ( .A(n5361), .B(n5362), .Z(n5327) );
  NAND U9440 ( .A(n5363), .B(n5364), .Z(n5362) );
  NANDN U9441 ( .A(n5365), .B(n5366), .Z(n5364) );
  NANDN U9442 ( .A(n5366), .B(n5365), .Z(n5361) );
  XOR U9443 ( .A(n5337), .B(n5367), .Z(n5329) );
  XNOR U9444 ( .A(n5334), .B(n5336), .Z(n5367) );
  AND U9445 ( .A(n5368), .B(n5369), .Z(n5336) );
  NANDN U9446 ( .A(n5370), .B(n5371), .Z(n5369) );
  NANDN U9447 ( .A(n5372), .B(n5373), .Z(n5371) );
  IV U9448 ( .A(n5374), .Z(n5373) );
  NAND U9449 ( .A(n5374), .B(n5372), .Z(n5368) );
  AND U9450 ( .A(n5375), .B(n5376), .Z(n5334) );
  NAND U9451 ( .A(n5377), .B(n5378), .Z(n5376) );
  OR U9452 ( .A(n5379), .B(n5380), .Z(n5378) );
  NAND U9453 ( .A(n5380), .B(n5379), .Z(n5375) );
  IV U9454 ( .A(n5381), .Z(n5380) );
  NAND U9455 ( .A(n5382), .B(n5383), .Z(n5337) );
  NANDN U9456 ( .A(n5384), .B(n5385), .Z(n5383) );
  NAND U9457 ( .A(n5386), .B(n5387), .Z(n5385) );
  OR U9458 ( .A(n5387), .B(n5386), .Z(n5382) );
  IV U9459 ( .A(n5388), .Z(n5386) );
  XOR U9460 ( .A(n5363), .B(n5389), .Z(N29706) );
  XNOR U9461 ( .A(n5366), .B(n5365), .Z(n5389) );
  XNOR U9462 ( .A(n5377), .B(n5390), .Z(n5365) );
  XOR U9463 ( .A(n5381), .B(n5379), .Z(n5390) );
  XOR U9464 ( .A(n5387), .B(n5391), .Z(n5379) );
  XOR U9465 ( .A(n5384), .B(n5388), .Z(n5391) );
  NAND U9466 ( .A(n5392), .B(n5393), .Z(n5388) );
  NAND U9467 ( .A(n5394), .B(n5395), .Z(n5393) );
  NAND U9468 ( .A(n5396), .B(n5397), .Z(n5392) );
  AND U9469 ( .A(n5398), .B(n5399), .Z(n5384) );
  NAND U9470 ( .A(n5400), .B(n5401), .Z(n5399) );
  NAND U9471 ( .A(n5402), .B(n5403), .Z(n5398) );
  NANDN U9472 ( .A(n5404), .B(n5405), .Z(n5387) );
  NANDN U9473 ( .A(n5406), .B(n5407), .Z(n5381) );
  XNOR U9474 ( .A(n5372), .B(n5408), .Z(n5377) );
  XOR U9475 ( .A(n5370), .B(n5374), .Z(n5408) );
  NAND U9476 ( .A(n5409), .B(n5410), .Z(n5374) );
  NAND U9477 ( .A(n5411), .B(n5412), .Z(n5410) );
  NAND U9478 ( .A(n5413), .B(n5414), .Z(n5409) );
  AND U9479 ( .A(n5415), .B(n5416), .Z(n5370) );
  NAND U9480 ( .A(n5417), .B(n5418), .Z(n5416) );
  NAND U9481 ( .A(n5419), .B(n5420), .Z(n5415) );
  AND U9482 ( .A(n5421), .B(n5422), .Z(n5372) );
  NAND U9483 ( .A(n5423), .B(n5424), .Z(n5366) );
  XNOR U9484 ( .A(n5349), .B(n5425), .Z(n5363) );
  XOR U9485 ( .A(n5353), .B(n5351), .Z(n5425) );
  XOR U9486 ( .A(n5359), .B(n5426), .Z(n5351) );
  XOR U9487 ( .A(n5356), .B(n5360), .Z(n5426) );
  NAND U9488 ( .A(n5427), .B(n5428), .Z(n5360) );
  NAND U9489 ( .A(n5429), .B(n5430), .Z(n5428) );
  NAND U9490 ( .A(n5431), .B(n5432), .Z(n5427) );
  AND U9491 ( .A(n5433), .B(n5434), .Z(n5356) );
  NAND U9492 ( .A(n5435), .B(n5436), .Z(n5434) );
  NAND U9493 ( .A(n5437), .B(n5438), .Z(n5433) );
  NANDN U9494 ( .A(n5439), .B(n5440), .Z(n5359) );
  NANDN U9495 ( .A(n5441), .B(n5442), .Z(n5353) );
  XNOR U9496 ( .A(n5344), .B(n5443), .Z(n5349) );
  XOR U9497 ( .A(n5342), .B(n5346), .Z(n5443) );
  NAND U9498 ( .A(n5444), .B(n5445), .Z(n5346) );
  NAND U9499 ( .A(n5446), .B(n5447), .Z(n5445) );
  NAND U9500 ( .A(n5448), .B(n5449), .Z(n5444) );
  AND U9501 ( .A(n5450), .B(n5451), .Z(n5342) );
  NAND U9502 ( .A(n5452), .B(n5453), .Z(n5451) );
  NAND U9503 ( .A(n5454), .B(n5455), .Z(n5450) );
  AND U9504 ( .A(n5456), .B(n5457), .Z(n5344) );
  XOR U9505 ( .A(n5424), .B(n5423), .Z(N29705) );
  XNOR U9506 ( .A(n5442), .B(n5441), .Z(n5423) );
  XNOR U9507 ( .A(n5456), .B(n5457), .Z(n5441) );
  XOR U9508 ( .A(n5453), .B(n5452), .Z(n5457) );
  XOR U9509 ( .A(y[3555]), .B(x[3555]), .Z(n5452) );
  XOR U9510 ( .A(n5455), .B(n5454), .Z(n5453) );
  XOR U9511 ( .A(y[3557]), .B(x[3557]), .Z(n5454) );
  XOR U9512 ( .A(y[3556]), .B(x[3556]), .Z(n5455) );
  XOR U9513 ( .A(n5447), .B(n5446), .Z(n5456) );
  XOR U9514 ( .A(n5449), .B(n5448), .Z(n5446) );
  XOR U9515 ( .A(y[3554]), .B(x[3554]), .Z(n5448) );
  XOR U9516 ( .A(y[3553]), .B(x[3553]), .Z(n5449) );
  XOR U9517 ( .A(y[3552]), .B(x[3552]), .Z(n5447) );
  XNOR U9518 ( .A(n5440), .B(n5439), .Z(n5442) );
  XNOR U9519 ( .A(n5436), .B(n5435), .Z(n5439) );
  XOR U9520 ( .A(n5438), .B(n5437), .Z(n5435) );
  XOR U9521 ( .A(y[3551]), .B(x[3551]), .Z(n5437) );
  XOR U9522 ( .A(y[3550]), .B(x[3550]), .Z(n5438) );
  XOR U9523 ( .A(y[3549]), .B(x[3549]), .Z(n5436) );
  XOR U9524 ( .A(n5430), .B(n5429), .Z(n5440) );
  XOR U9525 ( .A(n5432), .B(n5431), .Z(n5429) );
  XOR U9526 ( .A(y[3548]), .B(x[3548]), .Z(n5431) );
  XOR U9527 ( .A(y[3547]), .B(x[3547]), .Z(n5432) );
  XOR U9528 ( .A(y[3546]), .B(x[3546]), .Z(n5430) );
  XNOR U9529 ( .A(n5407), .B(n5406), .Z(n5424) );
  XNOR U9530 ( .A(n5421), .B(n5422), .Z(n5406) );
  XOR U9531 ( .A(n5418), .B(n5417), .Z(n5422) );
  XOR U9532 ( .A(y[3543]), .B(x[3543]), .Z(n5417) );
  XOR U9533 ( .A(n5420), .B(n5419), .Z(n5418) );
  XOR U9534 ( .A(y[3545]), .B(x[3545]), .Z(n5419) );
  XOR U9535 ( .A(y[3544]), .B(x[3544]), .Z(n5420) );
  XOR U9536 ( .A(n5412), .B(n5411), .Z(n5421) );
  XOR U9537 ( .A(n5414), .B(n5413), .Z(n5411) );
  XOR U9538 ( .A(y[3542]), .B(x[3542]), .Z(n5413) );
  XOR U9539 ( .A(y[3541]), .B(x[3541]), .Z(n5414) );
  XOR U9540 ( .A(y[3540]), .B(x[3540]), .Z(n5412) );
  XNOR U9541 ( .A(n5405), .B(n5404), .Z(n5407) );
  XNOR U9542 ( .A(n5401), .B(n5400), .Z(n5404) );
  XOR U9543 ( .A(n5403), .B(n5402), .Z(n5400) );
  XOR U9544 ( .A(y[3539]), .B(x[3539]), .Z(n5402) );
  XOR U9545 ( .A(y[3538]), .B(x[3538]), .Z(n5403) );
  XOR U9546 ( .A(y[3537]), .B(x[3537]), .Z(n5401) );
  XOR U9547 ( .A(n5395), .B(n5394), .Z(n5405) );
  XOR U9548 ( .A(n5397), .B(n5396), .Z(n5394) );
  XOR U9549 ( .A(y[3536]), .B(x[3536]), .Z(n5396) );
  XOR U9550 ( .A(y[3535]), .B(x[3535]), .Z(n5397) );
  XOR U9551 ( .A(y[3534]), .B(x[3534]), .Z(n5395) );
  NAND U9552 ( .A(n5458), .B(n5459), .Z(N29697) );
  NAND U9553 ( .A(n5460), .B(n5461), .Z(n5459) );
  NANDN U9554 ( .A(n5462), .B(n5463), .Z(n5461) );
  NANDN U9555 ( .A(n5463), .B(n5462), .Z(n5458) );
  XOR U9556 ( .A(n5462), .B(n5464), .Z(N29696) );
  XNOR U9557 ( .A(n5460), .B(n5463), .Z(n5464) );
  NAND U9558 ( .A(n5465), .B(n5466), .Z(n5463) );
  NAND U9559 ( .A(n5467), .B(n5468), .Z(n5466) );
  NANDN U9560 ( .A(n5469), .B(n5470), .Z(n5468) );
  NANDN U9561 ( .A(n5470), .B(n5469), .Z(n5465) );
  AND U9562 ( .A(n5471), .B(n5472), .Z(n5460) );
  NAND U9563 ( .A(n5473), .B(n5474), .Z(n5472) );
  OR U9564 ( .A(n5475), .B(n5476), .Z(n5474) );
  NAND U9565 ( .A(n5476), .B(n5475), .Z(n5471) );
  IV U9566 ( .A(n5477), .Z(n5476) );
  AND U9567 ( .A(n5478), .B(n5479), .Z(n5462) );
  NAND U9568 ( .A(n5480), .B(n5481), .Z(n5479) );
  NANDN U9569 ( .A(n5482), .B(n5483), .Z(n5481) );
  NANDN U9570 ( .A(n5483), .B(n5482), .Z(n5478) );
  XOR U9571 ( .A(n5475), .B(n5484), .Z(N29695) );
  XOR U9572 ( .A(n5473), .B(n5477), .Z(n5484) );
  XNOR U9573 ( .A(n5470), .B(n5485), .Z(n5477) );
  XNOR U9574 ( .A(n5467), .B(n5469), .Z(n5485) );
  AND U9575 ( .A(n5486), .B(n5487), .Z(n5469) );
  NANDN U9576 ( .A(n5488), .B(n5489), .Z(n5487) );
  NANDN U9577 ( .A(n5490), .B(n5491), .Z(n5489) );
  IV U9578 ( .A(n5492), .Z(n5491) );
  NAND U9579 ( .A(n5492), .B(n5490), .Z(n5486) );
  AND U9580 ( .A(n5493), .B(n5494), .Z(n5467) );
  NAND U9581 ( .A(n5495), .B(n5496), .Z(n5494) );
  OR U9582 ( .A(n5497), .B(n5498), .Z(n5496) );
  NAND U9583 ( .A(n5498), .B(n5497), .Z(n5493) );
  IV U9584 ( .A(n5499), .Z(n5498) );
  NAND U9585 ( .A(n5500), .B(n5501), .Z(n5470) );
  NANDN U9586 ( .A(n5502), .B(n5503), .Z(n5501) );
  NAND U9587 ( .A(n5504), .B(n5505), .Z(n5503) );
  OR U9588 ( .A(n5505), .B(n5504), .Z(n5500) );
  IV U9589 ( .A(n5506), .Z(n5504) );
  AND U9590 ( .A(n5507), .B(n5508), .Z(n5473) );
  NAND U9591 ( .A(n5509), .B(n5510), .Z(n5508) );
  NANDN U9592 ( .A(n5511), .B(n5512), .Z(n5510) );
  NANDN U9593 ( .A(n5512), .B(n5511), .Z(n5507) );
  XOR U9594 ( .A(n5483), .B(n5513), .Z(n5475) );
  XNOR U9595 ( .A(n5480), .B(n5482), .Z(n5513) );
  AND U9596 ( .A(n5514), .B(n5515), .Z(n5482) );
  NANDN U9597 ( .A(n5516), .B(n5517), .Z(n5515) );
  NANDN U9598 ( .A(n5518), .B(n5519), .Z(n5517) );
  IV U9599 ( .A(n5520), .Z(n5519) );
  NAND U9600 ( .A(n5520), .B(n5518), .Z(n5514) );
  AND U9601 ( .A(n5521), .B(n5522), .Z(n5480) );
  NAND U9602 ( .A(n5523), .B(n5524), .Z(n5522) );
  OR U9603 ( .A(n5525), .B(n5526), .Z(n5524) );
  NAND U9604 ( .A(n5526), .B(n5525), .Z(n5521) );
  IV U9605 ( .A(n5527), .Z(n5526) );
  NAND U9606 ( .A(n5528), .B(n5529), .Z(n5483) );
  NANDN U9607 ( .A(n5530), .B(n5531), .Z(n5529) );
  NAND U9608 ( .A(n5532), .B(n5533), .Z(n5531) );
  OR U9609 ( .A(n5533), .B(n5532), .Z(n5528) );
  IV U9610 ( .A(n5534), .Z(n5532) );
  XOR U9611 ( .A(n5509), .B(n5535), .Z(N29694) );
  XNOR U9612 ( .A(n5512), .B(n5511), .Z(n5535) );
  XNOR U9613 ( .A(n5523), .B(n5536), .Z(n5511) );
  XOR U9614 ( .A(n5527), .B(n5525), .Z(n5536) );
  XOR U9615 ( .A(n5533), .B(n5537), .Z(n5525) );
  XOR U9616 ( .A(n5530), .B(n5534), .Z(n5537) );
  NAND U9617 ( .A(n5538), .B(n5539), .Z(n5534) );
  NAND U9618 ( .A(n5540), .B(n5541), .Z(n5539) );
  NAND U9619 ( .A(n5542), .B(n5543), .Z(n5538) );
  AND U9620 ( .A(n5544), .B(n5545), .Z(n5530) );
  NAND U9621 ( .A(n5546), .B(n5547), .Z(n5545) );
  NAND U9622 ( .A(n5548), .B(n5549), .Z(n5544) );
  NANDN U9623 ( .A(n5550), .B(n5551), .Z(n5533) );
  NANDN U9624 ( .A(n5552), .B(n5553), .Z(n5527) );
  XNOR U9625 ( .A(n5518), .B(n5554), .Z(n5523) );
  XOR U9626 ( .A(n5516), .B(n5520), .Z(n5554) );
  NAND U9627 ( .A(n5555), .B(n5556), .Z(n5520) );
  NAND U9628 ( .A(n5557), .B(n5558), .Z(n5556) );
  NAND U9629 ( .A(n5559), .B(n5560), .Z(n5555) );
  AND U9630 ( .A(n5561), .B(n5562), .Z(n5516) );
  NAND U9631 ( .A(n5563), .B(n5564), .Z(n5562) );
  NAND U9632 ( .A(n5565), .B(n5566), .Z(n5561) );
  AND U9633 ( .A(n5567), .B(n5568), .Z(n5518) );
  NAND U9634 ( .A(n5569), .B(n5570), .Z(n5512) );
  XNOR U9635 ( .A(n5495), .B(n5571), .Z(n5509) );
  XOR U9636 ( .A(n5499), .B(n5497), .Z(n5571) );
  XOR U9637 ( .A(n5505), .B(n5572), .Z(n5497) );
  XOR U9638 ( .A(n5502), .B(n5506), .Z(n5572) );
  NAND U9639 ( .A(n5573), .B(n5574), .Z(n5506) );
  NAND U9640 ( .A(n5575), .B(n5576), .Z(n5574) );
  NAND U9641 ( .A(n5577), .B(n5578), .Z(n5573) );
  AND U9642 ( .A(n5579), .B(n5580), .Z(n5502) );
  NAND U9643 ( .A(n5581), .B(n5582), .Z(n5580) );
  NAND U9644 ( .A(n5583), .B(n5584), .Z(n5579) );
  NANDN U9645 ( .A(n5585), .B(n5586), .Z(n5505) );
  NANDN U9646 ( .A(n5587), .B(n5588), .Z(n5499) );
  XNOR U9647 ( .A(n5490), .B(n5589), .Z(n5495) );
  XOR U9648 ( .A(n5488), .B(n5492), .Z(n5589) );
  NAND U9649 ( .A(n5590), .B(n5591), .Z(n5492) );
  NAND U9650 ( .A(n5592), .B(n5593), .Z(n5591) );
  NAND U9651 ( .A(n5594), .B(n5595), .Z(n5590) );
  AND U9652 ( .A(n5596), .B(n5597), .Z(n5488) );
  NAND U9653 ( .A(n5598), .B(n5599), .Z(n5597) );
  NAND U9654 ( .A(n5600), .B(n5601), .Z(n5596) );
  AND U9655 ( .A(n5602), .B(n5603), .Z(n5490) );
  XOR U9656 ( .A(n5570), .B(n5569), .Z(N29693) );
  XNOR U9657 ( .A(n5588), .B(n5587), .Z(n5569) );
  XNOR U9658 ( .A(n5602), .B(n5603), .Z(n5587) );
  XOR U9659 ( .A(n5599), .B(n5598), .Z(n5603) );
  XOR U9660 ( .A(y[3531]), .B(x[3531]), .Z(n5598) );
  XOR U9661 ( .A(n5601), .B(n5600), .Z(n5599) );
  XOR U9662 ( .A(y[3533]), .B(x[3533]), .Z(n5600) );
  XOR U9663 ( .A(y[3532]), .B(x[3532]), .Z(n5601) );
  XOR U9664 ( .A(n5593), .B(n5592), .Z(n5602) );
  XOR U9665 ( .A(n5595), .B(n5594), .Z(n5592) );
  XOR U9666 ( .A(y[3530]), .B(x[3530]), .Z(n5594) );
  XOR U9667 ( .A(y[3529]), .B(x[3529]), .Z(n5595) );
  XOR U9668 ( .A(y[3528]), .B(x[3528]), .Z(n5593) );
  XNOR U9669 ( .A(n5586), .B(n5585), .Z(n5588) );
  XNOR U9670 ( .A(n5582), .B(n5581), .Z(n5585) );
  XOR U9671 ( .A(n5584), .B(n5583), .Z(n5581) );
  XOR U9672 ( .A(y[3527]), .B(x[3527]), .Z(n5583) );
  XOR U9673 ( .A(y[3526]), .B(x[3526]), .Z(n5584) );
  XOR U9674 ( .A(y[3525]), .B(x[3525]), .Z(n5582) );
  XOR U9675 ( .A(n5576), .B(n5575), .Z(n5586) );
  XOR U9676 ( .A(n5578), .B(n5577), .Z(n5575) );
  XOR U9677 ( .A(y[3524]), .B(x[3524]), .Z(n5577) );
  XOR U9678 ( .A(y[3523]), .B(x[3523]), .Z(n5578) );
  XOR U9679 ( .A(y[3522]), .B(x[3522]), .Z(n5576) );
  XNOR U9680 ( .A(n5553), .B(n5552), .Z(n5570) );
  XNOR U9681 ( .A(n5567), .B(n5568), .Z(n5552) );
  XOR U9682 ( .A(n5564), .B(n5563), .Z(n5568) );
  XOR U9683 ( .A(y[3519]), .B(x[3519]), .Z(n5563) );
  XOR U9684 ( .A(n5566), .B(n5565), .Z(n5564) );
  XOR U9685 ( .A(y[3521]), .B(x[3521]), .Z(n5565) );
  XOR U9686 ( .A(y[3520]), .B(x[3520]), .Z(n5566) );
  XOR U9687 ( .A(n5558), .B(n5557), .Z(n5567) );
  XOR U9688 ( .A(n5560), .B(n5559), .Z(n5557) );
  XOR U9689 ( .A(y[3518]), .B(x[3518]), .Z(n5559) );
  XOR U9690 ( .A(y[3517]), .B(x[3517]), .Z(n5560) );
  XOR U9691 ( .A(y[3516]), .B(x[3516]), .Z(n5558) );
  XNOR U9692 ( .A(n5551), .B(n5550), .Z(n5553) );
  XNOR U9693 ( .A(n5547), .B(n5546), .Z(n5550) );
  XOR U9694 ( .A(n5549), .B(n5548), .Z(n5546) );
  XOR U9695 ( .A(y[3515]), .B(x[3515]), .Z(n5548) );
  XOR U9696 ( .A(y[3514]), .B(x[3514]), .Z(n5549) );
  XOR U9697 ( .A(y[3513]), .B(x[3513]), .Z(n5547) );
  XOR U9698 ( .A(n5541), .B(n5540), .Z(n5551) );
  XOR U9699 ( .A(n5543), .B(n5542), .Z(n5540) );
  XOR U9700 ( .A(y[3512]), .B(x[3512]), .Z(n5542) );
  XOR U9701 ( .A(y[3511]), .B(x[3511]), .Z(n5543) );
  XOR U9702 ( .A(y[3510]), .B(x[3510]), .Z(n5541) );
  NAND U9703 ( .A(n5604), .B(n5605), .Z(N29685) );
  NAND U9704 ( .A(n5606), .B(n5607), .Z(n5605) );
  NANDN U9705 ( .A(n5608), .B(n5609), .Z(n5607) );
  NANDN U9706 ( .A(n5609), .B(n5608), .Z(n5604) );
  XOR U9707 ( .A(n5608), .B(n5610), .Z(N29684) );
  XNOR U9708 ( .A(n5606), .B(n5609), .Z(n5610) );
  NAND U9709 ( .A(n5611), .B(n5612), .Z(n5609) );
  NAND U9710 ( .A(n5613), .B(n5614), .Z(n5612) );
  NANDN U9711 ( .A(n5615), .B(n5616), .Z(n5614) );
  NANDN U9712 ( .A(n5616), .B(n5615), .Z(n5611) );
  AND U9713 ( .A(n5617), .B(n5618), .Z(n5606) );
  NAND U9714 ( .A(n5619), .B(n5620), .Z(n5618) );
  OR U9715 ( .A(n5621), .B(n5622), .Z(n5620) );
  NAND U9716 ( .A(n5622), .B(n5621), .Z(n5617) );
  IV U9717 ( .A(n5623), .Z(n5622) );
  AND U9718 ( .A(n5624), .B(n5625), .Z(n5608) );
  NAND U9719 ( .A(n5626), .B(n5627), .Z(n5625) );
  NANDN U9720 ( .A(n5628), .B(n5629), .Z(n5627) );
  NANDN U9721 ( .A(n5629), .B(n5628), .Z(n5624) );
  XOR U9722 ( .A(n5621), .B(n5630), .Z(N29683) );
  XOR U9723 ( .A(n5619), .B(n5623), .Z(n5630) );
  XNOR U9724 ( .A(n5616), .B(n5631), .Z(n5623) );
  XNOR U9725 ( .A(n5613), .B(n5615), .Z(n5631) );
  AND U9726 ( .A(n5632), .B(n5633), .Z(n5615) );
  NANDN U9727 ( .A(n5634), .B(n5635), .Z(n5633) );
  NANDN U9728 ( .A(n5636), .B(n5637), .Z(n5635) );
  IV U9729 ( .A(n5638), .Z(n5637) );
  NAND U9730 ( .A(n5638), .B(n5636), .Z(n5632) );
  AND U9731 ( .A(n5639), .B(n5640), .Z(n5613) );
  NAND U9732 ( .A(n5641), .B(n5642), .Z(n5640) );
  OR U9733 ( .A(n5643), .B(n5644), .Z(n5642) );
  NAND U9734 ( .A(n5644), .B(n5643), .Z(n5639) );
  IV U9735 ( .A(n5645), .Z(n5644) );
  NAND U9736 ( .A(n5646), .B(n5647), .Z(n5616) );
  NANDN U9737 ( .A(n5648), .B(n5649), .Z(n5647) );
  NAND U9738 ( .A(n5650), .B(n5651), .Z(n5649) );
  OR U9739 ( .A(n5651), .B(n5650), .Z(n5646) );
  IV U9740 ( .A(n5652), .Z(n5650) );
  AND U9741 ( .A(n5653), .B(n5654), .Z(n5619) );
  NAND U9742 ( .A(n5655), .B(n5656), .Z(n5654) );
  NANDN U9743 ( .A(n5657), .B(n5658), .Z(n5656) );
  NANDN U9744 ( .A(n5658), .B(n5657), .Z(n5653) );
  XOR U9745 ( .A(n5629), .B(n5659), .Z(n5621) );
  XNOR U9746 ( .A(n5626), .B(n5628), .Z(n5659) );
  AND U9747 ( .A(n5660), .B(n5661), .Z(n5628) );
  NANDN U9748 ( .A(n5662), .B(n5663), .Z(n5661) );
  NANDN U9749 ( .A(n5664), .B(n5665), .Z(n5663) );
  IV U9750 ( .A(n5666), .Z(n5665) );
  NAND U9751 ( .A(n5666), .B(n5664), .Z(n5660) );
  AND U9752 ( .A(n5667), .B(n5668), .Z(n5626) );
  NAND U9753 ( .A(n5669), .B(n5670), .Z(n5668) );
  OR U9754 ( .A(n5671), .B(n5672), .Z(n5670) );
  NAND U9755 ( .A(n5672), .B(n5671), .Z(n5667) );
  IV U9756 ( .A(n5673), .Z(n5672) );
  NAND U9757 ( .A(n5674), .B(n5675), .Z(n5629) );
  NANDN U9758 ( .A(n5676), .B(n5677), .Z(n5675) );
  NAND U9759 ( .A(n5678), .B(n5679), .Z(n5677) );
  OR U9760 ( .A(n5679), .B(n5678), .Z(n5674) );
  IV U9761 ( .A(n5680), .Z(n5678) );
  XOR U9762 ( .A(n5655), .B(n5681), .Z(N29682) );
  XNOR U9763 ( .A(n5658), .B(n5657), .Z(n5681) );
  XNOR U9764 ( .A(n5669), .B(n5682), .Z(n5657) );
  XOR U9765 ( .A(n5673), .B(n5671), .Z(n5682) );
  XOR U9766 ( .A(n5679), .B(n5683), .Z(n5671) );
  XOR U9767 ( .A(n5676), .B(n5680), .Z(n5683) );
  NAND U9768 ( .A(n5684), .B(n5685), .Z(n5680) );
  NAND U9769 ( .A(n5686), .B(n5687), .Z(n5685) );
  NAND U9770 ( .A(n5688), .B(n5689), .Z(n5684) );
  AND U9771 ( .A(n5690), .B(n5691), .Z(n5676) );
  NAND U9772 ( .A(n5692), .B(n5693), .Z(n5691) );
  NAND U9773 ( .A(n5694), .B(n5695), .Z(n5690) );
  NANDN U9774 ( .A(n5696), .B(n5697), .Z(n5679) );
  NANDN U9775 ( .A(n5698), .B(n5699), .Z(n5673) );
  XNOR U9776 ( .A(n5664), .B(n5700), .Z(n5669) );
  XOR U9777 ( .A(n5662), .B(n5666), .Z(n5700) );
  NAND U9778 ( .A(n5701), .B(n5702), .Z(n5666) );
  NAND U9779 ( .A(n5703), .B(n5704), .Z(n5702) );
  NAND U9780 ( .A(n5705), .B(n5706), .Z(n5701) );
  AND U9781 ( .A(n5707), .B(n5708), .Z(n5662) );
  NAND U9782 ( .A(n5709), .B(n5710), .Z(n5708) );
  NAND U9783 ( .A(n5711), .B(n5712), .Z(n5707) );
  AND U9784 ( .A(n5713), .B(n5714), .Z(n5664) );
  NAND U9785 ( .A(n5715), .B(n5716), .Z(n5658) );
  XNOR U9786 ( .A(n5641), .B(n5717), .Z(n5655) );
  XOR U9787 ( .A(n5645), .B(n5643), .Z(n5717) );
  XOR U9788 ( .A(n5651), .B(n5718), .Z(n5643) );
  XOR U9789 ( .A(n5648), .B(n5652), .Z(n5718) );
  NAND U9790 ( .A(n5719), .B(n5720), .Z(n5652) );
  NAND U9791 ( .A(n5721), .B(n5722), .Z(n5720) );
  NAND U9792 ( .A(n5723), .B(n5724), .Z(n5719) );
  AND U9793 ( .A(n5725), .B(n5726), .Z(n5648) );
  NAND U9794 ( .A(n5727), .B(n5728), .Z(n5726) );
  NAND U9795 ( .A(n5729), .B(n5730), .Z(n5725) );
  NANDN U9796 ( .A(n5731), .B(n5732), .Z(n5651) );
  NANDN U9797 ( .A(n5733), .B(n5734), .Z(n5645) );
  XNOR U9798 ( .A(n5636), .B(n5735), .Z(n5641) );
  XOR U9799 ( .A(n5634), .B(n5638), .Z(n5735) );
  NAND U9800 ( .A(n5736), .B(n5737), .Z(n5638) );
  NAND U9801 ( .A(n5738), .B(n5739), .Z(n5737) );
  NAND U9802 ( .A(n5740), .B(n5741), .Z(n5736) );
  AND U9803 ( .A(n5742), .B(n5743), .Z(n5634) );
  NAND U9804 ( .A(n5744), .B(n5745), .Z(n5743) );
  NAND U9805 ( .A(n5746), .B(n5747), .Z(n5742) );
  AND U9806 ( .A(n5748), .B(n5749), .Z(n5636) );
  XOR U9807 ( .A(n5716), .B(n5715), .Z(N29681) );
  XNOR U9808 ( .A(n5734), .B(n5733), .Z(n5715) );
  XNOR U9809 ( .A(n5748), .B(n5749), .Z(n5733) );
  XOR U9810 ( .A(n5745), .B(n5744), .Z(n5749) );
  XOR U9811 ( .A(y[3507]), .B(x[3507]), .Z(n5744) );
  XOR U9812 ( .A(n5747), .B(n5746), .Z(n5745) );
  XOR U9813 ( .A(y[3509]), .B(x[3509]), .Z(n5746) );
  XOR U9814 ( .A(y[3508]), .B(x[3508]), .Z(n5747) );
  XOR U9815 ( .A(n5739), .B(n5738), .Z(n5748) );
  XOR U9816 ( .A(n5741), .B(n5740), .Z(n5738) );
  XOR U9817 ( .A(y[3506]), .B(x[3506]), .Z(n5740) );
  XOR U9818 ( .A(y[3505]), .B(x[3505]), .Z(n5741) );
  XOR U9819 ( .A(y[3504]), .B(x[3504]), .Z(n5739) );
  XNOR U9820 ( .A(n5732), .B(n5731), .Z(n5734) );
  XNOR U9821 ( .A(n5728), .B(n5727), .Z(n5731) );
  XOR U9822 ( .A(n5730), .B(n5729), .Z(n5727) );
  XOR U9823 ( .A(y[3503]), .B(x[3503]), .Z(n5729) );
  XOR U9824 ( .A(y[3502]), .B(x[3502]), .Z(n5730) );
  XOR U9825 ( .A(y[3501]), .B(x[3501]), .Z(n5728) );
  XOR U9826 ( .A(n5722), .B(n5721), .Z(n5732) );
  XOR U9827 ( .A(n5724), .B(n5723), .Z(n5721) );
  XOR U9828 ( .A(y[3500]), .B(x[3500]), .Z(n5723) );
  XOR U9829 ( .A(y[3499]), .B(x[3499]), .Z(n5724) );
  XOR U9830 ( .A(y[3498]), .B(x[3498]), .Z(n5722) );
  XNOR U9831 ( .A(n5699), .B(n5698), .Z(n5716) );
  XNOR U9832 ( .A(n5713), .B(n5714), .Z(n5698) );
  XOR U9833 ( .A(n5710), .B(n5709), .Z(n5714) );
  XOR U9834 ( .A(y[3495]), .B(x[3495]), .Z(n5709) );
  XOR U9835 ( .A(n5712), .B(n5711), .Z(n5710) );
  XOR U9836 ( .A(y[3497]), .B(x[3497]), .Z(n5711) );
  XOR U9837 ( .A(y[3496]), .B(x[3496]), .Z(n5712) );
  XOR U9838 ( .A(n5704), .B(n5703), .Z(n5713) );
  XOR U9839 ( .A(n5706), .B(n5705), .Z(n5703) );
  XOR U9840 ( .A(y[3494]), .B(x[3494]), .Z(n5705) );
  XOR U9841 ( .A(y[3493]), .B(x[3493]), .Z(n5706) );
  XOR U9842 ( .A(y[3492]), .B(x[3492]), .Z(n5704) );
  XNOR U9843 ( .A(n5697), .B(n5696), .Z(n5699) );
  XNOR U9844 ( .A(n5693), .B(n5692), .Z(n5696) );
  XOR U9845 ( .A(n5695), .B(n5694), .Z(n5692) );
  XOR U9846 ( .A(y[3491]), .B(x[3491]), .Z(n5694) );
  XOR U9847 ( .A(y[3490]), .B(x[3490]), .Z(n5695) );
  XOR U9848 ( .A(y[3489]), .B(x[3489]), .Z(n5693) );
  XOR U9849 ( .A(n5687), .B(n5686), .Z(n5697) );
  XOR U9850 ( .A(n5689), .B(n5688), .Z(n5686) );
  XOR U9851 ( .A(y[3488]), .B(x[3488]), .Z(n5688) );
  XOR U9852 ( .A(y[3487]), .B(x[3487]), .Z(n5689) );
  XOR U9853 ( .A(y[3486]), .B(x[3486]), .Z(n5687) );
  NAND U9854 ( .A(n5750), .B(n5751), .Z(N29673) );
  NAND U9855 ( .A(n5752), .B(n5753), .Z(n5751) );
  NANDN U9856 ( .A(n5754), .B(n5755), .Z(n5753) );
  NANDN U9857 ( .A(n5755), .B(n5754), .Z(n5750) );
  XOR U9858 ( .A(n5754), .B(n5756), .Z(N29672) );
  XNOR U9859 ( .A(n5752), .B(n5755), .Z(n5756) );
  NAND U9860 ( .A(n5757), .B(n5758), .Z(n5755) );
  NAND U9861 ( .A(n5759), .B(n5760), .Z(n5758) );
  NANDN U9862 ( .A(n5761), .B(n5762), .Z(n5760) );
  NANDN U9863 ( .A(n5762), .B(n5761), .Z(n5757) );
  AND U9864 ( .A(n5763), .B(n5764), .Z(n5752) );
  NAND U9865 ( .A(n5765), .B(n5766), .Z(n5764) );
  OR U9866 ( .A(n5767), .B(n5768), .Z(n5766) );
  NAND U9867 ( .A(n5768), .B(n5767), .Z(n5763) );
  IV U9868 ( .A(n5769), .Z(n5768) );
  AND U9869 ( .A(n5770), .B(n5771), .Z(n5754) );
  NAND U9870 ( .A(n5772), .B(n5773), .Z(n5771) );
  NANDN U9871 ( .A(n5774), .B(n5775), .Z(n5773) );
  NANDN U9872 ( .A(n5775), .B(n5774), .Z(n5770) );
  XOR U9873 ( .A(n5767), .B(n5776), .Z(N29671) );
  XOR U9874 ( .A(n5765), .B(n5769), .Z(n5776) );
  XNOR U9875 ( .A(n5762), .B(n5777), .Z(n5769) );
  XNOR U9876 ( .A(n5759), .B(n5761), .Z(n5777) );
  AND U9877 ( .A(n5778), .B(n5779), .Z(n5761) );
  NANDN U9878 ( .A(n5780), .B(n5781), .Z(n5779) );
  NANDN U9879 ( .A(n5782), .B(n5783), .Z(n5781) );
  IV U9880 ( .A(n5784), .Z(n5783) );
  NAND U9881 ( .A(n5784), .B(n5782), .Z(n5778) );
  AND U9882 ( .A(n5785), .B(n5786), .Z(n5759) );
  NAND U9883 ( .A(n5787), .B(n5788), .Z(n5786) );
  OR U9884 ( .A(n5789), .B(n5790), .Z(n5788) );
  NAND U9885 ( .A(n5790), .B(n5789), .Z(n5785) );
  IV U9886 ( .A(n5791), .Z(n5790) );
  NAND U9887 ( .A(n5792), .B(n5793), .Z(n5762) );
  NANDN U9888 ( .A(n5794), .B(n5795), .Z(n5793) );
  NAND U9889 ( .A(n5796), .B(n5797), .Z(n5795) );
  OR U9890 ( .A(n5797), .B(n5796), .Z(n5792) );
  IV U9891 ( .A(n5798), .Z(n5796) );
  AND U9892 ( .A(n5799), .B(n5800), .Z(n5765) );
  NAND U9893 ( .A(n5801), .B(n5802), .Z(n5800) );
  NANDN U9894 ( .A(n5803), .B(n5804), .Z(n5802) );
  NANDN U9895 ( .A(n5804), .B(n5803), .Z(n5799) );
  XOR U9896 ( .A(n5775), .B(n5805), .Z(n5767) );
  XNOR U9897 ( .A(n5772), .B(n5774), .Z(n5805) );
  AND U9898 ( .A(n5806), .B(n5807), .Z(n5774) );
  NANDN U9899 ( .A(n5808), .B(n5809), .Z(n5807) );
  NANDN U9900 ( .A(n5810), .B(n5811), .Z(n5809) );
  IV U9901 ( .A(n5812), .Z(n5811) );
  NAND U9902 ( .A(n5812), .B(n5810), .Z(n5806) );
  AND U9903 ( .A(n5813), .B(n5814), .Z(n5772) );
  NAND U9904 ( .A(n5815), .B(n5816), .Z(n5814) );
  OR U9905 ( .A(n5817), .B(n5818), .Z(n5816) );
  NAND U9906 ( .A(n5818), .B(n5817), .Z(n5813) );
  IV U9907 ( .A(n5819), .Z(n5818) );
  NAND U9908 ( .A(n5820), .B(n5821), .Z(n5775) );
  NANDN U9909 ( .A(n5822), .B(n5823), .Z(n5821) );
  NAND U9910 ( .A(n5824), .B(n5825), .Z(n5823) );
  OR U9911 ( .A(n5825), .B(n5824), .Z(n5820) );
  IV U9912 ( .A(n5826), .Z(n5824) );
  XOR U9913 ( .A(n5801), .B(n5827), .Z(N29670) );
  XNOR U9914 ( .A(n5804), .B(n5803), .Z(n5827) );
  XNOR U9915 ( .A(n5815), .B(n5828), .Z(n5803) );
  XOR U9916 ( .A(n5819), .B(n5817), .Z(n5828) );
  XOR U9917 ( .A(n5825), .B(n5829), .Z(n5817) );
  XOR U9918 ( .A(n5822), .B(n5826), .Z(n5829) );
  NAND U9919 ( .A(n5830), .B(n5831), .Z(n5826) );
  NAND U9920 ( .A(n5832), .B(n5833), .Z(n5831) );
  NAND U9921 ( .A(n5834), .B(n5835), .Z(n5830) );
  AND U9922 ( .A(n5836), .B(n5837), .Z(n5822) );
  NAND U9923 ( .A(n5838), .B(n5839), .Z(n5837) );
  NAND U9924 ( .A(n5840), .B(n5841), .Z(n5836) );
  NANDN U9925 ( .A(n5842), .B(n5843), .Z(n5825) );
  NANDN U9926 ( .A(n5844), .B(n5845), .Z(n5819) );
  XNOR U9927 ( .A(n5810), .B(n5846), .Z(n5815) );
  XOR U9928 ( .A(n5808), .B(n5812), .Z(n5846) );
  NAND U9929 ( .A(n5847), .B(n5848), .Z(n5812) );
  NAND U9930 ( .A(n5849), .B(n5850), .Z(n5848) );
  NAND U9931 ( .A(n5851), .B(n5852), .Z(n5847) );
  AND U9932 ( .A(n5853), .B(n5854), .Z(n5808) );
  NAND U9933 ( .A(n5855), .B(n5856), .Z(n5854) );
  NAND U9934 ( .A(n5857), .B(n5858), .Z(n5853) );
  AND U9935 ( .A(n5859), .B(n5860), .Z(n5810) );
  NAND U9936 ( .A(n5861), .B(n5862), .Z(n5804) );
  XNOR U9937 ( .A(n5787), .B(n5863), .Z(n5801) );
  XOR U9938 ( .A(n5791), .B(n5789), .Z(n5863) );
  XOR U9939 ( .A(n5797), .B(n5864), .Z(n5789) );
  XOR U9940 ( .A(n5794), .B(n5798), .Z(n5864) );
  NAND U9941 ( .A(n5865), .B(n5866), .Z(n5798) );
  NAND U9942 ( .A(n5867), .B(n5868), .Z(n5866) );
  NAND U9943 ( .A(n5869), .B(n5870), .Z(n5865) );
  AND U9944 ( .A(n5871), .B(n5872), .Z(n5794) );
  NAND U9945 ( .A(n5873), .B(n5874), .Z(n5872) );
  NAND U9946 ( .A(n5875), .B(n5876), .Z(n5871) );
  NANDN U9947 ( .A(n5877), .B(n5878), .Z(n5797) );
  NANDN U9948 ( .A(n5879), .B(n5880), .Z(n5791) );
  XNOR U9949 ( .A(n5782), .B(n5881), .Z(n5787) );
  XOR U9950 ( .A(n5780), .B(n5784), .Z(n5881) );
  NAND U9951 ( .A(n5882), .B(n5883), .Z(n5784) );
  NAND U9952 ( .A(n5884), .B(n5885), .Z(n5883) );
  NAND U9953 ( .A(n5886), .B(n5887), .Z(n5882) );
  AND U9954 ( .A(n5888), .B(n5889), .Z(n5780) );
  NAND U9955 ( .A(n5890), .B(n5891), .Z(n5889) );
  NAND U9956 ( .A(n5892), .B(n5893), .Z(n5888) );
  AND U9957 ( .A(n5894), .B(n5895), .Z(n5782) );
  XOR U9958 ( .A(n5862), .B(n5861), .Z(N29669) );
  XNOR U9959 ( .A(n5880), .B(n5879), .Z(n5861) );
  XNOR U9960 ( .A(n5894), .B(n5895), .Z(n5879) );
  XOR U9961 ( .A(n5891), .B(n5890), .Z(n5895) );
  XOR U9962 ( .A(y[3483]), .B(x[3483]), .Z(n5890) );
  XOR U9963 ( .A(n5893), .B(n5892), .Z(n5891) );
  XOR U9964 ( .A(y[3485]), .B(x[3485]), .Z(n5892) );
  XOR U9965 ( .A(y[3484]), .B(x[3484]), .Z(n5893) );
  XOR U9966 ( .A(n5885), .B(n5884), .Z(n5894) );
  XOR U9967 ( .A(n5887), .B(n5886), .Z(n5884) );
  XOR U9968 ( .A(y[3482]), .B(x[3482]), .Z(n5886) );
  XOR U9969 ( .A(y[3481]), .B(x[3481]), .Z(n5887) );
  XOR U9970 ( .A(y[3480]), .B(x[3480]), .Z(n5885) );
  XNOR U9971 ( .A(n5878), .B(n5877), .Z(n5880) );
  XNOR U9972 ( .A(n5874), .B(n5873), .Z(n5877) );
  XOR U9973 ( .A(n5876), .B(n5875), .Z(n5873) );
  XOR U9974 ( .A(y[3479]), .B(x[3479]), .Z(n5875) );
  XOR U9975 ( .A(y[3478]), .B(x[3478]), .Z(n5876) );
  XOR U9976 ( .A(y[3477]), .B(x[3477]), .Z(n5874) );
  XOR U9977 ( .A(n5868), .B(n5867), .Z(n5878) );
  XOR U9978 ( .A(n5870), .B(n5869), .Z(n5867) );
  XOR U9979 ( .A(y[3476]), .B(x[3476]), .Z(n5869) );
  XOR U9980 ( .A(y[3475]), .B(x[3475]), .Z(n5870) );
  XOR U9981 ( .A(y[3474]), .B(x[3474]), .Z(n5868) );
  XNOR U9982 ( .A(n5845), .B(n5844), .Z(n5862) );
  XNOR U9983 ( .A(n5859), .B(n5860), .Z(n5844) );
  XOR U9984 ( .A(n5856), .B(n5855), .Z(n5860) );
  XOR U9985 ( .A(y[3471]), .B(x[3471]), .Z(n5855) );
  XOR U9986 ( .A(n5858), .B(n5857), .Z(n5856) );
  XOR U9987 ( .A(y[3473]), .B(x[3473]), .Z(n5857) );
  XOR U9988 ( .A(y[3472]), .B(x[3472]), .Z(n5858) );
  XOR U9989 ( .A(n5850), .B(n5849), .Z(n5859) );
  XOR U9990 ( .A(n5852), .B(n5851), .Z(n5849) );
  XOR U9991 ( .A(y[3470]), .B(x[3470]), .Z(n5851) );
  XOR U9992 ( .A(y[3469]), .B(x[3469]), .Z(n5852) );
  XOR U9993 ( .A(y[3468]), .B(x[3468]), .Z(n5850) );
  XNOR U9994 ( .A(n5843), .B(n5842), .Z(n5845) );
  XNOR U9995 ( .A(n5839), .B(n5838), .Z(n5842) );
  XOR U9996 ( .A(n5841), .B(n5840), .Z(n5838) );
  XOR U9997 ( .A(y[3467]), .B(x[3467]), .Z(n5840) );
  XOR U9998 ( .A(y[3466]), .B(x[3466]), .Z(n5841) );
  XOR U9999 ( .A(y[3465]), .B(x[3465]), .Z(n5839) );
  XOR U10000 ( .A(n5833), .B(n5832), .Z(n5843) );
  XOR U10001 ( .A(n5835), .B(n5834), .Z(n5832) );
  XOR U10002 ( .A(y[3464]), .B(x[3464]), .Z(n5834) );
  XOR U10003 ( .A(y[3463]), .B(x[3463]), .Z(n5835) );
  XOR U10004 ( .A(y[3462]), .B(x[3462]), .Z(n5833) );
  NAND U10005 ( .A(n5896), .B(n5897), .Z(N29661) );
  NAND U10006 ( .A(n5898), .B(n5899), .Z(n5897) );
  NANDN U10007 ( .A(n5900), .B(n5901), .Z(n5899) );
  NANDN U10008 ( .A(n5901), .B(n5900), .Z(n5896) );
  XOR U10009 ( .A(n5900), .B(n5902), .Z(N29660) );
  XNOR U10010 ( .A(n5898), .B(n5901), .Z(n5902) );
  NAND U10011 ( .A(n5903), .B(n5904), .Z(n5901) );
  NAND U10012 ( .A(n5905), .B(n5906), .Z(n5904) );
  NANDN U10013 ( .A(n5907), .B(n5908), .Z(n5906) );
  NANDN U10014 ( .A(n5908), .B(n5907), .Z(n5903) );
  AND U10015 ( .A(n5909), .B(n5910), .Z(n5898) );
  NAND U10016 ( .A(n5911), .B(n5912), .Z(n5910) );
  OR U10017 ( .A(n5913), .B(n5914), .Z(n5912) );
  NAND U10018 ( .A(n5914), .B(n5913), .Z(n5909) );
  IV U10019 ( .A(n5915), .Z(n5914) );
  AND U10020 ( .A(n5916), .B(n5917), .Z(n5900) );
  NAND U10021 ( .A(n5918), .B(n5919), .Z(n5917) );
  NANDN U10022 ( .A(n5920), .B(n5921), .Z(n5919) );
  NANDN U10023 ( .A(n5921), .B(n5920), .Z(n5916) );
  XOR U10024 ( .A(n5913), .B(n5922), .Z(N29659) );
  XOR U10025 ( .A(n5911), .B(n5915), .Z(n5922) );
  XNOR U10026 ( .A(n5908), .B(n5923), .Z(n5915) );
  XNOR U10027 ( .A(n5905), .B(n5907), .Z(n5923) );
  AND U10028 ( .A(n5924), .B(n5925), .Z(n5907) );
  NANDN U10029 ( .A(n5926), .B(n5927), .Z(n5925) );
  NANDN U10030 ( .A(n5928), .B(n5929), .Z(n5927) );
  IV U10031 ( .A(n5930), .Z(n5929) );
  NAND U10032 ( .A(n5930), .B(n5928), .Z(n5924) );
  AND U10033 ( .A(n5931), .B(n5932), .Z(n5905) );
  NAND U10034 ( .A(n5933), .B(n5934), .Z(n5932) );
  OR U10035 ( .A(n5935), .B(n5936), .Z(n5934) );
  NAND U10036 ( .A(n5936), .B(n5935), .Z(n5931) );
  IV U10037 ( .A(n5937), .Z(n5936) );
  NAND U10038 ( .A(n5938), .B(n5939), .Z(n5908) );
  NANDN U10039 ( .A(n5940), .B(n5941), .Z(n5939) );
  NAND U10040 ( .A(n5942), .B(n5943), .Z(n5941) );
  OR U10041 ( .A(n5943), .B(n5942), .Z(n5938) );
  IV U10042 ( .A(n5944), .Z(n5942) );
  AND U10043 ( .A(n5945), .B(n5946), .Z(n5911) );
  NAND U10044 ( .A(n5947), .B(n5948), .Z(n5946) );
  NANDN U10045 ( .A(n5949), .B(n5950), .Z(n5948) );
  NANDN U10046 ( .A(n5950), .B(n5949), .Z(n5945) );
  XOR U10047 ( .A(n5921), .B(n5951), .Z(n5913) );
  XNOR U10048 ( .A(n5918), .B(n5920), .Z(n5951) );
  AND U10049 ( .A(n5952), .B(n5953), .Z(n5920) );
  NANDN U10050 ( .A(n5954), .B(n5955), .Z(n5953) );
  NANDN U10051 ( .A(n5956), .B(n5957), .Z(n5955) );
  IV U10052 ( .A(n5958), .Z(n5957) );
  NAND U10053 ( .A(n5958), .B(n5956), .Z(n5952) );
  AND U10054 ( .A(n5959), .B(n5960), .Z(n5918) );
  NAND U10055 ( .A(n5961), .B(n5962), .Z(n5960) );
  OR U10056 ( .A(n5963), .B(n5964), .Z(n5962) );
  NAND U10057 ( .A(n5964), .B(n5963), .Z(n5959) );
  IV U10058 ( .A(n5965), .Z(n5964) );
  NAND U10059 ( .A(n5966), .B(n5967), .Z(n5921) );
  NANDN U10060 ( .A(n5968), .B(n5969), .Z(n5967) );
  NAND U10061 ( .A(n5970), .B(n5971), .Z(n5969) );
  OR U10062 ( .A(n5971), .B(n5970), .Z(n5966) );
  IV U10063 ( .A(n5972), .Z(n5970) );
  XOR U10064 ( .A(n5947), .B(n5973), .Z(N29658) );
  XNOR U10065 ( .A(n5950), .B(n5949), .Z(n5973) );
  XNOR U10066 ( .A(n5961), .B(n5974), .Z(n5949) );
  XOR U10067 ( .A(n5965), .B(n5963), .Z(n5974) );
  XOR U10068 ( .A(n5971), .B(n5975), .Z(n5963) );
  XOR U10069 ( .A(n5968), .B(n5972), .Z(n5975) );
  NAND U10070 ( .A(n5976), .B(n5977), .Z(n5972) );
  NAND U10071 ( .A(n5978), .B(n5979), .Z(n5977) );
  NAND U10072 ( .A(n5980), .B(n5981), .Z(n5976) );
  AND U10073 ( .A(n5982), .B(n5983), .Z(n5968) );
  NAND U10074 ( .A(n5984), .B(n5985), .Z(n5983) );
  NAND U10075 ( .A(n5986), .B(n5987), .Z(n5982) );
  NANDN U10076 ( .A(n5988), .B(n5989), .Z(n5971) );
  NANDN U10077 ( .A(n5990), .B(n5991), .Z(n5965) );
  XNOR U10078 ( .A(n5956), .B(n5992), .Z(n5961) );
  XOR U10079 ( .A(n5954), .B(n5958), .Z(n5992) );
  NAND U10080 ( .A(n5993), .B(n5994), .Z(n5958) );
  NAND U10081 ( .A(n5995), .B(n5996), .Z(n5994) );
  NAND U10082 ( .A(n5997), .B(n5998), .Z(n5993) );
  AND U10083 ( .A(n5999), .B(n6000), .Z(n5954) );
  NAND U10084 ( .A(n6001), .B(n6002), .Z(n6000) );
  NAND U10085 ( .A(n6003), .B(n6004), .Z(n5999) );
  AND U10086 ( .A(n6005), .B(n6006), .Z(n5956) );
  NAND U10087 ( .A(n6007), .B(n6008), .Z(n5950) );
  XNOR U10088 ( .A(n5933), .B(n6009), .Z(n5947) );
  XOR U10089 ( .A(n5937), .B(n5935), .Z(n6009) );
  XOR U10090 ( .A(n5943), .B(n6010), .Z(n5935) );
  XOR U10091 ( .A(n5940), .B(n5944), .Z(n6010) );
  NAND U10092 ( .A(n6011), .B(n6012), .Z(n5944) );
  NAND U10093 ( .A(n6013), .B(n6014), .Z(n6012) );
  NAND U10094 ( .A(n6015), .B(n6016), .Z(n6011) );
  AND U10095 ( .A(n6017), .B(n6018), .Z(n5940) );
  NAND U10096 ( .A(n6019), .B(n6020), .Z(n6018) );
  NAND U10097 ( .A(n6021), .B(n6022), .Z(n6017) );
  NANDN U10098 ( .A(n6023), .B(n6024), .Z(n5943) );
  NANDN U10099 ( .A(n6025), .B(n6026), .Z(n5937) );
  XNOR U10100 ( .A(n5928), .B(n6027), .Z(n5933) );
  XOR U10101 ( .A(n5926), .B(n5930), .Z(n6027) );
  NAND U10102 ( .A(n6028), .B(n6029), .Z(n5930) );
  NAND U10103 ( .A(n6030), .B(n6031), .Z(n6029) );
  NAND U10104 ( .A(n6032), .B(n6033), .Z(n6028) );
  AND U10105 ( .A(n6034), .B(n6035), .Z(n5926) );
  NAND U10106 ( .A(n6036), .B(n6037), .Z(n6035) );
  NAND U10107 ( .A(n6038), .B(n6039), .Z(n6034) );
  AND U10108 ( .A(n6040), .B(n6041), .Z(n5928) );
  XOR U10109 ( .A(n6008), .B(n6007), .Z(N29657) );
  XNOR U10110 ( .A(n6026), .B(n6025), .Z(n6007) );
  XNOR U10111 ( .A(n6040), .B(n6041), .Z(n6025) );
  XOR U10112 ( .A(n6037), .B(n6036), .Z(n6041) );
  XOR U10113 ( .A(y[3459]), .B(x[3459]), .Z(n6036) );
  XOR U10114 ( .A(n6039), .B(n6038), .Z(n6037) );
  XOR U10115 ( .A(y[3461]), .B(x[3461]), .Z(n6038) );
  XOR U10116 ( .A(y[3460]), .B(x[3460]), .Z(n6039) );
  XOR U10117 ( .A(n6031), .B(n6030), .Z(n6040) );
  XOR U10118 ( .A(n6033), .B(n6032), .Z(n6030) );
  XOR U10119 ( .A(y[3458]), .B(x[3458]), .Z(n6032) );
  XOR U10120 ( .A(y[3457]), .B(x[3457]), .Z(n6033) );
  XOR U10121 ( .A(y[3456]), .B(x[3456]), .Z(n6031) );
  XNOR U10122 ( .A(n6024), .B(n6023), .Z(n6026) );
  XNOR U10123 ( .A(n6020), .B(n6019), .Z(n6023) );
  XOR U10124 ( .A(n6022), .B(n6021), .Z(n6019) );
  XOR U10125 ( .A(y[3455]), .B(x[3455]), .Z(n6021) );
  XOR U10126 ( .A(y[3454]), .B(x[3454]), .Z(n6022) );
  XOR U10127 ( .A(y[3453]), .B(x[3453]), .Z(n6020) );
  XOR U10128 ( .A(n6014), .B(n6013), .Z(n6024) );
  XOR U10129 ( .A(n6016), .B(n6015), .Z(n6013) );
  XOR U10130 ( .A(y[3452]), .B(x[3452]), .Z(n6015) );
  XOR U10131 ( .A(y[3451]), .B(x[3451]), .Z(n6016) );
  XOR U10132 ( .A(y[3450]), .B(x[3450]), .Z(n6014) );
  XNOR U10133 ( .A(n5991), .B(n5990), .Z(n6008) );
  XNOR U10134 ( .A(n6005), .B(n6006), .Z(n5990) );
  XOR U10135 ( .A(n6002), .B(n6001), .Z(n6006) );
  XOR U10136 ( .A(y[3447]), .B(x[3447]), .Z(n6001) );
  XOR U10137 ( .A(n6004), .B(n6003), .Z(n6002) );
  XOR U10138 ( .A(y[3449]), .B(x[3449]), .Z(n6003) );
  XOR U10139 ( .A(y[3448]), .B(x[3448]), .Z(n6004) );
  XOR U10140 ( .A(n5996), .B(n5995), .Z(n6005) );
  XOR U10141 ( .A(n5998), .B(n5997), .Z(n5995) );
  XOR U10142 ( .A(y[3446]), .B(x[3446]), .Z(n5997) );
  XOR U10143 ( .A(y[3445]), .B(x[3445]), .Z(n5998) );
  XOR U10144 ( .A(y[3444]), .B(x[3444]), .Z(n5996) );
  XNOR U10145 ( .A(n5989), .B(n5988), .Z(n5991) );
  XNOR U10146 ( .A(n5985), .B(n5984), .Z(n5988) );
  XOR U10147 ( .A(n5987), .B(n5986), .Z(n5984) );
  XOR U10148 ( .A(y[3443]), .B(x[3443]), .Z(n5986) );
  XOR U10149 ( .A(y[3442]), .B(x[3442]), .Z(n5987) );
  XOR U10150 ( .A(y[3441]), .B(x[3441]), .Z(n5985) );
  XOR U10151 ( .A(n5979), .B(n5978), .Z(n5989) );
  XOR U10152 ( .A(n5981), .B(n5980), .Z(n5978) );
  XOR U10153 ( .A(y[3440]), .B(x[3440]), .Z(n5980) );
  XOR U10154 ( .A(y[3439]), .B(x[3439]), .Z(n5981) );
  XOR U10155 ( .A(y[3438]), .B(x[3438]), .Z(n5979) );
  NAND U10156 ( .A(n6042), .B(n6043), .Z(N29649) );
  NAND U10157 ( .A(n6044), .B(n6045), .Z(n6043) );
  NANDN U10158 ( .A(n6046), .B(n6047), .Z(n6045) );
  NANDN U10159 ( .A(n6047), .B(n6046), .Z(n6042) );
  XOR U10160 ( .A(n6046), .B(n6048), .Z(N29648) );
  XNOR U10161 ( .A(n6044), .B(n6047), .Z(n6048) );
  NAND U10162 ( .A(n6049), .B(n6050), .Z(n6047) );
  NAND U10163 ( .A(n6051), .B(n6052), .Z(n6050) );
  NANDN U10164 ( .A(n6053), .B(n6054), .Z(n6052) );
  NANDN U10165 ( .A(n6054), .B(n6053), .Z(n6049) );
  AND U10166 ( .A(n6055), .B(n6056), .Z(n6044) );
  NAND U10167 ( .A(n6057), .B(n6058), .Z(n6056) );
  OR U10168 ( .A(n6059), .B(n6060), .Z(n6058) );
  NAND U10169 ( .A(n6060), .B(n6059), .Z(n6055) );
  IV U10170 ( .A(n6061), .Z(n6060) );
  AND U10171 ( .A(n6062), .B(n6063), .Z(n6046) );
  NAND U10172 ( .A(n6064), .B(n6065), .Z(n6063) );
  NANDN U10173 ( .A(n6066), .B(n6067), .Z(n6065) );
  NANDN U10174 ( .A(n6067), .B(n6066), .Z(n6062) );
  XOR U10175 ( .A(n6059), .B(n6068), .Z(N29647) );
  XOR U10176 ( .A(n6057), .B(n6061), .Z(n6068) );
  XNOR U10177 ( .A(n6054), .B(n6069), .Z(n6061) );
  XNOR U10178 ( .A(n6051), .B(n6053), .Z(n6069) );
  AND U10179 ( .A(n6070), .B(n6071), .Z(n6053) );
  NANDN U10180 ( .A(n6072), .B(n6073), .Z(n6071) );
  NANDN U10181 ( .A(n6074), .B(n6075), .Z(n6073) );
  IV U10182 ( .A(n6076), .Z(n6075) );
  NAND U10183 ( .A(n6076), .B(n6074), .Z(n6070) );
  AND U10184 ( .A(n6077), .B(n6078), .Z(n6051) );
  NAND U10185 ( .A(n6079), .B(n6080), .Z(n6078) );
  OR U10186 ( .A(n6081), .B(n6082), .Z(n6080) );
  NAND U10187 ( .A(n6082), .B(n6081), .Z(n6077) );
  IV U10188 ( .A(n6083), .Z(n6082) );
  NAND U10189 ( .A(n6084), .B(n6085), .Z(n6054) );
  NANDN U10190 ( .A(n6086), .B(n6087), .Z(n6085) );
  NAND U10191 ( .A(n6088), .B(n6089), .Z(n6087) );
  OR U10192 ( .A(n6089), .B(n6088), .Z(n6084) );
  IV U10193 ( .A(n6090), .Z(n6088) );
  AND U10194 ( .A(n6091), .B(n6092), .Z(n6057) );
  NAND U10195 ( .A(n6093), .B(n6094), .Z(n6092) );
  NANDN U10196 ( .A(n6095), .B(n6096), .Z(n6094) );
  NANDN U10197 ( .A(n6096), .B(n6095), .Z(n6091) );
  XOR U10198 ( .A(n6067), .B(n6097), .Z(n6059) );
  XNOR U10199 ( .A(n6064), .B(n6066), .Z(n6097) );
  AND U10200 ( .A(n6098), .B(n6099), .Z(n6066) );
  NANDN U10201 ( .A(n6100), .B(n6101), .Z(n6099) );
  NANDN U10202 ( .A(n6102), .B(n6103), .Z(n6101) );
  IV U10203 ( .A(n6104), .Z(n6103) );
  NAND U10204 ( .A(n6104), .B(n6102), .Z(n6098) );
  AND U10205 ( .A(n6105), .B(n6106), .Z(n6064) );
  NAND U10206 ( .A(n6107), .B(n6108), .Z(n6106) );
  OR U10207 ( .A(n6109), .B(n6110), .Z(n6108) );
  NAND U10208 ( .A(n6110), .B(n6109), .Z(n6105) );
  IV U10209 ( .A(n6111), .Z(n6110) );
  NAND U10210 ( .A(n6112), .B(n6113), .Z(n6067) );
  NANDN U10211 ( .A(n6114), .B(n6115), .Z(n6113) );
  NAND U10212 ( .A(n6116), .B(n6117), .Z(n6115) );
  OR U10213 ( .A(n6117), .B(n6116), .Z(n6112) );
  IV U10214 ( .A(n6118), .Z(n6116) );
  XOR U10215 ( .A(n6093), .B(n6119), .Z(N29646) );
  XNOR U10216 ( .A(n6096), .B(n6095), .Z(n6119) );
  XNOR U10217 ( .A(n6107), .B(n6120), .Z(n6095) );
  XOR U10218 ( .A(n6111), .B(n6109), .Z(n6120) );
  XOR U10219 ( .A(n6117), .B(n6121), .Z(n6109) );
  XOR U10220 ( .A(n6114), .B(n6118), .Z(n6121) );
  NAND U10221 ( .A(n6122), .B(n6123), .Z(n6118) );
  NAND U10222 ( .A(n6124), .B(n6125), .Z(n6123) );
  NAND U10223 ( .A(n6126), .B(n6127), .Z(n6122) );
  AND U10224 ( .A(n6128), .B(n6129), .Z(n6114) );
  NAND U10225 ( .A(n6130), .B(n6131), .Z(n6129) );
  NAND U10226 ( .A(n6132), .B(n6133), .Z(n6128) );
  NANDN U10227 ( .A(n6134), .B(n6135), .Z(n6117) );
  NANDN U10228 ( .A(n6136), .B(n6137), .Z(n6111) );
  XNOR U10229 ( .A(n6102), .B(n6138), .Z(n6107) );
  XOR U10230 ( .A(n6100), .B(n6104), .Z(n6138) );
  NAND U10231 ( .A(n6139), .B(n6140), .Z(n6104) );
  NAND U10232 ( .A(n6141), .B(n6142), .Z(n6140) );
  NAND U10233 ( .A(n6143), .B(n6144), .Z(n6139) );
  AND U10234 ( .A(n6145), .B(n6146), .Z(n6100) );
  NAND U10235 ( .A(n6147), .B(n6148), .Z(n6146) );
  NAND U10236 ( .A(n6149), .B(n6150), .Z(n6145) );
  AND U10237 ( .A(n6151), .B(n6152), .Z(n6102) );
  NAND U10238 ( .A(n6153), .B(n6154), .Z(n6096) );
  XNOR U10239 ( .A(n6079), .B(n6155), .Z(n6093) );
  XOR U10240 ( .A(n6083), .B(n6081), .Z(n6155) );
  XOR U10241 ( .A(n6089), .B(n6156), .Z(n6081) );
  XOR U10242 ( .A(n6086), .B(n6090), .Z(n6156) );
  NAND U10243 ( .A(n6157), .B(n6158), .Z(n6090) );
  NAND U10244 ( .A(n6159), .B(n6160), .Z(n6158) );
  NAND U10245 ( .A(n6161), .B(n6162), .Z(n6157) );
  AND U10246 ( .A(n6163), .B(n6164), .Z(n6086) );
  NAND U10247 ( .A(n6165), .B(n6166), .Z(n6164) );
  NAND U10248 ( .A(n6167), .B(n6168), .Z(n6163) );
  NANDN U10249 ( .A(n6169), .B(n6170), .Z(n6089) );
  NANDN U10250 ( .A(n6171), .B(n6172), .Z(n6083) );
  XNOR U10251 ( .A(n6074), .B(n6173), .Z(n6079) );
  XOR U10252 ( .A(n6072), .B(n6076), .Z(n6173) );
  NAND U10253 ( .A(n6174), .B(n6175), .Z(n6076) );
  NAND U10254 ( .A(n6176), .B(n6177), .Z(n6175) );
  NAND U10255 ( .A(n6178), .B(n6179), .Z(n6174) );
  AND U10256 ( .A(n6180), .B(n6181), .Z(n6072) );
  NAND U10257 ( .A(n6182), .B(n6183), .Z(n6181) );
  NAND U10258 ( .A(n6184), .B(n6185), .Z(n6180) );
  AND U10259 ( .A(n6186), .B(n6187), .Z(n6074) );
  XOR U10260 ( .A(n6154), .B(n6153), .Z(N29645) );
  XNOR U10261 ( .A(n6172), .B(n6171), .Z(n6153) );
  XNOR U10262 ( .A(n6186), .B(n6187), .Z(n6171) );
  XOR U10263 ( .A(n6183), .B(n6182), .Z(n6187) );
  XOR U10264 ( .A(y[3435]), .B(x[3435]), .Z(n6182) );
  XOR U10265 ( .A(n6185), .B(n6184), .Z(n6183) );
  XOR U10266 ( .A(y[3437]), .B(x[3437]), .Z(n6184) );
  XOR U10267 ( .A(y[3436]), .B(x[3436]), .Z(n6185) );
  XOR U10268 ( .A(n6177), .B(n6176), .Z(n6186) );
  XOR U10269 ( .A(n6179), .B(n6178), .Z(n6176) );
  XOR U10270 ( .A(y[3434]), .B(x[3434]), .Z(n6178) );
  XOR U10271 ( .A(y[3433]), .B(x[3433]), .Z(n6179) );
  XOR U10272 ( .A(y[3432]), .B(x[3432]), .Z(n6177) );
  XNOR U10273 ( .A(n6170), .B(n6169), .Z(n6172) );
  XNOR U10274 ( .A(n6166), .B(n6165), .Z(n6169) );
  XOR U10275 ( .A(n6168), .B(n6167), .Z(n6165) );
  XOR U10276 ( .A(y[3431]), .B(x[3431]), .Z(n6167) );
  XOR U10277 ( .A(y[3430]), .B(x[3430]), .Z(n6168) );
  XOR U10278 ( .A(y[3429]), .B(x[3429]), .Z(n6166) );
  XOR U10279 ( .A(n6160), .B(n6159), .Z(n6170) );
  XOR U10280 ( .A(n6162), .B(n6161), .Z(n6159) );
  XOR U10281 ( .A(y[3428]), .B(x[3428]), .Z(n6161) );
  XOR U10282 ( .A(y[3427]), .B(x[3427]), .Z(n6162) );
  XOR U10283 ( .A(y[3426]), .B(x[3426]), .Z(n6160) );
  XNOR U10284 ( .A(n6137), .B(n6136), .Z(n6154) );
  XNOR U10285 ( .A(n6151), .B(n6152), .Z(n6136) );
  XOR U10286 ( .A(n6148), .B(n6147), .Z(n6152) );
  XOR U10287 ( .A(y[3423]), .B(x[3423]), .Z(n6147) );
  XOR U10288 ( .A(n6150), .B(n6149), .Z(n6148) );
  XOR U10289 ( .A(y[3425]), .B(x[3425]), .Z(n6149) );
  XOR U10290 ( .A(y[3424]), .B(x[3424]), .Z(n6150) );
  XOR U10291 ( .A(n6142), .B(n6141), .Z(n6151) );
  XOR U10292 ( .A(n6144), .B(n6143), .Z(n6141) );
  XOR U10293 ( .A(y[3422]), .B(x[3422]), .Z(n6143) );
  XOR U10294 ( .A(y[3421]), .B(x[3421]), .Z(n6144) );
  XOR U10295 ( .A(y[3420]), .B(x[3420]), .Z(n6142) );
  XNOR U10296 ( .A(n6135), .B(n6134), .Z(n6137) );
  XNOR U10297 ( .A(n6131), .B(n6130), .Z(n6134) );
  XOR U10298 ( .A(n6133), .B(n6132), .Z(n6130) );
  XOR U10299 ( .A(y[3419]), .B(x[3419]), .Z(n6132) );
  XOR U10300 ( .A(y[3418]), .B(x[3418]), .Z(n6133) );
  XOR U10301 ( .A(y[3417]), .B(x[3417]), .Z(n6131) );
  XOR U10302 ( .A(n6125), .B(n6124), .Z(n6135) );
  XOR U10303 ( .A(n6127), .B(n6126), .Z(n6124) );
  XOR U10304 ( .A(y[3416]), .B(x[3416]), .Z(n6126) );
  XOR U10305 ( .A(y[3415]), .B(x[3415]), .Z(n6127) );
  XOR U10306 ( .A(y[3414]), .B(x[3414]), .Z(n6125) );
  NAND U10307 ( .A(n6188), .B(n6189), .Z(N29637) );
  NAND U10308 ( .A(n6190), .B(n6191), .Z(n6189) );
  NANDN U10309 ( .A(n6192), .B(n6193), .Z(n6191) );
  NANDN U10310 ( .A(n6193), .B(n6192), .Z(n6188) );
  XOR U10311 ( .A(n6192), .B(n6194), .Z(N29636) );
  XNOR U10312 ( .A(n6190), .B(n6193), .Z(n6194) );
  NAND U10313 ( .A(n6195), .B(n6196), .Z(n6193) );
  NAND U10314 ( .A(n6197), .B(n6198), .Z(n6196) );
  NANDN U10315 ( .A(n6199), .B(n6200), .Z(n6198) );
  NANDN U10316 ( .A(n6200), .B(n6199), .Z(n6195) );
  AND U10317 ( .A(n6201), .B(n6202), .Z(n6190) );
  NAND U10318 ( .A(n6203), .B(n6204), .Z(n6202) );
  OR U10319 ( .A(n6205), .B(n6206), .Z(n6204) );
  NAND U10320 ( .A(n6206), .B(n6205), .Z(n6201) );
  IV U10321 ( .A(n6207), .Z(n6206) );
  AND U10322 ( .A(n6208), .B(n6209), .Z(n6192) );
  NAND U10323 ( .A(n6210), .B(n6211), .Z(n6209) );
  NANDN U10324 ( .A(n6212), .B(n6213), .Z(n6211) );
  NANDN U10325 ( .A(n6213), .B(n6212), .Z(n6208) );
  XOR U10326 ( .A(n6205), .B(n6214), .Z(N29635) );
  XOR U10327 ( .A(n6203), .B(n6207), .Z(n6214) );
  XNOR U10328 ( .A(n6200), .B(n6215), .Z(n6207) );
  XNOR U10329 ( .A(n6197), .B(n6199), .Z(n6215) );
  AND U10330 ( .A(n6216), .B(n6217), .Z(n6199) );
  NANDN U10331 ( .A(n6218), .B(n6219), .Z(n6217) );
  NANDN U10332 ( .A(n6220), .B(n6221), .Z(n6219) );
  IV U10333 ( .A(n6222), .Z(n6221) );
  NAND U10334 ( .A(n6222), .B(n6220), .Z(n6216) );
  AND U10335 ( .A(n6223), .B(n6224), .Z(n6197) );
  NAND U10336 ( .A(n6225), .B(n6226), .Z(n6224) );
  OR U10337 ( .A(n6227), .B(n6228), .Z(n6226) );
  NAND U10338 ( .A(n6228), .B(n6227), .Z(n6223) );
  IV U10339 ( .A(n6229), .Z(n6228) );
  NAND U10340 ( .A(n6230), .B(n6231), .Z(n6200) );
  NANDN U10341 ( .A(n6232), .B(n6233), .Z(n6231) );
  NAND U10342 ( .A(n6234), .B(n6235), .Z(n6233) );
  OR U10343 ( .A(n6235), .B(n6234), .Z(n6230) );
  IV U10344 ( .A(n6236), .Z(n6234) );
  AND U10345 ( .A(n6237), .B(n6238), .Z(n6203) );
  NAND U10346 ( .A(n6239), .B(n6240), .Z(n6238) );
  NANDN U10347 ( .A(n6241), .B(n6242), .Z(n6240) );
  NANDN U10348 ( .A(n6242), .B(n6241), .Z(n6237) );
  XOR U10349 ( .A(n6213), .B(n6243), .Z(n6205) );
  XNOR U10350 ( .A(n6210), .B(n6212), .Z(n6243) );
  AND U10351 ( .A(n6244), .B(n6245), .Z(n6212) );
  NANDN U10352 ( .A(n6246), .B(n6247), .Z(n6245) );
  NANDN U10353 ( .A(n6248), .B(n6249), .Z(n6247) );
  IV U10354 ( .A(n6250), .Z(n6249) );
  NAND U10355 ( .A(n6250), .B(n6248), .Z(n6244) );
  AND U10356 ( .A(n6251), .B(n6252), .Z(n6210) );
  NAND U10357 ( .A(n6253), .B(n6254), .Z(n6252) );
  OR U10358 ( .A(n6255), .B(n6256), .Z(n6254) );
  NAND U10359 ( .A(n6256), .B(n6255), .Z(n6251) );
  IV U10360 ( .A(n6257), .Z(n6256) );
  NAND U10361 ( .A(n6258), .B(n6259), .Z(n6213) );
  NANDN U10362 ( .A(n6260), .B(n6261), .Z(n6259) );
  NAND U10363 ( .A(n6262), .B(n6263), .Z(n6261) );
  OR U10364 ( .A(n6263), .B(n6262), .Z(n6258) );
  IV U10365 ( .A(n6264), .Z(n6262) );
  XOR U10366 ( .A(n6239), .B(n6265), .Z(N29634) );
  XNOR U10367 ( .A(n6242), .B(n6241), .Z(n6265) );
  XNOR U10368 ( .A(n6253), .B(n6266), .Z(n6241) );
  XOR U10369 ( .A(n6257), .B(n6255), .Z(n6266) );
  XOR U10370 ( .A(n6263), .B(n6267), .Z(n6255) );
  XOR U10371 ( .A(n6260), .B(n6264), .Z(n6267) );
  NAND U10372 ( .A(n6268), .B(n6269), .Z(n6264) );
  NAND U10373 ( .A(n6270), .B(n6271), .Z(n6269) );
  NAND U10374 ( .A(n6272), .B(n6273), .Z(n6268) );
  AND U10375 ( .A(n6274), .B(n6275), .Z(n6260) );
  NAND U10376 ( .A(n6276), .B(n6277), .Z(n6275) );
  NAND U10377 ( .A(n6278), .B(n6279), .Z(n6274) );
  NANDN U10378 ( .A(n6280), .B(n6281), .Z(n6263) );
  NANDN U10379 ( .A(n6282), .B(n6283), .Z(n6257) );
  XNOR U10380 ( .A(n6248), .B(n6284), .Z(n6253) );
  XOR U10381 ( .A(n6246), .B(n6250), .Z(n6284) );
  NAND U10382 ( .A(n6285), .B(n6286), .Z(n6250) );
  NAND U10383 ( .A(n6287), .B(n6288), .Z(n6286) );
  NAND U10384 ( .A(n6289), .B(n6290), .Z(n6285) );
  AND U10385 ( .A(n6291), .B(n6292), .Z(n6246) );
  NAND U10386 ( .A(n6293), .B(n6294), .Z(n6292) );
  NAND U10387 ( .A(n6295), .B(n6296), .Z(n6291) );
  AND U10388 ( .A(n6297), .B(n6298), .Z(n6248) );
  NAND U10389 ( .A(n6299), .B(n6300), .Z(n6242) );
  XNOR U10390 ( .A(n6225), .B(n6301), .Z(n6239) );
  XOR U10391 ( .A(n6229), .B(n6227), .Z(n6301) );
  XOR U10392 ( .A(n6235), .B(n6302), .Z(n6227) );
  XOR U10393 ( .A(n6232), .B(n6236), .Z(n6302) );
  NAND U10394 ( .A(n6303), .B(n6304), .Z(n6236) );
  NAND U10395 ( .A(n6305), .B(n6306), .Z(n6304) );
  NAND U10396 ( .A(n6307), .B(n6308), .Z(n6303) );
  AND U10397 ( .A(n6309), .B(n6310), .Z(n6232) );
  NAND U10398 ( .A(n6311), .B(n6312), .Z(n6310) );
  NAND U10399 ( .A(n6313), .B(n6314), .Z(n6309) );
  NANDN U10400 ( .A(n6315), .B(n6316), .Z(n6235) );
  NANDN U10401 ( .A(n6317), .B(n6318), .Z(n6229) );
  XNOR U10402 ( .A(n6220), .B(n6319), .Z(n6225) );
  XOR U10403 ( .A(n6218), .B(n6222), .Z(n6319) );
  NAND U10404 ( .A(n6320), .B(n6321), .Z(n6222) );
  NAND U10405 ( .A(n6322), .B(n6323), .Z(n6321) );
  NAND U10406 ( .A(n6324), .B(n6325), .Z(n6320) );
  AND U10407 ( .A(n6326), .B(n6327), .Z(n6218) );
  NAND U10408 ( .A(n6328), .B(n6329), .Z(n6327) );
  NAND U10409 ( .A(n6330), .B(n6331), .Z(n6326) );
  AND U10410 ( .A(n6332), .B(n6333), .Z(n6220) );
  XOR U10411 ( .A(n6300), .B(n6299), .Z(N29633) );
  XNOR U10412 ( .A(n6318), .B(n6317), .Z(n6299) );
  XNOR U10413 ( .A(n6332), .B(n6333), .Z(n6317) );
  XOR U10414 ( .A(n6329), .B(n6328), .Z(n6333) );
  XOR U10415 ( .A(y[3411]), .B(x[3411]), .Z(n6328) );
  XOR U10416 ( .A(n6331), .B(n6330), .Z(n6329) );
  XOR U10417 ( .A(y[3413]), .B(x[3413]), .Z(n6330) );
  XOR U10418 ( .A(y[3412]), .B(x[3412]), .Z(n6331) );
  XOR U10419 ( .A(n6323), .B(n6322), .Z(n6332) );
  XOR U10420 ( .A(n6325), .B(n6324), .Z(n6322) );
  XOR U10421 ( .A(y[3410]), .B(x[3410]), .Z(n6324) );
  XOR U10422 ( .A(y[3409]), .B(x[3409]), .Z(n6325) );
  XOR U10423 ( .A(y[3408]), .B(x[3408]), .Z(n6323) );
  XNOR U10424 ( .A(n6316), .B(n6315), .Z(n6318) );
  XNOR U10425 ( .A(n6312), .B(n6311), .Z(n6315) );
  XOR U10426 ( .A(n6314), .B(n6313), .Z(n6311) );
  XOR U10427 ( .A(y[3407]), .B(x[3407]), .Z(n6313) );
  XOR U10428 ( .A(y[3406]), .B(x[3406]), .Z(n6314) );
  XOR U10429 ( .A(y[3405]), .B(x[3405]), .Z(n6312) );
  XOR U10430 ( .A(n6306), .B(n6305), .Z(n6316) );
  XOR U10431 ( .A(n6308), .B(n6307), .Z(n6305) );
  XOR U10432 ( .A(y[3404]), .B(x[3404]), .Z(n6307) );
  XOR U10433 ( .A(y[3403]), .B(x[3403]), .Z(n6308) );
  XOR U10434 ( .A(y[3402]), .B(x[3402]), .Z(n6306) );
  XNOR U10435 ( .A(n6283), .B(n6282), .Z(n6300) );
  XNOR U10436 ( .A(n6297), .B(n6298), .Z(n6282) );
  XOR U10437 ( .A(n6294), .B(n6293), .Z(n6298) );
  XOR U10438 ( .A(y[3399]), .B(x[3399]), .Z(n6293) );
  XOR U10439 ( .A(n6296), .B(n6295), .Z(n6294) );
  XOR U10440 ( .A(y[3401]), .B(x[3401]), .Z(n6295) );
  XOR U10441 ( .A(y[3400]), .B(x[3400]), .Z(n6296) );
  XOR U10442 ( .A(n6288), .B(n6287), .Z(n6297) );
  XOR U10443 ( .A(n6290), .B(n6289), .Z(n6287) );
  XOR U10444 ( .A(y[3398]), .B(x[3398]), .Z(n6289) );
  XOR U10445 ( .A(y[3397]), .B(x[3397]), .Z(n6290) );
  XOR U10446 ( .A(y[3396]), .B(x[3396]), .Z(n6288) );
  XNOR U10447 ( .A(n6281), .B(n6280), .Z(n6283) );
  XNOR U10448 ( .A(n6277), .B(n6276), .Z(n6280) );
  XOR U10449 ( .A(n6279), .B(n6278), .Z(n6276) );
  XOR U10450 ( .A(y[3395]), .B(x[3395]), .Z(n6278) );
  XOR U10451 ( .A(y[3394]), .B(x[3394]), .Z(n6279) );
  XOR U10452 ( .A(y[3393]), .B(x[3393]), .Z(n6277) );
  XOR U10453 ( .A(n6271), .B(n6270), .Z(n6281) );
  XOR U10454 ( .A(n6273), .B(n6272), .Z(n6270) );
  XOR U10455 ( .A(y[3392]), .B(x[3392]), .Z(n6272) );
  XOR U10456 ( .A(y[3391]), .B(x[3391]), .Z(n6273) );
  XOR U10457 ( .A(y[3390]), .B(x[3390]), .Z(n6271) );
  NAND U10458 ( .A(n6334), .B(n6335), .Z(N29625) );
  NAND U10459 ( .A(n6336), .B(n6337), .Z(n6335) );
  NANDN U10460 ( .A(n6338), .B(n6339), .Z(n6337) );
  NANDN U10461 ( .A(n6339), .B(n6338), .Z(n6334) );
  XOR U10462 ( .A(n6338), .B(n6340), .Z(N29624) );
  XNOR U10463 ( .A(n6336), .B(n6339), .Z(n6340) );
  NAND U10464 ( .A(n6341), .B(n6342), .Z(n6339) );
  NAND U10465 ( .A(n6343), .B(n6344), .Z(n6342) );
  NANDN U10466 ( .A(n6345), .B(n6346), .Z(n6344) );
  NANDN U10467 ( .A(n6346), .B(n6345), .Z(n6341) );
  AND U10468 ( .A(n6347), .B(n6348), .Z(n6336) );
  NAND U10469 ( .A(n6349), .B(n6350), .Z(n6348) );
  OR U10470 ( .A(n6351), .B(n6352), .Z(n6350) );
  NAND U10471 ( .A(n6352), .B(n6351), .Z(n6347) );
  IV U10472 ( .A(n6353), .Z(n6352) );
  AND U10473 ( .A(n6354), .B(n6355), .Z(n6338) );
  NAND U10474 ( .A(n6356), .B(n6357), .Z(n6355) );
  NANDN U10475 ( .A(n6358), .B(n6359), .Z(n6357) );
  NANDN U10476 ( .A(n6359), .B(n6358), .Z(n6354) );
  XOR U10477 ( .A(n6351), .B(n6360), .Z(N29623) );
  XOR U10478 ( .A(n6349), .B(n6353), .Z(n6360) );
  XNOR U10479 ( .A(n6346), .B(n6361), .Z(n6353) );
  XNOR U10480 ( .A(n6343), .B(n6345), .Z(n6361) );
  AND U10481 ( .A(n6362), .B(n6363), .Z(n6345) );
  NANDN U10482 ( .A(n6364), .B(n6365), .Z(n6363) );
  NANDN U10483 ( .A(n6366), .B(n6367), .Z(n6365) );
  IV U10484 ( .A(n6368), .Z(n6367) );
  NAND U10485 ( .A(n6368), .B(n6366), .Z(n6362) );
  AND U10486 ( .A(n6369), .B(n6370), .Z(n6343) );
  NAND U10487 ( .A(n6371), .B(n6372), .Z(n6370) );
  OR U10488 ( .A(n6373), .B(n6374), .Z(n6372) );
  NAND U10489 ( .A(n6374), .B(n6373), .Z(n6369) );
  IV U10490 ( .A(n6375), .Z(n6374) );
  NAND U10491 ( .A(n6376), .B(n6377), .Z(n6346) );
  NANDN U10492 ( .A(n6378), .B(n6379), .Z(n6377) );
  NAND U10493 ( .A(n6380), .B(n6381), .Z(n6379) );
  OR U10494 ( .A(n6381), .B(n6380), .Z(n6376) );
  IV U10495 ( .A(n6382), .Z(n6380) );
  AND U10496 ( .A(n6383), .B(n6384), .Z(n6349) );
  NAND U10497 ( .A(n6385), .B(n6386), .Z(n6384) );
  NANDN U10498 ( .A(n6387), .B(n6388), .Z(n6386) );
  NANDN U10499 ( .A(n6388), .B(n6387), .Z(n6383) );
  XOR U10500 ( .A(n6359), .B(n6389), .Z(n6351) );
  XNOR U10501 ( .A(n6356), .B(n6358), .Z(n6389) );
  AND U10502 ( .A(n6390), .B(n6391), .Z(n6358) );
  NANDN U10503 ( .A(n6392), .B(n6393), .Z(n6391) );
  NANDN U10504 ( .A(n6394), .B(n6395), .Z(n6393) );
  IV U10505 ( .A(n6396), .Z(n6395) );
  NAND U10506 ( .A(n6396), .B(n6394), .Z(n6390) );
  AND U10507 ( .A(n6397), .B(n6398), .Z(n6356) );
  NAND U10508 ( .A(n6399), .B(n6400), .Z(n6398) );
  OR U10509 ( .A(n6401), .B(n6402), .Z(n6400) );
  NAND U10510 ( .A(n6402), .B(n6401), .Z(n6397) );
  IV U10511 ( .A(n6403), .Z(n6402) );
  NAND U10512 ( .A(n6404), .B(n6405), .Z(n6359) );
  NANDN U10513 ( .A(n6406), .B(n6407), .Z(n6405) );
  NAND U10514 ( .A(n6408), .B(n6409), .Z(n6407) );
  OR U10515 ( .A(n6409), .B(n6408), .Z(n6404) );
  IV U10516 ( .A(n6410), .Z(n6408) );
  XOR U10517 ( .A(n6385), .B(n6411), .Z(N29622) );
  XNOR U10518 ( .A(n6388), .B(n6387), .Z(n6411) );
  XNOR U10519 ( .A(n6399), .B(n6412), .Z(n6387) );
  XOR U10520 ( .A(n6403), .B(n6401), .Z(n6412) );
  XOR U10521 ( .A(n6409), .B(n6413), .Z(n6401) );
  XOR U10522 ( .A(n6406), .B(n6410), .Z(n6413) );
  NAND U10523 ( .A(n6414), .B(n6415), .Z(n6410) );
  NAND U10524 ( .A(n6416), .B(n6417), .Z(n6415) );
  NAND U10525 ( .A(n6418), .B(n6419), .Z(n6414) );
  AND U10526 ( .A(n6420), .B(n6421), .Z(n6406) );
  NAND U10527 ( .A(n6422), .B(n6423), .Z(n6421) );
  NAND U10528 ( .A(n6424), .B(n6425), .Z(n6420) );
  NANDN U10529 ( .A(n6426), .B(n6427), .Z(n6409) );
  NANDN U10530 ( .A(n6428), .B(n6429), .Z(n6403) );
  XNOR U10531 ( .A(n6394), .B(n6430), .Z(n6399) );
  XOR U10532 ( .A(n6392), .B(n6396), .Z(n6430) );
  NAND U10533 ( .A(n6431), .B(n6432), .Z(n6396) );
  NAND U10534 ( .A(n6433), .B(n6434), .Z(n6432) );
  NAND U10535 ( .A(n6435), .B(n6436), .Z(n6431) );
  AND U10536 ( .A(n6437), .B(n6438), .Z(n6392) );
  NAND U10537 ( .A(n6439), .B(n6440), .Z(n6438) );
  NAND U10538 ( .A(n6441), .B(n6442), .Z(n6437) );
  AND U10539 ( .A(n6443), .B(n6444), .Z(n6394) );
  NAND U10540 ( .A(n6445), .B(n6446), .Z(n6388) );
  XNOR U10541 ( .A(n6371), .B(n6447), .Z(n6385) );
  XOR U10542 ( .A(n6375), .B(n6373), .Z(n6447) );
  XOR U10543 ( .A(n6381), .B(n6448), .Z(n6373) );
  XOR U10544 ( .A(n6378), .B(n6382), .Z(n6448) );
  NAND U10545 ( .A(n6449), .B(n6450), .Z(n6382) );
  NAND U10546 ( .A(n6451), .B(n6452), .Z(n6450) );
  NAND U10547 ( .A(n6453), .B(n6454), .Z(n6449) );
  AND U10548 ( .A(n6455), .B(n6456), .Z(n6378) );
  NAND U10549 ( .A(n6457), .B(n6458), .Z(n6456) );
  NAND U10550 ( .A(n6459), .B(n6460), .Z(n6455) );
  NANDN U10551 ( .A(n6461), .B(n6462), .Z(n6381) );
  NANDN U10552 ( .A(n6463), .B(n6464), .Z(n6375) );
  XNOR U10553 ( .A(n6366), .B(n6465), .Z(n6371) );
  XOR U10554 ( .A(n6364), .B(n6368), .Z(n6465) );
  NAND U10555 ( .A(n6466), .B(n6467), .Z(n6368) );
  NAND U10556 ( .A(n6468), .B(n6469), .Z(n6467) );
  NAND U10557 ( .A(n6470), .B(n6471), .Z(n6466) );
  AND U10558 ( .A(n6472), .B(n6473), .Z(n6364) );
  NAND U10559 ( .A(n6474), .B(n6475), .Z(n6473) );
  NAND U10560 ( .A(n6476), .B(n6477), .Z(n6472) );
  AND U10561 ( .A(n6478), .B(n6479), .Z(n6366) );
  XOR U10562 ( .A(n6446), .B(n6445), .Z(N29621) );
  XNOR U10563 ( .A(n6464), .B(n6463), .Z(n6445) );
  XNOR U10564 ( .A(n6478), .B(n6479), .Z(n6463) );
  XOR U10565 ( .A(n6475), .B(n6474), .Z(n6479) );
  XOR U10566 ( .A(y[3387]), .B(x[3387]), .Z(n6474) );
  XOR U10567 ( .A(n6477), .B(n6476), .Z(n6475) );
  XOR U10568 ( .A(y[3389]), .B(x[3389]), .Z(n6476) );
  XOR U10569 ( .A(y[3388]), .B(x[3388]), .Z(n6477) );
  XOR U10570 ( .A(n6469), .B(n6468), .Z(n6478) );
  XOR U10571 ( .A(n6471), .B(n6470), .Z(n6468) );
  XOR U10572 ( .A(y[3386]), .B(x[3386]), .Z(n6470) );
  XOR U10573 ( .A(y[3385]), .B(x[3385]), .Z(n6471) );
  XOR U10574 ( .A(y[3384]), .B(x[3384]), .Z(n6469) );
  XNOR U10575 ( .A(n6462), .B(n6461), .Z(n6464) );
  XNOR U10576 ( .A(n6458), .B(n6457), .Z(n6461) );
  XOR U10577 ( .A(n6460), .B(n6459), .Z(n6457) );
  XOR U10578 ( .A(y[3383]), .B(x[3383]), .Z(n6459) );
  XOR U10579 ( .A(y[3382]), .B(x[3382]), .Z(n6460) );
  XOR U10580 ( .A(y[3381]), .B(x[3381]), .Z(n6458) );
  XOR U10581 ( .A(n6452), .B(n6451), .Z(n6462) );
  XOR U10582 ( .A(n6454), .B(n6453), .Z(n6451) );
  XOR U10583 ( .A(y[3380]), .B(x[3380]), .Z(n6453) );
  XOR U10584 ( .A(y[3379]), .B(x[3379]), .Z(n6454) );
  XOR U10585 ( .A(y[3378]), .B(x[3378]), .Z(n6452) );
  XNOR U10586 ( .A(n6429), .B(n6428), .Z(n6446) );
  XNOR U10587 ( .A(n6443), .B(n6444), .Z(n6428) );
  XOR U10588 ( .A(n6440), .B(n6439), .Z(n6444) );
  XOR U10589 ( .A(y[3375]), .B(x[3375]), .Z(n6439) );
  XOR U10590 ( .A(n6442), .B(n6441), .Z(n6440) );
  XOR U10591 ( .A(y[3377]), .B(x[3377]), .Z(n6441) );
  XOR U10592 ( .A(y[3376]), .B(x[3376]), .Z(n6442) );
  XOR U10593 ( .A(n6434), .B(n6433), .Z(n6443) );
  XOR U10594 ( .A(n6436), .B(n6435), .Z(n6433) );
  XOR U10595 ( .A(y[3374]), .B(x[3374]), .Z(n6435) );
  XOR U10596 ( .A(y[3373]), .B(x[3373]), .Z(n6436) );
  XOR U10597 ( .A(y[3372]), .B(x[3372]), .Z(n6434) );
  XNOR U10598 ( .A(n6427), .B(n6426), .Z(n6429) );
  XNOR U10599 ( .A(n6423), .B(n6422), .Z(n6426) );
  XOR U10600 ( .A(n6425), .B(n6424), .Z(n6422) );
  XOR U10601 ( .A(y[3371]), .B(x[3371]), .Z(n6424) );
  XOR U10602 ( .A(y[3370]), .B(x[3370]), .Z(n6425) );
  XOR U10603 ( .A(y[3369]), .B(x[3369]), .Z(n6423) );
  XOR U10604 ( .A(n6417), .B(n6416), .Z(n6427) );
  XOR U10605 ( .A(n6419), .B(n6418), .Z(n6416) );
  XOR U10606 ( .A(y[3368]), .B(x[3368]), .Z(n6418) );
  XOR U10607 ( .A(y[3367]), .B(x[3367]), .Z(n6419) );
  XOR U10608 ( .A(y[3366]), .B(x[3366]), .Z(n6417) );
  NAND U10609 ( .A(n6480), .B(n6481), .Z(N29613) );
  NAND U10610 ( .A(n6482), .B(n6483), .Z(n6481) );
  NANDN U10611 ( .A(n6484), .B(n6485), .Z(n6483) );
  NANDN U10612 ( .A(n6485), .B(n6484), .Z(n6480) );
  XOR U10613 ( .A(n6484), .B(n6486), .Z(N29612) );
  XNOR U10614 ( .A(n6482), .B(n6485), .Z(n6486) );
  NAND U10615 ( .A(n6487), .B(n6488), .Z(n6485) );
  NAND U10616 ( .A(n6489), .B(n6490), .Z(n6488) );
  NANDN U10617 ( .A(n6491), .B(n6492), .Z(n6490) );
  NANDN U10618 ( .A(n6492), .B(n6491), .Z(n6487) );
  AND U10619 ( .A(n6493), .B(n6494), .Z(n6482) );
  NAND U10620 ( .A(n6495), .B(n6496), .Z(n6494) );
  OR U10621 ( .A(n6497), .B(n6498), .Z(n6496) );
  NAND U10622 ( .A(n6498), .B(n6497), .Z(n6493) );
  IV U10623 ( .A(n6499), .Z(n6498) );
  AND U10624 ( .A(n6500), .B(n6501), .Z(n6484) );
  NAND U10625 ( .A(n6502), .B(n6503), .Z(n6501) );
  NANDN U10626 ( .A(n6504), .B(n6505), .Z(n6503) );
  NANDN U10627 ( .A(n6505), .B(n6504), .Z(n6500) );
  XOR U10628 ( .A(n6497), .B(n6506), .Z(N29611) );
  XOR U10629 ( .A(n6495), .B(n6499), .Z(n6506) );
  XNOR U10630 ( .A(n6492), .B(n6507), .Z(n6499) );
  XNOR U10631 ( .A(n6489), .B(n6491), .Z(n6507) );
  AND U10632 ( .A(n6508), .B(n6509), .Z(n6491) );
  NANDN U10633 ( .A(n6510), .B(n6511), .Z(n6509) );
  NANDN U10634 ( .A(n6512), .B(n6513), .Z(n6511) );
  IV U10635 ( .A(n6514), .Z(n6513) );
  NAND U10636 ( .A(n6514), .B(n6512), .Z(n6508) );
  AND U10637 ( .A(n6515), .B(n6516), .Z(n6489) );
  NAND U10638 ( .A(n6517), .B(n6518), .Z(n6516) );
  OR U10639 ( .A(n6519), .B(n6520), .Z(n6518) );
  NAND U10640 ( .A(n6520), .B(n6519), .Z(n6515) );
  IV U10641 ( .A(n6521), .Z(n6520) );
  NAND U10642 ( .A(n6522), .B(n6523), .Z(n6492) );
  NANDN U10643 ( .A(n6524), .B(n6525), .Z(n6523) );
  NAND U10644 ( .A(n6526), .B(n6527), .Z(n6525) );
  OR U10645 ( .A(n6527), .B(n6526), .Z(n6522) );
  IV U10646 ( .A(n6528), .Z(n6526) );
  AND U10647 ( .A(n6529), .B(n6530), .Z(n6495) );
  NAND U10648 ( .A(n6531), .B(n6532), .Z(n6530) );
  NANDN U10649 ( .A(n6533), .B(n6534), .Z(n6532) );
  NANDN U10650 ( .A(n6534), .B(n6533), .Z(n6529) );
  XOR U10651 ( .A(n6505), .B(n6535), .Z(n6497) );
  XNOR U10652 ( .A(n6502), .B(n6504), .Z(n6535) );
  AND U10653 ( .A(n6536), .B(n6537), .Z(n6504) );
  NANDN U10654 ( .A(n6538), .B(n6539), .Z(n6537) );
  NANDN U10655 ( .A(n6540), .B(n6541), .Z(n6539) );
  IV U10656 ( .A(n6542), .Z(n6541) );
  NAND U10657 ( .A(n6542), .B(n6540), .Z(n6536) );
  AND U10658 ( .A(n6543), .B(n6544), .Z(n6502) );
  NAND U10659 ( .A(n6545), .B(n6546), .Z(n6544) );
  OR U10660 ( .A(n6547), .B(n6548), .Z(n6546) );
  NAND U10661 ( .A(n6548), .B(n6547), .Z(n6543) );
  IV U10662 ( .A(n6549), .Z(n6548) );
  NAND U10663 ( .A(n6550), .B(n6551), .Z(n6505) );
  NANDN U10664 ( .A(n6552), .B(n6553), .Z(n6551) );
  NAND U10665 ( .A(n6554), .B(n6555), .Z(n6553) );
  OR U10666 ( .A(n6555), .B(n6554), .Z(n6550) );
  IV U10667 ( .A(n6556), .Z(n6554) );
  XOR U10668 ( .A(n6531), .B(n6557), .Z(N29610) );
  XNOR U10669 ( .A(n6534), .B(n6533), .Z(n6557) );
  XNOR U10670 ( .A(n6545), .B(n6558), .Z(n6533) );
  XOR U10671 ( .A(n6549), .B(n6547), .Z(n6558) );
  XOR U10672 ( .A(n6555), .B(n6559), .Z(n6547) );
  XOR U10673 ( .A(n6552), .B(n6556), .Z(n6559) );
  NAND U10674 ( .A(n6560), .B(n6561), .Z(n6556) );
  NAND U10675 ( .A(n6562), .B(n6563), .Z(n6561) );
  NAND U10676 ( .A(n6564), .B(n6565), .Z(n6560) );
  AND U10677 ( .A(n6566), .B(n6567), .Z(n6552) );
  NAND U10678 ( .A(n6568), .B(n6569), .Z(n6567) );
  NAND U10679 ( .A(n6570), .B(n6571), .Z(n6566) );
  NANDN U10680 ( .A(n6572), .B(n6573), .Z(n6555) );
  NANDN U10681 ( .A(n6574), .B(n6575), .Z(n6549) );
  XNOR U10682 ( .A(n6540), .B(n6576), .Z(n6545) );
  XOR U10683 ( .A(n6538), .B(n6542), .Z(n6576) );
  NAND U10684 ( .A(n6577), .B(n6578), .Z(n6542) );
  NAND U10685 ( .A(n6579), .B(n6580), .Z(n6578) );
  NAND U10686 ( .A(n6581), .B(n6582), .Z(n6577) );
  AND U10687 ( .A(n6583), .B(n6584), .Z(n6538) );
  NAND U10688 ( .A(n6585), .B(n6586), .Z(n6584) );
  NAND U10689 ( .A(n6587), .B(n6588), .Z(n6583) );
  AND U10690 ( .A(n6589), .B(n6590), .Z(n6540) );
  NAND U10691 ( .A(n6591), .B(n6592), .Z(n6534) );
  XNOR U10692 ( .A(n6517), .B(n6593), .Z(n6531) );
  XOR U10693 ( .A(n6521), .B(n6519), .Z(n6593) );
  XOR U10694 ( .A(n6527), .B(n6594), .Z(n6519) );
  XOR U10695 ( .A(n6524), .B(n6528), .Z(n6594) );
  NAND U10696 ( .A(n6595), .B(n6596), .Z(n6528) );
  NAND U10697 ( .A(n6597), .B(n6598), .Z(n6596) );
  NAND U10698 ( .A(n6599), .B(n6600), .Z(n6595) );
  AND U10699 ( .A(n6601), .B(n6602), .Z(n6524) );
  NAND U10700 ( .A(n6603), .B(n6604), .Z(n6602) );
  NAND U10701 ( .A(n6605), .B(n6606), .Z(n6601) );
  NANDN U10702 ( .A(n6607), .B(n6608), .Z(n6527) );
  NANDN U10703 ( .A(n6609), .B(n6610), .Z(n6521) );
  XNOR U10704 ( .A(n6512), .B(n6611), .Z(n6517) );
  XOR U10705 ( .A(n6510), .B(n6514), .Z(n6611) );
  NAND U10706 ( .A(n6612), .B(n6613), .Z(n6514) );
  NAND U10707 ( .A(n6614), .B(n6615), .Z(n6613) );
  NAND U10708 ( .A(n6616), .B(n6617), .Z(n6612) );
  AND U10709 ( .A(n6618), .B(n6619), .Z(n6510) );
  NAND U10710 ( .A(n6620), .B(n6621), .Z(n6619) );
  NAND U10711 ( .A(n6622), .B(n6623), .Z(n6618) );
  AND U10712 ( .A(n6624), .B(n6625), .Z(n6512) );
  XOR U10713 ( .A(n6592), .B(n6591), .Z(N29609) );
  XNOR U10714 ( .A(n6610), .B(n6609), .Z(n6591) );
  XNOR U10715 ( .A(n6624), .B(n6625), .Z(n6609) );
  XOR U10716 ( .A(n6621), .B(n6620), .Z(n6625) );
  XOR U10717 ( .A(y[3363]), .B(x[3363]), .Z(n6620) );
  XOR U10718 ( .A(n6623), .B(n6622), .Z(n6621) );
  XOR U10719 ( .A(y[3365]), .B(x[3365]), .Z(n6622) );
  XOR U10720 ( .A(y[3364]), .B(x[3364]), .Z(n6623) );
  XOR U10721 ( .A(n6615), .B(n6614), .Z(n6624) );
  XOR U10722 ( .A(n6617), .B(n6616), .Z(n6614) );
  XOR U10723 ( .A(y[3362]), .B(x[3362]), .Z(n6616) );
  XOR U10724 ( .A(y[3361]), .B(x[3361]), .Z(n6617) );
  XOR U10725 ( .A(y[3360]), .B(x[3360]), .Z(n6615) );
  XNOR U10726 ( .A(n6608), .B(n6607), .Z(n6610) );
  XNOR U10727 ( .A(n6604), .B(n6603), .Z(n6607) );
  XOR U10728 ( .A(n6606), .B(n6605), .Z(n6603) );
  XOR U10729 ( .A(y[3359]), .B(x[3359]), .Z(n6605) );
  XOR U10730 ( .A(y[3358]), .B(x[3358]), .Z(n6606) );
  XOR U10731 ( .A(y[3357]), .B(x[3357]), .Z(n6604) );
  XOR U10732 ( .A(n6598), .B(n6597), .Z(n6608) );
  XOR U10733 ( .A(n6600), .B(n6599), .Z(n6597) );
  XOR U10734 ( .A(y[3356]), .B(x[3356]), .Z(n6599) );
  XOR U10735 ( .A(y[3355]), .B(x[3355]), .Z(n6600) );
  XOR U10736 ( .A(y[3354]), .B(x[3354]), .Z(n6598) );
  XNOR U10737 ( .A(n6575), .B(n6574), .Z(n6592) );
  XNOR U10738 ( .A(n6589), .B(n6590), .Z(n6574) );
  XOR U10739 ( .A(n6586), .B(n6585), .Z(n6590) );
  XOR U10740 ( .A(y[3351]), .B(x[3351]), .Z(n6585) );
  XOR U10741 ( .A(n6588), .B(n6587), .Z(n6586) );
  XOR U10742 ( .A(y[3353]), .B(x[3353]), .Z(n6587) );
  XOR U10743 ( .A(y[3352]), .B(x[3352]), .Z(n6588) );
  XOR U10744 ( .A(n6580), .B(n6579), .Z(n6589) );
  XOR U10745 ( .A(n6582), .B(n6581), .Z(n6579) );
  XOR U10746 ( .A(y[3350]), .B(x[3350]), .Z(n6581) );
  XOR U10747 ( .A(y[3349]), .B(x[3349]), .Z(n6582) );
  XOR U10748 ( .A(y[3348]), .B(x[3348]), .Z(n6580) );
  XNOR U10749 ( .A(n6573), .B(n6572), .Z(n6575) );
  XNOR U10750 ( .A(n6569), .B(n6568), .Z(n6572) );
  XOR U10751 ( .A(n6571), .B(n6570), .Z(n6568) );
  XOR U10752 ( .A(y[3347]), .B(x[3347]), .Z(n6570) );
  XOR U10753 ( .A(y[3346]), .B(x[3346]), .Z(n6571) );
  XOR U10754 ( .A(y[3345]), .B(x[3345]), .Z(n6569) );
  XOR U10755 ( .A(n6563), .B(n6562), .Z(n6573) );
  XOR U10756 ( .A(n6565), .B(n6564), .Z(n6562) );
  XOR U10757 ( .A(y[3344]), .B(x[3344]), .Z(n6564) );
  XOR U10758 ( .A(y[3343]), .B(x[3343]), .Z(n6565) );
  XOR U10759 ( .A(y[3342]), .B(x[3342]), .Z(n6563) );
  NAND U10760 ( .A(n6626), .B(n6627), .Z(N29601) );
  NAND U10761 ( .A(n6628), .B(n6629), .Z(n6627) );
  NANDN U10762 ( .A(n6630), .B(n6631), .Z(n6629) );
  NANDN U10763 ( .A(n6631), .B(n6630), .Z(n6626) );
  XOR U10764 ( .A(n6630), .B(n6632), .Z(N29600) );
  XNOR U10765 ( .A(n6628), .B(n6631), .Z(n6632) );
  NAND U10766 ( .A(n6633), .B(n6634), .Z(n6631) );
  NAND U10767 ( .A(n6635), .B(n6636), .Z(n6634) );
  NANDN U10768 ( .A(n6637), .B(n6638), .Z(n6636) );
  NANDN U10769 ( .A(n6638), .B(n6637), .Z(n6633) );
  AND U10770 ( .A(n6639), .B(n6640), .Z(n6628) );
  NAND U10771 ( .A(n6641), .B(n6642), .Z(n6640) );
  OR U10772 ( .A(n6643), .B(n6644), .Z(n6642) );
  NAND U10773 ( .A(n6644), .B(n6643), .Z(n6639) );
  IV U10774 ( .A(n6645), .Z(n6644) );
  AND U10775 ( .A(n6646), .B(n6647), .Z(n6630) );
  NAND U10776 ( .A(n6648), .B(n6649), .Z(n6647) );
  NANDN U10777 ( .A(n6650), .B(n6651), .Z(n6649) );
  NANDN U10778 ( .A(n6651), .B(n6650), .Z(n6646) );
  XOR U10779 ( .A(n6643), .B(n6652), .Z(N29599) );
  XOR U10780 ( .A(n6641), .B(n6645), .Z(n6652) );
  XNOR U10781 ( .A(n6638), .B(n6653), .Z(n6645) );
  XNOR U10782 ( .A(n6635), .B(n6637), .Z(n6653) );
  AND U10783 ( .A(n6654), .B(n6655), .Z(n6637) );
  NANDN U10784 ( .A(n6656), .B(n6657), .Z(n6655) );
  NANDN U10785 ( .A(n6658), .B(n6659), .Z(n6657) );
  IV U10786 ( .A(n6660), .Z(n6659) );
  NAND U10787 ( .A(n6660), .B(n6658), .Z(n6654) );
  AND U10788 ( .A(n6661), .B(n6662), .Z(n6635) );
  NAND U10789 ( .A(n6663), .B(n6664), .Z(n6662) );
  OR U10790 ( .A(n6665), .B(n6666), .Z(n6664) );
  NAND U10791 ( .A(n6666), .B(n6665), .Z(n6661) );
  IV U10792 ( .A(n6667), .Z(n6666) );
  NAND U10793 ( .A(n6668), .B(n6669), .Z(n6638) );
  NANDN U10794 ( .A(n6670), .B(n6671), .Z(n6669) );
  NAND U10795 ( .A(n6672), .B(n6673), .Z(n6671) );
  OR U10796 ( .A(n6673), .B(n6672), .Z(n6668) );
  IV U10797 ( .A(n6674), .Z(n6672) );
  AND U10798 ( .A(n6675), .B(n6676), .Z(n6641) );
  NAND U10799 ( .A(n6677), .B(n6678), .Z(n6676) );
  NANDN U10800 ( .A(n6679), .B(n6680), .Z(n6678) );
  NANDN U10801 ( .A(n6680), .B(n6679), .Z(n6675) );
  XOR U10802 ( .A(n6651), .B(n6681), .Z(n6643) );
  XNOR U10803 ( .A(n6648), .B(n6650), .Z(n6681) );
  AND U10804 ( .A(n6682), .B(n6683), .Z(n6650) );
  NANDN U10805 ( .A(n6684), .B(n6685), .Z(n6683) );
  NANDN U10806 ( .A(n6686), .B(n6687), .Z(n6685) );
  IV U10807 ( .A(n6688), .Z(n6687) );
  NAND U10808 ( .A(n6688), .B(n6686), .Z(n6682) );
  AND U10809 ( .A(n6689), .B(n6690), .Z(n6648) );
  NAND U10810 ( .A(n6691), .B(n6692), .Z(n6690) );
  OR U10811 ( .A(n6693), .B(n6694), .Z(n6692) );
  NAND U10812 ( .A(n6694), .B(n6693), .Z(n6689) );
  IV U10813 ( .A(n6695), .Z(n6694) );
  NAND U10814 ( .A(n6696), .B(n6697), .Z(n6651) );
  NANDN U10815 ( .A(n6698), .B(n6699), .Z(n6697) );
  NAND U10816 ( .A(n6700), .B(n6701), .Z(n6699) );
  OR U10817 ( .A(n6701), .B(n6700), .Z(n6696) );
  IV U10818 ( .A(n6702), .Z(n6700) );
  XOR U10819 ( .A(n6677), .B(n6703), .Z(N29598) );
  XNOR U10820 ( .A(n6680), .B(n6679), .Z(n6703) );
  XNOR U10821 ( .A(n6691), .B(n6704), .Z(n6679) );
  XOR U10822 ( .A(n6695), .B(n6693), .Z(n6704) );
  XOR U10823 ( .A(n6701), .B(n6705), .Z(n6693) );
  XOR U10824 ( .A(n6698), .B(n6702), .Z(n6705) );
  NAND U10825 ( .A(n6706), .B(n6707), .Z(n6702) );
  NAND U10826 ( .A(n6708), .B(n6709), .Z(n6707) );
  NAND U10827 ( .A(n6710), .B(n6711), .Z(n6706) );
  AND U10828 ( .A(n6712), .B(n6713), .Z(n6698) );
  NAND U10829 ( .A(n6714), .B(n6715), .Z(n6713) );
  NAND U10830 ( .A(n6716), .B(n6717), .Z(n6712) );
  NANDN U10831 ( .A(n6718), .B(n6719), .Z(n6701) );
  NANDN U10832 ( .A(n6720), .B(n6721), .Z(n6695) );
  XNOR U10833 ( .A(n6686), .B(n6722), .Z(n6691) );
  XOR U10834 ( .A(n6684), .B(n6688), .Z(n6722) );
  NAND U10835 ( .A(n6723), .B(n6724), .Z(n6688) );
  NAND U10836 ( .A(n6725), .B(n6726), .Z(n6724) );
  NAND U10837 ( .A(n6727), .B(n6728), .Z(n6723) );
  AND U10838 ( .A(n6729), .B(n6730), .Z(n6684) );
  NAND U10839 ( .A(n6731), .B(n6732), .Z(n6730) );
  NAND U10840 ( .A(n6733), .B(n6734), .Z(n6729) );
  AND U10841 ( .A(n6735), .B(n6736), .Z(n6686) );
  NAND U10842 ( .A(n6737), .B(n6738), .Z(n6680) );
  XNOR U10843 ( .A(n6663), .B(n6739), .Z(n6677) );
  XOR U10844 ( .A(n6667), .B(n6665), .Z(n6739) );
  XOR U10845 ( .A(n6673), .B(n6740), .Z(n6665) );
  XOR U10846 ( .A(n6670), .B(n6674), .Z(n6740) );
  NAND U10847 ( .A(n6741), .B(n6742), .Z(n6674) );
  NAND U10848 ( .A(n6743), .B(n6744), .Z(n6742) );
  NAND U10849 ( .A(n6745), .B(n6746), .Z(n6741) );
  AND U10850 ( .A(n6747), .B(n6748), .Z(n6670) );
  NAND U10851 ( .A(n6749), .B(n6750), .Z(n6748) );
  NAND U10852 ( .A(n6751), .B(n6752), .Z(n6747) );
  NANDN U10853 ( .A(n6753), .B(n6754), .Z(n6673) );
  NANDN U10854 ( .A(n6755), .B(n6756), .Z(n6667) );
  XNOR U10855 ( .A(n6658), .B(n6757), .Z(n6663) );
  XOR U10856 ( .A(n6656), .B(n6660), .Z(n6757) );
  NAND U10857 ( .A(n6758), .B(n6759), .Z(n6660) );
  NAND U10858 ( .A(n6760), .B(n6761), .Z(n6759) );
  NAND U10859 ( .A(n6762), .B(n6763), .Z(n6758) );
  AND U10860 ( .A(n6764), .B(n6765), .Z(n6656) );
  NAND U10861 ( .A(n6766), .B(n6767), .Z(n6765) );
  NAND U10862 ( .A(n6768), .B(n6769), .Z(n6764) );
  AND U10863 ( .A(n6770), .B(n6771), .Z(n6658) );
  XOR U10864 ( .A(n6738), .B(n6737), .Z(N29597) );
  XNOR U10865 ( .A(n6756), .B(n6755), .Z(n6737) );
  XNOR U10866 ( .A(n6770), .B(n6771), .Z(n6755) );
  XOR U10867 ( .A(n6767), .B(n6766), .Z(n6771) );
  XOR U10868 ( .A(y[3339]), .B(x[3339]), .Z(n6766) );
  XOR U10869 ( .A(n6769), .B(n6768), .Z(n6767) );
  XOR U10870 ( .A(y[3341]), .B(x[3341]), .Z(n6768) );
  XOR U10871 ( .A(y[3340]), .B(x[3340]), .Z(n6769) );
  XOR U10872 ( .A(n6761), .B(n6760), .Z(n6770) );
  XOR U10873 ( .A(n6763), .B(n6762), .Z(n6760) );
  XOR U10874 ( .A(y[3338]), .B(x[3338]), .Z(n6762) );
  XOR U10875 ( .A(y[3337]), .B(x[3337]), .Z(n6763) );
  XOR U10876 ( .A(y[3336]), .B(x[3336]), .Z(n6761) );
  XNOR U10877 ( .A(n6754), .B(n6753), .Z(n6756) );
  XNOR U10878 ( .A(n6750), .B(n6749), .Z(n6753) );
  XOR U10879 ( .A(n6752), .B(n6751), .Z(n6749) );
  XOR U10880 ( .A(y[3335]), .B(x[3335]), .Z(n6751) );
  XOR U10881 ( .A(y[3334]), .B(x[3334]), .Z(n6752) );
  XOR U10882 ( .A(y[3333]), .B(x[3333]), .Z(n6750) );
  XOR U10883 ( .A(n6744), .B(n6743), .Z(n6754) );
  XOR U10884 ( .A(n6746), .B(n6745), .Z(n6743) );
  XOR U10885 ( .A(y[3332]), .B(x[3332]), .Z(n6745) );
  XOR U10886 ( .A(y[3331]), .B(x[3331]), .Z(n6746) );
  XOR U10887 ( .A(y[3330]), .B(x[3330]), .Z(n6744) );
  XNOR U10888 ( .A(n6721), .B(n6720), .Z(n6738) );
  XNOR U10889 ( .A(n6735), .B(n6736), .Z(n6720) );
  XOR U10890 ( .A(n6732), .B(n6731), .Z(n6736) );
  XOR U10891 ( .A(y[3327]), .B(x[3327]), .Z(n6731) );
  XOR U10892 ( .A(n6734), .B(n6733), .Z(n6732) );
  XOR U10893 ( .A(y[3329]), .B(x[3329]), .Z(n6733) );
  XOR U10894 ( .A(y[3328]), .B(x[3328]), .Z(n6734) );
  XOR U10895 ( .A(n6726), .B(n6725), .Z(n6735) );
  XOR U10896 ( .A(n6728), .B(n6727), .Z(n6725) );
  XOR U10897 ( .A(y[3326]), .B(x[3326]), .Z(n6727) );
  XOR U10898 ( .A(y[3325]), .B(x[3325]), .Z(n6728) );
  XOR U10899 ( .A(y[3324]), .B(x[3324]), .Z(n6726) );
  XNOR U10900 ( .A(n6719), .B(n6718), .Z(n6721) );
  XNOR U10901 ( .A(n6715), .B(n6714), .Z(n6718) );
  XOR U10902 ( .A(n6717), .B(n6716), .Z(n6714) );
  XOR U10903 ( .A(y[3323]), .B(x[3323]), .Z(n6716) );
  XOR U10904 ( .A(y[3322]), .B(x[3322]), .Z(n6717) );
  XOR U10905 ( .A(y[3321]), .B(x[3321]), .Z(n6715) );
  XOR U10906 ( .A(n6709), .B(n6708), .Z(n6719) );
  XOR U10907 ( .A(n6711), .B(n6710), .Z(n6708) );
  XOR U10908 ( .A(y[3320]), .B(x[3320]), .Z(n6710) );
  XOR U10909 ( .A(y[3319]), .B(x[3319]), .Z(n6711) );
  XOR U10910 ( .A(y[3318]), .B(x[3318]), .Z(n6709) );
  NAND U10911 ( .A(n6772), .B(n6773), .Z(N29589) );
  NAND U10912 ( .A(n6774), .B(n6775), .Z(n6773) );
  NANDN U10913 ( .A(n6776), .B(n6777), .Z(n6775) );
  NANDN U10914 ( .A(n6777), .B(n6776), .Z(n6772) );
  XOR U10915 ( .A(n6776), .B(n6778), .Z(N29588) );
  XNOR U10916 ( .A(n6774), .B(n6777), .Z(n6778) );
  NAND U10917 ( .A(n6779), .B(n6780), .Z(n6777) );
  NAND U10918 ( .A(n6781), .B(n6782), .Z(n6780) );
  NANDN U10919 ( .A(n6783), .B(n6784), .Z(n6782) );
  NANDN U10920 ( .A(n6784), .B(n6783), .Z(n6779) );
  AND U10921 ( .A(n6785), .B(n6786), .Z(n6774) );
  NAND U10922 ( .A(n6787), .B(n6788), .Z(n6786) );
  OR U10923 ( .A(n6789), .B(n6790), .Z(n6788) );
  NAND U10924 ( .A(n6790), .B(n6789), .Z(n6785) );
  IV U10925 ( .A(n6791), .Z(n6790) );
  AND U10926 ( .A(n6792), .B(n6793), .Z(n6776) );
  NAND U10927 ( .A(n6794), .B(n6795), .Z(n6793) );
  NANDN U10928 ( .A(n6796), .B(n6797), .Z(n6795) );
  NANDN U10929 ( .A(n6797), .B(n6796), .Z(n6792) );
  XOR U10930 ( .A(n6789), .B(n6798), .Z(N29587) );
  XOR U10931 ( .A(n6787), .B(n6791), .Z(n6798) );
  XNOR U10932 ( .A(n6784), .B(n6799), .Z(n6791) );
  XNOR U10933 ( .A(n6781), .B(n6783), .Z(n6799) );
  AND U10934 ( .A(n6800), .B(n6801), .Z(n6783) );
  NANDN U10935 ( .A(n6802), .B(n6803), .Z(n6801) );
  NANDN U10936 ( .A(n6804), .B(n6805), .Z(n6803) );
  IV U10937 ( .A(n6806), .Z(n6805) );
  NAND U10938 ( .A(n6806), .B(n6804), .Z(n6800) );
  AND U10939 ( .A(n6807), .B(n6808), .Z(n6781) );
  NAND U10940 ( .A(n6809), .B(n6810), .Z(n6808) );
  OR U10941 ( .A(n6811), .B(n6812), .Z(n6810) );
  NAND U10942 ( .A(n6812), .B(n6811), .Z(n6807) );
  IV U10943 ( .A(n6813), .Z(n6812) );
  NAND U10944 ( .A(n6814), .B(n6815), .Z(n6784) );
  NANDN U10945 ( .A(n6816), .B(n6817), .Z(n6815) );
  NAND U10946 ( .A(n6818), .B(n6819), .Z(n6817) );
  OR U10947 ( .A(n6819), .B(n6818), .Z(n6814) );
  IV U10948 ( .A(n6820), .Z(n6818) );
  AND U10949 ( .A(n6821), .B(n6822), .Z(n6787) );
  NAND U10950 ( .A(n6823), .B(n6824), .Z(n6822) );
  NANDN U10951 ( .A(n6825), .B(n6826), .Z(n6824) );
  NANDN U10952 ( .A(n6826), .B(n6825), .Z(n6821) );
  XOR U10953 ( .A(n6797), .B(n6827), .Z(n6789) );
  XNOR U10954 ( .A(n6794), .B(n6796), .Z(n6827) );
  AND U10955 ( .A(n6828), .B(n6829), .Z(n6796) );
  NANDN U10956 ( .A(n6830), .B(n6831), .Z(n6829) );
  NANDN U10957 ( .A(n6832), .B(n6833), .Z(n6831) );
  IV U10958 ( .A(n6834), .Z(n6833) );
  NAND U10959 ( .A(n6834), .B(n6832), .Z(n6828) );
  AND U10960 ( .A(n6835), .B(n6836), .Z(n6794) );
  NAND U10961 ( .A(n6837), .B(n6838), .Z(n6836) );
  OR U10962 ( .A(n6839), .B(n6840), .Z(n6838) );
  NAND U10963 ( .A(n6840), .B(n6839), .Z(n6835) );
  IV U10964 ( .A(n6841), .Z(n6840) );
  NAND U10965 ( .A(n6842), .B(n6843), .Z(n6797) );
  NANDN U10966 ( .A(n6844), .B(n6845), .Z(n6843) );
  NAND U10967 ( .A(n6846), .B(n6847), .Z(n6845) );
  OR U10968 ( .A(n6847), .B(n6846), .Z(n6842) );
  IV U10969 ( .A(n6848), .Z(n6846) );
  XOR U10970 ( .A(n6823), .B(n6849), .Z(N29586) );
  XNOR U10971 ( .A(n6826), .B(n6825), .Z(n6849) );
  XNOR U10972 ( .A(n6837), .B(n6850), .Z(n6825) );
  XOR U10973 ( .A(n6841), .B(n6839), .Z(n6850) );
  XOR U10974 ( .A(n6847), .B(n6851), .Z(n6839) );
  XOR U10975 ( .A(n6844), .B(n6848), .Z(n6851) );
  NAND U10976 ( .A(n6852), .B(n6853), .Z(n6848) );
  NAND U10977 ( .A(n6854), .B(n6855), .Z(n6853) );
  NAND U10978 ( .A(n6856), .B(n6857), .Z(n6852) );
  AND U10979 ( .A(n6858), .B(n6859), .Z(n6844) );
  NAND U10980 ( .A(n6860), .B(n6861), .Z(n6859) );
  NAND U10981 ( .A(n6862), .B(n6863), .Z(n6858) );
  NANDN U10982 ( .A(n6864), .B(n6865), .Z(n6847) );
  NANDN U10983 ( .A(n6866), .B(n6867), .Z(n6841) );
  XNOR U10984 ( .A(n6832), .B(n6868), .Z(n6837) );
  XOR U10985 ( .A(n6830), .B(n6834), .Z(n6868) );
  NAND U10986 ( .A(n6869), .B(n6870), .Z(n6834) );
  NAND U10987 ( .A(n6871), .B(n6872), .Z(n6870) );
  NAND U10988 ( .A(n6873), .B(n6874), .Z(n6869) );
  AND U10989 ( .A(n6875), .B(n6876), .Z(n6830) );
  NAND U10990 ( .A(n6877), .B(n6878), .Z(n6876) );
  NAND U10991 ( .A(n6879), .B(n6880), .Z(n6875) );
  AND U10992 ( .A(n6881), .B(n6882), .Z(n6832) );
  NAND U10993 ( .A(n6883), .B(n6884), .Z(n6826) );
  XNOR U10994 ( .A(n6809), .B(n6885), .Z(n6823) );
  XOR U10995 ( .A(n6813), .B(n6811), .Z(n6885) );
  XOR U10996 ( .A(n6819), .B(n6886), .Z(n6811) );
  XOR U10997 ( .A(n6816), .B(n6820), .Z(n6886) );
  NAND U10998 ( .A(n6887), .B(n6888), .Z(n6820) );
  NAND U10999 ( .A(n6889), .B(n6890), .Z(n6888) );
  NAND U11000 ( .A(n6891), .B(n6892), .Z(n6887) );
  AND U11001 ( .A(n6893), .B(n6894), .Z(n6816) );
  NAND U11002 ( .A(n6895), .B(n6896), .Z(n6894) );
  NAND U11003 ( .A(n6897), .B(n6898), .Z(n6893) );
  NANDN U11004 ( .A(n6899), .B(n6900), .Z(n6819) );
  NANDN U11005 ( .A(n6901), .B(n6902), .Z(n6813) );
  XNOR U11006 ( .A(n6804), .B(n6903), .Z(n6809) );
  XOR U11007 ( .A(n6802), .B(n6806), .Z(n6903) );
  NAND U11008 ( .A(n6904), .B(n6905), .Z(n6806) );
  NAND U11009 ( .A(n6906), .B(n6907), .Z(n6905) );
  NAND U11010 ( .A(n6908), .B(n6909), .Z(n6904) );
  AND U11011 ( .A(n6910), .B(n6911), .Z(n6802) );
  NAND U11012 ( .A(n6912), .B(n6913), .Z(n6911) );
  NAND U11013 ( .A(n6914), .B(n6915), .Z(n6910) );
  AND U11014 ( .A(n6916), .B(n6917), .Z(n6804) );
  XOR U11015 ( .A(n6884), .B(n6883), .Z(N29585) );
  XNOR U11016 ( .A(n6902), .B(n6901), .Z(n6883) );
  XNOR U11017 ( .A(n6916), .B(n6917), .Z(n6901) );
  XOR U11018 ( .A(n6913), .B(n6912), .Z(n6917) );
  XOR U11019 ( .A(y[3315]), .B(x[3315]), .Z(n6912) );
  XOR U11020 ( .A(n6915), .B(n6914), .Z(n6913) );
  XOR U11021 ( .A(y[3317]), .B(x[3317]), .Z(n6914) );
  XOR U11022 ( .A(y[3316]), .B(x[3316]), .Z(n6915) );
  XOR U11023 ( .A(n6907), .B(n6906), .Z(n6916) );
  XOR U11024 ( .A(n6909), .B(n6908), .Z(n6906) );
  XOR U11025 ( .A(y[3314]), .B(x[3314]), .Z(n6908) );
  XOR U11026 ( .A(y[3313]), .B(x[3313]), .Z(n6909) );
  XOR U11027 ( .A(y[3312]), .B(x[3312]), .Z(n6907) );
  XNOR U11028 ( .A(n6900), .B(n6899), .Z(n6902) );
  XNOR U11029 ( .A(n6896), .B(n6895), .Z(n6899) );
  XOR U11030 ( .A(n6898), .B(n6897), .Z(n6895) );
  XOR U11031 ( .A(y[3311]), .B(x[3311]), .Z(n6897) );
  XOR U11032 ( .A(y[3310]), .B(x[3310]), .Z(n6898) );
  XOR U11033 ( .A(y[3309]), .B(x[3309]), .Z(n6896) );
  XOR U11034 ( .A(n6890), .B(n6889), .Z(n6900) );
  XOR U11035 ( .A(n6892), .B(n6891), .Z(n6889) );
  XOR U11036 ( .A(y[3308]), .B(x[3308]), .Z(n6891) );
  XOR U11037 ( .A(y[3307]), .B(x[3307]), .Z(n6892) );
  XOR U11038 ( .A(y[3306]), .B(x[3306]), .Z(n6890) );
  XNOR U11039 ( .A(n6867), .B(n6866), .Z(n6884) );
  XNOR U11040 ( .A(n6881), .B(n6882), .Z(n6866) );
  XOR U11041 ( .A(n6878), .B(n6877), .Z(n6882) );
  XOR U11042 ( .A(y[3303]), .B(x[3303]), .Z(n6877) );
  XOR U11043 ( .A(n6880), .B(n6879), .Z(n6878) );
  XOR U11044 ( .A(y[3305]), .B(x[3305]), .Z(n6879) );
  XOR U11045 ( .A(y[3304]), .B(x[3304]), .Z(n6880) );
  XOR U11046 ( .A(n6872), .B(n6871), .Z(n6881) );
  XOR U11047 ( .A(n6874), .B(n6873), .Z(n6871) );
  XOR U11048 ( .A(y[3302]), .B(x[3302]), .Z(n6873) );
  XOR U11049 ( .A(y[3301]), .B(x[3301]), .Z(n6874) );
  XOR U11050 ( .A(y[3300]), .B(x[3300]), .Z(n6872) );
  XNOR U11051 ( .A(n6865), .B(n6864), .Z(n6867) );
  XNOR U11052 ( .A(n6861), .B(n6860), .Z(n6864) );
  XOR U11053 ( .A(n6863), .B(n6862), .Z(n6860) );
  XOR U11054 ( .A(y[3299]), .B(x[3299]), .Z(n6862) );
  XOR U11055 ( .A(y[3298]), .B(x[3298]), .Z(n6863) );
  XOR U11056 ( .A(y[3297]), .B(x[3297]), .Z(n6861) );
  XOR U11057 ( .A(n6855), .B(n6854), .Z(n6865) );
  XOR U11058 ( .A(n6857), .B(n6856), .Z(n6854) );
  XOR U11059 ( .A(y[3296]), .B(x[3296]), .Z(n6856) );
  XOR U11060 ( .A(y[3295]), .B(x[3295]), .Z(n6857) );
  XOR U11061 ( .A(y[3294]), .B(x[3294]), .Z(n6855) );
  NAND U11062 ( .A(n6918), .B(n6919), .Z(N29577) );
  NAND U11063 ( .A(n6920), .B(n6921), .Z(n6919) );
  NANDN U11064 ( .A(n6922), .B(n6923), .Z(n6921) );
  NANDN U11065 ( .A(n6923), .B(n6922), .Z(n6918) );
  XOR U11066 ( .A(n6922), .B(n6924), .Z(N29576) );
  XNOR U11067 ( .A(n6920), .B(n6923), .Z(n6924) );
  NAND U11068 ( .A(n6925), .B(n6926), .Z(n6923) );
  NAND U11069 ( .A(n6927), .B(n6928), .Z(n6926) );
  NANDN U11070 ( .A(n6929), .B(n6930), .Z(n6928) );
  NANDN U11071 ( .A(n6930), .B(n6929), .Z(n6925) );
  AND U11072 ( .A(n6931), .B(n6932), .Z(n6920) );
  NAND U11073 ( .A(n6933), .B(n6934), .Z(n6932) );
  OR U11074 ( .A(n6935), .B(n6936), .Z(n6934) );
  NAND U11075 ( .A(n6936), .B(n6935), .Z(n6931) );
  IV U11076 ( .A(n6937), .Z(n6936) );
  AND U11077 ( .A(n6938), .B(n6939), .Z(n6922) );
  NAND U11078 ( .A(n6940), .B(n6941), .Z(n6939) );
  NANDN U11079 ( .A(n6942), .B(n6943), .Z(n6941) );
  NANDN U11080 ( .A(n6943), .B(n6942), .Z(n6938) );
  XOR U11081 ( .A(n6935), .B(n6944), .Z(N29575) );
  XOR U11082 ( .A(n6933), .B(n6937), .Z(n6944) );
  XNOR U11083 ( .A(n6930), .B(n6945), .Z(n6937) );
  XNOR U11084 ( .A(n6927), .B(n6929), .Z(n6945) );
  AND U11085 ( .A(n6946), .B(n6947), .Z(n6929) );
  NANDN U11086 ( .A(n6948), .B(n6949), .Z(n6947) );
  NANDN U11087 ( .A(n6950), .B(n6951), .Z(n6949) );
  IV U11088 ( .A(n6952), .Z(n6951) );
  NAND U11089 ( .A(n6952), .B(n6950), .Z(n6946) );
  AND U11090 ( .A(n6953), .B(n6954), .Z(n6927) );
  NAND U11091 ( .A(n6955), .B(n6956), .Z(n6954) );
  OR U11092 ( .A(n6957), .B(n6958), .Z(n6956) );
  NAND U11093 ( .A(n6958), .B(n6957), .Z(n6953) );
  IV U11094 ( .A(n6959), .Z(n6958) );
  NAND U11095 ( .A(n6960), .B(n6961), .Z(n6930) );
  NANDN U11096 ( .A(n6962), .B(n6963), .Z(n6961) );
  NAND U11097 ( .A(n6964), .B(n6965), .Z(n6963) );
  OR U11098 ( .A(n6965), .B(n6964), .Z(n6960) );
  IV U11099 ( .A(n6966), .Z(n6964) );
  AND U11100 ( .A(n6967), .B(n6968), .Z(n6933) );
  NAND U11101 ( .A(n6969), .B(n6970), .Z(n6968) );
  NANDN U11102 ( .A(n6971), .B(n6972), .Z(n6970) );
  NANDN U11103 ( .A(n6972), .B(n6971), .Z(n6967) );
  XOR U11104 ( .A(n6943), .B(n6973), .Z(n6935) );
  XNOR U11105 ( .A(n6940), .B(n6942), .Z(n6973) );
  AND U11106 ( .A(n6974), .B(n6975), .Z(n6942) );
  NANDN U11107 ( .A(n6976), .B(n6977), .Z(n6975) );
  NANDN U11108 ( .A(n6978), .B(n6979), .Z(n6977) );
  IV U11109 ( .A(n6980), .Z(n6979) );
  NAND U11110 ( .A(n6980), .B(n6978), .Z(n6974) );
  AND U11111 ( .A(n6981), .B(n6982), .Z(n6940) );
  NAND U11112 ( .A(n6983), .B(n6984), .Z(n6982) );
  OR U11113 ( .A(n6985), .B(n6986), .Z(n6984) );
  NAND U11114 ( .A(n6986), .B(n6985), .Z(n6981) );
  IV U11115 ( .A(n6987), .Z(n6986) );
  NAND U11116 ( .A(n6988), .B(n6989), .Z(n6943) );
  NANDN U11117 ( .A(n6990), .B(n6991), .Z(n6989) );
  NAND U11118 ( .A(n6992), .B(n6993), .Z(n6991) );
  OR U11119 ( .A(n6993), .B(n6992), .Z(n6988) );
  IV U11120 ( .A(n6994), .Z(n6992) );
  XOR U11121 ( .A(n6969), .B(n6995), .Z(N29574) );
  XNOR U11122 ( .A(n6972), .B(n6971), .Z(n6995) );
  XNOR U11123 ( .A(n6983), .B(n6996), .Z(n6971) );
  XOR U11124 ( .A(n6987), .B(n6985), .Z(n6996) );
  XOR U11125 ( .A(n6993), .B(n6997), .Z(n6985) );
  XOR U11126 ( .A(n6990), .B(n6994), .Z(n6997) );
  NAND U11127 ( .A(n6998), .B(n6999), .Z(n6994) );
  NAND U11128 ( .A(n7000), .B(n7001), .Z(n6999) );
  NAND U11129 ( .A(n7002), .B(n7003), .Z(n6998) );
  AND U11130 ( .A(n7004), .B(n7005), .Z(n6990) );
  NAND U11131 ( .A(n7006), .B(n7007), .Z(n7005) );
  NAND U11132 ( .A(n7008), .B(n7009), .Z(n7004) );
  NANDN U11133 ( .A(n7010), .B(n7011), .Z(n6993) );
  NANDN U11134 ( .A(n7012), .B(n7013), .Z(n6987) );
  XNOR U11135 ( .A(n6978), .B(n7014), .Z(n6983) );
  XOR U11136 ( .A(n6976), .B(n6980), .Z(n7014) );
  NAND U11137 ( .A(n7015), .B(n7016), .Z(n6980) );
  NAND U11138 ( .A(n7017), .B(n7018), .Z(n7016) );
  NAND U11139 ( .A(n7019), .B(n7020), .Z(n7015) );
  AND U11140 ( .A(n7021), .B(n7022), .Z(n6976) );
  NAND U11141 ( .A(n7023), .B(n7024), .Z(n7022) );
  NAND U11142 ( .A(n7025), .B(n7026), .Z(n7021) );
  AND U11143 ( .A(n7027), .B(n7028), .Z(n6978) );
  NAND U11144 ( .A(n7029), .B(n7030), .Z(n6972) );
  XNOR U11145 ( .A(n6955), .B(n7031), .Z(n6969) );
  XOR U11146 ( .A(n6959), .B(n6957), .Z(n7031) );
  XOR U11147 ( .A(n6965), .B(n7032), .Z(n6957) );
  XOR U11148 ( .A(n6962), .B(n6966), .Z(n7032) );
  NAND U11149 ( .A(n7033), .B(n7034), .Z(n6966) );
  NAND U11150 ( .A(n7035), .B(n7036), .Z(n7034) );
  NAND U11151 ( .A(n7037), .B(n7038), .Z(n7033) );
  AND U11152 ( .A(n7039), .B(n7040), .Z(n6962) );
  NAND U11153 ( .A(n7041), .B(n7042), .Z(n7040) );
  NAND U11154 ( .A(n7043), .B(n7044), .Z(n7039) );
  NANDN U11155 ( .A(n7045), .B(n7046), .Z(n6965) );
  NANDN U11156 ( .A(n7047), .B(n7048), .Z(n6959) );
  XNOR U11157 ( .A(n6950), .B(n7049), .Z(n6955) );
  XOR U11158 ( .A(n6948), .B(n6952), .Z(n7049) );
  NAND U11159 ( .A(n7050), .B(n7051), .Z(n6952) );
  NAND U11160 ( .A(n7052), .B(n7053), .Z(n7051) );
  NAND U11161 ( .A(n7054), .B(n7055), .Z(n7050) );
  AND U11162 ( .A(n7056), .B(n7057), .Z(n6948) );
  NAND U11163 ( .A(n7058), .B(n7059), .Z(n7057) );
  NAND U11164 ( .A(n7060), .B(n7061), .Z(n7056) );
  AND U11165 ( .A(n7062), .B(n7063), .Z(n6950) );
  XOR U11166 ( .A(n7030), .B(n7029), .Z(N29573) );
  XNOR U11167 ( .A(n7048), .B(n7047), .Z(n7029) );
  XNOR U11168 ( .A(n7062), .B(n7063), .Z(n7047) );
  XOR U11169 ( .A(n7059), .B(n7058), .Z(n7063) );
  XOR U11170 ( .A(y[3291]), .B(x[3291]), .Z(n7058) );
  XOR U11171 ( .A(n7061), .B(n7060), .Z(n7059) );
  XOR U11172 ( .A(y[3293]), .B(x[3293]), .Z(n7060) );
  XOR U11173 ( .A(y[3292]), .B(x[3292]), .Z(n7061) );
  XOR U11174 ( .A(n7053), .B(n7052), .Z(n7062) );
  XOR U11175 ( .A(n7055), .B(n7054), .Z(n7052) );
  XOR U11176 ( .A(y[3290]), .B(x[3290]), .Z(n7054) );
  XOR U11177 ( .A(y[3289]), .B(x[3289]), .Z(n7055) );
  XOR U11178 ( .A(y[3288]), .B(x[3288]), .Z(n7053) );
  XNOR U11179 ( .A(n7046), .B(n7045), .Z(n7048) );
  XNOR U11180 ( .A(n7042), .B(n7041), .Z(n7045) );
  XOR U11181 ( .A(n7044), .B(n7043), .Z(n7041) );
  XOR U11182 ( .A(y[3287]), .B(x[3287]), .Z(n7043) );
  XOR U11183 ( .A(y[3286]), .B(x[3286]), .Z(n7044) );
  XOR U11184 ( .A(y[3285]), .B(x[3285]), .Z(n7042) );
  XOR U11185 ( .A(n7036), .B(n7035), .Z(n7046) );
  XOR U11186 ( .A(n7038), .B(n7037), .Z(n7035) );
  XOR U11187 ( .A(y[3284]), .B(x[3284]), .Z(n7037) );
  XOR U11188 ( .A(y[3283]), .B(x[3283]), .Z(n7038) );
  XOR U11189 ( .A(y[3282]), .B(x[3282]), .Z(n7036) );
  XNOR U11190 ( .A(n7013), .B(n7012), .Z(n7030) );
  XNOR U11191 ( .A(n7027), .B(n7028), .Z(n7012) );
  XOR U11192 ( .A(n7024), .B(n7023), .Z(n7028) );
  XOR U11193 ( .A(y[3279]), .B(x[3279]), .Z(n7023) );
  XOR U11194 ( .A(n7026), .B(n7025), .Z(n7024) );
  XOR U11195 ( .A(y[3281]), .B(x[3281]), .Z(n7025) );
  XOR U11196 ( .A(y[3280]), .B(x[3280]), .Z(n7026) );
  XOR U11197 ( .A(n7018), .B(n7017), .Z(n7027) );
  XOR U11198 ( .A(n7020), .B(n7019), .Z(n7017) );
  XOR U11199 ( .A(y[3278]), .B(x[3278]), .Z(n7019) );
  XOR U11200 ( .A(y[3277]), .B(x[3277]), .Z(n7020) );
  XOR U11201 ( .A(y[3276]), .B(x[3276]), .Z(n7018) );
  XNOR U11202 ( .A(n7011), .B(n7010), .Z(n7013) );
  XNOR U11203 ( .A(n7007), .B(n7006), .Z(n7010) );
  XOR U11204 ( .A(n7009), .B(n7008), .Z(n7006) );
  XOR U11205 ( .A(y[3275]), .B(x[3275]), .Z(n7008) );
  XOR U11206 ( .A(y[3274]), .B(x[3274]), .Z(n7009) );
  XOR U11207 ( .A(y[3273]), .B(x[3273]), .Z(n7007) );
  XOR U11208 ( .A(n7001), .B(n7000), .Z(n7011) );
  XOR U11209 ( .A(n7003), .B(n7002), .Z(n7000) );
  XOR U11210 ( .A(y[3272]), .B(x[3272]), .Z(n7002) );
  XOR U11211 ( .A(y[3271]), .B(x[3271]), .Z(n7003) );
  XOR U11212 ( .A(y[3270]), .B(x[3270]), .Z(n7001) );
  NAND U11213 ( .A(n7064), .B(n7065), .Z(N29565) );
  NAND U11214 ( .A(n7066), .B(n7067), .Z(n7065) );
  NANDN U11215 ( .A(n7068), .B(n7069), .Z(n7067) );
  NANDN U11216 ( .A(n7069), .B(n7068), .Z(n7064) );
  XOR U11217 ( .A(n7068), .B(n7070), .Z(N29564) );
  XNOR U11218 ( .A(n7066), .B(n7069), .Z(n7070) );
  NAND U11219 ( .A(n7071), .B(n7072), .Z(n7069) );
  NAND U11220 ( .A(n7073), .B(n7074), .Z(n7072) );
  NANDN U11221 ( .A(n7075), .B(n7076), .Z(n7074) );
  NANDN U11222 ( .A(n7076), .B(n7075), .Z(n7071) );
  AND U11223 ( .A(n7077), .B(n7078), .Z(n7066) );
  NAND U11224 ( .A(n7079), .B(n7080), .Z(n7078) );
  OR U11225 ( .A(n7081), .B(n7082), .Z(n7080) );
  NAND U11226 ( .A(n7082), .B(n7081), .Z(n7077) );
  IV U11227 ( .A(n7083), .Z(n7082) );
  AND U11228 ( .A(n7084), .B(n7085), .Z(n7068) );
  NAND U11229 ( .A(n7086), .B(n7087), .Z(n7085) );
  NANDN U11230 ( .A(n7088), .B(n7089), .Z(n7087) );
  NANDN U11231 ( .A(n7089), .B(n7088), .Z(n7084) );
  XOR U11232 ( .A(n7081), .B(n7090), .Z(N29563) );
  XOR U11233 ( .A(n7079), .B(n7083), .Z(n7090) );
  XNOR U11234 ( .A(n7076), .B(n7091), .Z(n7083) );
  XNOR U11235 ( .A(n7073), .B(n7075), .Z(n7091) );
  AND U11236 ( .A(n7092), .B(n7093), .Z(n7075) );
  NANDN U11237 ( .A(n7094), .B(n7095), .Z(n7093) );
  NANDN U11238 ( .A(n7096), .B(n7097), .Z(n7095) );
  IV U11239 ( .A(n7098), .Z(n7097) );
  NAND U11240 ( .A(n7098), .B(n7096), .Z(n7092) );
  AND U11241 ( .A(n7099), .B(n7100), .Z(n7073) );
  NAND U11242 ( .A(n7101), .B(n7102), .Z(n7100) );
  OR U11243 ( .A(n7103), .B(n7104), .Z(n7102) );
  NAND U11244 ( .A(n7104), .B(n7103), .Z(n7099) );
  IV U11245 ( .A(n7105), .Z(n7104) );
  NAND U11246 ( .A(n7106), .B(n7107), .Z(n7076) );
  NANDN U11247 ( .A(n7108), .B(n7109), .Z(n7107) );
  NAND U11248 ( .A(n7110), .B(n7111), .Z(n7109) );
  OR U11249 ( .A(n7111), .B(n7110), .Z(n7106) );
  IV U11250 ( .A(n7112), .Z(n7110) );
  AND U11251 ( .A(n7113), .B(n7114), .Z(n7079) );
  NAND U11252 ( .A(n7115), .B(n7116), .Z(n7114) );
  NANDN U11253 ( .A(n7117), .B(n7118), .Z(n7116) );
  NANDN U11254 ( .A(n7118), .B(n7117), .Z(n7113) );
  XOR U11255 ( .A(n7089), .B(n7119), .Z(n7081) );
  XNOR U11256 ( .A(n7086), .B(n7088), .Z(n7119) );
  AND U11257 ( .A(n7120), .B(n7121), .Z(n7088) );
  NANDN U11258 ( .A(n7122), .B(n7123), .Z(n7121) );
  NANDN U11259 ( .A(n7124), .B(n7125), .Z(n7123) );
  IV U11260 ( .A(n7126), .Z(n7125) );
  NAND U11261 ( .A(n7126), .B(n7124), .Z(n7120) );
  AND U11262 ( .A(n7127), .B(n7128), .Z(n7086) );
  NAND U11263 ( .A(n7129), .B(n7130), .Z(n7128) );
  OR U11264 ( .A(n7131), .B(n7132), .Z(n7130) );
  NAND U11265 ( .A(n7132), .B(n7131), .Z(n7127) );
  IV U11266 ( .A(n7133), .Z(n7132) );
  NAND U11267 ( .A(n7134), .B(n7135), .Z(n7089) );
  NANDN U11268 ( .A(n7136), .B(n7137), .Z(n7135) );
  NAND U11269 ( .A(n7138), .B(n7139), .Z(n7137) );
  OR U11270 ( .A(n7139), .B(n7138), .Z(n7134) );
  IV U11271 ( .A(n7140), .Z(n7138) );
  XOR U11272 ( .A(n7115), .B(n7141), .Z(N29562) );
  XNOR U11273 ( .A(n7118), .B(n7117), .Z(n7141) );
  XNOR U11274 ( .A(n7129), .B(n7142), .Z(n7117) );
  XOR U11275 ( .A(n7133), .B(n7131), .Z(n7142) );
  XOR U11276 ( .A(n7139), .B(n7143), .Z(n7131) );
  XOR U11277 ( .A(n7136), .B(n7140), .Z(n7143) );
  NAND U11278 ( .A(n7144), .B(n7145), .Z(n7140) );
  NAND U11279 ( .A(n7146), .B(n7147), .Z(n7145) );
  NAND U11280 ( .A(n7148), .B(n7149), .Z(n7144) );
  AND U11281 ( .A(n7150), .B(n7151), .Z(n7136) );
  NAND U11282 ( .A(n7152), .B(n7153), .Z(n7151) );
  NAND U11283 ( .A(n7154), .B(n7155), .Z(n7150) );
  NANDN U11284 ( .A(n7156), .B(n7157), .Z(n7139) );
  NANDN U11285 ( .A(n7158), .B(n7159), .Z(n7133) );
  XNOR U11286 ( .A(n7124), .B(n7160), .Z(n7129) );
  XOR U11287 ( .A(n7122), .B(n7126), .Z(n7160) );
  NAND U11288 ( .A(n7161), .B(n7162), .Z(n7126) );
  NAND U11289 ( .A(n7163), .B(n7164), .Z(n7162) );
  NAND U11290 ( .A(n7165), .B(n7166), .Z(n7161) );
  AND U11291 ( .A(n7167), .B(n7168), .Z(n7122) );
  NAND U11292 ( .A(n7169), .B(n7170), .Z(n7168) );
  NAND U11293 ( .A(n7171), .B(n7172), .Z(n7167) );
  AND U11294 ( .A(n7173), .B(n7174), .Z(n7124) );
  NAND U11295 ( .A(n7175), .B(n7176), .Z(n7118) );
  XNOR U11296 ( .A(n7101), .B(n7177), .Z(n7115) );
  XOR U11297 ( .A(n7105), .B(n7103), .Z(n7177) );
  XOR U11298 ( .A(n7111), .B(n7178), .Z(n7103) );
  XOR U11299 ( .A(n7108), .B(n7112), .Z(n7178) );
  NAND U11300 ( .A(n7179), .B(n7180), .Z(n7112) );
  NAND U11301 ( .A(n7181), .B(n7182), .Z(n7180) );
  NAND U11302 ( .A(n7183), .B(n7184), .Z(n7179) );
  AND U11303 ( .A(n7185), .B(n7186), .Z(n7108) );
  NAND U11304 ( .A(n7187), .B(n7188), .Z(n7186) );
  NAND U11305 ( .A(n7189), .B(n7190), .Z(n7185) );
  NANDN U11306 ( .A(n7191), .B(n7192), .Z(n7111) );
  NANDN U11307 ( .A(n7193), .B(n7194), .Z(n7105) );
  XNOR U11308 ( .A(n7096), .B(n7195), .Z(n7101) );
  XOR U11309 ( .A(n7094), .B(n7098), .Z(n7195) );
  NAND U11310 ( .A(n7196), .B(n7197), .Z(n7098) );
  NAND U11311 ( .A(n7198), .B(n7199), .Z(n7197) );
  NAND U11312 ( .A(n7200), .B(n7201), .Z(n7196) );
  AND U11313 ( .A(n7202), .B(n7203), .Z(n7094) );
  NAND U11314 ( .A(n7204), .B(n7205), .Z(n7203) );
  NAND U11315 ( .A(n7206), .B(n7207), .Z(n7202) );
  AND U11316 ( .A(n7208), .B(n7209), .Z(n7096) );
  XOR U11317 ( .A(n7176), .B(n7175), .Z(N29561) );
  XNOR U11318 ( .A(n7194), .B(n7193), .Z(n7175) );
  XNOR U11319 ( .A(n7208), .B(n7209), .Z(n7193) );
  XOR U11320 ( .A(n7205), .B(n7204), .Z(n7209) );
  XOR U11321 ( .A(y[3267]), .B(x[3267]), .Z(n7204) );
  XOR U11322 ( .A(n7207), .B(n7206), .Z(n7205) );
  XOR U11323 ( .A(y[3269]), .B(x[3269]), .Z(n7206) );
  XOR U11324 ( .A(y[3268]), .B(x[3268]), .Z(n7207) );
  XOR U11325 ( .A(n7199), .B(n7198), .Z(n7208) );
  XOR U11326 ( .A(n7201), .B(n7200), .Z(n7198) );
  XOR U11327 ( .A(y[3266]), .B(x[3266]), .Z(n7200) );
  XOR U11328 ( .A(y[3265]), .B(x[3265]), .Z(n7201) );
  XOR U11329 ( .A(y[3264]), .B(x[3264]), .Z(n7199) );
  XNOR U11330 ( .A(n7192), .B(n7191), .Z(n7194) );
  XNOR U11331 ( .A(n7188), .B(n7187), .Z(n7191) );
  XOR U11332 ( .A(n7190), .B(n7189), .Z(n7187) );
  XOR U11333 ( .A(y[3263]), .B(x[3263]), .Z(n7189) );
  XOR U11334 ( .A(y[3262]), .B(x[3262]), .Z(n7190) );
  XOR U11335 ( .A(y[3261]), .B(x[3261]), .Z(n7188) );
  XOR U11336 ( .A(n7182), .B(n7181), .Z(n7192) );
  XOR U11337 ( .A(n7184), .B(n7183), .Z(n7181) );
  XOR U11338 ( .A(y[3260]), .B(x[3260]), .Z(n7183) );
  XOR U11339 ( .A(y[3259]), .B(x[3259]), .Z(n7184) );
  XOR U11340 ( .A(y[3258]), .B(x[3258]), .Z(n7182) );
  XNOR U11341 ( .A(n7159), .B(n7158), .Z(n7176) );
  XNOR U11342 ( .A(n7173), .B(n7174), .Z(n7158) );
  XOR U11343 ( .A(n7170), .B(n7169), .Z(n7174) );
  XOR U11344 ( .A(y[3255]), .B(x[3255]), .Z(n7169) );
  XOR U11345 ( .A(n7172), .B(n7171), .Z(n7170) );
  XOR U11346 ( .A(y[3257]), .B(x[3257]), .Z(n7171) );
  XOR U11347 ( .A(y[3256]), .B(x[3256]), .Z(n7172) );
  XOR U11348 ( .A(n7164), .B(n7163), .Z(n7173) );
  XOR U11349 ( .A(n7166), .B(n7165), .Z(n7163) );
  XOR U11350 ( .A(y[3254]), .B(x[3254]), .Z(n7165) );
  XOR U11351 ( .A(y[3253]), .B(x[3253]), .Z(n7166) );
  XOR U11352 ( .A(y[3252]), .B(x[3252]), .Z(n7164) );
  XNOR U11353 ( .A(n7157), .B(n7156), .Z(n7159) );
  XNOR U11354 ( .A(n7153), .B(n7152), .Z(n7156) );
  XOR U11355 ( .A(n7155), .B(n7154), .Z(n7152) );
  XOR U11356 ( .A(y[3251]), .B(x[3251]), .Z(n7154) );
  XOR U11357 ( .A(y[3250]), .B(x[3250]), .Z(n7155) );
  XOR U11358 ( .A(y[3249]), .B(x[3249]), .Z(n7153) );
  XOR U11359 ( .A(n7147), .B(n7146), .Z(n7157) );
  XOR U11360 ( .A(n7149), .B(n7148), .Z(n7146) );
  XOR U11361 ( .A(y[3248]), .B(x[3248]), .Z(n7148) );
  XOR U11362 ( .A(y[3247]), .B(x[3247]), .Z(n7149) );
  XOR U11363 ( .A(y[3246]), .B(x[3246]), .Z(n7147) );
  NAND U11364 ( .A(n7210), .B(n7211), .Z(N29553) );
  NAND U11365 ( .A(n7212), .B(n7213), .Z(n7211) );
  NANDN U11366 ( .A(n7214), .B(n7215), .Z(n7213) );
  NANDN U11367 ( .A(n7215), .B(n7214), .Z(n7210) );
  XOR U11368 ( .A(n7214), .B(n7216), .Z(N29552) );
  XNOR U11369 ( .A(n7212), .B(n7215), .Z(n7216) );
  NAND U11370 ( .A(n7217), .B(n7218), .Z(n7215) );
  NAND U11371 ( .A(n7219), .B(n7220), .Z(n7218) );
  NANDN U11372 ( .A(n7221), .B(n7222), .Z(n7220) );
  NANDN U11373 ( .A(n7222), .B(n7221), .Z(n7217) );
  AND U11374 ( .A(n7223), .B(n7224), .Z(n7212) );
  NAND U11375 ( .A(n7225), .B(n7226), .Z(n7224) );
  OR U11376 ( .A(n7227), .B(n7228), .Z(n7226) );
  NAND U11377 ( .A(n7228), .B(n7227), .Z(n7223) );
  IV U11378 ( .A(n7229), .Z(n7228) );
  AND U11379 ( .A(n7230), .B(n7231), .Z(n7214) );
  NAND U11380 ( .A(n7232), .B(n7233), .Z(n7231) );
  NANDN U11381 ( .A(n7234), .B(n7235), .Z(n7233) );
  NANDN U11382 ( .A(n7235), .B(n7234), .Z(n7230) );
  XOR U11383 ( .A(n7227), .B(n7236), .Z(N29551) );
  XOR U11384 ( .A(n7225), .B(n7229), .Z(n7236) );
  XNOR U11385 ( .A(n7222), .B(n7237), .Z(n7229) );
  XNOR U11386 ( .A(n7219), .B(n7221), .Z(n7237) );
  AND U11387 ( .A(n7238), .B(n7239), .Z(n7221) );
  NANDN U11388 ( .A(n7240), .B(n7241), .Z(n7239) );
  NANDN U11389 ( .A(n7242), .B(n7243), .Z(n7241) );
  IV U11390 ( .A(n7244), .Z(n7243) );
  NAND U11391 ( .A(n7244), .B(n7242), .Z(n7238) );
  AND U11392 ( .A(n7245), .B(n7246), .Z(n7219) );
  NAND U11393 ( .A(n7247), .B(n7248), .Z(n7246) );
  OR U11394 ( .A(n7249), .B(n7250), .Z(n7248) );
  NAND U11395 ( .A(n7250), .B(n7249), .Z(n7245) );
  IV U11396 ( .A(n7251), .Z(n7250) );
  NAND U11397 ( .A(n7252), .B(n7253), .Z(n7222) );
  NANDN U11398 ( .A(n7254), .B(n7255), .Z(n7253) );
  NAND U11399 ( .A(n7256), .B(n7257), .Z(n7255) );
  OR U11400 ( .A(n7257), .B(n7256), .Z(n7252) );
  IV U11401 ( .A(n7258), .Z(n7256) );
  AND U11402 ( .A(n7259), .B(n7260), .Z(n7225) );
  NAND U11403 ( .A(n7261), .B(n7262), .Z(n7260) );
  NANDN U11404 ( .A(n7263), .B(n7264), .Z(n7262) );
  NANDN U11405 ( .A(n7264), .B(n7263), .Z(n7259) );
  XOR U11406 ( .A(n7235), .B(n7265), .Z(n7227) );
  XNOR U11407 ( .A(n7232), .B(n7234), .Z(n7265) );
  AND U11408 ( .A(n7266), .B(n7267), .Z(n7234) );
  NANDN U11409 ( .A(n7268), .B(n7269), .Z(n7267) );
  NANDN U11410 ( .A(n7270), .B(n7271), .Z(n7269) );
  IV U11411 ( .A(n7272), .Z(n7271) );
  NAND U11412 ( .A(n7272), .B(n7270), .Z(n7266) );
  AND U11413 ( .A(n7273), .B(n7274), .Z(n7232) );
  NAND U11414 ( .A(n7275), .B(n7276), .Z(n7274) );
  OR U11415 ( .A(n7277), .B(n7278), .Z(n7276) );
  NAND U11416 ( .A(n7278), .B(n7277), .Z(n7273) );
  IV U11417 ( .A(n7279), .Z(n7278) );
  NAND U11418 ( .A(n7280), .B(n7281), .Z(n7235) );
  NANDN U11419 ( .A(n7282), .B(n7283), .Z(n7281) );
  NAND U11420 ( .A(n7284), .B(n7285), .Z(n7283) );
  OR U11421 ( .A(n7285), .B(n7284), .Z(n7280) );
  IV U11422 ( .A(n7286), .Z(n7284) );
  XOR U11423 ( .A(n7261), .B(n7287), .Z(N29550) );
  XNOR U11424 ( .A(n7264), .B(n7263), .Z(n7287) );
  XNOR U11425 ( .A(n7275), .B(n7288), .Z(n7263) );
  XOR U11426 ( .A(n7279), .B(n7277), .Z(n7288) );
  XOR U11427 ( .A(n7285), .B(n7289), .Z(n7277) );
  XOR U11428 ( .A(n7282), .B(n7286), .Z(n7289) );
  NAND U11429 ( .A(n7290), .B(n7291), .Z(n7286) );
  NAND U11430 ( .A(n7292), .B(n7293), .Z(n7291) );
  NAND U11431 ( .A(n7294), .B(n7295), .Z(n7290) );
  AND U11432 ( .A(n7296), .B(n7297), .Z(n7282) );
  NAND U11433 ( .A(n7298), .B(n7299), .Z(n7297) );
  NAND U11434 ( .A(n7300), .B(n7301), .Z(n7296) );
  NANDN U11435 ( .A(n7302), .B(n7303), .Z(n7285) );
  NANDN U11436 ( .A(n7304), .B(n7305), .Z(n7279) );
  XNOR U11437 ( .A(n7270), .B(n7306), .Z(n7275) );
  XOR U11438 ( .A(n7268), .B(n7272), .Z(n7306) );
  NAND U11439 ( .A(n7307), .B(n7308), .Z(n7272) );
  NAND U11440 ( .A(n7309), .B(n7310), .Z(n7308) );
  NAND U11441 ( .A(n7311), .B(n7312), .Z(n7307) );
  AND U11442 ( .A(n7313), .B(n7314), .Z(n7268) );
  NAND U11443 ( .A(n7315), .B(n7316), .Z(n7314) );
  NAND U11444 ( .A(n7317), .B(n7318), .Z(n7313) );
  AND U11445 ( .A(n7319), .B(n7320), .Z(n7270) );
  NAND U11446 ( .A(n7321), .B(n7322), .Z(n7264) );
  XNOR U11447 ( .A(n7247), .B(n7323), .Z(n7261) );
  XOR U11448 ( .A(n7251), .B(n7249), .Z(n7323) );
  XOR U11449 ( .A(n7257), .B(n7324), .Z(n7249) );
  XOR U11450 ( .A(n7254), .B(n7258), .Z(n7324) );
  NAND U11451 ( .A(n7325), .B(n7326), .Z(n7258) );
  NAND U11452 ( .A(n7327), .B(n7328), .Z(n7326) );
  NAND U11453 ( .A(n7329), .B(n7330), .Z(n7325) );
  AND U11454 ( .A(n7331), .B(n7332), .Z(n7254) );
  NAND U11455 ( .A(n7333), .B(n7334), .Z(n7332) );
  NAND U11456 ( .A(n7335), .B(n7336), .Z(n7331) );
  NANDN U11457 ( .A(n7337), .B(n7338), .Z(n7257) );
  NANDN U11458 ( .A(n7339), .B(n7340), .Z(n7251) );
  XNOR U11459 ( .A(n7242), .B(n7341), .Z(n7247) );
  XOR U11460 ( .A(n7240), .B(n7244), .Z(n7341) );
  NAND U11461 ( .A(n7342), .B(n7343), .Z(n7244) );
  NAND U11462 ( .A(n7344), .B(n7345), .Z(n7343) );
  NAND U11463 ( .A(n7346), .B(n7347), .Z(n7342) );
  AND U11464 ( .A(n7348), .B(n7349), .Z(n7240) );
  NAND U11465 ( .A(n7350), .B(n7351), .Z(n7349) );
  NAND U11466 ( .A(n7352), .B(n7353), .Z(n7348) );
  AND U11467 ( .A(n7354), .B(n7355), .Z(n7242) );
  XOR U11468 ( .A(n7322), .B(n7321), .Z(N29549) );
  XNOR U11469 ( .A(n7340), .B(n7339), .Z(n7321) );
  XNOR U11470 ( .A(n7354), .B(n7355), .Z(n7339) );
  XOR U11471 ( .A(n7351), .B(n7350), .Z(n7355) );
  XOR U11472 ( .A(y[3243]), .B(x[3243]), .Z(n7350) );
  XOR U11473 ( .A(n7353), .B(n7352), .Z(n7351) );
  XOR U11474 ( .A(y[3245]), .B(x[3245]), .Z(n7352) );
  XOR U11475 ( .A(y[3244]), .B(x[3244]), .Z(n7353) );
  XOR U11476 ( .A(n7345), .B(n7344), .Z(n7354) );
  XOR U11477 ( .A(n7347), .B(n7346), .Z(n7344) );
  XOR U11478 ( .A(y[3242]), .B(x[3242]), .Z(n7346) );
  XOR U11479 ( .A(y[3241]), .B(x[3241]), .Z(n7347) );
  XOR U11480 ( .A(y[3240]), .B(x[3240]), .Z(n7345) );
  XNOR U11481 ( .A(n7338), .B(n7337), .Z(n7340) );
  XNOR U11482 ( .A(n7334), .B(n7333), .Z(n7337) );
  XOR U11483 ( .A(n7336), .B(n7335), .Z(n7333) );
  XOR U11484 ( .A(y[3239]), .B(x[3239]), .Z(n7335) );
  XOR U11485 ( .A(y[3238]), .B(x[3238]), .Z(n7336) );
  XOR U11486 ( .A(y[3237]), .B(x[3237]), .Z(n7334) );
  XOR U11487 ( .A(n7328), .B(n7327), .Z(n7338) );
  XOR U11488 ( .A(n7330), .B(n7329), .Z(n7327) );
  XOR U11489 ( .A(y[3236]), .B(x[3236]), .Z(n7329) );
  XOR U11490 ( .A(y[3235]), .B(x[3235]), .Z(n7330) );
  XOR U11491 ( .A(y[3234]), .B(x[3234]), .Z(n7328) );
  XNOR U11492 ( .A(n7305), .B(n7304), .Z(n7322) );
  XNOR U11493 ( .A(n7319), .B(n7320), .Z(n7304) );
  XOR U11494 ( .A(n7316), .B(n7315), .Z(n7320) );
  XOR U11495 ( .A(y[3231]), .B(x[3231]), .Z(n7315) );
  XOR U11496 ( .A(n7318), .B(n7317), .Z(n7316) );
  XOR U11497 ( .A(y[3233]), .B(x[3233]), .Z(n7317) );
  XOR U11498 ( .A(y[3232]), .B(x[3232]), .Z(n7318) );
  XOR U11499 ( .A(n7310), .B(n7309), .Z(n7319) );
  XOR U11500 ( .A(n7312), .B(n7311), .Z(n7309) );
  XOR U11501 ( .A(y[3230]), .B(x[3230]), .Z(n7311) );
  XOR U11502 ( .A(y[3229]), .B(x[3229]), .Z(n7312) );
  XOR U11503 ( .A(y[3228]), .B(x[3228]), .Z(n7310) );
  XNOR U11504 ( .A(n7303), .B(n7302), .Z(n7305) );
  XNOR U11505 ( .A(n7299), .B(n7298), .Z(n7302) );
  XOR U11506 ( .A(n7301), .B(n7300), .Z(n7298) );
  XOR U11507 ( .A(y[3227]), .B(x[3227]), .Z(n7300) );
  XOR U11508 ( .A(y[3226]), .B(x[3226]), .Z(n7301) );
  XOR U11509 ( .A(y[3225]), .B(x[3225]), .Z(n7299) );
  XOR U11510 ( .A(n7293), .B(n7292), .Z(n7303) );
  XOR U11511 ( .A(n7295), .B(n7294), .Z(n7292) );
  XOR U11512 ( .A(y[3224]), .B(x[3224]), .Z(n7294) );
  XOR U11513 ( .A(y[3223]), .B(x[3223]), .Z(n7295) );
  XOR U11514 ( .A(y[3222]), .B(x[3222]), .Z(n7293) );
  NAND U11515 ( .A(n7356), .B(n7357), .Z(N29541) );
  NAND U11516 ( .A(n7358), .B(n7359), .Z(n7357) );
  NANDN U11517 ( .A(n7360), .B(n7361), .Z(n7359) );
  NANDN U11518 ( .A(n7361), .B(n7360), .Z(n7356) );
  XOR U11519 ( .A(n7360), .B(n7362), .Z(N29540) );
  XNOR U11520 ( .A(n7358), .B(n7361), .Z(n7362) );
  NAND U11521 ( .A(n7363), .B(n7364), .Z(n7361) );
  NAND U11522 ( .A(n7365), .B(n7366), .Z(n7364) );
  NANDN U11523 ( .A(n7367), .B(n7368), .Z(n7366) );
  NANDN U11524 ( .A(n7368), .B(n7367), .Z(n7363) );
  AND U11525 ( .A(n7369), .B(n7370), .Z(n7358) );
  NAND U11526 ( .A(n7371), .B(n7372), .Z(n7370) );
  OR U11527 ( .A(n7373), .B(n7374), .Z(n7372) );
  NAND U11528 ( .A(n7374), .B(n7373), .Z(n7369) );
  IV U11529 ( .A(n7375), .Z(n7374) );
  AND U11530 ( .A(n7376), .B(n7377), .Z(n7360) );
  NAND U11531 ( .A(n7378), .B(n7379), .Z(n7377) );
  NANDN U11532 ( .A(n7380), .B(n7381), .Z(n7379) );
  NANDN U11533 ( .A(n7381), .B(n7380), .Z(n7376) );
  XOR U11534 ( .A(n7373), .B(n7382), .Z(N29539) );
  XOR U11535 ( .A(n7371), .B(n7375), .Z(n7382) );
  XNOR U11536 ( .A(n7368), .B(n7383), .Z(n7375) );
  XNOR U11537 ( .A(n7365), .B(n7367), .Z(n7383) );
  AND U11538 ( .A(n7384), .B(n7385), .Z(n7367) );
  NANDN U11539 ( .A(n7386), .B(n7387), .Z(n7385) );
  NANDN U11540 ( .A(n7388), .B(n7389), .Z(n7387) );
  IV U11541 ( .A(n7390), .Z(n7389) );
  NAND U11542 ( .A(n7390), .B(n7388), .Z(n7384) );
  AND U11543 ( .A(n7391), .B(n7392), .Z(n7365) );
  NAND U11544 ( .A(n7393), .B(n7394), .Z(n7392) );
  OR U11545 ( .A(n7395), .B(n7396), .Z(n7394) );
  NAND U11546 ( .A(n7396), .B(n7395), .Z(n7391) );
  IV U11547 ( .A(n7397), .Z(n7396) );
  NAND U11548 ( .A(n7398), .B(n7399), .Z(n7368) );
  NANDN U11549 ( .A(n7400), .B(n7401), .Z(n7399) );
  NAND U11550 ( .A(n7402), .B(n7403), .Z(n7401) );
  OR U11551 ( .A(n7403), .B(n7402), .Z(n7398) );
  IV U11552 ( .A(n7404), .Z(n7402) );
  AND U11553 ( .A(n7405), .B(n7406), .Z(n7371) );
  NAND U11554 ( .A(n7407), .B(n7408), .Z(n7406) );
  NANDN U11555 ( .A(n7409), .B(n7410), .Z(n7408) );
  NANDN U11556 ( .A(n7410), .B(n7409), .Z(n7405) );
  XOR U11557 ( .A(n7381), .B(n7411), .Z(n7373) );
  XNOR U11558 ( .A(n7378), .B(n7380), .Z(n7411) );
  AND U11559 ( .A(n7412), .B(n7413), .Z(n7380) );
  NANDN U11560 ( .A(n7414), .B(n7415), .Z(n7413) );
  NANDN U11561 ( .A(n7416), .B(n7417), .Z(n7415) );
  IV U11562 ( .A(n7418), .Z(n7417) );
  NAND U11563 ( .A(n7418), .B(n7416), .Z(n7412) );
  AND U11564 ( .A(n7419), .B(n7420), .Z(n7378) );
  NAND U11565 ( .A(n7421), .B(n7422), .Z(n7420) );
  OR U11566 ( .A(n7423), .B(n7424), .Z(n7422) );
  NAND U11567 ( .A(n7424), .B(n7423), .Z(n7419) );
  IV U11568 ( .A(n7425), .Z(n7424) );
  NAND U11569 ( .A(n7426), .B(n7427), .Z(n7381) );
  NANDN U11570 ( .A(n7428), .B(n7429), .Z(n7427) );
  NAND U11571 ( .A(n7430), .B(n7431), .Z(n7429) );
  OR U11572 ( .A(n7431), .B(n7430), .Z(n7426) );
  IV U11573 ( .A(n7432), .Z(n7430) );
  XOR U11574 ( .A(n7407), .B(n7433), .Z(N29538) );
  XNOR U11575 ( .A(n7410), .B(n7409), .Z(n7433) );
  XNOR U11576 ( .A(n7421), .B(n7434), .Z(n7409) );
  XOR U11577 ( .A(n7425), .B(n7423), .Z(n7434) );
  XOR U11578 ( .A(n7431), .B(n7435), .Z(n7423) );
  XOR U11579 ( .A(n7428), .B(n7432), .Z(n7435) );
  NAND U11580 ( .A(n7436), .B(n7437), .Z(n7432) );
  NAND U11581 ( .A(n7438), .B(n7439), .Z(n7437) );
  NAND U11582 ( .A(n7440), .B(n7441), .Z(n7436) );
  AND U11583 ( .A(n7442), .B(n7443), .Z(n7428) );
  NAND U11584 ( .A(n7444), .B(n7445), .Z(n7443) );
  NAND U11585 ( .A(n7446), .B(n7447), .Z(n7442) );
  NANDN U11586 ( .A(n7448), .B(n7449), .Z(n7431) );
  NANDN U11587 ( .A(n7450), .B(n7451), .Z(n7425) );
  XNOR U11588 ( .A(n7416), .B(n7452), .Z(n7421) );
  XOR U11589 ( .A(n7414), .B(n7418), .Z(n7452) );
  NAND U11590 ( .A(n7453), .B(n7454), .Z(n7418) );
  NAND U11591 ( .A(n7455), .B(n7456), .Z(n7454) );
  NAND U11592 ( .A(n7457), .B(n7458), .Z(n7453) );
  AND U11593 ( .A(n7459), .B(n7460), .Z(n7414) );
  NAND U11594 ( .A(n7461), .B(n7462), .Z(n7460) );
  NAND U11595 ( .A(n7463), .B(n7464), .Z(n7459) );
  AND U11596 ( .A(n7465), .B(n7466), .Z(n7416) );
  NAND U11597 ( .A(n7467), .B(n7468), .Z(n7410) );
  XNOR U11598 ( .A(n7393), .B(n7469), .Z(n7407) );
  XOR U11599 ( .A(n7397), .B(n7395), .Z(n7469) );
  XOR U11600 ( .A(n7403), .B(n7470), .Z(n7395) );
  XOR U11601 ( .A(n7400), .B(n7404), .Z(n7470) );
  NAND U11602 ( .A(n7471), .B(n7472), .Z(n7404) );
  NAND U11603 ( .A(n7473), .B(n7474), .Z(n7472) );
  NAND U11604 ( .A(n7475), .B(n7476), .Z(n7471) );
  AND U11605 ( .A(n7477), .B(n7478), .Z(n7400) );
  NAND U11606 ( .A(n7479), .B(n7480), .Z(n7478) );
  NAND U11607 ( .A(n7481), .B(n7482), .Z(n7477) );
  NANDN U11608 ( .A(n7483), .B(n7484), .Z(n7403) );
  NANDN U11609 ( .A(n7485), .B(n7486), .Z(n7397) );
  XNOR U11610 ( .A(n7388), .B(n7487), .Z(n7393) );
  XOR U11611 ( .A(n7386), .B(n7390), .Z(n7487) );
  NAND U11612 ( .A(n7488), .B(n7489), .Z(n7390) );
  NAND U11613 ( .A(n7490), .B(n7491), .Z(n7489) );
  NAND U11614 ( .A(n7492), .B(n7493), .Z(n7488) );
  AND U11615 ( .A(n7494), .B(n7495), .Z(n7386) );
  NAND U11616 ( .A(n7496), .B(n7497), .Z(n7495) );
  NAND U11617 ( .A(n7498), .B(n7499), .Z(n7494) );
  AND U11618 ( .A(n7500), .B(n7501), .Z(n7388) );
  XOR U11619 ( .A(n7468), .B(n7467), .Z(N29537) );
  XNOR U11620 ( .A(n7486), .B(n7485), .Z(n7467) );
  XNOR U11621 ( .A(n7500), .B(n7501), .Z(n7485) );
  XOR U11622 ( .A(n7497), .B(n7496), .Z(n7501) );
  XOR U11623 ( .A(y[3219]), .B(x[3219]), .Z(n7496) );
  XOR U11624 ( .A(n7499), .B(n7498), .Z(n7497) );
  XOR U11625 ( .A(y[3221]), .B(x[3221]), .Z(n7498) );
  XOR U11626 ( .A(y[3220]), .B(x[3220]), .Z(n7499) );
  XOR U11627 ( .A(n7491), .B(n7490), .Z(n7500) );
  XOR U11628 ( .A(n7493), .B(n7492), .Z(n7490) );
  XOR U11629 ( .A(y[3218]), .B(x[3218]), .Z(n7492) );
  XOR U11630 ( .A(y[3217]), .B(x[3217]), .Z(n7493) );
  XOR U11631 ( .A(y[3216]), .B(x[3216]), .Z(n7491) );
  XNOR U11632 ( .A(n7484), .B(n7483), .Z(n7486) );
  XNOR U11633 ( .A(n7480), .B(n7479), .Z(n7483) );
  XOR U11634 ( .A(n7482), .B(n7481), .Z(n7479) );
  XOR U11635 ( .A(y[3215]), .B(x[3215]), .Z(n7481) );
  XOR U11636 ( .A(y[3214]), .B(x[3214]), .Z(n7482) );
  XOR U11637 ( .A(y[3213]), .B(x[3213]), .Z(n7480) );
  XOR U11638 ( .A(n7474), .B(n7473), .Z(n7484) );
  XOR U11639 ( .A(n7476), .B(n7475), .Z(n7473) );
  XOR U11640 ( .A(y[3212]), .B(x[3212]), .Z(n7475) );
  XOR U11641 ( .A(y[3211]), .B(x[3211]), .Z(n7476) );
  XOR U11642 ( .A(y[3210]), .B(x[3210]), .Z(n7474) );
  XNOR U11643 ( .A(n7451), .B(n7450), .Z(n7468) );
  XNOR U11644 ( .A(n7465), .B(n7466), .Z(n7450) );
  XOR U11645 ( .A(n7462), .B(n7461), .Z(n7466) );
  XOR U11646 ( .A(y[3207]), .B(x[3207]), .Z(n7461) );
  XOR U11647 ( .A(n7464), .B(n7463), .Z(n7462) );
  XOR U11648 ( .A(y[3209]), .B(x[3209]), .Z(n7463) );
  XOR U11649 ( .A(y[3208]), .B(x[3208]), .Z(n7464) );
  XOR U11650 ( .A(n7456), .B(n7455), .Z(n7465) );
  XOR U11651 ( .A(n7458), .B(n7457), .Z(n7455) );
  XOR U11652 ( .A(y[3206]), .B(x[3206]), .Z(n7457) );
  XOR U11653 ( .A(y[3205]), .B(x[3205]), .Z(n7458) );
  XOR U11654 ( .A(y[3204]), .B(x[3204]), .Z(n7456) );
  XNOR U11655 ( .A(n7449), .B(n7448), .Z(n7451) );
  XNOR U11656 ( .A(n7445), .B(n7444), .Z(n7448) );
  XOR U11657 ( .A(n7447), .B(n7446), .Z(n7444) );
  XOR U11658 ( .A(y[3203]), .B(x[3203]), .Z(n7446) );
  XOR U11659 ( .A(y[3202]), .B(x[3202]), .Z(n7447) );
  XOR U11660 ( .A(y[3201]), .B(x[3201]), .Z(n7445) );
  XOR U11661 ( .A(n7439), .B(n7438), .Z(n7449) );
  XOR U11662 ( .A(n7441), .B(n7440), .Z(n7438) );
  XOR U11663 ( .A(y[3200]), .B(x[3200]), .Z(n7440) );
  XOR U11664 ( .A(y[3199]), .B(x[3199]), .Z(n7441) );
  XOR U11665 ( .A(y[3198]), .B(x[3198]), .Z(n7439) );
  NAND U11666 ( .A(n7502), .B(n7503), .Z(N29529) );
  NAND U11667 ( .A(n7504), .B(n7505), .Z(n7503) );
  NANDN U11668 ( .A(n7506), .B(n7507), .Z(n7505) );
  NANDN U11669 ( .A(n7507), .B(n7506), .Z(n7502) );
  XOR U11670 ( .A(n7506), .B(n7508), .Z(N29528) );
  XNOR U11671 ( .A(n7504), .B(n7507), .Z(n7508) );
  NAND U11672 ( .A(n7509), .B(n7510), .Z(n7507) );
  NAND U11673 ( .A(n7511), .B(n7512), .Z(n7510) );
  NANDN U11674 ( .A(n7513), .B(n7514), .Z(n7512) );
  NANDN U11675 ( .A(n7514), .B(n7513), .Z(n7509) );
  AND U11676 ( .A(n7515), .B(n7516), .Z(n7504) );
  NAND U11677 ( .A(n7517), .B(n7518), .Z(n7516) );
  OR U11678 ( .A(n7519), .B(n7520), .Z(n7518) );
  NAND U11679 ( .A(n7520), .B(n7519), .Z(n7515) );
  IV U11680 ( .A(n7521), .Z(n7520) );
  AND U11681 ( .A(n7522), .B(n7523), .Z(n7506) );
  NAND U11682 ( .A(n7524), .B(n7525), .Z(n7523) );
  NANDN U11683 ( .A(n7526), .B(n7527), .Z(n7525) );
  NANDN U11684 ( .A(n7527), .B(n7526), .Z(n7522) );
  XOR U11685 ( .A(n7519), .B(n7528), .Z(N29527) );
  XOR U11686 ( .A(n7517), .B(n7521), .Z(n7528) );
  XNOR U11687 ( .A(n7514), .B(n7529), .Z(n7521) );
  XNOR U11688 ( .A(n7511), .B(n7513), .Z(n7529) );
  AND U11689 ( .A(n7530), .B(n7531), .Z(n7513) );
  NANDN U11690 ( .A(n7532), .B(n7533), .Z(n7531) );
  NANDN U11691 ( .A(n7534), .B(n7535), .Z(n7533) );
  IV U11692 ( .A(n7536), .Z(n7535) );
  NAND U11693 ( .A(n7536), .B(n7534), .Z(n7530) );
  AND U11694 ( .A(n7537), .B(n7538), .Z(n7511) );
  NAND U11695 ( .A(n7539), .B(n7540), .Z(n7538) );
  OR U11696 ( .A(n7541), .B(n7542), .Z(n7540) );
  NAND U11697 ( .A(n7542), .B(n7541), .Z(n7537) );
  IV U11698 ( .A(n7543), .Z(n7542) );
  NAND U11699 ( .A(n7544), .B(n7545), .Z(n7514) );
  NANDN U11700 ( .A(n7546), .B(n7547), .Z(n7545) );
  NAND U11701 ( .A(n7548), .B(n7549), .Z(n7547) );
  OR U11702 ( .A(n7549), .B(n7548), .Z(n7544) );
  IV U11703 ( .A(n7550), .Z(n7548) );
  AND U11704 ( .A(n7551), .B(n7552), .Z(n7517) );
  NAND U11705 ( .A(n7553), .B(n7554), .Z(n7552) );
  NANDN U11706 ( .A(n7555), .B(n7556), .Z(n7554) );
  NANDN U11707 ( .A(n7556), .B(n7555), .Z(n7551) );
  XOR U11708 ( .A(n7527), .B(n7557), .Z(n7519) );
  XNOR U11709 ( .A(n7524), .B(n7526), .Z(n7557) );
  AND U11710 ( .A(n7558), .B(n7559), .Z(n7526) );
  NANDN U11711 ( .A(n7560), .B(n7561), .Z(n7559) );
  NANDN U11712 ( .A(n7562), .B(n7563), .Z(n7561) );
  IV U11713 ( .A(n7564), .Z(n7563) );
  NAND U11714 ( .A(n7564), .B(n7562), .Z(n7558) );
  AND U11715 ( .A(n7565), .B(n7566), .Z(n7524) );
  NAND U11716 ( .A(n7567), .B(n7568), .Z(n7566) );
  OR U11717 ( .A(n7569), .B(n7570), .Z(n7568) );
  NAND U11718 ( .A(n7570), .B(n7569), .Z(n7565) );
  IV U11719 ( .A(n7571), .Z(n7570) );
  NAND U11720 ( .A(n7572), .B(n7573), .Z(n7527) );
  NANDN U11721 ( .A(n7574), .B(n7575), .Z(n7573) );
  NAND U11722 ( .A(n7576), .B(n7577), .Z(n7575) );
  OR U11723 ( .A(n7577), .B(n7576), .Z(n7572) );
  IV U11724 ( .A(n7578), .Z(n7576) );
  XOR U11725 ( .A(n7553), .B(n7579), .Z(N29526) );
  XNOR U11726 ( .A(n7556), .B(n7555), .Z(n7579) );
  XNOR U11727 ( .A(n7567), .B(n7580), .Z(n7555) );
  XOR U11728 ( .A(n7571), .B(n7569), .Z(n7580) );
  XOR U11729 ( .A(n7577), .B(n7581), .Z(n7569) );
  XOR U11730 ( .A(n7574), .B(n7578), .Z(n7581) );
  NAND U11731 ( .A(n7582), .B(n7583), .Z(n7578) );
  NAND U11732 ( .A(n7584), .B(n7585), .Z(n7583) );
  NAND U11733 ( .A(n7586), .B(n7587), .Z(n7582) );
  AND U11734 ( .A(n7588), .B(n7589), .Z(n7574) );
  NAND U11735 ( .A(n7590), .B(n7591), .Z(n7589) );
  NAND U11736 ( .A(n7592), .B(n7593), .Z(n7588) );
  NANDN U11737 ( .A(n7594), .B(n7595), .Z(n7577) );
  NANDN U11738 ( .A(n7596), .B(n7597), .Z(n7571) );
  XNOR U11739 ( .A(n7562), .B(n7598), .Z(n7567) );
  XOR U11740 ( .A(n7560), .B(n7564), .Z(n7598) );
  NAND U11741 ( .A(n7599), .B(n7600), .Z(n7564) );
  NAND U11742 ( .A(n7601), .B(n7602), .Z(n7600) );
  NAND U11743 ( .A(n7603), .B(n7604), .Z(n7599) );
  AND U11744 ( .A(n7605), .B(n7606), .Z(n7560) );
  NAND U11745 ( .A(n7607), .B(n7608), .Z(n7606) );
  NAND U11746 ( .A(n7609), .B(n7610), .Z(n7605) );
  AND U11747 ( .A(n7611), .B(n7612), .Z(n7562) );
  NAND U11748 ( .A(n7613), .B(n7614), .Z(n7556) );
  XNOR U11749 ( .A(n7539), .B(n7615), .Z(n7553) );
  XOR U11750 ( .A(n7543), .B(n7541), .Z(n7615) );
  XOR U11751 ( .A(n7549), .B(n7616), .Z(n7541) );
  XOR U11752 ( .A(n7546), .B(n7550), .Z(n7616) );
  NAND U11753 ( .A(n7617), .B(n7618), .Z(n7550) );
  NAND U11754 ( .A(n7619), .B(n7620), .Z(n7618) );
  NAND U11755 ( .A(n7621), .B(n7622), .Z(n7617) );
  AND U11756 ( .A(n7623), .B(n7624), .Z(n7546) );
  NAND U11757 ( .A(n7625), .B(n7626), .Z(n7624) );
  NAND U11758 ( .A(n7627), .B(n7628), .Z(n7623) );
  NANDN U11759 ( .A(n7629), .B(n7630), .Z(n7549) );
  NANDN U11760 ( .A(n7631), .B(n7632), .Z(n7543) );
  XNOR U11761 ( .A(n7534), .B(n7633), .Z(n7539) );
  XOR U11762 ( .A(n7532), .B(n7536), .Z(n7633) );
  NAND U11763 ( .A(n7634), .B(n7635), .Z(n7536) );
  NAND U11764 ( .A(n7636), .B(n7637), .Z(n7635) );
  NAND U11765 ( .A(n7638), .B(n7639), .Z(n7634) );
  AND U11766 ( .A(n7640), .B(n7641), .Z(n7532) );
  NAND U11767 ( .A(n7642), .B(n7643), .Z(n7641) );
  NAND U11768 ( .A(n7644), .B(n7645), .Z(n7640) );
  AND U11769 ( .A(n7646), .B(n7647), .Z(n7534) );
  XOR U11770 ( .A(n7614), .B(n7613), .Z(N29525) );
  XNOR U11771 ( .A(n7632), .B(n7631), .Z(n7613) );
  XNOR U11772 ( .A(n7646), .B(n7647), .Z(n7631) );
  XOR U11773 ( .A(n7643), .B(n7642), .Z(n7647) );
  XOR U11774 ( .A(y[3195]), .B(x[3195]), .Z(n7642) );
  XOR U11775 ( .A(n7645), .B(n7644), .Z(n7643) );
  XOR U11776 ( .A(y[3197]), .B(x[3197]), .Z(n7644) );
  XOR U11777 ( .A(y[3196]), .B(x[3196]), .Z(n7645) );
  XOR U11778 ( .A(n7637), .B(n7636), .Z(n7646) );
  XOR U11779 ( .A(n7639), .B(n7638), .Z(n7636) );
  XOR U11780 ( .A(y[3194]), .B(x[3194]), .Z(n7638) );
  XOR U11781 ( .A(y[3193]), .B(x[3193]), .Z(n7639) );
  XOR U11782 ( .A(y[3192]), .B(x[3192]), .Z(n7637) );
  XNOR U11783 ( .A(n7630), .B(n7629), .Z(n7632) );
  XNOR U11784 ( .A(n7626), .B(n7625), .Z(n7629) );
  XOR U11785 ( .A(n7628), .B(n7627), .Z(n7625) );
  XOR U11786 ( .A(y[3191]), .B(x[3191]), .Z(n7627) );
  XOR U11787 ( .A(y[3190]), .B(x[3190]), .Z(n7628) );
  XOR U11788 ( .A(y[3189]), .B(x[3189]), .Z(n7626) );
  XOR U11789 ( .A(n7620), .B(n7619), .Z(n7630) );
  XOR U11790 ( .A(n7622), .B(n7621), .Z(n7619) );
  XOR U11791 ( .A(y[3188]), .B(x[3188]), .Z(n7621) );
  XOR U11792 ( .A(y[3187]), .B(x[3187]), .Z(n7622) );
  XOR U11793 ( .A(y[3186]), .B(x[3186]), .Z(n7620) );
  XNOR U11794 ( .A(n7597), .B(n7596), .Z(n7614) );
  XNOR U11795 ( .A(n7611), .B(n7612), .Z(n7596) );
  XOR U11796 ( .A(n7608), .B(n7607), .Z(n7612) );
  XOR U11797 ( .A(y[3183]), .B(x[3183]), .Z(n7607) );
  XOR U11798 ( .A(n7610), .B(n7609), .Z(n7608) );
  XOR U11799 ( .A(y[3185]), .B(x[3185]), .Z(n7609) );
  XOR U11800 ( .A(y[3184]), .B(x[3184]), .Z(n7610) );
  XOR U11801 ( .A(n7602), .B(n7601), .Z(n7611) );
  XOR U11802 ( .A(n7604), .B(n7603), .Z(n7601) );
  XOR U11803 ( .A(y[3182]), .B(x[3182]), .Z(n7603) );
  XOR U11804 ( .A(y[3181]), .B(x[3181]), .Z(n7604) );
  XOR U11805 ( .A(y[3180]), .B(x[3180]), .Z(n7602) );
  XNOR U11806 ( .A(n7595), .B(n7594), .Z(n7597) );
  XNOR U11807 ( .A(n7591), .B(n7590), .Z(n7594) );
  XOR U11808 ( .A(n7593), .B(n7592), .Z(n7590) );
  XOR U11809 ( .A(y[3179]), .B(x[3179]), .Z(n7592) );
  XOR U11810 ( .A(y[3178]), .B(x[3178]), .Z(n7593) );
  XOR U11811 ( .A(y[3177]), .B(x[3177]), .Z(n7591) );
  XOR U11812 ( .A(n7585), .B(n7584), .Z(n7595) );
  XOR U11813 ( .A(n7587), .B(n7586), .Z(n7584) );
  XOR U11814 ( .A(y[3176]), .B(x[3176]), .Z(n7586) );
  XOR U11815 ( .A(y[3175]), .B(x[3175]), .Z(n7587) );
  XOR U11816 ( .A(y[3174]), .B(x[3174]), .Z(n7585) );
  NAND U11817 ( .A(n7648), .B(n7649), .Z(N29517) );
  NAND U11818 ( .A(n7650), .B(n7651), .Z(n7649) );
  NANDN U11819 ( .A(n7652), .B(n7653), .Z(n7651) );
  NANDN U11820 ( .A(n7653), .B(n7652), .Z(n7648) );
  XOR U11821 ( .A(n7652), .B(n7654), .Z(N29516) );
  XNOR U11822 ( .A(n7650), .B(n7653), .Z(n7654) );
  NAND U11823 ( .A(n7655), .B(n7656), .Z(n7653) );
  NAND U11824 ( .A(n7657), .B(n7658), .Z(n7656) );
  NANDN U11825 ( .A(n7659), .B(n7660), .Z(n7658) );
  NANDN U11826 ( .A(n7660), .B(n7659), .Z(n7655) );
  AND U11827 ( .A(n7661), .B(n7662), .Z(n7650) );
  NAND U11828 ( .A(n7663), .B(n7664), .Z(n7662) );
  OR U11829 ( .A(n7665), .B(n7666), .Z(n7664) );
  NAND U11830 ( .A(n7666), .B(n7665), .Z(n7661) );
  IV U11831 ( .A(n7667), .Z(n7666) );
  AND U11832 ( .A(n7668), .B(n7669), .Z(n7652) );
  NAND U11833 ( .A(n7670), .B(n7671), .Z(n7669) );
  NANDN U11834 ( .A(n7672), .B(n7673), .Z(n7671) );
  NANDN U11835 ( .A(n7673), .B(n7672), .Z(n7668) );
  XOR U11836 ( .A(n7665), .B(n7674), .Z(N29515) );
  XOR U11837 ( .A(n7663), .B(n7667), .Z(n7674) );
  XNOR U11838 ( .A(n7660), .B(n7675), .Z(n7667) );
  XNOR U11839 ( .A(n7657), .B(n7659), .Z(n7675) );
  AND U11840 ( .A(n7676), .B(n7677), .Z(n7659) );
  NANDN U11841 ( .A(n7678), .B(n7679), .Z(n7677) );
  NANDN U11842 ( .A(n7680), .B(n7681), .Z(n7679) );
  IV U11843 ( .A(n7682), .Z(n7681) );
  NAND U11844 ( .A(n7682), .B(n7680), .Z(n7676) );
  AND U11845 ( .A(n7683), .B(n7684), .Z(n7657) );
  NAND U11846 ( .A(n7685), .B(n7686), .Z(n7684) );
  OR U11847 ( .A(n7687), .B(n7688), .Z(n7686) );
  NAND U11848 ( .A(n7688), .B(n7687), .Z(n7683) );
  IV U11849 ( .A(n7689), .Z(n7688) );
  NAND U11850 ( .A(n7690), .B(n7691), .Z(n7660) );
  NANDN U11851 ( .A(n7692), .B(n7693), .Z(n7691) );
  NAND U11852 ( .A(n7694), .B(n7695), .Z(n7693) );
  OR U11853 ( .A(n7695), .B(n7694), .Z(n7690) );
  IV U11854 ( .A(n7696), .Z(n7694) );
  AND U11855 ( .A(n7697), .B(n7698), .Z(n7663) );
  NAND U11856 ( .A(n7699), .B(n7700), .Z(n7698) );
  NANDN U11857 ( .A(n7701), .B(n7702), .Z(n7700) );
  NANDN U11858 ( .A(n7702), .B(n7701), .Z(n7697) );
  XOR U11859 ( .A(n7673), .B(n7703), .Z(n7665) );
  XNOR U11860 ( .A(n7670), .B(n7672), .Z(n7703) );
  AND U11861 ( .A(n7704), .B(n7705), .Z(n7672) );
  NANDN U11862 ( .A(n7706), .B(n7707), .Z(n7705) );
  NANDN U11863 ( .A(n7708), .B(n7709), .Z(n7707) );
  IV U11864 ( .A(n7710), .Z(n7709) );
  NAND U11865 ( .A(n7710), .B(n7708), .Z(n7704) );
  AND U11866 ( .A(n7711), .B(n7712), .Z(n7670) );
  NAND U11867 ( .A(n7713), .B(n7714), .Z(n7712) );
  OR U11868 ( .A(n7715), .B(n7716), .Z(n7714) );
  NAND U11869 ( .A(n7716), .B(n7715), .Z(n7711) );
  IV U11870 ( .A(n7717), .Z(n7716) );
  NAND U11871 ( .A(n7718), .B(n7719), .Z(n7673) );
  NANDN U11872 ( .A(n7720), .B(n7721), .Z(n7719) );
  NAND U11873 ( .A(n7722), .B(n7723), .Z(n7721) );
  OR U11874 ( .A(n7723), .B(n7722), .Z(n7718) );
  IV U11875 ( .A(n7724), .Z(n7722) );
  XOR U11876 ( .A(n7699), .B(n7725), .Z(N29514) );
  XNOR U11877 ( .A(n7702), .B(n7701), .Z(n7725) );
  XNOR U11878 ( .A(n7713), .B(n7726), .Z(n7701) );
  XOR U11879 ( .A(n7717), .B(n7715), .Z(n7726) );
  XOR U11880 ( .A(n7723), .B(n7727), .Z(n7715) );
  XOR U11881 ( .A(n7720), .B(n7724), .Z(n7727) );
  NAND U11882 ( .A(n7728), .B(n7729), .Z(n7724) );
  NAND U11883 ( .A(n7730), .B(n7731), .Z(n7729) );
  NAND U11884 ( .A(n7732), .B(n7733), .Z(n7728) );
  AND U11885 ( .A(n7734), .B(n7735), .Z(n7720) );
  NAND U11886 ( .A(n7736), .B(n7737), .Z(n7735) );
  NAND U11887 ( .A(n7738), .B(n7739), .Z(n7734) );
  NANDN U11888 ( .A(n7740), .B(n7741), .Z(n7723) );
  NANDN U11889 ( .A(n7742), .B(n7743), .Z(n7717) );
  XNOR U11890 ( .A(n7708), .B(n7744), .Z(n7713) );
  XOR U11891 ( .A(n7706), .B(n7710), .Z(n7744) );
  NAND U11892 ( .A(n7745), .B(n7746), .Z(n7710) );
  NAND U11893 ( .A(n7747), .B(n7748), .Z(n7746) );
  NAND U11894 ( .A(n7749), .B(n7750), .Z(n7745) );
  AND U11895 ( .A(n7751), .B(n7752), .Z(n7706) );
  NAND U11896 ( .A(n7753), .B(n7754), .Z(n7752) );
  NAND U11897 ( .A(n7755), .B(n7756), .Z(n7751) );
  AND U11898 ( .A(n7757), .B(n7758), .Z(n7708) );
  NAND U11899 ( .A(n7759), .B(n7760), .Z(n7702) );
  XNOR U11900 ( .A(n7685), .B(n7761), .Z(n7699) );
  XOR U11901 ( .A(n7689), .B(n7687), .Z(n7761) );
  XOR U11902 ( .A(n7695), .B(n7762), .Z(n7687) );
  XOR U11903 ( .A(n7692), .B(n7696), .Z(n7762) );
  NAND U11904 ( .A(n7763), .B(n7764), .Z(n7696) );
  NAND U11905 ( .A(n7765), .B(n7766), .Z(n7764) );
  NAND U11906 ( .A(n7767), .B(n7768), .Z(n7763) );
  AND U11907 ( .A(n7769), .B(n7770), .Z(n7692) );
  NAND U11908 ( .A(n7771), .B(n7772), .Z(n7770) );
  NAND U11909 ( .A(n7773), .B(n7774), .Z(n7769) );
  NANDN U11910 ( .A(n7775), .B(n7776), .Z(n7695) );
  NANDN U11911 ( .A(n7777), .B(n7778), .Z(n7689) );
  XNOR U11912 ( .A(n7680), .B(n7779), .Z(n7685) );
  XOR U11913 ( .A(n7678), .B(n7682), .Z(n7779) );
  NAND U11914 ( .A(n7780), .B(n7781), .Z(n7682) );
  NAND U11915 ( .A(n7782), .B(n7783), .Z(n7781) );
  NAND U11916 ( .A(n7784), .B(n7785), .Z(n7780) );
  AND U11917 ( .A(n7786), .B(n7787), .Z(n7678) );
  NAND U11918 ( .A(n7788), .B(n7789), .Z(n7787) );
  NAND U11919 ( .A(n7790), .B(n7791), .Z(n7786) );
  AND U11920 ( .A(n7792), .B(n7793), .Z(n7680) );
  XOR U11921 ( .A(n7760), .B(n7759), .Z(N29513) );
  XNOR U11922 ( .A(n7778), .B(n7777), .Z(n7759) );
  XNOR U11923 ( .A(n7792), .B(n7793), .Z(n7777) );
  XOR U11924 ( .A(n7789), .B(n7788), .Z(n7793) );
  XOR U11925 ( .A(y[3171]), .B(x[3171]), .Z(n7788) );
  XOR U11926 ( .A(n7791), .B(n7790), .Z(n7789) );
  XOR U11927 ( .A(y[3173]), .B(x[3173]), .Z(n7790) );
  XOR U11928 ( .A(y[3172]), .B(x[3172]), .Z(n7791) );
  XOR U11929 ( .A(n7783), .B(n7782), .Z(n7792) );
  XOR U11930 ( .A(n7785), .B(n7784), .Z(n7782) );
  XOR U11931 ( .A(y[3170]), .B(x[3170]), .Z(n7784) );
  XOR U11932 ( .A(y[3169]), .B(x[3169]), .Z(n7785) );
  XOR U11933 ( .A(y[3168]), .B(x[3168]), .Z(n7783) );
  XNOR U11934 ( .A(n7776), .B(n7775), .Z(n7778) );
  XNOR U11935 ( .A(n7772), .B(n7771), .Z(n7775) );
  XOR U11936 ( .A(n7774), .B(n7773), .Z(n7771) );
  XOR U11937 ( .A(y[3167]), .B(x[3167]), .Z(n7773) );
  XOR U11938 ( .A(y[3166]), .B(x[3166]), .Z(n7774) );
  XOR U11939 ( .A(y[3165]), .B(x[3165]), .Z(n7772) );
  XOR U11940 ( .A(n7766), .B(n7765), .Z(n7776) );
  XOR U11941 ( .A(n7768), .B(n7767), .Z(n7765) );
  XOR U11942 ( .A(y[3164]), .B(x[3164]), .Z(n7767) );
  XOR U11943 ( .A(y[3163]), .B(x[3163]), .Z(n7768) );
  XOR U11944 ( .A(y[3162]), .B(x[3162]), .Z(n7766) );
  XNOR U11945 ( .A(n7743), .B(n7742), .Z(n7760) );
  XNOR U11946 ( .A(n7757), .B(n7758), .Z(n7742) );
  XOR U11947 ( .A(n7754), .B(n7753), .Z(n7758) );
  XOR U11948 ( .A(y[3159]), .B(x[3159]), .Z(n7753) );
  XOR U11949 ( .A(n7756), .B(n7755), .Z(n7754) );
  XOR U11950 ( .A(y[3161]), .B(x[3161]), .Z(n7755) );
  XOR U11951 ( .A(y[3160]), .B(x[3160]), .Z(n7756) );
  XOR U11952 ( .A(n7748), .B(n7747), .Z(n7757) );
  XOR U11953 ( .A(n7750), .B(n7749), .Z(n7747) );
  XOR U11954 ( .A(y[3158]), .B(x[3158]), .Z(n7749) );
  XOR U11955 ( .A(y[3157]), .B(x[3157]), .Z(n7750) );
  XOR U11956 ( .A(y[3156]), .B(x[3156]), .Z(n7748) );
  XNOR U11957 ( .A(n7741), .B(n7740), .Z(n7743) );
  XNOR U11958 ( .A(n7737), .B(n7736), .Z(n7740) );
  XOR U11959 ( .A(n7739), .B(n7738), .Z(n7736) );
  XOR U11960 ( .A(y[3155]), .B(x[3155]), .Z(n7738) );
  XOR U11961 ( .A(y[3154]), .B(x[3154]), .Z(n7739) );
  XOR U11962 ( .A(y[3153]), .B(x[3153]), .Z(n7737) );
  XOR U11963 ( .A(n7731), .B(n7730), .Z(n7741) );
  XOR U11964 ( .A(n7733), .B(n7732), .Z(n7730) );
  XOR U11965 ( .A(y[3152]), .B(x[3152]), .Z(n7732) );
  XOR U11966 ( .A(y[3151]), .B(x[3151]), .Z(n7733) );
  XOR U11967 ( .A(y[3150]), .B(x[3150]), .Z(n7731) );
  NAND U11968 ( .A(n7794), .B(n7795), .Z(N29505) );
  NAND U11969 ( .A(n7796), .B(n7797), .Z(n7795) );
  NANDN U11970 ( .A(n7798), .B(n7799), .Z(n7797) );
  NANDN U11971 ( .A(n7799), .B(n7798), .Z(n7794) );
  XOR U11972 ( .A(n7798), .B(n7800), .Z(N29504) );
  XNOR U11973 ( .A(n7796), .B(n7799), .Z(n7800) );
  NAND U11974 ( .A(n7801), .B(n7802), .Z(n7799) );
  NAND U11975 ( .A(n7803), .B(n7804), .Z(n7802) );
  NANDN U11976 ( .A(n7805), .B(n7806), .Z(n7804) );
  NANDN U11977 ( .A(n7806), .B(n7805), .Z(n7801) );
  AND U11978 ( .A(n7807), .B(n7808), .Z(n7796) );
  NAND U11979 ( .A(n7809), .B(n7810), .Z(n7808) );
  OR U11980 ( .A(n7811), .B(n7812), .Z(n7810) );
  NAND U11981 ( .A(n7812), .B(n7811), .Z(n7807) );
  IV U11982 ( .A(n7813), .Z(n7812) );
  AND U11983 ( .A(n7814), .B(n7815), .Z(n7798) );
  NAND U11984 ( .A(n7816), .B(n7817), .Z(n7815) );
  NANDN U11985 ( .A(n7818), .B(n7819), .Z(n7817) );
  NANDN U11986 ( .A(n7819), .B(n7818), .Z(n7814) );
  XOR U11987 ( .A(n7811), .B(n7820), .Z(N29503) );
  XOR U11988 ( .A(n7809), .B(n7813), .Z(n7820) );
  XNOR U11989 ( .A(n7806), .B(n7821), .Z(n7813) );
  XNOR U11990 ( .A(n7803), .B(n7805), .Z(n7821) );
  AND U11991 ( .A(n7822), .B(n7823), .Z(n7805) );
  NANDN U11992 ( .A(n7824), .B(n7825), .Z(n7823) );
  NANDN U11993 ( .A(n7826), .B(n7827), .Z(n7825) );
  IV U11994 ( .A(n7828), .Z(n7827) );
  NAND U11995 ( .A(n7828), .B(n7826), .Z(n7822) );
  AND U11996 ( .A(n7829), .B(n7830), .Z(n7803) );
  NAND U11997 ( .A(n7831), .B(n7832), .Z(n7830) );
  OR U11998 ( .A(n7833), .B(n7834), .Z(n7832) );
  NAND U11999 ( .A(n7834), .B(n7833), .Z(n7829) );
  IV U12000 ( .A(n7835), .Z(n7834) );
  NAND U12001 ( .A(n7836), .B(n7837), .Z(n7806) );
  NANDN U12002 ( .A(n7838), .B(n7839), .Z(n7837) );
  NAND U12003 ( .A(n7840), .B(n7841), .Z(n7839) );
  OR U12004 ( .A(n7841), .B(n7840), .Z(n7836) );
  IV U12005 ( .A(n7842), .Z(n7840) );
  AND U12006 ( .A(n7843), .B(n7844), .Z(n7809) );
  NAND U12007 ( .A(n7845), .B(n7846), .Z(n7844) );
  NANDN U12008 ( .A(n7847), .B(n7848), .Z(n7846) );
  NANDN U12009 ( .A(n7848), .B(n7847), .Z(n7843) );
  XOR U12010 ( .A(n7819), .B(n7849), .Z(n7811) );
  XNOR U12011 ( .A(n7816), .B(n7818), .Z(n7849) );
  AND U12012 ( .A(n7850), .B(n7851), .Z(n7818) );
  NANDN U12013 ( .A(n7852), .B(n7853), .Z(n7851) );
  NANDN U12014 ( .A(n7854), .B(n7855), .Z(n7853) );
  IV U12015 ( .A(n7856), .Z(n7855) );
  NAND U12016 ( .A(n7856), .B(n7854), .Z(n7850) );
  AND U12017 ( .A(n7857), .B(n7858), .Z(n7816) );
  NAND U12018 ( .A(n7859), .B(n7860), .Z(n7858) );
  OR U12019 ( .A(n7861), .B(n7862), .Z(n7860) );
  NAND U12020 ( .A(n7862), .B(n7861), .Z(n7857) );
  IV U12021 ( .A(n7863), .Z(n7862) );
  NAND U12022 ( .A(n7864), .B(n7865), .Z(n7819) );
  NANDN U12023 ( .A(n7866), .B(n7867), .Z(n7865) );
  NAND U12024 ( .A(n7868), .B(n7869), .Z(n7867) );
  OR U12025 ( .A(n7869), .B(n7868), .Z(n7864) );
  IV U12026 ( .A(n7870), .Z(n7868) );
  XOR U12027 ( .A(n7845), .B(n7871), .Z(N29502) );
  XNOR U12028 ( .A(n7848), .B(n7847), .Z(n7871) );
  XNOR U12029 ( .A(n7859), .B(n7872), .Z(n7847) );
  XOR U12030 ( .A(n7863), .B(n7861), .Z(n7872) );
  XOR U12031 ( .A(n7869), .B(n7873), .Z(n7861) );
  XOR U12032 ( .A(n7866), .B(n7870), .Z(n7873) );
  NAND U12033 ( .A(n7874), .B(n7875), .Z(n7870) );
  NAND U12034 ( .A(n7876), .B(n7877), .Z(n7875) );
  NAND U12035 ( .A(n7878), .B(n7879), .Z(n7874) );
  AND U12036 ( .A(n7880), .B(n7881), .Z(n7866) );
  NAND U12037 ( .A(n7882), .B(n7883), .Z(n7881) );
  NAND U12038 ( .A(n7884), .B(n7885), .Z(n7880) );
  NANDN U12039 ( .A(n7886), .B(n7887), .Z(n7869) );
  NANDN U12040 ( .A(n7888), .B(n7889), .Z(n7863) );
  XNOR U12041 ( .A(n7854), .B(n7890), .Z(n7859) );
  XOR U12042 ( .A(n7852), .B(n7856), .Z(n7890) );
  NAND U12043 ( .A(n7891), .B(n7892), .Z(n7856) );
  NAND U12044 ( .A(n7893), .B(n7894), .Z(n7892) );
  NAND U12045 ( .A(n7895), .B(n7896), .Z(n7891) );
  AND U12046 ( .A(n7897), .B(n7898), .Z(n7852) );
  NAND U12047 ( .A(n7899), .B(n7900), .Z(n7898) );
  NAND U12048 ( .A(n7901), .B(n7902), .Z(n7897) );
  AND U12049 ( .A(n7903), .B(n7904), .Z(n7854) );
  NAND U12050 ( .A(n7905), .B(n7906), .Z(n7848) );
  XNOR U12051 ( .A(n7831), .B(n7907), .Z(n7845) );
  XOR U12052 ( .A(n7835), .B(n7833), .Z(n7907) );
  XOR U12053 ( .A(n7841), .B(n7908), .Z(n7833) );
  XOR U12054 ( .A(n7838), .B(n7842), .Z(n7908) );
  NAND U12055 ( .A(n7909), .B(n7910), .Z(n7842) );
  NAND U12056 ( .A(n7911), .B(n7912), .Z(n7910) );
  NAND U12057 ( .A(n7913), .B(n7914), .Z(n7909) );
  AND U12058 ( .A(n7915), .B(n7916), .Z(n7838) );
  NAND U12059 ( .A(n7917), .B(n7918), .Z(n7916) );
  NAND U12060 ( .A(n7919), .B(n7920), .Z(n7915) );
  NANDN U12061 ( .A(n7921), .B(n7922), .Z(n7841) );
  NANDN U12062 ( .A(n7923), .B(n7924), .Z(n7835) );
  XNOR U12063 ( .A(n7826), .B(n7925), .Z(n7831) );
  XOR U12064 ( .A(n7824), .B(n7828), .Z(n7925) );
  NAND U12065 ( .A(n7926), .B(n7927), .Z(n7828) );
  NAND U12066 ( .A(n7928), .B(n7929), .Z(n7927) );
  NAND U12067 ( .A(n7930), .B(n7931), .Z(n7926) );
  AND U12068 ( .A(n7932), .B(n7933), .Z(n7824) );
  NAND U12069 ( .A(n7934), .B(n7935), .Z(n7933) );
  NAND U12070 ( .A(n7936), .B(n7937), .Z(n7932) );
  AND U12071 ( .A(n7938), .B(n7939), .Z(n7826) );
  XOR U12072 ( .A(n7906), .B(n7905), .Z(N29501) );
  XNOR U12073 ( .A(n7924), .B(n7923), .Z(n7905) );
  XNOR U12074 ( .A(n7938), .B(n7939), .Z(n7923) );
  XOR U12075 ( .A(n7935), .B(n7934), .Z(n7939) );
  XOR U12076 ( .A(y[3147]), .B(x[3147]), .Z(n7934) );
  XOR U12077 ( .A(n7937), .B(n7936), .Z(n7935) );
  XOR U12078 ( .A(y[3149]), .B(x[3149]), .Z(n7936) );
  XOR U12079 ( .A(y[3148]), .B(x[3148]), .Z(n7937) );
  XOR U12080 ( .A(n7929), .B(n7928), .Z(n7938) );
  XOR U12081 ( .A(n7931), .B(n7930), .Z(n7928) );
  XOR U12082 ( .A(y[3146]), .B(x[3146]), .Z(n7930) );
  XOR U12083 ( .A(y[3145]), .B(x[3145]), .Z(n7931) );
  XOR U12084 ( .A(y[3144]), .B(x[3144]), .Z(n7929) );
  XNOR U12085 ( .A(n7922), .B(n7921), .Z(n7924) );
  XNOR U12086 ( .A(n7918), .B(n7917), .Z(n7921) );
  XOR U12087 ( .A(n7920), .B(n7919), .Z(n7917) );
  XOR U12088 ( .A(y[3143]), .B(x[3143]), .Z(n7919) );
  XOR U12089 ( .A(y[3142]), .B(x[3142]), .Z(n7920) );
  XOR U12090 ( .A(y[3141]), .B(x[3141]), .Z(n7918) );
  XOR U12091 ( .A(n7912), .B(n7911), .Z(n7922) );
  XOR U12092 ( .A(n7914), .B(n7913), .Z(n7911) );
  XOR U12093 ( .A(y[3140]), .B(x[3140]), .Z(n7913) );
  XOR U12094 ( .A(y[3139]), .B(x[3139]), .Z(n7914) );
  XOR U12095 ( .A(y[3138]), .B(x[3138]), .Z(n7912) );
  XNOR U12096 ( .A(n7889), .B(n7888), .Z(n7906) );
  XNOR U12097 ( .A(n7903), .B(n7904), .Z(n7888) );
  XOR U12098 ( .A(n7900), .B(n7899), .Z(n7904) );
  XOR U12099 ( .A(y[3135]), .B(x[3135]), .Z(n7899) );
  XOR U12100 ( .A(n7902), .B(n7901), .Z(n7900) );
  XOR U12101 ( .A(y[3137]), .B(x[3137]), .Z(n7901) );
  XOR U12102 ( .A(y[3136]), .B(x[3136]), .Z(n7902) );
  XOR U12103 ( .A(n7894), .B(n7893), .Z(n7903) );
  XOR U12104 ( .A(n7896), .B(n7895), .Z(n7893) );
  XOR U12105 ( .A(y[3134]), .B(x[3134]), .Z(n7895) );
  XOR U12106 ( .A(y[3133]), .B(x[3133]), .Z(n7896) );
  XOR U12107 ( .A(y[3132]), .B(x[3132]), .Z(n7894) );
  XNOR U12108 ( .A(n7887), .B(n7886), .Z(n7889) );
  XNOR U12109 ( .A(n7883), .B(n7882), .Z(n7886) );
  XOR U12110 ( .A(n7885), .B(n7884), .Z(n7882) );
  XOR U12111 ( .A(y[3131]), .B(x[3131]), .Z(n7884) );
  XOR U12112 ( .A(y[3130]), .B(x[3130]), .Z(n7885) );
  XOR U12113 ( .A(y[3129]), .B(x[3129]), .Z(n7883) );
  XOR U12114 ( .A(n7877), .B(n7876), .Z(n7887) );
  XOR U12115 ( .A(n7879), .B(n7878), .Z(n7876) );
  XOR U12116 ( .A(y[3128]), .B(x[3128]), .Z(n7878) );
  XOR U12117 ( .A(y[3127]), .B(x[3127]), .Z(n7879) );
  XOR U12118 ( .A(y[3126]), .B(x[3126]), .Z(n7877) );
  NAND U12119 ( .A(n7940), .B(n7941), .Z(N29493) );
  NAND U12120 ( .A(n7942), .B(n7943), .Z(n7941) );
  NANDN U12121 ( .A(n7944), .B(n7945), .Z(n7943) );
  NANDN U12122 ( .A(n7945), .B(n7944), .Z(n7940) );
  XOR U12123 ( .A(n7944), .B(n7946), .Z(N29492) );
  XNOR U12124 ( .A(n7942), .B(n7945), .Z(n7946) );
  NAND U12125 ( .A(n7947), .B(n7948), .Z(n7945) );
  NAND U12126 ( .A(n7949), .B(n7950), .Z(n7948) );
  NANDN U12127 ( .A(n7951), .B(n7952), .Z(n7950) );
  NANDN U12128 ( .A(n7952), .B(n7951), .Z(n7947) );
  AND U12129 ( .A(n7953), .B(n7954), .Z(n7942) );
  NAND U12130 ( .A(n7955), .B(n7956), .Z(n7954) );
  OR U12131 ( .A(n7957), .B(n7958), .Z(n7956) );
  NAND U12132 ( .A(n7958), .B(n7957), .Z(n7953) );
  IV U12133 ( .A(n7959), .Z(n7958) );
  AND U12134 ( .A(n7960), .B(n7961), .Z(n7944) );
  NAND U12135 ( .A(n7962), .B(n7963), .Z(n7961) );
  NANDN U12136 ( .A(n7964), .B(n7965), .Z(n7963) );
  NANDN U12137 ( .A(n7965), .B(n7964), .Z(n7960) );
  XOR U12138 ( .A(n7957), .B(n7966), .Z(N29491) );
  XOR U12139 ( .A(n7955), .B(n7959), .Z(n7966) );
  XNOR U12140 ( .A(n7952), .B(n7967), .Z(n7959) );
  XNOR U12141 ( .A(n7949), .B(n7951), .Z(n7967) );
  AND U12142 ( .A(n7968), .B(n7969), .Z(n7951) );
  NANDN U12143 ( .A(n7970), .B(n7971), .Z(n7969) );
  NANDN U12144 ( .A(n7972), .B(n7973), .Z(n7971) );
  IV U12145 ( .A(n7974), .Z(n7973) );
  NAND U12146 ( .A(n7974), .B(n7972), .Z(n7968) );
  AND U12147 ( .A(n7975), .B(n7976), .Z(n7949) );
  NAND U12148 ( .A(n7977), .B(n7978), .Z(n7976) );
  OR U12149 ( .A(n7979), .B(n7980), .Z(n7978) );
  NAND U12150 ( .A(n7980), .B(n7979), .Z(n7975) );
  IV U12151 ( .A(n7981), .Z(n7980) );
  NAND U12152 ( .A(n7982), .B(n7983), .Z(n7952) );
  NANDN U12153 ( .A(n7984), .B(n7985), .Z(n7983) );
  NAND U12154 ( .A(n7986), .B(n7987), .Z(n7985) );
  OR U12155 ( .A(n7987), .B(n7986), .Z(n7982) );
  IV U12156 ( .A(n7988), .Z(n7986) );
  AND U12157 ( .A(n7989), .B(n7990), .Z(n7955) );
  NAND U12158 ( .A(n7991), .B(n7992), .Z(n7990) );
  NANDN U12159 ( .A(n7993), .B(n7994), .Z(n7992) );
  NANDN U12160 ( .A(n7994), .B(n7993), .Z(n7989) );
  XOR U12161 ( .A(n7965), .B(n7995), .Z(n7957) );
  XNOR U12162 ( .A(n7962), .B(n7964), .Z(n7995) );
  AND U12163 ( .A(n7996), .B(n7997), .Z(n7964) );
  NANDN U12164 ( .A(n7998), .B(n7999), .Z(n7997) );
  NANDN U12165 ( .A(n8000), .B(n8001), .Z(n7999) );
  IV U12166 ( .A(n8002), .Z(n8001) );
  NAND U12167 ( .A(n8002), .B(n8000), .Z(n7996) );
  AND U12168 ( .A(n8003), .B(n8004), .Z(n7962) );
  NAND U12169 ( .A(n8005), .B(n8006), .Z(n8004) );
  OR U12170 ( .A(n8007), .B(n8008), .Z(n8006) );
  NAND U12171 ( .A(n8008), .B(n8007), .Z(n8003) );
  IV U12172 ( .A(n8009), .Z(n8008) );
  NAND U12173 ( .A(n8010), .B(n8011), .Z(n7965) );
  NANDN U12174 ( .A(n8012), .B(n8013), .Z(n8011) );
  NAND U12175 ( .A(n8014), .B(n8015), .Z(n8013) );
  OR U12176 ( .A(n8015), .B(n8014), .Z(n8010) );
  IV U12177 ( .A(n8016), .Z(n8014) );
  XOR U12178 ( .A(n7991), .B(n8017), .Z(N29490) );
  XNOR U12179 ( .A(n7994), .B(n7993), .Z(n8017) );
  XNOR U12180 ( .A(n8005), .B(n8018), .Z(n7993) );
  XOR U12181 ( .A(n8009), .B(n8007), .Z(n8018) );
  XOR U12182 ( .A(n8015), .B(n8019), .Z(n8007) );
  XOR U12183 ( .A(n8012), .B(n8016), .Z(n8019) );
  NAND U12184 ( .A(n8020), .B(n8021), .Z(n8016) );
  NAND U12185 ( .A(n8022), .B(n8023), .Z(n8021) );
  NAND U12186 ( .A(n8024), .B(n8025), .Z(n8020) );
  AND U12187 ( .A(n8026), .B(n8027), .Z(n8012) );
  NAND U12188 ( .A(n8028), .B(n8029), .Z(n8027) );
  NAND U12189 ( .A(n8030), .B(n8031), .Z(n8026) );
  NANDN U12190 ( .A(n8032), .B(n8033), .Z(n8015) );
  NANDN U12191 ( .A(n8034), .B(n8035), .Z(n8009) );
  XNOR U12192 ( .A(n8000), .B(n8036), .Z(n8005) );
  XOR U12193 ( .A(n7998), .B(n8002), .Z(n8036) );
  NAND U12194 ( .A(n8037), .B(n8038), .Z(n8002) );
  NAND U12195 ( .A(n8039), .B(n8040), .Z(n8038) );
  NAND U12196 ( .A(n8041), .B(n8042), .Z(n8037) );
  AND U12197 ( .A(n8043), .B(n8044), .Z(n7998) );
  NAND U12198 ( .A(n8045), .B(n8046), .Z(n8044) );
  NAND U12199 ( .A(n8047), .B(n8048), .Z(n8043) );
  AND U12200 ( .A(n8049), .B(n8050), .Z(n8000) );
  NAND U12201 ( .A(n8051), .B(n8052), .Z(n7994) );
  XNOR U12202 ( .A(n7977), .B(n8053), .Z(n7991) );
  XOR U12203 ( .A(n7981), .B(n7979), .Z(n8053) );
  XOR U12204 ( .A(n7987), .B(n8054), .Z(n7979) );
  XOR U12205 ( .A(n7984), .B(n7988), .Z(n8054) );
  NAND U12206 ( .A(n8055), .B(n8056), .Z(n7988) );
  NAND U12207 ( .A(n8057), .B(n8058), .Z(n8056) );
  NAND U12208 ( .A(n8059), .B(n8060), .Z(n8055) );
  AND U12209 ( .A(n8061), .B(n8062), .Z(n7984) );
  NAND U12210 ( .A(n8063), .B(n8064), .Z(n8062) );
  NAND U12211 ( .A(n8065), .B(n8066), .Z(n8061) );
  NANDN U12212 ( .A(n8067), .B(n8068), .Z(n7987) );
  NANDN U12213 ( .A(n8069), .B(n8070), .Z(n7981) );
  XNOR U12214 ( .A(n7972), .B(n8071), .Z(n7977) );
  XOR U12215 ( .A(n7970), .B(n7974), .Z(n8071) );
  NAND U12216 ( .A(n8072), .B(n8073), .Z(n7974) );
  NAND U12217 ( .A(n8074), .B(n8075), .Z(n8073) );
  NAND U12218 ( .A(n8076), .B(n8077), .Z(n8072) );
  AND U12219 ( .A(n8078), .B(n8079), .Z(n7970) );
  NAND U12220 ( .A(n8080), .B(n8081), .Z(n8079) );
  NAND U12221 ( .A(n8082), .B(n8083), .Z(n8078) );
  AND U12222 ( .A(n8084), .B(n8085), .Z(n7972) );
  XOR U12223 ( .A(n8052), .B(n8051), .Z(N29489) );
  XNOR U12224 ( .A(n8070), .B(n8069), .Z(n8051) );
  XNOR U12225 ( .A(n8084), .B(n8085), .Z(n8069) );
  XOR U12226 ( .A(n8081), .B(n8080), .Z(n8085) );
  XOR U12227 ( .A(y[3123]), .B(x[3123]), .Z(n8080) );
  XOR U12228 ( .A(n8083), .B(n8082), .Z(n8081) );
  XOR U12229 ( .A(y[3125]), .B(x[3125]), .Z(n8082) );
  XOR U12230 ( .A(y[3124]), .B(x[3124]), .Z(n8083) );
  XOR U12231 ( .A(n8075), .B(n8074), .Z(n8084) );
  XOR U12232 ( .A(n8077), .B(n8076), .Z(n8074) );
  XOR U12233 ( .A(y[3122]), .B(x[3122]), .Z(n8076) );
  XOR U12234 ( .A(y[3121]), .B(x[3121]), .Z(n8077) );
  XOR U12235 ( .A(y[3120]), .B(x[3120]), .Z(n8075) );
  XNOR U12236 ( .A(n8068), .B(n8067), .Z(n8070) );
  XNOR U12237 ( .A(n8064), .B(n8063), .Z(n8067) );
  XOR U12238 ( .A(n8066), .B(n8065), .Z(n8063) );
  XOR U12239 ( .A(y[3119]), .B(x[3119]), .Z(n8065) );
  XOR U12240 ( .A(y[3118]), .B(x[3118]), .Z(n8066) );
  XOR U12241 ( .A(y[3117]), .B(x[3117]), .Z(n8064) );
  XOR U12242 ( .A(n8058), .B(n8057), .Z(n8068) );
  XOR U12243 ( .A(n8060), .B(n8059), .Z(n8057) );
  XOR U12244 ( .A(y[3116]), .B(x[3116]), .Z(n8059) );
  XOR U12245 ( .A(y[3115]), .B(x[3115]), .Z(n8060) );
  XOR U12246 ( .A(y[3114]), .B(x[3114]), .Z(n8058) );
  XNOR U12247 ( .A(n8035), .B(n8034), .Z(n8052) );
  XNOR U12248 ( .A(n8049), .B(n8050), .Z(n8034) );
  XOR U12249 ( .A(n8046), .B(n8045), .Z(n8050) );
  XOR U12250 ( .A(y[3111]), .B(x[3111]), .Z(n8045) );
  XOR U12251 ( .A(n8048), .B(n8047), .Z(n8046) );
  XOR U12252 ( .A(y[3113]), .B(x[3113]), .Z(n8047) );
  XOR U12253 ( .A(y[3112]), .B(x[3112]), .Z(n8048) );
  XOR U12254 ( .A(n8040), .B(n8039), .Z(n8049) );
  XOR U12255 ( .A(n8042), .B(n8041), .Z(n8039) );
  XOR U12256 ( .A(y[3110]), .B(x[3110]), .Z(n8041) );
  XOR U12257 ( .A(y[3109]), .B(x[3109]), .Z(n8042) );
  XOR U12258 ( .A(y[3108]), .B(x[3108]), .Z(n8040) );
  XNOR U12259 ( .A(n8033), .B(n8032), .Z(n8035) );
  XNOR U12260 ( .A(n8029), .B(n8028), .Z(n8032) );
  XOR U12261 ( .A(n8031), .B(n8030), .Z(n8028) );
  XOR U12262 ( .A(y[3107]), .B(x[3107]), .Z(n8030) );
  XOR U12263 ( .A(y[3106]), .B(x[3106]), .Z(n8031) );
  XOR U12264 ( .A(y[3105]), .B(x[3105]), .Z(n8029) );
  XOR U12265 ( .A(n8023), .B(n8022), .Z(n8033) );
  XOR U12266 ( .A(n8025), .B(n8024), .Z(n8022) );
  XOR U12267 ( .A(y[3104]), .B(x[3104]), .Z(n8024) );
  XOR U12268 ( .A(y[3103]), .B(x[3103]), .Z(n8025) );
  XOR U12269 ( .A(y[3102]), .B(x[3102]), .Z(n8023) );
  NAND U12270 ( .A(n8086), .B(n8087), .Z(N29481) );
  NAND U12271 ( .A(n8088), .B(n8089), .Z(n8087) );
  NANDN U12272 ( .A(n8090), .B(n8091), .Z(n8089) );
  NANDN U12273 ( .A(n8091), .B(n8090), .Z(n8086) );
  XOR U12274 ( .A(n8090), .B(n8092), .Z(N29480) );
  XNOR U12275 ( .A(n8088), .B(n8091), .Z(n8092) );
  NAND U12276 ( .A(n8093), .B(n8094), .Z(n8091) );
  NAND U12277 ( .A(n8095), .B(n8096), .Z(n8094) );
  NANDN U12278 ( .A(n8097), .B(n8098), .Z(n8096) );
  NANDN U12279 ( .A(n8098), .B(n8097), .Z(n8093) );
  AND U12280 ( .A(n8099), .B(n8100), .Z(n8088) );
  NAND U12281 ( .A(n8101), .B(n8102), .Z(n8100) );
  OR U12282 ( .A(n8103), .B(n8104), .Z(n8102) );
  NAND U12283 ( .A(n8104), .B(n8103), .Z(n8099) );
  IV U12284 ( .A(n8105), .Z(n8104) );
  AND U12285 ( .A(n8106), .B(n8107), .Z(n8090) );
  NAND U12286 ( .A(n8108), .B(n8109), .Z(n8107) );
  NANDN U12287 ( .A(n8110), .B(n8111), .Z(n8109) );
  NANDN U12288 ( .A(n8111), .B(n8110), .Z(n8106) );
  XOR U12289 ( .A(n8103), .B(n8112), .Z(N29479) );
  XOR U12290 ( .A(n8101), .B(n8105), .Z(n8112) );
  XNOR U12291 ( .A(n8098), .B(n8113), .Z(n8105) );
  XNOR U12292 ( .A(n8095), .B(n8097), .Z(n8113) );
  AND U12293 ( .A(n8114), .B(n8115), .Z(n8097) );
  NANDN U12294 ( .A(n8116), .B(n8117), .Z(n8115) );
  NANDN U12295 ( .A(n8118), .B(n8119), .Z(n8117) );
  IV U12296 ( .A(n8120), .Z(n8119) );
  NAND U12297 ( .A(n8120), .B(n8118), .Z(n8114) );
  AND U12298 ( .A(n8121), .B(n8122), .Z(n8095) );
  NAND U12299 ( .A(n8123), .B(n8124), .Z(n8122) );
  OR U12300 ( .A(n8125), .B(n8126), .Z(n8124) );
  NAND U12301 ( .A(n8126), .B(n8125), .Z(n8121) );
  IV U12302 ( .A(n8127), .Z(n8126) );
  NAND U12303 ( .A(n8128), .B(n8129), .Z(n8098) );
  NANDN U12304 ( .A(n8130), .B(n8131), .Z(n8129) );
  NAND U12305 ( .A(n8132), .B(n8133), .Z(n8131) );
  OR U12306 ( .A(n8133), .B(n8132), .Z(n8128) );
  IV U12307 ( .A(n8134), .Z(n8132) );
  AND U12308 ( .A(n8135), .B(n8136), .Z(n8101) );
  NAND U12309 ( .A(n8137), .B(n8138), .Z(n8136) );
  NANDN U12310 ( .A(n8139), .B(n8140), .Z(n8138) );
  NANDN U12311 ( .A(n8140), .B(n8139), .Z(n8135) );
  XOR U12312 ( .A(n8111), .B(n8141), .Z(n8103) );
  XNOR U12313 ( .A(n8108), .B(n8110), .Z(n8141) );
  AND U12314 ( .A(n8142), .B(n8143), .Z(n8110) );
  NANDN U12315 ( .A(n8144), .B(n8145), .Z(n8143) );
  NANDN U12316 ( .A(n8146), .B(n8147), .Z(n8145) );
  IV U12317 ( .A(n8148), .Z(n8147) );
  NAND U12318 ( .A(n8148), .B(n8146), .Z(n8142) );
  AND U12319 ( .A(n8149), .B(n8150), .Z(n8108) );
  NAND U12320 ( .A(n8151), .B(n8152), .Z(n8150) );
  OR U12321 ( .A(n8153), .B(n8154), .Z(n8152) );
  NAND U12322 ( .A(n8154), .B(n8153), .Z(n8149) );
  IV U12323 ( .A(n8155), .Z(n8154) );
  NAND U12324 ( .A(n8156), .B(n8157), .Z(n8111) );
  NANDN U12325 ( .A(n8158), .B(n8159), .Z(n8157) );
  NAND U12326 ( .A(n8160), .B(n8161), .Z(n8159) );
  OR U12327 ( .A(n8161), .B(n8160), .Z(n8156) );
  IV U12328 ( .A(n8162), .Z(n8160) );
  XOR U12329 ( .A(n8137), .B(n8163), .Z(N29478) );
  XNOR U12330 ( .A(n8140), .B(n8139), .Z(n8163) );
  XNOR U12331 ( .A(n8151), .B(n8164), .Z(n8139) );
  XOR U12332 ( .A(n8155), .B(n8153), .Z(n8164) );
  XOR U12333 ( .A(n8161), .B(n8165), .Z(n8153) );
  XOR U12334 ( .A(n8158), .B(n8162), .Z(n8165) );
  NAND U12335 ( .A(n8166), .B(n8167), .Z(n8162) );
  NAND U12336 ( .A(n8168), .B(n8169), .Z(n8167) );
  NAND U12337 ( .A(n8170), .B(n8171), .Z(n8166) );
  AND U12338 ( .A(n8172), .B(n8173), .Z(n8158) );
  NAND U12339 ( .A(n8174), .B(n8175), .Z(n8173) );
  NAND U12340 ( .A(n8176), .B(n8177), .Z(n8172) );
  NANDN U12341 ( .A(n8178), .B(n8179), .Z(n8161) );
  NANDN U12342 ( .A(n8180), .B(n8181), .Z(n8155) );
  XNOR U12343 ( .A(n8146), .B(n8182), .Z(n8151) );
  XOR U12344 ( .A(n8144), .B(n8148), .Z(n8182) );
  NAND U12345 ( .A(n8183), .B(n8184), .Z(n8148) );
  NAND U12346 ( .A(n8185), .B(n8186), .Z(n8184) );
  NAND U12347 ( .A(n8187), .B(n8188), .Z(n8183) );
  AND U12348 ( .A(n8189), .B(n8190), .Z(n8144) );
  NAND U12349 ( .A(n8191), .B(n8192), .Z(n8190) );
  NAND U12350 ( .A(n8193), .B(n8194), .Z(n8189) );
  AND U12351 ( .A(n8195), .B(n8196), .Z(n8146) );
  NAND U12352 ( .A(n8197), .B(n8198), .Z(n8140) );
  XNOR U12353 ( .A(n8123), .B(n8199), .Z(n8137) );
  XOR U12354 ( .A(n8127), .B(n8125), .Z(n8199) );
  XOR U12355 ( .A(n8133), .B(n8200), .Z(n8125) );
  XOR U12356 ( .A(n8130), .B(n8134), .Z(n8200) );
  NAND U12357 ( .A(n8201), .B(n8202), .Z(n8134) );
  NAND U12358 ( .A(n8203), .B(n8204), .Z(n8202) );
  NAND U12359 ( .A(n8205), .B(n8206), .Z(n8201) );
  AND U12360 ( .A(n8207), .B(n8208), .Z(n8130) );
  NAND U12361 ( .A(n8209), .B(n8210), .Z(n8208) );
  NAND U12362 ( .A(n8211), .B(n8212), .Z(n8207) );
  NANDN U12363 ( .A(n8213), .B(n8214), .Z(n8133) );
  NANDN U12364 ( .A(n8215), .B(n8216), .Z(n8127) );
  XNOR U12365 ( .A(n8118), .B(n8217), .Z(n8123) );
  XOR U12366 ( .A(n8116), .B(n8120), .Z(n8217) );
  NAND U12367 ( .A(n8218), .B(n8219), .Z(n8120) );
  NAND U12368 ( .A(n8220), .B(n8221), .Z(n8219) );
  NAND U12369 ( .A(n8222), .B(n8223), .Z(n8218) );
  AND U12370 ( .A(n8224), .B(n8225), .Z(n8116) );
  NAND U12371 ( .A(n8226), .B(n8227), .Z(n8225) );
  NAND U12372 ( .A(n8228), .B(n8229), .Z(n8224) );
  AND U12373 ( .A(n8230), .B(n8231), .Z(n8118) );
  XOR U12374 ( .A(n8198), .B(n8197), .Z(N29477) );
  XNOR U12375 ( .A(n8216), .B(n8215), .Z(n8197) );
  XNOR U12376 ( .A(n8230), .B(n8231), .Z(n8215) );
  XOR U12377 ( .A(n8227), .B(n8226), .Z(n8231) );
  XOR U12378 ( .A(y[3099]), .B(x[3099]), .Z(n8226) );
  XOR U12379 ( .A(n8229), .B(n8228), .Z(n8227) );
  XOR U12380 ( .A(y[3101]), .B(x[3101]), .Z(n8228) );
  XOR U12381 ( .A(y[3100]), .B(x[3100]), .Z(n8229) );
  XOR U12382 ( .A(n8221), .B(n8220), .Z(n8230) );
  XOR U12383 ( .A(n8223), .B(n8222), .Z(n8220) );
  XOR U12384 ( .A(y[3098]), .B(x[3098]), .Z(n8222) );
  XOR U12385 ( .A(y[3097]), .B(x[3097]), .Z(n8223) );
  XOR U12386 ( .A(y[3096]), .B(x[3096]), .Z(n8221) );
  XNOR U12387 ( .A(n8214), .B(n8213), .Z(n8216) );
  XNOR U12388 ( .A(n8210), .B(n8209), .Z(n8213) );
  XOR U12389 ( .A(n8212), .B(n8211), .Z(n8209) );
  XOR U12390 ( .A(y[3095]), .B(x[3095]), .Z(n8211) );
  XOR U12391 ( .A(y[3094]), .B(x[3094]), .Z(n8212) );
  XOR U12392 ( .A(y[3093]), .B(x[3093]), .Z(n8210) );
  XOR U12393 ( .A(n8204), .B(n8203), .Z(n8214) );
  XOR U12394 ( .A(n8206), .B(n8205), .Z(n8203) );
  XOR U12395 ( .A(y[3092]), .B(x[3092]), .Z(n8205) );
  XOR U12396 ( .A(y[3091]), .B(x[3091]), .Z(n8206) );
  XOR U12397 ( .A(y[3090]), .B(x[3090]), .Z(n8204) );
  XNOR U12398 ( .A(n8181), .B(n8180), .Z(n8198) );
  XNOR U12399 ( .A(n8195), .B(n8196), .Z(n8180) );
  XOR U12400 ( .A(n8192), .B(n8191), .Z(n8196) );
  XOR U12401 ( .A(y[3087]), .B(x[3087]), .Z(n8191) );
  XOR U12402 ( .A(n8194), .B(n8193), .Z(n8192) );
  XOR U12403 ( .A(y[3089]), .B(x[3089]), .Z(n8193) );
  XOR U12404 ( .A(y[3088]), .B(x[3088]), .Z(n8194) );
  XOR U12405 ( .A(n8186), .B(n8185), .Z(n8195) );
  XOR U12406 ( .A(n8188), .B(n8187), .Z(n8185) );
  XOR U12407 ( .A(y[3086]), .B(x[3086]), .Z(n8187) );
  XOR U12408 ( .A(y[3085]), .B(x[3085]), .Z(n8188) );
  XOR U12409 ( .A(y[3084]), .B(x[3084]), .Z(n8186) );
  XNOR U12410 ( .A(n8179), .B(n8178), .Z(n8181) );
  XNOR U12411 ( .A(n8175), .B(n8174), .Z(n8178) );
  XOR U12412 ( .A(n8177), .B(n8176), .Z(n8174) );
  XOR U12413 ( .A(y[3083]), .B(x[3083]), .Z(n8176) );
  XOR U12414 ( .A(y[3082]), .B(x[3082]), .Z(n8177) );
  XOR U12415 ( .A(y[3081]), .B(x[3081]), .Z(n8175) );
  XOR U12416 ( .A(n8169), .B(n8168), .Z(n8179) );
  XOR U12417 ( .A(n8171), .B(n8170), .Z(n8168) );
  XOR U12418 ( .A(y[3080]), .B(x[3080]), .Z(n8170) );
  XOR U12419 ( .A(y[3079]), .B(x[3079]), .Z(n8171) );
  XOR U12420 ( .A(y[3078]), .B(x[3078]), .Z(n8169) );
  NAND U12421 ( .A(n8232), .B(n8233), .Z(N29469) );
  NAND U12422 ( .A(n8234), .B(n8235), .Z(n8233) );
  NANDN U12423 ( .A(n8236), .B(n8237), .Z(n8235) );
  NANDN U12424 ( .A(n8237), .B(n8236), .Z(n8232) );
  XOR U12425 ( .A(n8236), .B(n8238), .Z(N29468) );
  XNOR U12426 ( .A(n8234), .B(n8237), .Z(n8238) );
  NAND U12427 ( .A(n8239), .B(n8240), .Z(n8237) );
  NAND U12428 ( .A(n8241), .B(n8242), .Z(n8240) );
  NANDN U12429 ( .A(n8243), .B(n8244), .Z(n8242) );
  NANDN U12430 ( .A(n8244), .B(n8243), .Z(n8239) );
  AND U12431 ( .A(n8245), .B(n8246), .Z(n8234) );
  NAND U12432 ( .A(n8247), .B(n8248), .Z(n8246) );
  OR U12433 ( .A(n8249), .B(n8250), .Z(n8248) );
  NAND U12434 ( .A(n8250), .B(n8249), .Z(n8245) );
  IV U12435 ( .A(n8251), .Z(n8250) );
  AND U12436 ( .A(n8252), .B(n8253), .Z(n8236) );
  NAND U12437 ( .A(n8254), .B(n8255), .Z(n8253) );
  NANDN U12438 ( .A(n8256), .B(n8257), .Z(n8255) );
  NANDN U12439 ( .A(n8257), .B(n8256), .Z(n8252) );
  XOR U12440 ( .A(n8249), .B(n8258), .Z(N29467) );
  XOR U12441 ( .A(n8247), .B(n8251), .Z(n8258) );
  XNOR U12442 ( .A(n8244), .B(n8259), .Z(n8251) );
  XNOR U12443 ( .A(n8241), .B(n8243), .Z(n8259) );
  AND U12444 ( .A(n8260), .B(n8261), .Z(n8243) );
  NANDN U12445 ( .A(n8262), .B(n8263), .Z(n8261) );
  NANDN U12446 ( .A(n8264), .B(n8265), .Z(n8263) );
  IV U12447 ( .A(n8266), .Z(n8265) );
  NAND U12448 ( .A(n8266), .B(n8264), .Z(n8260) );
  AND U12449 ( .A(n8267), .B(n8268), .Z(n8241) );
  NAND U12450 ( .A(n8269), .B(n8270), .Z(n8268) );
  OR U12451 ( .A(n8271), .B(n8272), .Z(n8270) );
  NAND U12452 ( .A(n8272), .B(n8271), .Z(n8267) );
  IV U12453 ( .A(n8273), .Z(n8272) );
  NAND U12454 ( .A(n8274), .B(n8275), .Z(n8244) );
  NANDN U12455 ( .A(n8276), .B(n8277), .Z(n8275) );
  NAND U12456 ( .A(n8278), .B(n8279), .Z(n8277) );
  OR U12457 ( .A(n8279), .B(n8278), .Z(n8274) );
  IV U12458 ( .A(n8280), .Z(n8278) );
  AND U12459 ( .A(n8281), .B(n8282), .Z(n8247) );
  NAND U12460 ( .A(n8283), .B(n8284), .Z(n8282) );
  NANDN U12461 ( .A(n8285), .B(n8286), .Z(n8284) );
  NANDN U12462 ( .A(n8286), .B(n8285), .Z(n8281) );
  XOR U12463 ( .A(n8257), .B(n8287), .Z(n8249) );
  XNOR U12464 ( .A(n8254), .B(n8256), .Z(n8287) );
  AND U12465 ( .A(n8288), .B(n8289), .Z(n8256) );
  NANDN U12466 ( .A(n8290), .B(n8291), .Z(n8289) );
  NANDN U12467 ( .A(n8292), .B(n8293), .Z(n8291) );
  IV U12468 ( .A(n8294), .Z(n8293) );
  NAND U12469 ( .A(n8294), .B(n8292), .Z(n8288) );
  AND U12470 ( .A(n8295), .B(n8296), .Z(n8254) );
  NAND U12471 ( .A(n8297), .B(n8298), .Z(n8296) );
  OR U12472 ( .A(n8299), .B(n8300), .Z(n8298) );
  NAND U12473 ( .A(n8300), .B(n8299), .Z(n8295) );
  IV U12474 ( .A(n8301), .Z(n8300) );
  NAND U12475 ( .A(n8302), .B(n8303), .Z(n8257) );
  NANDN U12476 ( .A(n8304), .B(n8305), .Z(n8303) );
  NAND U12477 ( .A(n8306), .B(n8307), .Z(n8305) );
  OR U12478 ( .A(n8307), .B(n8306), .Z(n8302) );
  IV U12479 ( .A(n8308), .Z(n8306) );
  XOR U12480 ( .A(n8283), .B(n8309), .Z(N29466) );
  XNOR U12481 ( .A(n8286), .B(n8285), .Z(n8309) );
  XNOR U12482 ( .A(n8297), .B(n8310), .Z(n8285) );
  XOR U12483 ( .A(n8301), .B(n8299), .Z(n8310) );
  XOR U12484 ( .A(n8307), .B(n8311), .Z(n8299) );
  XOR U12485 ( .A(n8304), .B(n8308), .Z(n8311) );
  NAND U12486 ( .A(n8312), .B(n8313), .Z(n8308) );
  NAND U12487 ( .A(n8314), .B(n8315), .Z(n8313) );
  NAND U12488 ( .A(n8316), .B(n8317), .Z(n8312) );
  AND U12489 ( .A(n8318), .B(n8319), .Z(n8304) );
  NAND U12490 ( .A(n8320), .B(n8321), .Z(n8319) );
  NAND U12491 ( .A(n8322), .B(n8323), .Z(n8318) );
  NANDN U12492 ( .A(n8324), .B(n8325), .Z(n8307) );
  NANDN U12493 ( .A(n8326), .B(n8327), .Z(n8301) );
  XNOR U12494 ( .A(n8292), .B(n8328), .Z(n8297) );
  XOR U12495 ( .A(n8290), .B(n8294), .Z(n8328) );
  NAND U12496 ( .A(n8329), .B(n8330), .Z(n8294) );
  NAND U12497 ( .A(n8331), .B(n8332), .Z(n8330) );
  NAND U12498 ( .A(n8333), .B(n8334), .Z(n8329) );
  AND U12499 ( .A(n8335), .B(n8336), .Z(n8290) );
  NAND U12500 ( .A(n8337), .B(n8338), .Z(n8336) );
  NAND U12501 ( .A(n8339), .B(n8340), .Z(n8335) );
  AND U12502 ( .A(n8341), .B(n8342), .Z(n8292) );
  NAND U12503 ( .A(n8343), .B(n8344), .Z(n8286) );
  XNOR U12504 ( .A(n8269), .B(n8345), .Z(n8283) );
  XOR U12505 ( .A(n8273), .B(n8271), .Z(n8345) );
  XOR U12506 ( .A(n8279), .B(n8346), .Z(n8271) );
  XOR U12507 ( .A(n8276), .B(n8280), .Z(n8346) );
  NAND U12508 ( .A(n8347), .B(n8348), .Z(n8280) );
  NAND U12509 ( .A(n8349), .B(n8350), .Z(n8348) );
  NAND U12510 ( .A(n8351), .B(n8352), .Z(n8347) );
  AND U12511 ( .A(n8353), .B(n8354), .Z(n8276) );
  NAND U12512 ( .A(n8355), .B(n8356), .Z(n8354) );
  NAND U12513 ( .A(n8357), .B(n8358), .Z(n8353) );
  NANDN U12514 ( .A(n8359), .B(n8360), .Z(n8279) );
  NANDN U12515 ( .A(n8361), .B(n8362), .Z(n8273) );
  XNOR U12516 ( .A(n8264), .B(n8363), .Z(n8269) );
  XOR U12517 ( .A(n8262), .B(n8266), .Z(n8363) );
  NAND U12518 ( .A(n8364), .B(n8365), .Z(n8266) );
  NAND U12519 ( .A(n8366), .B(n8367), .Z(n8365) );
  NAND U12520 ( .A(n8368), .B(n8369), .Z(n8364) );
  AND U12521 ( .A(n8370), .B(n8371), .Z(n8262) );
  NAND U12522 ( .A(n8372), .B(n8373), .Z(n8371) );
  NAND U12523 ( .A(n8374), .B(n8375), .Z(n8370) );
  AND U12524 ( .A(n8376), .B(n8377), .Z(n8264) );
  XOR U12525 ( .A(n8344), .B(n8343), .Z(N29465) );
  XNOR U12526 ( .A(n8362), .B(n8361), .Z(n8343) );
  XNOR U12527 ( .A(n8376), .B(n8377), .Z(n8361) );
  XOR U12528 ( .A(n8373), .B(n8372), .Z(n8377) );
  XOR U12529 ( .A(y[3075]), .B(x[3075]), .Z(n8372) );
  XOR U12530 ( .A(n8375), .B(n8374), .Z(n8373) );
  XOR U12531 ( .A(y[3077]), .B(x[3077]), .Z(n8374) );
  XOR U12532 ( .A(y[3076]), .B(x[3076]), .Z(n8375) );
  XOR U12533 ( .A(n8367), .B(n8366), .Z(n8376) );
  XOR U12534 ( .A(n8369), .B(n8368), .Z(n8366) );
  XOR U12535 ( .A(y[3074]), .B(x[3074]), .Z(n8368) );
  XOR U12536 ( .A(y[3073]), .B(x[3073]), .Z(n8369) );
  XOR U12537 ( .A(y[3072]), .B(x[3072]), .Z(n8367) );
  XNOR U12538 ( .A(n8360), .B(n8359), .Z(n8362) );
  XNOR U12539 ( .A(n8356), .B(n8355), .Z(n8359) );
  XOR U12540 ( .A(n8358), .B(n8357), .Z(n8355) );
  XOR U12541 ( .A(y[3071]), .B(x[3071]), .Z(n8357) );
  XOR U12542 ( .A(y[3070]), .B(x[3070]), .Z(n8358) );
  XOR U12543 ( .A(y[3069]), .B(x[3069]), .Z(n8356) );
  XOR U12544 ( .A(n8350), .B(n8349), .Z(n8360) );
  XOR U12545 ( .A(n8352), .B(n8351), .Z(n8349) );
  XOR U12546 ( .A(y[3068]), .B(x[3068]), .Z(n8351) );
  XOR U12547 ( .A(y[3067]), .B(x[3067]), .Z(n8352) );
  XOR U12548 ( .A(y[3066]), .B(x[3066]), .Z(n8350) );
  XNOR U12549 ( .A(n8327), .B(n8326), .Z(n8344) );
  XNOR U12550 ( .A(n8341), .B(n8342), .Z(n8326) );
  XOR U12551 ( .A(n8338), .B(n8337), .Z(n8342) );
  XOR U12552 ( .A(y[3063]), .B(x[3063]), .Z(n8337) );
  XOR U12553 ( .A(n8340), .B(n8339), .Z(n8338) );
  XOR U12554 ( .A(y[3065]), .B(x[3065]), .Z(n8339) );
  XOR U12555 ( .A(y[3064]), .B(x[3064]), .Z(n8340) );
  XOR U12556 ( .A(n8332), .B(n8331), .Z(n8341) );
  XOR U12557 ( .A(n8334), .B(n8333), .Z(n8331) );
  XOR U12558 ( .A(y[3062]), .B(x[3062]), .Z(n8333) );
  XOR U12559 ( .A(y[3061]), .B(x[3061]), .Z(n8334) );
  XOR U12560 ( .A(y[3060]), .B(x[3060]), .Z(n8332) );
  XNOR U12561 ( .A(n8325), .B(n8324), .Z(n8327) );
  XNOR U12562 ( .A(n8321), .B(n8320), .Z(n8324) );
  XOR U12563 ( .A(n8323), .B(n8322), .Z(n8320) );
  XOR U12564 ( .A(y[3059]), .B(x[3059]), .Z(n8322) );
  XOR U12565 ( .A(y[3058]), .B(x[3058]), .Z(n8323) );
  XOR U12566 ( .A(y[3057]), .B(x[3057]), .Z(n8321) );
  XOR U12567 ( .A(n8315), .B(n8314), .Z(n8325) );
  XOR U12568 ( .A(n8317), .B(n8316), .Z(n8314) );
  XOR U12569 ( .A(y[3056]), .B(x[3056]), .Z(n8316) );
  XOR U12570 ( .A(y[3055]), .B(x[3055]), .Z(n8317) );
  XOR U12571 ( .A(y[3054]), .B(x[3054]), .Z(n8315) );
  NAND U12572 ( .A(n8378), .B(n8379), .Z(N29457) );
  NAND U12573 ( .A(n8380), .B(n8381), .Z(n8379) );
  NANDN U12574 ( .A(n8382), .B(n8383), .Z(n8381) );
  NANDN U12575 ( .A(n8383), .B(n8382), .Z(n8378) );
  XOR U12576 ( .A(n8382), .B(n8384), .Z(N29456) );
  XNOR U12577 ( .A(n8380), .B(n8383), .Z(n8384) );
  NAND U12578 ( .A(n8385), .B(n8386), .Z(n8383) );
  NAND U12579 ( .A(n8387), .B(n8388), .Z(n8386) );
  NANDN U12580 ( .A(n8389), .B(n8390), .Z(n8388) );
  NANDN U12581 ( .A(n8390), .B(n8389), .Z(n8385) );
  AND U12582 ( .A(n8391), .B(n8392), .Z(n8380) );
  NAND U12583 ( .A(n8393), .B(n8394), .Z(n8392) );
  OR U12584 ( .A(n8395), .B(n8396), .Z(n8394) );
  NAND U12585 ( .A(n8396), .B(n8395), .Z(n8391) );
  IV U12586 ( .A(n8397), .Z(n8396) );
  AND U12587 ( .A(n8398), .B(n8399), .Z(n8382) );
  NAND U12588 ( .A(n8400), .B(n8401), .Z(n8399) );
  NANDN U12589 ( .A(n8402), .B(n8403), .Z(n8401) );
  NANDN U12590 ( .A(n8403), .B(n8402), .Z(n8398) );
  XOR U12591 ( .A(n8395), .B(n8404), .Z(N29455) );
  XOR U12592 ( .A(n8393), .B(n8397), .Z(n8404) );
  XNOR U12593 ( .A(n8390), .B(n8405), .Z(n8397) );
  XNOR U12594 ( .A(n8387), .B(n8389), .Z(n8405) );
  AND U12595 ( .A(n8406), .B(n8407), .Z(n8389) );
  NANDN U12596 ( .A(n8408), .B(n8409), .Z(n8407) );
  NANDN U12597 ( .A(n8410), .B(n8411), .Z(n8409) );
  IV U12598 ( .A(n8412), .Z(n8411) );
  NAND U12599 ( .A(n8412), .B(n8410), .Z(n8406) );
  AND U12600 ( .A(n8413), .B(n8414), .Z(n8387) );
  NAND U12601 ( .A(n8415), .B(n8416), .Z(n8414) );
  OR U12602 ( .A(n8417), .B(n8418), .Z(n8416) );
  NAND U12603 ( .A(n8418), .B(n8417), .Z(n8413) );
  IV U12604 ( .A(n8419), .Z(n8418) );
  NAND U12605 ( .A(n8420), .B(n8421), .Z(n8390) );
  NANDN U12606 ( .A(n8422), .B(n8423), .Z(n8421) );
  NAND U12607 ( .A(n8424), .B(n8425), .Z(n8423) );
  OR U12608 ( .A(n8425), .B(n8424), .Z(n8420) );
  IV U12609 ( .A(n8426), .Z(n8424) );
  AND U12610 ( .A(n8427), .B(n8428), .Z(n8393) );
  NAND U12611 ( .A(n8429), .B(n8430), .Z(n8428) );
  NANDN U12612 ( .A(n8431), .B(n8432), .Z(n8430) );
  NANDN U12613 ( .A(n8432), .B(n8431), .Z(n8427) );
  XOR U12614 ( .A(n8403), .B(n8433), .Z(n8395) );
  XNOR U12615 ( .A(n8400), .B(n8402), .Z(n8433) );
  AND U12616 ( .A(n8434), .B(n8435), .Z(n8402) );
  NANDN U12617 ( .A(n8436), .B(n8437), .Z(n8435) );
  NANDN U12618 ( .A(n8438), .B(n8439), .Z(n8437) );
  IV U12619 ( .A(n8440), .Z(n8439) );
  NAND U12620 ( .A(n8440), .B(n8438), .Z(n8434) );
  AND U12621 ( .A(n8441), .B(n8442), .Z(n8400) );
  NAND U12622 ( .A(n8443), .B(n8444), .Z(n8442) );
  OR U12623 ( .A(n8445), .B(n8446), .Z(n8444) );
  NAND U12624 ( .A(n8446), .B(n8445), .Z(n8441) );
  IV U12625 ( .A(n8447), .Z(n8446) );
  NAND U12626 ( .A(n8448), .B(n8449), .Z(n8403) );
  NANDN U12627 ( .A(n8450), .B(n8451), .Z(n8449) );
  NAND U12628 ( .A(n8452), .B(n8453), .Z(n8451) );
  OR U12629 ( .A(n8453), .B(n8452), .Z(n8448) );
  IV U12630 ( .A(n8454), .Z(n8452) );
  XOR U12631 ( .A(n8429), .B(n8455), .Z(N29454) );
  XNOR U12632 ( .A(n8432), .B(n8431), .Z(n8455) );
  XNOR U12633 ( .A(n8443), .B(n8456), .Z(n8431) );
  XOR U12634 ( .A(n8447), .B(n8445), .Z(n8456) );
  XOR U12635 ( .A(n8453), .B(n8457), .Z(n8445) );
  XOR U12636 ( .A(n8450), .B(n8454), .Z(n8457) );
  NAND U12637 ( .A(n8458), .B(n8459), .Z(n8454) );
  NAND U12638 ( .A(n8460), .B(n8461), .Z(n8459) );
  NAND U12639 ( .A(n8462), .B(n8463), .Z(n8458) );
  AND U12640 ( .A(n8464), .B(n8465), .Z(n8450) );
  NAND U12641 ( .A(n8466), .B(n8467), .Z(n8465) );
  NAND U12642 ( .A(n8468), .B(n8469), .Z(n8464) );
  NANDN U12643 ( .A(n8470), .B(n8471), .Z(n8453) );
  NANDN U12644 ( .A(n8472), .B(n8473), .Z(n8447) );
  XNOR U12645 ( .A(n8438), .B(n8474), .Z(n8443) );
  XOR U12646 ( .A(n8436), .B(n8440), .Z(n8474) );
  NAND U12647 ( .A(n8475), .B(n8476), .Z(n8440) );
  NAND U12648 ( .A(n8477), .B(n8478), .Z(n8476) );
  NAND U12649 ( .A(n8479), .B(n8480), .Z(n8475) );
  AND U12650 ( .A(n8481), .B(n8482), .Z(n8436) );
  NAND U12651 ( .A(n8483), .B(n8484), .Z(n8482) );
  NAND U12652 ( .A(n8485), .B(n8486), .Z(n8481) );
  AND U12653 ( .A(n8487), .B(n8488), .Z(n8438) );
  NAND U12654 ( .A(n8489), .B(n8490), .Z(n8432) );
  XNOR U12655 ( .A(n8415), .B(n8491), .Z(n8429) );
  XOR U12656 ( .A(n8419), .B(n8417), .Z(n8491) );
  XOR U12657 ( .A(n8425), .B(n8492), .Z(n8417) );
  XOR U12658 ( .A(n8422), .B(n8426), .Z(n8492) );
  NAND U12659 ( .A(n8493), .B(n8494), .Z(n8426) );
  NAND U12660 ( .A(n8495), .B(n8496), .Z(n8494) );
  NAND U12661 ( .A(n8497), .B(n8498), .Z(n8493) );
  AND U12662 ( .A(n8499), .B(n8500), .Z(n8422) );
  NAND U12663 ( .A(n8501), .B(n8502), .Z(n8500) );
  NAND U12664 ( .A(n8503), .B(n8504), .Z(n8499) );
  NANDN U12665 ( .A(n8505), .B(n8506), .Z(n8425) );
  NANDN U12666 ( .A(n8507), .B(n8508), .Z(n8419) );
  XNOR U12667 ( .A(n8410), .B(n8509), .Z(n8415) );
  XOR U12668 ( .A(n8408), .B(n8412), .Z(n8509) );
  NAND U12669 ( .A(n8510), .B(n8511), .Z(n8412) );
  NAND U12670 ( .A(n8512), .B(n8513), .Z(n8511) );
  NAND U12671 ( .A(n8514), .B(n8515), .Z(n8510) );
  AND U12672 ( .A(n8516), .B(n8517), .Z(n8408) );
  NAND U12673 ( .A(n8518), .B(n8519), .Z(n8517) );
  NAND U12674 ( .A(n8520), .B(n8521), .Z(n8516) );
  AND U12675 ( .A(n8522), .B(n8523), .Z(n8410) );
  XOR U12676 ( .A(n8490), .B(n8489), .Z(N29453) );
  XNOR U12677 ( .A(n8508), .B(n8507), .Z(n8489) );
  XNOR U12678 ( .A(n8522), .B(n8523), .Z(n8507) );
  XOR U12679 ( .A(n8519), .B(n8518), .Z(n8523) );
  XOR U12680 ( .A(y[3051]), .B(x[3051]), .Z(n8518) );
  XOR U12681 ( .A(n8521), .B(n8520), .Z(n8519) );
  XOR U12682 ( .A(y[3053]), .B(x[3053]), .Z(n8520) );
  XOR U12683 ( .A(y[3052]), .B(x[3052]), .Z(n8521) );
  XOR U12684 ( .A(n8513), .B(n8512), .Z(n8522) );
  XOR U12685 ( .A(n8515), .B(n8514), .Z(n8512) );
  XOR U12686 ( .A(y[3050]), .B(x[3050]), .Z(n8514) );
  XOR U12687 ( .A(y[3049]), .B(x[3049]), .Z(n8515) );
  XOR U12688 ( .A(y[3048]), .B(x[3048]), .Z(n8513) );
  XNOR U12689 ( .A(n8506), .B(n8505), .Z(n8508) );
  XNOR U12690 ( .A(n8502), .B(n8501), .Z(n8505) );
  XOR U12691 ( .A(n8504), .B(n8503), .Z(n8501) );
  XOR U12692 ( .A(y[3047]), .B(x[3047]), .Z(n8503) );
  XOR U12693 ( .A(y[3046]), .B(x[3046]), .Z(n8504) );
  XOR U12694 ( .A(y[3045]), .B(x[3045]), .Z(n8502) );
  XOR U12695 ( .A(n8496), .B(n8495), .Z(n8506) );
  XOR U12696 ( .A(n8498), .B(n8497), .Z(n8495) );
  XOR U12697 ( .A(y[3044]), .B(x[3044]), .Z(n8497) );
  XOR U12698 ( .A(y[3043]), .B(x[3043]), .Z(n8498) );
  XOR U12699 ( .A(y[3042]), .B(x[3042]), .Z(n8496) );
  XNOR U12700 ( .A(n8473), .B(n8472), .Z(n8490) );
  XNOR U12701 ( .A(n8487), .B(n8488), .Z(n8472) );
  XOR U12702 ( .A(n8484), .B(n8483), .Z(n8488) );
  XOR U12703 ( .A(y[3039]), .B(x[3039]), .Z(n8483) );
  XOR U12704 ( .A(n8486), .B(n8485), .Z(n8484) );
  XOR U12705 ( .A(y[3041]), .B(x[3041]), .Z(n8485) );
  XOR U12706 ( .A(y[3040]), .B(x[3040]), .Z(n8486) );
  XOR U12707 ( .A(n8478), .B(n8477), .Z(n8487) );
  XOR U12708 ( .A(n8480), .B(n8479), .Z(n8477) );
  XOR U12709 ( .A(y[3038]), .B(x[3038]), .Z(n8479) );
  XOR U12710 ( .A(y[3037]), .B(x[3037]), .Z(n8480) );
  XOR U12711 ( .A(y[3036]), .B(x[3036]), .Z(n8478) );
  XNOR U12712 ( .A(n8471), .B(n8470), .Z(n8473) );
  XNOR U12713 ( .A(n8467), .B(n8466), .Z(n8470) );
  XOR U12714 ( .A(n8469), .B(n8468), .Z(n8466) );
  XOR U12715 ( .A(y[3035]), .B(x[3035]), .Z(n8468) );
  XOR U12716 ( .A(y[3034]), .B(x[3034]), .Z(n8469) );
  XOR U12717 ( .A(y[3033]), .B(x[3033]), .Z(n8467) );
  XOR U12718 ( .A(n8461), .B(n8460), .Z(n8471) );
  XOR U12719 ( .A(n8463), .B(n8462), .Z(n8460) );
  XOR U12720 ( .A(y[3032]), .B(x[3032]), .Z(n8462) );
  XOR U12721 ( .A(y[3031]), .B(x[3031]), .Z(n8463) );
  XOR U12722 ( .A(y[3030]), .B(x[3030]), .Z(n8461) );
  NAND U12723 ( .A(n8524), .B(n8525), .Z(N29445) );
  NAND U12724 ( .A(n8526), .B(n8527), .Z(n8525) );
  NANDN U12725 ( .A(n8528), .B(n8529), .Z(n8527) );
  NANDN U12726 ( .A(n8529), .B(n8528), .Z(n8524) );
  XOR U12727 ( .A(n8528), .B(n8530), .Z(N29444) );
  XNOR U12728 ( .A(n8526), .B(n8529), .Z(n8530) );
  NAND U12729 ( .A(n8531), .B(n8532), .Z(n8529) );
  NAND U12730 ( .A(n8533), .B(n8534), .Z(n8532) );
  NANDN U12731 ( .A(n8535), .B(n8536), .Z(n8534) );
  NANDN U12732 ( .A(n8536), .B(n8535), .Z(n8531) );
  AND U12733 ( .A(n8537), .B(n8538), .Z(n8526) );
  NAND U12734 ( .A(n8539), .B(n8540), .Z(n8538) );
  OR U12735 ( .A(n8541), .B(n8542), .Z(n8540) );
  NAND U12736 ( .A(n8542), .B(n8541), .Z(n8537) );
  IV U12737 ( .A(n8543), .Z(n8542) );
  AND U12738 ( .A(n8544), .B(n8545), .Z(n8528) );
  NAND U12739 ( .A(n8546), .B(n8547), .Z(n8545) );
  NANDN U12740 ( .A(n8548), .B(n8549), .Z(n8547) );
  NANDN U12741 ( .A(n8549), .B(n8548), .Z(n8544) );
  XOR U12742 ( .A(n8541), .B(n8550), .Z(N29443) );
  XOR U12743 ( .A(n8539), .B(n8543), .Z(n8550) );
  XNOR U12744 ( .A(n8536), .B(n8551), .Z(n8543) );
  XNOR U12745 ( .A(n8533), .B(n8535), .Z(n8551) );
  AND U12746 ( .A(n8552), .B(n8553), .Z(n8535) );
  NANDN U12747 ( .A(n8554), .B(n8555), .Z(n8553) );
  NANDN U12748 ( .A(n8556), .B(n8557), .Z(n8555) );
  IV U12749 ( .A(n8558), .Z(n8557) );
  NAND U12750 ( .A(n8558), .B(n8556), .Z(n8552) );
  AND U12751 ( .A(n8559), .B(n8560), .Z(n8533) );
  NAND U12752 ( .A(n8561), .B(n8562), .Z(n8560) );
  OR U12753 ( .A(n8563), .B(n8564), .Z(n8562) );
  NAND U12754 ( .A(n8564), .B(n8563), .Z(n8559) );
  IV U12755 ( .A(n8565), .Z(n8564) );
  NAND U12756 ( .A(n8566), .B(n8567), .Z(n8536) );
  NANDN U12757 ( .A(n8568), .B(n8569), .Z(n8567) );
  NAND U12758 ( .A(n8570), .B(n8571), .Z(n8569) );
  OR U12759 ( .A(n8571), .B(n8570), .Z(n8566) );
  IV U12760 ( .A(n8572), .Z(n8570) );
  AND U12761 ( .A(n8573), .B(n8574), .Z(n8539) );
  NAND U12762 ( .A(n8575), .B(n8576), .Z(n8574) );
  NANDN U12763 ( .A(n8577), .B(n8578), .Z(n8576) );
  NANDN U12764 ( .A(n8578), .B(n8577), .Z(n8573) );
  XOR U12765 ( .A(n8549), .B(n8579), .Z(n8541) );
  XNOR U12766 ( .A(n8546), .B(n8548), .Z(n8579) );
  AND U12767 ( .A(n8580), .B(n8581), .Z(n8548) );
  NANDN U12768 ( .A(n8582), .B(n8583), .Z(n8581) );
  NANDN U12769 ( .A(n8584), .B(n8585), .Z(n8583) );
  IV U12770 ( .A(n8586), .Z(n8585) );
  NAND U12771 ( .A(n8586), .B(n8584), .Z(n8580) );
  AND U12772 ( .A(n8587), .B(n8588), .Z(n8546) );
  NAND U12773 ( .A(n8589), .B(n8590), .Z(n8588) );
  OR U12774 ( .A(n8591), .B(n8592), .Z(n8590) );
  NAND U12775 ( .A(n8592), .B(n8591), .Z(n8587) );
  IV U12776 ( .A(n8593), .Z(n8592) );
  NAND U12777 ( .A(n8594), .B(n8595), .Z(n8549) );
  NANDN U12778 ( .A(n8596), .B(n8597), .Z(n8595) );
  NAND U12779 ( .A(n8598), .B(n8599), .Z(n8597) );
  OR U12780 ( .A(n8599), .B(n8598), .Z(n8594) );
  IV U12781 ( .A(n8600), .Z(n8598) );
  XOR U12782 ( .A(n8575), .B(n8601), .Z(N29442) );
  XNOR U12783 ( .A(n8578), .B(n8577), .Z(n8601) );
  XNOR U12784 ( .A(n8589), .B(n8602), .Z(n8577) );
  XOR U12785 ( .A(n8593), .B(n8591), .Z(n8602) );
  XOR U12786 ( .A(n8599), .B(n8603), .Z(n8591) );
  XOR U12787 ( .A(n8596), .B(n8600), .Z(n8603) );
  NAND U12788 ( .A(n8604), .B(n8605), .Z(n8600) );
  NAND U12789 ( .A(n8606), .B(n8607), .Z(n8605) );
  NAND U12790 ( .A(n8608), .B(n8609), .Z(n8604) );
  AND U12791 ( .A(n8610), .B(n8611), .Z(n8596) );
  NAND U12792 ( .A(n8612), .B(n8613), .Z(n8611) );
  NAND U12793 ( .A(n8614), .B(n8615), .Z(n8610) );
  NANDN U12794 ( .A(n8616), .B(n8617), .Z(n8599) );
  NANDN U12795 ( .A(n8618), .B(n8619), .Z(n8593) );
  XNOR U12796 ( .A(n8584), .B(n8620), .Z(n8589) );
  XOR U12797 ( .A(n8582), .B(n8586), .Z(n8620) );
  NAND U12798 ( .A(n8621), .B(n8622), .Z(n8586) );
  NAND U12799 ( .A(n8623), .B(n8624), .Z(n8622) );
  NAND U12800 ( .A(n8625), .B(n8626), .Z(n8621) );
  AND U12801 ( .A(n8627), .B(n8628), .Z(n8582) );
  NAND U12802 ( .A(n8629), .B(n8630), .Z(n8628) );
  NAND U12803 ( .A(n8631), .B(n8632), .Z(n8627) );
  AND U12804 ( .A(n8633), .B(n8634), .Z(n8584) );
  NAND U12805 ( .A(n8635), .B(n8636), .Z(n8578) );
  XNOR U12806 ( .A(n8561), .B(n8637), .Z(n8575) );
  XOR U12807 ( .A(n8565), .B(n8563), .Z(n8637) );
  XOR U12808 ( .A(n8571), .B(n8638), .Z(n8563) );
  XOR U12809 ( .A(n8568), .B(n8572), .Z(n8638) );
  NAND U12810 ( .A(n8639), .B(n8640), .Z(n8572) );
  NAND U12811 ( .A(n8641), .B(n8642), .Z(n8640) );
  NAND U12812 ( .A(n8643), .B(n8644), .Z(n8639) );
  AND U12813 ( .A(n8645), .B(n8646), .Z(n8568) );
  NAND U12814 ( .A(n8647), .B(n8648), .Z(n8646) );
  NAND U12815 ( .A(n8649), .B(n8650), .Z(n8645) );
  NANDN U12816 ( .A(n8651), .B(n8652), .Z(n8571) );
  NANDN U12817 ( .A(n8653), .B(n8654), .Z(n8565) );
  XNOR U12818 ( .A(n8556), .B(n8655), .Z(n8561) );
  XOR U12819 ( .A(n8554), .B(n8558), .Z(n8655) );
  NAND U12820 ( .A(n8656), .B(n8657), .Z(n8558) );
  NAND U12821 ( .A(n8658), .B(n8659), .Z(n8657) );
  NAND U12822 ( .A(n8660), .B(n8661), .Z(n8656) );
  AND U12823 ( .A(n8662), .B(n8663), .Z(n8554) );
  NAND U12824 ( .A(n8664), .B(n8665), .Z(n8663) );
  NAND U12825 ( .A(n8666), .B(n8667), .Z(n8662) );
  AND U12826 ( .A(n8668), .B(n8669), .Z(n8556) );
  XOR U12827 ( .A(n8636), .B(n8635), .Z(N29441) );
  XNOR U12828 ( .A(n8654), .B(n8653), .Z(n8635) );
  XNOR U12829 ( .A(n8668), .B(n8669), .Z(n8653) );
  XOR U12830 ( .A(n8665), .B(n8664), .Z(n8669) );
  XOR U12831 ( .A(y[3027]), .B(x[3027]), .Z(n8664) );
  XOR U12832 ( .A(n8667), .B(n8666), .Z(n8665) );
  XOR U12833 ( .A(y[3029]), .B(x[3029]), .Z(n8666) );
  XOR U12834 ( .A(y[3028]), .B(x[3028]), .Z(n8667) );
  XOR U12835 ( .A(n8659), .B(n8658), .Z(n8668) );
  XOR U12836 ( .A(n8661), .B(n8660), .Z(n8658) );
  XOR U12837 ( .A(y[3026]), .B(x[3026]), .Z(n8660) );
  XOR U12838 ( .A(y[3025]), .B(x[3025]), .Z(n8661) );
  XOR U12839 ( .A(y[3024]), .B(x[3024]), .Z(n8659) );
  XNOR U12840 ( .A(n8652), .B(n8651), .Z(n8654) );
  XNOR U12841 ( .A(n8648), .B(n8647), .Z(n8651) );
  XOR U12842 ( .A(n8650), .B(n8649), .Z(n8647) );
  XOR U12843 ( .A(y[3023]), .B(x[3023]), .Z(n8649) );
  XOR U12844 ( .A(y[3022]), .B(x[3022]), .Z(n8650) );
  XOR U12845 ( .A(y[3021]), .B(x[3021]), .Z(n8648) );
  XOR U12846 ( .A(n8642), .B(n8641), .Z(n8652) );
  XOR U12847 ( .A(n8644), .B(n8643), .Z(n8641) );
  XOR U12848 ( .A(y[3020]), .B(x[3020]), .Z(n8643) );
  XOR U12849 ( .A(y[3019]), .B(x[3019]), .Z(n8644) );
  XOR U12850 ( .A(y[3018]), .B(x[3018]), .Z(n8642) );
  XNOR U12851 ( .A(n8619), .B(n8618), .Z(n8636) );
  XNOR U12852 ( .A(n8633), .B(n8634), .Z(n8618) );
  XOR U12853 ( .A(n8630), .B(n8629), .Z(n8634) );
  XOR U12854 ( .A(y[3015]), .B(x[3015]), .Z(n8629) );
  XOR U12855 ( .A(n8632), .B(n8631), .Z(n8630) );
  XOR U12856 ( .A(y[3017]), .B(x[3017]), .Z(n8631) );
  XOR U12857 ( .A(y[3016]), .B(x[3016]), .Z(n8632) );
  XOR U12858 ( .A(n8624), .B(n8623), .Z(n8633) );
  XOR U12859 ( .A(n8626), .B(n8625), .Z(n8623) );
  XOR U12860 ( .A(y[3014]), .B(x[3014]), .Z(n8625) );
  XOR U12861 ( .A(y[3013]), .B(x[3013]), .Z(n8626) );
  XOR U12862 ( .A(y[3012]), .B(x[3012]), .Z(n8624) );
  XNOR U12863 ( .A(n8617), .B(n8616), .Z(n8619) );
  XNOR U12864 ( .A(n8613), .B(n8612), .Z(n8616) );
  XOR U12865 ( .A(n8615), .B(n8614), .Z(n8612) );
  XOR U12866 ( .A(y[3011]), .B(x[3011]), .Z(n8614) );
  XOR U12867 ( .A(y[3010]), .B(x[3010]), .Z(n8615) );
  XOR U12868 ( .A(y[3009]), .B(x[3009]), .Z(n8613) );
  XOR U12869 ( .A(n8607), .B(n8606), .Z(n8617) );
  XOR U12870 ( .A(n8609), .B(n8608), .Z(n8606) );
  XOR U12871 ( .A(y[3008]), .B(x[3008]), .Z(n8608) );
  XOR U12872 ( .A(y[3007]), .B(x[3007]), .Z(n8609) );
  XOR U12873 ( .A(y[3006]), .B(x[3006]), .Z(n8607) );
  NAND U12874 ( .A(n8670), .B(n8671), .Z(N29433) );
  NAND U12875 ( .A(n8672), .B(n8673), .Z(n8671) );
  NANDN U12876 ( .A(n8674), .B(n8675), .Z(n8673) );
  NANDN U12877 ( .A(n8675), .B(n8674), .Z(n8670) );
  XOR U12878 ( .A(n8674), .B(n8676), .Z(N29432) );
  XNOR U12879 ( .A(n8672), .B(n8675), .Z(n8676) );
  NAND U12880 ( .A(n8677), .B(n8678), .Z(n8675) );
  NAND U12881 ( .A(n8679), .B(n8680), .Z(n8678) );
  NANDN U12882 ( .A(n8681), .B(n8682), .Z(n8680) );
  NANDN U12883 ( .A(n8682), .B(n8681), .Z(n8677) );
  AND U12884 ( .A(n8683), .B(n8684), .Z(n8672) );
  NAND U12885 ( .A(n8685), .B(n8686), .Z(n8684) );
  OR U12886 ( .A(n8687), .B(n8688), .Z(n8686) );
  NAND U12887 ( .A(n8688), .B(n8687), .Z(n8683) );
  IV U12888 ( .A(n8689), .Z(n8688) );
  AND U12889 ( .A(n8690), .B(n8691), .Z(n8674) );
  NAND U12890 ( .A(n8692), .B(n8693), .Z(n8691) );
  NANDN U12891 ( .A(n8694), .B(n8695), .Z(n8693) );
  NANDN U12892 ( .A(n8695), .B(n8694), .Z(n8690) );
  XOR U12893 ( .A(n8687), .B(n8696), .Z(N29431) );
  XOR U12894 ( .A(n8685), .B(n8689), .Z(n8696) );
  XNOR U12895 ( .A(n8682), .B(n8697), .Z(n8689) );
  XNOR U12896 ( .A(n8679), .B(n8681), .Z(n8697) );
  AND U12897 ( .A(n8698), .B(n8699), .Z(n8681) );
  NANDN U12898 ( .A(n8700), .B(n8701), .Z(n8699) );
  NANDN U12899 ( .A(n8702), .B(n8703), .Z(n8701) );
  IV U12900 ( .A(n8704), .Z(n8703) );
  NAND U12901 ( .A(n8704), .B(n8702), .Z(n8698) );
  AND U12902 ( .A(n8705), .B(n8706), .Z(n8679) );
  NAND U12903 ( .A(n8707), .B(n8708), .Z(n8706) );
  OR U12904 ( .A(n8709), .B(n8710), .Z(n8708) );
  NAND U12905 ( .A(n8710), .B(n8709), .Z(n8705) );
  IV U12906 ( .A(n8711), .Z(n8710) );
  NAND U12907 ( .A(n8712), .B(n8713), .Z(n8682) );
  NANDN U12908 ( .A(n8714), .B(n8715), .Z(n8713) );
  NAND U12909 ( .A(n8716), .B(n8717), .Z(n8715) );
  OR U12910 ( .A(n8717), .B(n8716), .Z(n8712) );
  IV U12911 ( .A(n8718), .Z(n8716) );
  AND U12912 ( .A(n8719), .B(n8720), .Z(n8685) );
  NAND U12913 ( .A(n8721), .B(n8722), .Z(n8720) );
  NANDN U12914 ( .A(n8723), .B(n8724), .Z(n8722) );
  NANDN U12915 ( .A(n8724), .B(n8723), .Z(n8719) );
  XOR U12916 ( .A(n8695), .B(n8725), .Z(n8687) );
  XNOR U12917 ( .A(n8692), .B(n8694), .Z(n8725) );
  AND U12918 ( .A(n8726), .B(n8727), .Z(n8694) );
  NANDN U12919 ( .A(n8728), .B(n8729), .Z(n8727) );
  NANDN U12920 ( .A(n8730), .B(n8731), .Z(n8729) );
  IV U12921 ( .A(n8732), .Z(n8731) );
  NAND U12922 ( .A(n8732), .B(n8730), .Z(n8726) );
  AND U12923 ( .A(n8733), .B(n8734), .Z(n8692) );
  NAND U12924 ( .A(n8735), .B(n8736), .Z(n8734) );
  OR U12925 ( .A(n8737), .B(n8738), .Z(n8736) );
  NAND U12926 ( .A(n8738), .B(n8737), .Z(n8733) );
  IV U12927 ( .A(n8739), .Z(n8738) );
  NAND U12928 ( .A(n8740), .B(n8741), .Z(n8695) );
  NANDN U12929 ( .A(n8742), .B(n8743), .Z(n8741) );
  NAND U12930 ( .A(n8744), .B(n8745), .Z(n8743) );
  OR U12931 ( .A(n8745), .B(n8744), .Z(n8740) );
  IV U12932 ( .A(n8746), .Z(n8744) );
  XOR U12933 ( .A(n8721), .B(n8747), .Z(N29430) );
  XNOR U12934 ( .A(n8724), .B(n8723), .Z(n8747) );
  XNOR U12935 ( .A(n8735), .B(n8748), .Z(n8723) );
  XOR U12936 ( .A(n8739), .B(n8737), .Z(n8748) );
  XOR U12937 ( .A(n8745), .B(n8749), .Z(n8737) );
  XOR U12938 ( .A(n8742), .B(n8746), .Z(n8749) );
  NAND U12939 ( .A(n8750), .B(n8751), .Z(n8746) );
  NAND U12940 ( .A(n8752), .B(n8753), .Z(n8751) );
  NAND U12941 ( .A(n8754), .B(n8755), .Z(n8750) );
  AND U12942 ( .A(n8756), .B(n8757), .Z(n8742) );
  NAND U12943 ( .A(n8758), .B(n8759), .Z(n8757) );
  NAND U12944 ( .A(n8760), .B(n8761), .Z(n8756) );
  NANDN U12945 ( .A(n8762), .B(n8763), .Z(n8745) );
  NANDN U12946 ( .A(n8764), .B(n8765), .Z(n8739) );
  XNOR U12947 ( .A(n8730), .B(n8766), .Z(n8735) );
  XOR U12948 ( .A(n8728), .B(n8732), .Z(n8766) );
  NAND U12949 ( .A(n8767), .B(n8768), .Z(n8732) );
  NAND U12950 ( .A(n8769), .B(n8770), .Z(n8768) );
  NAND U12951 ( .A(n8771), .B(n8772), .Z(n8767) );
  AND U12952 ( .A(n8773), .B(n8774), .Z(n8728) );
  NAND U12953 ( .A(n8775), .B(n8776), .Z(n8774) );
  NAND U12954 ( .A(n8777), .B(n8778), .Z(n8773) );
  AND U12955 ( .A(n8779), .B(n8780), .Z(n8730) );
  NAND U12956 ( .A(n8781), .B(n8782), .Z(n8724) );
  XNOR U12957 ( .A(n8707), .B(n8783), .Z(n8721) );
  XOR U12958 ( .A(n8711), .B(n8709), .Z(n8783) );
  XOR U12959 ( .A(n8717), .B(n8784), .Z(n8709) );
  XOR U12960 ( .A(n8714), .B(n8718), .Z(n8784) );
  NAND U12961 ( .A(n8785), .B(n8786), .Z(n8718) );
  NAND U12962 ( .A(n8787), .B(n8788), .Z(n8786) );
  NAND U12963 ( .A(n8789), .B(n8790), .Z(n8785) );
  AND U12964 ( .A(n8791), .B(n8792), .Z(n8714) );
  NAND U12965 ( .A(n8793), .B(n8794), .Z(n8792) );
  NAND U12966 ( .A(n8795), .B(n8796), .Z(n8791) );
  NANDN U12967 ( .A(n8797), .B(n8798), .Z(n8717) );
  NANDN U12968 ( .A(n8799), .B(n8800), .Z(n8711) );
  XNOR U12969 ( .A(n8702), .B(n8801), .Z(n8707) );
  XOR U12970 ( .A(n8700), .B(n8704), .Z(n8801) );
  NAND U12971 ( .A(n8802), .B(n8803), .Z(n8704) );
  NAND U12972 ( .A(n8804), .B(n8805), .Z(n8803) );
  NAND U12973 ( .A(n8806), .B(n8807), .Z(n8802) );
  AND U12974 ( .A(n8808), .B(n8809), .Z(n8700) );
  NAND U12975 ( .A(n8810), .B(n8811), .Z(n8809) );
  NAND U12976 ( .A(n8812), .B(n8813), .Z(n8808) );
  AND U12977 ( .A(n8814), .B(n8815), .Z(n8702) );
  XOR U12978 ( .A(n8782), .B(n8781), .Z(N29429) );
  XNOR U12979 ( .A(n8800), .B(n8799), .Z(n8781) );
  XNOR U12980 ( .A(n8814), .B(n8815), .Z(n8799) );
  XOR U12981 ( .A(n8811), .B(n8810), .Z(n8815) );
  XOR U12982 ( .A(y[3003]), .B(x[3003]), .Z(n8810) );
  XOR U12983 ( .A(n8813), .B(n8812), .Z(n8811) );
  XOR U12984 ( .A(y[3005]), .B(x[3005]), .Z(n8812) );
  XOR U12985 ( .A(y[3004]), .B(x[3004]), .Z(n8813) );
  XOR U12986 ( .A(n8805), .B(n8804), .Z(n8814) );
  XOR U12987 ( .A(n8807), .B(n8806), .Z(n8804) );
  XOR U12988 ( .A(y[3002]), .B(x[3002]), .Z(n8806) );
  XOR U12989 ( .A(y[3001]), .B(x[3001]), .Z(n8807) );
  XOR U12990 ( .A(y[3000]), .B(x[3000]), .Z(n8805) );
  XNOR U12991 ( .A(n8798), .B(n8797), .Z(n8800) );
  XNOR U12992 ( .A(n8794), .B(n8793), .Z(n8797) );
  XOR U12993 ( .A(n8796), .B(n8795), .Z(n8793) );
  XOR U12994 ( .A(y[2999]), .B(x[2999]), .Z(n8795) );
  XOR U12995 ( .A(y[2998]), .B(x[2998]), .Z(n8796) );
  XOR U12996 ( .A(y[2997]), .B(x[2997]), .Z(n8794) );
  XOR U12997 ( .A(n8788), .B(n8787), .Z(n8798) );
  XOR U12998 ( .A(n8790), .B(n8789), .Z(n8787) );
  XOR U12999 ( .A(y[2996]), .B(x[2996]), .Z(n8789) );
  XOR U13000 ( .A(y[2995]), .B(x[2995]), .Z(n8790) );
  XOR U13001 ( .A(y[2994]), .B(x[2994]), .Z(n8788) );
  XNOR U13002 ( .A(n8765), .B(n8764), .Z(n8782) );
  XNOR U13003 ( .A(n8779), .B(n8780), .Z(n8764) );
  XOR U13004 ( .A(n8776), .B(n8775), .Z(n8780) );
  XOR U13005 ( .A(y[2991]), .B(x[2991]), .Z(n8775) );
  XOR U13006 ( .A(n8778), .B(n8777), .Z(n8776) );
  XOR U13007 ( .A(y[2993]), .B(x[2993]), .Z(n8777) );
  XOR U13008 ( .A(y[2992]), .B(x[2992]), .Z(n8778) );
  XOR U13009 ( .A(n8770), .B(n8769), .Z(n8779) );
  XOR U13010 ( .A(n8772), .B(n8771), .Z(n8769) );
  XOR U13011 ( .A(y[2990]), .B(x[2990]), .Z(n8771) );
  XOR U13012 ( .A(y[2989]), .B(x[2989]), .Z(n8772) );
  XOR U13013 ( .A(y[2988]), .B(x[2988]), .Z(n8770) );
  XNOR U13014 ( .A(n8763), .B(n8762), .Z(n8765) );
  XNOR U13015 ( .A(n8759), .B(n8758), .Z(n8762) );
  XOR U13016 ( .A(n8761), .B(n8760), .Z(n8758) );
  XOR U13017 ( .A(y[2987]), .B(x[2987]), .Z(n8760) );
  XOR U13018 ( .A(y[2986]), .B(x[2986]), .Z(n8761) );
  XOR U13019 ( .A(y[2985]), .B(x[2985]), .Z(n8759) );
  XOR U13020 ( .A(n8753), .B(n8752), .Z(n8763) );
  XOR U13021 ( .A(n8755), .B(n8754), .Z(n8752) );
  XOR U13022 ( .A(y[2984]), .B(x[2984]), .Z(n8754) );
  XOR U13023 ( .A(y[2983]), .B(x[2983]), .Z(n8755) );
  XOR U13024 ( .A(y[2982]), .B(x[2982]), .Z(n8753) );
  NAND U13025 ( .A(n8816), .B(n8817), .Z(N29421) );
  NAND U13026 ( .A(n8818), .B(n8819), .Z(n8817) );
  NANDN U13027 ( .A(n8820), .B(n8821), .Z(n8819) );
  NANDN U13028 ( .A(n8821), .B(n8820), .Z(n8816) );
  XOR U13029 ( .A(n8820), .B(n8822), .Z(N29420) );
  XNOR U13030 ( .A(n8818), .B(n8821), .Z(n8822) );
  NAND U13031 ( .A(n8823), .B(n8824), .Z(n8821) );
  NAND U13032 ( .A(n8825), .B(n8826), .Z(n8824) );
  NANDN U13033 ( .A(n8827), .B(n8828), .Z(n8826) );
  NANDN U13034 ( .A(n8828), .B(n8827), .Z(n8823) );
  AND U13035 ( .A(n8829), .B(n8830), .Z(n8818) );
  NAND U13036 ( .A(n8831), .B(n8832), .Z(n8830) );
  OR U13037 ( .A(n8833), .B(n8834), .Z(n8832) );
  NAND U13038 ( .A(n8834), .B(n8833), .Z(n8829) );
  IV U13039 ( .A(n8835), .Z(n8834) );
  AND U13040 ( .A(n8836), .B(n8837), .Z(n8820) );
  NAND U13041 ( .A(n8838), .B(n8839), .Z(n8837) );
  NANDN U13042 ( .A(n8840), .B(n8841), .Z(n8839) );
  NANDN U13043 ( .A(n8841), .B(n8840), .Z(n8836) );
  XOR U13044 ( .A(n8833), .B(n8842), .Z(N29419) );
  XOR U13045 ( .A(n8831), .B(n8835), .Z(n8842) );
  XNOR U13046 ( .A(n8828), .B(n8843), .Z(n8835) );
  XNOR U13047 ( .A(n8825), .B(n8827), .Z(n8843) );
  AND U13048 ( .A(n8844), .B(n8845), .Z(n8827) );
  NANDN U13049 ( .A(n8846), .B(n8847), .Z(n8845) );
  NANDN U13050 ( .A(n8848), .B(n8849), .Z(n8847) );
  IV U13051 ( .A(n8850), .Z(n8849) );
  NAND U13052 ( .A(n8850), .B(n8848), .Z(n8844) );
  AND U13053 ( .A(n8851), .B(n8852), .Z(n8825) );
  NAND U13054 ( .A(n8853), .B(n8854), .Z(n8852) );
  OR U13055 ( .A(n8855), .B(n8856), .Z(n8854) );
  NAND U13056 ( .A(n8856), .B(n8855), .Z(n8851) );
  IV U13057 ( .A(n8857), .Z(n8856) );
  NAND U13058 ( .A(n8858), .B(n8859), .Z(n8828) );
  NANDN U13059 ( .A(n8860), .B(n8861), .Z(n8859) );
  NAND U13060 ( .A(n8862), .B(n8863), .Z(n8861) );
  OR U13061 ( .A(n8863), .B(n8862), .Z(n8858) );
  IV U13062 ( .A(n8864), .Z(n8862) );
  AND U13063 ( .A(n8865), .B(n8866), .Z(n8831) );
  NAND U13064 ( .A(n8867), .B(n8868), .Z(n8866) );
  NANDN U13065 ( .A(n8869), .B(n8870), .Z(n8868) );
  NANDN U13066 ( .A(n8870), .B(n8869), .Z(n8865) );
  XOR U13067 ( .A(n8841), .B(n8871), .Z(n8833) );
  XNOR U13068 ( .A(n8838), .B(n8840), .Z(n8871) );
  AND U13069 ( .A(n8872), .B(n8873), .Z(n8840) );
  NANDN U13070 ( .A(n8874), .B(n8875), .Z(n8873) );
  NANDN U13071 ( .A(n8876), .B(n8877), .Z(n8875) );
  IV U13072 ( .A(n8878), .Z(n8877) );
  NAND U13073 ( .A(n8878), .B(n8876), .Z(n8872) );
  AND U13074 ( .A(n8879), .B(n8880), .Z(n8838) );
  NAND U13075 ( .A(n8881), .B(n8882), .Z(n8880) );
  OR U13076 ( .A(n8883), .B(n8884), .Z(n8882) );
  NAND U13077 ( .A(n8884), .B(n8883), .Z(n8879) );
  IV U13078 ( .A(n8885), .Z(n8884) );
  NAND U13079 ( .A(n8886), .B(n8887), .Z(n8841) );
  NANDN U13080 ( .A(n8888), .B(n8889), .Z(n8887) );
  NAND U13081 ( .A(n8890), .B(n8891), .Z(n8889) );
  OR U13082 ( .A(n8891), .B(n8890), .Z(n8886) );
  IV U13083 ( .A(n8892), .Z(n8890) );
  XOR U13084 ( .A(n8867), .B(n8893), .Z(N29418) );
  XNOR U13085 ( .A(n8870), .B(n8869), .Z(n8893) );
  XNOR U13086 ( .A(n8881), .B(n8894), .Z(n8869) );
  XOR U13087 ( .A(n8885), .B(n8883), .Z(n8894) );
  XOR U13088 ( .A(n8891), .B(n8895), .Z(n8883) );
  XOR U13089 ( .A(n8888), .B(n8892), .Z(n8895) );
  NAND U13090 ( .A(n8896), .B(n8897), .Z(n8892) );
  NAND U13091 ( .A(n8898), .B(n8899), .Z(n8897) );
  NAND U13092 ( .A(n8900), .B(n8901), .Z(n8896) );
  AND U13093 ( .A(n8902), .B(n8903), .Z(n8888) );
  NAND U13094 ( .A(n8904), .B(n8905), .Z(n8903) );
  NAND U13095 ( .A(n8906), .B(n8907), .Z(n8902) );
  NANDN U13096 ( .A(n8908), .B(n8909), .Z(n8891) );
  NANDN U13097 ( .A(n8910), .B(n8911), .Z(n8885) );
  XNOR U13098 ( .A(n8876), .B(n8912), .Z(n8881) );
  XOR U13099 ( .A(n8874), .B(n8878), .Z(n8912) );
  NAND U13100 ( .A(n8913), .B(n8914), .Z(n8878) );
  NAND U13101 ( .A(n8915), .B(n8916), .Z(n8914) );
  NAND U13102 ( .A(n8917), .B(n8918), .Z(n8913) );
  AND U13103 ( .A(n8919), .B(n8920), .Z(n8874) );
  NAND U13104 ( .A(n8921), .B(n8922), .Z(n8920) );
  NAND U13105 ( .A(n8923), .B(n8924), .Z(n8919) );
  AND U13106 ( .A(n8925), .B(n8926), .Z(n8876) );
  NAND U13107 ( .A(n8927), .B(n8928), .Z(n8870) );
  XNOR U13108 ( .A(n8853), .B(n8929), .Z(n8867) );
  XOR U13109 ( .A(n8857), .B(n8855), .Z(n8929) );
  XOR U13110 ( .A(n8863), .B(n8930), .Z(n8855) );
  XOR U13111 ( .A(n8860), .B(n8864), .Z(n8930) );
  NAND U13112 ( .A(n8931), .B(n8932), .Z(n8864) );
  NAND U13113 ( .A(n8933), .B(n8934), .Z(n8932) );
  NAND U13114 ( .A(n8935), .B(n8936), .Z(n8931) );
  AND U13115 ( .A(n8937), .B(n8938), .Z(n8860) );
  NAND U13116 ( .A(n8939), .B(n8940), .Z(n8938) );
  NAND U13117 ( .A(n8941), .B(n8942), .Z(n8937) );
  NANDN U13118 ( .A(n8943), .B(n8944), .Z(n8863) );
  NANDN U13119 ( .A(n8945), .B(n8946), .Z(n8857) );
  XNOR U13120 ( .A(n8848), .B(n8947), .Z(n8853) );
  XOR U13121 ( .A(n8846), .B(n8850), .Z(n8947) );
  NAND U13122 ( .A(n8948), .B(n8949), .Z(n8850) );
  NAND U13123 ( .A(n8950), .B(n8951), .Z(n8949) );
  NAND U13124 ( .A(n8952), .B(n8953), .Z(n8948) );
  AND U13125 ( .A(n8954), .B(n8955), .Z(n8846) );
  NAND U13126 ( .A(n8956), .B(n8957), .Z(n8955) );
  NAND U13127 ( .A(n8958), .B(n8959), .Z(n8954) );
  AND U13128 ( .A(n8960), .B(n8961), .Z(n8848) );
  XOR U13129 ( .A(n8928), .B(n8927), .Z(N29417) );
  XNOR U13130 ( .A(n8946), .B(n8945), .Z(n8927) );
  XNOR U13131 ( .A(n8960), .B(n8961), .Z(n8945) );
  XOR U13132 ( .A(n8957), .B(n8956), .Z(n8961) );
  XOR U13133 ( .A(y[2979]), .B(x[2979]), .Z(n8956) );
  XOR U13134 ( .A(n8959), .B(n8958), .Z(n8957) );
  XOR U13135 ( .A(y[2981]), .B(x[2981]), .Z(n8958) );
  XOR U13136 ( .A(y[2980]), .B(x[2980]), .Z(n8959) );
  XOR U13137 ( .A(n8951), .B(n8950), .Z(n8960) );
  XOR U13138 ( .A(n8953), .B(n8952), .Z(n8950) );
  XOR U13139 ( .A(y[2978]), .B(x[2978]), .Z(n8952) );
  XOR U13140 ( .A(y[2977]), .B(x[2977]), .Z(n8953) );
  XOR U13141 ( .A(y[2976]), .B(x[2976]), .Z(n8951) );
  XNOR U13142 ( .A(n8944), .B(n8943), .Z(n8946) );
  XNOR U13143 ( .A(n8940), .B(n8939), .Z(n8943) );
  XOR U13144 ( .A(n8942), .B(n8941), .Z(n8939) );
  XOR U13145 ( .A(y[2975]), .B(x[2975]), .Z(n8941) );
  XOR U13146 ( .A(y[2974]), .B(x[2974]), .Z(n8942) );
  XOR U13147 ( .A(y[2973]), .B(x[2973]), .Z(n8940) );
  XOR U13148 ( .A(n8934), .B(n8933), .Z(n8944) );
  XOR U13149 ( .A(n8936), .B(n8935), .Z(n8933) );
  XOR U13150 ( .A(y[2972]), .B(x[2972]), .Z(n8935) );
  XOR U13151 ( .A(y[2971]), .B(x[2971]), .Z(n8936) );
  XOR U13152 ( .A(y[2970]), .B(x[2970]), .Z(n8934) );
  XNOR U13153 ( .A(n8911), .B(n8910), .Z(n8928) );
  XNOR U13154 ( .A(n8925), .B(n8926), .Z(n8910) );
  XOR U13155 ( .A(n8922), .B(n8921), .Z(n8926) );
  XOR U13156 ( .A(y[2967]), .B(x[2967]), .Z(n8921) );
  XOR U13157 ( .A(n8924), .B(n8923), .Z(n8922) );
  XOR U13158 ( .A(y[2969]), .B(x[2969]), .Z(n8923) );
  XOR U13159 ( .A(y[2968]), .B(x[2968]), .Z(n8924) );
  XOR U13160 ( .A(n8916), .B(n8915), .Z(n8925) );
  XOR U13161 ( .A(n8918), .B(n8917), .Z(n8915) );
  XOR U13162 ( .A(y[2966]), .B(x[2966]), .Z(n8917) );
  XOR U13163 ( .A(y[2965]), .B(x[2965]), .Z(n8918) );
  XOR U13164 ( .A(y[2964]), .B(x[2964]), .Z(n8916) );
  XNOR U13165 ( .A(n8909), .B(n8908), .Z(n8911) );
  XNOR U13166 ( .A(n8905), .B(n8904), .Z(n8908) );
  XOR U13167 ( .A(n8907), .B(n8906), .Z(n8904) );
  XOR U13168 ( .A(y[2963]), .B(x[2963]), .Z(n8906) );
  XOR U13169 ( .A(y[2962]), .B(x[2962]), .Z(n8907) );
  XOR U13170 ( .A(y[2961]), .B(x[2961]), .Z(n8905) );
  XOR U13171 ( .A(n8899), .B(n8898), .Z(n8909) );
  XOR U13172 ( .A(n8901), .B(n8900), .Z(n8898) );
  XOR U13173 ( .A(y[2960]), .B(x[2960]), .Z(n8900) );
  XOR U13174 ( .A(y[2959]), .B(x[2959]), .Z(n8901) );
  XOR U13175 ( .A(y[2958]), .B(x[2958]), .Z(n8899) );
  NAND U13176 ( .A(n8962), .B(n8963), .Z(N29409) );
  NAND U13177 ( .A(n8964), .B(n8965), .Z(n8963) );
  NANDN U13178 ( .A(n8966), .B(n8967), .Z(n8965) );
  NANDN U13179 ( .A(n8967), .B(n8966), .Z(n8962) );
  XOR U13180 ( .A(n8966), .B(n8968), .Z(N29408) );
  XNOR U13181 ( .A(n8964), .B(n8967), .Z(n8968) );
  NAND U13182 ( .A(n8969), .B(n8970), .Z(n8967) );
  NAND U13183 ( .A(n8971), .B(n8972), .Z(n8970) );
  NANDN U13184 ( .A(n8973), .B(n8974), .Z(n8972) );
  NANDN U13185 ( .A(n8974), .B(n8973), .Z(n8969) );
  AND U13186 ( .A(n8975), .B(n8976), .Z(n8964) );
  NAND U13187 ( .A(n8977), .B(n8978), .Z(n8976) );
  OR U13188 ( .A(n8979), .B(n8980), .Z(n8978) );
  NAND U13189 ( .A(n8980), .B(n8979), .Z(n8975) );
  IV U13190 ( .A(n8981), .Z(n8980) );
  AND U13191 ( .A(n8982), .B(n8983), .Z(n8966) );
  NAND U13192 ( .A(n8984), .B(n8985), .Z(n8983) );
  NANDN U13193 ( .A(n8986), .B(n8987), .Z(n8985) );
  NANDN U13194 ( .A(n8987), .B(n8986), .Z(n8982) );
  XOR U13195 ( .A(n8979), .B(n8988), .Z(N29407) );
  XOR U13196 ( .A(n8977), .B(n8981), .Z(n8988) );
  XNOR U13197 ( .A(n8974), .B(n8989), .Z(n8981) );
  XNOR U13198 ( .A(n8971), .B(n8973), .Z(n8989) );
  AND U13199 ( .A(n8990), .B(n8991), .Z(n8973) );
  NANDN U13200 ( .A(n8992), .B(n8993), .Z(n8991) );
  NANDN U13201 ( .A(n8994), .B(n8995), .Z(n8993) );
  IV U13202 ( .A(n8996), .Z(n8995) );
  NAND U13203 ( .A(n8996), .B(n8994), .Z(n8990) );
  AND U13204 ( .A(n8997), .B(n8998), .Z(n8971) );
  NAND U13205 ( .A(n8999), .B(n9000), .Z(n8998) );
  OR U13206 ( .A(n9001), .B(n9002), .Z(n9000) );
  NAND U13207 ( .A(n9002), .B(n9001), .Z(n8997) );
  IV U13208 ( .A(n9003), .Z(n9002) );
  NAND U13209 ( .A(n9004), .B(n9005), .Z(n8974) );
  NANDN U13210 ( .A(n9006), .B(n9007), .Z(n9005) );
  NAND U13211 ( .A(n9008), .B(n9009), .Z(n9007) );
  OR U13212 ( .A(n9009), .B(n9008), .Z(n9004) );
  IV U13213 ( .A(n9010), .Z(n9008) );
  AND U13214 ( .A(n9011), .B(n9012), .Z(n8977) );
  NAND U13215 ( .A(n9013), .B(n9014), .Z(n9012) );
  NANDN U13216 ( .A(n9015), .B(n9016), .Z(n9014) );
  NANDN U13217 ( .A(n9016), .B(n9015), .Z(n9011) );
  XOR U13218 ( .A(n8987), .B(n9017), .Z(n8979) );
  XNOR U13219 ( .A(n8984), .B(n8986), .Z(n9017) );
  AND U13220 ( .A(n9018), .B(n9019), .Z(n8986) );
  NANDN U13221 ( .A(n9020), .B(n9021), .Z(n9019) );
  NANDN U13222 ( .A(n9022), .B(n9023), .Z(n9021) );
  IV U13223 ( .A(n9024), .Z(n9023) );
  NAND U13224 ( .A(n9024), .B(n9022), .Z(n9018) );
  AND U13225 ( .A(n9025), .B(n9026), .Z(n8984) );
  NAND U13226 ( .A(n9027), .B(n9028), .Z(n9026) );
  OR U13227 ( .A(n9029), .B(n9030), .Z(n9028) );
  NAND U13228 ( .A(n9030), .B(n9029), .Z(n9025) );
  IV U13229 ( .A(n9031), .Z(n9030) );
  NAND U13230 ( .A(n9032), .B(n9033), .Z(n8987) );
  NANDN U13231 ( .A(n9034), .B(n9035), .Z(n9033) );
  NAND U13232 ( .A(n9036), .B(n9037), .Z(n9035) );
  OR U13233 ( .A(n9037), .B(n9036), .Z(n9032) );
  IV U13234 ( .A(n9038), .Z(n9036) );
  XOR U13235 ( .A(n9013), .B(n9039), .Z(N29406) );
  XNOR U13236 ( .A(n9016), .B(n9015), .Z(n9039) );
  XNOR U13237 ( .A(n9027), .B(n9040), .Z(n9015) );
  XOR U13238 ( .A(n9031), .B(n9029), .Z(n9040) );
  XOR U13239 ( .A(n9037), .B(n9041), .Z(n9029) );
  XOR U13240 ( .A(n9034), .B(n9038), .Z(n9041) );
  NAND U13241 ( .A(n9042), .B(n9043), .Z(n9038) );
  NAND U13242 ( .A(n9044), .B(n9045), .Z(n9043) );
  NAND U13243 ( .A(n9046), .B(n9047), .Z(n9042) );
  AND U13244 ( .A(n9048), .B(n9049), .Z(n9034) );
  NAND U13245 ( .A(n9050), .B(n9051), .Z(n9049) );
  NAND U13246 ( .A(n9052), .B(n9053), .Z(n9048) );
  NANDN U13247 ( .A(n9054), .B(n9055), .Z(n9037) );
  NANDN U13248 ( .A(n9056), .B(n9057), .Z(n9031) );
  XNOR U13249 ( .A(n9022), .B(n9058), .Z(n9027) );
  XOR U13250 ( .A(n9020), .B(n9024), .Z(n9058) );
  NAND U13251 ( .A(n9059), .B(n9060), .Z(n9024) );
  NAND U13252 ( .A(n9061), .B(n9062), .Z(n9060) );
  NAND U13253 ( .A(n9063), .B(n9064), .Z(n9059) );
  AND U13254 ( .A(n9065), .B(n9066), .Z(n9020) );
  NAND U13255 ( .A(n9067), .B(n9068), .Z(n9066) );
  NAND U13256 ( .A(n9069), .B(n9070), .Z(n9065) );
  AND U13257 ( .A(n9071), .B(n9072), .Z(n9022) );
  NAND U13258 ( .A(n9073), .B(n9074), .Z(n9016) );
  XNOR U13259 ( .A(n8999), .B(n9075), .Z(n9013) );
  XOR U13260 ( .A(n9003), .B(n9001), .Z(n9075) );
  XOR U13261 ( .A(n9009), .B(n9076), .Z(n9001) );
  XOR U13262 ( .A(n9006), .B(n9010), .Z(n9076) );
  NAND U13263 ( .A(n9077), .B(n9078), .Z(n9010) );
  NAND U13264 ( .A(n9079), .B(n9080), .Z(n9078) );
  NAND U13265 ( .A(n9081), .B(n9082), .Z(n9077) );
  AND U13266 ( .A(n9083), .B(n9084), .Z(n9006) );
  NAND U13267 ( .A(n9085), .B(n9086), .Z(n9084) );
  NAND U13268 ( .A(n9087), .B(n9088), .Z(n9083) );
  NANDN U13269 ( .A(n9089), .B(n9090), .Z(n9009) );
  NANDN U13270 ( .A(n9091), .B(n9092), .Z(n9003) );
  XNOR U13271 ( .A(n8994), .B(n9093), .Z(n8999) );
  XOR U13272 ( .A(n8992), .B(n8996), .Z(n9093) );
  NAND U13273 ( .A(n9094), .B(n9095), .Z(n8996) );
  NAND U13274 ( .A(n9096), .B(n9097), .Z(n9095) );
  NAND U13275 ( .A(n9098), .B(n9099), .Z(n9094) );
  AND U13276 ( .A(n9100), .B(n9101), .Z(n8992) );
  NAND U13277 ( .A(n9102), .B(n9103), .Z(n9101) );
  NAND U13278 ( .A(n9104), .B(n9105), .Z(n9100) );
  AND U13279 ( .A(n9106), .B(n9107), .Z(n8994) );
  XOR U13280 ( .A(n9074), .B(n9073), .Z(N29405) );
  XNOR U13281 ( .A(n9092), .B(n9091), .Z(n9073) );
  XNOR U13282 ( .A(n9106), .B(n9107), .Z(n9091) );
  XOR U13283 ( .A(n9103), .B(n9102), .Z(n9107) );
  XOR U13284 ( .A(y[2955]), .B(x[2955]), .Z(n9102) );
  XOR U13285 ( .A(n9105), .B(n9104), .Z(n9103) );
  XOR U13286 ( .A(y[2957]), .B(x[2957]), .Z(n9104) );
  XOR U13287 ( .A(y[2956]), .B(x[2956]), .Z(n9105) );
  XOR U13288 ( .A(n9097), .B(n9096), .Z(n9106) );
  XOR U13289 ( .A(n9099), .B(n9098), .Z(n9096) );
  XOR U13290 ( .A(y[2954]), .B(x[2954]), .Z(n9098) );
  XOR U13291 ( .A(y[2953]), .B(x[2953]), .Z(n9099) );
  XOR U13292 ( .A(y[2952]), .B(x[2952]), .Z(n9097) );
  XNOR U13293 ( .A(n9090), .B(n9089), .Z(n9092) );
  XNOR U13294 ( .A(n9086), .B(n9085), .Z(n9089) );
  XOR U13295 ( .A(n9088), .B(n9087), .Z(n9085) );
  XOR U13296 ( .A(y[2951]), .B(x[2951]), .Z(n9087) );
  XOR U13297 ( .A(y[2950]), .B(x[2950]), .Z(n9088) );
  XOR U13298 ( .A(y[2949]), .B(x[2949]), .Z(n9086) );
  XOR U13299 ( .A(n9080), .B(n9079), .Z(n9090) );
  XOR U13300 ( .A(n9082), .B(n9081), .Z(n9079) );
  XOR U13301 ( .A(y[2948]), .B(x[2948]), .Z(n9081) );
  XOR U13302 ( .A(y[2947]), .B(x[2947]), .Z(n9082) );
  XOR U13303 ( .A(y[2946]), .B(x[2946]), .Z(n9080) );
  XNOR U13304 ( .A(n9057), .B(n9056), .Z(n9074) );
  XNOR U13305 ( .A(n9071), .B(n9072), .Z(n9056) );
  XOR U13306 ( .A(n9068), .B(n9067), .Z(n9072) );
  XOR U13307 ( .A(y[2943]), .B(x[2943]), .Z(n9067) );
  XOR U13308 ( .A(n9070), .B(n9069), .Z(n9068) );
  XOR U13309 ( .A(y[2945]), .B(x[2945]), .Z(n9069) );
  XOR U13310 ( .A(y[2944]), .B(x[2944]), .Z(n9070) );
  XOR U13311 ( .A(n9062), .B(n9061), .Z(n9071) );
  XOR U13312 ( .A(n9064), .B(n9063), .Z(n9061) );
  XOR U13313 ( .A(y[2942]), .B(x[2942]), .Z(n9063) );
  XOR U13314 ( .A(y[2941]), .B(x[2941]), .Z(n9064) );
  XOR U13315 ( .A(y[2940]), .B(x[2940]), .Z(n9062) );
  XNOR U13316 ( .A(n9055), .B(n9054), .Z(n9057) );
  XNOR U13317 ( .A(n9051), .B(n9050), .Z(n9054) );
  XOR U13318 ( .A(n9053), .B(n9052), .Z(n9050) );
  XOR U13319 ( .A(y[2939]), .B(x[2939]), .Z(n9052) );
  XOR U13320 ( .A(y[2938]), .B(x[2938]), .Z(n9053) );
  XOR U13321 ( .A(y[2937]), .B(x[2937]), .Z(n9051) );
  XOR U13322 ( .A(n9045), .B(n9044), .Z(n9055) );
  XOR U13323 ( .A(n9047), .B(n9046), .Z(n9044) );
  XOR U13324 ( .A(y[2936]), .B(x[2936]), .Z(n9046) );
  XOR U13325 ( .A(y[2935]), .B(x[2935]), .Z(n9047) );
  XOR U13326 ( .A(y[2934]), .B(x[2934]), .Z(n9045) );
  NAND U13327 ( .A(n9108), .B(n9109), .Z(N29397) );
  NAND U13328 ( .A(n9110), .B(n9111), .Z(n9109) );
  NANDN U13329 ( .A(n9112), .B(n9113), .Z(n9111) );
  NANDN U13330 ( .A(n9113), .B(n9112), .Z(n9108) );
  XOR U13331 ( .A(n9112), .B(n9114), .Z(N29396) );
  XNOR U13332 ( .A(n9110), .B(n9113), .Z(n9114) );
  NAND U13333 ( .A(n9115), .B(n9116), .Z(n9113) );
  NAND U13334 ( .A(n9117), .B(n9118), .Z(n9116) );
  NANDN U13335 ( .A(n9119), .B(n9120), .Z(n9118) );
  NANDN U13336 ( .A(n9120), .B(n9119), .Z(n9115) );
  AND U13337 ( .A(n9121), .B(n9122), .Z(n9110) );
  NAND U13338 ( .A(n9123), .B(n9124), .Z(n9122) );
  OR U13339 ( .A(n9125), .B(n9126), .Z(n9124) );
  NAND U13340 ( .A(n9126), .B(n9125), .Z(n9121) );
  IV U13341 ( .A(n9127), .Z(n9126) );
  AND U13342 ( .A(n9128), .B(n9129), .Z(n9112) );
  NAND U13343 ( .A(n9130), .B(n9131), .Z(n9129) );
  NANDN U13344 ( .A(n9132), .B(n9133), .Z(n9131) );
  NANDN U13345 ( .A(n9133), .B(n9132), .Z(n9128) );
  XOR U13346 ( .A(n9125), .B(n9134), .Z(N29395) );
  XOR U13347 ( .A(n9123), .B(n9127), .Z(n9134) );
  XNOR U13348 ( .A(n9120), .B(n9135), .Z(n9127) );
  XNOR U13349 ( .A(n9117), .B(n9119), .Z(n9135) );
  AND U13350 ( .A(n9136), .B(n9137), .Z(n9119) );
  NANDN U13351 ( .A(n9138), .B(n9139), .Z(n9137) );
  NANDN U13352 ( .A(n9140), .B(n9141), .Z(n9139) );
  IV U13353 ( .A(n9142), .Z(n9141) );
  NAND U13354 ( .A(n9142), .B(n9140), .Z(n9136) );
  AND U13355 ( .A(n9143), .B(n9144), .Z(n9117) );
  NAND U13356 ( .A(n9145), .B(n9146), .Z(n9144) );
  OR U13357 ( .A(n9147), .B(n9148), .Z(n9146) );
  NAND U13358 ( .A(n9148), .B(n9147), .Z(n9143) );
  IV U13359 ( .A(n9149), .Z(n9148) );
  NAND U13360 ( .A(n9150), .B(n9151), .Z(n9120) );
  NANDN U13361 ( .A(n9152), .B(n9153), .Z(n9151) );
  NAND U13362 ( .A(n9154), .B(n9155), .Z(n9153) );
  OR U13363 ( .A(n9155), .B(n9154), .Z(n9150) );
  IV U13364 ( .A(n9156), .Z(n9154) );
  AND U13365 ( .A(n9157), .B(n9158), .Z(n9123) );
  NAND U13366 ( .A(n9159), .B(n9160), .Z(n9158) );
  NANDN U13367 ( .A(n9161), .B(n9162), .Z(n9160) );
  NANDN U13368 ( .A(n9162), .B(n9161), .Z(n9157) );
  XOR U13369 ( .A(n9133), .B(n9163), .Z(n9125) );
  XNOR U13370 ( .A(n9130), .B(n9132), .Z(n9163) );
  AND U13371 ( .A(n9164), .B(n9165), .Z(n9132) );
  NANDN U13372 ( .A(n9166), .B(n9167), .Z(n9165) );
  NANDN U13373 ( .A(n9168), .B(n9169), .Z(n9167) );
  IV U13374 ( .A(n9170), .Z(n9169) );
  NAND U13375 ( .A(n9170), .B(n9168), .Z(n9164) );
  AND U13376 ( .A(n9171), .B(n9172), .Z(n9130) );
  NAND U13377 ( .A(n9173), .B(n9174), .Z(n9172) );
  OR U13378 ( .A(n9175), .B(n9176), .Z(n9174) );
  NAND U13379 ( .A(n9176), .B(n9175), .Z(n9171) );
  IV U13380 ( .A(n9177), .Z(n9176) );
  NAND U13381 ( .A(n9178), .B(n9179), .Z(n9133) );
  NANDN U13382 ( .A(n9180), .B(n9181), .Z(n9179) );
  NAND U13383 ( .A(n9182), .B(n9183), .Z(n9181) );
  OR U13384 ( .A(n9183), .B(n9182), .Z(n9178) );
  IV U13385 ( .A(n9184), .Z(n9182) );
  XOR U13386 ( .A(n9159), .B(n9185), .Z(N29394) );
  XNOR U13387 ( .A(n9162), .B(n9161), .Z(n9185) );
  XNOR U13388 ( .A(n9173), .B(n9186), .Z(n9161) );
  XOR U13389 ( .A(n9177), .B(n9175), .Z(n9186) );
  XOR U13390 ( .A(n9183), .B(n9187), .Z(n9175) );
  XOR U13391 ( .A(n9180), .B(n9184), .Z(n9187) );
  NAND U13392 ( .A(n9188), .B(n9189), .Z(n9184) );
  NAND U13393 ( .A(n9190), .B(n9191), .Z(n9189) );
  NAND U13394 ( .A(n9192), .B(n9193), .Z(n9188) );
  AND U13395 ( .A(n9194), .B(n9195), .Z(n9180) );
  NAND U13396 ( .A(n9196), .B(n9197), .Z(n9195) );
  NAND U13397 ( .A(n9198), .B(n9199), .Z(n9194) );
  NANDN U13398 ( .A(n9200), .B(n9201), .Z(n9183) );
  NANDN U13399 ( .A(n9202), .B(n9203), .Z(n9177) );
  XNOR U13400 ( .A(n9168), .B(n9204), .Z(n9173) );
  XOR U13401 ( .A(n9166), .B(n9170), .Z(n9204) );
  NAND U13402 ( .A(n9205), .B(n9206), .Z(n9170) );
  NAND U13403 ( .A(n9207), .B(n9208), .Z(n9206) );
  NAND U13404 ( .A(n9209), .B(n9210), .Z(n9205) );
  AND U13405 ( .A(n9211), .B(n9212), .Z(n9166) );
  NAND U13406 ( .A(n9213), .B(n9214), .Z(n9212) );
  NAND U13407 ( .A(n9215), .B(n9216), .Z(n9211) );
  AND U13408 ( .A(n9217), .B(n9218), .Z(n9168) );
  NAND U13409 ( .A(n9219), .B(n9220), .Z(n9162) );
  XNOR U13410 ( .A(n9145), .B(n9221), .Z(n9159) );
  XOR U13411 ( .A(n9149), .B(n9147), .Z(n9221) );
  XOR U13412 ( .A(n9155), .B(n9222), .Z(n9147) );
  XOR U13413 ( .A(n9152), .B(n9156), .Z(n9222) );
  NAND U13414 ( .A(n9223), .B(n9224), .Z(n9156) );
  NAND U13415 ( .A(n9225), .B(n9226), .Z(n9224) );
  NAND U13416 ( .A(n9227), .B(n9228), .Z(n9223) );
  AND U13417 ( .A(n9229), .B(n9230), .Z(n9152) );
  NAND U13418 ( .A(n9231), .B(n9232), .Z(n9230) );
  NAND U13419 ( .A(n9233), .B(n9234), .Z(n9229) );
  NANDN U13420 ( .A(n9235), .B(n9236), .Z(n9155) );
  NANDN U13421 ( .A(n9237), .B(n9238), .Z(n9149) );
  XNOR U13422 ( .A(n9140), .B(n9239), .Z(n9145) );
  XOR U13423 ( .A(n9138), .B(n9142), .Z(n9239) );
  NAND U13424 ( .A(n9240), .B(n9241), .Z(n9142) );
  NAND U13425 ( .A(n9242), .B(n9243), .Z(n9241) );
  NAND U13426 ( .A(n9244), .B(n9245), .Z(n9240) );
  AND U13427 ( .A(n9246), .B(n9247), .Z(n9138) );
  NAND U13428 ( .A(n9248), .B(n9249), .Z(n9247) );
  NAND U13429 ( .A(n9250), .B(n9251), .Z(n9246) );
  AND U13430 ( .A(n9252), .B(n9253), .Z(n9140) );
  XOR U13431 ( .A(n9220), .B(n9219), .Z(N29393) );
  XNOR U13432 ( .A(n9238), .B(n9237), .Z(n9219) );
  XNOR U13433 ( .A(n9252), .B(n9253), .Z(n9237) );
  XOR U13434 ( .A(n9249), .B(n9248), .Z(n9253) );
  XOR U13435 ( .A(y[2931]), .B(x[2931]), .Z(n9248) );
  XOR U13436 ( .A(n9251), .B(n9250), .Z(n9249) );
  XOR U13437 ( .A(y[2933]), .B(x[2933]), .Z(n9250) );
  XOR U13438 ( .A(y[2932]), .B(x[2932]), .Z(n9251) );
  XOR U13439 ( .A(n9243), .B(n9242), .Z(n9252) );
  XOR U13440 ( .A(n9245), .B(n9244), .Z(n9242) );
  XOR U13441 ( .A(y[2930]), .B(x[2930]), .Z(n9244) );
  XOR U13442 ( .A(y[2929]), .B(x[2929]), .Z(n9245) );
  XOR U13443 ( .A(y[2928]), .B(x[2928]), .Z(n9243) );
  XNOR U13444 ( .A(n9236), .B(n9235), .Z(n9238) );
  XNOR U13445 ( .A(n9232), .B(n9231), .Z(n9235) );
  XOR U13446 ( .A(n9234), .B(n9233), .Z(n9231) );
  XOR U13447 ( .A(y[2927]), .B(x[2927]), .Z(n9233) );
  XOR U13448 ( .A(y[2926]), .B(x[2926]), .Z(n9234) );
  XOR U13449 ( .A(y[2925]), .B(x[2925]), .Z(n9232) );
  XOR U13450 ( .A(n9226), .B(n9225), .Z(n9236) );
  XOR U13451 ( .A(n9228), .B(n9227), .Z(n9225) );
  XOR U13452 ( .A(y[2924]), .B(x[2924]), .Z(n9227) );
  XOR U13453 ( .A(y[2923]), .B(x[2923]), .Z(n9228) );
  XOR U13454 ( .A(y[2922]), .B(x[2922]), .Z(n9226) );
  XNOR U13455 ( .A(n9203), .B(n9202), .Z(n9220) );
  XNOR U13456 ( .A(n9217), .B(n9218), .Z(n9202) );
  XOR U13457 ( .A(n9214), .B(n9213), .Z(n9218) );
  XOR U13458 ( .A(y[2919]), .B(x[2919]), .Z(n9213) );
  XOR U13459 ( .A(n9216), .B(n9215), .Z(n9214) );
  XOR U13460 ( .A(y[2921]), .B(x[2921]), .Z(n9215) );
  XOR U13461 ( .A(y[2920]), .B(x[2920]), .Z(n9216) );
  XOR U13462 ( .A(n9208), .B(n9207), .Z(n9217) );
  XOR U13463 ( .A(n9210), .B(n9209), .Z(n9207) );
  XOR U13464 ( .A(y[2918]), .B(x[2918]), .Z(n9209) );
  XOR U13465 ( .A(y[2917]), .B(x[2917]), .Z(n9210) );
  XOR U13466 ( .A(y[2916]), .B(x[2916]), .Z(n9208) );
  XNOR U13467 ( .A(n9201), .B(n9200), .Z(n9203) );
  XNOR U13468 ( .A(n9197), .B(n9196), .Z(n9200) );
  XOR U13469 ( .A(n9199), .B(n9198), .Z(n9196) );
  XOR U13470 ( .A(y[2915]), .B(x[2915]), .Z(n9198) );
  XOR U13471 ( .A(y[2914]), .B(x[2914]), .Z(n9199) );
  XOR U13472 ( .A(y[2913]), .B(x[2913]), .Z(n9197) );
  XOR U13473 ( .A(n9191), .B(n9190), .Z(n9201) );
  XOR U13474 ( .A(n9193), .B(n9192), .Z(n9190) );
  XOR U13475 ( .A(y[2912]), .B(x[2912]), .Z(n9192) );
  XOR U13476 ( .A(y[2911]), .B(x[2911]), .Z(n9193) );
  XOR U13477 ( .A(y[2910]), .B(x[2910]), .Z(n9191) );
  NAND U13478 ( .A(n9254), .B(n9255), .Z(N29385) );
  NAND U13479 ( .A(n9256), .B(n9257), .Z(n9255) );
  NANDN U13480 ( .A(n9258), .B(n9259), .Z(n9257) );
  NANDN U13481 ( .A(n9259), .B(n9258), .Z(n9254) );
  XOR U13482 ( .A(n9258), .B(n9260), .Z(N29384) );
  XNOR U13483 ( .A(n9256), .B(n9259), .Z(n9260) );
  NAND U13484 ( .A(n9261), .B(n9262), .Z(n9259) );
  NAND U13485 ( .A(n9263), .B(n9264), .Z(n9262) );
  NANDN U13486 ( .A(n9265), .B(n9266), .Z(n9264) );
  NANDN U13487 ( .A(n9266), .B(n9265), .Z(n9261) );
  AND U13488 ( .A(n9267), .B(n9268), .Z(n9256) );
  NAND U13489 ( .A(n9269), .B(n9270), .Z(n9268) );
  OR U13490 ( .A(n9271), .B(n9272), .Z(n9270) );
  NAND U13491 ( .A(n9272), .B(n9271), .Z(n9267) );
  IV U13492 ( .A(n9273), .Z(n9272) );
  AND U13493 ( .A(n9274), .B(n9275), .Z(n9258) );
  NAND U13494 ( .A(n9276), .B(n9277), .Z(n9275) );
  NANDN U13495 ( .A(n9278), .B(n9279), .Z(n9277) );
  NANDN U13496 ( .A(n9279), .B(n9278), .Z(n9274) );
  XOR U13497 ( .A(n9271), .B(n9280), .Z(N29383) );
  XOR U13498 ( .A(n9269), .B(n9273), .Z(n9280) );
  XNOR U13499 ( .A(n9266), .B(n9281), .Z(n9273) );
  XNOR U13500 ( .A(n9263), .B(n9265), .Z(n9281) );
  AND U13501 ( .A(n9282), .B(n9283), .Z(n9265) );
  NANDN U13502 ( .A(n9284), .B(n9285), .Z(n9283) );
  NANDN U13503 ( .A(n9286), .B(n9287), .Z(n9285) );
  IV U13504 ( .A(n9288), .Z(n9287) );
  NAND U13505 ( .A(n9288), .B(n9286), .Z(n9282) );
  AND U13506 ( .A(n9289), .B(n9290), .Z(n9263) );
  NAND U13507 ( .A(n9291), .B(n9292), .Z(n9290) );
  OR U13508 ( .A(n9293), .B(n9294), .Z(n9292) );
  NAND U13509 ( .A(n9294), .B(n9293), .Z(n9289) );
  IV U13510 ( .A(n9295), .Z(n9294) );
  NAND U13511 ( .A(n9296), .B(n9297), .Z(n9266) );
  NANDN U13512 ( .A(n9298), .B(n9299), .Z(n9297) );
  NAND U13513 ( .A(n9300), .B(n9301), .Z(n9299) );
  OR U13514 ( .A(n9301), .B(n9300), .Z(n9296) );
  IV U13515 ( .A(n9302), .Z(n9300) );
  AND U13516 ( .A(n9303), .B(n9304), .Z(n9269) );
  NAND U13517 ( .A(n9305), .B(n9306), .Z(n9304) );
  NANDN U13518 ( .A(n9307), .B(n9308), .Z(n9306) );
  NANDN U13519 ( .A(n9308), .B(n9307), .Z(n9303) );
  XOR U13520 ( .A(n9279), .B(n9309), .Z(n9271) );
  XNOR U13521 ( .A(n9276), .B(n9278), .Z(n9309) );
  AND U13522 ( .A(n9310), .B(n9311), .Z(n9278) );
  NANDN U13523 ( .A(n9312), .B(n9313), .Z(n9311) );
  NANDN U13524 ( .A(n9314), .B(n9315), .Z(n9313) );
  IV U13525 ( .A(n9316), .Z(n9315) );
  NAND U13526 ( .A(n9316), .B(n9314), .Z(n9310) );
  AND U13527 ( .A(n9317), .B(n9318), .Z(n9276) );
  NAND U13528 ( .A(n9319), .B(n9320), .Z(n9318) );
  OR U13529 ( .A(n9321), .B(n9322), .Z(n9320) );
  NAND U13530 ( .A(n9322), .B(n9321), .Z(n9317) );
  IV U13531 ( .A(n9323), .Z(n9322) );
  NAND U13532 ( .A(n9324), .B(n9325), .Z(n9279) );
  NANDN U13533 ( .A(n9326), .B(n9327), .Z(n9325) );
  NAND U13534 ( .A(n9328), .B(n9329), .Z(n9327) );
  OR U13535 ( .A(n9329), .B(n9328), .Z(n9324) );
  IV U13536 ( .A(n9330), .Z(n9328) );
  XOR U13537 ( .A(n9305), .B(n9331), .Z(N29382) );
  XNOR U13538 ( .A(n9308), .B(n9307), .Z(n9331) );
  XNOR U13539 ( .A(n9319), .B(n9332), .Z(n9307) );
  XOR U13540 ( .A(n9323), .B(n9321), .Z(n9332) );
  XOR U13541 ( .A(n9329), .B(n9333), .Z(n9321) );
  XOR U13542 ( .A(n9326), .B(n9330), .Z(n9333) );
  NAND U13543 ( .A(n9334), .B(n9335), .Z(n9330) );
  NAND U13544 ( .A(n9336), .B(n9337), .Z(n9335) );
  NAND U13545 ( .A(n9338), .B(n9339), .Z(n9334) );
  AND U13546 ( .A(n9340), .B(n9341), .Z(n9326) );
  NAND U13547 ( .A(n9342), .B(n9343), .Z(n9341) );
  NAND U13548 ( .A(n9344), .B(n9345), .Z(n9340) );
  NANDN U13549 ( .A(n9346), .B(n9347), .Z(n9329) );
  NANDN U13550 ( .A(n9348), .B(n9349), .Z(n9323) );
  XNOR U13551 ( .A(n9314), .B(n9350), .Z(n9319) );
  XOR U13552 ( .A(n9312), .B(n9316), .Z(n9350) );
  NAND U13553 ( .A(n9351), .B(n9352), .Z(n9316) );
  NAND U13554 ( .A(n9353), .B(n9354), .Z(n9352) );
  NAND U13555 ( .A(n9355), .B(n9356), .Z(n9351) );
  AND U13556 ( .A(n9357), .B(n9358), .Z(n9312) );
  NAND U13557 ( .A(n9359), .B(n9360), .Z(n9358) );
  NAND U13558 ( .A(n9361), .B(n9362), .Z(n9357) );
  AND U13559 ( .A(n9363), .B(n9364), .Z(n9314) );
  NAND U13560 ( .A(n9365), .B(n9366), .Z(n9308) );
  XNOR U13561 ( .A(n9291), .B(n9367), .Z(n9305) );
  XOR U13562 ( .A(n9295), .B(n9293), .Z(n9367) );
  XOR U13563 ( .A(n9301), .B(n9368), .Z(n9293) );
  XOR U13564 ( .A(n9298), .B(n9302), .Z(n9368) );
  NAND U13565 ( .A(n9369), .B(n9370), .Z(n9302) );
  NAND U13566 ( .A(n9371), .B(n9372), .Z(n9370) );
  NAND U13567 ( .A(n9373), .B(n9374), .Z(n9369) );
  AND U13568 ( .A(n9375), .B(n9376), .Z(n9298) );
  NAND U13569 ( .A(n9377), .B(n9378), .Z(n9376) );
  NAND U13570 ( .A(n9379), .B(n9380), .Z(n9375) );
  NANDN U13571 ( .A(n9381), .B(n9382), .Z(n9301) );
  NANDN U13572 ( .A(n9383), .B(n9384), .Z(n9295) );
  XNOR U13573 ( .A(n9286), .B(n9385), .Z(n9291) );
  XOR U13574 ( .A(n9284), .B(n9288), .Z(n9385) );
  NAND U13575 ( .A(n9386), .B(n9387), .Z(n9288) );
  NAND U13576 ( .A(n9388), .B(n9389), .Z(n9387) );
  NAND U13577 ( .A(n9390), .B(n9391), .Z(n9386) );
  AND U13578 ( .A(n9392), .B(n9393), .Z(n9284) );
  NAND U13579 ( .A(n9394), .B(n9395), .Z(n9393) );
  NAND U13580 ( .A(n9396), .B(n9397), .Z(n9392) );
  AND U13581 ( .A(n9398), .B(n9399), .Z(n9286) );
  XOR U13582 ( .A(n9366), .B(n9365), .Z(N29381) );
  XNOR U13583 ( .A(n9384), .B(n9383), .Z(n9365) );
  XNOR U13584 ( .A(n9398), .B(n9399), .Z(n9383) );
  XOR U13585 ( .A(n9395), .B(n9394), .Z(n9399) );
  XOR U13586 ( .A(y[2907]), .B(x[2907]), .Z(n9394) );
  XOR U13587 ( .A(n9397), .B(n9396), .Z(n9395) );
  XOR U13588 ( .A(y[2909]), .B(x[2909]), .Z(n9396) );
  XOR U13589 ( .A(y[2908]), .B(x[2908]), .Z(n9397) );
  XOR U13590 ( .A(n9389), .B(n9388), .Z(n9398) );
  XOR U13591 ( .A(n9391), .B(n9390), .Z(n9388) );
  XOR U13592 ( .A(y[2906]), .B(x[2906]), .Z(n9390) );
  XOR U13593 ( .A(y[2905]), .B(x[2905]), .Z(n9391) );
  XOR U13594 ( .A(y[2904]), .B(x[2904]), .Z(n9389) );
  XNOR U13595 ( .A(n9382), .B(n9381), .Z(n9384) );
  XNOR U13596 ( .A(n9378), .B(n9377), .Z(n9381) );
  XOR U13597 ( .A(n9380), .B(n9379), .Z(n9377) );
  XOR U13598 ( .A(y[2903]), .B(x[2903]), .Z(n9379) );
  XOR U13599 ( .A(y[2902]), .B(x[2902]), .Z(n9380) );
  XOR U13600 ( .A(y[2901]), .B(x[2901]), .Z(n9378) );
  XOR U13601 ( .A(n9372), .B(n9371), .Z(n9382) );
  XOR U13602 ( .A(n9374), .B(n9373), .Z(n9371) );
  XOR U13603 ( .A(y[2900]), .B(x[2900]), .Z(n9373) );
  XOR U13604 ( .A(y[2899]), .B(x[2899]), .Z(n9374) );
  XOR U13605 ( .A(y[2898]), .B(x[2898]), .Z(n9372) );
  XNOR U13606 ( .A(n9349), .B(n9348), .Z(n9366) );
  XNOR U13607 ( .A(n9363), .B(n9364), .Z(n9348) );
  XOR U13608 ( .A(n9360), .B(n9359), .Z(n9364) );
  XOR U13609 ( .A(y[2895]), .B(x[2895]), .Z(n9359) );
  XOR U13610 ( .A(n9362), .B(n9361), .Z(n9360) );
  XOR U13611 ( .A(y[2897]), .B(x[2897]), .Z(n9361) );
  XOR U13612 ( .A(y[2896]), .B(x[2896]), .Z(n9362) );
  XOR U13613 ( .A(n9354), .B(n9353), .Z(n9363) );
  XOR U13614 ( .A(n9356), .B(n9355), .Z(n9353) );
  XOR U13615 ( .A(y[2894]), .B(x[2894]), .Z(n9355) );
  XOR U13616 ( .A(y[2893]), .B(x[2893]), .Z(n9356) );
  XOR U13617 ( .A(y[2892]), .B(x[2892]), .Z(n9354) );
  XNOR U13618 ( .A(n9347), .B(n9346), .Z(n9349) );
  XNOR U13619 ( .A(n9343), .B(n9342), .Z(n9346) );
  XOR U13620 ( .A(n9345), .B(n9344), .Z(n9342) );
  XOR U13621 ( .A(y[2891]), .B(x[2891]), .Z(n9344) );
  XOR U13622 ( .A(y[2890]), .B(x[2890]), .Z(n9345) );
  XOR U13623 ( .A(y[2889]), .B(x[2889]), .Z(n9343) );
  XOR U13624 ( .A(n9337), .B(n9336), .Z(n9347) );
  XOR U13625 ( .A(n9339), .B(n9338), .Z(n9336) );
  XOR U13626 ( .A(y[2888]), .B(x[2888]), .Z(n9338) );
  XOR U13627 ( .A(y[2887]), .B(x[2887]), .Z(n9339) );
  XOR U13628 ( .A(y[2886]), .B(x[2886]), .Z(n9337) );
  NAND U13629 ( .A(n9400), .B(n9401), .Z(N29373) );
  NAND U13630 ( .A(n9402), .B(n9403), .Z(n9401) );
  NANDN U13631 ( .A(n9404), .B(n9405), .Z(n9403) );
  NANDN U13632 ( .A(n9405), .B(n9404), .Z(n9400) );
  XOR U13633 ( .A(n9404), .B(n9406), .Z(N29372) );
  XNOR U13634 ( .A(n9402), .B(n9405), .Z(n9406) );
  NAND U13635 ( .A(n9407), .B(n9408), .Z(n9405) );
  NAND U13636 ( .A(n9409), .B(n9410), .Z(n9408) );
  NANDN U13637 ( .A(n9411), .B(n9412), .Z(n9410) );
  NANDN U13638 ( .A(n9412), .B(n9411), .Z(n9407) );
  AND U13639 ( .A(n9413), .B(n9414), .Z(n9402) );
  NAND U13640 ( .A(n9415), .B(n9416), .Z(n9414) );
  OR U13641 ( .A(n9417), .B(n9418), .Z(n9416) );
  NAND U13642 ( .A(n9418), .B(n9417), .Z(n9413) );
  IV U13643 ( .A(n9419), .Z(n9418) );
  AND U13644 ( .A(n9420), .B(n9421), .Z(n9404) );
  NAND U13645 ( .A(n9422), .B(n9423), .Z(n9421) );
  NANDN U13646 ( .A(n9424), .B(n9425), .Z(n9423) );
  NANDN U13647 ( .A(n9425), .B(n9424), .Z(n9420) );
  XOR U13648 ( .A(n9417), .B(n9426), .Z(N29371) );
  XOR U13649 ( .A(n9415), .B(n9419), .Z(n9426) );
  XNOR U13650 ( .A(n9412), .B(n9427), .Z(n9419) );
  XNOR U13651 ( .A(n9409), .B(n9411), .Z(n9427) );
  AND U13652 ( .A(n9428), .B(n9429), .Z(n9411) );
  NANDN U13653 ( .A(n9430), .B(n9431), .Z(n9429) );
  NANDN U13654 ( .A(n9432), .B(n9433), .Z(n9431) );
  IV U13655 ( .A(n9434), .Z(n9433) );
  NAND U13656 ( .A(n9434), .B(n9432), .Z(n9428) );
  AND U13657 ( .A(n9435), .B(n9436), .Z(n9409) );
  NAND U13658 ( .A(n9437), .B(n9438), .Z(n9436) );
  OR U13659 ( .A(n9439), .B(n9440), .Z(n9438) );
  NAND U13660 ( .A(n9440), .B(n9439), .Z(n9435) );
  IV U13661 ( .A(n9441), .Z(n9440) );
  NAND U13662 ( .A(n9442), .B(n9443), .Z(n9412) );
  NANDN U13663 ( .A(n9444), .B(n9445), .Z(n9443) );
  NAND U13664 ( .A(n9446), .B(n9447), .Z(n9445) );
  OR U13665 ( .A(n9447), .B(n9446), .Z(n9442) );
  IV U13666 ( .A(n9448), .Z(n9446) );
  AND U13667 ( .A(n9449), .B(n9450), .Z(n9415) );
  NAND U13668 ( .A(n9451), .B(n9452), .Z(n9450) );
  NANDN U13669 ( .A(n9453), .B(n9454), .Z(n9452) );
  NANDN U13670 ( .A(n9454), .B(n9453), .Z(n9449) );
  XOR U13671 ( .A(n9425), .B(n9455), .Z(n9417) );
  XNOR U13672 ( .A(n9422), .B(n9424), .Z(n9455) );
  AND U13673 ( .A(n9456), .B(n9457), .Z(n9424) );
  NANDN U13674 ( .A(n9458), .B(n9459), .Z(n9457) );
  NANDN U13675 ( .A(n9460), .B(n9461), .Z(n9459) );
  IV U13676 ( .A(n9462), .Z(n9461) );
  NAND U13677 ( .A(n9462), .B(n9460), .Z(n9456) );
  AND U13678 ( .A(n9463), .B(n9464), .Z(n9422) );
  NAND U13679 ( .A(n9465), .B(n9466), .Z(n9464) );
  OR U13680 ( .A(n9467), .B(n9468), .Z(n9466) );
  NAND U13681 ( .A(n9468), .B(n9467), .Z(n9463) );
  IV U13682 ( .A(n9469), .Z(n9468) );
  NAND U13683 ( .A(n9470), .B(n9471), .Z(n9425) );
  NANDN U13684 ( .A(n9472), .B(n9473), .Z(n9471) );
  NAND U13685 ( .A(n9474), .B(n9475), .Z(n9473) );
  OR U13686 ( .A(n9475), .B(n9474), .Z(n9470) );
  IV U13687 ( .A(n9476), .Z(n9474) );
  XOR U13688 ( .A(n9451), .B(n9477), .Z(N29370) );
  XNOR U13689 ( .A(n9454), .B(n9453), .Z(n9477) );
  XNOR U13690 ( .A(n9465), .B(n9478), .Z(n9453) );
  XOR U13691 ( .A(n9469), .B(n9467), .Z(n9478) );
  XOR U13692 ( .A(n9475), .B(n9479), .Z(n9467) );
  XOR U13693 ( .A(n9472), .B(n9476), .Z(n9479) );
  NAND U13694 ( .A(n9480), .B(n9481), .Z(n9476) );
  NAND U13695 ( .A(n9482), .B(n9483), .Z(n9481) );
  NAND U13696 ( .A(n9484), .B(n9485), .Z(n9480) );
  AND U13697 ( .A(n9486), .B(n9487), .Z(n9472) );
  NAND U13698 ( .A(n9488), .B(n9489), .Z(n9487) );
  NAND U13699 ( .A(n9490), .B(n9491), .Z(n9486) );
  NANDN U13700 ( .A(n9492), .B(n9493), .Z(n9475) );
  NANDN U13701 ( .A(n9494), .B(n9495), .Z(n9469) );
  XNOR U13702 ( .A(n9460), .B(n9496), .Z(n9465) );
  XOR U13703 ( .A(n9458), .B(n9462), .Z(n9496) );
  NAND U13704 ( .A(n9497), .B(n9498), .Z(n9462) );
  NAND U13705 ( .A(n9499), .B(n9500), .Z(n9498) );
  NAND U13706 ( .A(n9501), .B(n9502), .Z(n9497) );
  AND U13707 ( .A(n9503), .B(n9504), .Z(n9458) );
  NAND U13708 ( .A(n9505), .B(n9506), .Z(n9504) );
  NAND U13709 ( .A(n9507), .B(n9508), .Z(n9503) );
  AND U13710 ( .A(n9509), .B(n9510), .Z(n9460) );
  NAND U13711 ( .A(n9511), .B(n9512), .Z(n9454) );
  XNOR U13712 ( .A(n9437), .B(n9513), .Z(n9451) );
  XOR U13713 ( .A(n9441), .B(n9439), .Z(n9513) );
  XOR U13714 ( .A(n9447), .B(n9514), .Z(n9439) );
  XOR U13715 ( .A(n9444), .B(n9448), .Z(n9514) );
  NAND U13716 ( .A(n9515), .B(n9516), .Z(n9448) );
  NAND U13717 ( .A(n9517), .B(n9518), .Z(n9516) );
  NAND U13718 ( .A(n9519), .B(n9520), .Z(n9515) );
  AND U13719 ( .A(n9521), .B(n9522), .Z(n9444) );
  NAND U13720 ( .A(n9523), .B(n9524), .Z(n9522) );
  NAND U13721 ( .A(n9525), .B(n9526), .Z(n9521) );
  NANDN U13722 ( .A(n9527), .B(n9528), .Z(n9447) );
  NANDN U13723 ( .A(n9529), .B(n9530), .Z(n9441) );
  XNOR U13724 ( .A(n9432), .B(n9531), .Z(n9437) );
  XOR U13725 ( .A(n9430), .B(n9434), .Z(n9531) );
  NAND U13726 ( .A(n9532), .B(n9533), .Z(n9434) );
  NAND U13727 ( .A(n9534), .B(n9535), .Z(n9533) );
  NAND U13728 ( .A(n9536), .B(n9537), .Z(n9532) );
  AND U13729 ( .A(n9538), .B(n9539), .Z(n9430) );
  NAND U13730 ( .A(n9540), .B(n9541), .Z(n9539) );
  NAND U13731 ( .A(n9542), .B(n9543), .Z(n9538) );
  AND U13732 ( .A(n9544), .B(n9545), .Z(n9432) );
  XOR U13733 ( .A(n9512), .B(n9511), .Z(N29369) );
  XNOR U13734 ( .A(n9530), .B(n9529), .Z(n9511) );
  XNOR U13735 ( .A(n9544), .B(n9545), .Z(n9529) );
  XOR U13736 ( .A(n9541), .B(n9540), .Z(n9545) );
  XOR U13737 ( .A(y[2883]), .B(x[2883]), .Z(n9540) );
  XOR U13738 ( .A(n9543), .B(n9542), .Z(n9541) );
  XOR U13739 ( .A(y[2885]), .B(x[2885]), .Z(n9542) );
  XOR U13740 ( .A(y[2884]), .B(x[2884]), .Z(n9543) );
  XOR U13741 ( .A(n9535), .B(n9534), .Z(n9544) );
  XOR U13742 ( .A(n9537), .B(n9536), .Z(n9534) );
  XOR U13743 ( .A(y[2882]), .B(x[2882]), .Z(n9536) );
  XOR U13744 ( .A(y[2881]), .B(x[2881]), .Z(n9537) );
  XOR U13745 ( .A(y[2880]), .B(x[2880]), .Z(n9535) );
  XNOR U13746 ( .A(n9528), .B(n9527), .Z(n9530) );
  XNOR U13747 ( .A(n9524), .B(n9523), .Z(n9527) );
  XOR U13748 ( .A(n9526), .B(n9525), .Z(n9523) );
  XOR U13749 ( .A(y[2879]), .B(x[2879]), .Z(n9525) );
  XOR U13750 ( .A(y[2878]), .B(x[2878]), .Z(n9526) );
  XOR U13751 ( .A(y[2877]), .B(x[2877]), .Z(n9524) );
  XOR U13752 ( .A(n9518), .B(n9517), .Z(n9528) );
  XOR U13753 ( .A(n9520), .B(n9519), .Z(n9517) );
  XOR U13754 ( .A(y[2876]), .B(x[2876]), .Z(n9519) );
  XOR U13755 ( .A(y[2875]), .B(x[2875]), .Z(n9520) );
  XOR U13756 ( .A(y[2874]), .B(x[2874]), .Z(n9518) );
  XNOR U13757 ( .A(n9495), .B(n9494), .Z(n9512) );
  XNOR U13758 ( .A(n9509), .B(n9510), .Z(n9494) );
  XOR U13759 ( .A(n9506), .B(n9505), .Z(n9510) );
  XOR U13760 ( .A(y[2871]), .B(x[2871]), .Z(n9505) );
  XOR U13761 ( .A(n9508), .B(n9507), .Z(n9506) );
  XOR U13762 ( .A(y[2873]), .B(x[2873]), .Z(n9507) );
  XOR U13763 ( .A(y[2872]), .B(x[2872]), .Z(n9508) );
  XOR U13764 ( .A(n9500), .B(n9499), .Z(n9509) );
  XOR U13765 ( .A(n9502), .B(n9501), .Z(n9499) );
  XOR U13766 ( .A(y[2870]), .B(x[2870]), .Z(n9501) );
  XOR U13767 ( .A(y[2869]), .B(x[2869]), .Z(n9502) );
  XOR U13768 ( .A(y[2868]), .B(x[2868]), .Z(n9500) );
  XNOR U13769 ( .A(n9493), .B(n9492), .Z(n9495) );
  XNOR U13770 ( .A(n9489), .B(n9488), .Z(n9492) );
  XOR U13771 ( .A(n9491), .B(n9490), .Z(n9488) );
  XOR U13772 ( .A(y[2867]), .B(x[2867]), .Z(n9490) );
  XOR U13773 ( .A(y[2866]), .B(x[2866]), .Z(n9491) );
  XOR U13774 ( .A(y[2865]), .B(x[2865]), .Z(n9489) );
  XOR U13775 ( .A(n9483), .B(n9482), .Z(n9493) );
  XOR U13776 ( .A(n9485), .B(n9484), .Z(n9482) );
  XOR U13777 ( .A(y[2864]), .B(x[2864]), .Z(n9484) );
  XOR U13778 ( .A(y[2863]), .B(x[2863]), .Z(n9485) );
  XOR U13779 ( .A(y[2862]), .B(x[2862]), .Z(n9483) );
  NAND U13780 ( .A(n9546), .B(n9547), .Z(N29361) );
  NAND U13781 ( .A(n9548), .B(n9549), .Z(n9547) );
  NANDN U13782 ( .A(n9550), .B(n9551), .Z(n9549) );
  NANDN U13783 ( .A(n9551), .B(n9550), .Z(n9546) );
  XOR U13784 ( .A(n9550), .B(n9552), .Z(N29360) );
  XNOR U13785 ( .A(n9548), .B(n9551), .Z(n9552) );
  NAND U13786 ( .A(n9553), .B(n9554), .Z(n9551) );
  NAND U13787 ( .A(n9555), .B(n9556), .Z(n9554) );
  NANDN U13788 ( .A(n9557), .B(n9558), .Z(n9556) );
  NANDN U13789 ( .A(n9558), .B(n9557), .Z(n9553) );
  AND U13790 ( .A(n9559), .B(n9560), .Z(n9548) );
  NAND U13791 ( .A(n9561), .B(n9562), .Z(n9560) );
  OR U13792 ( .A(n9563), .B(n9564), .Z(n9562) );
  NAND U13793 ( .A(n9564), .B(n9563), .Z(n9559) );
  IV U13794 ( .A(n9565), .Z(n9564) );
  AND U13795 ( .A(n9566), .B(n9567), .Z(n9550) );
  NAND U13796 ( .A(n9568), .B(n9569), .Z(n9567) );
  NANDN U13797 ( .A(n9570), .B(n9571), .Z(n9569) );
  NANDN U13798 ( .A(n9571), .B(n9570), .Z(n9566) );
  XOR U13799 ( .A(n9563), .B(n9572), .Z(N29359) );
  XOR U13800 ( .A(n9561), .B(n9565), .Z(n9572) );
  XNOR U13801 ( .A(n9558), .B(n9573), .Z(n9565) );
  XNOR U13802 ( .A(n9555), .B(n9557), .Z(n9573) );
  AND U13803 ( .A(n9574), .B(n9575), .Z(n9557) );
  NANDN U13804 ( .A(n9576), .B(n9577), .Z(n9575) );
  NANDN U13805 ( .A(n9578), .B(n9579), .Z(n9577) );
  IV U13806 ( .A(n9580), .Z(n9579) );
  NAND U13807 ( .A(n9580), .B(n9578), .Z(n9574) );
  AND U13808 ( .A(n9581), .B(n9582), .Z(n9555) );
  NAND U13809 ( .A(n9583), .B(n9584), .Z(n9582) );
  OR U13810 ( .A(n9585), .B(n9586), .Z(n9584) );
  NAND U13811 ( .A(n9586), .B(n9585), .Z(n9581) );
  IV U13812 ( .A(n9587), .Z(n9586) );
  NAND U13813 ( .A(n9588), .B(n9589), .Z(n9558) );
  NANDN U13814 ( .A(n9590), .B(n9591), .Z(n9589) );
  NAND U13815 ( .A(n9592), .B(n9593), .Z(n9591) );
  OR U13816 ( .A(n9593), .B(n9592), .Z(n9588) );
  IV U13817 ( .A(n9594), .Z(n9592) );
  AND U13818 ( .A(n9595), .B(n9596), .Z(n9561) );
  NAND U13819 ( .A(n9597), .B(n9598), .Z(n9596) );
  NANDN U13820 ( .A(n9599), .B(n9600), .Z(n9598) );
  NANDN U13821 ( .A(n9600), .B(n9599), .Z(n9595) );
  XOR U13822 ( .A(n9571), .B(n9601), .Z(n9563) );
  XNOR U13823 ( .A(n9568), .B(n9570), .Z(n9601) );
  AND U13824 ( .A(n9602), .B(n9603), .Z(n9570) );
  NANDN U13825 ( .A(n9604), .B(n9605), .Z(n9603) );
  NANDN U13826 ( .A(n9606), .B(n9607), .Z(n9605) );
  IV U13827 ( .A(n9608), .Z(n9607) );
  NAND U13828 ( .A(n9608), .B(n9606), .Z(n9602) );
  AND U13829 ( .A(n9609), .B(n9610), .Z(n9568) );
  NAND U13830 ( .A(n9611), .B(n9612), .Z(n9610) );
  OR U13831 ( .A(n9613), .B(n9614), .Z(n9612) );
  NAND U13832 ( .A(n9614), .B(n9613), .Z(n9609) );
  IV U13833 ( .A(n9615), .Z(n9614) );
  NAND U13834 ( .A(n9616), .B(n9617), .Z(n9571) );
  NANDN U13835 ( .A(n9618), .B(n9619), .Z(n9617) );
  NAND U13836 ( .A(n9620), .B(n9621), .Z(n9619) );
  OR U13837 ( .A(n9621), .B(n9620), .Z(n9616) );
  IV U13838 ( .A(n9622), .Z(n9620) );
  XOR U13839 ( .A(n9597), .B(n9623), .Z(N29358) );
  XNOR U13840 ( .A(n9600), .B(n9599), .Z(n9623) );
  XNOR U13841 ( .A(n9611), .B(n9624), .Z(n9599) );
  XOR U13842 ( .A(n9615), .B(n9613), .Z(n9624) );
  XOR U13843 ( .A(n9621), .B(n9625), .Z(n9613) );
  XOR U13844 ( .A(n9618), .B(n9622), .Z(n9625) );
  NAND U13845 ( .A(n9626), .B(n9627), .Z(n9622) );
  NAND U13846 ( .A(n9628), .B(n9629), .Z(n9627) );
  NAND U13847 ( .A(n9630), .B(n9631), .Z(n9626) );
  AND U13848 ( .A(n9632), .B(n9633), .Z(n9618) );
  NAND U13849 ( .A(n9634), .B(n9635), .Z(n9633) );
  NAND U13850 ( .A(n9636), .B(n9637), .Z(n9632) );
  NANDN U13851 ( .A(n9638), .B(n9639), .Z(n9621) );
  NANDN U13852 ( .A(n9640), .B(n9641), .Z(n9615) );
  XNOR U13853 ( .A(n9606), .B(n9642), .Z(n9611) );
  XOR U13854 ( .A(n9604), .B(n9608), .Z(n9642) );
  NAND U13855 ( .A(n9643), .B(n9644), .Z(n9608) );
  NAND U13856 ( .A(n9645), .B(n9646), .Z(n9644) );
  NAND U13857 ( .A(n9647), .B(n9648), .Z(n9643) );
  AND U13858 ( .A(n9649), .B(n9650), .Z(n9604) );
  NAND U13859 ( .A(n9651), .B(n9652), .Z(n9650) );
  NAND U13860 ( .A(n9653), .B(n9654), .Z(n9649) );
  AND U13861 ( .A(n9655), .B(n9656), .Z(n9606) );
  NAND U13862 ( .A(n9657), .B(n9658), .Z(n9600) );
  XNOR U13863 ( .A(n9583), .B(n9659), .Z(n9597) );
  XOR U13864 ( .A(n9587), .B(n9585), .Z(n9659) );
  XOR U13865 ( .A(n9593), .B(n9660), .Z(n9585) );
  XOR U13866 ( .A(n9590), .B(n9594), .Z(n9660) );
  NAND U13867 ( .A(n9661), .B(n9662), .Z(n9594) );
  NAND U13868 ( .A(n9663), .B(n9664), .Z(n9662) );
  NAND U13869 ( .A(n9665), .B(n9666), .Z(n9661) );
  AND U13870 ( .A(n9667), .B(n9668), .Z(n9590) );
  NAND U13871 ( .A(n9669), .B(n9670), .Z(n9668) );
  NAND U13872 ( .A(n9671), .B(n9672), .Z(n9667) );
  NANDN U13873 ( .A(n9673), .B(n9674), .Z(n9593) );
  NANDN U13874 ( .A(n9675), .B(n9676), .Z(n9587) );
  XNOR U13875 ( .A(n9578), .B(n9677), .Z(n9583) );
  XOR U13876 ( .A(n9576), .B(n9580), .Z(n9677) );
  NAND U13877 ( .A(n9678), .B(n9679), .Z(n9580) );
  NAND U13878 ( .A(n9680), .B(n9681), .Z(n9679) );
  NAND U13879 ( .A(n9682), .B(n9683), .Z(n9678) );
  AND U13880 ( .A(n9684), .B(n9685), .Z(n9576) );
  NAND U13881 ( .A(n9686), .B(n9687), .Z(n9685) );
  NAND U13882 ( .A(n9688), .B(n9689), .Z(n9684) );
  AND U13883 ( .A(n9690), .B(n9691), .Z(n9578) );
  XOR U13884 ( .A(n9658), .B(n9657), .Z(N29357) );
  XNOR U13885 ( .A(n9676), .B(n9675), .Z(n9657) );
  XNOR U13886 ( .A(n9690), .B(n9691), .Z(n9675) );
  XOR U13887 ( .A(n9687), .B(n9686), .Z(n9691) );
  XOR U13888 ( .A(y[2859]), .B(x[2859]), .Z(n9686) );
  XOR U13889 ( .A(n9689), .B(n9688), .Z(n9687) );
  XOR U13890 ( .A(y[2861]), .B(x[2861]), .Z(n9688) );
  XOR U13891 ( .A(y[2860]), .B(x[2860]), .Z(n9689) );
  XOR U13892 ( .A(n9681), .B(n9680), .Z(n9690) );
  XOR U13893 ( .A(n9683), .B(n9682), .Z(n9680) );
  XOR U13894 ( .A(y[2858]), .B(x[2858]), .Z(n9682) );
  XOR U13895 ( .A(y[2857]), .B(x[2857]), .Z(n9683) );
  XOR U13896 ( .A(y[2856]), .B(x[2856]), .Z(n9681) );
  XNOR U13897 ( .A(n9674), .B(n9673), .Z(n9676) );
  XNOR U13898 ( .A(n9670), .B(n9669), .Z(n9673) );
  XOR U13899 ( .A(n9672), .B(n9671), .Z(n9669) );
  XOR U13900 ( .A(y[2855]), .B(x[2855]), .Z(n9671) );
  XOR U13901 ( .A(y[2854]), .B(x[2854]), .Z(n9672) );
  XOR U13902 ( .A(y[2853]), .B(x[2853]), .Z(n9670) );
  XOR U13903 ( .A(n9664), .B(n9663), .Z(n9674) );
  XOR U13904 ( .A(n9666), .B(n9665), .Z(n9663) );
  XOR U13905 ( .A(y[2852]), .B(x[2852]), .Z(n9665) );
  XOR U13906 ( .A(y[2851]), .B(x[2851]), .Z(n9666) );
  XOR U13907 ( .A(y[2850]), .B(x[2850]), .Z(n9664) );
  XNOR U13908 ( .A(n9641), .B(n9640), .Z(n9658) );
  XNOR U13909 ( .A(n9655), .B(n9656), .Z(n9640) );
  XOR U13910 ( .A(n9652), .B(n9651), .Z(n9656) );
  XOR U13911 ( .A(y[2847]), .B(x[2847]), .Z(n9651) );
  XOR U13912 ( .A(n9654), .B(n9653), .Z(n9652) );
  XOR U13913 ( .A(y[2849]), .B(x[2849]), .Z(n9653) );
  XOR U13914 ( .A(y[2848]), .B(x[2848]), .Z(n9654) );
  XOR U13915 ( .A(n9646), .B(n9645), .Z(n9655) );
  XOR U13916 ( .A(n9648), .B(n9647), .Z(n9645) );
  XOR U13917 ( .A(y[2846]), .B(x[2846]), .Z(n9647) );
  XOR U13918 ( .A(y[2845]), .B(x[2845]), .Z(n9648) );
  XOR U13919 ( .A(y[2844]), .B(x[2844]), .Z(n9646) );
  XNOR U13920 ( .A(n9639), .B(n9638), .Z(n9641) );
  XNOR U13921 ( .A(n9635), .B(n9634), .Z(n9638) );
  XOR U13922 ( .A(n9637), .B(n9636), .Z(n9634) );
  XOR U13923 ( .A(y[2843]), .B(x[2843]), .Z(n9636) );
  XOR U13924 ( .A(y[2842]), .B(x[2842]), .Z(n9637) );
  XOR U13925 ( .A(y[2841]), .B(x[2841]), .Z(n9635) );
  XOR U13926 ( .A(n9629), .B(n9628), .Z(n9639) );
  XOR U13927 ( .A(n9631), .B(n9630), .Z(n9628) );
  XOR U13928 ( .A(y[2840]), .B(x[2840]), .Z(n9630) );
  XOR U13929 ( .A(y[2839]), .B(x[2839]), .Z(n9631) );
  XOR U13930 ( .A(y[2838]), .B(x[2838]), .Z(n9629) );
  NAND U13931 ( .A(n9692), .B(n9693), .Z(N29349) );
  NAND U13932 ( .A(n9694), .B(n9695), .Z(n9693) );
  NANDN U13933 ( .A(n9696), .B(n9697), .Z(n9695) );
  NANDN U13934 ( .A(n9697), .B(n9696), .Z(n9692) );
  XOR U13935 ( .A(n9696), .B(n9698), .Z(N29348) );
  XNOR U13936 ( .A(n9694), .B(n9697), .Z(n9698) );
  NAND U13937 ( .A(n9699), .B(n9700), .Z(n9697) );
  NAND U13938 ( .A(n9701), .B(n9702), .Z(n9700) );
  NANDN U13939 ( .A(n9703), .B(n9704), .Z(n9702) );
  NANDN U13940 ( .A(n9704), .B(n9703), .Z(n9699) );
  AND U13941 ( .A(n9705), .B(n9706), .Z(n9694) );
  NAND U13942 ( .A(n9707), .B(n9708), .Z(n9706) );
  OR U13943 ( .A(n9709), .B(n9710), .Z(n9708) );
  NAND U13944 ( .A(n9710), .B(n9709), .Z(n9705) );
  IV U13945 ( .A(n9711), .Z(n9710) );
  AND U13946 ( .A(n9712), .B(n9713), .Z(n9696) );
  NAND U13947 ( .A(n9714), .B(n9715), .Z(n9713) );
  NANDN U13948 ( .A(n9716), .B(n9717), .Z(n9715) );
  NANDN U13949 ( .A(n9717), .B(n9716), .Z(n9712) );
  XOR U13950 ( .A(n9709), .B(n9718), .Z(N29347) );
  XOR U13951 ( .A(n9707), .B(n9711), .Z(n9718) );
  XNOR U13952 ( .A(n9704), .B(n9719), .Z(n9711) );
  XNOR U13953 ( .A(n9701), .B(n9703), .Z(n9719) );
  AND U13954 ( .A(n9720), .B(n9721), .Z(n9703) );
  NANDN U13955 ( .A(n9722), .B(n9723), .Z(n9721) );
  NANDN U13956 ( .A(n9724), .B(n9725), .Z(n9723) );
  IV U13957 ( .A(n9726), .Z(n9725) );
  NAND U13958 ( .A(n9726), .B(n9724), .Z(n9720) );
  AND U13959 ( .A(n9727), .B(n9728), .Z(n9701) );
  NAND U13960 ( .A(n9729), .B(n9730), .Z(n9728) );
  OR U13961 ( .A(n9731), .B(n9732), .Z(n9730) );
  NAND U13962 ( .A(n9732), .B(n9731), .Z(n9727) );
  IV U13963 ( .A(n9733), .Z(n9732) );
  NAND U13964 ( .A(n9734), .B(n9735), .Z(n9704) );
  NANDN U13965 ( .A(n9736), .B(n9737), .Z(n9735) );
  NAND U13966 ( .A(n9738), .B(n9739), .Z(n9737) );
  OR U13967 ( .A(n9739), .B(n9738), .Z(n9734) );
  IV U13968 ( .A(n9740), .Z(n9738) );
  AND U13969 ( .A(n9741), .B(n9742), .Z(n9707) );
  NAND U13970 ( .A(n9743), .B(n9744), .Z(n9742) );
  NANDN U13971 ( .A(n9745), .B(n9746), .Z(n9744) );
  NANDN U13972 ( .A(n9746), .B(n9745), .Z(n9741) );
  XOR U13973 ( .A(n9717), .B(n9747), .Z(n9709) );
  XNOR U13974 ( .A(n9714), .B(n9716), .Z(n9747) );
  AND U13975 ( .A(n9748), .B(n9749), .Z(n9716) );
  NANDN U13976 ( .A(n9750), .B(n9751), .Z(n9749) );
  NANDN U13977 ( .A(n9752), .B(n9753), .Z(n9751) );
  IV U13978 ( .A(n9754), .Z(n9753) );
  NAND U13979 ( .A(n9754), .B(n9752), .Z(n9748) );
  AND U13980 ( .A(n9755), .B(n9756), .Z(n9714) );
  NAND U13981 ( .A(n9757), .B(n9758), .Z(n9756) );
  OR U13982 ( .A(n9759), .B(n9760), .Z(n9758) );
  NAND U13983 ( .A(n9760), .B(n9759), .Z(n9755) );
  IV U13984 ( .A(n9761), .Z(n9760) );
  NAND U13985 ( .A(n9762), .B(n9763), .Z(n9717) );
  NANDN U13986 ( .A(n9764), .B(n9765), .Z(n9763) );
  NAND U13987 ( .A(n9766), .B(n9767), .Z(n9765) );
  OR U13988 ( .A(n9767), .B(n9766), .Z(n9762) );
  IV U13989 ( .A(n9768), .Z(n9766) );
  XOR U13990 ( .A(n9743), .B(n9769), .Z(N29346) );
  XNOR U13991 ( .A(n9746), .B(n9745), .Z(n9769) );
  XNOR U13992 ( .A(n9757), .B(n9770), .Z(n9745) );
  XOR U13993 ( .A(n9761), .B(n9759), .Z(n9770) );
  XOR U13994 ( .A(n9767), .B(n9771), .Z(n9759) );
  XOR U13995 ( .A(n9764), .B(n9768), .Z(n9771) );
  NAND U13996 ( .A(n9772), .B(n9773), .Z(n9768) );
  NAND U13997 ( .A(n9774), .B(n9775), .Z(n9773) );
  NAND U13998 ( .A(n9776), .B(n9777), .Z(n9772) );
  AND U13999 ( .A(n9778), .B(n9779), .Z(n9764) );
  NAND U14000 ( .A(n9780), .B(n9781), .Z(n9779) );
  NAND U14001 ( .A(n9782), .B(n9783), .Z(n9778) );
  NANDN U14002 ( .A(n9784), .B(n9785), .Z(n9767) );
  NANDN U14003 ( .A(n9786), .B(n9787), .Z(n9761) );
  XNOR U14004 ( .A(n9752), .B(n9788), .Z(n9757) );
  XOR U14005 ( .A(n9750), .B(n9754), .Z(n9788) );
  NAND U14006 ( .A(n9789), .B(n9790), .Z(n9754) );
  NAND U14007 ( .A(n9791), .B(n9792), .Z(n9790) );
  NAND U14008 ( .A(n9793), .B(n9794), .Z(n9789) );
  AND U14009 ( .A(n9795), .B(n9796), .Z(n9750) );
  NAND U14010 ( .A(n9797), .B(n9798), .Z(n9796) );
  NAND U14011 ( .A(n9799), .B(n9800), .Z(n9795) );
  AND U14012 ( .A(n9801), .B(n9802), .Z(n9752) );
  NAND U14013 ( .A(n9803), .B(n9804), .Z(n9746) );
  XNOR U14014 ( .A(n9729), .B(n9805), .Z(n9743) );
  XOR U14015 ( .A(n9733), .B(n9731), .Z(n9805) );
  XOR U14016 ( .A(n9739), .B(n9806), .Z(n9731) );
  XOR U14017 ( .A(n9736), .B(n9740), .Z(n9806) );
  NAND U14018 ( .A(n9807), .B(n9808), .Z(n9740) );
  NAND U14019 ( .A(n9809), .B(n9810), .Z(n9808) );
  NAND U14020 ( .A(n9811), .B(n9812), .Z(n9807) );
  AND U14021 ( .A(n9813), .B(n9814), .Z(n9736) );
  NAND U14022 ( .A(n9815), .B(n9816), .Z(n9814) );
  NAND U14023 ( .A(n9817), .B(n9818), .Z(n9813) );
  NANDN U14024 ( .A(n9819), .B(n9820), .Z(n9739) );
  NANDN U14025 ( .A(n9821), .B(n9822), .Z(n9733) );
  XNOR U14026 ( .A(n9724), .B(n9823), .Z(n9729) );
  XOR U14027 ( .A(n9722), .B(n9726), .Z(n9823) );
  NAND U14028 ( .A(n9824), .B(n9825), .Z(n9726) );
  NAND U14029 ( .A(n9826), .B(n9827), .Z(n9825) );
  NAND U14030 ( .A(n9828), .B(n9829), .Z(n9824) );
  AND U14031 ( .A(n9830), .B(n9831), .Z(n9722) );
  NAND U14032 ( .A(n9832), .B(n9833), .Z(n9831) );
  NAND U14033 ( .A(n9834), .B(n9835), .Z(n9830) );
  AND U14034 ( .A(n9836), .B(n9837), .Z(n9724) );
  XOR U14035 ( .A(n9804), .B(n9803), .Z(N29345) );
  XNOR U14036 ( .A(n9822), .B(n9821), .Z(n9803) );
  XNOR U14037 ( .A(n9836), .B(n9837), .Z(n9821) );
  XOR U14038 ( .A(n9833), .B(n9832), .Z(n9837) );
  XOR U14039 ( .A(y[2835]), .B(x[2835]), .Z(n9832) );
  XOR U14040 ( .A(n9835), .B(n9834), .Z(n9833) );
  XOR U14041 ( .A(y[2837]), .B(x[2837]), .Z(n9834) );
  XOR U14042 ( .A(y[2836]), .B(x[2836]), .Z(n9835) );
  XOR U14043 ( .A(n9827), .B(n9826), .Z(n9836) );
  XOR U14044 ( .A(n9829), .B(n9828), .Z(n9826) );
  XOR U14045 ( .A(y[2834]), .B(x[2834]), .Z(n9828) );
  XOR U14046 ( .A(y[2833]), .B(x[2833]), .Z(n9829) );
  XOR U14047 ( .A(y[2832]), .B(x[2832]), .Z(n9827) );
  XNOR U14048 ( .A(n9820), .B(n9819), .Z(n9822) );
  XNOR U14049 ( .A(n9816), .B(n9815), .Z(n9819) );
  XOR U14050 ( .A(n9818), .B(n9817), .Z(n9815) );
  XOR U14051 ( .A(y[2831]), .B(x[2831]), .Z(n9817) );
  XOR U14052 ( .A(y[2830]), .B(x[2830]), .Z(n9818) );
  XOR U14053 ( .A(y[2829]), .B(x[2829]), .Z(n9816) );
  XOR U14054 ( .A(n9810), .B(n9809), .Z(n9820) );
  XOR U14055 ( .A(n9812), .B(n9811), .Z(n9809) );
  XOR U14056 ( .A(y[2828]), .B(x[2828]), .Z(n9811) );
  XOR U14057 ( .A(y[2827]), .B(x[2827]), .Z(n9812) );
  XOR U14058 ( .A(y[2826]), .B(x[2826]), .Z(n9810) );
  XNOR U14059 ( .A(n9787), .B(n9786), .Z(n9804) );
  XNOR U14060 ( .A(n9801), .B(n9802), .Z(n9786) );
  XOR U14061 ( .A(n9798), .B(n9797), .Z(n9802) );
  XOR U14062 ( .A(y[2823]), .B(x[2823]), .Z(n9797) );
  XOR U14063 ( .A(n9800), .B(n9799), .Z(n9798) );
  XOR U14064 ( .A(y[2825]), .B(x[2825]), .Z(n9799) );
  XOR U14065 ( .A(y[2824]), .B(x[2824]), .Z(n9800) );
  XOR U14066 ( .A(n9792), .B(n9791), .Z(n9801) );
  XOR U14067 ( .A(n9794), .B(n9793), .Z(n9791) );
  XOR U14068 ( .A(y[2822]), .B(x[2822]), .Z(n9793) );
  XOR U14069 ( .A(y[2821]), .B(x[2821]), .Z(n9794) );
  XOR U14070 ( .A(y[2820]), .B(x[2820]), .Z(n9792) );
  XNOR U14071 ( .A(n9785), .B(n9784), .Z(n9787) );
  XNOR U14072 ( .A(n9781), .B(n9780), .Z(n9784) );
  XOR U14073 ( .A(n9783), .B(n9782), .Z(n9780) );
  XOR U14074 ( .A(y[2819]), .B(x[2819]), .Z(n9782) );
  XOR U14075 ( .A(y[2818]), .B(x[2818]), .Z(n9783) );
  XOR U14076 ( .A(y[2817]), .B(x[2817]), .Z(n9781) );
  XOR U14077 ( .A(n9775), .B(n9774), .Z(n9785) );
  XOR U14078 ( .A(n9777), .B(n9776), .Z(n9774) );
  XOR U14079 ( .A(y[2816]), .B(x[2816]), .Z(n9776) );
  XOR U14080 ( .A(y[2815]), .B(x[2815]), .Z(n9777) );
  XOR U14081 ( .A(y[2814]), .B(x[2814]), .Z(n9775) );
  NAND U14082 ( .A(n9838), .B(n9839), .Z(N29337) );
  NAND U14083 ( .A(n9840), .B(n9841), .Z(n9839) );
  NANDN U14084 ( .A(n9842), .B(n9843), .Z(n9841) );
  NANDN U14085 ( .A(n9843), .B(n9842), .Z(n9838) );
  XOR U14086 ( .A(n9842), .B(n9844), .Z(N29336) );
  XNOR U14087 ( .A(n9840), .B(n9843), .Z(n9844) );
  NAND U14088 ( .A(n9845), .B(n9846), .Z(n9843) );
  NAND U14089 ( .A(n9847), .B(n9848), .Z(n9846) );
  NANDN U14090 ( .A(n9849), .B(n9850), .Z(n9848) );
  NANDN U14091 ( .A(n9850), .B(n9849), .Z(n9845) );
  AND U14092 ( .A(n9851), .B(n9852), .Z(n9840) );
  NAND U14093 ( .A(n9853), .B(n9854), .Z(n9852) );
  OR U14094 ( .A(n9855), .B(n9856), .Z(n9854) );
  NAND U14095 ( .A(n9856), .B(n9855), .Z(n9851) );
  IV U14096 ( .A(n9857), .Z(n9856) );
  AND U14097 ( .A(n9858), .B(n9859), .Z(n9842) );
  NAND U14098 ( .A(n9860), .B(n9861), .Z(n9859) );
  NANDN U14099 ( .A(n9862), .B(n9863), .Z(n9861) );
  NANDN U14100 ( .A(n9863), .B(n9862), .Z(n9858) );
  XOR U14101 ( .A(n9855), .B(n9864), .Z(N29335) );
  XOR U14102 ( .A(n9853), .B(n9857), .Z(n9864) );
  XNOR U14103 ( .A(n9850), .B(n9865), .Z(n9857) );
  XNOR U14104 ( .A(n9847), .B(n9849), .Z(n9865) );
  AND U14105 ( .A(n9866), .B(n9867), .Z(n9849) );
  NANDN U14106 ( .A(n9868), .B(n9869), .Z(n9867) );
  NANDN U14107 ( .A(n9870), .B(n9871), .Z(n9869) );
  IV U14108 ( .A(n9872), .Z(n9871) );
  NAND U14109 ( .A(n9872), .B(n9870), .Z(n9866) );
  AND U14110 ( .A(n9873), .B(n9874), .Z(n9847) );
  NAND U14111 ( .A(n9875), .B(n9876), .Z(n9874) );
  OR U14112 ( .A(n9877), .B(n9878), .Z(n9876) );
  NAND U14113 ( .A(n9878), .B(n9877), .Z(n9873) );
  IV U14114 ( .A(n9879), .Z(n9878) );
  NAND U14115 ( .A(n9880), .B(n9881), .Z(n9850) );
  NANDN U14116 ( .A(n9882), .B(n9883), .Z(n9881) );
  NAND U14117 ( .A(n9884), .B(n9885), .Z(n9883) );
  OR U14118 ( .A(n9885), .B(n9884), .Z(n9880) );
  IV U14119 ( .A(n9886), .Z(n9884) );
  AND U14120 ( .A(n9887), .B(n9888), .Z(n9853) );
  NAND U14121 ( .A(n9889), .B(n9890), .Z(n9888) );
  NANDN U14122 ( .A(n9891), .B(n9892), .Z(n9890) );
  NANDN U14123 ( .A(n9892), .B(n9891), .Z(n9887) );
  XOR U14124 ( .A(n9863), .B(n9893), .Z(n9855) );
  XNOR U14125 ( .A(n9860), .B(n9862), .Z(n9893) );
  AND U14126 ( .A(n9894), .B(n9895), .Z(n9862) );
  NANDN U14127 ( .A(n9896), .B(n9897), .Z(n9895) );
  NANDN U14128 ( .A(n9898), .B(n9899), .Z(n9897) );
  IV U14129 ( .A(n9900), .Z(n9899) );
  NAND U14130 ( .A(n9900), .B(n9898), .Z(n9894) );
  AND U14131 ( .A(n9901), .B(n9902), .Z(n9860) );
  NAND U14132 ( .A(n9903), .B(n9904), .Z(n9902) );
  OR U14133 ( .A(n9905), .B(n9906), .Z(n9904) );
  NAND U14134 ( .A(n9906), .B(n9905), .Z(n9901) );
  IV U14135 ( .A(n9907), .Z(n9906) );
  NAND U14136 ( .A(n9908), .B(n9909), .Z(n9863) );
  NANDN U14137 ( .A(n9910), .B(n9911), .Z(n9909) );
  NAND U14138 ( .A(n9912), .B(n9913), .Z(n9911) );
  OR U14139 ( .A(n9913), .B(n9912), .Z(n9908) );
  IV U14140 ( .A(n9914), .Z(n9912) );
  XOR U14141 ( .A(n9889), .B(n9915), .Z(N29334) );
  XNOR U14142 ( .A(n9892), .B(n9891), .Z(n9915) );
  XNOR U14143 ( .A(n9903), .B(n9916), .Z(n9891) );
  XOR U14144 ( .A(n9907), .B(n9905), .Z(n9916) );
  XOR U14145 ( .A(n9913), .B(n9917), .Z(n9905) );
  XOR U14146 ( .A(n9910), .B(n9914), .Z(n9917) );
  NAND U14147 ( .A(n9918), .B(n9919), .Z(n9914) );
  NAND U14148 ( .A(n9920), .B(n9921), .Z(n9919) );
  NAND U14149 ( .A(n9922), .B(n9923), .Z(n9918) );
  AND U14150 ( .A(n9924), .B(n9925), .Z(n9910) );
  NAND U14151 ( .A(n9926), .B(n9927), .Z(n9925) );
  NAND U14152 ( .A(n9928), .B(n9929), .Z(n9924) );
  NANDN U14153 ( .A(n9930), .B(n9931), .Z(n9913) );
  NANDN U14154 ( .A(n9932), .B(n9933), .Z(n9907) );
  XNOR U14155 ( .A(n9898), .B(n9934), .Z(n9903) );
  XOR U14156 ( .A(n9896), .B(n9900), .Z(n9934) );
  NAND U14157 ( .A(n9935), .B(n9936), .Z(n9900) );
  NAND U14158 ( .A(n9937), .B(n9938), .Z(n9936) );
  NAND U14159 ( .A(n9939), .B(n9940), .Z(n9935) );
  AND U14160 ( .A(n9941), .B(n9942), .Z(n9896) );
  NAND U14161 ( .A(n9943), .B(n9944), .Z(n9942) );
  NAND U14162 ( .A(n9945), .B(n9946), .Z(n9941) );
  AND U14163 ( .A(n9947), .B(n9948), .Z(n9898) );
  NAND U14164 ( .A(n9949), .B(n9950), .Z(n9892) );
  XNOR U14165 ( .A(n9875), .B(n9951), .Z(n9889) );
  XOR U14166 ( .A(n9879), .B(n9877), .Z(n9951) );
  XOR U14167 ( .A(n9885), .B(n9952), .Z(n9877) );
  XOR U14168 ( .A(n9882), .B(n9886), .Z(n9952) );
  NAND U14169 ( .A(n9953), .B(n9954), .Z(n9886) );
  NAND U14170 ( .A(n9955), .B(n9956), .Z(n9954) );
  NAND U14171 ( .A(n9957), .B(n9958), .Z(n9953) );
  AND U14172 ( .A(n9959), .B(n9960), .Z(n9882) );
  NAND U14173 ( .A(n9961), .B(n9962), .Z(n9960) );
  NAND U14174 ( .A(n9963), .B(n9964), .Z(n9959) );
  NANDN U14175 ( .A(n9965), .B(n9966), .Z(n9885) );
  NANDN U14176 ( .A(n9967), .B(n9968), .Z(n9879) );
  XNOR U14177 ( .A(n9870), .B(n9969), .Z(n9875) );
  XOR U14178 ( .A(n9868), .B(n9872), .Z(n9969) );
  NAND U14179 ( .A(n9970), .B(n9971), .Z(n9872) );
  NAND U14180 ( .A(n9972), .B(n9973), .Z(n9971) );
  NAND U14181 ( .A(n9974), .B(n9975), .Z(n9970) );
  AND U14182 ( .A(n9976), .B(n9977), .Z(n9868) );
  NAND U14183 ( .A(n9978), .B(n9979), .Z(n9977) );
  NAND U14184 ( .A(n9980), .B(n9981), .Z(n9976) );
  AND U14185 ( .A(n9982), .B(n9983), .Z(n9870) );
  XOR U14186 ( .A(n9950), .B(n9949), .Z(N29333) );
  XNOR U14187 ( .A(n9968), .B(n9967), .Z(n9949) );
  XNOR U14188 ( .A(n9982), .B(n9983), .Z(n9967) );
  XOR U14189 ( .A(n9979), .B(n9978), .Z(n9983) );
  XOR U14190 ( .A(y[2811]), .B(x[2811]), .Z(n9978) );
  XOR U14191 ( .A(n9981), .B(n9980), .Z(n9979) );
  XOR U14192 ( .A(y[2813]), .B(x[2813]), .Z(n9980) );
  XOR U14193 ( .A(y[2812]), .B(x[2812]), .Z(n9981) );
  XOR U14194 ( .A(n9973), .B(n9972), .Z(n9982) );
  XOR U14195 ( .A(n9975), .B(n9974), .Z(n9972) );
  XOR U14196 ( .A(y[2810]), .B(x[2810]), .Z(n9974) );
  XOR U14197 ( .A(y[2809]), .B(x[2809]), .Z(n9975) );
  XOR U14198 ( .A(y[2808]), .B(x[2808]), .Z(n9973) );
  XNOR U14199 ( .A(n9966), .B(n9965), .Z(n9968) );
  XNOR U14200 ( .A(n9962), .B(n9961), .Z(n9965) );
  XOR U14201 ( .A(n9964), .B(n9963), .Z(n9961) );
  XOR U14202 ( .A(y[2807]), .B(x[2807]), .Z(n9963) );
  XOR U14203 ( .A(y[2806]), .B(x[2806]), .Z(n9964) );
  XOR U14204 ( .A(y[2805]), .B(x[2805]), .Z(n9962) );
  XOR U14205 ( .A(n9956), .B(n9955), .Z(n9966) );
  XOR U14206 ( .A(n9958), .B(n9957), .Z(n9955) );
  XOR U14207 ( .A(y[2804]), .B(x[2804]), .Z(n9957) );
  XOR U14208 ( .A(y[2803]), .B(x[2803]), .Z(n9958) );
  XOR U14209 ( .A(y[2802]), .B(x[2802]), .Z(n9956) );
  XNOR U14210 ( .A(n9933), .B(n9932), .Z(n9950) );
  XNOR U14211 ( .A(n9947), .B(n9948), .Z(n9932) );
  XOR U14212 ( .A(n9944), .B(n9943), .Z(n9948) );
  XOR U14213 ( .A(y[2799]), .B(x[2799]), .Z(n9943) );
  XOR U14214 ( .A(n9946), .B(n9945), .Z(n9944) );
  XOR U14215 ( .A(y[2801]), .B(x[2801]), .Z(n9945) );
  XOR U14216 ( .A(y[2800]), .B(x[2800]), .Z(n9946) );
  XOR U14217 ( .A(n9938), .B(n9937), .Z(n9947) );
  XOR U14218 ( .A(n9940), .B(n9939), .Z(n9937) );
  XOR U14219 ( .A(y[2798]), .B(x[2798]), .Z(n9939) );
  XOR U14220 ( .A(y[2797]), .B(x[2797]), .Z(n9940) );
  XOR U14221 ( .A(y[2796]), .B(x[2796]), .Z(n9938) );
  XNOR U14222 ( .A(n9931), .B(n9930), .Z(n9933) );
  XNOR U14223 ( .A(n9927), .B(n9926), .Z(n9930) );
  XOR U14224 ( .A(n9929), .B(n9928), .Z(n9926) );
  XOR U14225 ( .A(y[2795]), .B(x[2795]), .Z(n9928) );
  XOR U14226 ( .A(y[2794]), .B(x[2794]), .Z(n9929) );
  XOR U14227 ( .A(y[2793]), .B(x[2793]), .Z(n9927) );
  XOR U14228 ( .A(n9921), .B(n9920), .Z(n9931) );
  XOR U14229 ( .A(n9923), .B(n9922), .Z(n9920) );
  XOR U14230 ( .A(y[2792]), .B(x[2792]), .Z(n9922) );
  XOR U14231 ( .A(y[2791]), .B(x[2791]), .Z(n9923) );
  XOR U14232 ( .A(y[2790]), .B(x[2790]), .Z(n9921) );
  NAND U14233 ( .A(n9984), .B(n9985), .Z(N29325) );
  NAND U14234 ( .A(n9986), .B(n9987), .Z(n9985) );
  NANDN U14235 ( .A(n9988), .B(n9989), .Z(n9987) );
  NANDN U14236 ( .A(n9989), .B(n9988), .Z(n9984) );
  XOR U14237 ( .A(n9988), .B(n9990), .Z(N29324) );
  XNOR U14238 ( .A(n9986), .B(n9989), .Z(n9990) );
  NAND U14239 ( .A(n9991), .B(n9992), .Z(n9989) );
  NAND U14240 ( .A(n9993), .B(n9994), .Z(n9992) );
  NANDN U14241 ( .A(n9995), .B(n9996), .Z(n9994) );
  NANDN U14242 ( .A(n9996), .B(n9995), .Z(n9991) );
  AND U14243 ( .A(n9997), .B(n9998), .Z(n9986) );
  NAND U14244 ( .A(n9999), .B(n10000), .Z(n9998) );
  OR U14245 ( .A(n10001), .B(n10002), .Z(n10000) );
  NAND U14246 ( .A(n10002), .B(n10001), .Z(n9997) );
  IV U14247 ( .A(n10003), .Z(n10002) );
  AND U14248 ( .A(n10004), .B(n10005), .Z(n9988) );
  NAND U14249 ( .A(n10006), .B(n10007), .Z(n10005) );
  NANDN U14250 ( .A(n10008), .B(n10009), .Z(n10007) );
  NANDN U14251 ( .A(n10009), .B(n10008), .Z(n10004) );
  XOR U14252 ( .A(n10001), .B(n10010), .Z(N29323) );
  XOR U14253 ( .A(n9999), .B(n10003), .Z(n10010) );
  XNOR U14254 ( .A(n9996), .B(n10011), .Z(n10003) );
  XNOR U14255 ( .A(n9993), .B(n9995), .Z(n10011) );
  AND U14256 ( .A(n10012), .B(n10013), .Z(n9995) );
  NANDN U14257 ( .A(n10014), .B(n10015), .Z(n10013) );
  NANDN U14258 ( .A(n10016), .B(n10017), .Z(n10015) );
  IV U14259 ( .A(n10018), .Z(n10017) );
  NAND U14260 ( .A(n10018), .B(n10016), .Z(n10012) );
  AND U14261 ( .A(n10019), .B(n10020), .Z(n9993) );
  NAND U14262 ( .A(n10021), .B(n10022), .Z(n10020) );
  OR U14263 ( .A(n10023), .B(n10024), .Z(n10022) );
  NAND U14264 ( .A(n10024), .B(n10023), .Z(n10019) );
  IV U14265 ( .A(n10025), .Z(n10024) );
  NAND U14266 ( .A(n10026), .B(n10027), .Z(n9996) );
  NANDN U14267 ( .A(n10028), .B(n10029), .Z(n10027) );
  NAND U14268 ( .A(n10030), .B(n10031), .Z(n10029) );
  OR U14269 ( .A(n10031), .B(n10030), .Z(n10026) );
  IV U14270 ( .A(n10032), .Z(n10030) );
  AND U14271 ( .A(n10033), .B(n10034), .Z(n9999) );
  NAND U14272 ( .A(n10035), .B(n10036), .Z(n10034) );
  NANDN U14273 ( .A(n10037), .B(n10038), .Z(n10036) );
  NANDN U14274 ( .A(n10038), .B(n10037), .Z(n10033) );
  XOR U14275 ( .A(n10009), .B(n10039), .Z(n10001) );
  XNOR U14276 ( .A(n10006), .B(n10008), .Z(n10039) );
  AND U14277 ( .A(n10040), .B(n10041), .Z(n10008) );
  NANDN U14278 ( .A(n10042), .B(n10043), .Z(n10041) );
  NANDN U14279 ( .A(n10044), .B(n10045), .Z(n10043) );
  IV U14280 ( .A(n10046), .Z(n10045) );
  NAND U14281 ( .A(n10046), .B(n10044), .Z(n10040) );
  AND U14282 ( .A(n10047), .B(n10048), .Z(n10006) );
  NAND U14283 ( .A(n10049), .B(n10050), .Z(n10048) );
  OR U14284 ( .A(n10051), .B(n10052), .Z(n10050) );
  NAND U14285 ( .A(n10052), .B(n10051), .Z(n10047) );
  IV U14286 ( .A(n10053), .Z(n10052) );
  NAND U14287 ( .A(n10054), .B(n10055), .Z(n10009) );
  NANDN U14288 ( .A(n10056), .B(n10057), .Z(n10055) );
  NAND U14289 ( .A(n10058), .B(n10059), .Z(n10057) );
  OR U14290 ( .A(n10059), .B(n10058), .Z(n10054) );
  IV U14291 ( .A(n10060), .Z(n10058) );
  XOR U14292 ( .A(n10035), .B(n10061), .Z(N29322) );
  XNOR U14293 ( .A(n10038), .B(n10037), .Z(n10061) );
  XNOR U14294 ( .A(n10049), .B(n10062), .Z(n10037) );
  XOR U14295 ( .A(n10053), .B(n10051), .Z(n10062) );
  XOR U14296 ( .A(n10059), .B(n10063), .Z(n10051) );
  XOR U14297 ( .A(n10056), .B(n10060), .Z(n10063) );
  NAND U14298 ( .A(n10064), .B(n10065), .Z(n10060) );
  NAND U14299 ( .A(n10066), .B(n10067), .Z(n10065) );
  NAND U14300 ( .A(n10068), .B(n10069), .Z(n10064) );
  AND U14301 ( .A(n10070), .B(n10071), .Z(n10056) );
  NAND U14302 ( .A(n10072), .B(n10073), .Z(n10071) );
  NAND U14303 ( .A(n10074), .B(n10075), .Z(n10070) );
  NANDN U14304 ( .A(n10076), .B(n10077), .Z(n10059) );
  NANDN U14305 ( .A(n10078), .B(n10079), .Z(n10053) );
  XNOR U14306 ( .A(n10044), .B(n10080), .Z(n10049) );
  XOR U14307 ( .A(n10042), .B(n10046), .Z(n10080) );
  NAND U14308 ( .A(n10081), .B(n10082), .Z(n10046) );
  NAND U14309 ( .A(n10083), .B(n10084), .Z(n10082) );
  NAND U14310 ( .A(n10085), .B(n10086), .Z(n10081) );
  AND U14311 ( .A(n10087), .B(n10088), .Z(n10042) );
  NAND U14312 ( .A(n10089), .B(n10090), .Z(n10088) );
  NAND U14313 ( .A(n10091), .B(n10092), .Z(n10087) );
  AND U14314 ( .A(n10093), .B(n10094), .Z(n10044) );
  NAND U14315 ( .A(n10095), .B(n10096), .Z(n10038) );
  XNOR U14316 ( .A(n10021), .B(n10097), .Z(n10035) );
  XOR U14317 ( .A(n10025), .B(n10023), .Z(n10097) );
  XOR U14318 ( .A(n10031), .B(n10098), .Z(n10023) );
  XOR U14319 ( .A(n10028), .B(n10032), .Z(n10098) );
  NAND U14320 ( .A(n10099), .B(n10100), .Z(n10032) );
  NAND U14321 ( .A(n10101), .B(n10102), .Z(n10100) );
  NAND U14322 ( .A(n10103), .B(n10104), .Z(n10099) );
  AND U14323 ( .A(n10105), .B(n10106), .Z(n10028) );
  NAND U14324 ( .A(n10107), .B(n10108), .Z(n10106) );
  NAND U14325 ( .A(n10109), .B(n10110), .Z(n10105) );
  NANDN U14326 ( .A(n10111), .B(n10112), .Z(n10031) );
  NANDN U14327 ( .A(n10113), .B(n10114), .Z(n10025) );
  XNOR U14328 ( .A(n10016), .B(n10115), .Z(n10021) );
  XOR U14329 ( .A(n10014), .B(n10018), .Z(n10115) );
  NAND U14330 ( .A(n10116), .B(n10117), .Z(n10018) );
  NAND U14331 ( .A(n10118), .B(n10119), .Z(n10117) );
  NAND U14332 ( .A(n10120), .B(n10121), .Z(n10116) );
  AND U14333 ( .A(n10122), .B(n10123), .Z(n10014) );
  NAND U14334 ( .A(n10124), .B(n10125), .Z(n10123) );
  NAND U14335 ( .A(n10126), .B(n10127), .Z(n10122) );
  AND U14336 ( .A(n10128), .B(n10129), .Z(n10016) );
  XOR U14337 ( .A(n10096), .B(n10095), .Z(N29321) );
  XNOR U14338 ( .A(n10114), .B(n10113), .Z(n10095) );
  XNOR U14339 ( .A(n10128), .B(n10129), .Z(n10113) );
  XOR U14340 ( .A(n10125), .B(n10124), .Z(n10129) );
  XOR U14341 ( .A(y[2787]), .B(x[2787]), .Z(n10124) );
  XOR U14342 ( .A(n10127), .B(n10126), .Z(n10125) );
  XOR U14343 ( .A(y[2789]), .B(x[2789]), .Z(n10126) );
  XOR U14344 ( .A(y[2788]), .B(x[2788]), .Z(n10127) );
  XOR U14345 ( .A(n10119), .B(n10118), .Z(n10128) );
  XOR U14346 ( .A(n10121), .B(n10120), .Z(n10118) );
  XOR U14347 ( .A(y[2786]), .B(x[2786]), .Z(n10120) );
  XOR U14348 ( .A(y[2785]), .B(x[2785]), .Z(n10121) );
  XOR U14349 ( .A(y[2784]), .B(x[2784]), .Z(n10119) );
  XNOR U14350 ( .A(n10112), .B(n10111), .Z(n10114) );
  XNOR U14351 ( .A(n10108), .B(n10107), .Z(n10111) );
  XOR U14352 ( .A(n10110), .B(n10109), .Z(n10107) );
  XOR U14353 ( .A(y[2783]), .B(x[2783]), .Z(n10109) );
  XOR U14354 ( .A(y[2782]), .B(x[2782]), .Z(n10110) );
  XOR U14355 ( .A(y[2781]), .B(x[2781]), .Z(n10108) );
  XOR U14356 ( .A(n10102), .B(n10101), .Z(n10112) );
  XOR U14357 ( .A(n10104), .B(n10103), .Z(n10101) );
  XOR U14358 ( .A(y[2780]), .B(x[2780]), .Z(n10103) );
  XOR U14359 ( .A(y[2779]), .B(x[2779]), .Z(n10104) );
  XOR U14360 ( .A(y[2778]), .B(x[2778]), .Z(n10102) );
  XNOR U14361 ( .A(n10079), .B(n10078), .Z(n10096) );
  XNOR U14362 ( .A(n10093), .B(n10094), .Z(n10078) );
  XOR U14363 ( .A(n10090), .B(n10089), .Z(n10094) );
  XOR U14364 ( .A(y[2775]), .B(x[2775]), .Z(n10089) );
  XOR U14365 ( .A(n10092), .B(n10091), .Z(n10090) );
  XOR U14366 ( .A(y[2777]), .B(x[2777]), .Z(n10091) );
  XOR U14367 ( .A(y[2776]), .B(x[2776]), .Z(n10092) );
  XOR U14368 ( .A(n10084), .B(n10083), .Z(n10093) );
  XOR U14369 ( .A(n10086), .B(n10085), .Z(n10083) );
  XOR U14370 ( .A(y[2774]), .B(x[2774]), .Z(n10085) );
  XOR U14371 ( .A(y[2773]), .B(x[2773]), .Z(n10086) );
  XOR U14372 ( .A(y[2772]), .B(x[2772]), .Z(n10084) );
  XNOR U14373 ( .A(n10077), .B(n10076), .Z(n10079) );
  XNOR U14374 ( .A(n10073), .B(n10072), .Z(n10076) );
  XOR U14375 ( .A(n10075), .B(n10074), .Z(n10072) );
  XOR U14376 ( .A(y[2771]), .B(x[2771]), .Z(n10074) );
  XOR U14377 ( .A(y[2770]), .B(x[2770]), .Z(n10075) );
  XOR U14378 ( .A(y[2769]), .B(x[2769]), .Z(n10073) );
  XOR U14379 ( .A(n10067), .B(n10066), .Z(n10077) );
  XOR U14380 ( .A(n10069), .B(n10068), .Z(n10066) );
  XOR U14381 ( .A(y[2768]), .B(x[2768]), .Z(n10068) );
  XOR U14382 ( .A(y[2767]), .B(x[2767]), .Z(n10069) );
  XOR U14383 ( .A(y[2766]), .B(x[2766]), .Z(n10067) );
  NAND U14384 ( .A(n10130), .B(n10131), .Z(N29313) );
  NAND U14385 ( .A(n10132), .B(n10133), .Z(n10131) );
  NANDN U14386 ( .A(n10134), .B(n10135), .Z(n10133) );
  NANDN U14387 ( .A(n10135), .B(n10134), .Z(n10130) );
  XOR U14388 ( .A(n10134), .B(n10136), .Z(N29312) );
  XNOR U14389 ( .A(n10132), .B(n10135), .Z(n10136) );
  NAND U14390 ( .A(n10137), .B(n10138), .Z(n10135) );
  NAND U14391 ( .A(n10139), .B(n10140), .Z(n10138) );
  NANDN U14392 ( .A(n10141), .B(n10142), .Z(n10140) );
  NANDN U14393 ( .A(n10142), .B(n10141), .Z(n10137) );
  AND U14394 ( .A(n10143), .B(n10144), .Z(n10132) );
  NAND U14395 ( .A(n10145), .B(n10146), .Z(n10144) );
  OR U14396 ( .A(n10147), .B(n10148), .Z(n10146) );
  NAND U14397 ( .A(n10148), .B(n10147), .Z(n10143) );
  IV U14398 ( .A(n10149), .Z(n10148) );
  AND U14399 ( .A(n10150), .B(n10151), .Z(n10134) );
  NAND U14400 ( .A(n10152), .B(n10153), .Z(n10151) );
  NANDN U14401 ( .A(n10154), .B(n10155), .Z(n10153) );
  NANDN U14402 ( .A(n10155), .B(n10154), .Z(n10150) );
  XOR U14403 ( .A(n10147), .B(n10156), .Z(N29311) );
  XOR U14404 ( .A(n10145), .B(n10149), .Z(n10156) );
  XNOR U14405 ( .A(n10142), .B(n10157), .Z(n10149) );
  XNOR U14406 ( .A(n10139), .B(n10141), .Z(n10157) );
  AND U14407 ( .A(n10158), .B(n10159), .Z(n10141) );
  NANDN U14408 ( .A(n10160), .B(n10161), .Z(n10159) );
  NANDN U14409 ( .A(n10162), .B(n10163), .Z(n10161) );
  IV U14410 ( .A(n10164), .Z(n10163) );
  NAND U14411 ( .A(n10164), .B(n10162), .Z(n10158) );
  AND U14412 ( .A(n10165), .B(n10166), .Z(n10139) );
  NAND U14413 ( .A(n10167), .B(n10168), .Z(n10166) );
  OR U14414 ( .A(n10169), .B(n10170), .Z(n10168) );
  NAND U14415 ( .A(n10170), .B(n10169), .Z(n10165) );
  IV U14416 ( .A(n10171), .Z(n10170) );
  NAND U14417 ( .A(n10172), .B(n10173), .Z(n10142) );
  NANDN U14418 ( .A(n10174), .B(n10175), .Z(n10173) );
  NAND U14419 ( .A(n10176), .B(n10177), .Z(n10175) );
  OR U14420 ( .A(n10177), .B(n10176), .Z(n10172) );
  IV U14421 ( .A(n10178), .Z(n10176) );
  AND U14422 ( .A(n10179), .B(n10180), .Z(n10145) );
  NAND U14423 ( .A(n10181), .B(n10182), .Z(n10180) );
  NANDN U14424 ( .A(n10183), .B(n10184), .Z(n10182) );
  NANDN U14425 ( .A(n10184), .B(n10183), .Z(n10179) );
  XOR U14426 ( .A(n10155), .B(n10185), .Z(n10147) );
  XNOR U14427 ( .A(n10152), .B(n10154), .Z(n10185) );
  AND U14428 ( .A(n10186), .B(n10187), .Z(n10154) );
  NANDN U14429 ( .A(n10188), .B(n10189), .Z(n10187) );
  NANDN U14430 ( .A(n10190), .B(n10191), .Z(n10189) );
  IV U14431 ( .A(n10192), .Z(n10191) );
  NAND U14432 ( .A(n10192), .B(n10190), .Z(n10186) );
  AND U14433 ( .A(n10193), .B(n10194), .Z(n10152) );
  NAND U14434 ( .A(n10195), .B(n10196), .Z(n10194) );
  OR U14435 ( .A(n10197), .B(n10198), .Z(n10196) );
  NAND U14436 ( .A(n10198), .B(n10197), .Z(n10193) );
  IV U14437 ( .A(n10199), .Z(n10198) );
  NAND U14438 ( .A(n10200), .B(n10201), .Z(n10155) );
  NANDN U14439 ( .A(n10202), .B(n10203), .Z(n10201) );
  NAND U14440 ( .A(n10204), .B(n10205), .Z(n10203) );
  OR U14441 ( .A(n10205), .B(n10204), .Z(n10200) );
  IV U14442 ( .A(n10206), .Z(n10204) );
  XOR U14443 ( .A(n10181), .B(n10207), .Z(N29310) );
  XNOR U14444 ( .A(n10184), .B(n10183), .Z(n10207) );
  XNOR U14445 ( .A(n10195), .B(n10208), .Z(n10183) );
  XOR U14446 ( .A(n10199), .B(n10197), .Z(n10208) );
  XOR U14447 ( .A(n10205), .B(n10209), .Z(n10197) );
  XOR U14448 ( .A(n10202), .B(n10206), .Z(n10209) );
  NAND U14449 ( .A(n10210), .B(n10211), .Z(n10206) );
  NAND U14450 ( .A(n10212), .B(n10213), .Z(n10211) );
  NAND U14451 ( .A(n10214), .B(n10215), .Z(n10210) );
  AND U14452 ( .A(n10216), .B(n10217), .Z(n10202) );
  NAND U14453 ( .A(n10218), .B(n10219), .Z(n10217) );
  NAND U14454 ( .A(n10220), .B(n10221), .Z(n10216) );
  NANDN U14455 ( .A(n10222), .B(n10223), .Z(n10205) );
  NANDN U14456 ( .A(n10224), .B(n10225), .Z(n10199) );
  XNOR U14457 ( .A(n10190), .B(n10226), .Z(n10195) );
  XOR U14458 ( .A(n10188), .B(n10192), .Z(n10226) );
  NAND U14459 ( .A(n10227), .B(n10228), .Z(n10192) );
  NAND U14460 ( .A(n10229), .B(n10230), .Z(n10228) );
  NAND U14461 ( .A(n10231), .B(n10232), .Z(n10227) );
  AND U14462 ( .A(n10233), .B(n10234), .Z(n10188) );
  NAND U14463 ( .A(n10235), .B(n10236), .Z(n10234) );
  NAND U14464 ( .A(n10237), .B(n10238), .Z(n10233) );
  AND U14465 ( .A(n10239), .B(n10240), .Z(n10190) );
  NAND U14466 ( .A(n10241), .B(n10242), .Z(n10184) );
  XNOR U14467 ( .A(n10167), .B(n10243), .Z(n10181) );
  XOR U14468 ( .A(n10171), .B(n10169), .Z(n10243) );
  XOR U14469 ( .A(n10177), .B(n10244), .Z(n10169) );
  XOR U14470 ( .A(n10174), .B(n10178), .Z(n10244) );
  NAND U14471 ( .A(n10245), .B(n10246), .Z(n10178) );
  NAND U14472 ( .A(n10247), .B(n10248), .Z(n10246) );
  NAND U14473 ( .A(n10249), .B(n10250), .Z(n10245) );
  AND U14474 ( .A(n10251), .B(n10252), .Z(n10174) );
  NAND U14475 ( .A(n10253), .B(n10254), .Z(n10252) );
  NAND U14476 ( .A(n10255), .B(n10256), .Z(n10251) );
  NANDN U14477 ( .A(n10257), .B(n10258), .Z(n10177) );
  NANDN U14478 ( .A(n10259), .B(n10260), .Z(n10171) );
  XNOR U14479 ( .A(n10162), .B(n10261), .Z(n10167) );
  XOR U14480 ( .A(n10160), .B(n10164), .Z(n10261) );
  NAND U14481 ( .A(n10262), .B(n10263), .Z(n10164) );
  NAND U14482 ( .A(n10264), .B(n10265), .Z(n10263) );
  NAND U14483 ( .A(n10266), .B(n10267), .Z(n10262) );
  AND U14484 ( .A(n10268), .B(n10269), .Z(n10160) );
  NAND U14485 ( .A(n10270), .B(n10271), .Z(n10269) );
  NAND U14486 ( .A(n10272), .B(n10273), .Z(n10268) );
  AND U14487 ( .A(n10274), .B(n10275), .Z(n10162) );
  XOR U14488 ( .A(n10242), .B(n10241), .Z(N29309) );
  XNOR U14489 ( .A(n10260), .B(n10259), .Z(n10241) );
  XNOR U14490 ( .A(n10274), .B(n10275), .Z(n10259) );
  XOR U14491 ( .A(n10271), .B(n10270), .Z(n10275) );
  XOR U14492 ( .A(y[2763]), .B(x[2763]), .Z(n10270) );
  XOR U14493 ( .A(n10273), .B(n10272), .Z(n10271) );
  XOR U14494 ( .A(y[2765]), .B(x[2765]), .Z(n10272) );
  XOR U14495 ( .A(y[2764]), .B(x[2764]), .Z(n10273) );
  XOR U14496 ( .A(n10265), .B(n10264), .Z(n10274) );
  XOR U14497 ( .A(n10267), .B(n10266), .Z(n10264) );
  XOR U14498 ( .A(y[2762]), .B(x[2762]), .Z(n10266) );
  XOR U14499 ( .A(y[2761]), .B(x[2761]), .Z(n10267) );
  XOR U14500 ( .A(y[2760]), .B(x[2760]), .Z(n10265) );
  XNOR U14501 ( .A(n10258), .B(n10257), .Z(n10260) );
  XNOR U14502 ( .A(n10254), .B(n10253), .Z(n10257) );
  XOR U14503 ( .A(n10256), .B(n10255), .Z(n10253) );
  XOR U14504 ( .A(y[2759]), .B(x[2759]), .Z(n10255) );
  XOR U14505 ( .A(y[2758]), .B(x[2758]), .Z(n10256) );
  XOR U14506 ( .A(y[2757]), .B(x[2757]), .Z(n10254) );
  XOR U14507 ( .A(n10248), .B(n10247), .Z(n10258) );
  XOR U14508 ( .A(n10250), .B(n10249), .Z(n10247) );
  XOR U14509 ( .A(y[2756]), .B(x[2756]), .Z(n10249) );
  XOR U14510 ( .A(y[2755]), .B(x[2755]), .Z(n10250) );
  XOR U14511 ( .A(y[2754]), .B(x[2754]), .Z(n10248) );
  XNOR U14512 ( .A(n10225), .B(n10224), .Z(n10242) );
  XNOR U14513 ( .A(n10239), .B(n10240), .Z(n10224) );
  XOR U14514 ( .A(n10236), .B(n10235), .Z(n10240) );
  XOR U14515 ( .A(y[2751]), .B(x[2751]), .Z(n10235) );
  XOR U14516 ( .A(n10238), .B(n10237), .Z(n10236) );
  XOR U14517 ( .A(y[2753]), .B(x[2753]), .Z(n10237) );
  XOR U14518 ( .A(y[2752]), .B(x[2752]), .Z(n10238) );
  XOR U14519 ( .A(n10230), .B(n10229), .Z(n10239) );
  XOR U14520 ( .A(n10232), .B(n10231), .Z(n10229) );
  XOR U14521 ( .A(y[2750]), .B(x[2750]), .Z(n10231) );
  XOR U14522 ( .A(y[2749]), .B(x[2749]), .Z(n10232) );
  XOR U14523 ( .A(y[2748]), .B(x[2748]), .Z(n10230) );
  XNOR U14524 ( .A(n10223), .B(n10222), .Z(n10225) );
  XNOR U14525 ( .A(n10219), .B(n10218), .Z(n10222) );
  XOR U14526 ( .A(n10221), .B(n10220), .Z(n10218) );
  XOR U14527 ( .A(y[2747]), .B(x[2747]), .Z(n10220) );
  XOR U14528 ( .A(y[2746]), .B(x[2746]), .Z(n10221) );
  XOR U14529 ( .A(y[2745]), .B(x[2745]), .Z(n10219) );
  XOR U14530 ( .A(n10213), .B(n10212), .Z(n10223) );
  XOR U14531 ( .A(n10215), .B(n10214), .Z(n10212) );
  XOR U14532 ( .A(y[2744]), .B(x[2744]), .Z(n10214) );
  XOR U14533 ( .A(y[2743]), .B(x[2743]), .Z(n10215) );
  XOR U14534 ( .A(y[2742]), .B(x[2742]), .Z(n10213) );
  NAND U14535 ( .A(n10276), .B(n10277), .Z(N29301) );
  NAND U14536 ( .A(n10278), .B(n10279), .Z(n10277) );
  NANDN U14537 ( .A(n10280), .B(n10281), .Z(n10279) );
  NANDN U14538 ( .A(n10281), .B(n10280), .Z(n10276) );
  XOR U14539 ( .A(n10280), .B(n10282), .Z(N29300) );
  XNOR U14540 ( .A(n10278), .B(n10281), .Z(n10282) );
  NAND U14541 ( .A(n10283), .B(n10284), .Z(n10281) );
  NAND U14542 ( .A(n10285), .B(n10286), .Z(n10284) );
  NANDN U14543 ( .A(n10287), .B(n10288), .Z(n10286) );
  NANDN U14544 ( .A(n10288), .B(n10287), .Z(n10283) );
  AND U14545 ( .A(n10289), .B(n10290), .Z(n10278) );
  NAND U14546 ( .A(n10291), .B(n10292), .Z(n10290) );
  OR U14547 ( .A(n10293), .B(n10294), .Z(n10292) );
  NAND U14548 ( .A(n10294), .B(n10293), .Z(n10289) );
  IV U14549 ( .A(n10295), .Z(n10294) );
  AND U14550 ( .A(n10296), .B(n10297), .Z(n10280) );
  NAND U14551 ( .A(n10298), .B(n10299), .Z(n10297) );
  NANDN U14552 ( .A(n10300), .B(n10301), .Z(n10299) );
  NANDN U14553 ( .A(n10301), .B(n10300), .Z(n10296) );
  XOR U14554 ( .A(n10293), .B(n10302), .Z(N29299) );
  XOR U14555 ( .A(n10291), .B(n10295), .Z(n10302) );
  XNOR U14556 ( .A(n10288), .B(n10303), .Z(n10295) );
  XNOR U14557 ( .A(n10285), .B(n10287), .Z(n10303) );
  AND U14558 ( .A(n10304), .B(n10305), .Z(n10287) );
  NANDN U14559 ( .A(n10306), .B(n10307), .Z(n10305) );
  NANDN U14560 ( .A(n10308), .B(n10309), .Z(n10307) );
  IV U14561 ( .A(n10310), .Z(n10309) );
  NAND U14562 ( .A(n10310), .B(n10308), .Z(n10304) );
  AND U14563 ( .A(n10311), .B(n10312), .Z(n10285) );
  NAND U14564 ( .A(n10313), .B(n10314), .Z(n10312) );
  OR U14565 ( .A(n10315), .B(n10316), .Z(n10314) );
  NAND U14566 ( .A(n10316), .B(n10315), .Z(n10311) );
  IV U14567 ( .A(n10317), .Z(n10316) );
  NAND U14568 ( .A(n10318), .B(n10319), .Z(n10288) );
  NANDN U14569 ( .A(n10320), .B(n10321), .Z(n10319) );
  NAND U14570 ( .A(n10322), .B(n10323), .Z(n10321) );
  OR U14571 ( .A(n10323), .B(n10322), .Z(n10318) );
  IV U14572 ( .A(n10324), .Z(n10322) );
  AND U14573 ( .A(n10325), .B(n10326), .Z(n10291) );
  NAND U14574 ( .A(n10327), .B(n10328), .Z(n10326) );
  NANDN U14575 ( .A(n10329), .B(n10330), .Z(n10328) );
  NANDN U14576 ( .A(n10330), .B(n10329), .Z(n10325) );
  XOR U14577 ( .A(n10301), .B(n10331), .Z(n10293) );
  XNOR U14578 ( .A(n10298), .B(n10300), .Z(n10331) );
  AND U14579 ( .A(n10332), .B(n10333), .Z(n10300) );
  NANDN U14580 ( .A(n10334), .B(n10335), .Z(n10333) );
  NANDN U14581 ( .A(n10336), .B(n10337), .Z(n10335) );
  IV U14582 ( .A(n10338), .Z(n10337) );
  NAND U14583 ( .A(n10338), .B(n10336), .Z(n10332) );
  AND U14584 ( .A(n10339), .B(n10340), .Z(n10298) );
  NAND U14585 ( .A(n10341), .B(n10342), .Z(n10340) );
  OR U14586 ( .A(n10343), .B(n10344), .Z(n10342) );
  NAND U14587 ( .A(n10344), .B(n10343), .Z(n10339) );
  IV U14588 ( .A(n10345), .Z(n10344) );
  NAND U14589 ( .A(n10346), .B(n10347), .Z(n10301) );
  NANDN U14590 ( .A(n10348), .B(n10349), .Z(n10347) );
  NAND U14591 ( .A(n10350), .B(n10351), .Z(n10349) );
  OR U14592 ( .A(n10351), .B(n10350), .Z(n10346) );
  IV U14593 ( .A(n10352), .Z(n10350) );
  XOR U14594 ( .A(n10327), .B(n10353), .Z(N29298) );
  XNOR U14595 ( .A(n10330), .B(n10329), .Z(n10353) );
  XNOR U14596 ( .A(n10341), .B(n10354), .Z(n10329) );
  XOR U14597 ( .A(n10345), .B(n10343), .Z(n10354) );
  XOR U14598 ( .A(n10351), .B(n10355), .Z(n10343) );
  XOR U14599 ( .A(n10348), .B(n10352), .Z(n10355) );
  NAND U14600 ( .A(n10356), .B(n10357), .Z(n10352) );
  NAND U14601 ( .A(n10358), .B(n10359), .Z(n10357) );
  NAND U14602 ( .A(n10360), .B(n10361), .Z(n10356) );
  AND U14603 ( .A(n10362), .B(n10363), .Z(n10348) );
  NAND U14604 ( .A(n10364), .B(n10365), .Z(n10363) );
  NAND U14605 ( .A(n10366), .B(n10367), .Z(n10362) );
  NANDN U14606 ( .A(n10368), .B(n10369), .Z(n10351) );
  NANDN U14607 ( .A(n10370), .B(n10371), .Z(n10345) );
  XNOR U14608 ( .A(n10336), .B(n10372), .Z(n10341) );
  XOR U14609 ( .A(n10334), .B(n10338), .Z(n10372) );
  NAND U14610 ( .A(n10373), .B(n10374), .Z(n10338) );
  NAND U14611 ( .A(n10375), .B(n10376), .Z(n10374) );
  NAND U14612 ( .A(n10377), .B(n10378), .Z(n10373) );
  AND U14613 ( .A(n10379), .B(n10380), .Z(n10334) );
  NAND U14614 ( .A(n10381), .B(n10382), .Z(n10380) );
  NAND U14615 ( .A(n10383), .B(n10384), .Z(n10379) );
  AND U14616 ( .A(n10385), .B(n10386), .Z(n10336) );
  NAND U14617 ( .A(n10387), .B(n10388), .Z(n10330) );
  XNOR U14618 ( .A(n10313), .B(n10389), .Z(n10327) );
  XOR U14619 ( .A(n10317), .B(n10315), .Z(n10389) );
  XOR U14620 ( .A(n10323), .B(n10390), .Z(n10315) );
  XOR U14621 ( .A(n10320), .B(n10324), .Z(n10390) );
  NAND U14622 ( .A(n10391), .B(n10392), .Z(n10324) );
  NAND U14623 ( .A(n10393), .B(n10394), .Z(n10392) );
  NAND U14624 ( .A(n10395), .B(n10396), .Z(n10391) );
  AND U14625 ( .A(n10397), .B(n10398), .Z(n10320) );
  NAND U14626 ( .A(n10399), .B(n10400), .Z(n10398) );
  NAND U14627 ( .A(n10401), .B(n10402), .Z(n10397) );
  NANDN U14628 ( .A(n10403), .B(n10404), .Z(n10323) );
  NANDN U14629 ( .A(n10405), .B(n10406), .Z(n10317) );
  XNOR U14630 ( .A(n10308), .B(n10407), .Z(n10313) );
  XOR U14631 ( .A(n10306), .B(n10310), .Z(n10407) );
  NAND U14632 ( .A(n10408), .B(n10409), .Z(n10310) );
  NAND U14633 ( .A(n10410), .B(n10411), .Z(n10409) );
  NAND U14634 ( .A(n10412), .B(n10413), .Z(n10408) );
  AND U14635 ( .A(n10414), .B(n10415), .Z(n10306) );
  NAND U14636 ( .A(n10416), .B(n10417), .Z(n10415) );
  NAND U14637 ( .A(n10418), .B(n10419), .Z(n10414) );
  AND U14638 ( .A(n10420), .B(n10421), .Z(n10308) );
  XOR U14639 ( .A(n10388), .B(n10387), .Z(N29297) );
  XNOR U14640 ( .A(n10406), .B(n10405), .Z(n10387) );
  XNOR U14641 ( .A(n10420), .B(n10421), .Z(n10405) );
  XOR U14642 ( .A(n10417), .B(n10416), .Z(n10421) );
  XOR U14643 ( .A(y[2739]), .B(x[2739]), .Z(n10416) );
  XOR U14644 ( .A(n10419), .B(n10418), .Z(n10417) );
  XOR U14645 ( .A(y[2741]), .B(x[2741]), .Z(n10418) );
  XOR U14646 ( .A(y[2740]), .B(x[2740]), .Z(n10419) );
  XOR U14647 ( .A(n10411), .B(n10410), .Z(n10420) );
  XOR U14648 ( .A(n10413), .B(n10412), .Z(n10410) );
  XOR U14649 ( .A(y[2738]), .B(x[2738]), .Z(n10412) );
  XOR U14650 ( .A(y[2737]), .B(x[2737]), .Z(n10413) );
  XOR U14651 ( .A(y[2736]), .B(x[2736]), .Z(n10411) );
  XNOR U14652 ( .A(n10404), .B(n10403), .Z(n10406) );
  XNOR U14653 ( .A(n10400), .B(n10399), .Z(n10403) );
  XOR U14654 ( .A(n10402), .B(n10401), .Z(n10399) );
  XOR U14655 ( .A(y[2735]), .B(x[2735]), .Z(n10401) );
  XOR U14656 ( .A(y[2734]), .B(x[2734]), .Z(n10402) );
  XOR U14657 ( .A(y[2733]), .B(x[2733]), .Z(n10400) );
  XOR U14658 ( .A(n10394), .B(n10393), .Z(n10404) );
  XOR U14659 ( .A(n10396), .B(n10395), .Z(n10393) );
  XOR U14660 ( .A(y[2732]), .B(x[2732]), .Z(n10395) );
  XOR U14661 ( .A(y[2731]), .B(x[2731]), .Z(n10396) );
  XOR U14662 ( .A(y[2730]), .B(x[2730]), .Z(n10394) );
  XNOR U14663 ( .A(n10371), .B(n10370), .Z(n10388) );
  XNOR U14664 ( .A(n10385), .B(n10386), .Z(n10370) );
  XOR U14665 ( .A(n10382), .B(n10381), .Z(n10386) );
  XOR U14666 ( .A(y[2727]), .B(x[2727]), .Z(n10381) );
  XOR U14667 ( .A(n10384), .B(n10383), .Z(n10382) );
  XOR U14668 ( .A(y[2729]), .B(x[2729]), .Z(n10383) );
  XOR U14669 ( .A(y[2728]), .B(x[2728]), .Z(n10384) );
  XOR U14670 ( .A(n10376), .B(n10375), .Z(n10385) );
  XOR U14671 ( .A(n10378), .B(n10377), .Z(n10375) );
  XOR U14672 ( .A(y[2726]), .B(x[2726]), .Z(n10377) );
  XOR U14673 ( .A(y[2725]), .B(x[2725]), .Z(n10378) );
  XOR U14674 ( .A(y[2724]), .B(x[2724]), .Z(n10376) );
  XNOR U14675 ( .A(n10369), .B(n10368), .Z(n10371) );
  XNOR U14676 ( .A(n10365), .B(n10364), .Z(n10368) );
  XOR U14677 ( .A(n10367), .B(n10366), .Z(n10364) );
  XOR U14678 ( .A(y[2723]), .B(x[2723]), .Z(n10366) );
  XOR U14679 ( .A(y[2722]), .B(x[2722]), .Z(n10367) );
  XOR U14680 ( .A(y[2721]), .B(x[2721]), .Z(n10365) );
  XOR U14681 ( .A(n10359), .B(n10358), .Z(n10369) );
  XOR U14682 ( .A(n10361), .B(n10360), .Z(n10358) );
  XOR U14683 ( .A(y[2720]), .B(x[2720]), .Z(n10360) );
  XOR U14684 ( .A(y[2719]), .B(x[2719]), .Z(n10361) );
  XOR U14685 ( .A(y[2718]), .B(x[2718]), .Z(n10359) );
  NAND U14686 ( .A(n10422), .B(n10423), .Z(N29289) );
  NAND U14687 ( .A(n10424), .B(n10425), .Z(n10423) );
  NANDN U14688 ( .A(n10426), .B(n10427), .Z(n10425) );
  NANDN U14689 ( .A(n10427), .B(n10426), .Z(n10422) );
  XOR U14690 ( .A(n10426), .B(n10428), .Z(N29288) );
  XNOR U14691 ( .A(n10424), .B(n10427), .Z(n10428) );
  NAND U14692 ( .A(n10429), .B(n10430), .Z(n10427) );
  NAND U14693 ( .A(n10431), .B(n10432), .Z(n10430) );
  NANDN U14694 ( .A(n10433), .B(n10434), .Z(n10432) );
  NANDN U14695 ( .A(n10434), .B(n10433), .Z(n10429) );
  AND U14696 ( .A(n10435), .B(n10436), .Z(n10424) );
  NAND U14697 ( .A(n10437), .B(n10438), .Z(n10436) );
  OR U14698 ( .A(n10439), .B(n10440), .Z(n10438) );
  NAND U14699 ( .A(n10440), .B(n10439), .Z(n10435) );
  IV U14700 ( .A(n10441), .Z(n10440) );
  AND U14701 ( .A(n10442), .B(n10443), .Z(n10426) );
  NAND U14702 ( .A(n10444), .B(n10445), .Z(n10443) );
  NANDN U14703 ( .A(n10446), .B(n10447), .Z(n10445) );
  NANDN U14704 ( .A(n10447), .B(n10446), .Z(n10442) );
  XOR U14705 ( .A(n10439), .B(n10448), .Z(N29287) );
  XOR U14706 ( .A(n10437), .B(n10441), .Z(n10448) );
  XNOR U14707 ( .A(n10434), .B(n10449), .Z(n10441) );
  XNOR U14708 ( .A(n10431), .B(n10433), .Z(n10449) );
  AND U14709 ( .A(n10450), .B(n10451), .Z(n10433) );
  NANDN U14710 ( .A(n10452), .B(n10453), .Z(n10451) );
  NANDN U14711 ( .A(n10454), .B(n10455), .Z(n10453) );
  IV U14712 ( .A(n10456), .Z(n10455) );
  NAND U14713 ( .A(n10456), .B(n10454), .Z(n10450) );
  AND U14714 ( .A(n10457), .B(n10458), .Z(n10431) );
  NAND U14715 ( .A(n10459), .B(n10460), .Z(n10458) );
  OR U14716 ( .A(n10461), .B(n10462), .Z(n10460) );
  NAND U14717 ( .A(n10462), .B(n10461), .Z(n10457) );
  IV U14718 ( .A(n10463), .Z(n10462) );
  NAND U14719 ( .A(n10464), .B(n10465), .Z(n10434) );
  NANDN U14720 ( .A(n10466), .B(n10467), .Z(n10465) );
  NAND U14721 ( .A(n10468), .B(n10469), .Z(n10467) );
  OR U14722 ( .A(n10469), .B(n10468), .Z(n10464) );
  IV U14723 ( .A(n10470), .Z(n10468) );
  AND U14724 ( .A(n10471), .B(n10472), .Z(n10437) );
  NAND U14725 ( .A(n10473), .B(n10474), .Z(n10472) );
  NANDN U14726 ( .A(n10475), .B(n10476), .Z(n10474) );
  NANDN U14727 ( .A(n10476), .B(n10475), .Z(n10471) );
  XOR U14728 ( .A(n10447), .B(n10477), .Z(n10439) );
  XNOR U14729 ( .A(n10444), .B(n10446), .Z(n10477) );
  AND U14730 ( .A(n10478), .B(n10479), .Z(n10446) );
  NANDN U14731 ( .A(n10480), .B(n10481), .Z(n10479) );
  NANDN U14732 ( .A(n10482), .B(n10483), .Z(n10481) );
  IV U14733 ( .A(n10484), .Z(n10483) );
  NAND U14734 ( .A(n10484), .B(n10482), .Z(n10478) );
  AND U14735 ( .A(n10485), .B(n10486), .Z(n10444) );
  NAND U14736 ( .A(n10487), .B(n10488), .Z(n10486) );
  OR U14737 ( .A(n10489), .B(n10490), .Z(n10488) );
  NAND U14738 ( .A(n10490), .B(n10489), .Z(n10485) );
  IV U14739 ( .A(n10491), .Z(n10490) );
  NAND U14740 ( .A(n10492), .B(n10493), .Z(n10447) );
  NANDN U14741 ( .A(n10494), .B(n10495), .Z(n10493) );
  NAND U14742 ( .A(n10496), .B(n10497), .Z(n10495) );
  OR U14743 ( .A(n10497), .B(n10496), .Z(n10492) );
  IV U14744 ( .A(n10498), .Z(n10496) );
  XOR U14745 ( .A(n10473), .B(n10499), .Z(N29286) );
  XNOR U14746 ( .A(n10476), .B(n10475), .Z(n10499) );
  XNOR U14747 ( .A(n10487), .B(n10500), .Z(n10475) );
  XOR U14748 ( .A(n10491), .B(n10489), .Z(n10500) );
  XOR U14749 ( .A(n10497), .B(n10501), .Z(n10489) );
  XOR U14750 ( .A(n10494), .B(n10498), .Z(n10501) );
  NAND U14751 ( .A(n10502), .B(n10503), .Z(n10498) );
  NAND U14752 ( .A(n10504), .B(n10505), .Z(n10503) );
  NAND U14753 ( .A(n10506), .B(n10507), .Z(n10502) );
  AND U14754 ( .A(n10508), .B(n10509), .Z(n10494) );
  NAND U14755 ( .A(n10510), .B(n10511), .Z(n10509) );
  NAND U14756 ( .A(n10512), .B(n10513), .Z(n10508) );
  NANDN U14757 ( .A(n10514), .B(n10515), .Z(n10497) );
  NANDN U14758 ( .A(n10516), .B(n10517), .Z(n10491) );
  XNOR U14759 ( .A(n10482), .B(n10518), .Z(n10487) );
  XOR U14760 ( .A(n10480), .B(n10484), .Z(n10518) );
  NAND U14761 ( .A(n10519), .B(n10520), .Z(n10484) );
  NAND U14762 ( .A(n10521), .B(n10522), .Z(n10520) );
  NAND U14763 ( .A(n10523), .B(n10524), .Z(n10519) );
  AND U14764 ( .A(n10525), .B(n10526), .Z(n10480) );
  NAND U14765 ( .A(n10527), .B(n10528), .Z(n10526) );
  NAND U14766 ( .A(n10529), .B(n10530), .Z(n10525) );
  AND U14767 ( .A(n10531), .B(n10532), .Z(n10482) );
  NAND U14768 ( .A(n10533), .B(n10534), .Z(n10476) );
  XNOR U14769 ( .A(n10459), .B(n10535), .Z(n10473) );
  XOR U14770 ( .A(n10463), .B(n10461), .Z(n10535) );
  XOR U14771 ( .A(n10469), .B(n10536), .Z(n10461) );
  XOR U14772 ( .A(n10466), .B(n10470), .Z(n10536) );
  NAND U14773 ( .A(n10537), .B(n10538), .Z(n10470) );
  NAND U14774 ( .A(n10539), .B(n10540), .Z(n10538) );
  NAND U14775 ( .A(n10541), .B(n10542), .Z(n10537) );
  AND U14776 ( .A(n10543), .B(n10544), .Z(n10466) );
  NAND U14777 ( .A(n10545), .B(n10546), .Z(n10544) );
  NAND U14778 ( .A(n10547), .B(n10548), .Z(n10543) );
  NANDN U14779 ( .A(n10549), .B(n10550), .Z(n10469) );
  NANDN U14780 ( .A(n10551), .B(n10552), .Z(n10463) );
  XNOR U14781 ( .A(n10454), .B(n10553), .Z(n10459) );
  XOR U14782 ( .A(n10452), .B(n10456), .Z(n10553) );
  NAND U14783 ( .A(n10554), .B(n10555), .Z(n10456) );
  NAND U14784 ( .A(n10556), .B(n10557), .Z(n10555) );
  NAND U14785 ( .A(n10558), .B(n10559), .Z(n10554) );
  AND U14786 ( .A(n10560), .B(n10561), .Z(n10452) );
  NAND U14787 ( .A(n10562), .B(n10563), .Z(n10561) );
  NAND U14788 ( .A(n10564), .B(n10565), .Z(n10560) );
  AND U14789 ( .A(n10566), .B(n10567), .Z(n10454) );
  XOR U14790 ( .A(n10534), .B(n10533), .Z(N29285) );
  XNOR U14791 ( .A(n10552), .B(n10551), .Z(n10533) );
  XNOR U14792 ( .A(n10566), .B(n10567), .Z(n10551) );
  XOR U14793 ( .A(n10563), .B(n10562), .Z(n10567) );
  XOR U14794 ( .A(y[2715]), .B(x[2715]), .Z(n10562) );
  XOR U14795 ( .A(n10565), .B(n10564), .Z(n10563) );
  XOR U14796 ( .A(y[2717]), .B(x[2717]), .Z(n10564) );
  XOR U14797 ( .A(y[2716]), .B(x[2716]), .Z(n10565) );
  XOR U14798 ( .A(n10557), .B(n10556), .Z(n10566) );
  XOR U14799 ( .A(n10559), .B(n10558), .Z(n10556) );
  XOR U14800 ( .A(y[2714]), .B(x[2714]), .Z(n10558) );
  XOR U14801 ( .A(y[2713]), .B(x[2713]), .Z(n10559) );
  XOR U14802 ( .A(y[2712]), .B(x[2712]), .Z(n10557) );
  XNOR U14803 ( .A(n10550), .B(n10549), .Z(n10552) );
  XNOR U14804 ( .A(n10546), .B(n10545), .Z(n10549) );
  XOR U14805 ( .A(n10548), .B(n10547), .Z(n10545) );
  XOR U14806 ( .A(y[2711]), .B(x[2711]), .Z(n10547) );
  XOR U14807 ( .A(y[2710]), .B(x[2710]), .Z(n10548) );
  XOR U14808 ( .A(y[2709]), .B(x[2709]), .Z(n10546) );
  XOR U14809 ( .A(n10540), .B(n10539), .Z(n10550) );
  XOR U14810 ( .A(n10542), .B(n10541), .Z(n10539) );
  XOR U14811 ( .A(y[2708]), .B(x[2708]), .Z(n10541) );
  XOR U14812 ( .A(y[2707]), .B(x[2707]), .Z(n10542) );
  XOR U14813 ( .A(y[2706]), .B(x[2706]), .Z(n10540) );
  XNOR U14814 ( .A(n10517), .B(n10516), .Z(n10534) );
  XNOR U14815 ( .A(n10531), .B(n10532), .Z(n10516) );
  XOR U14816 ( .A(n10528), .B(n10527), .Z(n10532) );
  XOR U14817 ( .A(y[2703]), .B(x[2703]), .Z(n10527) );
  XOR U14818 ( .A(n10530), .B(n10529), .Z(n10528) );
  XOR U14819 ( .A(y[2705]), .B(x[2705]), .Z(n10529) );
  XOR U14820 ( .A(y[2704]), .B(x[2704]), .Z(n10530) );
  XOR U14821 ( .A(n10522), .B(n10521), .Z(n10531) );
  XOR U14822 ( .A(n10524), .B(n10523), .Z(n10521) );
  XOR U14823 ( .A(y[2702]), .B(x[2702]), .Z(n10523) );
  XOR U14824 ( .A(y[2701]), .B(x[2701]), .Z(n10524) );
  XOR U14825 ( .A(y[2700]), .B(x[2700]), .Z(n10522) );
  XNOR U14826 ( .A(n10515), .B(n10514), .Z(n10517) );
  XNOR U14827 ( .A(n10511), .B(n10510), .Z(n10514) );
  XOR U14828 ( .A(n10513), .B(n10512), .Z(n10510) );
  XOR U14829 ( .A(y[2699]), .B(x[2699]), .Z(n10512) );
  XOR U14830 ( .A(y[2698]), .B(x[2698]), .Z(n10513) );
  XOR U14831 ( .A(y[2697]), .B(x[2697]), .Z(n10511) );
  XOR U14832 ( .A(n10505), .B(n10504), .Z(n10515) );
  XOR U14833 ( .A(n10507), .B(n10506), .Z(n10504) );
  XOR U14834 ( .A(y[2696]), .B(x[2696]), .Z(n10506) );
  XOR U14835 ( .A(y[2695]), .B(x[2695]), .Z(n10507) );
  XOR U14836 ( .A(y[2694]), .B(x[2694]), .Z(n10505) );
  NAND U14837 ( .A(n10568), .B(n10569), .Z(N29277) );
  NAND U14838 ( .A(n10570), .B(n10571), .Z(n10569) );
  NANDN U14839 ( .A(n10572), .B(n10573), .Z(n10571) );
  NANDN U14840 ( .A(n10573), .B(n10572), .Z(n10568) );
  XOR U14841 ( .A(n10572), .B(n10574), .Z(N29276) );
  XNOR U14842 ( .A(n10570), .B(n10573), .Z(n10574) );
  NAND U14843 ( .A(n10575), .B(n10576), .Z(n10573) );
  NAND U14844 ( .A(n10577), .B(n10578), .Z(n10576) );
  NANDN U14845 ( .A(n10579), .B(n10580), .Z(n10578) );
  NANDN U14846 ( .A(n10580), .B(n10579), .Z(n10575) );
  AND U14847 ( .A(n10581), .B(n10582), .Z(n10570) );
  NAND U14848 ( .A(n10583), .B(n10584), .Z(n10582) );
  OR U14849 ( .A(n10585), .B(n10586), .Z(n10584) );
  NAND U14850 ( .A(n10586), .B(n10585), .Z(n10581) );
  IV U14851 ( .A(n10587), .Z(n10586) );
  AND U14852 ( .A(n10588), .B(n10589), .Z(n10572) );
  NAND U14853 ( .A(n10590), .B(n10591), .Z(n10589) );
  NANDN U14854 ( .A(n10592), .B(n10593), .Z(n10591) );
  NANDN U14855 ( .A(n10593), .B(n10592), .Z(n10588) );
  XOR U14856 ( .A(n10585), .B(n10594), .Z(N29275) );
  XOR U14857 ( .A(n10583), .B(n10587), .Z(n10594) );
  XNOR U14858 ( .A(n10580), .B(n10595), .Z(n10587) );
  XNOR U14859 ( .A(n10577), .B(n10579), .Z(n10595) );
  AND U14860 ( .A(n10596), .B(n10597), .Z(n10579) );
  NANDN U14861 ( .A(n10598), .B(n10599), .Z(n10597) );
  NANDN U14862 ( .A(n10600), .B(n10601), .Z(n10599) );
  IV U14863 ( .A(n10602), .Z(n10601) );
  NAND U14864 ( .A(n10602), .B(n10600), .Z(n10596) );
  AND U14865 ( .A(n10603), .B(n10604), .Z(n10577) );
  NAND U14866 ( .A(n10605), .B(n10606), .Z(n10604) );
  OR U14867 ( .A(n10607), .B(n10608), .Z(n10606) );
  NAND U14868 ( .A(n10608), .B(n10607), .Z(n10603) );
  IV U14869 ( .A(n10609), .Z(n10608) );
  NAND U14870 ( .A(n10610), .B(n10611), .Z(n10580) );
  NANDN U14871 ( .A(n10612), .B(n10613), .Z(n10611) );
  NAND U14872 ( .A(n10614), .B(n10615), .Z(n10613) );
  OR U14873 ( .A(n10615), .B(n10614), .Z(n10610) );
  IV U14874 ( .A(n10616), .Z(n10614) );
  AND U14875 ( .A(n10617), .B(n10618), .Z(n10583) );
  NAND U14876 ( .A(n10619), .B(n10620), .Z(n10618) );
  NANDN U14877 ( .A(n10621), .B(n10622), .Z(n10620) );
  NANDN U14878 ( .A(n10622), .B(n10621), .Z(n10617) );
  XOR U14879 ( .A(n10593), .B(n10623), .Z(n10585) );
  XNOR U14880 ( .A(n10590), .B(n10592), .Z(n10623) );
  AND U14881 ( .A(n10624), .B(n10625), .Z(n10592) );
  NANDN U14882 ( .A(n10626), .B(n10627), .Z(n10625) );
  NANDN U14883 ( .A(n10628), .B(n10629), .Z(n10627) );
  IV U14884 ( .A(n10630), .Z(n10629) );
  NAND U14885 ( .A(n10630), .B(n10628), .Z(n10624) );
  AND U14886 ( .A(n10631), .B(n10632), .Z(n10590) );
  NAND U14887 ( .A(n10633), .B(n10634), .Z(n10632) );
  OR U14888 ( .A(n10635), .B(n10636), .Z(n10634) );
  NAND U14889 ( .A(n10636), .B(n10635), .Z(n10631) );
  IV U14890 ( .A(n10637), .Z(n10636) );
  NAND U14891 ( .A(n10638), .B(n10639), .Z(n10593) );
  NANDN U14892 ( .A(n10640), .B(n10641), .Z(n10639) );
  NAND U14893 ( .A(n10642), .B(n10643), .Z(n10641) );
  OR U14894 ( .A(n10643), .B(n10642), .Z(n10638) );
  IV U14895 ( .A(n10644), .Z(n10642) );
  XOR U14896 ( .A(n10619), .B(n10645), .Z(N29274) );
  XNOR U14897 ( .A(n10622), .B(n10621), .Z(n10645) );
  XNOR U14898 ( .A(n10633), .B(n10646), .Z(n10621) );
  XOR U14899 ( .A(n10637), .B(n10635), .Z(n10646) );
  XOR U14900 ( .A(n10643), .B(n10647), .Z(n10635) );
  XOR U14901 ( .A(n10640), .B(n10644), .Z(n10647) );
  NAND U14902 ( .A(n10648), .B(n10649), .Z(n10644) );
  NAND U14903 ( .A(n10650), .B(n10651), .Z(n10649) );
  NAND U14904 ( .A(n10652), .B(n10653), .Z(n10648) );
  AND U14905 ( .A(n10654), .B(n10655), .Z(n10640) );
  NAND U14906 ( .A(n10656), .B(n10657), .Z(n10655) );
  NAND U14907 ( .A(n10658), .B(n10659), .Z(n10654) );
  NANDN U14908 ( .A(n10660), .B(n10661), .Z(n10643) );
  NANDN U14909 ( .A(n10662), .B(n10663), .Z(n10637) );
  XNOR U14910 ( .A(n10628), .B(n10664), .Z(n10633) );
  XOR U14911 ( .A(n10626), .B(n10630), .Z(n10664) );
  NAND U14912 ( .A(n10665), .B(n10666), .Z(n10630) );
  NAND U14913 ( .A(n10667), .B(n10668), .Z(n10666) );
  NAND U14914 ( .A(n10669), .B(n10670), .Z(n10665) );
  AND U14915 ( .A(n10671), .B(n10672), .Z(n10626) );
  NAND U14916 ( .A(n10673), .B(n10674), .Z(n10672) );
  NAND U14917 ( .A(n10675), .B(n10676), .Z(n10671) );
  AND U14918 ( .A(n10677), .B(n10678), .Z(n10628) );
  NAND U14919 ( .A(n10679), .B(n10680), .Z(n10622) );
  XNOR U14920 ( .A(n10605), .B(n10681), .Z(n10619) );
  XOR U14921 ( .A(n10609), .B(n10607), .Z(n10681) );
  XOR U14922 ( .A(n10615), .B(n10682), .Z(n10607) );
  XOR U14923 ( .A(n10612), .B(n10616), .Z(n10682) );
  NAND U14924 ( .A(n10683), .B(n10684), .Z(n10616) );
  NAND U14925 ( .A(n10685), .B(n10686), .Z(n10684) );
  NAND U14926 ( .A(n10687), .B(n10688), .Z(n10683) );
  AND U14927 ( .A(n10689), .B(n10690), .Z(n10612) );
  NAND U14928 ( .A(n10691), .B(n10692), .Z(n10690) );
  NAND U14929 ( .A(n10693), .B(n10694), .Z(n10689) );
  NANDN U14930 ( .A(n10695), .B(n10696), .Z(n10615) );
  NANDN U14931 ( .A(n10697), .B(n10698), .Z(n10609) );
  XNOR U14932 ( .A(n10600), .B(n10699), .Z(n10605) );
  XOR U14933 ( .A(n10598), .B(n10602), .Z(n10699) );
  NAND U14934 ( .A(n10700), .B(n10701), .Z(n10602) );
  NAND U14935 ( .A(n10702), .B(n10703), .Z(n10701) );
  NAND U14936 ( .A(n10704), .B(n10705), .Z(n10700) );
  AND U14937 ( .A(n10706), .B(n10707), .Z(n10598) );
  NAND U14938 ( .A(n10708), .B(n10709), .Z(n10707) );
  NAND U14939 ( .A(n10710), .B(n10711), .Z(n10706) );
  AND U14940 ( .A(n10712), .B(n10713), .Z(n10600) );
  XOR U14941 ( .A(n10680), .B(n10679), .Z(N29273) );
  XNOR U14942 ( .A(n10698), .B(n10697), .Z(n10679) );
  XNOR U14943 ( .A(n10712), .B(n10713), .Z(n10697) );
  XOR U14944 ( .A(n10709), .B(n10708), .Z(n10713) );
  XOR U14945 ( .A(y[2691]), .B(x[2691]), .Z(n10708) );
  XOR U14946 ( .A(n10711), .B(n10710), .Z(n10709) );
  XOR U14947 ( .A(y[2693]), .B(x[2693]), .Z(n10710) );
  XOR U14948 ( .A(y[2692]), .B(x[2692]), .Z(n10711) );
  XOR U14949 ( .A(n10703), .B(n10702), .Z(n10712) );
  XOR U14950 ( .A(n10705), .B(n10704), .Z(n10702) );
  XOR U14951 ( .A(y[2690]), .B(x[2690]), .Z(n10704) );
  XOR U14952 ( .A(y[2689]), .B(x[2689]), .Z(n10705) );
  XOR U14953 ( .A(y[2688]), .B(x[2688]), .Z(n10703) );
  XNOR U14954 ( .A(n10696), .B(n10695), .Z(n10698) );
  XNOR U14955 ( .A(n10692), .B(n10691), .Z(n10695) );
  XOR U14956 ( .A(n10694), .B(n10693), .Z(n10691) );
  XOR U14957 ( .A(y[2687]), .B(x[2687]), .Z(n10693) );
  XOR U14958 ( .A(y[2686]), .B(x[2686]), .Z(n10694) );
  XOR U14959 ( .A(y[2685]), .B(x[2685]), .Z(n10692) );
  XOR U14960 ( .A(n10686), .B(n10685), .Z(n10696) );
  XOR U14961 ( .A(n10688), .B(n10687), .Z(n10685) );
  XOR U14962 ( .A(y[2684]), .B(x[2684]), .Z(n10687) );
  XOR U14963 ( .A(y[2683]), .B(x[2683]), .Z(n10688) );
  XOR U14964 ( .A(y[2682]), .B(x[2682]), .Z(n10686) );
  XNOR U14965 ( .A(n10663), .B(n10662), .Z(n10680) );
  XNOR U14966 ( .A(n10677), .B(n10678), .Z(n10662) );
  XOR U14967 ( .A(n10674), .B(n10673), .Z(n10678) );
  XOR U14968 ( .A(y[2679]), .B(x[2679]), .Z(n10673) );
  XOR U14969 ( .A(n10676), .B(n10675), .Z(n10674) );
  XOR U14970 ( .A(y[2681]), .B(x[2681]), .Z(n10675) );
  XOR U14971 ( .A(y[2680]), .B(x[2680]), .Z(n10676) );
  XOR U14972 ( .A(n10668), .B(n10667), .Z(n10677) );
  XOR U14973 ( .A(n10670), .B(n10669), .Z(n10667) );
  XOR U14974 ( .A(y[2678]), .B(x[2678]), .Z(n10669) );
  XOR U14975 ( .A(y[2677]), .B(x[2677]), .Z(n10670) );
  XOR U14976 ( .A(y[2676]), .B(x[2676]), .Z(n10668) );
  XNOR U14977 ( .A(n10661), .B(n10660), .Z(n10663) );
  XNOR U14978 ( .A(n10657), .B(n10656), .Z(n10660) );
  XOR U14979 ( .A(n10659), .B(n10658), .Z(n10656) );
  XOR U14980 ( .A(y[2675]), .B(x[2675]), .Z(n10658) );
  XOR U14981 ( .A(y[2674]), .B(x[2674]), .Z(n10659) );
  XOR U14982 ( .A(y[2673]), .B(x[2673]), .Z(n10657) );
  XOR U14983 ( .A(n10651), .B(n10650), .Z(n10661) );
  XOR U14984 ( .A(n10653), .B(n10652), .Z(n10650) );
  XOR U14985 ( .A(y[2672]), .B(x[2672]), .Z(n10652) );
  XOR U14986 ( .A(y[2671]), .B(x[2671]), .Z(n10653) );
  XOR U14987 ( .A(y[2670]), .B(x[2670]), .Z(n10651) );
  NAND U14988 ( .A(n10714), .B(n10715), .Z(N29265) );
  NAND U14989 ( .A(n10716), .B(n10717), .Z(n10715) );
  NANDN U14990 ( .A(n10718), .B(n10719), .Z(n10717) );
  NANDN U14991 ( .A(n10719), .B(n10718), .Z(n10714) );
  XOR U14992 ( .A(n10718), .B(n10720), .Z(N29264) );
  XNOR U14993 ( .A(n10716), .B(n10719), .Z(n10720) );
  NAND U14994 ( .A(n10721), .B(n10722), .Z(n10719) );
  NAND U14995 ( .A(n10723), .B(n10724), .Z(n10722) );
  NANDN U14996 ( .A(n10725), .B(n10726), .Z(n10724) );
  NANDN U14997 ( .A(n10726), .B(n10725), .Z(n10721) );
  AND U14998 ( .A(n10727), .B(n10728), .Z(n10716) );
  NAND U14999 ( .A(n10729), .B(n10730), .Z(n10728) );
  OR U15000 ( .A(n10731), .B(n10732), .Z(n10730) );
  NAND U15001 ( .A(n10732), .B(n10731), .Z(n10727) );
  IV U15002 ( .A(n10733), .Z(n10732) );
  AND U15003 ( .A(n10734), .B(n10735), .Z(n10718) );
  NAND U15004 ( .A(n10736), .B(n10737), .Z(n10735) );
  NANDN U15005 ( .A(n10738), .B(n10739), .Z(n10737) );
  NANDN U15006 ( .A(n10739), .B(n10738), .Z(n10734) );
  XOR U15007 ( .A(n10731), .B(n10740), .Z(N29263) );
  XOR U15008 ( .A(n10729), .B(n10733), .Z(n10740) );
  XNOR U15009 ( .A(n10726), .B(n10741), .Z(n10733) );
  XNOR U15010 ( .A(n10723), .B(n10725), .Z(n10741) );
  AND U15011 ( .A(n10742), .B(n10743), .Z(n10725) );
  NANDN U15012 ( .A(n10744), .B(n10745), .Z(n10743) );
  NANDN U15013 ( .A(n10746), .B(n10747), .Z(n10745) );
  IV U15014 ( .A(n10748), .Z(n10747) );
  NAND U15015 ( .A(n10748), .B(n10746), .Z(n10742) );
  AND U15016 ( .A(n10749), .B(n10750), .Z(n10723) );
  NAND U15017 ( .A(n10751), .B(n10752), .Z(n10750) );
  OR U15018 ( .A(n10753), .B(n10754), .Z(n10752) );
  NAND U15019 ( .A(n10754), .B(n10753), .Z(n10749) );
  IV U15020 ( .A(n10755), .Z(n10754) );
  NAND U15021 ( .A(n10756), .B(n10757), .Z(n10726) );
  NANDN U15022 ( .A(n10758), .B(n10759), .Z(n10757) );
  NAND U15023 ( .A(n10760), .B(n10761), .Z(n10759) );
  OR U15024 ( .A(n10761), .B(n10760), .Z(n10756) );
  IV U15025 ( .A(n10762), .Z(n10760) );
  AND U15026 ( .A(n10763), .B(n10764), .Z(n10729) );
  NAND U15027 ( .A(n10765), .B(n10766), .Z(n10764) );
  NANDN U15028 ( .A(n10767), .B(n10768), .Z(n10766) );
  NANDN U15029 ( .A(n10768), .B(n10767), .Z(n10763) );
  XOR U15030 ( .A(n10739), .B(n10769), .Z(n10731) );
  XNOR U15031 ( .A(n10736), .B(n10738), .Z(n10769) );
  AND U15032 ( .A(n10770), .B(n10771), .Z(n10738) );
  NANDN U15033 ( .A(n10772), .B(n10773), .Z(n10771) );
  NANDN U15034 ( .A(n10774), .B(n10775), .Z(n10773) );
  IV U15035 ( .A(n10776), .Z(n10775) );
  NAND U15036 ( .A(n10776), .B(n10774), .Z(n10770) );
  AND U15037 ( .A(n10777), .B(n10778), .Z(n10736) );
  NAND U15038 ( .A(n10779), .B(n10780), .Z(n10778) );
  OR U15039 ( .A(n10781), .B(n10782), .Z(n10780) );
  NAND U15040 ( .A(n10782), .B(n10781), .Z(n10777) );
  IV U15041 ( .A(n10783), .Z(n10782) );
  NAND U15042 ( .A(n10784), .B(n10785), .Z(n10739) );
  NANDN U15043 ( .A(n10786), .B(n10787), .Z(n10785) );
  NAND U15044 ( .A(n10788), .B(n10789), .Z(n10787) );
  OR U15045 ( .A(n10789), .B(n10788), .Z(n10784) );
  IV U15046 ( .A(n10790), .Z(n10788) );
  XOR U15047 ( .A(n10765), .B(n10791), .Z(N29262) );
  XNOR U15048 ( .A(n10768), .B(n10767), .Z(n10791) );
  XNOR U15049 ( .A(n10779), .B(n10792), .Z(n10767) );
  XOR U15050 ( .A(n10783), .B(n10781), .Z(n10792) );
  XOR U15051 ( .A(n10789), .B(n10793), .Z(n10781) );
  XOR U15052 ( .A(n10786), .B(n10790), .Z(n10793) );
  NAND U15053 ( .A(n10794), .B(n10795), .Z(n10790) );
  NAND U15054 ( .A(n10796), .B(n10797), .Z(n10795) );
  NAND U15055 ( .A(n10798), .B(n10799), .Z(n10794) );
  AND U15056 ( .A(n10800), .B(n10801), .Z(n10786) );
  NAND U15057 ( .A(n10802), .B(n10803), .Z(n10801) );
  NAND U15058 ( .A(n10804), .B(n10805), .Z(n10800) );
  NANDN U15059 ( .A(n10806), .B(n10807), .Z(n10789) );
  NANDN U15060 ( .A(n10808), .B(n10809), .Z(n10783) );
  XNOR U15061 ( .A(n10774), .B(n10810), .Z(n10779) );
  XOR U15062 ( .A(n10772), .B(n10776), .Z(n10810) );
  NAND U15063 ( .A(n10811), .B(n10812), .Z(n10776) );
  NAND U15064 ( .A(n10813), .B(n10814), .Z(n10812) );
  NAND U15065 ( .A(n10815), .B(n10816), .Z(n10811) );
  AND U15066 ( .A(n10817), .B(n10818), .Z(n10772) );
  NAND U15067 ( .A(n10819), .B(n10820), .Z(n10818) );
  NAND U15068 ( .A(n10821), .B(n10822), .Z(n10817) );
  AND U15069 ( .A(n10823), .B(n10824), .Z(n10774) );
  NAND U15070 ( .A(n10825), .B(n10826), .Z(n10768) );
  XNOR U15071 ( .A(n10751), .B(n10827), .Z(n10765) );
  XOR U15072 ( .A(n10755), .B(n10753), .Z(n10827) );
  XOR U15073 ( .A(n10761), .B(n10828), .Z(n10753) );
  XOR U15074 ( .A(n10758), .B(n10762), .Z(n10828) );
  NAND U15075 ( .A(n10829), .B(n10830), .Z(n10762) );
  NAND U15076 ( .A(n10831), .B(n10832), .Z(n10830) );
  NAND U15077 ( .A(n10833), .B(n10834), .Z(n10829) );
  AND U15078 ( .A(n10835), .B(n10836), .Z(n10758) );
  NAND U15079 ( .A(n10837), .B(n10838), .Z(n10836) );
  NAND U15080 ( .A(n10839), .B(n10840), .Z(n10835) );
  NANDN U15081 ( .A(n10841), .B(n10842), .Z(n10761) );
  NANDN U15082 ( .A(n10843), .B(n10844), .Z(n10755) );
  XNOR U15083 ( .A(n10746), .B(n10845), .Z(n10751) );
  XOR U15084 ( .A(n10744), .B(n10748), .Z(n10845) );
  NAND U15085 ( .A(n10846), .B(n10847), .Z(n10748) );
  NAND U15086 ( .A(n10848), .B(n10849), .Z(n10847) );
  NAND U15087 ( .A(n10850), .B(n10851), .Z(n10846) );
  AND U15088 ( .A(n10852), .B(n10853), .Z(n10744) );
  NAND U15089 ( .A(n10854), .B(n10855), .Z(n10853) );
  NAND U15090 ( .A(n10856), .B(n10857), .Z(n10852) );
  AND U15091 ( .A(n10858), .B(n10859), .Z(n10746) );
  XOR U15092 ( .A(n10826), .B(n10825), .Z(N29261) );
  XNOR U15093 ( .A(n10844), .B(n10843), .Z(n10825) );
  XNOR U15094 ( .A(n10858), .B(n10859), .Z(n10843) );
  XOR U15095 ( .A(n10855), .B(n10854), .Z(n10859) );
  XOR U15096 ( .A(y[2667]), .B(x[2667]), .Z(n10854) );
  XOR U15097 ( .A(n10857), .B(n10856), .Z(n10855) );
  XOR U15098 ( .A(y[2669]), .B(x[2669]), .Z(n10856) );
  XOR U15099 ( .A(y[2668]), .B(x[2668]), .Z(n10857) );
  XOR U15100 ( .A(n10849), .B(n10848), .Z(n10858) );
  XOR U15101 ( .A(n10851), .B(n10850), .Z(n10848) );
  XOR U15102 ( .A(y[2666]), .B(x[2666]), .Z(n10850) );
  XOR U15103 ( .A(y[2665]), .B(x[2665]), .Z(n10851) );
  XOR U15104 ( .A(y[2664]), .B(x[2664]), .Z(n10849) );
  XNOR U15105 ( .A(n10842), .B(n10841), .Z(n10844) );
  XNOR U15106 ( .A(n10838), .B(n10837), .Z(n10841) );
  XOR U15107 ( .A(n10840), .B(n10839), .Z(n10837) );
  XOR U15108 ( .A(y[2663]), .B(x[2663]), .Z(n10839) );
  XOR U15109 ( .A(y[2662]), .B(x[2662]), .Z(n10840) );
  XOR U15110 ( .A(y[2661]), .B(x[2661]), .Z(n10838) );
  XOR U15111 ( .A(n10832), .B(n10831), .Z(n10842) );
  XOR U15112 ( .A(n10834), .B(n10833), .Z(n10831) );
  XOR U15113 ( .A(y[2660]), .B(x[2660]), .Z(n10833) );
  XOR U15114 ( .A(y[2659]), .B(x[2659]), .Z(n10834) );
  XOR U15115 ( .A(y[2658]), .B(x[2658]), .Z(n10832) );
  XNOR U15116 ( .A(n10809), .B(n10808), .Z(n10826) );
  XNOR U15117 ( .A(n10823), .B(n10824), .Z(n10808) );
  XOR U15118 ( .A(n10820), .B(n10819), .Z(n10824) );
  XOR U15119 ( .A(y[2655]), .B(x[2655]), .Z(n10819) );
  XOR U15120 ( .A(n10822), .B(n10821), .Z(n10820) );
  XOR U15121 ( .A(y[2657]), .B(x[2657]), .Z(n10821) );
  XOR U15122 ( .A(y[2656]), .B(x[2656]), .Z(n10822) );
  XOR U15123 ( .A(n10814), .B(n10813), .Z(n10823) );
  XOR U15124 ( .A(n10816), .B(n10815), .Z(n10813) );
  XOR U15125 ( .A(y[2654]), .B(x[2654]), .Z(n10815) );
  XOR U15126 ( .A(y[2653]), .B(x[2653]), .Z(n10816) );
  XOR U15127 ( .A(y[2652]), .B(x[2652]), .Z(n10814) );
  XNOR U15128 ( .A(n10807), .B(n10806), .Z(n10809) );
  XNOR U15129 ( .A(n10803), .B(n10802), .Z(n10806) );
  XOR U15130 ( .A(n10805), .B(n10804), .Z(n10802) );
  XOR U15131 ( .A(y[2651]), .B(x[2651]), .Z(n10804) );
  XOR U15132 ( .A(y[2650]), .B(x[2650]), .Z(n10805) );
  XOR U15133 ( .A(y[2649]), .B(x[2649]), .Z(n10803) );
  XOR U15134 ( .A(n10797), .B(n10796), .Z(n10807) );
  XOR U15135 ( .A(n10799), .B(n10798), .Z(n10796) );
  XOR U15136 ( .A(y[2648]), .B(x[2648]), .Z(n10798) );
  XOR U15137 ( .A(y[2647]), .B(x[2647]), .Z(n10799) );
  XOR U15138 ( .A(y[2646]), .B(x[2646]), .Z(n10797) );
  NAND U15139 ( .A(n10860), .B(n10861), .Z(N29253) );
  NAND U15140 ( .A(n10862), .B(n10863), .Z(n10861) );
  NANDN U15141 ( .A(n10864), .B(n10865), .Z(n10863) );
  NANDN U15142 ( .A(n10865), .B(n10864), .Z(n10860) );
  XOR U15143 ( .A(n10864), .B(n10866), .Z(N29252) );
  XNOR U15144 ( .A(n10862), .B(n10865), .Z(n10866) );
  NAND U15145 ( .A(n10867), .B(n10868), .Z(n10865) );
  NAND U15146 ( .A(n10869), .B(n10870), .Z(n10868) );
  NANDN U15147 ( .A(n10871), .B(n10872), .Z(n10870) );
  NANDN U15148 ( .A(n10872), .B(n10871), .Z(n10867) );
  AND U15149 ( .A(n10873), .B(n10874), .Z(n10862) );
  NAND U15150 ( .A(n10875), .B(n10876), .Z(n10874) );
  OR U15151 ( .A(n10877), .B(n10878), .Z(n10876) );
  NAND U15152 ( .A(n10878), .B(n10877), .Z(n10873) );
  IV U15153 ( .A(n10879), .Z(n10878) );
  AND U15154 ( .A(n10880), .B(n10881), .Z(n10864) );
  NAND U15155 ( .A(n10882), .B(n10883), .Z(n10881) );
  NANDN U15156 ( .A(n10884), .B(n10885), .Z(n10883) );
  NANDN U15157 ( .A(n10885), .B(n10884), .Z(n10880) );
  XOR U15158 ( .A(n10877), .B(n10886), .Z(N29251) );
  XOR U15159 ( .A(n10875), .B(n10879), .Z(n10886) );
  XNOR U15160 ( .A(n10872), .B(n10887), .Z(n10879) );
  XNOR U15161 ( .A(n10869), .B(n10871), .Z(n10887) );
  AND U15162 ( .A(n10888), .B(n10889), .Z(n10871) );
  NANDN U15163 ( .A(n10890), .B(n10891), .Z(n10889) );
  NANDN U15164 ( .A(n10892), .B(n10893), .Z(n10891) );
  IV U15165 ( .A(n10894), .Z(n10893) );
  NAND U15166 ( .A(n10894), .B(n10892), .Z(n10888) );
  AND U15167 ( .A(n10895), .B(n10896), .Z(n10869) );
  NAND U15168 ( .A(n10897), .B(n10898), .Z(n10896) );
  OR U15169 ( .A(n10899), .B(n10900), .Z(n10898) );
  NAND U15170 ( .A(n10900), .B(n10899), .Z(n10895) );
  IV U15171 ( .A(n10901), .Z(n10900) );
  NAND U15172 ( .A(n10902), .B(n10903), .Z(n10872) );
  NANDN U15173 ( .A(n10904), .B(n10905), .Z(n10903) );
  NAND U15174 ( .A(n10906), .B(n10907), .Z(n10905) );
  OR U15175 ( .A(n10907), .B(n10906), .Z(n10902) );
  IV U15176 ( .A(n10908), .Z(n10906) );
  AND U15177 ( .A(n10909), .B(n10910), .Z(n10875) );
  NAND U15178 ( .A(n10911), .B(n10912), .Z(n10910) );
  NANDN U15179 ( .A(n10913), .B(n10914), .Z(n10912) );
  NANDN U15180 ( .A(n10914), .B(n10913), .Z(n10909) );
  XOR U15181 ( .A(n10885), .B(n10915), .Z(n10877) );
  XNOR U15182 ( .A(n10882), .B(n10884), .Z(n10915) );
  AND U15183 ( .A(n10916), .B(n10917), .Z(n10884) );
  NANDN U15184 ( .A(n10918), .B(n10919), .Z(n10917) );
  NANDN U15185 ( .A(n10920), .B(n10921), .Z(n10919) );
  IV U15186 ( .A(n10922), .Z(n10921) );
  NAND U15187 ( .A(n10922), .B(n10920), .Z(n10916) );
  AND U15188 ( .A(n10923), .B(n10924), .Z(n10882) );
  NAND U15189 ( .A(n10925), .B(n10926), .Z(n10924) );
  OR U15190 ( .A(n10927), .B(n10928), .Z(n10926) );
  NAND U15191 ( .A(n10928), .B(n10927), .Z(n10923) );
  IV U15192 ( .A(n10929), .Z(n10928) );
  NAND U15193 ( .A(n10930), .B(n10931), .Z(n10885) );
  NANDN U15194 ( .A(n10932), .B(n10933), .Z(n10931) );
  NAND U15195 ( .A(n10934), .B(n10935), .Z(n10933) );
  OR U15196 ( .A(n10935), .B(n10934), .Z(n10930) );
  IV U15197 ( .A(n10936), .Z(n10934) );
  XOR U15198 ( .A(n10911), .B(n10937), .Z(N29250) );
  XNOR U15199 ( .A(n10914), .B(n10913), .Z(n10937) );
  XNOR U15200 ( .A(n10925), .B(n10938), .Z(n10913) );
  XOR U15201 ( .A(n10929), .B(n10927), .Z(n10938) );
  XOR U15202 ( .A(n10935), .B(n10939), .Z(n10927) );
  XOR U15203 ( .A(n10932), .B(n10936), .Z(n10939) );
  NAND U15204 ( .A(n10940), .B(n10941), .Z(n10936) );
  NAND U15205 ( .A(n10942), .B(n10943), .Z(n10941) );
  NAND U15206 ( .A(n10944), .B(n10945), .Z(n10940) );
  AND U15207 ( .A(n10946), .B(n10947), .Z(n10932) );
  NAND U15208 ( .A(n10948), .B(n10949), .Z(n10947) );
  NAND U15209 ( .A(n10950), .B(n10951), .Z(n10946) );
  NANDN U15210 ( .A(n10952), .B(n10953), .Z(n10935) );
  NANDN U15211 ( .A(n10954), .B(n10955), .Z(n10929) );
  XNOR U15212 ( .A(n10920), .B(n10956), .Z(n10925) );
  XOR U15213 ( .A(n10918), .B(n10922), .Z(n10956) );
  NAND U15214 ( .A(n10957), .B(n10958), .Z(n10922) );
  NAND U15215 ( .A(n10959), .B(n10960), .Z(n10958) );
  NAND U15216 ( .A(n10961), .B(n10962), .Z(n10957) );
  AND U15217 ( .A(n10963), .B(n10964), .Z(n10918) );
  NAND U15218 ( .A(n10965), .B(n10966), .Z(n10964) );
  NAND U15219 ( .A(n10967), .B(n10968), .Z(n10963) );
  AND U15220 ( .A(n10969), .B(n10970), .Z(n10920) );
  NAND U15221 ( .A(n10971), .B(n10972), .Z(n10914) );
  XNOR U15222 ( .A(n10897), .B(n10973), .Z(n10911) );
  XOR U15223 ( .A(n10901), .B(n10899), .Z(n10973) );
  XOR U15224 ( .A(n10907), .B(n10974), .Z(n10899) );
  XOR U15225 ( .A(n10904), .B(n10908), .Z(n10974) );
  NAND U15226 ( .A(n10975), .B(n10976), .Z(n10908) );
  NAND U15227 ( .A(n10977), .B(n10978), .Z(n10976) );
  NAND U15228 ( .A(n10979), .B(n10980), .Z(n10975) );
  AND U15229 ( .A(n10981), .B(n10982), .Z(n10904) );
  NAND U15230 ( .A(n10983), .B(n10984), .Z(n10982) );
  NAND U15231 ( .A(n10985), .B(n10986), .Z(n10981) );
  NANDN U15232 ( .A(n10987), .B(n10988), .Z(n10907) );
  NANDN U15233 ( .A(n10989), .B(n10990), .Z(n10901) );
  XNOR U15234 ( .A(n10892), .B(n10991), .Z(n10897) );
  XOR U15235 ( .A(n10890), .B(n10894), .Z(n10991) );
  NAND U15236 ( .A(n10992), .B(n10993), .Z(n10894) );
  NAND U15237 ( .A(n10994), .B(n10995), .Z(n10993) );
  NAND U15238 ( .A(n10996), .B(n10997), .Z(n10992) );
  AND U15239 ( .A(n10998), .B(n10999), .Z(n10890) );
  NAND U15240 ( .A(n11000), .B(n11001), .Z(n10999) );
  NAND U15241 ( .A(n11002), .B(n11003), .Z(n10998) );
  AND U15242 ( .A(n11004), .B(n11005), .Z(n10892) );
  XOR U15243 ( .A(n10972), .B(n10971), .Z(N29249) );
  XNOR U15244 ( .A(n10990), .B(n10989), .Z(n10971) );
  XNOR U15245 ( .A(n11004), .B(n11005), .Z(n10989) );
  XOR U15246 ( .A(n11001), .B(n11000), .Z(n11005) );
  XOR U15247 ( .A(y[2643]), .B(x[2643]), .Z(n11000) );
  XOR U15248 ( .A(n11003), .B(n11002), .Z(n11001) );
  XOR U15249 ( .A(y[2645]), .B(x[2645]), .Z(n11002) );
  XOR U15250 ( .A(y[2644]), .B(x[2644]), .Z(n11003) );
  XOR U15251 ( .A(n10995), .B(n10994), .Z(n11004) );
  XOR U15252 ( .A(n10997), .B(n10996), .Z(n10994) );
  XOR U15253 ( .A(y[2642]), .B(x[2642]), .Z(n10996) );
  XOR U15254 ( .A(y[2641]), .B(x[2641]), .Z(n10997) );
  XOR U15255 ( .A(y[2640]), .B(x[2640]), .Z(n10995) );
  XNOR U15256 ( .A(n10988), .B(n10987), .Z(n10990) );
  XNOR U15257 ( .A(n10984), .B(n10983), .Z(n10987) );
  XOR U15258 ( .A(n10986), .B(n10985), .Z(n10983) );
  XOR U15259 ( .A(y[2639]), .B(x[2639]), .Z(n10985) );
  XOR U15260 ( .A(y[2638]), .B(x[2638]), .Z(n10986) );
  XOR U15261 ( .A(y[2637]), .B(x[2637]), .Z(n10984) );
  XOR U15262 ( .A(n10978), .B(n10977), .Z(n10988) );
  XOR U15263 ( .A(n10980), .B(n10979), .Z(n10977) );
  XOR U15264 ( .A(y[2636]), .B(x[2636]), .Z(n10979) );
  XOR U15265 ( .A(y[2635]), .B(x[2635]), .Z(n10980) );
  XOR U15266 ( .A(y[2634]), .B(x[2634]), .Z(n10978) );
  XNOR U15267 ( .A(n10955), .B(n10954), .Z(n10972) );
  XNOR U15268 ( .A(n10969), .B(n10970), .Z(n10954) );
  XOR U15269 ( .A(n10966), .B(n10965), .Z(n10970) );
  XOR U15270 ( .A(y[2631]), .B(x[2631]), .Z(n10965) );
  XOR U15271 ( .A(n10968), .B(n10967), .Z(n10966) );
  XOR U15272 ( .A(y[2633]), .B(x[2633]), .Z(n10967) );
  XOR U15273 ( .A(y[2632]), .B(x[2632]), .Z(n10968) );
  XOR U15274 ( .A(n10960), .B(n10959), .Z(n10969) );
  XOR U15275 ( .A(n10962), .B(n10961), .Z(n10959) );
  XOR U15276 ( .A(y[2630]), .B(x[2630]), .Z(n10961) );
  XOR U15277 ( .A(y[2629]), .B(x[2629]), .Z(n10962) );
  XOR U15278 ( .A(y[2628]), .B(x[2628]), .Z(n10960) );
  XNOR U15279 ( .A(n10953), .B(n10952), .Z(n10955) );
  XNOR U15280 ( .A(n10949), .B(n10948), .Z(n10952) );
  XOR U15281 ( .A(n10951), .B(n10950), .Z(n10948) );
  XOR U15282 ( .A(y[2627]), .B(x[2627]), .Z(n10950) );
  XOR U15283 ( .A(y[2626]), .B(x[2626]), .Z(n10951) );
  XOR U15284 ( .A(y[2625]), .B(x[2625]), .Z(n10949) );
  XOR U15285 ( .A(n10943), .B(n10942), .Z(n10953) );
  XOR U15286 ( .A(n10945), .B(n10944), .Z(n10942) );
  XOR U15287 ( .A(y[2624]), .B(x[2624]), .Z(n10944) );
  XOR U15288 ( .A(y[2623]), .B(x[2623]), .Z(n10945) );
  XOR U15289 ( .A(y[2622]), .B(x[2622]), .Z(n10943) );
  NAND U15290 ( .A(n11006), .B(n11007), .Z(N29241) );
  NAND U15291 ( .A(n11008), .B(n11009), .Z(n11007) );
  NANDN U15292 ( .A(n11010), .B(n11011), .Z(n11009) );
  NANDN U15293 ( .A(n11011), .B(n11010), .Z(n11006) );
  XOR U15294 ( .A(n11010), .B(n11012), .Z(N29240) );
  XNOR U15295 ( .A(n11008), .B(n11011), .Z(n11012) );
  NAND U15296 ( .A(n11013), .B(n11014), .Z(n11011) );
  NAND U15297 ( .A(n11015), .B(n11016), .Z(n11014) );
  NANDN U15298 ( .A(n11017), .B(n11018), .Z(n11016) );
  NANDN U15299 ( .A(n11018), .B(n11017), .Z(n11013) );
  AND U15300 ( .A(n11019), .B(n11020), .Z(n11008) );
  NAND U15301 ( .A(n11021), .B(n11022), .Z(n11020) );
  OR U15302 ( .A(n11023), .B(n11024), .Z(n11022) );
  NAND U15303 ( .A(n11024), .B(n11023), .Z(n11019) );
  IV U15304 ( .A(n11025), .Z(n11024) );
  AND U15305 ( .A(n11026), .B(n11027), .Z(n11010) );
  NAND U15306 ( .A(n11028), .B(n11029), .Z(n11027) );
  NANDN U15307 ( .A(n11030), .B(n11031), .Z(n11029) );
  NANDN U15308 ( .A(n11031), .B(n11030), .Z(n11026) );
  XOR U15309 ( .A(n11023), .B(n11032), .Z(N29239) );
  XOR U15310 ( .A(n11021), .B(n11025), .Z(n11032) );
  XNOR U15311 ( .A(n11018), .B(n11033), .Z(n11025) );
  XNOR U15312 ( .A(n11015), .B(n11017), .Z(n11033) );
  AND U15313 ( .A(n11034), .B(n11035), .Z(n11017) );
  NANDN U15314 ( .A(n11036), .B(n11037), .Z(n11035) );
  NANDN U15315 ( .A(n11038), .B(n11039), .Z(n11037) );
  IV U15316 ( .A(n11040), .Z(n11039) );
  NAND U15317 ( .A(n11040), .B(n11038), .Z(n11034) );
  AND U15318 ( .A(n11041), .B(n11042), .Z(n11015) );
  NAND U15319 ( .A(n11043), .B(n11044), .Z(n11042) );
  OR U15320 ( .A(n11045), .B(n11046), .Z(n11044) );
  NAND U15321 ( .A(n11046), .B(n11045), .Z(n11041) );
  IV U15322 ( .A(n11047), .Z(n11046) );
  NAND U15323 ( .A(n11048), .B(n11049), .Z(n11018) );
  NANDN U15324 ( .A(n11050), .B(n11051), .Z(n11049) );
  NAND U15325 ( .A(n11052), .B(n11053), .Z(n11051) );
  OR U15326 ( .A(n11053), .B(n11052), .Z(n11048) );
  IV U15327 ( .A(n11054), .Z(n11052) );
  AND U15328 ( .A(n11055), .B(n11056), .Z(n11021) );
  NAND U15329 ( .A(n11057), .B(n11058), .Z(n11056) );
  NANDN U15330 ( .A(n11059), .B(n11060), .Z(n11058) );
  NANDN U15331 ( .A(n11060), .B(n11059), .Z(n11055) );
  XOR U15332 ( .A(n11031), .B(n11061), .Z(n11023) );
  XNOR U15333 ( .A(n11028), .B(n11030), .Z(n11061) );
  AND U15334 ( .A(n11062), .B(n11063), .Z(n11030) );
  NANDN U15335 ( .A(n11064), .B(n11065), .Z(n11063) );
  NANDN U15336 ( .A(n11066), .B(n11067), .Z(n11065) );
  IV U15337 ( .A(n11068), .Z(n11067) );
  NAND U15338 ( .A(n11068), .B(n11066), .Z(n11062) );
  AND U15339 ( .A(n11069), .B(n11070), .Z(n11028) );
  NAND U15340 ( .A(n11071), .B(n11072), .Z(n11070) );
  OR U15341 ( .A(n11073), .B(n11074), .Z(n11072) );
  NAND U15342 ( .A(n11074), .B(n11073), .Z(n11069) );
  IV U15343 ( .A(n11075), .Z(n11074) );
  NAND U15344 ( .A(n11076), .B(n11077), .Z(n11031) );
  NANDN U15345 ( .A(n11078), .B(n11079), .Z(n11077) );
  NAND U15346 ( .A(n11080), .B(n11081), .Z(n11079) );
  OR U15347 ( .A(n11081), .B(n11080), .Z(n11076) );
  IV U15348 ( .A(n11082), .Z(n11080) );
  XOR U15349 ( .A(n11057), .B(n11083), .Z(N29238) );
  XNOR U15350 ( .A(n11060), .B(n11059), .Z(n11083) );
  XNOR U15351 ( .A(n11071), .B(n11084), .Z(n11059) );
  XOR U15352 ( .A(n11075), .B(n11073), .Z(n11084) );
  XOR U15353 ( .A(n11081), .B(n11085), .Z(n11073) );
  XOR U15354 ( .A(n11078), .B(n11082), .Z(n11085) );
  NAND U15355 ( .A(n11086), .B(n11087), .Z(n11082) );
  NAND U15356 ( .A(n11088), .B(n11089), .Z(n11087) );
  NAND U15357 ( .A(n11090), .B(n11091), .Z(n11086) );
  AND U15358 ( .A(n11092), .B(n11093), .Z(n11078) );
  NAND U15359 ( .A(n11094), .B(n11095), .Z(n11093) );
  NAND U15360 ( .A(n11096), .B(n11097), .Z(n11092) );
  NANDN U15361 ( .A(n11098), .B(n11099), .Z(n11081) );
  NANDN U15362 ( .A(n11100), .B(n11101), .Z(n11075) );
  XNOR U15363 ( .A(n11066), .B(n11102), .Z(n11071) );
  XOR U15364 ( .A(n11064), .B(n11068), .Z(n11102) );
  NAND U15365 ( .A(n11103), .B(n11104), .Z(n11068) );
  NAND U15366 ( .A(n11105), .B(n11106), .Z(n11104) );
  NAND U15367 ( .A(n11107), .B(n11108), .Z(n11103) );
  AND U15368 ( .A(n11109), .B(n11110), .Z(n11064) );
  NAND U15369 ( .A(n11111), .B(n11112), .Z(n11110) );
  NAND U15370 ( .A(n11113), .B(n11114), .Z(n11109) );
  AND U15371 ( .A(n11115), .B(n11116), .Z(n11066) );
  NAND U15372 ( .A(n11117), .B(n11118), .Z(n11060) );
  XNOR U15373 ( .A(n11043), .B(n11119), .Z(n11057) );
  XOR U15374 ( .A(n11047), .B(n11045), .Z(n11119) );
  XOR U15375 ( .A(n11053), .B(n11120), .Z(n11045) );
  XOR U15376 ( .A(n11050), .B(n11054), .Z(n11120) );
  NAND U15377 ( .A(n11121), .B(n11122), .Z(n11054) );
  NAND U15378 ( .A(n11123), .B(n11124), .Z(n11122) );
  NAND U15379 ( .A(n11125), .B(n11126), .Z(n11121) );
  AND U15380 ( .A(n11127), .B(n11128), .Z(n11050) );
  NAND U15381 ( .A(n11129), .B(n11130), .Z(n11128) );
  NAND U15382 ( .A(n11131), .B(n11132), .Z(n11127) );
  NANDN U15383 ( .A(n11133), .B(n11134), .Z(n11053) );
  NANDN U15384 ( .A(n11135), .B(n11136), .Z(n11047) );
  XNOR U15385 ( .A(n11038), .B(n11137), .Z(n11043) );
  XOR U15386 ( .A(n11036), .B(n11040), .Z(n11137) );
  NAND U15387 ( .A(n11138), .B(n11139), .Z(n11040) );
  NAND U15388 ( .A(n11140), .B(n11141), .Z(n11139) );
  NAND U15389 ( .A(n11142), .B(n11143), .Z(n11138) );
  AND U15390 ( .A(n11144), .B(n11145), .Z(n11036) );
  NAND U15391 ( .A(n11146), .B(n11147), .Z(n11145) );
  NAND U15392 ( .A(n11148), .B(n11149), .Z(n11144) );
  AND U15393 ( .A(n11150), .B(n11151), .Z(n11038) );
  XOR U15394 ( .A(n11118), .B(n11117), .Z(N29237) );
  XNOR U15395 ( .A(n11136), .B(n11135), .Z(n11117) );
  XNOR U15396 ( .A(n11150), .B(n11151), .Z(n11135) );
  XOR U15397 ( .A(n11147), .B(n11146), .Z(n11151) );
  XOR U15398 ( .A(y[2619]), .B(x[2619]), .Z(n11146) );
  XOR U15399 ( .A(n11149), .B(n11148), .Z(n11147) );
  XOR U15400 ( .A(y[2621]), .B(x[2621]), .Z(n11148) );
  XOR U15401 ( .A(y[2620]), .B(x[2620]), .Z(n11149) );
  XOR U15402 ( .A(n11141), .B(n11140), .Z(n11150) );
  XOR U15403 ( .A(n11143), .B(n11142), .Z(n11140) );
  XOR U15404 ( .A(y[2618]), .B(x[2618]), .Z(n11142) );
  XOR U15405 ( .A(y[2617]), .B(x[2617]), .Z(n11143) );
  XOR U15406 ( .A(y[2616]), .B(x[2616]), .Z(n11141) );
  XNOR U15407 ( .A(n11134), .B(n11133), .Z(n11136) );
  XNOR U15408 ( .A(n11130), .B(n11129), .Z(n11133) );
  XOR U15409 ( .A(n11132), .B(n11131), .Z(n11129) );
  XOR U15410 ( .A(y[2615]), .B(x[2615]), .Z(n11131) );
  XOR U15411 ( .A(y[2614]), .B(x[2614]), .Z(n11132) );
  XOR U15412 ( .A(y[2613]), .B(x[2613]), .Z(n11130) );
  XOR U15413 ( .A(n11124), .B(n11123), .Z(n11134) );
  XOR U15414 ( .A(n11126), .B(n11125), .Z(n11123) );
  XOR U15415 ( .A(y[2612]), .B(x[2612]), .Z(n11125) );
  XOR U15416 ( .A(y[2611]), .B(x[2611]), .Z(n11126) );
  XOR U15417 ( .A(y[2610]), .B(x[2610]), .Z(n11124) );
  XNOR U15418 ( .A(n11101), .B(n11100), .Z(n11118) );
  XNOR U15419 ( .A(n11115), .B(n11116), .Z(n11100) );
  XOR U15420 ( .A(n11112), .B(n11111), .Z(n11116) );
  XOR U15421 ( .A(y[2607]), .B(x[2607]), .Z(n11111) );
  XOR U15422 ( .A(n11114), .B(n11113), .Z(n11112) );
  XOR U15423 ( .A(y[2609]), .B(x[2609]), .Z(n11113) );
  XOR U15424 ( .A(y[2608]), .B(x[2608]), .Z(n11114) );
  XOR U15425 ( .A(n11106), .B(n11105), .Z(n11115) );
  XOR U15426 ( .A(n11108), .B(n11107), .Z(n11105) );
  XOR U15427 ( .A(y[2606]), .B(x[2606]), .Z(n11107) );
  XOR U15428 ( .A(y[2605]), .B(x[2605]), .Z(n11108) );
  XOR U15429 ( .A(y[2604]), .B(x[2604]), .Z(n11106) );
  XNOR U15430 ( .A(n11099), .B(n11098), .Z(n11101) );
  XNOR U15431 ( .A(n11095), .B(n11094), .Z(n11098) );
  XOR U15432 ( .A(n11097), .B(n11096), .Z(n11094) );
  XOR U15433 ( .A(y[2603]), .B(x[2603]), .Z(n11096) );
  XOR U15434 ( .A(y[2602]), .B(x[2602]), .Z(n11097) );
  XOR U15435 ( .A(y[2601]), .B(x[2601]), .Z(n11095) );
  XOR U15436 ( .A(n11089), .B(n11088), .Z(n11099) );
  XOR U15437 ( .A(n11091), .B(n11090), .Z(n11088) );
  XOR U15438 ( .A(y[2600]), .B(x[2600]), .Z(n11090) );
  XOR U15439 ( .A(y[2599]), .B(x[2599]), .Z(n11091) );
  XOR U15440 ( .A(y[2598]), .B(x[2598]), .Z(n11089) );
  NAND U15441 ( .A(n11152), .B(n11153), .Z(N29229) );
  NAND U15442 ( .A(n11154), .B(n11155), .Z(n11153) );
  NANDN U15443 ( .A(n11156), .B(n11157), .Z(n11155) );
  NANDN U15444 ( .A(n11157), .B(n11156), .Z(n11152) );
  XOR U15445 ( .A(n11156), .B(n11158), .Z(N29228) );
  XNOR U15446 ( .A(n11154), .B(n11157), .Z(n11158) );
  NAND U15447 ( .A(n11159), .B(n11160), .Z(n11157) );
  NAND U15448 ( .A(n11161), .B(n11162), .Z(n11160) );
  NANDN U15449 ( .A(n11163), .B(n11164), .Z(n11162) );
  NANDN U15450 ( .A(n11164), .B(n11163), .Z(n11159) );
  AND U15451 ( .A(n11165), .B(n11166), .Z(n11154) );
  NAND U15452 ( .A(n11167), .B(n11168), .Z(n11166) );
  OR U15453 ( .A(n11169), .B(n11170), .Z(n11168) );
  NAND U15454 ( .A(n11170), .B(n11169), .Z(n11165) );
  IV U15455 ( .A(n11171), .Z(n11170) );
  AND U15456 ( .A(n11172), .B(n11173), .Z(n11156) );
  NAND U15457 ( .A(n11174), .B(n11175), .Z(n11173) );
  NANDN U15458 ( .A(n11176), .B(n11177), .Z(n11175) );
  NANDN U15459 ( .A(n11177), .B(n11176), .Z(n11172) );
  XOR U15460 ( .A(n11169), .B(n11178), .Z(N29227) );
  XOR U15461 ( .A(n11167), .B(n11171), .Z(n11178) );
  XNOR U15462 ( .A(n11164), .B(n11179), .Z(n11171) );
  XNOR U15463 ( .A(n11161), .B(n11163), .Z(n11179) );
  AND U15464 ( .A(n11180), .B(n11181), .Z(n11163) );
  NANDN U15465 ( .A(n11182), .B(n11183), .Z(n11181) );
  NANDN U15466 ( .A(n11184), .B(n11185), .Z(n11183) );
  IV U15467 ( .A(n11186), .Z(n11185) );
  NAND U15468 ( .A(n11186), .B(n11184), .Z(n11180) );
  AND U15469 ( .A(n11187), .B(n11188), .Z(n11161) );
  NAND U15470 ( .A(n11189), .B(n11190), .Z(n11188) );
  OR U15471 ( .A(n11191), .B(n11192), .Z(n11190) );
  NAND U15472 ( .A(n11192), .B(n11191), .Z(n11187) );
  IV U15473 ( .A(n11193), .Z(n11192) );
  NAND U15474 ( .A(n11194), .B(n11195), .Z(n11164) );
  NANDN U15475 ( .A(n11196), .B(n11197), .Z(n11195) );
  NAND U15476 ( .A(n11198), .B(n11199), .Z(n11197) );
  OR U15477 ( .A(n11199), .B(n11198), .Z(n11194) );
  IV U15478 ( .A(n11200), .Z(n11198) );
  AND U15479 ( .A(n11201), .B(n11202), .Z(n11167) );
  NAND U15480 ( .A(n11203), .B(n11204), .Z(n11202) );
  NANDN U15481 ( .A(n11205), .B(n11206), .Z(n11204) );
  NANDN U15482 ( .A(n11206), .B(n11205), .Z(n11201) );
  XOR U15483 ( .A(n11177), .B(n11207), .Z(n11169) );
  XNOR U15484 ( .A(n11174), .B(n11176), .Z(n11207) );
  AND U15485 ( .A(n11208), .B(n11209), .Z(n11176) );
  NANDN U15486 ( .A(n11210), .B(n11211), .Z(n11209) );
  NANDN U15487 ( .A(n11212), .B(n11213), .Z(n11211) );
  IV U15488 ( .A(n11214), .Z(n11213) );
  NAND U15489 ( .A(n11214), .B(n11212), .Z(n11208) );
  AND U15490 ( .A(n11215), .B(n11216), .Z(n11174) );
  NAND U15491 ( .A(n11217), .B(n11218), .Z(n11216) );
  OR U15492 ( .A(n11219), .B(n11220), .Z(n11218) );
  NAND U15493 ( .A(n11220), .B(n11219), .Z(n11215) );
  IV U15494 ( .A(n11221), .Z(n11220) );
  NAND U15495 ( .A(n11222), .B(n11223), .Z(n11177) );
  NANDN U15496 ( .A(n11224), .B(n11225), .Z(n11223) );
  NAND U15497 ( .A(n11226), .B(n11227), .Z(n11225) );
  OR U15498 ( .A(n11227), .B(n11226), .Z(n11222) );
  IV U15499 ( .A(n11228), .Z(n11226) );
  XOR U15500 ( .A(n11203), .B(n11229), .Z(N29226) );
  XNOR U15501 ( .A(n11206), .B(n11205), .Z(n11229) );
  XNOR U15502 ( .A(n11217), .B(n11230), .Z(n11205) );
  XOR U15503 ( .A(n11221), .B(n11219), .Z(n11230) );
  XOR U15504 ( .A(n11227), .B(n11231), .Z(n11219) );
  XOR U15505 ( .A(n11224), .B(n11228), .Z(n11231) );
  NAND U15506 ( .A(n11232), .B(n11233), .Z(n11228) );
  NAND U15507 ( .A(n11234), .B(n11235), .Z(n11233) );
  NAND U15508 ( .A(n11236), .B(n11237), .Z(n11232) );
  AND U15509 ( .A(n11238), .B(n11239), .Z(n11224) );
  NAND U15510 ( .A(n11240), .B(n11241), .Z(n11239) );
  NAND U15511 ( .A(n11242), .B(n11243), .Z(n11238) );
  NANDN U15512 ( .A(n11244), .B(n11245), .Z(n11227) );
  NANDN U15513 ( .A(n11246), .B(n11247), .Z(n11221) );
  XNOR U15514 ( .A(n11212), .B(n11248), .Z(n11217) );
  XOR U15515 ( .A(n11210), .B(n11214), .Z(n11248) );
  NAND U15516 ( .A(n11249), .B(n11250), .Z(n11214) );
  NAND U15517 ( .A(n11251), .B(n11252), .Z(n11250) );
  NAND U15518 ( .A(n11253), .B(n11254), .Z(n11249) );
  AND U15519 ( .A(n11255), .B(n11256), .Z(n11210) );
  NAND U15520 ( .A(n11257), .B(n11258), .Z(n11256) );
  NAND U15521 ( .A(n11259), .B(n11260), .Z(n11255) );
  AND U15522 ( .A(n11261), .B(n11262), .Z(n11212) );
  NAND U15523 ( .A(n11263), .B(n11264), .Z(n11206) );
  XNOR U15524 ( .A(n11189), .B(n11265), .Z(n11203) );
  XOR U15525 ( .A(n11193), .B(n11191), .Z(n11265) );
  XOR U15526 ( .A(n11199), .B(n11266), .Z(n11191) );
  XOR U15527 ( .A(n11196), .B(n11200), .Z(n11266) );
  NAND U15528 ( .A(n11267), .B(n11268), .Z(n11200) );
  NAND U15529 ( .A(n11269), .B(n11270), .Z(n11268) );
  NAND U15530 ( .A(n11271), .B(n11272), .Z(n11267) );
  AND U15531 ( .A(n11273), .B(n11274), .Z(n11196) );
  NAND U15532 ( .A(n11275), .B(n11276), .Z(n11274) );
  NAND U15533 ( .A(n11277), .B(n11278), .Z(n11273) );
  NANDN U15534 ( .A(n11279), .B(n11280), .Z(n11199) );
  NANDN U15535 ( .A(n11281), .B(n11282), .Z(n11193) );
  XNOR U15536 ( .A(n11184), .B(n11283), .Z(n11189) );
  XOR U15537 ( .A(n11182), .B(n11186), .Z(n11283) );
  NAND U15538 ( .A(n11284), .B(n11285), .Z(n11186) );
  NAND U15539 ( .A(n11286), .B(n11287), .Z(n11285) );
  NAND U15540 ( .A(n11288), .B(n11289), .Z(n11284) );
  AND U15541 ( .A(n11290), .B(n11291), .Z(n11182) );
  NAND U15542 ( .A(n11292), .B(n11293), .Z(n11291) );
  NAND U15543 ( .A(n11294), .B(n11295), .Z(n11290) );
  AND U15544 ( .A(n11296), .B(n11297), .Z(n11184) );
  XOR U15545 ( .A(n11264), .B(n11263), .Z(N29225) );
  XNOR U15546 ( .A(n11282), .B(n11281), .Z(n11263) );
  XNOR U15547 ( .A(n11296), .B(n11297), .Z(n11281) );
  XOR U15548 ( .A(n11293), .B(n11292), .Z(n11297) );
  XOR U15549 ( .A(y[2595]), .B(x[2595]), .Z(n11292) );
  XOR U15550 ( .A(n11295), .B(n11294), .Z(n11293) );
  XOR U15551 ( .A(y[2597]), .B(x[2597]), .Z(n11294) );
  XOR U15552 ( .A(y[2596]), .B(x[2596]), .Z(n11295) );
  XOR U15553 ( .A(n11287), .B(n11286), .Z(n11296) );
  XOR U15554 ( .A(n11289), .B(n11288), .Z(n11286) );
  XOR U15555 ( .A(y[2594]), .B(x[2594]), .Z(n11288) );
  XOR U15556 ( .A(y[2593]), .B(x[2593]), .Z(n11289) );
  XOR U15557 ( .A(y[2592]), .B(x[2592]), .Z(n11287) );
  XNOR U15558 ( .A(n11280), .B(n11279), .Z(n11282) );
  XNOR U15559 ( .A(n11276), .B(n11275), .Z(n11279) );
  XOR U15560 ( .A(n11278), .B(n11277), .Z(n11275) );
  XOR U15561 ( .A(y[2591]), .B(x[2591]), .Z(n11277) );
  XOR U15562 ( .A(y[2590]), .B(x[2590]), .Z(n11278) );
  XOR U15563 ( .A(y[2589]), .B(x[2589]), .Z(n11276) );
  XOR U15564 ( .A(n11270), .B(n11269), .Z(n11280) );
  XOR U15565 ( .A(n11272), .B(n11271), .Z(n11269) );
  XOR U15566 ( .A(y[2588]), .B(x[2588]), .Z(n11271) );
  XOR U15567 ( .A(y[2587]), .B(x[2587]), .Z(n11272) );
  XOR U15568 ( .A(y[2586]), .B(x[2586]), .Z(n11270) );
  XNOR U15569 ( .A(n11247), .B(n11246), .Z(n11264) );
  XNOR U15570 ( .A(n11261), .B(n11262), .Z(n11246) );
  XOR U15571 ( .A(n11258), .B(n11257), .Z(n11262) );
  XOR U15572 ( .A(y[2583]), .B(x[2583]), .Z(n11257) );
  XOR U15573 ( .A(n11260), .B(n11259), .Z(n11258) );
  XOR U15574 ( .A(y[2585]), .B(x[2585]), .Z(n11259) );
  XOR U15575 ( .A(y[2584]), .B(x[2584]), .Z(n11260) );
  XOR U15576 ( .A(n11252), .B(n11251), .Z(n11261) );
  XOR U15577 ( .A(n11254), .B(n11253), .Z(n11251) );
  XOR U15578 ( .A(y[2582]), .B(x[2582]), .Z(n11253) );
  XOR U15579 ( .A(y[2581]), .B(x[2581]), .Z(n11254) );
  XOR U15580 ( .A(y[2580]), .B(x[2580]), .Z(n11252) );
  XNOR U15581 ( .A(n11245), .B(n11244), .Z(n11247) );
  XNOR U15582 ( .A(n11241), .B(n11240), .Z(n11244) );
  XOR U15583 ( .A(n11243), .B(n11242), .Z(n11240) );
  XOR U15584 ( .A(y[2579]), .B(x[2579]), .Z(n11242) );
  XOR U15585 ( .A(y[2578]), .B(x[2578]), .Z(n11243) );
  XOR U15586 ( .A(y[2577]), .B(x[2577]), .Z(n11241) );
  XOR U15587 ( .A(n11235), .B(n11234), .Z(n11245) );
  XOR U15588 ( .A(n11237), .B(n11236), .Z(n11234) );
  XOR U15589 ( .A(y[2576]), .B(x[2576]), .Z(n11236) );
  XOR U15590 ( .A(y[2575]), .B(x[2575]), .Z(n11237) );
  XOR U15591 ( .A(y[2574]), .B(x[2574]), .Z(n11235) );
  NAND U15592 ( .A(n11298), .B(n11299), .Z(N29217) );
  NAND U15593 ( .A(n11300), .B(n11301), .Z(n11299) );
  NANDN U15594 ( .A(n11302), .B(n11303), .Z(n11301) );
  NANDN U15595 ( .A(n11303), .B(n11302), .Z(n11298) );
  XOR U15596 ( .A(n11302), .B(n11304), .Z(N29216) );
  XNOR U15597 ( .A(n11300), .B(n11303), .Z(n11304) );
  NAND U15598 ( .A(n11305), .B(n11306), .Z(n11303) );
  NAND U15599 ( .A(n11307), .B(n11308), .Z(n11306) );
  NANDN U15600 ( .A(n11309), .B(n11310), .Z(n11308) );
  NANDN U15601 ( .A(n11310), .B(n11309), .Z(n11305) );
  AND U15602 ( .A(n11311), .B(n11312), .Z(n11300) );
  NAND U15603 ( .A(n11313), .B(n11314), .Z(n11312) );
  OR U15604 ( .A(n11315), .B(n11316), .Z(n11314) );
  NAND U15605 ( .A(n11316), .B(n11315), .Z(n11311) );
  IV U15606 ( .A(n11317), .Z(n11316) );
  AND U15607 ( .A(n11318), .B(n11319), .Z(n11302) );
  NAND U15608 ( .A(n11320), .B(n11321), .Z(n11319) );
  NANDN U15609 ( .A(n11322), .B(n11323), .Z(n11321) );
  NANDN U15610 ( .A(n11323), .B(n11322), .Z(n11318) );
  XOR U15611 ( .A(n11315), .B(n11324), .Z(N29215) );
  XOR U15612 ( .A(n11313), .B(n11317), .Z(n11324) );
  XNOR U15613 ( .A(n11310), .B(n11325), .Z(n11317) );
  XNOR U15614 ( .A(n11307), .B(n11309), .Z(n11325) );
  AND U15615 ( .A(n11326), .B(n11327), .Z(n11309) );
  NANDN U15616 ( .A(n11328), .B(n11329), .Z(n11327) );
  NANDN U15617 ( .A(n11330), .B(n11331), .Z(n11329) );
  IV U15618 ( .A(n11332), .Z(n11331) );
  NAND U15619 ( .A(n11332), .B(n11330), .Z(n11326) );
  AND U15620 ( .A(n11333), .B(n11334), .Z(n11307) );
  NAND U15621 ( .A(n11335), .B(n11336), .Z(n11334) );
  OR U15622 ( .A(n11337), .B(n11338), .Z(n11336) );
  NAND U15623 ( .A(n11338), .B(n11337), .Z(n11333) );
  IV U15624 ( .A(n11339), .Z(n11338) );
  NAND U15625 ( .A(n11340), .B(n11341), .Z(n11310) );
  NANDN U15626 ( .A(n11342), .B(n11343), .Z(n11341) );
  NAND U15627 ( .A(n11344), .B(n11345), .Z(n11343) );
  OR U15628 ( .A(n11345), .B(n11344), .Z(n11340) );
  IV U15629 ( .A(n11346), .Z(n11344) );
  AND U15630 ( .A(n11347), .B(n11348), .Z(n11313) );
  NAND U15631 ( .A(n11349), .B(n11350), .Z(n11348) );
  NANDN U15632 ( .A(n11351), .B(n11352), .Z(n11350) );
  NANDN U15633 ( .A(n11352), .B(n11351), .Z(n11347) );
  XOR U15634 ( .A(n11323), .B(n11353), .Z(n11315) );
  XNOR U15635 ( .A(n11320), .B(n11322), .Z(n11353) );
  AND U15636 ( .A(n11354), .B(n11355), .Z(n11322) );
  NANDN U15637 ( .A(n11356), .B(n11357), .Z(n11355) );
  NANDN U15638 ( .A(n11358), .B(n11359), .Z(n11357) );
  IV U15639 ( .A(n11360), .Z(n11359) );
  NAND U15640 ( .A(n11360), .B(n11358), .Z(n11354) );
  AND U15641 ( .A(n11361), .B(n11362), .Z(n11320) );
  NAND U15642 ( .A(n11363), .B(n11364), .Z(n11362) );
  OR U15643 ( .A(n11365), .B(n11366), .Z(n11364) );
  NAND U15644 ( .A(n11366), .B(n11365), .Z(n11361) );
  IV U15645 ( .A(n11367), .Z(n11366) );
  NAND U15646 ( .A(n11368), .B(n11369), .Z(n11323) );
  NANDN U15647 ( .A(n11370), .B(n11371), .Z(n11369) );
  NAND U15648 ( .A(n11372), .B(n11373), .Z(n11371) );
  OR U15649 ( .A(n11373), .B(n11372), .Z(n11368) );
  IV U15650 ( .A(n11374), .Z(n11372) );
  XOR U15651 ( .A(n11349), .B(n11375), .Z(N29214) );
  XNOR U15652 ( .A(n11352), .B(n11351), .Z(n11375) );
  XNOR U15653 ( .A(n11363), .B(n11376), .Z(n11351) );
  XOR U15654 ( .A(n11367), .B(n11365), .Z(n11376) );
  XOR U15655 ( .A(n11373), .B(n11377), .Z(n11365) );
  XOR U15656 ( .A(n11370), .B(n11374), .Z(n11377) );
  NAND U15657 ( .A(n11378), .B(n11379), .Z(n11374) );
  NAND U15658 ( .A(n11380), .B(n11381), .Z(n11379) );
  NAND U15659 ( .A(n11382), .B(n11383), .Z(n11378) );
  AND U15660 ( .A(n11384), .B(n11385), .Z(n11370) );
  NAND U15661 ( .A(n11386), .B(n11387), .Z(n11385) );
  NAND U15662 ( .A(n11388), .B(n11389), .Z(n11384) );
  NANDN U15663 ( .A(n11390), .B(n11391), .Z(n11373) );
  NANDN U15664 ( .A(n11392), .B(n11393), .Z(n11367) );
  XNOR U15665 ( .A(n11358), .B(n11394), .Z(n11363) );
  XOR U15666 ( .A(n11356), .B(n11360), .Z(n11394) );
  NAND U15667 ( .A(n11395), .B(n11396), .Z(n11360) );
  NAND U15668 ( .A(n11397), .B(n11398), .Z(n11396) );
  NAND U15669 ( .A(n11399), .B(n11400), .Z(n11395) );
  AND U15670 ( .A(n11401), .B(n11402), .Z(n11356) );
  NAND U15671 ( .A(n11403), .B(n11404), .Z(n11402) );
  NAND U15672 ( .A(n11405), .B(n11406), .Z(n11401) );
  AND U15673 ( .A(n11407), .B(n11408), .Z(n11358) );
  NAND U15674 ( .A(n11409), .B(n11410), .Z(n11352) );
  XNOR U15675 ( .A(n11335), .B(n11411), .Z(n11349) );
  XOR U15676 ( .A(n11339), .B(n11337), .Z(n11411) );
  XOR U15677 ( .A(n11345), .B(n11412), .Z(n11337) );
  XOR U15678 ( .A(n11342), .B(n11346), .Z(n11412) );
  NAND U15679 ( .A(n11413), .B(n11414), .Z(n11346) );
  NAND U15680 ( .A(n11415), .B(n11416), .Z(n11414) );
  NAND U15681 ( .A(n11417), .B(n11418), .Z(n11413) );
  AND U15682 ( .A(n11419), .B(n11420), .Z(n11342) );
  NAND U15683 ( .A(n11421), .B(n11422), .Z(n11420) );
  NAND U15684 ( .A(n11423), .B(n11424), .Z(n11419) );
  NANDN U15685 ( .A(n11425), .B(n11426), .Z(n11345) );
  NANDN U15686 ( .A(n11427), .B(n11428), .Z(n11339) );
  XNOR U15687 ( .A(n11330), .B(n11429), .Z(n11335) );
  XOR U15688 ( .A(n11328), .B(n11332), .Z(n11429) );
  NAND U15689 ( .A(n11430), .B(n11431), .Z(n11332) );
  NAND U15690 ( .A(n11432), .B(n11433), .Z(n11431) );
  NAND U15691 ( .A(n11434), .B(n11435), .Z(n11430) );
  AND U15692 ( .A(n11436), .B(n11437), .Z(n11328) );
  NAND U15693 ( .A(n11438), .B(n11439), .Z(n11437) );
  NAND U15694 ( .A(n11440), .B(n11441), .Z(n11436) );
  AND U15695 ( .A(n11442), .B(n11443), .Z(n11330) );
  XOR U15696 ( .A(n11410), .B(n11409), .Z(N29213) );
  XNOR U15697 ( .A(n11428), .B(n11427), .Z(n11409) );
  XNOR U15698 ( .A(n11442), .B(n11443), .Z(n11427) );
  XOR U15699 ( .A(n11439), .B(n11438), .Z(n11443) );
  XOR U15700 ( .A(y[2571]), .B(x[2571]), .Z(n11438) );
  XOR U15701 ( .A(n11441), .B(n11440), .Z(n11439) );
  XOR U15702 ( .A(y[2573]), .B(x[2573]), .Z(n11440) );
  XOR U15703 ( .A(y[2572]), .B(x[2572]), .Z(n11441) );
  XOR U15704 ( .A(n11433), .B(n11432), .Z(n11442) );
  XOR U15705 ( .A(n11435), .B(n11434), .Z(n11432) );
  XOR U15706 ( .A(y[2570]), .B(x[2570]), .Z(n11434) );
  XOR U15707 ( .A(y[2569]), .B(x[2569]), .Z(n11435) );
  XOR U15708 ( .A(y[2568]), .B(x[2568]), .Z(n11433) );
  XNOR U15709 ( .A(n11426), .B(n11425), .Z(n11428) );
  XNOR U15710 ( .A(n11422), .B(n11421), .Z(n11425) );
  XOR U15711 ( .A(n11424), .B(n11423), .Z(n11421) );
  XOR U15712 ( .A(y[2567]), .B(x[2567]), .Z(n11423) );
  XOR U15713 ( .A(y[2566]), .B(x[2566]), .Z(n11424) );
  XOR U15714 ( .A(y[2565]), .B(x[2565]), .Z(n11422) );
  XOR U15715 ( .A(n11416), .B(n11415), .Z(n11426) );
  XOR U15716 ( .A(n11418), .B(n11417), .Z(n11415) );
  XOR U15717 ( .A(y[2564]), .B(x[2564]), .Z(n11417) );
  XOR U15718 ( .A(y[2563]), .B(x[2563]), .Z(n11418) );
  XOR U15719 ( .A(y[2562]), .B(x[2562]), .Z(n11416) );
  XNOR U15720 ( .A(n11393), .B(n11392), .Z(n11410) );
  XNOR U15721 ( .A(n11407), .B(n11408), .Z(n11392) );
  XOR U15722 ( .A(n11404), .B(n11403), .Z(n11408) );
  XOR U15723 ( .A(y[2559]), .B(x[2559]), .Z(n11403) );
  XOR U15724 ( .A(n11406), .B(n11405), .Z(n11404) );
  XOR U15725 ( .A(y[2561]), .B(x[2561]), .Z(n11405) );
  XOR U15726 ( .A(y[2560]), .B(x[2560]), .Z(n11406) );
  XOR U15727 ( .A(n11398), .B(n11397), .Z(n11407) );
  XOR U15728 ( .A(n11400), .B(n11399), .Z(n11397) );
  XOR U15729 ( .A(y[2558]), .B(x[2558]), .Z(n11399) );
  XOR U15730 ( .A(y[2557]), .B(x[2557]), .Z(n11400) );
  XOR U15731 ( .A(y[2556]), .B(x[2556]), .Z(n11398) );
  XNOR U15732 ( .A(n11391), .B(n11390), .Z(n11393) );
  XNOR U15733 ( .A(n11387), .B(n11386), .Z(n11390) );
  XOR U15734 ( .A(n11389), .B(n11388), .Z(n11386) );
  XOR U15735 ( .A(y[2555]), .B(x[2555]), .Z(n11388) );
  XOR U15736 ( .A(y[2554]), .B(x[2554]), .Z(n11389) );
  XOR U15737 ( .A(y[2553]), .B(x[2553]), .Z(n11387) );
  XOR U15738 ( .A(n11381), .B(n11380), .Z(n11391) );
  XOR U15739 ( .A(n11383), .B(n11382), .Z(n11380) );
  XOR U15740 ( .A(y[2552]), .B(x[2552]), .Z(n11382) );
  XOR U15741 ( .A(y[2551]), .B(x[2551]), .Z(n11383) );
  XOR U15742 ( .A(y[2550]), .B(x[2550]), .Z(n11381) );
  NAND U15743 ( .A(n11444), .B(n11445), .Z(N29205) );
  NAND U15744 ( .A(n11446), .B(n11447), .Z(n11445) );
  NANDN U15745 ( .A(n11448), .B(n11449), .Z(n11447) );
  NANDN U15746 ( .A(n11449), .B(n11448), .Z(n11444) );
  XOR U15747 ( .A(n11448), .B(n11450), .Z(N29204) );
  XNOR U15748 ( .A(n11446), .B(n11449), .Z(n11450) );
  NAND U15749 ( .A(n11451), .B(n11452), .Z(n11449) );
  NAND U15750 ( .A(n11453), .B(n11454), .Z(n11452) );
  NANDN U15751 ( .A(n11455), .B(n11456), .Z(n11454) );
  NANDN U15752 ( .A(n11456), .B(n11455), .Z(n11451) );
  AND U15753 ( .A(n11457), .B(n11458), .Z(n11446) );
  NAND U15754 ( .A(n11459), .B(n11460), .Z(n11458) );
  OR U15755 ( .A(n11461), .B(n11462), .Z(n11460) );
  NAND U15756 ( .A(n11462), .B(n11461), .Z(n11457) );
  IV U15757 ( .A(n11463), .Z(n11462) );
  AND U15758 ( .A(n11464), .B(n11465), .Z(n11448) );
  NAND U15759 ( .A(n11466), .B(n11467), .Z(n11465) );
  NANDN U15760 ( .A(n11468), .B(n11469), .Z(n11467) );
  NANDN U15761 ( .A(n11469), .B(n11468), .Z(n11464) );
  XOR U15762 ( .A(n11461), .B(n11470), .Z(N29203) );
  XOR U15763 ( .A(n11459), .B(n11463), .Z(n11470) );
  XNOR U15764 ( .A(n11456), .B(n11471), .Z(n11463) );
  XNOR U15765 ( .A(n11453), .B(n11455), .Z(n11471) );
  AND U15766 ( .A(n11472), .B(n11473), .Z(n11455) );
  NANDN U15767 ( .A(n11474), .B(n11475), .Z(n11473) );
  NANDN U15768 ( .A(n11476), .B(n11477), .Z(n11475) );
  IV U15769 ( .A(n11478), .Z(n11477) );
  NAND U15770 ( .A(n11478), .B(n11476), .Z(n11472) );
  AND U15771 ( .A(n11479), .B(n11480), .Z(n11453) );
  NAND U15772 ( .A(n11481), .B(n11482), .Z(n11480) );
  OR U15773 ( .A(n11483), .B(n11484), .Z(n11482) );
  NAND U15774 ( .A(n11484), .B(n11483), .Z(n11479) );
  IV U15775 ( .A(n11485), .Z(n11484) );
  NAND U15776 ( .A(n11486), .B(n11487), .Z(n11456) );
  NANDN U15777 ( .A(n11488), .B(n11489), .Z(n11487) );
  NAND U15778 ( .A(n11490), .B(n11491), .Z(n11489) );
  OR U15779 ( .A(n11491), .B(n11490), .Z(n11486) );
  IV U15780 ( .A(n11492), .Z(n11490) );
  AND U15781 ( .A(n11493), .B(n11494), .Z(n11459) );
  NAND U15782 ( .A(n11495), .B(n11496), .Z(n11494) );
  NANDN U15783 ( .A(n11497), .B(n11498), .Z(n11496) );
  NANDN U15784 ( .A(n11498), .B(n11497), .Z(n11493) );
  XOR U15785 ( .A(n11469), .B(n11499), .Z(n11461) );
  XNOR U15786 ( .A(n11466), .B(n11468), .Z(n11499) );
  AND U15787 ( .A(n11500), .B(n11501), .Z(n11468) );
  NANDN U15788 ( .A(n11502), .B(n11503), .Z(n11501) );
  NANDN U15789 ( .A(n11504), .B(n11505), .Z(n11503) );
  IV U15790 ( .A(n11506), .Z(n11505) );
  NAND U15791 ( .A(n11506), .B(n11504), .Z(n11500) );
  AND U15792 ( .A(n11507), .B(n11508), .Z(n11466) );
  NAND U15793 ( .A(n11509), .B(n11510), .Z(n11508) );
  OR U15794 ( .A(n11511), .B(n11512), .Z(n11510) );
  NAND U15795 ( .A(n11512), .B(n11511), .Z(n11507) );
  IV U15796 ( .A(n11513), .Z(n11512) );
  NAND U15797 ( .A(n11514), .B(n11515), .Z(n11469) );
  NANDN U15798 ( .A(n11516), .B(n11517), .Z(n11515) );
  NAND U15799 ( .A(n11518), .B(n11519), .Z(n11517) );
  OR U15800 ( .A(n11519), .B(n11518), .Z(n11514) );
  IV U15801 ( .A(n11520), .Z(n11518) );
  XOR U15802 ( .A(n11495), .B(n11521), .Z(N29202) );
  XNOR U15803 ( .A(n11498), .B(n11497), .Z(n11521) );
  XNOR U15804 ( .A(n11509), .B(n11522), .Z(n11497) );
  XOR U15805 ( .A(n11513), .B(n11511), .Z(n11522) );
  XOR U15806 ( .A(n11519), .B(n11523), .Z(n11511) );
  XOR U15807 ( .A(n11516), .B(n11520), .Z(n11523) );
  NAND U15808 ( .A(n11524), .B(n11525), .Z(n11520) );
  NAND U15809 ( .A(n11526), .B(n11527), .Z(n11525) );
  NAND U15810 ( .A(n11528), .B(n11529), .Z(n11524) );
  AND U15811 ( .A(n11530), .B(n11531), .Z(n11516) );
  NAND U15812 ( .A(n11532), .B(n11533), .Z(n11531) );
  NAND U15813 ( .A(n11534), .B(n11535), .Z(n11530) );
  NANDN U15814 ( .A(n11536), .B(n11537), .Z(n11519) );
  NANDN U15815 ( .A(n11538), .B(n11539), .Z(n11513) );
  XNOR U15816 ( .A(n11504), .B(n11540), .Z(n11509) );
  XOR U15817 ( .A(n11502), .B(n11506), .Z(n11540) );
  NAND U15818 ( .A(n11541), .B(n11542), .Z(n11506) );
  NAND U15819 ( .A(n11543), .B(n11544), .Z(n11542) );
  NAND U15820 ( .A(n11545), .B(n11546), .Z(n11541) );
  AND U15821 ( .A(n11547), .B(n11548), .Z(n11502) );
  NAND U15822 ( .A(n11549), .B(n11550), .Z(n11548) );
  NAND U15823 ( .A(n11551), .B(n11552), .Z(n11547) );
  AND U15824 ( .A(n11553), .B(n11554), .Z(n11504) );
  NAND U15825 ( .A(n11555), .B(n11556), .Z(n11498) );
  XNOR U15826 ( .A(n11481), .B(n11557), .Z(n11495) );
  XOR U15827 ( .A(n11485), .B(n11483), .Z(n11557) );
  XOR U15828 ( .A(n11491), .B(n11558), .Z(n11483) );
  XOR U15829 ( .A(n11488), .B(n11492), .Z(n11558) );
  NAND U15830 ( .A(n11559), .B(n11560), .Z(n11492) );
  NAND U15831 ( .A(n11561), .B(n11562), .Z(n11560) );
  NAND U15832 ( .A(n11563), .B(n11564), .Z(n11559) );
  AND U15833 ( .A(n11565), .B(n11566), .Z(n11488) );
  NAND U15834 ( .A(n11567), .B(n11568), .Z(n11566) );
  NAND U15835 ( .A(n11569), .B(n11570), .Z(n11565) );
  NANDN U15836 ( .A(n11571), .B(n11572), .Z(n11491) );
  NANDN U15837 ( .A(n11573), .B(n11574), .Z(n11485) );
  XNOR U15838 ( .A(n11476), .B(n11575), .Z(n11481) );
  XOR U15839 ( .A(n11474), .B(n11478), .Z(n11575) );
  NAND U15840 ( .A(n11576), .B(n11577), .Z(n11478) );
  NAND U15841 ( .A(n11578), .B(n11579), .Z(n11577) );
  NAND U15842 ( .A(n11580), .B(n11581), .Z(n11576) );
  AND U15843 ( .A(n11582), .B(n11583), .Z(n11474) );
  NAND U15844 ( .A(n11584), .B(n11585), .Z(n11583) );
  NAND U15845 ( .A(n11586), .B(n11587), .Z(n11582) );
  AND U15846 ( .A(n11588), .B(n11589), .Z(n11476) );
  XOR U15847 ( .A(n11556), .B(n11555), .Z(N29201) );
  XNOR U15848 ( .A(n11574), .B(n11573), .Z(n11555) );
  XNOR U15849 ( .A(n11588), .B(n11589), .Z(n11573) );
  XOR U15850 ( .A(n11585), .B(n11584), .Z(n11589) );
  XOR U15851 ( .A(y[2547]), .B(x[2547]), .Z(n11584) );
  XOR U15852 ( .A(n11587), .B(n11586), .Z(n11585) );
  XOR U15853 ( .A(y[2549]), .B(x[2549]), .Z(n11586) );
  XOR U15854 ( .A(y[2548]), .B(x[2548]), .Z(n11587) );
  XOR U15855 ( .A(n11579), .B(n11578), .Z(n11588) );
  XOR U15856 ( .A(n11581), .B(n11580), .Z(n11578) );
  XOR U15857 ( .A(y[2546]), .B(x[2546]), .Z(n11580) );
  XOR U15858 ( .A(y[2545]), .B(x[2545]), .Z(n11581) );
  XOR U15859 ( .A(y[2544]), .B(x[2544]), .Z(n11579) );
  XNOR U15860 ( .A(n11572), .B(n11571), .Z(n11574) );
  XNOR U15861 ( .A(n11568), .B(n11567), .Z(n11571) );
  XOR U15862 ( .A(n11570), .B(n11569), .Z(n11567) );
  XOR U15863 ( .A(y[2543]), .B(x[2543]), .Z(n11569) );
  XOR U15864 ( .A(y[2542]), .B(x[2542]), .Z(n11570) );
  XOR U15865 ( .A(y[2541]), .B(x[2541]), .Z(n11568) );
  XOR U15866 ( .A(n11562), .B(n11561), .Z(n11572) );
  XOR U15867 ( .A(n11564), .B(n11563), .Z(n11561) );
  XOR U15868 ( .A(y[2540]), .B(x[2540]), .Z(n11563) );
  XOR U15869 ( .A(y[2539]), .B(x[2539]), .Z(n11564) );
  XOR U15870 ( .A(y[2538]), .B(x[2538]), .Z(n11562) );
  XNOR U15871 ( .A(n11539), .B(n11538), .Z(n11556) );
  XNOR U15872 ( .A(n11553), .B(n11554), .Z(n11538) );
  XOR U15873 ( .A(n11550), .B(n11549), .Z(n11554) );
  XOR U15874 ( .A(y[2535]), .B(x[2535]), .Z(n11549) );
  XOR U15875 ( .A(n11552), .B(n11551), .Z(n11550) );
  XOR U15876 ( .A(y[2537]), .B(x[2537]), .Z(n11551) );
  XOR U15877 ( .A(y[2536]), .B(x[2536]), .Z(n11552) );
  XOR U15878 ( .A(n11544), .B(n11543), .Z(n11553) );
  XOR U15879 ( .A(n11546), .B(n11545), .Z(n11543) );
  XOR U15880 ( .A(y[2534]), .B(x[2534]), .Z(n11545) );
  XOR U15881 ( .A(y[2533]), .B(x[2533]), .Z(n11546) );
  XOR U15882 ( .A(y[2532]), .B(x[2532]), .Z(n11544) );
  XNOR U15883 ( .A(n11537), .B(n11536), .Z(n11539) );
  XNOR U15884 ( .A(n11533), .B(n11532), .Z(n11536) );
  XOR U15885 ( .A(n11535), .B(n11534), .Z(n11532) );
  XOR U15886 ( .A(y[2531]), .B(x[2531]), .Z(n11534) );
  XOR U15887 ( .A(y[2530]), .B(x[2530]), .Z(n11535) );
  XOR U15888 ( .A(y[2529]), .B(x[2529]), .Z(n11533) );
  XOR U15889 ( .A(n11527), .B(n11526), .Z(n11537) );
  XOR U15890 ( .A(n11529), .B(n11528), .Z(n11526) );
  XOR U15891 ( .A(y[2528]), .B(x[2528]), .Z(n11528) );
  XOR U15892 ( .A(y[2527]), .B(x[2527]), .Z(n11529) );
  XOR U15893 ( .A(y[2526]), .B(x[2526]), .Z(n11527) );
  NAND U15894 ( .A(n11590), .B(n11591), .Z(N29193) );
  NAND U15895 ( .A(n11592), .B(n11593), .Z(n11591) );
  NANDN U15896 ( .A(n11594), .B(n11595), .Z(n11593) );
  NANDN U15897 ( .A(n11595), .B(n11594), .Z(n11590) );
  XOR U15898 ( .A(n11594), .B(n11596), .Z(N29192) );
  XNOR U15899 ( .A(n11592), .B(n11595), .Z(n11596) );
  NAND U15900 ( .A(n11597), .B(n11598), .Z(n11595) );
  NAND U15901 ( .A(n11599), .B(n11600), .Z(n11598) );
  NANDN U15902 ( .A(n11601), .B(n11602), .Z(n11600) );
  NANDN U15903 ( .A(n11602), .B(n11601), .Z(n11597) );
  AND U15904 ( .A(n11603), .B(n11604), .Z(n11592) );
  NAND U15905 ( .A(n11605), .B(n11606), .Z(n11604) );
  OR U15906 ( .A(n11607), .B(n11608), .Z(n11606) );
  NAND U15907 ( .A(n11608), .B(n11607), .Z(n11603) );
  IV U15908 ( .A(n11609), .Z(n11608) );
  AND U15909 ( .A(n11610), .B(n11611), .Z(n11594) );
  NAND U15910 ( .A(n11612), .B(n11613), .Z(n11611) );
  NANDN U15911 ( .A(n11614), .B(n11615), .Z(n11613) );
  NANDN U15912 ( .A(n11615), .B(n11614), .Z(n11610) );
  XOR U15913 ( .A(n11607), .B(n11616), .Z(N29191) );
  XOR U15914 ( .A(n11605), .B(n11609), .Z(n11616) );
  XNOR U15915 ( .A(n11602), .B(n11617), .Z(n11609) );
  XNOR U15916 ( .A(n11599), .B(n11601), .Z(n11617) );
  AND U15917 ( .A(n11618), .B(n11619), .Z(n11601) );
  NANDN U15918 ( .A(n11620), .B(n11621), .Z(n11619) );
  NANDN U15919 ( .A(n11622), .B(n11623), .Z(n11621) );
  IV U15920 ( .A(n11624), .Z(n11623) );
  NAND U15921 ( .A(n11624), .B(n11622), .Z(n11618) );
  AND U15922 ( .A(n11625), .B(n11626), .Z(n11599) );
  NAND U15923 ( .A(n11627), .B(n11628), .Z(n11626) );
  OR U15924 ( .A(n11629), .B(n11630), .Z(n11628) );
  NAND U15925 ( .A(n11630), .B(n11629), .Z(n11625) );
  IV U15926 ( .A(n11631), .Z(n11630) );
  NAND U15927 ( .A(n11632), .B(n11633), .Z(n11602) );
  NANDN U15928 ( .A(n11634), .B(n11635), .Z(n11633) );
  NAND U15929 ( .A(n11636), .B(n11637), .Z(n11635) );
  OR U15930 ( .A(n11637), .B(n11636), .Z(n11632) );
  IV U15931 ( .A(n11638), .Z(n11636) );
  AND U15932 ( .A(n11639), .B(n11640), .Z(n11605) );
  NAND U15933 ( .A(n11641), .B(n11642), .Z(n11640) );
  NANDN U15934 ( .A(n11643), .B(n11644), .Z(n11642) );
  NANDN U15935 ( .A(n11644), .B(n11643), .Z(n11639) );
  XOR U15936 ( .A(n11615), .B(n11645), .Z(n11607) );
  XNOR U15937 ( .A(n11612), .B(n11614), .Z(n11645) );
  AND U15938 ( .A(n11646), .B(n11647), .Z(n11614) );
  NANDN U15939 ( .A(n11648), .B(n11649), .Z(n11647) );
  NANDN U15940 ( .A(n11650), .B(n11651), .Z(n11649) );
  IV U15941 ( .A(n11652), .Z(n11651) );
  NAND U15942 ( .A(n11652), .B(n11650), .Z(n11646) );
  AND U15943 ( .A(n11653), .B(n11654), .Z(n11612) );
  NAND U15944 ( .A(n11655), .B(n11656), .Z(n11654) );
  OR U15945 ( .A(n11657), .B(n11658), .Z(n11656) );
  NAND U15946 ( .A(n11658), .B(n11657), .Z(n11653) );
  IV U15947 ( .A(n11659), .Z(n11658) );
  NAND U15948 ( .A(n11660), .B(n11661), .Z(n11615) );
  NANDN U15949 ( .A(n11662), .B(n11663), .Z(n11661) );
  NAND U15950 ( .A(n11664), .B(n11665), .Z(n11663) );
  OR U15951 ( .A(n11665), .B(n11664), .Z(n11660) );
  IV U15952 ( .A(n11666), .Z(n11664) );
  XOR U15953 ( .A(n11641), .B(n11667), .Z(N29190) );
  XNOR U15954 ( .A(n11644), .B(n11643), .Z(n11667) );
  XNOR U15955 ( .A(n11655), .B(n11668), .Z(n11643) );
  XOR U15956 ( .A(n11659), .B(n11657), .Z(n11668) );
  XOR U15957 ( .A(n11665), .B(n11669), .Z(n11657) );
  XOR U15958 ( .A(n11662), .B(n11666), .Z(n11669) );
  NAND U15959 ( .A(n11670), .B(n11671), .Z(n11666) );
  NAND U15960 ( .A(n11672), .B(n11673), .Z(n11671) );
  NAND U15961 ( .A(n11674), .B(n11675), .Z(n11670) );
  AND U15962 ( .A(n11676), .B(n11677), .Z(n11662) );
  NAND U15963 ( .A(n11678), .B(n11679), .Z(n11677) );
  NAND U15964 ( .A(n11680), .B(n11681), .Z(n11676) );
  NANDN U15965 ( .A(n11682), .B(n11683), .Z(n11665) );
  NANDN U15966 ( .A(n11684), .B(n11685), .Z(n11659) );
  XNOR U15967 ( .A(n11650), .B(n11686), .Z(n11655) );
  XOR U15968 ( .A(n11648), .B(n11652), .Z(n11686) );
  NAND U15969 ( .A(n11687), .B(n11688), .Z(n11652) );
  NAND U15970 ( .A(n11689), .B(n11690), .Z(n11688) );
  NAND U15971 ( .A(n11691), .B(n11692), .Z(n11687) );
  AND U15972 ( .A(n11693), .B(n11694), .Z(n11648) );
  NAND U15973 ( .A(n11695), .B(n11696), .Z(n11694) );
  NAND U15974 ( .A(n11697), .B(n11698), .Z(n11693) );
  AND U15975 ( .A(n11699), .B(n11700), .Z(n11650) );
  NAND U15976 ( .A(n11701), .B(n11702), .Z(n11644) );
  XNOR U15977 ( .A(n11627), .B(n11703), .Z(n11641) );
  XOR U15978 ( .A(n11631), .B(n11629), .Z(n11703) );
  XOR U15979 ( .A(n11637), .B(n11704), .Z(n11629) );
  XOR U15980 ( .A(n11634), .B(n11638), .Z(n11704) );
  NAND U15981 ( .A(n11705), .B(n11706), .Z(n11638) );
  NAND U15982 ( .A(n11707), .B(n11708), .Z(n11706) );
  NAND U15983 ( .A(n11709), .B(n11710), .Z(n11705) );
  AND U15984 ( .A(n11711), .B(n11712), .Z(n11634) );
  NAND U15985 ( .A(n11713), .B(n11714), .Z(n11712) );
  NAND U15986 ( .A(n11715), .B(n11716), .Z(n11711) );
  NANDN U15987 ( .A(n11717), .B(n11718), .Z(n11637) );
  NANDN U15988 ( .A(n11719), .B(n11720), .Z(n11631) );
  XNOR U15989 ( .A(n11622), .B(n11721), .Z(n11627) );
  XOR U15990 ( .A(n11620), .B(n11624), .Z(n11721) );
  NAND U15991 ( .A(n11722), .B(n11723), .Z(n11624) );
  NAND U15992 ( .A(n11724), .B(n11725), .Z(n11723) );
  NAND U15993 ( .A(n11726), .B(n11727), .Z(n11722) );
  AND U15994 ( .A(n11728), .B(n11729), .Z(n11620) );
  NAND U15995 ( .A(n11730), .B(n11731), .Z(n11729) );
  NAND U15996 ( .A(n11732), .B(n11733), .Z(n11728) );
  AND U15997 ( .A(n11734), .B(n11735), .Z(n11622) );
  XOR U15998 ( .A(n11702), .B(n11701), .Z(N29189) );
  XNOR U15999 ( .A(n11720), .B(n11719), .Z(n11701) );
  XNOR U16000 ( .A(n11734), .B(n11735), .Z(n11719) );
  XOR U16001 ( .A(n11731), .B(n11730), .Z(n11735) );
  XOR U16002 ( .A(y[2523]), .B(x[2523]), .Z(n11730) );
  XOR U16003 ( .A(n11733), .B(n11732), .Z(n11731) );
  XOR U16004 ( .A(y[2525]), .B(x[2525]), .Z(n11732) );
  XOR U16005 ( .A(y[2524]), .B(x[2524]), .Z(n11733) );
  XOR U16006 ( .A(n11725), .B(n11724), .Z(n11734) );
  XOR U16007 ( .A(n11727), .B(n11726), .Z(n11724) );
  XOR U16008 ( .A(y[2522]), .B(x[2522]), .Z(n11726) );
  XOR U16009 ( .A(y[2521]), .B(x[2521]), .Z(n11727) );
  XOR U16010 ( .A(y[2520]), .B(x[2520]), .Z(n11725) );
  XNOR U16011 ( .A(n11718), .B(n11717), .Z(n11720) );
  XNOR U16012 ( .A(n11714), .B(n11713), .Z(n11717) );
  XOR U16013 ( .A(n11716), .B(n11715), .Z(n11713) );
  XOR U16014 ( .A(y[2519]), .B(x[2519]), .Z(n11715) );
  XOR U16015 ( .A(y[2518]), .B(x[2518]), .Z(n11716) );
  XOR U16016 ( .A(y[2517]), .B(x[2517]), .Z(n11714) );
  XOR U16017 ( .A(n11708), .B(n11707), .Z(n11718) );
  XOR U16018 ( .A(n11710), .B(n11709), .Z(n11707) );
  XOR U16019 ( .A(y[2516]), .B(x[2516]), .Z(n11709) );
  XOR U16020 ( .A(y[2515]), .B(x[2515]), .Z(n11710) );
  XOR U16021 ( .A(y[2514]), .B(x[2514]), .Z(n11708) );
  XNOR U16022 ( .A(n11685), .B(n11684), .Z(n11702) );
  XNOR U16023 ( .A(n11699), .B(n11700), .Z(n11684) );
  XOR U16024 ( .A(n11696), .B(n11695), .Z(n11700) );
  XOR U16025 ( .A(y[2511]), .B(x[2511]), .Z(n11695) );
  XOR U16026 ( .A(n11698), .B(n11697), .Z(n11696) );
  XOR U16027 ( .A(y[2513]), .B(x[2513]), .Z(n11697) );
  XOR U16028 ( .A(y[2512]), .B(x[2512]), .Z(n11698) );
  XOR U16029 ( .A(n11690), .B(n11689), .Z(n11699) );
  XOR U16030 ( .A(n11692), .B(n11691), .Z(n11689) );
  XOR U16031 ( .A(y[2510]), .B(x[2510]), .Z(n11691) );
  XOR U16032 ( .A(y[2509]), .B(x[2509]), .Z(n11692) );
  XOR U16033 ( .A(y[2508]), .B(x[2508]), .Z(n11690) );
  XNOR U16034 ( .A(n11683), .B(n11682), .Z(n11685) );
  XNOR U16035 ( .A(n11679), .B(n11678), .Z(n11682) );
  XOR U16036 ( .A(n11681), .B(n11680), .Z(n11678) );
  XOR U16037 ( .A(y[2507]), .B(x[2507]), .Z(n11680) );
  XOR U16038 ( .A(y[2506]), .B(x[2506]), .Z(n11681) );
  XOR U16039 ( .A(y[2505]), .B(x[2505]), .Z(n11679) );
  XOR U16040 ( .A(n11673), .B(n11672), .Z(n11683) );
  XOR U16041 ( .A(n11675), .B(n11674), .Z(n11672) );
  XOR U16042 ( .A(y[2504]), .B(x[2504]), .Z(n11674) );
  XOR U16043 ( .A(y[2503]), .B(x[2503]), .Z(n11675) );
  XOR U16044 ( .A(y[2502]), .B(x[2502]), .Z(n11673) );
  NAND U16045 ( .A(n11736), .B(n11737), .Z(N29181) );
  NAND U16046 ( .A(n11738), .B(n11739), .Z(n11737) );
  NANDN U16047 ( .A(n11740), .B(n11741), .Z(n11739) );
  NANDN U16048 ( .A(n11741), .B(n11740), .Z(n11736) );
  XOR U16049 ( .A(n11740), .B(n11742), .Z(N29180) );
  XNOR U16050 ( .A(n11738), .B(n11741), .Z(n11742) );
  NAND U16051 ( .A(n11743), .B(n11744), .Z(n11741) );
  NAND U16052 ( .A(n11745), .B(n11746), .Z(n11744) );
  NANDN U16053 ( .A(n11747), .B(n11748), .Z(n11746) );
  NANDN U16054 ( .A(n11748), .B(n11747), .Z(n11743) );
  AND U16055 ( .A(n11749), .B(n11750), .Z(n11738) );
  NAND U16056 ( .A(n11751), .B(n11752), .Z(n11750) );
  OR U16057 ( .A(n11753), .B(n11754), .Z(n11752) );
  NAND U16058 ( .A(n11754), .B(n11753), .Z(n11749) );
  IV U16059 ( .A(n11755), .Z(n11754) );
  AND U16060 ( .A(n11756), .B(n11757), .Z(n11740) );
  NAND U16061 ( .A(n11758), .B(n11759), .Z(n11757) );
  NANDN U16062 ( .A(n11760), .B(n11761), .Z(n11759) );
  NANDN U16063 ( .A(n11761), .B(n11760), .Z(n11756) );
  XOR U16064 ( .A(n11753), .B(n11762), .Z(N29179) );
  XOR U16065 ( .A(n11751), .B(n11755), .Z(n11762) );
  XNOR U16066 ( .A(n11748), .B(n11763), .Z(n11755) );
  XNOR U16067 ( .A(n11745), .B(n11747), .Z(n11763) );
  AND U16068 ( .A(n11764), .B(n11765), .Z(n11747) );
  NANDN U16069 ( .A(n11766), .B(n11767), .Z(n11765) );
  NANDN U16070 ( .A(n11768), .B(n11769), .Z(n11767) );
  IV U16071 ( .A(n11770), .Z(n11769) );
  NAND U16072 ( .A(n11770), .B(n11768), .Z(n11764) );
  AND U16073 ( .A(n11771), .B(n11772), .Z(n11745) );
  NAND U16074 ( .A(n11773), .B(n11774), .Z(n11772) );
  OR U16075 ( .A(n11775), .B(n11776), .Z(n11774) );
  NAND U16076 ( .A(n11776), .B(n11775), .Z(n11771) );
  IV U16077 ( .A(n11777), .Z(n11776) );
  NAND U16078 ( .A(n11778), .B(n11779), .Z(n11748) );
  NANDN U16079 ( .A(n11780), .B(n11781), .Z(n11779) );
  NAND U16080 ( .A(n11782), .B(n11783), .Z(n11781) );
  OR U16081 ( .A(n11783), .B(n11782), .Z(n11778) );
  IV U16082 ( .A(n11784), .Z(n11782) );
  AND U16083 ( .A(n11785), .B(n11786), .Z(n11751) );
  NAND U16084 ( .A(n11787), .B(n11788), .Z(n11786) );
  NANDN U16085 ( .A(n11789), .B(n11790), .Z(n11788) );
  NANDN U16086 ( .A(n11790), .B(n11789), .Z(n11785) );
  XOR U16087 ( .A(n11761), .B(n11791), .Z(n11753) );
  XNOR U16088 ( .A(n11758), .B(n11760), .Z(n11791) );
  AND U16089 ( .A(n11792), .B(n11793), .Z(n11760) );
  NANDN U16090 ( .A(n11794), .B(n11795), .Z(n11793) );
  NANDN U16091 ( .A(n11796), .B(n11797), .Z(n11795) );
  IV U16092 ( .A(n11798), .Z(n11797) );
  NAND U16093 ( .A(n11798), .B(n11796), .Z(n11792) );
  AND U16094 ( .A(n11799), .B(n11800), .Z(n11758) );
  NAND U16095 ( .A(n11801), .B(n11802), .Z(n11800) );
  OR U16096 ( .A(n11803), .B(n11804), .Z(n11802) );
  NAND U16097 ( .A(n11804), .B(n11803), .Z(n11799) );
  IV U16098 ( .A(n11805), .Z(n11804) );
  NAND U16099 ( .A(n11806), .B(n11807), .Z(n11761) );
  NANDN U16100 ( .A(n11808), .B(n11809), .Z(n11807) );
  NAND U16101 ( .A(n11810), .B(n11811), .Z(n11809) );
  OR U16102 ( .A(n11811), .B(n11810), .Z(n11806) );
  IV U16103 ( .A(n11812), .Z(n11810) );
  XOR U16104 ( .A(n11787), .B(n11813), .Z(N29178) );
  XNOR U16105 ( .A(n11790), .B(n11789), .Z(n11813) );
  XNOR U16106 ( .A(n11801), .B(n11814), .Z(n11789) );
  XOR U16107 ( .A(n11805), .B(n11803), .Z(n11814) );
  XOR U16108 ( .A(n11811), .B(n11815), .Z(n11803) );
  XOR U16109 ( .A(n11808), .B(n11812), .Z(n11815) );
  NAND U16110 ( .A(n11816), .B(n11817), .Z(n11812) );
  NAND U16111 ( .A(n11818), .B(n11819), .Z(n11817) );
  NAND U16112 ( .A(n11820), .B(n11821), .Z(n11816) );
  AND U16113 ( .A(n11822), .B(n11823), .Z(n11808) );
  NAND U16114 ( .A(n11824), .B(n11825), .Z(n11823) );
  NAND U16115 ( .A(n11826), .B(n11827), .Z(n11822) );
  NANDN U16116 ( .A(n11828), .B(n11829), .Z(n11811) );
  NANDN U16117 ( .A(n11830), .B(n11831), .Z(n11805) );
  XNOR U16118 ( .A(n11796), .B(n11832), .Z(n11801) );
  XOR U16119 ( .A(n11794), .B(n11798), .Z(n11832) );
  NAND U16120 ( .A(n11833), .B(n11834), .Z(n11798) );
  NAND U16121 ( .A(n11835), .B(n11836), .Z(n11834) );
  NAND U16122 ( .A(n11837), .B(n11838), .Z(n11833) );
  AND U16123 ( .A(n11839), .B(n11840), .Z(n11794) );
  NAND U16124 ( .A(n11841), .B(n11842), .Z(n11840) );
  NAND U16125 ( .A(n11843), .B(n11844), .Z(n11839) );
  AND U16126 ( .A(n11845), .B(n11846), .Z(n11796) );
  NAND U16127 ( .A(n11847), .B(n11848), .Z(n11790) );
  XNOR U16128 ( .A(n11773), .B(n11849), .Z(n11787) );
  XOR U16129 ( .A(n11777), .B(n11775), .Z(n11849) );
  XOR U16130 ( .A(n11783), .B(n11850), .Z(n11775) );
  XOR U16131 ( .A(n11780), .B(n11784), .Z(n11850) );
  NAND U16132 ( .A(n11851), .B(n11852), .Z(n11784) );
  NAND U16133 ( .A(n11853), .B(n11854), .Z(n11852) );
  NAND U16134 ( .A(n11855), .B(n11856), .Z(n11851) );
  AND U16135 ( .A(n11857), .B(n11858), .Z(n11780) );
  NAND U16136 ( .A(n11859), .B(n11860), .Z(n11858) );
  NAND U16137 ( .A(n11861), .B(n11862), .Z(n11857) );
  NANDN U16138 ( .A(n11863), .B(n11864), .Z(n11783) );
  NANDN U16139 ( .A(n11865), .B(n11866), .Z(n11777) );
  XNOR U16140 ( .A(n11768), .B(n11867), .Z(n11773) );
  XOR U16141 ( .A(n11766), .B(n11770), .Z(n11867) );
  NAND U16142 ( .A(n11868), .B(n11869), .Z(n11770) );
  NAND U16143 ( .A(n11870), .B(n11871), .Z(n11869) );
  NAND U16144 ( .A(n11872), .B(n11873), .Z(n11868) );
  AND U16145 ( .A(n11874), .B(n11875), .Z(n11766) );
  NAND U16146 ( .A(n11876), .B(n11877), .Z(n11875) );
  NAND U16147 ( .A(n11878), .B(n11879), .Z(n11874) );
  AND U16148 ( .A(n11880), .B(n11881), .Z(n11768) );
  XOR U16149 ( .A(n11848), .B(n11847), .Z(N29177) );
  XNOR U16150 ( .A(n11866), .B(n11865), .Z(n11847) );
  XNOR U16151 ( .A(n11880), .B(n11881), .Z(n11865) );
  XOR U16152 ( .A(n11877), .B(n11876), .Z(n11881) );
  XOR U16153 ( .A(y[2499]), .B(x[2499]), .Z(n11876) );
  XOR U16154 ( .A(n11879), .B(n11878), .Z(n11877) );
  XOR U16155 ( .A(y[2501]), .B(x[2501]), .Z(n11878) );
  XOR U16156 ( .A(y[2500]), .B(x[2500]), .Z(n11879) );
  XOR U16157 ( .A(n11871), .B(n11870), .Z(n11880) );
  XOR U16158 ( .A(n11873), .B(n11872), .Z(n11870) );
  XOR U16159 ( .A(y[2498]), .B(x[2498]), .Z(n11872) );
  XOR U16160 ( .A(y[2497]), .B(x[2497]), .Z(n11873) );
  XOR U16161 ( .A(y[2496]), .B(x[2496]), .Z(n11871) );
  XNOR U16162 ( .A(n11864), .B(n11863), .Z(n11866) );
  XNOR U16163 ( .A(n11860), .B(n11859), .Z(n11863) );
  XOR U16164 ( .A(n11862), .B(n11861), .Z(n11859) );
  XOR U16165 ( .A(y[2495]), .B(x[2495]), .Z(n11861) );
  XOR U16166 ( .A(y[2494]), .B(x[2494]), .Z(n11862) );
  XOR U16167 ( .A(y[2493]), .B(x[2493]), .Z(n11860) );
  XOR U16168 ( .A(n11854), .B(n11853), .Z(n11864) );
  XOR U16169 ( .A(n11856), .B(n11855), .Z(n11853) );
  XOR U16170 ( .A(y[2492]), .B(x[2492]), .Z(n11855) );
  XOR U16171 ( .A(y[2491]), .B(x[2491]), .Z(n11856) );
  XOR U16172 ( .A(y[2490]), .B(x[2490]), .Z(n11854) );
  XNOR U16173 ( .A(n11831), .B(n11830), .Z(n11848) );
  XNOR U16174 ( .A(n11845), .B(n11846), .Z(n11830) );
  XOR U16175 ( .A(n11842), .B(n11841), .Z(n11846) );
  XOR U16176 ( .A(y[2487]), .B(x[2487]), .Z(n11841) );
  XOR U16177 ( .A(n11844), .B(n11843), .Z(n11842) );
  XOR U16178 ( .A(y[2489]), .B(x[2489]), .Z(n11843) );
  XOR U16179 ( .A(y[2488]), .B(x[2488]), .Z(n11844) );
  XOR U16180 ( .A(n11836), .B(n11835), .Z(n11845) );
  XOR U16181 ( .A(n11838), .B(n11837), .Z(n11835) );
  XOR U16182 ( .A(y[2486]), .B(x[2486]), .Z(n11837) );
  XOR U16183 ( .A(y[2485]), .B(x[2485]), .Z(n11838) );
  XOR U16184 ( .A(y[2484]), .B(x[2484]), .Z(n11836) );
  XNOR U16185 ( .A(n11829), .B(n11828), .Z(n11831) );
  XNOR U16186 ( .A(n11825), .B(n11824), .Z(n11828) );
  XOR U16187 ( .A(n11827), .B(n11826), .Z(n11824) );
  XOR U16188 ( .A(y[2483]), .B(x[2483]), .Z(n11826) );
  XOR U16189 ( .A(y[2482]), .B(x[2482]), .Z(n11827) );
  XOR U16190 ( .A(y[2481]), .B(x[2481]), .Z(n11825) );
  XOR U16191 ( .A(n11819), .B(n11818), .Z(n11829) );
  XOR U16192 ( .A(n11821), .B(n11820), .Z(n11818) );
  XOR U16193 ( .A(y[2480]), .B(x[2480]), .Z(n11820) );
  XOR U16194 ( .A(y[2479]), .B(x[2479]), .Z(n11821) );
  XOR U16195 ( .A(y[2478]), .B(x[2478]), .Z(n11819) );
  NAND U16196 ( .A(n11882), .B(n11883), .Z(N29169) );
  NAND U16197 ( .A(n11884), .B(n11885), .Z(n11883) );
  NANDN U16198 ( .A(n11886), .B(n11887), .Z(n11885) );
  NANDN U16199 ( .A(n11887), .B(n11886), .Z(n11882) );
  XOR U16200 ( .A(n11886), .B(n11888), .Z(N29168) );
  XNOR U16201 ( .A(n11884), .B(n11887), .Z(n11888) );
  NAND U16202 ( .A(n11889), .B(n11890), .Z(n11887) );
  NAND U16203 ( .A(n11891), .B(n11892), .Z(n11890) );
  NANDN U16204 ( .A(n11893), .B(n11894), .Z(n11892) );
  NANDN U16205 ( .A(n11894), .B(n11893), .Z(n11889) );
  AND U16206 ( .A(n11895), .B(n11896), .Z(n11884) );
  NAND U16207 ( .A(n11897), .B(n11898), .Z(n11896) );
  OR U16208 ( .A(n11899), .B(n11900), .Z(n11898) );
  NAND U16209 ( .A(n11900), .B(n11899), .Z(n11895) );
  IV U16210 ( .A(n11901), .Z(n11900) );
  AND U16211 ( .A(n11902), .B(n11903), .Z(n11886) );
  NAND U16212 ( .A(n11904), .B(n11905), .Z(n11903) );
  NANDN U16213 ( .A(n11906), .B(n11907), .Z(n11905) );
  NANDN U16214 ( .A(n11907), .B(n11906), .Z(n11902) );
  XOR U16215 ( .A(n11899), .B(n11908), .Z(N29167) );
  XOR U16216 ( .A(n11897), .B(n11901), .Z(n11908) );
  XNOR U16217 ( .A(n11894), .B(n11909), .Z(n11901) );
  XNOR U16218 ( .A(n11891), .B(n11893), .Z(n11909) );
  AND U16219 ( .A(n11910), .B(n11911), .Z(n11893) );
  NANDN U16220 ( .A(n11912), .B(n11913), .Z(n11911) );
  NANDN U16221 ( .A(n11914), .B(n11915), .Z(n11913) );
  IV U16222 ( .A(n11916), .Z(n11915) );
  NAND U16223 ( .A(n11916), .B(n11914), .Z(n11910) );
  AND U16224 ( .A(n11917), .B(n11918), .Z(n11891) );
  NAND U16225 ( .A(n11919), .B(n11920), .Z(n11918) );
  OR U16226 ( .A(n11921), .B(n11922), .Z(n11920) );
  NAND U16227 ( .A(n11922), .B(n11921), .Z(n11917) );
  IV U16228 ( .A(n11923), .Z(n11922) );
  NAND U16229 ( .A(n11924), .B(n11925), .Z(n11894) );
  NANDN U16230 ( .A(n11926), .B(n11927), .Z(n11925) );
  NAND U16231 ( .A(n11928), .B(n11929), .Z(n11927) );
  OR U16232 ( .A(n11929), .B(n11928), .Z(n11924) );
  IV U16233 ( .A(n11930), .Z(n11928) );
  AND U16234 ( .A(n11931), .B(n11932), .Z(n11897) );
  NAND U16235 ( .A(n11933), .B(n11934), .Z(n11932) );
  NANDN U16236 ( .A(n11935), .B(n11936), .Z(n11934) );
  NANDN U16237 ( .A(n11936), .B(n11935), .Z(n11931) );
  XOR U16238 ( .A(n11907), .B(n11937), .Z(n11899) );
  XNOR U16239 ( .A(n11904), .B(n11906), .Z(n11937) );
  AND U16240 ( .A(n11938), .B(n11939), .Z(n11906) );
  NANDN U16241 ( .A(n11940), .B(n11941), .Z(n11939) );
  NANDN U16242 ( .A(n11942), .B(n11943), .Z(n11941) );
  IV U16243 ( .A(n11944), .Z(n11943) );
  NAND U16244 ( .A(n11944), .B(n11942), .Z(n11938) );
  AND U16245 ( .A(n11945), .B(n11946), .Z(n11904) );
  NAND U16246 ( .A(n11947), .B(n11948), .Z(n11946) );
  OR U16247 ( .A(n11949), .B(n11950), .Z(n11948) );
  NAND U16248 ( .A(n11950), .B(n11949), .Z(n11945) );
  IV U16249 ( .A(n11951), .Z(n11950) );
  NAND U16250 ( .A(n11952), .B(n11953), .Z(n11907) );
  NANDN U16251 ( .A(n11954), .B(n11955), .Z(n11953) );
  NAND U16252 ( .A(n11956), .B(n11957), .Z(n11955) );
  OR U16253 ( .A(n11957), .B(n11956), .Z(n11952) );
  IV U16254 ( .A(n11958), .Z(n11956) );
  XOR U16255 ( .A(n11933), .B(n11959), .Z(N29166) );
  XNOR U16256 ( .A(n11936), .B(n11935), .Z(n11959) );
  XNOR U16257 ( .A(n11947), .B(n11960), .Z(n11935) );
  XOR U16258 ( .A(n11951), .B(n11949), .Z(n11960) );
  XOR U16259 ( .A(n11957), .B(n11961), .Z(n11949) );
  XOR U16260 ( .A(n11954), .B(n11958), .Z(n11961) );
  NAND U16261 ( .A(n11962), .B(n11963), .Z(n11958) );
  NAND U16262 ( .A(n11964), .B(n11965), .Z(n11963) );
  NAND U16263 ( .A(n11966), .B(n11967), .Z(n11962) );
  AND U16264 ( .A(n11968), .B(n11969), .Z(n11954) );
  NAND U16265 ( .A(n11970), .B(n11971), .Z(n11969) );
  NAND U16266 ( .A(n11972), .B(n11973), .Z(n11968) );
  NANDN U16267 ( .A(n11974), .B(n11975), .Z(n11957) );
  NANDN U16268 ( .A(n11976), .B(n11977), .Z(n11951) );
  XNOR U16269 ( .A(n11942), .B(n11978), .Z(n11947) );
  XOR U16270 ( .A(n11940), .B(n11944), .Z(n11978) );
  NAND U16271 ( .A(n11979), .B(n11980), .Z(n11944) );
  NAND U16272 ( .A(n11981), .B(n11982), .Z(n11980) );
  NAND U16273 ( .A(n11983), .B(n11984), .Z(n11979) );
  AND U16274 ( .A(n11985), .B(n11986), .Z(n11940) );
  NAND U16275 ( .A(n11987), .B(n11988), .Z(n11986) );
  NAND U16276 ( .A(n11989), .B(n11990), .Z(n11985) );
  AND U16277 ( .A(n11991), .B(n11992), .Z(n11942) );
  NAND U16278 ( .A(n11993), .B(n11994), .Z(n11936) );
  XNOR U16279 ( .A(n11919), .B(n11995), .Z(n11933) );
  XOR U16280 ( .A(n11923), .B(n11921), .Z(n11995) );
  XOR U16281 ( .A(n11929), .B(n11996), .Z(n11921) );
  XOR U16282 ( .A(n11926), .B(n11930), .Z(n11996) );
  NAND U16283 ( .A(n11997), .B(n11998), .Z(n11930) );
  NAND U16284 ( .A(n11999), .B(n12000), .Z(n11998) );
  NAND U16285 ( .A(n12001), .B(n12002), .Z(n11997) );
  AND U16286 ( .A(n12003), .B(n12004), .Z(n11926) );
  NAND U16287 ( .A(n12005), .B(n12006), .Z(n12004) );
  NAND U16288 ( .A(n12007), .B(n12008), .Z(n12003) );
  NANDN U16289 ( .A(n12009), .B(n12010), .Z(n11929) );
  NANDN U16290 ( .A(n12011), .B(n12012), .Z(n11923) );
  XNOR U16291 ( .A(n11914), .B(n12013), .Z(n11919) );
  XOR U16292 ( .A(n11912), .B(n11916), .Z(n12013) );
  NAND U16293 ( .A(n12014), .B(n12015), .Z(n11916) );
  NAND U16294 ( .A(n12016), .B(n12017), .Z(n12015) );
  NAND U16295 ( .A(n12018), .B(n12019), .Z(n12014) );
  AND U16296 ( .A(n12020), .B(n12021), .Z(n11912) );
  NAND U16297 ( .A(n12022), .B(n12023), .Z(n12021) );
  NAND U16298 ( .A(n12024), .B(n12025), .Z(n12020) );
  AND U16299 ( .A(n12026), .B(n12027), .Z(n11914) );
  XOR U16300 ( .A(n11994), .B(n11993), .Z(N29165) );
  XNOR U16301 ( .A(n12012), .B(n12011), .Z(n11993) );
  XNOR U16302 ( .A(n12026), .B(n12027), .Z(n12011) );
  XOR U16303 ( .A(n12023), .B(n12022), .Z(n12027) );
  XOR U16304 ( .A(y[2475]), .B(x[2475]), .Z(n12022) );
  XOR U16305 ( .A(n12025), .B(n12024), .Z(n12023) );
  XOR U16306 ( .A(y[2477]), .B(x[2477]), .Z(n12024) );
  XOR U16307 ( .A(y[2476]), .B(x[2476]), .Z(n12025) );
  XOR U16308 ( .A(n12017), .B(n12016), .Z(n12026) );
  XOR U16309 ( .A(n12019), .B(n12018), .Z(n12016) );
  XOR U16310 ( .A(y[2474]), .B(x[2474]), .Z(n12018) );
  XOR U16311 ( .A(y[2473]), .B(x[2473]), .Z(n12019) );
  XOR U16312 ( .A(y[2472]), .B(x[2472]), .Z(n12017) );
  XNOR U16313 ( .A(n12010), .B(n12009), .Z(n12012) );
  XNOR U16314 ( .A(n12006), .B(n12005), .Z(n12009) );
  XOR U16315 ( .A(n12008), .B(n12007), .Z(n12005) );
  XOR U16316 ( .A(y[2471]), .B(x[2471]), .Z(n12007) );
  XOR U16317 ( .A(y[2470]), .B(x[2470]), .Z(n12008) );
  XOR U16318 ( .A(y[2469]), .B(x[2469]), .Z(n12006) );
  XOR U16319 ( .A(n12000), .B(n11999), .Z(n12010) );
  XOR U16320 ( .A(n12002), .B(n12001), .Z(n11999) );
  XOR U16321 ( .A(y[2468]), .B(x[2468]), .Z(n12001) );
  XOR U16322 ( .A(y[2467]), .B(x[2467]), .Z(n12002) );
  XOR U16323 ( .A(y[2466]), .B(x[2466]), .Z(n12000) );
  XNOR U16324 ( .A(n11977), .B(n11976), .Z(n11994) );
  XNOR U16325 ( .A(n11991), .B(n11992), .Z(n11976) );
  XOR U16326 ( .A(n11988), .B(n11987), .Z(n11992) );
  XOR U16327 ( .A(y[2463]), .B(x[2463]), .Z(n11987) );
  XOR U16328 ( .A(n11990), .B(n11989), .Z(n11988) );
  XOR U16329 ( .A(y[2465]), .B(x[2465]), .Z(n11989) );
  XOR U16330 ( .A(y[2464]), .B(x[2464]), .Z(n11990) );
  XOR U16331 ( .A(n11982), .B(n11981), .Z(n11991) );
  XOR U16332 ( .A(n11984), .B(n11983), .Z(n11981) );
  XOR U16333 ( .A(y[2462]), .B(x[2462]), .Z(n11983) );
  XOR U16334 ( .A(y[2461]), .B(x[2461]), .Z(n11984) );
  XOR U16335 ( .A(y[2460]), .B(x[2460]), .Z(n11982) );
  XNOR U16336 ( .A(n11975), .B(n11974), .Z(n11977) );
  XNOR U16337 ( .A(n11971), .B(n11970), .Z(n11974) );
  XOR U16338 ( .A(n11973), .B(n11972), .Z(n11970) );
  XOR U16339 ( .A(y[2459]), .B(x[2459]), .Z(n11972) );
  XOR U16340 ( .A(y[2458]), .B(x[2458]), .Z(n11973) );
  XOR U16341 ( .A(y[2457]), .B(x[2457]), .Z(n11971) );
  XOR U16342 ( .A(n11965), .B(n11964), .Z(n11975) );
  XOR U16343 ( .A(n11967), .B(n11966), .Z(n11964) );
  XOR U16344 ( .A(y[2456]), .B(x[2456]), .Z(n11966) );
  XOR U16345 ( .A(y[2455]), .B(x[2455]), .Z(n11967) );
  XOR U16346 ( .A(y[2454]), .B(x[2454]), .Z(n11965) );
  NAND U16347 ( .A(n12028), .B(n12029), .Z(N29157) );
  NAND U16348 ( .A(n12030), .B(n12031), .Z(n12029) );
  NANDN U16349 ( .A(n12032), .B(n12033), .Z(n12031) );
  NANDN U16350 ( .A(n12033), .B(n12032), .Z(n12028) );
  XOR U16351 ( .A(n12032), .B(n12034), .Z(N29156) );
  XNOR U16352 ( .A(n12030), .B(n12033), .Z(n12034) );
  NAND U16353 ( .A(n12035), .B(n12036), .Z(n12033) );
  NAND U16354 ( .A(n12037), .B(n12038), .Z(n12036) );
  NANDN U16355 ( .A(n12039), .B(n12040), .Z(n12038) );
  NANDN U16356 ( .A(n12040), .B(n12039), .Z(n12035) );
  AND U16357 ( .A(n12041), .B(n12042), .Z(n12030) );
  NAND U16358 ( .A(n12043), .B(n12044), .Z(n12042) );
  OR U16359 ( .A(n12045), .B(n12046), .Z(n12044) );
  NAND U16360 ( .A(n12046), .B(n12045), .Z(n12041) );
  IV U16361 ( .A(n12047), .Z(n12046) );
  AND U16362 ( .A(n12048), .B(n12049), .Z(n12032) );
  NAND U16363 ( .A(n12050), .B(n12051), .Z(n12049) );
  NANDN U16364 ( .A(n12052), .B(n12053), .Z(n12051) );
  NANDN U16365 ( .A(n12053), .B(n12052), .Z(n12048) );
  XOR U16366 ( .A(n12045), .B(n12054), .Z(N29155) );
  XOR U16367 ( .A(n12043), .B(n12047), .Z(n12054) );
  XNOR U16368 ( .A(n12040), .B(n12055), .Z(n12047) );
  XNOR U16369 ( .A(n12037), .B(n12039), .Z(n12055) );
  AND U16370 ( .A(n12056), .B(n12057), .Z(n12039) );
  NANDN U16371 ( .A(n12058), .B(n12059), .Z(n12057) );
  NANDN U16372 ( .A(n12060), .B(n12061), .Z(n12059) );
  IV U16373 ( .A(n12062), .Z(n12061) );
  NAND U16374 ( .A(n12062), .B(n12060), .Z(n12056) );
  AND U16375 ( .A(n12063), .B(n12064), .Z(n12037) );
  NAND U16376 ( .A(n12065), .B(n12066), .Z(n12064) );
  OR U16377 ( .A(n12067), .B(n12068), .Z(n12066) );
  NAND U16378 ( .A(n12068), .B(n12067), .Z(n12063) );
  IV U16379 ( .A(n12069), .Z(n12068) );
  NAND U16380 ( .A(n12070), .B(n12071), .Z(n12040) );
  NANDN U16381 ( .A(n12072), .B(n12073), .Z(n12071) );
  NAND U16382 ( .A(n12074), .B(n12075), .Z(n12073) );
  OR U16383 ( .A(n12075), .B(n12074), .Z(n12070) );
  IV U16384 ( .A(n12076), .Z(n12074) );
  AND U16385 ( .A(n12077), .B(n12078), .Z(n12043) );
  NAND U16386 ( .A(n12079), .B(n12080), .Z(n12078) );
  NANDN U16387 ( .A(n12081), .B(n12082), .Z(n12080) );
  NANDN U16388 ( .A(n12082), .B(n12081), .Z(n12077) );
  XOR U16389 ( .A(n12053), .B(n12083), .Z(n12045) );
  XNOR U16390 ( .A(n12050), .B(n12052), .Z(n12083) );
  AND U16391 ( .A(n12084), .B(n12085), .Z(n12052) );
  NANDN U16392 ( .A(n12086), .B(n12087), .Z(n12085) );
  NANDN U16393 ( .A(n12088), .B(n12089), .Z(n12087) );
  IV U16394 ( .A(n12090), .Z(n12089) );
  NAND U16395 ( .A(n12090), .B(n12088), .Z(n12084) );
  AND U16396 ( .A(n12091), .B(n12092), .Z(n12050) );
  NAND U16397 ( .A(n12093), .B(n12094), .Z(n12092) );
  OR U16398 ( .A(n12095), .B(n12096), .Z(n12094) );
  NAND U16399 ( .A(n12096), .B(n12095), .Z(n12091) );
  IV U16400 ( .A(n12097), .Z(n12096) );
  NAND U16401 ( .A(n12098), .B(n12099), .Z(n12053) );
  NANDN U16402 ( .A(n12100), .B(n12101), .Z(n12099) );
  NAND U16403 ( .A(n12102), .B(n12103), .Z(n12101) );
  OR U16404 ( .A(n12103), .B(n12102), .Z(n12098) );
  IV U16405 ( .A(n12104), .Z(n12102) );
  XOR U16406 ( .A(n12079), .B(n12105), .Z(N29154) );
  XNOR U16407 ( .A(n12082), .B(n12081), .Z(n12105) );
  XNOR U16408 ( .A(n12093), .B(n12106), .Z(n12081) );
  XOR U16409 ( .A(n12097), .B(n12095), .Z(n12106) );
  XOR U16410 ( .A(n12103), .B(n12107), .Z(n12095) );
  XOR U16411 ( .A(n12100), .B(n12104), .Z(n12107) );
  NAND U16412 ( .A(n12108), .B(n12109), .Z(n12104) );
  NAND U16413 ( .A(n12110), .B(n12111), .Z(n12109) );
  NAND U16414 ( .A(n12112), .B(n12113), .Z(n12108) );
  AND U16415 ( .A(n12114), .B(n12115), .Z(n12100) );
  NAND U16416 ( .A(n12116), .B(n12117), .Z(n12115) );
  NAND U16417 ( .A(n12118), .B(n12119), .Z(n12114) );
  NANDN U16418 ( .A(n12120), .B(n12121), .Z(n12103) );
  NANDN U16419 ( .A(n12122), .B(n12123), .Z(n12097) );
  XNOR U16420 ( .A(n12088), .B(n12124), .Z(n12093) );
  XOR U16421 ( .A(n12086), .B(n12090), .Z(n12124) );
  NAND U16422 ( .A(n12125), .B(n12126), .Z(n12090) );
  NAND U16423 ( .A(n12127), .B(n12128), .Z(n12126) );
  NAND U16424 ( .A(n12129), .B(n12130), .Z(n12125) );
  AND U16425 ( .A(n12131), .B(n12132), .Z(n12086) );
  NAND U16426 ( .A(n12133), .B(n12134), .Z(n12132) );
  NAND U16427 ( .A(n12135), .B(n12136), .Z(n12131) );
  AND U16428 ( .A(n12137), .B(n12138), .Z(n12088) );
  NAND U16429 ( .A(n12139), .B(n12140), .Z(n12082) );
  XNOR U16430 ( .A(n12065), .B(n12141), .Z(n12079) );
  XOR U16431 ( .A(n12069), .B(n12067), .Z(n12141) );
  XOR U16432 ( .A(n12075), .B(n12142), .Z(n12067) );
  XOR U16433 ( .A(n12072), .B(n12076), .Z(n12142) );
  NAND U16434 ( .A(n12143), .B(n12144), .Z(n12076) );
  NAND U16435 ( .A(n12145), .B(n12146), .Z(n12144) );
  NAND U16436 ( .A(n12147), .B(n12148), .Z(n12143) );
  AND U16437 ( .A(n12149), .B(n12150), .Z(n12072) );
  NAND U16438 ( .A(n12151), .B(n12152), .Z(n12150) );
  NAND U16439 ( .A(n12153), .B(n12154), .Z(n12149) );
  NANDN U16440 ( .A(n12155), .B(n12156), .Z(n12075) );
  NANDN U16441 ( .A(n12157), .B(n12158), .Z(n12069) );
  XNOR U16442 ( .A(n12060), .B(n12159), .Z(n12065) );
  XOR U16443 ( .A(n12058), .B(n12062), .Z(n12159) );
  NAND U16444 ( .A(n12160), .B(n12161), .Z(n12062) );
  NAND U16445 ( .A(n12162), .B(n12163), .Z(n12161) );
  NAND U16446 ( .A(n12164), .B(n12165), .Z(n12160) );
  AND U16447 ( .A(n12166), .B(n12167), .Z(n12058) );
  NAND U16448 ( .A(n12168), .B(n12169), .Z(n12167) );
  NAND U16449 ( .A(n12170), .B(n12171), .Z(n12166) );
  AND U16450 ( .A(n12172), .B(n12173), .Z(n12060) );
  XOR U16451 ( .A(n12140), .B(n12139), .Z(N29153) );
  XNOR U16452 ( .A(n12158), .B(n12157), .Z(n12139) );
  XNOR U16453 ( .A(n12172), .B(n12173), .Z(n12157) );
  XOR U16454 ( .A(n12169), .B(n12168), .Z(n12173) );
  XOR U16455 ( .A(y[2451]), .B(x[2451]), .Z(n12168) );
  XOR U16456 ( .A(n12171), .B(n12170), .Z(n12169) );
  XOR U16457 ( .A(y[2453]), .B(x[2453]), .Z(n12170) );
  XOR U16458 ( .A(y[2452]), .B(x[2452]), .Z(n12171) );
  XOR U16459 ( .A(n12163), .B(n12162), .Z(n12172) );
  XOR U16460 ( .A(n12165), .B(n12164), .Z(n12162) );
  XOR U16461 ( .A(y[2450]), .B(x[2450]), .Z(n12164) );
  XOR U16462 ( .A(y[2449]), .B(x[2449]), .Z(n12165) );
  XOR U16463 ( .A(y[2448]), .B(x[2448]), .Z(n12163) );
  XNOR U16464 ( .A(n12156), .B(n12155), .Z(n12158) );
  XNOR U16465 ( .A(n12152), .B(n12151), .Z(n12155) );
  XOR U16466 ( .A(n12154), .B(n12153), .Z(n12151) );
  XOR U16467 ( .A(y[2447]), .B(x[2447]), .Z(n12153) );
  XOR U16468 ( .A(y[2446]), .B(x[2446]), .Z(n12154) );
  XOR U16469 ( .A(y[2445]), .B(x[2445]), .Z(n12152) );
  XOR U16470 ( .A(n12146), .B(n12145), .Z(n12156) );
  XOR U16471 ( .A(n12148), .B(n12147), .Z(n12145) );
  XOR U16472 ( .A(y[2444]), .B(x[2444]), .Z(n12147) );
  XOR U16473 ( .A(y[2443]), .B(x[2443]), .Z(n12148) );
  XOR U16474 ( .A(y[2442]), .B(x[2442]), .Z(n12146) );
  XNOR U16475 ( .A(n12123), .B(n12122), .Z(n12140) );
  XNOR U16476 ( .A(n12137), .B(n12138), .Z(n12122) );
  XOR U16477 ( .A(n12134), .B(n12133), .Z(n12138) );
  XOR U16478 ( .A(y[2439]), .B(x[2439]), .Z(n12133) );
  XOR U16479 ( .A(n12136), .B(n12135), .Z(n12134) );
  XOR U16480 ( .A(y[2441]), .B(x[2441]), .Z(n12135) );
  XOR U16481 ( .A(y[2440]), .B(x[2440]), .Z(n12136) );
  XOR U16482 ( .A(n12128), .B(n12127), .Z(n12137) );
  XOR U16483 ( .A(n12130), .B(n12129), .Z(n12127) );
  XOR U16484 ( .A(y[2438]), .B(x[2438]), .Z(n12129) );
  XOR U16485 ( .A(y[2437]), .B(x[2437]), .Z(n12130) );
  XOR U16486 ( .A(y[2436]), .B(x[2436]), .Z(n12128) );
  XNOR U16487 ( .A(n12121), .B(n12120), .Z(n12123) );
  XNOR U16488 ( .A(n12117), .B(n12116), .Z(n12120) );
  XOR U16489 ( .A(n12119), .B(n12118), .Z(n12116) );
  XOR U16490 ( .A(y[2435]), .B(x[2435]), .Z(n12118) );
  XOR U16491 ( .A(y[2434]), .B(x[2434]), .Z(n12119) );
  XOR U16492 ( .A(y[2433]), .B(x[2433]), .Z(n12117) );
  XOR U16493 ( .A(n12111), .B(n12110), .Z(n12121) );
  XOR U16494 ( .A(n12113), .B(n12112), .Z(n12110) );
  XOR U16495 ( .A(y[2432]), .B(x[2432]), .Z(n12112) );
  XOR U16496 ( .A(y[2431]), .B(x[2431]), .Z(n12113) );
  XOR U16497 ( .A(y[2430]), .B(x[2430]), .Z(n12111) );
  NAND U16498 ( .A(n12174), .B(n12175), .Z(N29145) );
  NAND U16499 ( .A(n12176), .B(n12177), .Z(n12175) );
  NANDN U16500 ( .A(n12178), .B(n12179), .Z(n12177) );
  NANDN U16501 ( .A(n12179), .B(n12178), .Z(n12174) );
  XOR U16502 ( .A(n12178), .B(n12180), .Z(N29144) );
  XNOR U16503 ( .A(n12176), .B(n12179), .Z(n12180) );
  NAND U16504 ( .A(n12181), .B(n12182), .Z(n12179) );
  NAND U16505 ( .A(n12183), .B(n12184), .Z(n12182) );
  NANDN U16506 ( .A(n12185), .B(n12186), .Z(n12184) );
  NANDN U16507 ( .A(n12186), .B(n12185), .Z(n12181) );
  AND U16508 ( .A(n12187), .B(n12188), .Z(n12176) );
  NAND U16509 ( .A(n12189), .B(n12190), .Z(n12188) );
  OR U16510 ( .A(n12191), .B(n12192), .Z(n12190) );
  NAND U16511 ( .A(n12192), .B(n12191), .Z(n12187) );
  IV U16512 ( .A(n12193), .Z(n12192) );
  AND U16513 ( .A(n12194), .B(n12195), .Z(n12178) );
  NAND U16514 ( .A(n12196), .B(n12197), .Z(n12195) );
  NANDN U16515 ( .A(n12198), .B(n12199), .Z(n12197) );
  NANDN U16516 ( .A(n12199), .B(n12198), .Z(n12194) );
  XOR U16517 ( .A(n12191), .B(n12200), .Z(N29143) );
  XOR U16518 ( .A(n12189), .B(n12193), .Z(n12200) );
  XNOR U16519 ( .A(n12186), .B(n12201), .Z(n12193) );
  XNOR U16520 ( .A(n12183), .B(n12185), .Z(n12201) );
  AND U16521 ( .A(n12202), .B(n12203), .Z(n12185) );
  NANDN U16522 ( .A(n12204), .B(n12205), .Z(n12203) );
  NANDN U16523 ( .A(n12206), .B(n12207), .Z(n12205) );
  IV U16524 ( .A(n12208), .Z(n12207) );
  NAND U16525 ( .A(n12208), .B(n12206), .Z(n12202) );
  AND U16526 ( .A(n12209), .B(n12210), .Z(n12183) );
  NAND U16527 ( .A(n12211), .B(n12212), .Z(n12210) );
  OR U16528 ( .A(n12213), .B(n12214), .Z(n12212) );
  NAND U16529 ( .A(n12214), .B(n12213), .Z(n12209) );
  IV U16530 ( .A(n12215), .Z(n12214) );
  NAND U16531 ( .A(n12216), .B(n12217), .Z(n12186) );
  NANDN U16532 ( .A(n12218), .B(n12219), .Z(n12217) );
  NAND U16533 ( .A(n12220), .B(n12221), .Z(n12219) );
  OR U16534 ( .A(n12221), .B(n12220), .Z(n12216) );
  IV U16535 ( .A(n12222), .Z(n12220) );
  AND U16536 ( .A(n12223), .B(n12224), .Z(n12189) );
  NAND U16537 ( .A(n12225), .B(n12226), .Z(n12224) );
  NANDN U16538 ( .A(n12227), .B(n12228), .Z(n12226) );
  NANDN U16539 ( .A(n12228), .B(n12227), .Z(n12223) );
  XOR U16540 ( .A(n12199), .B(n12229), .Z(n12191) );
  XNOR U16541 ( .A(n12196), .B(n12198), .Z(n12229) );
  AND U16542 ( .A(n12230), .B(n12231), .Z(n12198) );
  NANDN U16543 ( .A(n12232), .B(n12233), .Z(n12231) );
  NANDN U16544 ( .A(n12234), .B(n12235), .Z(n12233) );
  IV U16545 ( .A(n12236), .Z(n12235) );
  NAND U16546 ( .A(n12236), .B(n12234), .Z(n12230) );
  AND U16547 ( .A(n12237), .B(n12238), .Z(n12196) );
  NAND U16548 ( .A(n12239), .B(n12240), .Z(n12238) );
  OR U16549 ( .A(n12241), .B(n12242), .Z(n12240) );
  NAND U16550 ( .A(n12242), .B(n12241), .Z(n12237) );
  IV U16551 ( .A(n12243), .Z(n12242) );
  NAND U16552 ( .A(n12244), .B(n12245), .Z(n12199) );
  NANDN U16553 ( .A(n12246), .B(n12247), .Z(n12245) );
  NAND U16554 ( .A(n12248), .B(n12249), .Z(n12247) );
  OR U16555 ( .A(n12249), .B(n12248), .Z(n12244) );
  IV U16556 ( .A(n12250), .Z(n12248) );
  XOR U16557 ( .A(n12225), .B(n12251), .Z(N29142) );
  XNOR U16558 ( .A(n12228), .B(n12227), .Z(n12251) );
  XNOR U16559 ( .A(n12239), .B(n12252), .Z(n12227) );
  XOR U16560 ( .A(n12243), .B(n12241), .Z(n12252) );
  XOR U16561 ( .A(n12249), .B(n12253), .Z(n12241) );
  XOR U16562 ( .A(n12246), .B(n12250), .Z(n12253) );
  NAND U16563 ( .A(n12254), .B(n12255), .Z(n12250) );
  NAND U16564 ( .A(n12256), .B(n12257), .Z(n12255) );
  NAND U16565 ( .A(n12258), .B(n12259), .Z(n12254) );
  AND U16566 ( .A(n12260), .B(n12261), .Z(n12246) );
  NAND U16567 ( .A(n12262), .B(n12263), .Z(n12261) );
  NAND U16568 ( .A(n12264), .B(n12265), .Z(n12260) );
  NANDN U16569 ( .A(n12266), .B(n12267), .Z(n12249) );
  NANDN U16570 ( .A(n12268), .B(n12269), .Z(n12243) );
  XNOR U16571 ( .A(n12234), .B(n12270), .Z(n12239) );
  XOR U16572 ( .A(n12232), .B(n12236), .Z(n12270) );
  NAND U16573 ( .A(n12271), .B(n12272), .Z(n12236) );
  NAND U16574 ( .A(n12273), .B(n12274), .Z(n12272) );
  NAND U16575 ( .A(n12275), .B(n12276), .Z(n12271) );
  AND U16576 ( .A(n12277), .B(n12278), .Z(n12232) );
  NAND U16577 ( .A(n12279), .B(n12280), .Z(n12278) );
  NAND U16578 ( .A(n12281), .B(n12282), .Z(n12277) );
  AND U16579 ( .A(n12283), .B(n12284), .Z(n12234) );
  NAND U16580 ( .A(n12285), .B(n12286), .Z(n12228) );
  XNOR U16581 ( .A(n12211), .B(n12287), .Z(n12225) );
  XOR U16582 ( .A(n12215), .B(n12213), .Z(n12287) );
  XOR U16583 ( .A(n12221), .B(n12288), .Z(n12213) );
  XOR U16584 ( .A(n12218), .B(n12222), .Z(n12288) );
  NAND U16585 ( .A(n12289), .B(n12290), .Z(n12222) );
  NAND U16586 ( .A(n12291), .B(n12292), .Z(n12290) );
  NAND U16587 ( .A(n12293), .B(n12294), .Z(n12289) );
  AND U16588 ( .A(n12295), .B(n12296), .Z(n12218) );
  NAND U16589 ( .A(n12297), .B(n12298), .Z(n12296) );
  NAND U16590 ( .A(n12299), .B(n12300), .Z(n12295) );
  NANDN U16591 ( .A(n12301), .B(n12302), .Z(n12221) );
  NANDN U16592 ( .A(n12303), .B(n12304), .Z(n12215) );
  XNOR U16593 ( .A(n12206), .B(n12305), .Z(n12211) );
  XOR U16594 ( .A(n12204), .B(n12208), .Z(n12305) );
  NAND U16595 ( .A(n12306), .B(n12307), .Z(n12208) );
  NAND U16596 ( .A(n12308), .B(n12309), .Z(n12307) );
  NAND U16597 ( .A(n12310), .B(n12311), .Z(n12306) );
  AND U16598 ( .A(n12312), .B(n12313), .Z(n12204) );
  NAND U16599 ( .A(n12314), .B(n12315), .Z(n12313) );
  NAND U16600 ( .A(n12316), .B(n12317), .Z(n12312) );
  AND U16601 ( .A(n12318), .B(n12319), .Z(n12206) );
  XOR U16602 ( .A(n12286), .B(n12285), .Z(N29141) );
  XNOR U16603 ( .A(n12304), .B(n12303), .Z(n12285) );
  XNOR U16604 ( .A(n12318), .B(n12319), .Z(n12303) );
  XOR U16605 ( .A(n12315), .B(n12314), .Z(n12319) );
  XOR U16606 ( .A(y[2427]), .B(x[2427]), .Z(n12314) );
  XOR U16607 ( .A(n12317), .B(n12316), .Z(n12315) );
  XOR U16608 ( .A(y[2429]), .B(x[2429]), .Z(n12316) );
  XOR U16609 ( .A(y[2428]), .B(x[2428]), .Z(n12317) );
  XOR U16610 ( .A(n12309), .B(n12308), .Z(n12318) );
  XOR U16611 ( .A(n12311), .B(n12310), .Z(n12308) );
  XOR U16612 ( .A(y[2426]), .B(x[2426]), .Z(n12310) );
  XOR U16613 ( .A(y[2425]), .B(x[2425]), .Z(n12311) );
  XOR U16614 ( .A(y[2424]), .B(x[2424]), .Z(n12309) );
  XNOR U16615 ( .A(n12302), .B(n12301), .Z(n12304) );
  XNOR U16616 ( .A(n12298), .B(n12297), .Z(n12301) );
  XOR U16617 ( .A(n12300), .B(n12299), .Z(n12297) );
  XOR U16618 ( .A(y[2423]), .B(x[2423]), .Z(n12299) );
  XOR U16619 ( .A(y[2422]), .B(x[2422]), .Z(n12300) );
  XOR U16620 ( .A(y[2421]), .B(x[2421]), .Z(n12298) );
  XOR U16621 ( .A(n12292), .B(n12291), .Z(n12302) );
  XOR U16622 ( .A(n12294), .B(n12293), .Z(n12291) );
  XOR U16623 ( .A(y[2420]), .B(x[2420]), .Z(n12293) );
  XOR U16624 ( .A(y[2419]), .B(x[2419]), .Z(n12294) );
  XOR U16625 ( .A(y[2418]), .B(x[2418]), .Z(n12292) );
  XNOR U16626 ( .A(n12269), .B(n12268), .Z(n12286) );
  XNOR U16627 ( .A(n12283), .B(n12284), .Z(n12268) );
  XOR U16628 ( .A(n12280), .B(n12279), .Z(n12284) );
  XOR U16629 ( .A(y[2415]), .B(x[2415]), .Z(n12279) );
  XOR U16630 ( .A(n12282), .B(n12281), .Z(n12280) );
  XOR U16631 ( .A(y[2417]), .B(x[2417]), .Z(n12281) );
  XOR U16632 ( .A(y[2416]), .B(x[2416]), .Z(n12282) );
  XOR U16633 ( .A(n12274), .B(n12273), .Z(n12283) );
  XOR U16634 ( .A(n12276), .B(n12275), .Z(n12273) );
  XOR U16635 ( .A(y[2414]), .B(x[2414]), .Z(n12275) );
  XOR U16636 ( .A(y[2413]), .B(x[2413]), .Z(n12276) );
  XOR U16637 ( .A(y[2412]), .B(x[2412]), .Z(n12274) );
  XNOR U16638 ( .A(n12267), .B(n12266), .Z(n12269) );
  XNOR U16639 ( .A(n12263), .B(n12262), .Z(n12266) );
  XOR U16640 ( .A(n12265), .B(n12264), .Z(n12262) );
  XOR U16641 ( .A(y[2411]), .B(x[2411]), .Z(n12264) );
  XOR U16642 ( .A(y[2410]), .B(x[2410]), .Z(n12265) );
  XOR U16643 ( .A(y[2409]), .B(x[2409]), .Z(n12263) );
  XOR U16644 ( .A(n12257), .B(n12256), .Z(n12267) );
  XOR U16645 ( .A(n12259), .B(n12258), .Z(n12256) );
  XOR U16646 ( .A(y[2408]), .B(x[2408]), .Z(n12258) );
  XOR U16647 ( .A(y[2407]), .B(x[2407]), .Z(n12259) );
  XOR U16648 ( .A(y[2406]), .B(x[2406]), .Z(n12257) );
  NAND U16649 ( .A(n12320), .B(n12321), .Z(N29133) );
  NAND U16650 ( .A(n12322), .B(n12323), .Z(n12321) );
  NANDN U16651 ( .A(n12324), .B(n12325), .Z(n12323) );
  NANDN U16652 ( .A(n12325), .B(n12324), .Z(n12320) );
  XOR U16653 ( .A(n12324), .B(n12326), .Z(N29132) );
  XNOR U16654 ( .A(n12322), .B(n12325), .Z(n12326) );
  NAND U16655 ( .A(n12327), .B(n12328), .Z(n12325) );
  NAND U16656 ( .A(n12329), .B(n12330), .Z(n12328) );
  NANDN U16657 ( .A(n12331), .B(n12332), .Z(n12330) );
  NANDN U16658 ( .A(n12332), .B(n12331), .Z(n12327) );
  AND U16659 ( .A(n12333), .B(n12334), .Z(n12322) );
  NAND U16660 ( .A(n12335), .B(n12336), .Z(n12334) );
  OR U16661 ( .A(n12337), .B(n12338), .Z(n12336) );
  NAND U16662 ( .A(n12338), .B(n12337), .Z(n12333) );
  IV U16663 ( .A(n12339), .Z(n12338) );
  AND U16664 ( .A(n12340), .B(n12341), .Z(n12324) );
  NAND U16665 ( .A(n12342), .B(n12343), .Z(n12341) );
  NANDN U16666 ( .A(n12344), .B(n12345), .Z(n12343) );
  NANDN U16667 ( .A(n12345), .B(n12344), .Z(n12340) );
  XOR U16668 ( .A(n12337), .B(n12346), .Z(N29131) );
  XOR U16669 ( .A(n12335), .B(n12339), .Z(n12346) );
  XNOR U16670 ( .A(n12332), .B(n12347), .Z(n12339) );
  XNOR U16671 ( .A(n12329), .B(n12331), .Z(n12347) );
  AND U16672 ( .A(n12348), .B(n12349), .Z(n12331) );
  NANDN U16673 ( .A(n12350), .B(n12351), .Z(n12349) );
  NANDN U16674 ( .A(n12352), .B(n12353), .Z(n12351) );
  IV U16675 ( .A(n12354), .Z(n12353) );
  NAND U16676 ( .A(n12354), .B(n12352), .Z(n12348) );
  AND U16677 ( .A(n12355), .B(n12356), .Z(n12329) );
  NAND U16678 ( .A(n12357), .B(n12358), .Z(n12356) );
  OR U16679 ( .A(n12359), .B(n12360), .Z(n12358) );
  NAND U16680 ( .A(n12360), .B(n12359), .Z(n12355) );
  IV U16681 ( .A(n12361), .Z(n12360) );
  NAND U16682 ( .A(n12362), .B(n12363), .Z(n12332) );
  NANDN U16683 ( .A(n12364), .B(n12365), .Z(n12363) );
  NAND U16684 ( .A(n12366), .B(n12367), .Z(n12365) );
  OR U16685 ( .A(n12367), .B(n12366), .Z(n12362) );
  IV U16686 ( .A(n12368), .Z(n12366) );
  AND U16687 ( .A(n12369), .B(n12370), .Z(n12335) );
  NAND U16688 ( .A(n12371), .B(n12372), .Z(n12370) );
  NANDN U16689 ( .A(n12373), .B(n12374), .Z(n12372) );
  NANDN U16690 ( .A(n12374), .B(n12373), .Z(n12369) );
  XOR U16691 ( .A(n12345), .B(n12375), .Z(n12337) );
  XNOR U16692 ( .A(n12342), .B(n12344), .Z(n12375) );
  AND U16693 ( .A(n12376), .B(n12377), .Z(n12344) );
  NANDN U16694 ( .A(n12378), .B(n12379), .Z(n12377) );
  NANDN U16695 ( .A(n12380), .B(n12381), .Z(n12379) );
  IV U16696 ( .A(n12382), .Z(n12381) );
  NAND U16697 ( .A(n12382), .B(n12380), .Z(n12376) );
  AND U16698 ( .A(n12383), .B(n12384), .Z(n12342) );
  NAND U16699 ( .A(n12385), .B(n12386), .Z(n12384) );
  OR U16700 ( .A(n12387), .B(n12388), .Z(n12386) );
  NAND U16701 ( .A(n12388), .B(n12387), .Z(n12383) );
  IV U16702 ( .A(n12389), .Z(n12388) );
  NAND U16703 ( .A(n12390), .B(n12391), .Z(n12345) );
  NANDN U16704 ( .A(n12392), .B(n12393), .Z(n12391) );
  NAND U16705 ( .A(n12394), .B(n12395), .Z(n12393) );
  OR U16706 ( .A(n12395), .B(n12394), .Z(n12390) );
  IV U16707 ( .A(n12396), .Z(n12394) );
  XOR U16708 ( .A(n12371), .B(n12397), .Z(N29130) );
  XNOR U16709 ( .A(n12374), .B(n12373), .Z(n12397) );
  XNOR U16710 ( .A(n12385), .B(n12398), .Z(n12373) );
  XOR U16711 ( .A(n12389), .B(n12387), .Z(n12398) );
  XOR U16712 ( .A(n12395), .B(n12399), .Z(n12387) );
  XOR U16713 ( .A(n12392), .B(n12396), .Z(n12399) );
  NAND U16714 ( .A(n12400), .B(n12401), .Z(n12396) );
  NAND U16715 ( .A(n12402), .B(n12403), .Z(n12401) );
  NAND U16716 ( .A(n12404), .B(n12405), .Z(n12400) );
  AND U16717 ( .A(n12406), .B(n12407), .Z(n12392) );
  NAND U16718 ( .A(n12408), .B(n12409), .Z(n12407) );
  NAND U16719 ( .A(n12410), .B(n12411), .Z(n12406) );
  NANDN U16720 ( .A(n12412), .B(n12413), .Z(n12395) );
  NANDN U16721 ( .A(n12414), .B(n12415), .Z(n12389) );
  XNOR U16722 ( .A(n12380), .B(n12416), .Z(n12385) );
  XOR U16723 ( .A(n12378), .B(n12382), .Z(n12416) );
  NAND U16724 ( .A(n12417), .B(n12418), .Z(n12382) );
  NAND U16725 ( .A(n12419), .B(n12420), .Z(n12418) );
  NAND U16726 ( .A(n12421), .B(n12422), .Z(n12417) );
  AND U16727 ( .A(n12423), .B(n12424), .Z(n12378) );
  NAND U16728 ( .A(n12425), .B(n12426), .Z(n12424) );
  NAND U16729 ( .A(n12427), .B(n12428), .Z(n12423) );
  AND U16730 ( .A(n12429), .B(n12430), .Z(n12380) );
  NAND U16731 ( .A(n12431), .B(n12432), .Z(n12374) );
  XNOR U16732 ( .A(n12357), .B(n12433), .Z(n12371) );
  XOR U16733 ( .A(n12361), .B(n12359), .Z(n12433) );
  XOR U16734 ( .A(n12367), .B(n12434), .Z(n12359) );
  XOR U16735 ( .A(n12364), .B(n12368), .Z(n12434) );
  NAND U16736 ( .A(n12435), .B(n12436), .Z(n12368) );
  NAND U16737 ( .A(n12437), .B(n12438), .Z(n12436) );
  NAND U16738 ( .A(n12439), .B(n12440), .Z(n12435) );
  AND U16739 ( .A(n12441), .B(n12442), .Z(n12364) );
  NAND U16740 ( .A(n12443), .B(n12444), .Z(n12442) );
  NAND U16741 ( .A(n12445), .B(n12446), .Z(n12441) );
  NANDN U16742 ( .A(n12447), .B(n12448), .Z(n12367) );
  NANDN U16743 ( .A(n12449), .B(n12450), .Z(n12361) );
  XNOR U16744 ( .A(n12352), .B(n12451), .Z(n12357) );
  XOR U16745 ( .A(n12350), .B(n12354), .Z(n12451) );
  NAND U16746 ( .A(n12452), .B(n12453), .Z(n12354) );
  NAND U16747 ( .A(n12454), .B(n12455), .Z(n12453) );
  NAND U16748 ( .A(n12456), .B(n12457), .Z(n12452) );
  AND U16749 ( .A(n12458), .B(n12459), .Z(n12350) );
  NAND U16750 ( .A(n12460), .B(n12461), .Z(n12459) );
  NAND U16751 ( .A(n12462), .B(n12463), .Z(n12458) );
  AND U16752 ( .A(n12464), .B(n12465), .Z(n12352) );
  XOR U16753 ( .A(n12432), .B(n12431), .Z(N29129) );
  XNOR U16754 ( .A(n12450), .B(n12449), .Z(n12431) );
  XNOR U16755 ( .A(n12464), .B(n12465), .Z(n12449) );
  XOR U16756 ( .A(n12461), .B(n12460), .Z(n12465) );
  XOR U16757 ( .A(y[2403]), .B(x[2403]), .Z(n12460) );
  XOR U16758 ( .A(n12463), .B(n12462), .Z(n12461) );
  XOR U16759 ( .A(y[2405]), .B(x[2405]), .Z(n12462) );
  XOR U16760 ( .A(y[2404]), .B(x[2404]), .Z(n12463) );
  XOR U16761 ( .A(n12455), .B(n12454), .Z(n12464) );
  XOR U16762 ( .A(n12457), .B(n12456), .Z(n12454) );
  XOR U16763 ( .A(y[2402]), .B(x[2402]), .Z(n12456) );
  XOR U16764 ( .A(y[2401]), .B(x[2401]), .Z(n12457) );
  XOR U16765 ( .A(y[2400]), .B(x[2400]), .Z(n12455) );
  XNOR U16766 ( .A(n12448), .B(n12447), .Z(n12450) );
  XNOR U16767 ( .A(n12444), .B(n12443), .Z(n12447) );
  XOR U16768 ( .A(n12446), .B(n12445), .Z(n12443) );
  XOR U16769 ( .A(y[2399]), .B(x[2399]), .Z(n12445) );
  XOR U16770 ( .A(y[2398]), .B(x[2398]), .Z(n12446) );
  XOR U16771 ( .A(y[2397]), .B(x[2397]), .Z(n12444) );
  XOR U16772 ( .A(n12438), .B(n12437), .Z(n12448) );
  XOR U16773 ( .A(n12440), .B(n12439), .Z(n12437) );
  XOR U16774 ( .A(y[2396]), .B(x[2396]), .Z(n12439) );
  XOR U16775 ( .A(y[2395]), .B(x[2395]), .Z(n12440) );
  XOR U16776 ( .A(y[2394]), .B(x[2394]), .Z(n12438) );
  XNOR U16777 ( .A(n12415), .B(n12414), .Z(n12432) );
  XNOR U16778 ( .A(n12429), .B(n12430), .Z(n12414) );
  XOR U16779 ( .A(n12426), .B(n12425), .Z(n12430) );
  XOR U16780 ( .A(y[2391]), .B(x[2391]), .Z(n12425) );
  XOR U16781 ( .A(n12428), .B(n12427), .Z(n12426) );
  XOR U16782 ( .A(y[2393]), .B(x[2393]), .Z(n12427) );
  XOR U16783 ( .A(y[2392]), .B(x[2392]), .Z(n12428) );
  XOR U16784 ( .A(n12420), .B(n12419), .Z(n12429) );
  XOR U16785 ( .A(n12422), .B(n12421), .Z(n12419) );
  XOR U16786 ( .A(y[2390]), .B(x[2390]), .Z(n12421) );
  XOR U16787 ( .A(y[2389]), .B(x[2389]), .Z(n12422) );
  XOR U16788 ( .A(y[2388]), .B(x[2388]), .Z(n12420) );
  XNOR U16789 ( .A(n12413), .B(n12412), .Z(n12415) );
  XNOR U16790 ( .A(n12409), .B(n12408), .Z(n12412) );
  XOR U16791 ( .A(n12411), .B(n12410), .Z(n12408) );
  XOR U16792 ( .A(y[2387]), .B(x[2387]), .Z(n12410) );
  XOR U16793 ( .A(y[2386]), .B(x[2386]), .Z(n12411) );
  XOR U16794 ( .A(y[2385]), .B(x[2385]), .Z(n12409) );
  XOR U16795 ( .A(n12403), .B(n12402), .Z(n12413) );
  XOR U16796 ( .A(n12405), .B(n12404), .Z(n12402) );
  XOR U16797 ( .A(y[2384]), .B(x[2384]), .Z(n12404) );
  XOR U16798 ( .A(y[2383]), .B(x[2383]), .Z(n12405) );
  XOR U16799 ( .A(y[2382]), .B(x[2382]), .Z(n12403) );
  NAND U16800 ( .A(n12466), .B(n12467), .Z(N29121) );
  NAND U16801 ( .A(n12468), .B(n12469), .Z(n12467) );
  NANDN U16802 ( .A(n12470), .B(n12471), .Z(n12469) );
  NANDN U16803 ( .A(n12471), .B(n12470), .Z(n12466) );
  XOR U16804 ( .A(n12470), .B(n12472), .Z(N29120) );
  XNOR U16805 ( .A(n12468), .B(n12471), .Z(n12472) );
  NAND U16806 ( .A(n12473), .B(n12474), .Z(n12471) );
  NAND U16807 ( .A(n12475), .B(n12476), .Z(n12474) );
  NANDN U16808 ( .A(n12477), .B(n12478), .Z(n12476) );
  NANDN U16809 ( .A(n12478), .B(n12477), .Z(n12473) );
  AND U16810 ( .A(n12479), .B(n12480), .Z(n12468) );
  NAND U16811 ( .A(n12481), .B(n12482), .Z(n12480) );
  OR U16812 ( .A(n12483), .B(n12484), .Z(n12482) );
  NAND U16813 ( .A(n12484), .B(n12483), .Z(n12479) );
  IV U16814 ( .A(n12485), .Z(n12484) );
  AND U16815 ( .A(n12486), .B(n12487), .Z(n12470) );
  NAND U16816 ( .A(n12488), .B(n12489), .Z(n12487) );
  NANDN U16817 ( .A(n12490), .B(n12491), .Z(n12489) );
  NANDN U16818 ( .A(n12491), .B(n12490), .Z(n12486) );
  XOR U16819 ( .A(n12483), .B(n12492), .Z(N29119) );
  XOR U16820 ( .A(n12481), .B(n12485), .Z(n12492) );
  XNOR U16821 ( .A(n12478), .B(n12493), .Z(n12485) );
  XNOR U16822 ( .A(n12475), .B(n12477), .Z(n12493) );
  AND U16823 ( .A(n12494), .B(n12495), .Z(n12477) );
  NANDN U16824 ( .A(n12496), .B(n12497), .Z(n12495) );
  NANDN U16825 ( .A(n12498), .B(n12499), .Z(n12497) );
  IV U16826 ( .A(n12500), .Z(n12499) );
  NAND U16827 ( .A(n12500), .B(n12498), .Z(n12494) );
  AND U16828 ( .A(n12501), .B(n12502), .Z(n12475) );
  NAND U16829 ( .A(n12503), .B(n12504), .Z(n12502) );
  OR U16830 ( .A(n12505), .B(n12506), .Z(n12504) );
  NAND U16831 ( .A(n12506), .B(n12505), .Z(n12501) );
  IV U16832 ( .A(n12507), .Z(n12506) );
  NAND U16833 ( .A(n12508), .B(n12509), .Z(n12478) );
  NANDN U16834 ( .A(n12510), .B(n12511), .Z(n12509) );
  NAND U16835 ( .A(n12512), .B(n12513), .Z(n12511) );
  OR U16836 ( .A(n12513), .B(n12512), .Z(n12508) );
  IV U16837 ( .A(n12514), .Z(n12512) );
  AND U16838 ( .A(n12515), .B(n12516), .Z(n12481) );
  NAND U16839 ( .A(n12517), .B(n12518), .Z(n12516) );
  NANDN U16840 ( .A(n12519), .B(n12520), .Z(n12518) );
  NANDN U16841 ( .A(n12520), .B(n12519), .Z(n12515) );
  XOR U16842 ( .A(n12491), .B(n12521), .Z(n12483) );
  XNOR U16843 ( .A(n12488), .B(n12490), .Z(n12521) );
  AND U16844 ( .A(n12522), .B(n12523), .Z(n12490) );
  NANDN U16845 ( .A(n12524), .B(n12525), .Z(n12523) );
  NANDN U16846 ( .A(n12526), .B(n12527), .Z(n12525) );
  IV U16847 ( .A(n12528), .Z(n12527) );
  NAND U16848 ( .A(n12528), .B(n12526), .Z(n12522) );
  AND U16849 ( .A(n12529), .B(n12530), .Z(n12488) );
  NAND U16850 ( .A(n12531), .B(n12532), .Z(n12530) );
  OR U16851 ( .A(n12533), .B(n12534), .Z(n12532) );
  NAND U16852 ( .A(n12534), .B(n12533), .Z(n12529) );
  IV U16853 ( .A(n12535), .Z(n12534) );
  NAND U16854 ( .A(n12536), .B(n12537), .Z(n12491) );
  NANDN U16855 ( .A(n12538), .B(n12539), .Z(n12537) );
  NAND U16856 ( .A(n12540), .B(n12541), .Z(n12539) );
  OR U16857 ( .A(n12541), .B(n12540), .Z(n12536) );
  IV U16858 ( .A(n12542), .Z(n12540) );
  XOR U16859 ( .A(n12517), .B(n12543), .Z(N29118) );
  XNOR U16860 ( .A(n12520), .B(n12519), .Z(n12543) );
  XNOR U16861 ( .A(n12531), .B(n12544), .Z(n12519) );
  XOR U16862 ( .A(n12535), .B(n12533), .Z(n12544) );
  XOR U16863 ( .A(n12541), .B(n12545), .Z(n12533) );
  XOR U16864 ( .A(n12538), .B(n12542), .Z(n12545) );
  NAND U16865 ( .A(n12546), .B(n12547), .Z(n12542) );
  NAND U16866 ( .A(n12548), .B(n12549), .Z(n12547) );
  NAND U16867 ( .A(n12550), .B(n12551), .Z(n12546) );
  AND U16868 ( .A(n12552), .B(n12553), .Z(n12538) );
  NAND U16869 ( .A(n12554), .B(n12555), .Z(n12553) );
  NAND U16870 ( .A(n12556), .B(n12557), .Z(n12552) );
  NANDN U16871 ( .A(n12558), .B(n12559), .Z(n12541) );
  NANDN U16872 ( .A(n12560), .B(n12561), .Z(n12535) );
  XNOR U16873 ( .A(n12526), .B(n12562), .Z(n12531) );
  XOR U16874 ( .A(n12524), .B(n12528), .Z(n12562) );
  NAND U16875 ( .A(n12563), .B(n12564), .Z(n12528) );
  NAND U16876 ( .A(n12565), .B(n12566), .Z(n12564) );
  NAND U16877 ( .A(n12567), .B(n12568), .Z(n12563) );
  AND U16878 ( .A(n12569), .B(n12570), .Z(n12524) );
  NAND U16879 ( .A(n12571), .B(n12572), .Z(n12570) );
  NAND U16880 ( .A(n12573), .B(n12574), .Z(n12569) );
  AND U16881 ( .A(n12575), .B(n12576), .Z(n12526) );
  NAND U16882 ( .A(n12577), .B(n12578), .Z(n12520) );
  XNOR U16883 ( .A(n12503), .B(n12579), .Z(n12517) );
  XOR U16884 ( .A(n12507), .B(n12505), .Z(n12579) );
  XOR U16885 ( .A(n12513), .B(n12580), .Z(n12505) );
  XOR U16886 ( .A(n12510), .B(n12514), .Z(n12580) );
  NAND U16887 ( .A(n12581), .B(n12582), .Z(n12514) );
  NAND U16888 ( .A(n12583), .B(n12584), .Z(n12582) );
  NAND U16889 ( .A(n12585), .B(n12586), .Z(n12581) );
  AND U16890 ( .A(n12587), .B(n12588), .Z(n12510) );
  NAND U16891 ( .A(n12589), .B(n12590), .Z(n12588) );
  NAND U16892 ( .A(n12591), .B(n12592), .Z(n12587) );
  NANDN U16893 ( .A(n12593), .B(n12594), .Z(n12513) );
  NANDN U16894 ( .A(n12595), .B(n12596), .Z(n12507) );
  XNOR U16895 ( .A(n12498), .B(n12597), .Z(n12503) );
  XOR U16896 ( .A(n12496), .B(n12500), .Z(n12597) );
  NAND U16897 ( .A(n12598), .B(n12599), .Z(n12500) );
  NAND U16898 ( .A(n12600), .B(n12601), .Z(n12599) );
  NAND U16899 ( .A(n12602), .B(n12603), .Z(n12598) );
  AND U16900 ( .A(n12604), .B(n12605), .Z(n12496) );
  NAND U16901 ( .A(n12606), .B(n12607), .Z(n12605) );
  NAND U16902 ( .A(n12608), .B(n12609), .Z(n12604) );
  AND U16903 ( .A(n12610), .B(n12611), .Z(n12498) );
  XOR U16904 ( .A(n12578), .B(n12577), .Z(N29117) );
  XNOR U16905 ( .A(n12596), .B(n12595), .Z(n12577) );
  XNOR U16906 ( .A(n12610), .B(n12611), .Z(n12595) );
  XOR U16907 ( .A(n12607), .B(n12606), .Z(n12611) );
  XOR U16908 ( .A(y[2379]), .B(x[2379]), .Z(n12606) );
  XOR U16909 ( .A(n12609), .B(n12608), .Z(n12607) );
  XOR U16910 ( .A(y[2381]), .B(x[2381]), .Z(n12608) );
  XOR U16911 ( .A(y[2380]), .B(x[2380]), .Z(n12609) );
  XOR U16912 ( .A(n12601), .B(n12600), .Z(n12610) );
  XOR U16913 ( .A(n12603), .B(n12602), .Z(n12600) );
  XOR U16914 ( .A(y[2378]), .B(x[2378]), .Z(n12602) );
  XOR U16915 ( .A(y[2377]), .B(x[2377]), .Z(n12603) );
  XOR U16916 ( .A(y[2376]), .B(x[2376]), .Z(n12601) );
  XNOR U16917 ( .A(n12594), .B(n12593), .Z(n12596) );
  XNOR U16918 ( .A(n12590), .B(n12589), .Z(n12593) );
  XOR U16919 ( .A(n12592), .B(n12591), .Z(n12589) );
  XOR U16920 ( .A(y[2375]), .B(x[2375]), .Z(n12591) );
  XOR U16921 ( .A(y[2374]), .B(x[2374]), .Z(n12592) );
  XOR U16922 ( .A(y[2373]), .B(x[2373]), .Z(n12590) );
  XOR U16923 ( .A(n12584), .B(n12583), .Z(n12594) );
  XOR U16924 ( .A(n12586), .B(n12585), .Z(n12583) );
  XOR U16925 ( .A(y[2372]), .B(x[2372]), .Z(n12585) );
  XOR U16926 ( .A(y[2371]), .B(x[2371]), .Z(n12586) );
  XOR U16927 ( .A(y[2370]), .B(x[2370]), .Z(n12584) );
  XNOR U16928 ( .A(n12561), .B(n12560), .Z(n12578) );
  XNOR U16929 ( .A(n12575), .B(n12576), .Z(n12560) );
  XOR U16930 ( .A(n12572), .B(n12571), .Z(n12576) );
  XOR U16931 ( .A(y[2367]), .B(x[2367]), .Z(n12571) );
  XOR U16932 ( .A(n12574), .B(n12573), .Z(n12572) );
  XOR U16933 ( .A(y[2369]), .B(x[2369]), .Z(n12573) );
  XOR U16934 ( .A(y[2368]), .B(x[2368]), .Z(n12574) );
  XOR U16935 ( .A(n12566), .B(n12565), .Z(n12575) );
  XOR U16936 ( .A(n12568), .B(n12567), .Z(n12565) );
  XOR U16937 ( .A(y[2366]), .B(x[2366]), .Z(n12567) );
  XOR U16938 ( .A(y[2365]), .B(x[2365]), .Z(n12568) );
  XOR U16939 ( .A(y[2364]), .B(x[2364]), .Z(n12566) );
  XNOR U16940 ( .A(n12559), .B(n12558), .Z(n12561) );
  XNOR U16941 ( .A(n12555), .B(n12554), .Z(n12558) );
  XOR U16942 ( .A(n12557), .B(n12556), .Z(n12554) );
  XOR U16943 ( .A(y[2363]), .B(x[2363]), .Z(n12556) );
  XOR U16944 ( .A(y[2362]), .B(x[2362]), .Z(n12557) );
  XOR U16945 ( .A(y[2361]), .B(x[2361]), .Z(n12555) );
  XOR U16946 ( .A(n12549), .B(n12548), .Z(n12559) );
  XOR U16947 ( .A(n12551), .B(n12550), .Z(n12548) );
  XOR U16948 ( .A(y[2360]), .B(x[2360]), .Z(n12550) );
  XOR U16949 ( .A(y[2359]), .B(x[2359]), .Z(n12551) );
  XOR U16950 ( .A(y[2358]), .B(x[2358]), .Z(n12549) );
  NAND U16951 ( .A(n12612), .B(n12613), .Z(N29109) );
  NAND U16952 ( .A(n12614), .B(n12615), .Z(n12613) );
  NANDN U16953 ( .A(n12616), .B(n12617), .Z(n12615) );
  NANDN U16954 ( .A(n12617), .B(n12616), .Z(n12612) );
  XOR U16955 ( .A(n12616), .B(n12618), .Z(N29108) );
  XNOR U16956 ( .A(n12614), .B(n12617), .Z(n12618) );
  NAND U16957 ( .A(n12619), .B(n12620), .Z(n12617) );
  NAND U16958 ( .A(n12621), .B(n12622), .Z(n12620) );
  NANDN U16959 ( .A(n12623), .B(n12624), .Z(n12622) );
  NANDN U16960 ( .A(n12624), .B(n12623), .Z(n12619) );
  AND U16961 ( .A(n12625), .B(n12626), .Z(n12614) );
  NAND U16962 ( .A(n12627), .B(n12628), .Z(n12626) );
  OR U16963 ( .A(n12629), .B(n12630), .Z(n12628) );
  NAND U16964 ( .A(n12630), .B(n12629), .Z(n12625) );
  IV U16965 ( .A(n12631), .Z(n12630) );
  AND U16966 ( .A(n12632), .B(n12633), .Z(n12616) );
  NAND U16967 ( .A(n12634), .B(n12635), .Z(n12633) );
  NANDN U16968 ( .A(n12636), .B(n12637), .Z(n12635) );
  NANDN U16969 ( .A(n12637), .B(n12636), .Z(n12632) );
  XOR U16970 ( .A(n12629), .B(n12638), .Z(N29107) );
  XOR U16971 ( .A(n12627), .B(n12631), .Z(n12638) );
  XNOR U16972 ( .A(n12624), .B(n12639), .Z(n12631) );
  XNOR U16973 ( .A(n12621), .B(n12623), .Z(n12639) );
  AND U16974 ( .A(n12640), .B(n12641), .Z(n12623) );
  NANDN U16975 ( .A(n12642), .B(n12643), .Z(n12641) );
  NANDN U16976 ( .A(n12644), .B(n12645), .Z(n12643) );
  IV U16977 ( .A(n12646), .Z(n12645) );
  NAND U16978 ( .A(n12646), .B(n12644), .Z(n12640) );
  AND U16979 ( .A(n12647), .B(n12648), .Z(n12621) );
  NAND U16980 ( .A(n12649), .B(n12650), .Z(n12648) );
  OR U16981 ( .A(n12651), .B(n12652), .Z(n12650) );
  NAND U16982 ( .A(n12652), .B(n12651), .Z(n12647) );
  IV U16983 ( .A(n12653), .Z(n12652) );
  NAND U16984 ( .A(n12654), .B(n12655), .Z(n12624) );
  NANDN U16985 ( .A(n12656), .B(n12657), .Z(n12655) );
  NAND U16986 ( .A(n12658), .B(n12659), .Z(n12657) );
  OR U16987 ( .A(n12659), .B(n12658), .Z(n12654) );
  IV U16988 ( .A(n12660), .Z(n12658) );
  AND U16989 ( .A(n12661), .B(n12662), .Z(n12627) );
  NAND U16990 ( .A(n12663), .B(n12664), .Z(n12662) );
  NANDN U16991 ( .A(n12665), .B(n12666), .Z(n12664) );
  NANDN U16992 ( .A(n12666), .B(n12665), .Z(n12661) );
  XOR U16993 ( .A(n12637), .B(n12667), .Z(n12629) );
  XNOR U16994 ( .A(n12634), .B(n12636), .Z(n12667) );
  AND U16995 ( .A(n12668), .B(n12669), .Z(n12636) );
  NANDN U16996 ( .A(n12670), .B(n12671), .Z(n12669) );
  NANDN U16997 ( .A(n12672), .B(n12673), .Z(n12671) );
  IV U16998 ( .A(n12674), .Z(n12673) );
  NAND U16999 ( .A(n12674), .B(n12672), .Z(n12668) );
  AND U17000 ( .A(n12675), .B(n12676), .Z(n12634) );
  NAND U17001 ( .A(n12677), .B(n12678), .Z(n12676) );
  OR U17002 ( .A(n12679), .B(n12680), .Z(n12678) );
  NAND U17003 ( .A(n12680), .B(n12679), .Z(n12675) );
  IV U17004 ( .A(n12681), .Z(n12680) );
  NAND U17005 ( .A(n12682), .B(n12683), .Z(n12637) );
  NANDN U17006 ( .A(n12684), .B(n12685), .Z(n12683) );
  NAND U17007 ( .A(n12686), .B(n12687), .Z(n12685) );
  OR U17008 ( .A(n12687), .B(n12686), .Z(n12682) );
  IV U17009 ( .A(n12688), .Z(n12686) );
  XOR U17010 ( .A(n12663), .B(n12689), .Z(N29106) );
  XNOR U17011 ( .A(n12666), .B(n12665), .Z(n12689) );
  XNOR U17012 ( .A(n12677), .B(n12690), .Z(n12665) );
  XOR U17013 ( .A(n12681), .B(n12679), .Z(n12690) );
  XOR U17014 ( .A(n12687), .B(n12691), .Z(n12679) );
  XOR U17015 ( .A(n12684), .B(n12688), .Z(n12691) );
  NAND U17016 ( .A(n12692), .B(n12693), .Z(n12688) );
  NAND U17017 ( .A(n12694), .B(n12695), .Z(n12693) );
  NAND U17018 ( .A(n12696), .B(n12697), .Z(n12692) );
  AND U17019 ( .A(n12698), .B(n12699), .Z(n12684) );
  NAND U17020 ( .A(n12700), .B(n12701), .Z(n12699) );
  NAND U17021 ( .A(n12702), .B(n12703), .Z(n12698) );
  NANDN U17022 ( .A(n12704), .B(n12705), .Z(n12687) );
  NANDN U17023 ( .A(n12706), .B(n12707), .Z(n12681) );
  XNOR U17024 ( .A(n12672), .B(n12708), .Z(n12677) );
  XOR U17025 ( .A(n12670), .B(n12674), .Z(n12708) );
  NAND U17026 ( .A(n12709), .B(n12710), .Z(n12674) );
  NAND U17027 ( .A(n12711), .B(n12712), .Z(n12710) );
  NAND U17028 ( .A(n12713), .B(n12714), .Z(n12709) );
  AND U17029 ( .A(n12715), .B(n12716), .Z(n12670) );
  NAND U17030 ( .A(n12717), .B(n12718), .Z(n12716) );
  NAND U17031 ( .A(n12719), .B(n12720), .Z(n12715) );
  AND U17032 ( .A(n12721), .B(n12722), .Z(n12672) );
  NAND U17033 ( .A(n12723), .B(n12724), .Z(n12666) );
  XNOR U17034 ( .A(n12649), .B(n12725), .Z(n12663) );
  XOR U17035 ( .A(n12653), .B(n12651), .Z(n12725) );
  XOR U17036 ( .A(n12659), .B(n12726), .Z(n12651) );
  XOR U17037 ( .A(n12656), .B(n12660), .Z(n12726) );
  NAND U17038 ( .A(n12727), .B(n12728), .Z(n12660) );
  NAND U17039 ( .A(n12729), .B(n12730), .Z(n12728) );
  NAND U17040 ( .A(n12731), .B(n12732), .Z(n12727) );
  AND U17041 ( .A(n12733), .B(n12734), .Z(n12656) );
  NAND U17042 ( .A(n12735), .B(n12736), .Z(n12734) );
  NAND U17043 ( .A(n12737), .B(n12738), .Z(n12733) );
  NANDN U17044 ( .A(n12739), .B(n12740), .Z(n12659) );
  NANDN U17045 ( .A(n12741), .B(n12742), .Z(n12653) );
  XNOR U17046 ( .A(n12644), .B(n12743), .Z(n12649) );
  XOR U17047 ( .A(n12642), .B(n12646), .Z(n12743) );
  NAND U17048 ( .A(n12744), .B(n12745), .Z(n12646) );
  NAND U17049 ( .A(n12746), .B(n12747), .Z(n12745) );
  NAND U17050 ( .A(n12748), .B(n12749), .Z(n12744) );
  AND U17051 ( .A(n12750), .B(n12751), .Z(n12642) );
  NAND U17052 ( .A(n12752), .B(n12753), .Z(n12751) );
  NAND U17053 ( .A(n12754), .B(n12755), .Z(n12750) );
  AND U17054 ( .A(n12756), .B(n12757), .Z(n12644) );
  XOR U17055 ( .A(n12724), .B(n12723), .Z(N29105) );
  XNOR U17056 ( .A(n12742), .B(n12741), .Z(n12723) );
  XNOR U17057 ( .A(n12756), .B(n12757), .Z(n12741) );
  XOR U17058 ( .A(n12753), .B(n12752), .Z(n12757) );
  XOR U17059 ( .A(y[2355]), .B(x[2355]), .Z(n12752) );
  XOR U17060 ( .A(n12755), .B(n12754), .Z(n12753) );
  XOR U17061 ( .A(y[2357]), .B(x[2357]), .Z(n12754) );
  XOR U17062 ( .A(y[2356]), .B(x[2356]), .Z(n12755) );
  XOR U17063 ( .A(n12747), .B(n12746), .Z(n12756) );
  XOR U17064 ( .A(n12749), .B(n12748), .Z(n12746) );
  XOR U17065 ( .A(y[2354]), .B(x[2354]), .Z(n12748) );
  XOR U17066 ( .A(y[2353]), .B(x[2353]), .Z(n12749) );
  XOR U17067 ( .A(y[2352]), .B(x[2352]), .Z(n12747) );
  XNOR U17068 ( .A(n12740), .B(n12739), .Z(n12742) );
  XNOR U17069 ( .A(n12736), .B(n12735), .Z(n12739) );
  XOR U17070 ( .A(n12738), .B(n12737), .Z(n12735) );
  XOR U17071 ( .A(y[2351]), .B(x[2351]), .Z(n12737) );
  XOR U17072 ( .A(y[2350]), .B(x[2350]), .Z(n12738) );
  XOR U17073 ( .A(y[2349]), .B(x[2349]), .Z(n12736) );
  XOR U17074 ( .A(n12730), .B(n12729), .Z(n12740) );
  XOR U17075 ( .A(n12732), .B(n12731), .Z(n12729) );
  XOR U17076 ( .A(y[2348]), .B(x[2348]), .Z(n12731) );
  XOR U17077 ( .A(y[2347]), .B(x[2347]), .Z(n12732) );
  XOR U17078 ( .A(y[2346]), .B(x[2346]), .Z(n12730) );
  XNOR U17079 ( .A(n12707), .B(n12706), .Z(n12724) );
  XNOR U17080 ( .A(n12721), .B(n12722), .Z(n12706) );
  XOR U17081 ( .A(n12718), .B(n12717), .Z(n12722) );
  XOR U17082 ( .A(y[2343]), .B(x[2343]), .Z(n12717) );
  XOR U17083 ( .A(n12720), .B(n12719), .Z(n12718) );
  XOR U17084 ( .A(y[2345]), .B(x[2345]), .Z(n12719) );
  XOR U17085 ( .A(y[2344]), .B(x[2344]), .Z(n12720) );
  XOR U17086 ( .A(n12712), .B(n12711), .Z(n12721) );
  XOR U17087 ( .A(n12714), .B(n12713), .Z(n12711) );
  XOR U17088 ( .A(y[2342]), .B(x[2342]), .Z(n12713) );
  XOR U17089 ( .A(y[2341]), .B(x[2341]), .Z(n12714) );
  XOR U17090 ( .A(y[2340]), .B(x[2340]), .Z(n12712) );
  XNOR U17091 ( .A(n12705), .B(n12704), .Z(n12707) );
  XNOR U17092 ( .A(n12701), .B(n12700), .Z(n12704) );
  XOR U17093 ( .A(n12703), .B(n12702), .Z(n12700) );
  XOR U17094 ( .A(y[2339]), .B(x[2339]), .Z(n12702) );
  XOR U17095 ( .A(y[2338]), .B(x[2338]), .Z(n12703) );
  XOR U17096 ( .A(y[2337]), .B(x[2337]), .Z(n12701) );
  XOR U17097 ( .A(n12695), .B(n12694), .Z(n12705) );
  XOR U17098 ( .A(n12697), .B(n12696), .Z(n12694) );
  XOR U17099 ( .A(y[2336]), .B(x[2336]), .Z(n12696) );
  XOR U17100 ( .A(y[2335]), .B(x[2335]), .Z(n12697) );
  XOR U17101 ( .A(y[2334]), .B(x[2334]), .Z(n12695) );
  NAND U17102 ( .A(n12758), .B(n12759), .Z(N29097) );
  NAND U17103 ( .A(n12760), .B(n12761), .Z(n12759) );
  NANDN U17104 ( .A(n12762), .B(n12763), .Z(n12761) );
  NANDN U17105 ( .A(n12763), .B(n12762), .Z(n12758) );
  XOR U17106 ( .A(n12762), .B(n12764), .Z(N29096) );
  XNOR U17107 ( .A(n12760), .B(n12763), .Z(n12764) );
  NAND U17108 ( .A(n12765), .B(n12766), .Z(n12763) );
  NAND U17109 ( .A(n12767), .B(n12768), .Z(n12766) );
  NANDN U17110 ( .A(n12769), .B(n12770), .Z(n12768) );
  NANDN U17111 ( .A(n12770), .B(n12769), .Z(n12765) );
  AND U17112 ( .A(n12771), .B(n12772), .Z(n12760) );
  NAND U17113 ( .A(n12773), .B(n12774), .Z(n12772) );
  OR U17114 ( .A(n12775), .B(n12776), .Z(n12774) );
  NAND U17115 ( .A(n12776), .B(n12775), .Z(n12771) );
  IV U17116 ( .A(n12777), .Z(n12776) );
  AND U17117 ( .A(n12778), .B(n12779), .Z(n12762) );
  NAND U17118 ( .A(n12780), .B(n12781), .Z(n12779) );
  NANDN U17119 ( .A(n12782), .B(n12783), .Z(n12781) );
  NANDN U17120 ( .A(n12783), .B(n12782), .Z(n12778) );
  XOR U17121 ( .A(n12775), .B(n12784), .Z(N29095) );
  XOR U17122 ( .A(n12773), .B(n12777), .Z(n12784) );
  XNOR U17123 ( .A(n12770), .B(n12785), .Z(n12777) );
  XNOR U17124 ( .A(n12767), .B(n12769), .Z(n12785) );
  AND U17125 ( .A(n12786), .B(n12787), .Z(n12769) );
  NANDN U17126 ( .A(n12788), .B(n12789), .Z(n12787) );
  NANDN U17127 ( .A(n12790), .B(n12791), .Z(n12789) );
  IV U17128 ( .A(n12792), .Z(n12791) );
  NAND U17129 ( .A(n12792), .B(n12790), .Z(n12786) );
  AND U17130 ( .A(n12793), .B(n12794), .Z(n12767) );
  NAND U17131 ( .A(n12795), .B(n12796), .Z(n12794) );
  OR U17132 ( .A(n12797), .B(n12798), .Z(n12796) );
  NAND U17133 ( .A(n12798), .B(n12797), .Z(n12793) );
  IV U17134 ( .A(n12799), .Z(n12798) );
  NAND U17135 ( .A(n12800), .B(n12801), .Z(n12770) );
  NANDN U17136 ( .A(n12802), .B(n12803), .Z(n12801) );
  NAND U17137 ( .A(n12804), .B(n12805), .Z(n12803) );
  OR U17138 ( .A(n12805), .B(n12804), .Z(n12800) );
  IV U17139 ( .A(n12806), .Z(n12804) );
  AND U17140 ( .A(n12807), .B(n12808), .Z(n12773) );
  NAND U17141 ( .A(n12809), .B(n12810), .Z(n12808) );
  NANDN U17142 ( .A(n12811), .B(n12812), .Z(n12810) );
  NANDN U17143 ( .A(n12812), .B(n12811), .Z(n12807) );
  XOR U17144 ( .A(n12783), .B(n12813), .Z(n12775) );
  XNOR U17145 ( .A(n12780), .B(n12782), .Z(n12813) );
  AND U17146 ( .A(n12814), .B(n12815), .Z(n12782) );
  NANDN U17147 ( .A(n12816), .B(n12817), .Z(n12815) );
  NANDN U17148 ( .A(n12818), .B(n12819), .Z(n12817) );
  IV U17149 ( .A(n12820), .Z(n12819) );
  NAND U17150 ( .A(n12820), .B(n12818), .Z(n12814) );
  AND U17151 ( .A(n12821), .B(n12822), .Z(n12780) );
  NAND U17152 ( .A(n12823), .B(n12824), .Z(n12822) );
  OR U17153 ( .A(n12825), .B(n12826), .Z(n12824) );
  NAND U17154 ( .A(n12826), .B(n12825), .Z(n12821) );
  IV U17155 ( .A(n12827), .Z(n12826) );
  NAND U17156 ( .A(n12828), .B(n12829), .Z(n12783) );
  NANDN U17157 ( .A(n12830), .B(n12831), .Z(n12829) );
  NAND U17158 ( .A(n12832), .B(n12833), .Z(n12831) );
  OR U17159 ( .A(n12833), .B(n12832), .Z(n12828) );
  IV U17160 ( .A(n12834), .Z(n12832) );
  XOR U17161 ( .A(n12809), .B(n12835), .Z(N29094) );
  XNOR U17162 ( .A(n12812), .B(n12811), .Z(n12835) );
  XNOR U17163 ( .A(n12823), .B(n12836), .Z(n12811) );
  XOR U17164 ( .A(n12827), .B(n12825), .Z(n12836) );
  XOR U17165 ( .A(n12833), .B(n12837), .Z(n12825) );
  XOR U17166 ( .A(n12830), .B(n12834), .Z(n12837) );
  NAND U17167 ( .A(n12838), .B(n12839), .Z(n12834) );
  NAND U17168 ( .A(n12840), .B(n12841), .Z(n12839) );
  NAND U17169 ( .A(n12842), .B(n12843), .Z(n12838) );
  AND U17170 ( .A(n12844), .B(n12845), .Z(n12830) );
  NAND U17171 ( .A(n12846), .B(n12847), .Z(n12845) );
  NAND U17172 ( .A(n12848), .B(n12849), .Z(n12844) );
  NANDN U17173 ( .A(n12850), .B(n12851), .Z(n12833) );
  NANDN U17174 ( .A(n12852), .B(n12853), .Z(n12827) );
  XNOR U17175 ( .A(n12818), .B(n12854), .Z(n12823) );
  XOR U17176 ( .A(n12816), .B(n12820), .Z(n12854) );
  NAND U17177 ( .A(n12855), .B(n12856), .Z(n12820) );
  NAND U17178 ( .A(n12857), .B(n12858), .Z(n12856) );
  NAND U17179 ( .A(n12859), .B(n12860), .Z(n12855) );
  AND U17180 ( .A(n12861), .B(n12862), .Z(n12816) );
  NAND U17181 ( .A(n12863), .B(n12864), .Z(n12862) );
  NAND U17182 ( .A(n12865), .B(n12866), .Z(n12861) );
  AND U17183 ( .A(n12867), .B(n12868), .Z(n12818) );
  NAND U17184 ( .A(n12869), .B(n12870), .Z(n12812) );
  XNOR U17185 ( .A(n12795), .B(n12871), .Z(n12809) );
  XOR U17186 ( .A(n12799), .B(n12797), .Z(n12871) );
  XOR U17187 ( .A(n12805), .B(n12872), .Z(n12797) );
  XOR U17188 ( .A(n12802), .B(n12806), .Z(n12872) );
  NAND U17189 ( .A(n12873), .B(n12874), .Z(n12806) );
  NAND U17190 ( .A(n12875), .B(n12876), .Z(n12874) );
  NAND U17191 ( .A(n12877), .B(n12878), .Z(n12873) );
  AND U17192 ( .A(n12879), .B(n12880), .Z(n12802) );
  NAND U17193 ( .A(n12881), .B(n12882), .Z(n12880) );
  NAND U17194 ( .A(n12883), .B(n12884), .Z(n12879) );
  NANDN U17195 ( .A(n12885), .B(n12886), .Z(n12805) );
  NANDN U17196 ( .A(n12887), .B(n12888), .Z(n12799) );
  XNOR U17197 ( .A(n12790), .B(n12889), .Z(n12795) );
  XOR U17198 ( .A(n12788), .B(n12792), .Z(n12889) );
  NAND U17199 ( .A(n12890), .B(n12891), .Z(n12792) );
  NAND U17200 ( .A(n12892), .B(n12893), .Z(n12891) );
  NAND U17201 ( .A(n12894), .B(n12895), .Z(n12890) );
  AND U17202 ( .A(n12896), .B(n12897), .Z(n12788) );
  NAND U17203 ( .A(n12898), .B(n12899), .Z(n12897) );
  NAND U17204 ( .A(n12900), .B(n12901), .Z(n12896) );
  AND U17205 ( .A(n12902), .B(n12903), .Z(n12790) );
  XOR U17206 ( .A(n12870), .B(n12869), .Z(N29093) );
  XNOR U17207 ( .A(n12888), .B(n12887), .Z(n12869) );
  XNOR U17208 ( .A(n12902), .B(n12903), .Z(n12887) );
  XOR U17209 ( .A(n12899), .B(n12898), .Z(n12903) );
  XOR U17210 ( .A(y[2331]), .B(x[2331]), .Z(n12898) );
  XOR U17211 ( .A(n12901), .B(n12900), .Z(n12899) );
  XOR U17212 ( .A(y[2333]), .B(x[2333]), .Z(n12900) );
  XOR U17213 ( .A(y[2332]), .B(x[2332]), .Z(n12901) );
  XOR U17214 ( .A(n12893), .B(n12892), .Z(n12902) );
  XOR U17215 ( .A(n12895), .B(n12894), .Z(n12892) );
  XOR U17216 ( .A(y[2330]), .B(x[2330]), .Z(n12894) );
  XOR U17217 ( .A(y[2329]), .B(x[2329]), .Z(n12895) );
  XOR U17218 ( .A(y[2328]), .B(x[2328]), .Z(n12893) );
  XNOR U17219 ( .A(n12886), .B(n12885), .Z(n12888) );
  XNOR U17220 ( .A(n12882), .B(n12881), .Z(n12885) );
  XOR U17221 ( .A(n12884), .B(n12883), .Z(n12881) );
  XOR U17222 ( .A(y[2327]), .B(x[2327]), .Z(n12883) );
  XOR U17223 ( .A(y[2326]), .B(x[2326]), .Z(n12884) );
  XOR U17224 ( .A(y[2325]), .B(x[2325]), .Z(n12882) );
  XOR U17225 ( .A(n12876), .B(n12875), .Z(n12886) );
  XOR U17226 ( .A(n12878), .B(n12877), .Z(n12875) );
  XOR U17227 ( .A(y[2324]), .B(x[2324]), .Z(n12877) );
  XOR U17228 ( .A(y[2323]), .B(x[2323]), .Z(n12878) );
  XOR U17229 ( .A(y[2322]), .B(x[2322]), .Z(n12876) );
  XNOR U17230 ( .A(n12853), .B(n12852), .Z(n12870) );
  XNOR U17231 ( .A(n12867), .B(n12868), .Z(n12852) );
  XOR U17232 ( .A(n12864), .B(n12863), .Z(n12868) );
  XOR U17233 ( .A(y[2319]), .B(x[2319]), .Z(n12863) );
  XOR U17234 ( .A(n12866), .B(n12865), .Z(n12864) );
  XOR U17235 ( .A(y[2321]), .B(x[2321]), .Z(n12865) );
  XOR U17236 ( .A(y[2320]), .B(x[2320]), .Z(n12866) );
  XOR U17237 ( .A(n12858), .B(n12857), .Z(n12867) );
  XOR U17238 ( .A(n12860), .B(n12859), .Z(n12857) );
  XOR U17239 ( .A(y[2318]), .B(x[2318]), .Z(n12859) );
  XOR U17240 ( .A(y[2317]), .B(x[2317]), .Z(n12860) );
  XOR U17241 ( .A(y[2316]), .B(x[2316]), .Z(n12858) );
  XNOR U17242 ( .A(n12851), .B(n12850), .Z(n12853) );
  XNOR U17243 ( .A(n12847), .B(n12846), .Z(n12850) );
  XOR U17244 ( .A(n12849), .B(n12848), .Z(n12846) );
  XOR U17245 ( .A(y[2315]), .B(x[2315]), .Z(n12848) );
  XOR U17246 ( .A(y[2314]), .B(x[2314]), .Z(n12849) );
  XOR U17247 ( .A(y[2313]), .B(x[2313]), .Z(n12847) );
  XOR U17248 ( .A(n12841), .B(n12840), .Z(n12851) );
  XOR U17249 ( .A(n12843), .B(n12842), .Z(n12840) );
  XOR U17250 ( .A(y[2312]), .B(x[2312]), .Z(n12842) );
  XOR U17251 ( .A(y[2311]), .B(x[2311]), .Z(n12843) );
  XOR U17252 ( .A(y[2310]), .B(x[2310]), .Z(n12841) );
  NAND U17253 ( .A(n12904), .B(n12905), .Z(N29085) );
  NAND U17254 ( .A(n12906), .B(n12907), .Z(n12905) );
  NANDN U17255 ( .A(n12908), .B(n12909), .Z(n12907) );
  NANDN U17256 ( .A(n12909), .B(n12908), .Z(n12904) );
  XOR U17257 ( .A(n12908), .B(n12910), .Z(N29084) );
  XNOR U17258 ( .A(n12906), .B(n12909), .Z(n12910) );
  NAND U17259 ( .A(n12911), .B(n12912), .Z(n12909) );
  NAND U17260 ( .A(n12913), .B(n12914), .Z(n12912) );
  NANDN U17261 ( .A(n12915), .B(n12916), .Z(n12914) );
  NANDN U17262 ( .A(n12916), .B(n12915), .Z(n12911) );
  AND U17263 ( .A(n12917), .B(n12918), .Z(n12906) );
  NAND U17264 ( .A(n12919), .B(n12920), .Z(n12918) );
  OR U17265 ( .A(n12921), .B(n12922), .Z(n12920) );
  NAND U17266 ( .A(n12922), .B(n12921), .Z(n12917) );
  IV U17267 ( .A(n12923), .Z(n12922) );
  AND U17268 ( .A(n12924), .B(n12925), .Z(n12908) );
  NAND U17269 ( .A(n12926), .B(n12927), .Z(n12925) );
  NANDN U17270 ( .A(n12928), .B(n12929), .Z(n12927) );
  NANDN U17271 ( .A(n12929), .B(n12928), .Z(n12924) );
  XOR U17272 ( .A(n12921), .B(n12930), .Z(N29083) );
  XOR U17273 ( .A(n12919), .B(n12923), .Z(n12930) );
  XNOR U17274 ( .A(n12916), .B(n12931), .Z(n12923) );
  XNOR U17275 ( .A(n12913), .B(n12915), .Z(n12931) );
  AND U17276 ( .A(n12932), .B(n12933), .Z(n12915) );
  NANDN U17277 ( .A(n12934), .B(n12935), .Z(n12933) );
  NANDN U17278 ( .A(n12936), .B(n12937), .Z(n12935) );
  IV U17279 ( .A(n12938), .Z(n12937) );
  NAND U17280 ( .A(n12938), .B(n12936), .Z(n12932) );
  AND U17281 ( .A(n12939), .B(n12940), .Z(n12913) );
  NAND U17282 ( .A(n12941), .B(n12942), .Z(n12940) );
  OR U17283 ( .A(n12943), .B(n12944), .Z(n12942) );
  NAND U17284 ( .A(n12944), .B(n12943), .Z(n12939) );
  IV U17285 ( .A(n12945), .Z(n12944) );
  NAND U17286 ( .A(n12946), .B(n12947), .Z(n12916) );
  NANDN U17287 ( .A(n12948), .B(n12949), .Z(n12947) );
  NAND U17288 ( .A(n12950), .B(n12951), .Z(n12949) );
  OR U17289 ( .A(n12951), .B(n12950), .Z(n12946) );
  IV U17290 ( .A(n12952), .Z(n12950) );
  AND U17291 ( .A(n12953), .B(n12954), .Z(n12919) );
  NAND U17292 ( .A(n12955), .B(n12956), .Z(n12954) );
  NANDN U17293 ( .A(n12957), .B(n12958), .Z(n12956) );
  NANDN U17294 ( .A(n12958), .B(n12957), .Z(n12953) );
  XOR U17295 ( .A(n12929), .B(n12959), .Z(n12921) );
  XNOR U17296 ( .A(n12926), .B(n12928), .Z(n12959) );
  AND U17297 ( .A(n12960), .B(n12961), .Z(n12928) );
  NANDN U17298 ( .A(n12962), .B(n12963), .Z(n12961) );
  NANDN U17299 ( .A(n12964), .B(n12965), .Z(n12963) );
  IV U17300 ( .A(n12966), .Z(n12965) );
  NAND U17301 ( .A(n12966), .B(n12964), .Z(n12960) );
  AND U17302 ( .A(n12967), .B(n12968), .Z(n12926) );
  NAND U17303 ( .A(n12969), .B(n12970), .Z(n12968) );
  OR U17304 ( .A(n12971), .B(n12972), .Z(n12970) );
  NAND U17305 ( .A(n12972), .B(n12971), .Z(n12967) );
  IV U17306 ( .A(n12973), .Z(n12972) );
  NAND U17307 ( .A(n12974), .B(n12975), .Z(n12929) );
  NANDN U17308 ( .A(n12976), .B(n12977), .Z(n12975) );
  NAND U17309 ( .A(n12978), .B(n12979), .Z(n12977) );
  OR U17310 ( .A(n12979), .B(n12978), .Z(n12974) );
  IV U17311 ( .A(n12980), .Z(n12978) );
  XOR U17312 ( .A(n12955), .B(n12981), .Z(N29082) );
  XNOR U17313 ( .A(n12958), .B(n12957), .Z(n12981) );
  XNOR U17314 ( .A(n12969), .B(n12982), .Z(n12957) );
  XOR U17315 ( .A(n12973), .B(n12971), .Z(n12982) );
  XOR U17316 ( .A(n12979), .B(n12983), .Z(n12971) );
  XOR U17317 ( .A(n12976), .B(n12980), .Z(n12983) );
  NAND U17318 ( .A(n12984), .B(n12985), .Z(n12980) );
  NAND U17319 ( .A(n12986), .B(n12987), .Z(n12985) );
  NAND U17320 ( .A(n12988), .B(n12989), .Z(n12984) );
  AND U17321 ( .A(n12990), .B(n12991), .Z(n12976) );
  NAND U17322 ( .A(n12992), .B(n12993), .Z(n12991) );
  NAND U17323 ( .A(n12994), .B(n12995), .Z(n12990) );
  NANDN U17324 ( .A(n12996), .B(n12997), .Z(n12979) );
  NANDN U17325 ( .A(n12998), .B(n12999), .Z(n12973) );
  XNOR U17326 ( .A(n12964), .B(n13000), .Z(n12969) );
  XOR U17327 ( .A(n12962), .B(n12966), .Z(n13000) );
  NAND U17328 ( .A(n13001), .B(n13002), .Z(n12966) );
  NAND U17329 ( .A(n13003), .B(n13004), .Z(n13002) );
  NAND U17330 ( .A(n13005), .B(n13006), .Z(n13001) );
  AND U17331 ( .A(n13007), .B(n13008), .Z(n12962) );
  NAND U17332 ( .A(n13009), .B(n13010), .Z(n13008) );
  NAND U17333 ( .A(n13011), .B(n13012), .Z(n13007) );
  AND U17334 ( .A(n13013), .B(n13014), .Z(n12964) );
  NAND U17335 ( .A(n13015), .B(n13016), .Z(n12958) );
  XNOR U17336 ( .A(n12941), .B(n13017), .Z(n12955) );
  XOR U17337 ( .A(n12945), .B(n12943), .Z(n13017) );
  XOR U17338 ( .A(n12951), .B(n13018), .Z(n12943) );
  XOR U17339 ( .A(n12948), .B(n12952), .Z(n13018) );
  NAND U17340 ( .A(n13019), .B(n13020), .Z(n12952) );
  NAND U17341 ( .A(n13021), .B(n13022), .Z(n13020) );
  NAND U17342 ( .A(n13023), .B(n13024), .Z(n13019) );
  AND U17343 ( .A(n13025), .B(n13026), .Z(n12948) );
  NAND U17344 ( .A(n13027), .B(n13028), .Z(n13026) );
  NAND U17345 ( .A(n13029), .B(n13030), .Z(n13025) );
  NANDN U17346 ( .A(n13031), .B(n13032), .Z(n12951) );
  NANDN U17347 ( .A(n13033), .B(n13034), .Z(n12945) );
  XNOR U17348 ( .A(n12936), .B(n13035), .Z(n12941) );
  XOR U17349 ( .A(n12934), .B(n12938), .Z(n13035) );
  NAND U17350 ( .A(n13036), .B(n13037), .Z(n12938) );
  NAND U17351 ( .A(n13038), .B(n13039), .Z(n13037) );
  NAND U17352 ( .A(n13040), .B(n13041), .Z(n13036) );
  AND U17353 ( .A(n13042), .B(n13043), .Z(n12934) );
  NAND U17354 ( .A(n13044), .B(n13045), .Z(n13043) );
  NAND U17355 ( .A(n13046), .B(n13047), .Z(n13042) );
  AND U17356 ( .A(n13048), .B(n13049), .Z(n12936) );
  XOR U17357 ( .A(n13016), .B(n13015), .Z(N29081) );
  XNOR U17358 ( .A(n13034), .B(n13033), .Z(n13015) );
  XNOR U17359 ( .A(n13048), .B(n13049), .Z(n13033) );
  XOR U17360 ( .A(n13045), .B(n13044), .Z(n13049) );
  XOR U17361 ( .A(y[2307]), .B(x[2307]), .Z(n13044) );
  XOR U17362 ( .A(n13047), .B(n13046), .Z(n13045) );
  XOR U17363 ( .A(y[2309]), .B(x[2309]), .Z(n13046) );
  XOR U17364 ( .A(y[2308]), .B(x[2308]), .Z(n13047) );
  XOR U17365 ( .A(n13039), .B(n13038), .Z(n13048) );
  XOR U17366 ( .A(n13041), .B(n13040), .Z(n13038) );
  XOR U17367 ( .A(y[2306]), .B(x[2306]), .Z(n13040) );
  XOR U17368 ( .A(y[2305]), .B(x[2305]), .Z(n13041) );
  XOR U17369 ( .A(y[2304]), .B(x[2304]), .Z(n13039) );
  XNOR U17370 ( .A(n13032), .B(n13031), .Z(n13034) );
  XNOR U17371 ( .A(n13028), .B(n13027), .Z(n13031) );
  XOR U17372 ( .A(n13030), .B(n13029), .Z(n13027) );
  XOR U17373 ( .A(y[2303]), .B(x[2303]), .Z(n13029) );
  XOR U17374 ( .A(y[2302]), .B(x[2302]), .Z(n13030) );
  XOR U17375 ( .A(y[2301]), .B(x[2301]), .Z(n13028) );
  XOR U17376 ( .A(n13022), .B(n13021), .Z(n13032) );
  XOR U17377 ( .A(n13024), .B(n13023), .Z(n13021) );
  XOR U17378 ( .A(y[2300]), .B(x[2300]), .Z(n13023) );
  XOR U17379 ( .A(y[2299]), .B(x[2299]), .Z(n13024) );
  XOR U17380 ( .A(y[2298]), .B(x[2298]), .Z(n13022) );
  XNOR U17381 ( .A(n12999), .B(n12998), .Z(n13016) );
  XNOR U17382 ( .A(n13013), .B(n13014), .Z(n12998) );
  XOR U17383 ( .A(n13010), .B(n13009), .Z(n13014) );
  XOR U17384 ( .A(y[2295]), .B(x[2295]), .Z(n13009) );
  XOR U17385 ( .A(n13012), .B(n13011), .Z(n13010) );
  XOR U17386 ( .A(y[2297]), .B(x[2297]), .Z(n13011) );
  XOR U17387 ( .A(y[2296]), .B(x[2296]), .Z(n13012) );
  XOR U17388 ( .A(n13004), .B(n13003), .Z(n13013) );
  XOR U17389 ( .A(n13006), .B(n13005), .Z(n13003) );
  XOR U17390 ( .A(y[2294]), .B(x[2294]), .Z(n13005) );
  XOR U17391 ( .A(y[2293]), .B(x[2293]), .Z(n13006) );
  XOR U17392 ( .A(y[2292]), .B(x[2292]), .Z(n13004) );
  XNOR U17393 ( .A(n12997), .B(n12996), .Z(n12999) );
  XNOR U17394 ( .A(n12993), .B(n12992), .Z(n12996) );
  XOR U17395 ( .A(n12995), .B(n12994), .Z(n12992) );
  XOR U17396 ( .A(y[2291]), .B(x[2291]), .Z(n12994) );
  XOR U17397 ( .A(y[2290]), .B(x[2290]), .Z(n12995) );
  XOR U17398 ( .A(y[2289]), .B(x[2289]), .Z(n12993) );
  XOR U17399 ( .A(n12987), .B(n12986), .Z(n12997) );
  XOR U17400 ( .A(n12989), .B(n12988), .Z(n12986) );
  XOR U17401 ( .A(y[2288]), .B(x[2288]), .Z(n12988) );
  XOR U17402 ( .A(y[2287]), .B(x[2287]), .Z(n12989) );
  XOR U17403 ( .A(y[2286]), .B(x[2286]), .Z(n12987) );
  NAND U17404 ( .A(n13050), .B(n13051), .Z(N29073) );
  NAND U17405 ( .A(n13052), .B(n13053), .Z(n13051) );
  NANDN U17406 ( .A(n13054), .B(n13055), .Z(n13053) );
  NANDN U17407 ( .A(n13055), .B(n13054), .Z(n13050) );
  XOR U17408 ( .A(n13054), .B(n13056), .Z(N29072) );
  XNOR U17409 ( .A(n13052), .B(n13055), .Z(n13056) );
  NAND U17410 ( .A(n13057), .B(n13058), .Z(n13055) );
  NAND U17411 ( .A(n13059), .B(n13060), .Z(n13058) );
  NANDN U17412 ( .A(n13061), .B(n13062), .Z(n13060) );
  NANDN U17413 ( .A(n13062), .B(n13061), .Z(n13057) );
  AND U17414 ( .A(n13063), .B(n13064), .Z(n13052) );
  NAND U17415 ( .A(n13065), .B(n13066), .Z(n13064) );
  OR U17416 ( .A(n13067), .B(n13068), .Z(n13066) );
  NAND U17417 ( .A(n13068), .B(n13067), .Z(n13063) );
  IV U17418 ( .A(n13069), .Z(n13068) );
  AND U17419 ( .A(n13070), .B(n13071), .Z(n13054) );
  NAND U17420 ( .A(n13072), .B(n13073), .Z(n13071) );
  NANDN U17421 ( .A(n13074), .B(n13075), .Z(n13073) );
  NANDN U17422 ( .A(n13075), .B(n13074), .Z(n13070) );
  XOR U17423 ( .A(n13067), .B(n13076), .Z(N29071) );
  XOR U17424 ( .A(n13065), .B(n13069), .Z(n13076) );
  XNOR U17425 ( .A(n13062), .B(n13077), .Z(n13069) );
  XNOR U17426 ( .A(n13059), .B(n13061), .Z(n13077) );
  AND U17427 ( .A(n13078), .B(n13079), .Z(n13061) );
  NANDN U17428 ( .A(n13080), .B(n13081), .Z(n13079) );
  NANDN U17429 ( .A(n13082), .B(n13083), .Z(n13081) );
  IV U17430 ( .A(n13084), .Z(n13083) );
  NAND U17431 ( .A(n13084), .B(n13082), .Z(n13078) );
  AND U17432 ( .A(n13085), .B(n13086), .Z(n13059) );
  NAND U17433 ( .A(n13087), .B(n13088), .Z(n13086) );
  OR U17434 ( .A(n13089), .B(n13090), .Z(n13088) );
  NAND U17435 ( .A(n13090), .B(n13089), .Z(n13085) );
  IV U17436 ( .A(n13091), .Z(n13090) );
  NAND U17437 ( .A(n13092), .B(n13093), .Z(n13062) );
  NANDN U17438 ( .A(n13094), .B(n13095), .Z(n13093) );
  NAND U17439 ( .A(n13096), .B(n13097), .Z(n13095) );
  OR U17440 ( .A(n13097), .B(n13096), .Z(n13092) );
  IV U17441 ( .A(n13098), .Z(n13096) );
  AND U17442 ( .A(n13099), .B(n13100), .Z(n13065) );
  NAND U17443 ( .A(n13101), .B(n13102), .Z(n13100) );
  NANDN U17444 ( .A(n13103), .B(n13104), .Z(n13102) );
  NANDN U17445 ( .A(n13104), .B(n13103), .Z(n13099) );
  XOR U17446 ( .A(n13075), .B(n13105), .Z(n13067) );
  XNOR U17447 ( .A(n13072), .B(n13074), .Z(n13105) );
  AND U17448 ( .A(n13106), .B(n13107), .Z(n13074) );
  NANDN U17449 ( .A(n13108), .B(n13109), .Z(n13107) );
  NANDN U17450 ( .A(n13110), .B(n13111), .Z(n13109) );
  IV U17451 ( .A(n13112), .Z(n13111) );
  NAND U17452 ( .A(n13112), .B(n13110), .Z(n13106) );
  AND U17453 ( .A(n13113), .B(n13114), .Z(n13072) );
  NAND U17454 ( .A(n13115), .B(n13116), .Z(n13114) );
  OR U17455 ( .A(n13117), .B(n13118), .Z(n13116) );
  NAND U17456 ( .A(n13118), .B(n13117), .Z(n13113) );
  IV U17457 ( .A(n13119), .Z(n13118) );
  NAND U17458 ( .A(n13120), .B(n13121), .Z(n13075) );
  NANDN U17459 ( .A(n13122), .B(n13123), .Z(n13121) );
  NAND U17460 ( .A(n13124), .B(n13125), .Z(n13123) );
  OR U17461 ( .A(n13125), .B(n13124), .Z(n13120) );
  IV U17462 ( .A(n13126), .Z(n13124) );
  XOR U17463 ( .A(n13101), .B(n13127), .Z(N29070) );
  XNOR U17464 ( .A(n13104), .B(n13103), .Z(n13127) );
  XNOR U17465 ( .A(n13115), .B(n13128), .Z(n13103) );
  XOR U17466 ( .A(n13119), .B(n13117), .Z(n13128) );
  XOR U17467 ( .A(n13125), .B(n13129), .Z(n13117) );
  XOR U17468 ( .A(n13122), .B(n13126), .Z(n13129) );
  NAND U17469 ( .A(n13130), .B(n13131), .Z(n13126) );
  NAND U17470 ( .A(n13132), .B(n13133), .Z(n13131) );
  NAND U17471 ( .A(n13134), .B(n13135), .Z(n13130) );
  AND U17472 ( .A(n13136), .B(n13137), .Z(n13122) );
  NAND U17473 ( .A(n13138), .B(n13139), .Z(n13137) );
  NAND U17474 ( .A(n13140), .B(n13141), .Z(n13136) );
  NANDN U17475 ( .A(n13142), .B(n13143), .Z(n13125) );
  NANDN U17476 ( .A(n13144), .B(n13145), .Z(n13119) );
  XNOR U17477 ( .A(n13110), .B(n13146), .Z(n13115) );
  XOR U17478 ( .A(n13108), .B(n13112), .Z(n13146) );
  NAND U17479 ( .A(n13147), .B(n13148), .Z(n13112) );
  NAND U17480 ( .A(n13149), .B(n13150), .Z(n13148) );
  NAND U17481 ( .A(n13151), .B(n13152), .Z(n13147) );
  AND U17482 ( .A(n13153), .B(n13154), .Z(n13108) );
  NAND U17483 ( .A(n13155), .B(n13156), .Z(n13154) );
  NAND U17484 ( .A(n13157), .B(n13158), .Z(n13153) );
  AND U17485 ( .A(n13159), .B(n13160), .Z(n13110) );
  NAND U17486 ( .A(n13161), .B(n13162), .Z(n13104) );
  XNOR U17487 ( .A(n13087), .B(n13163), .Z(n13101) );
  XOR U17488 ( .A(n13091), .B(n13089), .Z(n13163) );
  XOR U17489 ( .A(n13097), .B(n13164), .Z(n13089) );
  XOR U17490 ( .A(n13094), .B(n13098), .Z(n13164) );
  NAND U17491 ( .A(n13165), .B(n13166), .Z(n13098) );
  NAND U17492 ( .A(n13167), .B(n13168), .Z(n13166) );
  NAND U17493 ( .A(n13169), .B(n13170), .Z(n13165) );
  AND U17494 ( .A(n13171), .B(n13172), .Z(n13094) );
  NAND U17495 ( .A(n13173), .B(n13174), .Z(n13172) );
  NAND U17496 ( .A(n13175), .B(n13176), .Z(n13171) );
  NANDN U17497 ( .A(n13177), .B(n13178), .Z(n13097) );
  NANDN U17498 ( .A(n13179), .B(n13180), .Z(n13091) );
  XNOR U17499 ( .A(n13082), .B(n13181), .Z(n13087) );
  XOR U17500 ( .A(n13080), .B(n13084), .Z(n13181) );
  NAND U17501 ( .A(n13182), .B(n13183), .Z(n13084) );
  NAND U17502 ( .A(n13184), .B(n13185), .Z(n13183) );
  NAND U17503 ( .A(n13186), .B(n13187), .Z(n13182) );
  AND U17504 ( .A(n13188), .B(n13189), .Z(n13080) );
  NAND U17505 ( .A(n13190), .B(n13191), .Z(n13189) );
  NAND U17506 ( .A(n13192), .B(n13193), .Z(n13188) );
  AND U17507 ( .A(n13194), .B(n13195), .Z(n13082) );
  XOR U17508 ( .A(n13162), .B(n13161), .Z(N29069) );
  XNOR U17509 ( .A(n13180), .B(n13179), .Z(n13161) );
  XNOR U17510 ( .A(n13194), .B(n13195), .Z(n13179) );
  XOR U17511 ( .A(n13191), .B(n13190), .Z(n13195) );
  XOR U17512 ( .A(y[2283]), .B(x[2283]), .Z(n13190) );
  XOR U17513 ( .A(n13193), .B(n13192), .Z(n13191) );
  XOR U17514 ( .A(y[2285]), .B(x[2285]), .Z(n13192) );
  XOR U17515 ( .A(y[2284]), .B(x[2284]), .Z(n13193) );
  XOR U17516 ( .A(n13185), .B(n13184), .Z(n13194) );
  XOR U17517 ( .A(n13187), .B(n13186), .Z(n13184) );
  XOR U17518 ( .A(y[2282]), .B(x[2282]), .Z(n13186) );
  XOR U17519 ( .A(y[2281]), .B(x[2281]), .Z(n13187) );
  XOR U17520 ( .A(y[2280]), .B(x[2280]), .Z(n13185) );
  XNOR U17521 ( .A(n13178), .B(n13177), .Z(n13180) );
  XNOR U17522 ( .A(n13174), .B(n13173), .Z(n13177) );
  XOR U17523 ( .A(n13176), .B(n13175), .Z(n13173) );
  XOR U17524 ( .A(y[2279]), .B(x[2279]), .Z(n13175) );
  XOR U17525 ( .A(y[2278]), .B(x[2278]), .Z(n13176) );
  XOR U17526 ( .A(y[2277]), .B(x[2277]), .Z(n13174) );
  XOR U17527 ( .A(n13168), .B(n13167), .Z(n13178) );
  XOR U17528 ( .A(n13170), .B(n13169), .Z(n13167) );
  XOR U17529 ( .A(y[2276]), .B(x[2276]), .Z(n13169) );
  XOR U17530 ( .A(y[2275]), .B(x[2275]), .Z(n13170) );
  XOR U17531 ( .A(y[2274]), .B(x[2274]), .Z(n13168) );
  XNOR U17532 ( .A(n13145), .B(n13144), .Z(n13162) );
  XNOR U17533 ( .A(n13159), .B(n13160), .Z(n13144) );
  XOR U17534 ( .A(n13156), .B(n13155), .Z(n13160) );
  XOR U17535 ( .A(y[2271]), .B(x[2271]), .Z(n13155) );
  XOR U17536 ( .A(n13158), .B(n13157), .Z(n13156) );
  XOR U17537 ( .A(y[2273]), .B(x[2273]), .Z(n13157) );
  XOR U17538 ( .A(y[2272]), .B(x[2272]), .Z(n13158) );
  XOR U17539 ( .A(n13150), .B(n13149), .Z(n13159) );
  XOR U17540 ( .A(n13152), .B(n13151), .Z(n13149) );
  XOR U17541 ( .A(y[2270]), .B(x[2270]), .Z(n13151) );
  XOR U17542 ( .A(y[2269]), .B(x[2269]), .Z(n13152) );
  XOR U17543 ( .A(y[2268]), .B(x[2268]), .Z(n13150) );
  XNOR U17544 ( .A(n13143), .B(n13142), .Z(n13145) );
  XNOR U17545 ( .A(n13139), .B(n13138), .Z(n13142) );
  XOR U17546 ( .A(n13141), .B(n13140), .Z(n13138) );
  XOR U17547 ( .A(y[2267]), .B(x[2267]), .Z(n13140) );
  XOR U17548 ( .A(y[2266]), .B(x[2266]), .Z(n13141) );
  XOR U17549 ( .A(y[2265]), .B(x[2265]), .Z(n13139) );
  XOR U17550 ( .A(n13133), .B(n13132), .Z(n13143) );
  XOR U17551 ( .A(n13135), .B(n13134), .Z(n13132) );
  XOR U17552 ( .A(y[2264]), .B(x[2264]), .Z(n13134) );
  XOR U17553 ( .A(y[2263]), .B(x[2263]), .Z(n13135) );
  XOR U17554 ( .A(y[2262]), .B(x[2262]), .Z(n13133) );
  NAND U17555 ( .A(n13196), .B(n13197), .Z(N29061) );
  NAND U17556 ( .A(n13198), .B(n13199), .Z(n13197) );
  NANDN U17557 ( .A(n13200), .B(n13201), .Z(n13199) );
  NANDN U17558 ( .A(n13201), .B(n13200), .Z(n13196) );
  XOR U17559 ( .A(n13200), .B(n13202), .Z(N29060) );
  XNOR U17560 ( .A(n13198), .B(n13201), .Z(n13202) );
  NAND U17561 ( .A(n13203), .B(n13204), .Z(n13201) );
  NAND U17562 ( .A(n13205), .B(n13206), .Z(n13204) );
  NANDN U17563 ( .A(n13207), .B(n13208), .Z(n13206) );
  NANDN U17564 ( .A(n13208), .B(n13207), .Z(n13203) );
  AND U17565 ( .A(n13209), .B(n13210), .Z(n13198) );
  NAND U17566 ( .A(n13211), .B(n13212), .Z(n13210) );
  OR U17567 ( .A(n13213), .B(n13214), .Z(n13212) );
  NAND U17568 ( .A(n13214), .B(n13213), .Z(n13209) );
  IV U17569 ( .A(n13215), .Z(n13214) );
  AND U17570 ( .A(n13216), .B(n13217), .Z(n13200) );
  NAND U17571 ( .A(n13218), .B(n13219), .Z(n13217) );
  NANDN U17572 ( .A(n13220), .B(n13221), .Z(n13219) );
  NANDN U17573 ( .A(n13221), .B(n13220), .Z(n13216) );
  XOR U17574 ( .A(n13213), .B(n13222), .Z(N29059) );
  XOR U17575 ( .A(n13211), .B(n13215), .Z(n13222) );
  XNOR U17576 ( .A(n13208), .B(n13223), .Z(n13215) );
  XNOR U17577 ( .A(n13205), .B(n13207), .Z(n13223) );
  AND U17578 ( .A(n13224), .B(n13225), .Z(n13207) );
  NANDN U17579 ( .A(n13226), .B(n13227), .Z(n13225) );
  NANDN U17580 ( .A(n13228), .B(n13229), .Z(n13227) );
  IV U17581 ( .A(n13230), .Z(n13229) );
  NAND U17582 ( .A(n13230), .B(n13228), .Z(n13224) );
  AND U17583 ( .A(n13231), .B(n13232), .Z(n13205) );
  NAND U17584 ( .A(n13233), .B(n13234), .Z(n13232) );
  OR U17585 ( .A(n13235), .B(n13236), .Z(n13234) );
  NAND U17586 ( .A(n13236), .B(n13235), .Z(n13231) );
  IV U17587 ( .A(n13237), .Z(n13236) );
  NAND U17588 ( .A(n13238), .B(n13239), .Z(n13208) );
  NANDN U17589 ( .A(n13240), .B(n13241), .Z(n13239) );
  NAND U17590 ( .A(n13242), .B(n13243), .Z(n13241) );
  OR U17591 ( .A(n13243), .B(n13242), .Z(n13238) );
  IV U17592 ( .A(n13244), .Z(n13242) );
  AND U17593 ( .A(n13245), .B(n13246), .Z(n13211) );
  NAND U17594 ( .A(n13247), .B(n13248), .Z(n13246) );
  NANDN U17595 ( .A(n13249), .B(n13250), .Z(n13248) );
  NANDN U17596 ( .A(n13250), .B(n13249), .Z(n13245) );
  XOR U17597 ( .A(n13221), .B(n13251), .Z(n13213) );
  XNOR U17598 ( .A(n13218), .B(n13220), .Z(n13251) );
  AND U17599 ( .A(n13252), .B(n13253), .Z(n13220) );
  NANDN U17600 ( .A(n13254), .B(n13255), .Z(n13253) );
  NANDN U17601 ( .A(n13256), .B(n13257), .Z(n13255) );
  IV U17602 ( .A(n13258), .Z(n13257) );
  NAND U17603 ( .A(n13258), .B(n13256), .Z(n13252) );
  AND U17604 ( .A(n13259), .B(n13260), .Z(n13218) );
  NAND U17605 ( .A(n13261), .B(n13262), .Z(n13260) );
  OR U17606 ( .A(n13263), .B(n13264), .Z(n13262) );
  NAND U17607 ( .A(n13264), .B(n13263), .Z(n13259) );
  IV U17608 ( .A(n13265), .Z(n13264) );
  NAND U17609 ( .A(n13266), .B(n13267), .Z(n13221) );
  NANDN U17610 ( .A(n13268), .B(n13269), .Z(n13267) );
  NAND U17611 ( .A(n13270), .B(n13271), .Z(n13269) );
  OR U17612 ( .A(n13271), .B(n13270), .Z(n13266) );
  IV U17613 ( .A(n13272), .Z(n13270) );
  XOR U17614 ( .A(n13247), .B(n13273), .Z(N29058) );
  XNOR U17615 ( .A(n13250), .B(n13249), .Z(n13273) );
  XNOR U17616 ( .A(n13261), .B(n13274), .Z(n13249) );
  XOR U17617 ( .A(n13265), .B(n13263), .Z(n13274) );
  XOR U17618 ( .A(n13271), .B(n13275), .Z(n13263) );
  XOR U17619 ( .A(n13268), .B(n13272), .Z(n13275) );
  NAND U17620 ( .A(n13276), .B(n13277), .Z(n13272) );
  NAND U17621 ( .A(n13278), .B(n13279), .Z(n13277) );
  NAND U17622 ( .A(n13280), .B(n13281), .Z(n13276) );
  AND U17623 ( .A(n13282), .B(n13283), .Z(n13268) );
  NAND U17624 ( .A(n13284), .B(n13285), .Z(n13283) );
  NAND U17625 ( .A(n13286), .B(n13287), .Z(n13282) );
  NANDN U17626 ( .A(n13288), .B(n13289), .Z(n13271) );
  NANDN U17627 ( .A(n13290), .B(n13291), .Z(n13265) );
  XNOR U17628 ( .A(n13256), .B(n13292), .Z(n13261) );
  XOR U17629 ( .A(n13254), .B(n13258), .Z(n13292) );
  NAND U17630 ( .A(n13293), .B(n13294), .Z(n13258) );
  NAND U17631 ( .A(n13295), .B(n13296), .Z(n13294) );
  NAND U17632 ( .A(n13297), .B(n13298), .Z(n13293) );
  AND U17633 ( .A(n13299), .B(n13300), .Z(n13254) );
  NAND U17634 ( .A(n13301), .B(n13302), .Z(n13300) );
  NAND U17635 ( .A(n13303), .B(n13304), .Z(n13299) );
  AND U17636 ( .A(n13305), .B(n13306), .Z(n13256) );
  NAND U17637 ( .A(n13307), .B(n13308), .Z(n13250) );
  XNOR U17638 ( .A(n13233), .B(n13309), .Z(n13247) );
  XOR U17639 ( .A(n13237), .B(n13235), .Z(n13309) );
  XOR U17640 ( .A(n13243), .B(n13310), .Z(n13235) );
  XOR U17641 ( .A(n13240), .B(n13244), .Z(n13310) );
  NAND U17642 ( .A(n13311), .B(n13312), .Z(n13244) );
  NAND U17643 ( .A(n13313), .B(n13314), .Z(n13312) );
  NAND U17644 ( .A(n13315), .B(n13316), .Z(n13311) );
  AND U17645 ( .A(n13317), .B(n13318), .Z(n13240) );
  NAND U17646 ( .A(n13319), .B(n13320), .Z(n13318) );
  NAND U17647 ( .A(n13321), .B(n13322), .Z(n13317) );
  NANDN U17648 ( .A(n13323), .B(n13324), .Z(n13243) );
  NANDN U17649 ( .A(n13325), .B(n13326), .Z(n13237) );
  XNOR U17650 ( .A(n13228), .B(n13327), .Z(n13233) );
  XOR U17651 ( .A(n13226), .B(n13230), .Z(n13327) );
  NAND U17652 ( .A(n13328), .B(n13329), .Z(n13230) );
  NAND U17653 ( .A(n13330), .B(n13331), .Z(n13329) );
  NAND U17654 ( .A(n13332), .B(n13333), .Z(n13328) );
  AND U17655 ( .A(n13334), .B(n13335), .Z(n13226) );
  NAND U17656 ( .A(n13336), .B(n13337), .Z(n13335) );
  NAND U17657 ( .A(n13338), .B(n13339), .Z(n13334) );
  AND U17658 ( .A(n13340), .B(n13341), .Z(n13228) );
  XOR U17659 ( .A(n13308), .B(n13307), .Z(N29057) );
  XNOR U17660 ( .A(n13326), .B(n13325), .Z(n13307) );
  XNOR U17661 ( .A(n13340), .B(n13341), .Z(n13325) );
  XOR U17662 ( .A(n13337), .B(n13336), .Z(n13341) );
  XOR U17663 ( .A(y[2259]), .B(x[2259]), .Z(n13336) );
  XOR U17664 ( .A(n13339), .B(n13338), .Z(n13337) );
  XOR U17665 ( .A(y[2261]), .B(x[2261]), .Z(n13338) );
  XOR U17666 ( .A(y[2260]), .B(x[2260]), .Z(n13339) );
  XOR U17667 ( .A(n13331), .B(n13330), .Z(n13340) );
  XOR U17668 ( .A(n13333), .B(n13332), .Z(n13330) );
  XOR U17669 ( .A(y[2258]), .B(x[2258]), .Z(n13332) );
  XOR U17670 ( .A(y[2257]), .B(x[2257]), .Z(n13333) );
  XOR U17671 ( .A(y[2256]), .B(x[2256]), .Z(n13331) );
  XNOR U17672 ( .A(n13324), .B(n13323), .Z(n13326) );
  XNOR U17673 ( .A(n13320), .B(n13319), .Z(n13323) );
  XOR U17674 ( .A(n13322), .B(n13321), .Z(n13319) );
  XOR U17675 ( .A(y[2255]), .B(x[2255]), .Z(n13321) );
  XOR U17676 ( .A(y[2254]), .B(x[2254]), .Z(n13322) );
  XOR U17677 ( .A(y[2253]), .B(x[2253]), .Z(n13320) );
  XOR U17678 ( .A(n13314), .B(n13313), .Z(n13324) );
  XOR U17679 ( .A(n13316), .B(n13315), .Z(n13313) );
  XOR U17680 ( .A(y[2252]), .B(x[2252]), .Z(n13315) );
  XOR U17681 ( .A(y[2251]), .B(x[2251]), .Z(n13316) );
  XOR U17682 ( .A(y[2250]), .B(x[2250]), .Z(n13314) );
  XNOR U17683 ( .A(n13291), .B(n13290), .Z(n13308) );
  XNOR U17684 ( .A(n13305), .B(n13306), .Z(n13290) );
  XOR U17685 ( .A(n13302), .B(n13301), .Z(n13306) );
  XOR U17686 ( .A(y[2247]), .B(x[2247]), .Z(n13301) );
  XOR U17687 ( .A(n13304), .B(n13303), .Z(n13302) );
  XOR U17688 ( .A(y[2249]), .B(x[2249]), .Z(n13303) );
  XOR U17689 ( .A(y[2248]), .B(x[2248]), .Z(n13304) );
  XOR U17690 ( .A(n13296), .B(n13295), .Z(n13305) );
  XOR U17691 ( .A(n13298), .B(n13297), .Z(n13295) );
  XOR U17692 ( .A(y[2246]), .B(x[2246]), .Z(n13297) );
  XOR U17693 ( .A(y[2245]), .B(x[2245]), .Z(n13298) );
  XOR U17694 ( .A(y[2244]), .B(x[2244]), .Z(n13296) );
  XNOR U17695 ( .A(n13289), .B(n13288), .Z(n13291) );
  XNOR U17696 ( .A(n13285), .B(n13284), .Z(n13288) );
  XOR U17697 ( .A(n13287), .B(n13286), .Z(n13284) );
  XOR U17698 ( .A(y[2243]), .B(x[2243]), .Z(n13286) );
  XOR U17699 ( .A(y[2242]), .B(x[2242]), .Z(n13287) );
  XOR U17700 ( .A(y[2241]), .B(x[2241]), .Z(n13285) );
  XOR U17701 ( .A(n13279), .B(n13278), .Z(n13289) );
  XOR U17702 ( .A(n13281), .B(n13280), .Z(n13278) );
  XOR U17703 ( .A(y[2240]), .B(x[2240]), .Z(n13280) );
  XOR U17704 ( .A(y[2239]), .B(x[2239]), .Z(n13281) );
  XOR U17705 ( .A(y[2238]), .B(x[2238]), .Z(n13279) );
  NAND U17706 ( .A(n13342), .B(n13343), .Z(N29049) );
  NAND U17707 ( .A(n13344), .B(n13345), .Z(n13343) );
  NANDN U17708 ( .A(n13346), .B(n13347), .Z(n13345) );
  NANDN U17709 ( .A(n13347), .B(n13346), .Z(n13342) );
  XOR U17710 ( .A(n13346), .B(n13348), .Z(N29048) );
  XNOR U17711 ( .A(n13344), .B(n13347), .Z(n13348) );
  NAND U17712 ( .A(n13349), .B(n13350), .Z(n13347) );
  NAND U17713 ( .A(n13351), .B(n13352), .Z(n13350) );
  NANDN U17714 ( .A(n13353), .B(n13354), .Z(n13352) );
  NANDN U17715 ( .A(n13354), .B(n13353), .Z(n13349) );
  AND U17716 ( .A(n13355), .B(n13356), .Z(n13344) );
  NAND U17717 ( .A(n13357), .B(n13358), .Z(n13356) );
  OR U17718 ( .A(n13359), .B(n13360), .Z(n13358) );
  NAND U17719 ( .A(n13360), .B(n13359), .Z(n13355) );
  IV U17720 ( .A(n13361), .Z(n13360) );
  AND U17721 ( .A(n13362), .B(n13363), .Z(n13346) );
  NAND U17722 ( .A(n13364), .B(n13365), .Z(n13363) );
  NANDN U17723 ( .A(n13366), .B(n13367), .Z(n13365) );
  NANDN U17724 ( .A(n13367), .B(n13366), .Z(n13362) );
  XOR U17725 ( .A(n13359), .B(n13368), .Z(N29047) );
  XOR U17726 ( .A(n13357), .B(n13361), .Z(n13368) );
  XNOR U17727 ( .A(n13354), .B(n13369), .Z(n13361) );
  XNOR U17728 ( .A(n13351), .B(n13353), .Z(n13369) );
  AND U17729 ( .A(n13370), .B(n13371), .Z(n13353) );
  NANDN U17730 ( .A(n13372), .B(n13373), .Z(n13371) );
  NANDN U17731 ( .A(n13374), .B(n13375), .Z(n13373) );
  IV U17732 ( .A(n13376), .Z(n13375) );
  NAND U17733 ( .A(n13376), .B(n13374), .Z(n13370) );
  AND U17734 ( .A(n13377), .B(n13378), .Z(n13351) );
  NAND U17735 ( .A(n13379), .B(n13380), .Z(n13378) );
  OR U17736 ( .A(n13381), .B(n13382), .Z(n13380) );
  NAND U17737 ( .A(n13382), .B(n13381), .Z(n13377) );
  IV U17738 ( .A(n13383), .Z(n13382) );
  NAND U17739 ( .A(n13384), .B(n13385), .Z(n13354) );
  NANDN U17740 ( .A(n13386), .B(n13387), .Z(n13385) );
  NAND U17741 ( .A(n13388), .B(n13389), .Z(n13387) );
  OR U17742 ( .A(n13389), .B(n13388), .Z(n13384) );
  IV U17743 ( .A(n13390), .Z(n13388) );
  AND U17744 ( .A(n13391), .B(n13392), .Z(n13357) );
  NAND U17745 ( .A(n13393), .B(n13394), .Z(n13392) );
  NANDN U17746 ( .A(n13395), .B(n13396), .Z(n13394) );
  NANDN U17747 ( .A(n13396), .B(n13395), .Z(n13391) );
  XOR U17748 ( .A(n13367), .B(n13397), .Z(n13359) );
  XNOR U17749 ( .A(n13364), .B(n13366), .Z(n13397) );
  AND U17750 ( .A(n13398), .B(n13399), .Z(n13366) );
  NANDN U17751 ( .A(n13400), .B(n13401), .Z(n13399) );
  NANDN U17752 ( .A(n13402), .B(n13403), .Z(n13401) );
  IV U17753 ( .A(n13404), .Z(n13403) );
  NAND U17754 ( .A(n13404), .B(n13402), .Z(n13398) );
  AND U17755 ( .A(n13405), .B(n13406), .Z(n13364) );
  NAND U17756 ( .A(n13407), .B(n13408), .Z(n13406) );
  OR U17757 ( .A(n13409), .B(n13410), .Z(n13408) );
  NAND U17758 ( .A(n13410), .B(n13409), .Z(n13405) );
  IV U17759 ( .A(n13411), .Z(n13410) );
  NAND U17760 ( .A(n13412), .B(n13413), .Z(n13367) );
  NANDN U17761 ( .A(n13414), .B(n13415), .Z(n13413) );
  NAND U17762 ( .A(n13416), .B(n13417), .Z(n13415) );
  OR U17763 ( .A(n13417), .B(n13416), .Z(n13412) );
  IV U17764 ( .A(n13418), .Z(n13416) );
  XOR U17765 ( .A(n13393), .B(n13419), .Z(N29046) );
  XNOR U17766 ( .A(n13396), .B(n13395), .Z(n13419) );
  XNOR U17767 ( .A(n13407), .B(n13420), .Z(n13395) );
  XOR U17768 ( .A(n13411), .B(n13409), .Z(n13420) );
  XOR U17769 ( .A(n13417), .B(n13421), .Z(n13409) );
  XOR U17770 ( .A(n13414), .B(n13418), .Z(n13421) );
  NAND U17771 ( .A(n13422), .B(n13423), .Z(n13418) );
  NAND U17772 ( .A(n13424), .B(n13425), .Z(n13423) );
  NAND U17773 ( .A(n13426), .B(n13427), .Z(n13422) );
  AND U17774 ( .A(n13428), .B(n13429), .Z(n13414) );
  NAND U17775 ( .A(n13430), .B(n13431), .Z(n13429) );
  NAND U17776 ( .A(n13432), .B(n13433), .Z(n13428) );
  NANDN U17777 ( .A(n13434), .B(n13435), .Z(n13417) );
  NANDN U17778 ( .A(n13436), .B(n13437), .Z(n13411) );
  XNOR U17779 ( .A(n13402), .B(n13438), .Z(n13407) );
  XOR U17780 ( .A(n13400), .B(n13404), .Z(n13438) );
  NAND U17781 ( .A(n13439), .B(n13440), .Z(n13404) );
  NAND U17782 ( .A(n13441), .B(n13442), .Z(n13440) );
  NAND U17783 ( .A(n13443), .B(n13444), .Z(n13439) );
  AND U17784 ( .A(n13445), .B(n13446), .Z(n13400) );
  NAND U17785 ( .A(n13447), .B(n13448), .Z(n13446) );
  NAND U17786 ( .A(n13449), .B(n13450), .Z(n13445) );
  AND U17787 ( .A(n13451), .B(n13452), .Z(n13402) );
  NAND U17788 ( .A(n13453), .B(n13454), .Z(n13396) );
  XNOR U17789 ( .A(n13379), .B(n13455), .Z(n13393) );
  XOR U17790 ( .A(n13383), .B(n13381), .Z(n13455) );
  XOR U17791 ( .A(n13389), .B(n13456), .Z(n13381) );
  XOR U17792 ( .A(n13386), .B(n13390), .Z(n13456) );
  NAND U17793 ( .A(n13457), .B(n13458), .Z(n13390) );
  NAND U17794 ( .A(n13459), .B(n13460), .Z(n13458) );
  NAND U17795 ( .A(n13461), .B(n13462), .Z(n13457) );
  AND U17796 ( .A(n13463), .B(n13464), .Z(n13386) );
  NAND U17797 ( .A(n13465), .B(n13466), .Z(n13464) );
  NAND U17798 ( .A(n13467), .B(n13468), .Z(n13463) );
  NANDN U17799 ( .A(n13469), .B(n13470), .Z(n13389) );
  NANDN U17800 ( .A(n13471), .B(n13472), .Z(n13383) );
  XNOR U17801 ( .A(n13374), .B(n13473), .Z(n13379) );
  XOR U17802 ( .A(n13372), .B(n13376), .Z(n13473) );
  NAND U17803 ( .A(n13474), .B(n13475), .Z(n13376) );
  NAND U17804 ( .A(n13476), .B(n13477), .Z(n13475) );
  NAND U17805 ( .A(n13478), .B(n13479), .Z(n13474) );
  AND U17806 ( .A(n13480), .B(n13481), .Z(n13372) );
  NAND U17807 ( .A(n13482), .B(n13483), .Z(n13481) );
  NAND U17808 ( .A(n13484), .B(n13485), .Z(n13480) );
  AND U17809 ( .A(n13486), .B(n13487), .Z(n13374) );
  XOR U17810 ( .A(n13454), .B(n13453), .Z(N29045) );
  XNOR U17811 ( .A(n13472), .B(n13471), .Z(n13453) );
  XNOR U17812 ( .A(n13486), .B(n13487), .Z(n13471) );
  XOR U17813 ( .A(n13483), .B(n13482), .Z(n13487) );
  XOR U17814 ( .A(y[2235]), .B(x[2235]), .Z(n13482) );
  XOR U17815 ( .A(n13485), .B(n13484), .Z(n13483) );
  XOR U17816 ( .A(y[2237]), .B(x[2237]), .Z(n13484) );
  XOR U17817 ( .A(y[2236]), .B(x[2236]), .Z(n13485) );
  XOR U17818 ( .A(n13477), .B(n13476), .Z(n13486) );
  XOR U17819 ( .A(n13479), .B(n13478), .Z(n13476) );
  XOR U17820 ( .A(y[2234]), .B(x[2234]), .Z(n13478) );
  XOR U17821 ( .A(y[2233]), .B(x[2233]), .Z(n13479) );
  XOR U17822 ( .A(y[2232]), .B(x[2232]), .Z(n13477) );
  XNOR U17823 ( .A(n13470), .B(n13469), .Z(n13472) );
  XNOR U17824 ( .A(n13466), .B(n13465), .Z(n13469) );
  XOR U17825 ( .A(n13468), .B(n13467), .Z(n13465) );
  XOR U17826 ( .A(y[2231]), .B(x[2231]), .Z(n13467) );
  XOR U17827 ( .A(y[2230]), .B(x[2230]), .Z(n13468) );
  XOR U17828 ( .A(y[2229]), .B(x[2229]), .Z(n13466) );
  XOR U17829 ( .A(n13460), .B(n13459), .Z(n13470) );
  XOR U17830 ( .A(n13462), .B(n13461), .Z(n13459) );
  XOR U17831 ( .A(y[2228]), .B(x[2228]), .Z(n13461) );
  XOR U17832 ( .A(y[2227]), .B(x[2227]), .Z(n13462) );
  XOR U17833 ( .A(y[2226]), .B(x[2226]), .Z(n13460) );
  XNOR U17834 ( .A(n13437), .B(n13436), .Z(n13454) );
  XNOR U17835 ( .A(n13451), .B(n13452), .Z(n13436) );
  XOR U17836 ( .A(n13448), .B(n13447), .Z(n13452) );
  XOR U17837 ( .A(y[2223]), .B(x[2223]), .Z(n13447) );
  XOR U17838 ( .A(n13450), .B(n13449), .Z(n13448) );
  XOR U17839 ( .A(y[2225]), .B(x[2225]), .Z(n13449) );
  XOR U17840 ( .A(y[2224]), .B(x[2224]), .Z(n13450) );
  XOR U17841 ( .A(n13442), .B(n13441), .Z(n13451) );
  XOR U17842 ( .A(n13444), .B(n13443), .Z(n13441) );
  XOR U17843 ( .A(y[2222]), .B(x[2222]), .Z(n13443) );
  XOR U17844 ( .A(y[2221]), .B(x[2221]), .Z(n13444) );
  XOR U17845 ( .A(y[2220]), .B(x[2220]), .Z(n13442) );
  XNOR U17846 ( .A(n13435), .B(n13434), .Z(n13437) );
  XNOR U17847 ( .A(n13431), .B(n13430), .Z(n13434) );
  XOR U17848 ( .A(n13433), .B(n13432), .Z(n13430) );
  XOR U17849 ( .A(y[2219]), .B(x[2219]), .Z(n13432) );
  XOR U17850 ( .A(y[2218]), .B(x[2218]), .Z(n13433) );
  XOR U17851 ( .A(y[2217]), .B(x[2217]), .Z(n13431) );
  XOR U17852 ( .A(n13425), .B(n13424), .Z(n13435) );
  XOR U17853 ( .A(n13427), .B(n13426), .Z(n13424) );
  XOR U17854 ( .A(y[2216]), .B(x[2216]), .Z(n13426) );
  XOR U17855 ( .A(y[2215]), .B(x[2215]), .Z(n13427) );
  XOR U17856 ( .A(y[2214]), .B(x[2214]), .Z(n13425) );
  NAND U17857 ( .A(n13488), .B(n13489), .Z(N29037) );
  NAND U17858 ( .A(n13490), .B(n13491), .Z(n13489) );
  NANDN U17859 ( .A(n13492), .B(n13493), .Z(n13491) );
  NANDN U17860 ( .A(n13493), .B(n13492), .Z(n13488) );
  XOR U17861 ( .A(n13492), .B(n13494), .Z(N29036) );
  XNOR U17862 ( .A(n13490), .B(n13493), .Z(n13494) );
  NAND U17863 ( .A(n13495), .B(n13496), .Z(n13493) );
  NAND U17864 ( .A(n13497), .B(n13498), .Z(n13496) );
  NANDN U17865 ( .A(n13499), .B(n13500), .Z(n13498) );
  NANDN U17866 ( .A(n13500), .B(n13499), .Z(n13495) );
  AND U17867 ( .A(n13501), .B(n13502), .Z(n13490) );
  NAND U17868 ( .A(n13503), .B(n13504), .Z(n13502) );
  OR U17869 ( .A(n13505), .B(n13506), .Z(n13504) );
  NAND U17870 ( .A(n13506), .B(n13505), .Z(n13501) );
  IV U17871 ( .A(n13507), .Z(n13506) );
  AND U17872 ( .A(n13508), .B(n13509), .Z(n13492) );
  NAND U17873 ( .A(n13510), .B(n13511), .Z(n13509) );
  NANDN U17874 ( .A(n13512), .B(n13513), .Z(n13511) );
  NANDN U17875 ( .A(n13513), .B(n13512), .Z(n13508) );
  XOR U17876 ( .A(n13505), .B(n13514), .Z(N29035) );
  XOR U17877 ( .A(n13503), .B(n13507), .Z(n13514) );
  XNOR U17878 ( .A(n13500), .B(n13515), .Z(n13507) );
  XNOR U17879 ( .A(n13497), .B(n13499), .Z(n13515) );
  AND U17880 ( .A(n13516), .B(n13517), .Z(n13499) );
  NANDN U17881 ( .A(n13518), .B(n13519), .Z(n13517) );
  NANDN U17882 ( .A(n13520), .B(n13521), .Z(n13519) );
  IV U17883 ( .A(n13522), .Z(n13521) );
  NAND U17884 ( .A(n13522), .B(n13520), .Z(n13516) );
  AND U17885 ( .A(n13523), .B(n13524), .Z(n13497) );
  NAND U17886 ( .A(n13525), .B(n13526), .Z(n13524) );
  OR U17887 ( .A(n13527), .B(n13528), .Z(n13526) );
  NAND U17888 ( .A(n13528), .B(n13527), .Z(n13523) );
  IV U17889 ( .A(n13529), .Z(n13528) );
  NAND U17890 ( .A(n13530), .B(n13531), .Z(n13500) );
  NANDN U17891 ( .A(n13532), .B(n13533), .Z(n13531) );
  NAND U17892 ( .A(n13534), .B(n13535), .Z(n13533) );
  OR U17893 ( .A(n13535), .B(n13534), .Z(n13530) );
  IV U17894 ( .A(n13536), .Z(n13534) );
  AND U17895 ( .A(n13537), .B(n13538), .Z(n13503) );
  NAND U17896 ( .A(n13539), .B(n13540), .Z(n13538) );
  NANDN U17897 ( .A(n13541), .B(n13542), .Z(n13540) );
  NANDN U17898 ( .A(n13542), .B(n13541), .Z(n13537) );
  XOR U17899 ( .A(n13513), .B(n13543), .Z(n13505) );
  XNOR U17900 ( .A(n13510), .B(n13512), .Z(n13543) );
  AND U17901 ( .A(n13544), .B(n13545), .Z(n13512) );
  NANDN U17902 ( .A(n13546), .B(n13547), .Z(n13545) );
  NANDN U17903 ( .A(n13548), .B(n13549), .Z(n13547) );
  IV U17904 ( .A(n13550), .Z(n13549) );
  NAND U17905 ( .A(n13550), .B(n13548), .Z(n13544) );
  AND U17906 ( .A(n13551), .B(n13552), .Z(n13510) );
  NAND U17907 ( .A(n13553), .B(n13554), .Z(n13552) );
  OR U17908 ( .A(n13555), .B(n13556), .Z(n13554) );
  NAND U17909 ( .A(n13556), .B(n13555), .Z(n13551) );
  IV U17910 ( .A(n13557), .Z(n13556) );
  NAND U17911 ( .A(n13558), .B(n13559), .Z(n13513) );
  NANDN U17912 ( .A(n13560), .B(n13561), .Z(n13559) );
  NAND U17913 ( .A(n13562), .B(n13563), .Z(n13561) );
  OR U17914 ( .A(n13563), .B(n13562), .Z(n13558) );
  IV U17915 ( .A(n13564), .Z(n13562) );
  XOR U17916 ( .A(n13539), .B(n13565), .Z(N29034) );
  XNOR U17917 ( .A(n13542), .B(n13541), .Z(n13565) );
  XNOR U17918 ( .A(n13553), .B(n13566), .Z(n13541) );
  XOR U17919 ( .A(n13557), .B(n13555), .Z(n13566) );
  XOR U17920 ( .A(n13563), .B(n13567), .Z(n13555) );
  XOR U17921 ( .A(n13560), .B(n13564), .Z(n13567) );
  NAND U17922 ( .A(n13568), .B(n13569), .Z(n13564) );
  NAND U17923 ( .A(n13570), .B(n13571), .Z(n13569) );
  NAND U17924 ( .A(n13572), .B(n13573), .Z(n13568) );
  AND U17925 ( .A(n13574), .B(n13575), .Z(n13560) );
  NAND U17926 ( .A(n13576), .B(n13577), .Z(n13575) );
  NAND U17927 ( .A(n13578), .B(n13579), .Z(n13574) );
  NANDN U17928 ( .A(n13580), .B(n13581), .Z(n13563) );
  NANDN U17929 ( .A(n13582), .B(n13583), .Z(n13557) );
  XNOR U17930 ( .A(n13548), .B(n13584), .Z(n13553) );
  XOR U17931 ( .A(n13546), .B(n13550), .Z(n13584) );
  NAND U17932 ( .A(n13585), .B(n13586), .Z(n13550) );
  NAND U17933 ( .A(n13587), .B(n13588), .Z(n13586) );
  NAND U17934 ( .A(n13589), .B(n13590), .Z(n13585) );
  AND U17935 ( .A(n13591), .B(n13592), .Z(n13546) );
  NAND U17936 ( .A(n13593), .B(n13594), .Z(n13592) );
  NAND U17937 ( .A(n13595), .B(n13596), .Z(n13591) );
  AND U17938 ( .A(n13597), .B(n13598), .Z(n13548) );
  NAND U17939 ( .A(n13599), .B(n13600), .Z(n13542) );
  XNOR U17940 ( .A(n13525), .B(n13601), .Z(n13539) );
  XOR U17941 ( .A(n13529), .B(n13527), .Z(n13601) );
  XOR U17942 ( .A(n13535), .B(n13602), .Z(n13527) );
  XOR U17943 ( .A(n13532), .B(n13536), .Z(n13602) );
  NAND U17944 ( .A(n13603), .B(n13604), .Z(n13536) );
  NAND U17945 ( .A(n13605), .B(n13606), .Z(n13604) );
  NAND U17946 ( .A(n13607), .B(n13608), .Z(n13603) );
  AND U17947 ( .A(n13609), .B(n13610), .Z(n13532) );
  NAND U17948 ( .A(n13611), .B(n13612), .Z(n13610) );
  NAND U17949 ( .A(n13613), .B(n13614), .Z(n13609) );
  NANDN U17950 ( .A(n13615), .B(n13616), .Z(n13535) );
  NANDN U17951 ( .A(n13617), .B(n13618), .Z(n13529) );
  XNOR U17952 ( .A(n13520), .B(n13619), .Z(n13525) );
  XOR U17953 ( .A(n13518), .B(n13522), .Z(n13619) );
  NAND U17954 ( .A(n13620), .B(n13621), .Z(n13522) );
  NAND U17955 ( .A(n13622), .B(n13623), .Z(n13621) );
  NAND U17956 ( .A(n13624), .B(n13625), .Z(n13620) );
  AND U17957 ( .A(n13626), .B(n13627), .Z(n13518) );
  NAND U17958 ( .A(n13628), .B(n13629), .Z(n13627) );
  NAND U17959 ( .A(n13630), .B(n13631), .Z(n13626) );
  AND U17960 ( .A(n13632), .B(n13633), .Z(n13520) );
  XOR U17961 ( .A(n13600), .B(n13599), .Z(N29033) );
  XNOR U17962 ( .A(n13618), .B(n13617), .Z(n13599) );
  XNOR U17963 ( .A(n13632), .B(n13633), .Z(n13617) );
  XOR U17964 ( .A(n13629), .B(n13628), .Z(n13633) );
  XOR U17965 ( .A(y[2211]), .B(x[2211]), .Z(n13628) );
  XOR U17966 ( .A(n13631), .B(n13630), .Z(n13629) );
  XOR U17967 ( .A(y[2213]), .B(x[2213]), .Z(n13630) );
  XOR U17968 ( .A(y[2212]), .B(x[2212]), .Z(n13631) );
  XOR U17969 ( .A(n13623), .B(n13622), .Z(n13632) );
  XOR U17970 ( .A(n13625), .B(n13624), .Z(n13622) );
  XOR U17971 ( .A(y[2210]), .B(x[2210]), .Z(n13624) );
  XOR U17972 ( .A(y[2209]), .B(x[2209]), .Z(n13625) );
  XOR U17973 ( .A(y[2208]), .B(x[2208]), .Z(n13623) );
  XNOR U17974 ( .A(n13616), .B(n13615), .Z(n13618) );
  XNOR U17975 ( .A(n13612), .B(n13611), .Z(n13615) );
  XOR U17976 ( .A(n13614), .B(n13613), .Z(n13611) );
  XOR U17977 ( .A(y[2207]), .B(x[2207]), .Z(n13613) );
  XOR U17978 ( .A(y[2206]), .B(x[2206]), .Z(n13614) );
  XOR U17979 ( .A(y[2205]), .B(x[2205]), .Z(n13612) );
  XOR U17980 ( .A(n13606), .B(n13605), .Z(n13616) );
  XOR U17981 ( .A(n13608), .B(n13607), .Z(n13605) );
  XOR U17982 ( .A(y[2204]), .B(x[2204]), .Z(n13607) );
  XOR U17983 ( .A(y[2203]), .B(x[2203]), .Z(n13608) );
  XOR U17984 ( .A(y[2202]), .B(x[2202]), .Z(n13606) );
  XNOR U17985 ( .A(n13583), .B(n13582), .Z(n13600) );
  XNOR U17986 ( .A(n13597), .B(n13598), .Z(n13582) );
  XOR U17987 ( .A(n13594), .B(n13593), .Z(n13598) );
  XOR U17988 ( .A(y[2199]), .B(x[2199]), .Z(n13593) );
  XOR U17989 ( .A(n13596), .B(n13595), .Z(n13594) );
  XOR U17990 ( .A(y[2201]), .B(x[2201]), .Z(n13595) );
  XOR U17991 ( .A(y[2200]), .B(x[2200]), .Z(n13596) );
  XOR U17992 ( .A(n13588), .B(n13587), .Z(n13597) );
  XOR U17993 ( .A(n13590), .B(n13589), .Z(n13587) );
  XOR U17994 ( .A(y[2198]), .B(x[2198]), .Z(n13589) );
  XOR U17995 ( .A(y[2197]), .B(x[2197]), .Z(n13590) );
  XOR U17996 ( .A(y[2196]), .B(x[2196]), .Z(n13588) );
  XNOR U17997 ( .A(n13581), .B(n13580), .Z(n13583) );
  XNOR U17998 ( .A(n13577), .B(n13576), .Z(n13580) );
  XOR U17999 ( .A(n13579), .B(n13578), .Z(n13576) );
  XOR U18000 ( .A(y[2195]), .B(x[2195]), .Z(n13578) );
  XOR U18001 ( .A(y[2194]), .B(x[2194]), .Z(n13579) );
  XOR U18002 ( .A(y[2193]), .B(x[2193]), .Z(n13577) );
  XOR U18003 ( .A(n13571), .B(n13570), .Z(n13581) );
  XOR U18004 ( .A(n13573), .B(n13572), .Z(n13570) );
  XOR U18005 ( .A(y[2192]), .B(x[2192]), .Z(n13572) );
  XOR U18006 ( .A(y[2191]), .B(x[2191]), .Z(n13573) );
  XOR U18007 ( .A(y[2190]), .B(x[2190]), .Z(n13571) );
  NAND U18008 ( .A(n13634), .B(n13635), .Z(N29025) );
  NAND U18009 ( .A(n13636), .B(n13637), .Z(n13635) );
  NANDN U18010 ( .A(n13638), .B(n13639), .Z(n13637) );
  NANDN U18011 ( .A(n13639), .B(n13638), .Z(n13634) );
  XOR U18012 ( .A(n13638), .B(n13640), .Z(N29024) );
  XNOR U18013 ( .A(n13636), .B(n13639), .Z(n13640) );
  NAND U18014 ( .A(n13641), .B(n13642), .Z(n13639) );
  NAND U18015 ( .A(n13643), .B(n13644), .Z(n13642) );
  NANDN U18016 ( .A(n13645), .B(n13646), .Z(n13644) );
  NANDN U18017 ( .A(n13646), .B(n13645), .Z(n13641) );
  AND U18018 ( .A(n13647), .B(n13648), .Z(n13636) );
  NAND U18019 ( .A(n13649), .B(n13650), .Z(n13648) );
  OR U18020 ( .A(n13651), .B(n13652), .Z(n13650) );
  NAND U18021 ( .A(n13652), .B(n13651), .Z(n13647) );
  IV U18022 ( .A(n13653), .Z(n13652) );
  AND U18023 ( .A(n13654), .B(n13655), .Z(n13638) );
  NAND U18024 ( .A(n13656), .B(n13657), .Z(n13655) );
  NANDN U18025 ( .A(n13658), .B(n13659), .Z(n13657) );
  NANDN U18026 ( .A(n13659), .B(n13658), .Z(n13654) );
  XOR U18027 ( .A(n13651), .B(n13660), .Z(N29023) );
  XOR U18028 ( .A(n13649), .B(n13653), .Z(n13660) );
  XNOR U18029 ( .A(n13646), .B(n13661), .Z(n13653) );
  XNOR U18030 ( .A(n13643), .B(n13645), .Z(n13661) );
  AND U18031 ( .A(n13662), .B(n13663), .Z(n13645) );
  NANDN U18032 ( .A(n13664), .B(n13665), .Z(n13663) );
  NANDN U18033 ( .A(n13666), .B(n13667), .Z(n13665) );
  IV U18034 ( .A(n13668), .Z(n13667) );
  NAND U18035 ( .A(n13668), .B(n13666), .Z(n13662) );
  AND U18036 ( .A(n13669), .B(n13670), .Z(n13643) );
  NAND U18037 ( .A(n13671), .B(n13672), .Z(n13670) );
  OR U18038 ( .A(n13673), .B(n13674), .Z(n13672) );
  NAND U18039 ( .A(n13674), .B(n13673), .Z(n13669) );
  IV U18040 ( .A(n13675), .Z(n13674) );
  NAND U18041 ( .A(n13676), .B(n13677), .Z(n13646) );
  NANDN U18042 ( .A(n13678), .B(n13679), .Z(n13677) );
  NAND U18043 ( .A(n13680), .B(n13681), .Z(n13679) );
  OR U18044 ( .A(n13681), .B(n13680), .Z(n13676) );
  IV U18045 ( .A(n13682), .Z(n13680) );
  AND U18046 ( .A(n13683), .B(n13684), .Z(n13649) );
  NAND U18047 ( .A(n13685), .B(n13686), .Z(n13684) );
  NANDN U18048 ( .A(n13687), .B(n13688), .Z(n13686) );
  NANDN U18049 ( .A(n13688), .B(n13687), .Z(n13683) );
  XOR U18050 ( .A(n13659), .B(n13689), .Z(n13651) );
  XNOR U18051 ( .A(n13656), .B(n13658), .Z(n13689) );
  AND U18052 ( .A(n13690), .B(n13691), .Z(n13658) );
  NANDN U18053 ( .A(n13692), .B(n13693), .Z(n13691) );
  NANDN U18054 ( .A(n13694), .B(n13695), .Z(n13693) );
  IV U18055 ( .A(n13696), .Z(n13695) );
  NAND U18056 ( .A(n13696), .B(n13694), .Z(n13690) );
  AND U18057 ( .A(n13697), .B(n13698), .Z(n13656) );
  NAND U18058 ( .A(n13699), .B(n13700), .Z(n13698) );
  OR U18059 ( .A(n13701), .B(n13702), .Z(n13700) );
  NAND U18060 ( .A(n13702), .B(n13701), .Z(n13697) );
  IV U18061 ( .A(n13703), .Z(n13702) );
  NAND U18062 ( .A(n13704), .B(n13705), .Z(n13659) );
  NANDN U18063 ( .A(n13706), .B(n13707), .Z(n13705) );
  NAND U18064 ( .A(n13708), .B(n13709), .Z(n13707) );
  OR U18065 ( .A(n13709), .B(n13708), .Z(n13704) );
  IV U18066 ( .A(n13710), .Z(n13708) );
  XOR U18067 ( .A(n13685), .B(n13711), .Z(N29022) );
  XNOR U18068 ( .A(n13688), .B(n13687), .Z(n13711) );
  XNOR U18069 ( .A(n13699), .B(n13712), .Z(n13687) );
  XOR U18070 ( .A(n13703), .B(n13701), .Z(n13712) );
  XOR U18071 ( .A(n13709), .B(n13713), .Z(n13701) );
  XOR U18072 ( .A(n13706), .B(n13710), .Z(n13713) );
  NAND U18073 ( .A(n13714), .B(n13715), .Z(n13710) );
  NAND U18074 ( .A(n13716), .B(n13717), .Z(n13715) );
  NAND U18075 ( .A(n13718), .B(n13719), .Z(n13714) );
  AND U18076 ( .A(n13720), .B(n13721), .Z(n13706) );
  NAND U18077 ( .A(n13722), .B(n13723), .Z(n13721) );
  NAND U18078 ( .A(n13724), .B(n13725), .Z(n13720) );
  NANDN U18079 ( .A(n13726), .B(n13727), .Z(n13709) );
  NANDN U18080 ( .A(n13728), .B(n13729), .Z(n13703) );
  XNOR U18081 ( .A(n13694), .B(n13730), .Z(n13699) );
  XOR U18082 ( .A(n13692), .B(n13696), .Z(n13730) );
  NAND U18083 ( .A(n13731), .B(n13732), .Z(n13696) );
  NAND U18084 ( .A(n13733), .B(n13734), .Z(n13732) );
  NAND U18085 ( .A(n13735), .B(n13736), .Z(n13731) );
  AND U18086 ( .A(n13737), .B(n13738), .Z(n13692) );
  NAND U18087 ( .A(n13739), .B(n13740), .Z(n13738) );
  NAND U18088 ( .A(n13741), .B(n13742), .Z(n13737) );
  AND U18089 ( .A(n13743), .B(n13744), .Z(n13694) );
  NAND U18090 ( .A(n13745), .B(n13746), .Z(n13688) );
  XNOR U18091 ( .A(n13671), .B(n13747), .Z(n13685) );
  XOR U18092 ( .A(n13675), .B(n13673), .Z(n13747) );
  XOR U18093 ( .A(n13681), .B(n13748), .Z(n13673) );
  XOR U18094 ( .A(n13678), .B(n13682), .Z(n13748) );
  NAND U18095 ( .A(n13749), .B(n13750), .Z(n13682) );
  NAND U18096 ( .A(n13751), .B(n13752), .Z(n13750) );
  NAND U18097 ( .A(n13753), .B(n13754), .Z(n13749) );
  AND U18098 ( .A(n13755), .B(n13756), .Z(n13678) );
  NAND U18099 ( .A(n13757), .B(n13758), .Z(n13756) );
  NAND U18100 ( .A(n13759), .B(n13760), .Z(n13755) );
  NANDN U18101 ( .A(n13761), .B(n13762), .Z(n13681) );
  NANDN U18102 ( .A(n13763), .B(n13764), .Z(n13675) );
  XNOR U18103 ( .A(n13666), .B(n13765), .Z(n13671) );
  XOR U18104 ( .A(n13664), .B(n13668), .Z(n13765) );
  NAND U18105 ( .A(n13766), .B(n13767), .Z(n13668) );
  NAND U18106 ( .A(n13768), .B(n13769), .Z(n13767) );
  NAND U18107 ( .A(n13770), .B(n13771), .Z(n13766) );
  AND U18108 ( .A(n13772), .B(n13773), .Z(n13664) );
  NAND U18109 ( .A(n13774), .B(n13775), .Z(n13773) );
  NAND U18110 ( .A(n13776), .B(n13777), .Z(n13772) );
  AND U18111 ( .A(n13778), .B(n13779), .Z(n13666) );
  XOR U18112 ( .A(n13746), .B(n13745), .Z(N29021) );
  XNOR U18113 ( .A(n13764), .B(n13763), .Z(n13745) );
  XNOR U18114 ( .A(n13778), .B(n13779), .Z(n13763) );
  XOR U18115 ( .A(n13775), .B(n13774), .Z(n13779) );
  XOR U18116 ( .A(y[2187]), .B(x[2187]), .Z(n13774) );
  XOR U18117 ( .A(n13777), .B(n13776), .Z(n13775) );
  XOR U18118 ( .A(y[2189]), .B(x[2189]), .Z(n13776) );
  XOR U18119 ( .A(y[2188]), .B(x[2188]), .Z(n13777) );
  XOR U18120 ( .A(n13769), .B(n13768), .Z(n13778) );
  XOR U18121 ( .A(n13771), .B(n13770), .Z(n13768) );
  XOR U18122 ( .A(y[2186]), .B(x[2186]), .Z(n13770) );
  XOR U18123 ( .A(y[2185]), .B(x[2185]), .Z(n13771) );
  XOR U18124 ( .A(y[2184]), .B(x[2184]), .Z(n13769) );
  XNOR U18125 ( .A(n13762), .B(n13761), .Z(n13764) );
  XNOR U18126 ( .A(n13758), .B(n13757), .Z(n13761) );
  XOR U18127 ( .A(n13760), .B(n13759), .Z(n13757) );
  XOR U18128 ( .A(y[2183]), .B(x[2183]), .Z(n13759) );
  XOR U18129 ( .A(y[2182]), .B(x[2182]), .Z(n13760) );
  XOR U18130 ( .A(y[2181]), .B(x[2181]), .Z(n13758) );
  XOR U18131 ( .A(n13752), .B(n13751), .Z(n13762) );
  XOR U18132 ( .A(n13754), .B(n13753), .Z(n13751) );
  XOR U18133 ( .A(y[2180]), .B(x[2180]), .Z(n13753) );
  XOR U18134 ( .A(y[2179]), .B(x[2179]), .Z(n13754) );
  XOR U18135 ( .A(y[2178]), .B(x[2178]), .Z(n13752) );
  XNOR U18136 ( .A(n13729), .B(n13728), .Z(n13746) );
  XNOR U18137 ( .A(n13743), .B(n13744), .Z(n13728) );
  XOR U18138 ( .A(n13740), .B(n13739), .Z(n13744) );
  XOR U18139 ( .A(y[2175]), .B(x[2175]), .Z(n13739) );
  XOR U18140 ( .A(n13742), .B(n13741), .Z(n13740) );
  XOR U18141 ( .A(y[2177]), .B(x[2177]), .Z(n13741) );
  XOR U18142 ( .A(y[2176]), .B(x[2176]), .Z(n13742) );
  XOR U18143 ( .A(n13734), .B(n13733), .Z(n13743) );
  XOR U18144 ( .A(n13736), .B(n13735), .Z(n13733) );
  XOR U18145 ( .A(y[2174]), .B(x[2174]), .Z(n13735) );
  XOR U18146 ( .A(y[2173]), .B(x[2173]), .Z(n13736) );
  XOR U18147 ( .A(y[2172]), .B(x[2172]), .Z(n13734) );
  XNOR U18148 ( .A(n13727), .B(n13726), .Z(n13729) );
  XNOR U18149 ( .A(n13723), .B(n13722), .Z(n13726) );
  XOR U18150 ( .A(n13725), .B(n13724), .Z(n13722) );
  XOR U18151 ( .A(y[2171]), .B(x[2171]), .Z(n13724) );
  XOR U18152 ( .A(y[2170]), .B(x[2170]), .Z(n13725) );
  XOR U18153 ( .A(y[2169]), .B(x[2169]), .Z(n13723) );
  XOR U18154 ( .A(n13717), .B(n13716), .Z(n13727) );
  XOR U18155 ( .A(n13719), .B(n13718), .Z(n13716) );
  XOR U18156 ( .A(y[2168]), .B(x[2168]), .Z(n13718) );
  XOR U18157 ( .A(y[2167]), .B(x[2167]), .Z(n13719) );
  XOR U18158 ( .A(y[2166]), .B(x[2166]), .Z(n13717) );
  NAND U18159 ( .A(n13780), .B(n13781), .Z(N29013) );
  NAND U18160 ( .A(n13782), .B(n13783), .Z(n13781) );
  NANDN U18161 ( .A(n13784), .B(n13785), .Z(n13783) );
  NANDN U18162 ( .A(n13785), .B(n13784), .Z(n13780) );
  XOR U18163 ( .A(n13784), .B(n13786), .Z(N29012) );
  XNOR U18164 ( .A(n13782), .B(n13785), .Z(n13786) );
  NAND U18165 ( .A(n13787), .B(n13788), .Z(n13785) );
  NAND U18166 ( .A(n13789), .B(n13790), .Z(n13788) );
  NANDN U18167 ( .A(n13791), .B(n13792), .Z(n13790) );
  NANDN U18168 ( .A(n13792), .B(n13791), .Z(n13787) );
  AND U18169 ( .A(n13793), .B(n13794), .Z(n13782) );
  NAND U18170 ( .A(n13795), .B(n13796), .Z(n13794) );
  OR U18171 ( .A(n13797), .B(n13798), .Z(n13796) );
  NAND U18172 ( .A(n13798), .B(n13797), .Z(n13793) );
  IV U18173 ( .A(n13799), .Z(n13798) );
  AND U18174 ( .A(n13800), .B(n13801), .Z(n13784) );
  NAND U18175 ( .A(n13802), .B(n13803), .Z(n13801) );
  NANDN U18176 ( .A(n13804), .B(n13805), .Z(n13803) );
  NANDN U18177 ( .A(n13805), .B(n13804), .Z(n13800) );
  XOR U18178 ( .A(n13797), .B(n13806), .Z(N29011) );
  XOR U18179 ( .A(n13795), .B(n13799), .Z(n13806) );
  XNOR U18180 ( .A(n13792), .B(n13807), .Z(n13799) );
  XNOR U18181 ( .A(n13789), .B(n13791), .Z(n13807) );
  AND U18182 ( .A(n13808), .B(n13809), .Z(n13791) );
  NANDN U18183 ( .A(n13810), .B(n13811), .Z(n13809) );
  NANDN U18184 ( .A(n13812), .B(n13813), .Z(n13811) );
  IV U18185 ( .A(n13814), .Z(n13813) );
  NAND U18186 ( .A(n13814), .B(n13812), .Z(n13808) );
  AND U18187 ( .A(n13815), .B(n13816), .Z(n13789) );
  NAND U18188 ( .A(n13817), .B(n13818), .Z(n13816) );
  OR U18189 ( .A(n13819), .B(n13820), .Z(n13818) );
  NAND U18190 ( .A(n13820), .B(n13819), .Z(n13815) );
  IV U18191 ( .A(n13821), .Z(n13820) );
  NAND U18192 ( .A(n13822), .B(n13823), .Z(n13792) );
  NANDN U18193 ( .A(n13824), .B(n13825), .Z(n13823) );
  NAND U18194 ( .A(n13826), .B(n13827), .Z(n13825) );
  OR U18195 ( .A(n13827), .B(n13826), .Z(n13822) );
  IV U18196 ( .A(n13828), .Z(n13826) );
  AND U18197 ( .A(n13829), .B(n13830), .Z(n13795) );
  NAND U18198 ( .A(n13831), .B(n13832), .Z(n13830) );
  NANDN U18199 ( .A(n13833), .B(n13834), .Z(n13832) );
  NANDN U18200 ( .A(n13834), .B(n13833), .Z(n13829) );
  XOR U18201 ( .A(n13805), .B(n13835), .Z(n13797) );
  XNOR U18202 ( .A(n13802), .B(n13804), .Z(n13835) );
  AND U18203 ( .A(n13836), .B(n13837), .Z(n13804) );
  NANDN U18204 ( .A(n13838), .B(n13839), .Z(n13837) );
  NANDN U18205 ( .A(n13840), .B(n13841), .Z(n13839) );
  IV U18206 ( .A(n13842), .Z(n13841) );
  NAND U18207 ( .A(n13842), .B(n13840), .Z(n13836) );
  AND U18208 ( .A(n13843), .B(n13844), .Z(n13802) );
  NAND U18209 ( .A(n13845), .B(n13846), .Z(n13844) );
  OR U18210 ( .A(n13847), .B(n13848), .Z(n13846) );
  NAND U18211 ( .A(n13848), .B(n13847), .Z(n13843) );
  IV U18212 ( .A(n13849), .Z(n13848) );
  NAND U18213 ( .A(n13850), .B(n13851), .Z(n13805) );
  NANDN U18214 ( .A(n13852), .B(n13853), .Z(n13851) );
  NAND U18215 ( .A(n13854), .B(n13855), .Z(n13853) );
  OR U18216 ( .A(n13855), .B(n13854), .Z(n13850) );
  IV U18217 ( .A(n13856), .Z(n13854) );
  XOR U18218 ( .A(n13831), .B(n13857), .Z(N29010) );
  XNOR U18219 ( .A(n13834), .B(n13833), .Z(n13857) );
  XNOR U18220 ( .A(n13845), .B(n13858), .Z(n13833) );
  XOR U18221 ( .A(n13849), .B(n13847), .Z(n13858) );
  XOR U18222 ( .A(n13855), .B(n13859), .Z(n13847) );
  XOR U18223 ( .A(n13852), .B(n13856), .Z(n13859) );
  NAND U18224 ( .A(n13860), .B(n13861), .Z(n13856) );
  NAND U18225 ( .A(n13862), .B(n13863), .Z(n13861) );
  NAND U18226 ( .A(n13864), .B(n13865), .Z(n13860) );
  AND U18227 ( .A(n13866), .B(n13867), .Z(n13852) );
  NAND U18228 ( .A(n13868), .B(n13869), .Z(n13867) );
  NAND U18229 ( .A(n13870), .B(n13871), .Z(n13866) );
  NANDN U18230 ( .A(n13872), .B(n13873), .Z(n13855) );
  NANDN U18231 ( .A(n13874), .B(n13875), .Z(n13849) );
  XNOR U18232 ( .A(n13840), .B(n13876), .Z(n13845) );
  XOR U18233 ( .A(n13838), .B(n13842), .Z(n13876) );
  NAND U18234 ( .A(n13877), .B(n13878), .Z(n13842) );
  NAND U18235 ( .A(n13879), .B(n13880), .Z(n13878) );
  NAND U18236 ( .A(n13881), .B(n13882), .Z(n13877) );
  AND U18237 ( .A(n13883), .B(n13884), .Z(n13838) );
  NAND U18238 ( .A(n13885), .B(n13886), .Z(n13884) );
  NAND U18239 ( .A(n13887), .B(n13888), .Z(n13883) );
  AND U18240 ( .A(n13889), .B(n13890), .Z(n13840) );
  NAND U18241 ( .A(n13891), .B(n13892), .Z(n13834) );
  XNOR U18242 ( .A(n13817), .B(n13893), .Z(n13831) );
  XOR U18243 ( .A(n13821), .B(n13819), .Z(n13893) );
  XOR U18244 ( .A(n13827), .B(n13894), .Z(n13819) );
  XOR U18245 ( .A(n13824), .B(n13828), .Z(n13894) );
  NAND U18246 ( .A(n13895), .B(n13896), .Z(n13828) );
  NAND U18247 ( .A(n13897), .B(n13898), .Z(n13896) );
  NAND U18248 ( .A(n13899), .B(n13900), .Z(n13895) );
  AND U18249 ( .A(n13901), .B(n13902), .Z(n13824) );
  NAND U18250 ( .A(n13903), .B(n13904), .Z(n13902) );
  NAND U18251 ( .A(n13905), .B(n13906), .Z(n13901) );
  NANDN U18252 ( .A(n13907), .B(n13908), .Z(n13827) );
  NANDN U18253 ( .A(n13909), .B(n13910), .Z(n13821) );
  XNOR U18254 ( .A(n13812), .B(n13911), .Z(n13817) );
  XOR U18255 ( .A(n13810), .B(n13814), .Z(n13911) );
  NAND U18256 ( .A(n13912), .B(n13913), .Z(n13814) );
  NAND U18257 ( .A(n13914), .B(n13915), .Z(n13913) );
  NAND U18258 ( .A(n13916), .B(n13917), .Z(n13912) );
  AND U18259 ( .A(n13918), .B(n13919), .Z(n13810) );
  NAND U18260 ( .A(n13920), .B(n13921), .Z(n13919) );
  NAND U18261 ( .A(n13922), .B(n13923), .Z(n13918) );
  AND U18262 ( .A(n13924), .B(n13925), .Z(n13812) );
  XOR U18263 ( .A(n13892), .B(n13891), .Z(N29009) );
  XNOR U18264 ( .A(n13910), .B(n13909), .Z(n13891) );
  XNOR U18265 ( .A(n13924), .B(n13925), .Z(n13909) );
  XOR U18266 ( .A(n13921), .B(n13920), .Z(n13925) );
  XOR U18267 ( .A(y[2163]), .B(x[2163]), .Z(n13920) );
  XOR U18268 ( .A(n13923), .B(n13922), .Z(n13921) );
  XOR U18269 ( .A(y[2165]), .B(x[2165]), .Z(n13922) );
  XOR U18270 ( .A(y[2164]), .B(x[2164]), .Z(n13923) );
  XOR U18271 ( .A(n13915), .B(n13914), .Z(n13924) );
  XOR U18272 ( .A(n13917), .B(n13916), .Z(n13914) );
  XOR U18273 ( .A(y[2162]), .B(x[2162]), .Z(n13916) );
  XOR U18274 ( .A(y[2161]), .B(x[2161]), .Z(n13917) );
  XOR U18275 ( .A(y[2160]), .B(x[2160]), .Z(n13915) );
  XNOR U18276 ( .A(n13908), .B(n13907), .Z(n13910) );
  XNOR U18277 ( .A(n13904), .B(n13903), .Z(n13907) );
  XOR U18278 ( .A(n13906), .B(n13905), .Z(n13903) );
  XOR U18279 ( .A(y[2159]), .B(x[2159]), .Z(n13905) );
  XOR U18280 ( .A(y[2158]), .B(x[2158]), .Z(n13906) );
  XOR U18281 ( .A(y[2157]), .B(x[2157]), .Z(n13904) );
  XOR U18282 ( .A(n13898), .B(n13897), .Z(n13908) );
  XOR U18283 ( .A(n13900), .B(n13899), .Z(n13897) );
  XOR U18284 ( .A(y[2156]), .B(x[2156]), .Z(n13899) );
  XOR U18285 ( .A(y[2155]), .B(x[2155]), .Z(n13900) );
  XOR U18286 ( .A(y[2154]), .B(x[2154]), .Z(n13898) );
  XNOR U18287 ( .A(n13875), .B(n13874), .Z(n13892) );
  XNOR U18288 ( .A(n13889), .B(n13890), .Z(n13874) );
  XOR U18289 ( .A(n13886), .B(n13885), .Z(n13890) );
  XOR U18290 ( .A(y[2151]), .B(x[2151]), .Z(n13885) );
  XOR U18291 ( .A(n13888), .B(n13887), .Z(n13886) );
  XOR U18292 ( .A(y[2153]), .B(x[2153]), .Z(n13887) );
  XOR U18293 ( .A(y[2152]), .B(x[2152]), .Z(n13888) );
  XOR U18294 ( .A(n13880), .B(n13879), .Z(n13889) );
  XOR U18295 ( .A(n13882), .B(n13881), .Z(n13879) );
  XOR U18296 ( .A(y[2150]), .B(x[2150]), .Z(n13881) );
  XOR U18297 ( .A(y[2149]), .B(x[2149]), .Z(n13882) );
  XOR U18298 ( .A(y[2148]), .B(x[2148]), .Z(n13880) );
  XNOR U18299 ( .A(n13873), .B(n13872), .Z(n13875) );
  XNOR U18300 ( .A(n13869), .B(n13868), .Z(n13872) );
  XOR U18301 ( .A(n13871), .B(n13870), .Z(n13868) );
  XOR U18302 ( .A(y[2147]), .B(x[2147]), .Z(n13870) );
  XOR U18303 ( .A(y[2146]), .B(x[2146]), .Z(n13871) );
  XOR U18304 ( .A(y[2145]), .B(x[2145]), .Z(n13869) );
  XOR U18305 ( .A(n13863), .B(n13862), .Z(n13873) );
  XOR U18306 ( .A(n13865), .B(n13864), .Z(n13862) );
  XOR U18307 ( .A(y[2144]), .B(x[2144]), .Z(n13864) );
  XOR U18308 ( .A(y[2143]), .B(x[2143]), .Z(n13865) );
  XOR U18309 ( .A(y[2142]), .B(x[2142]), .Z(n13863) );
  NAND U18310 ( .A(n13926), .B(n13927), .Z(N29001) );
  NAND U18311 ( .A(n13928), .B(n13929), .Z(n13927) );
  NANDN U18312 ( .A(n13930), .B(n13931), .Z(n13929) );
  NANDN U18313 ( .A(n13931), .B(n13930), .Z(n13926) );
  XOR U18314 ( .A(n13930), .B(n13932), .Z(N29000) );
  XNOR U18315 ( .A(n13928), .B(n13931), .Z(n13932) );
  NAND U18316 ( .A(n13933), .B(n13934), .Z(n13931) );
  NAND U18317 ( .A(n13935), .B(n13936), .Z(n13934) );
  NANDN U18318 ( .A(n13937), .B(n13938), .Z(n13936) );
  NANDN U18319 ( .A(n13938), .B(n13937), .Z(n13933) );
  AND U18320 ( .A(n13939), .B(n13940), .Z(n13928) );
  NAND U18321 ( .A(n13941), .B(n13942), .Z(n13940) );
  OR U18322 ( .A(n13943), .B(n13944), .Z(n13942) );
  NAND U18323 ( .A(n13944), .B(n13943), .Z(n13939) );
  IV U18324 ( .A(n13945), .Z(n13944) );
  AND U18325 ( .A(n13946), .B(n13947), .Z(n13930) );
  NAND U18326 ( .A(n13948), .B(n13949), .Z(n13947) );
  NANDN U18327 ( .A(n13950), .B(n13951), .Z(n13949) );
  NANDN U18328 ( .A(n13951), .B(n13950), .Z(n13946) );
  XOR U18329 ( .A(n13943), .B(n13952), .Z(N28999) );
  XOR U18330 ( .A(n13941), .B(n13945), .Z(n13952) );
  XNOR U18331 ( .A(n13938), .B(n13953), .Z(n13945) );
  XNOR U18332 ( .A(n13935), .B(n13937), .Z(n13953) );
  AND U18333 ( .A(n13954), .B(n13955), .Z(n13937) );
  NANDN U18334 ( .A(n13956), .B(n13957), .Z(n13955) );
  NANDN U18335 ( .A(n13958), .B(n13959), .Z(n13957) );
  IV U18336 ( .A(n13960), .Z(n13959) );
  NAND U18337 ( .A(n13960), .B(n13958), .Z(n13954) );
  AND U18338 ( .A(n13961), .B(n13962), .Z(n13935) );
  NAND U18339 ( .A(n13963), .B(n13964), .Z(n13962) );
  OR U18340 ( .A(n13965), .B(n13966), .Z(n13964) );
  NAND U18341 ( .A(n13966), .B(n13965), .Z(n13961) );
  IV U18342 ( .A(n13967), .Z(n13966) );
  NAND U18343 ( .A(n13968), .B(n13969), .Z(n13938) );
  NANDN U18344 ( .A(n13970), .B(n13971), .Z(n13969) );
  NAND U18345 ( .A(n13972), .B(n13973), .Z(n13971) );
  OR U18346 ( .A(n13973), .B(n13972), .Z(n13968) );
  IV U18347 ( .A(n13974), .Z(n13972) );
  AND U18348 ( .A(n13975), .B(n13976), .Z(n13941) );
  NAND U18349 ( .A(n13977), .B(n13978), .Z(n13976) );
  NANDN U18350 ( .A(n13979), .B(n13980), .Z(n13978) );
  NANDN U18351 ( .A(n13980), .B(n13979), .Z(n13975) );
  XOR U18352 ( .A(n13951), .B(n13981), .Z(n13943) );
  XNOR U18353 ( .A(n13948), .B(n13950), .Z(n13981) );
  AND U18354 ( .A(n13982), .B(n13983), .Z(n13950) );
  NANDN U18355 ( .A(n13984), .B(n13985), .Z(n13983) );
  NANDN U18356 ( .A(n13986), .B(n13987), .Z(n13985) );
  IV U18357 ( .A(n13988), .Z(n13987) );
  NAND U18358 ( .A(n13988), .B(n13986), .Z(n13982) );
  AND U18359 ( .A(n13989), .B(n13990), .Z(n13948) );
  NAND U18360 ( .A(n13991), .B(n13992), .Z(n13990) );
  OR U18361 ( .A(n13993), .B(n13994), .Z(n13992) );
  NAND U18362 ( .A(n13994), .B(n13993), .Z(n13989) );
  IV U18363 ( .A(n13995), .Z(n13994) );
  NAND U18364 ( .A(n13996), .B(n13997), .Z(n13951) );
  NANDN U18365 ( .A(n13998), .B(n13999), .Z(n13997) );
  NAND U18366 ( .A(n14000), .B(n14001), .Z(n13999) );
  OR U18367 ( .A(n14001), .B(n14000), .Z(n13996) );
  IV U18368 ( .A(n14002), .Z(n14000) );
  XOR U18369 ( .A(n13977), .B(n14003), .Z(N28998) );
  XNOR U18370 ( .A(n13980), .B(n13979), .Z(n14003) );
  XNOR U18371 ( .A(n13991), .B(n14004), .Z(n13979) );
  XOR U18372 ( .A(n13995), .B(n13993), .Z(n14004) );
  XOR U18373 ( .A(n14001), .B(n14005), .Z(n13993) );
  XOR U18374 ( .A(n13998), .B(n14002), .Z(n14005) );
  NAND U18375 ( .A(n14006), .B(n14007), .Z(n14002) );
  NAND U18376 ( .A(n14008), .B(n14009), .Z(n14007) );
  NAND U18377 ( .A(n14010), .B(n14011), .Z(n14006) );
  AND U18378 ( .A(n14012), .B(n14013), .Z(n13998) );
  NAND U18379 ( .A(n14014), .B(n14015), .Z(n14013) );
  NAND U18380 ( .A(n14016), .B(n14017), .Z(n14012) );
  NANDN U18381 ( .A(n14018), .B(n14019), .Z(n14001) );
  NANDN U18382 ( .A(n14020), .B(n14021), .Z(n13995) );
  XNOR U18383 ( .A(n13986), .B(n14022), .Z(n13991) );
  XOR U18384 ( .A(n13984), .B(n13988), .Z(n14022) );
  NAND U18385 ( .A(n14023), .B(n14024), .Z(n13988) );
  NAND U18386 ( .A(n14025), .B(n14026), .Z(n14024) );
  NAND U18387 ( .A(n14027), .B(n14028), .Z(n14023) );
  AND U18388 ( .A(n14029), .B(n14030), .Z(n13984) );
  NAND U18389 ( .A(n14031), .B(n14032), .Z(n14030) );
  NAND U18390 ( .A(n14033), .B(n14034), .Z(n14029) );
  AND U18391 ( .A(n14035), .B(n14036), .Z(n13986) );
  NAND U18392 ( .A(n14037), .B(n14038), .Z(n13980) );
  XNOR U18393 ( .A(n13963), .B(n14039), .Z(n13977) );
  XOR U18394 ( .A(n13967), .B(n13965), .Z(n14039) );
  XOR U18395 ( .A(n13973), .B(n14040), .Z(n13965) );
  XOR U18396 ( .A(n13970), .B(n13974), .Z(n14040) );
  NAND U18397 ( .A(n14041), .B(n14042), .Z(n13974) );
  NAND U18398 ( .A(n14043), .B(n14044), .Z(n14042) );
  NAND U18399 ( .A(n14045), .B(n14046), .Z(n14041) );
  AND U18400 ( .A(n14047), .B(n14048), .Z(n13970) );
  NAND U18401 ( .A(n14049), .B(n14050), .Z(n14048) );
  NAND U18402 ( .A(n14051), .B(n14052), .Z(n14047) );
  NANDN U18403 ( .A(n14053), .B(n14054), .Z(n13973) );
  NANDN U18404 ( .A(n14055), .B(n14056), .Z(n13967) );
  XNOR U18405 ( .A(n13958), .B(n14057), .Z(n13963) );
  XOR U18406 ( .A(n13956), .B(n13960), .Z(n14057) );
  NAND U18407 ( .A(n14058), .B(n14059), .Z(n13960) );
  NAND U18408 ( .A(n14060), .B(n14061), .Z(n14059) );
  NAND U18409 ( .A(n14062), .B(n14063), .Z(n14058) );
  AND U18410 ( .A(n14064), .B(n14065), .Z(n13956) );
  NAND U18411 ( .A(n14066), .B(n14067), .Z(n14065) );
  NAND U18412 ( .A(n14068), .B(n14069), .Z(n14064) );
  AND U18413 ( .A(n14070), .B(n14071), .Z(n13958) );
  XOR U18414 ( .A(n14038), .B(n14037), .Z(N28997) );
  XNOR U18415 ( .A(n14056), .B(n14055), .Z(n14037) );
  XNOR U18416 ( .A(n14070), .B(n14071), .Z(n14055) );
  XOR U18417 ( .A(n14067), .B(n14066), .Z(n14071) );
  XOR U18418 ( .A(y[2139]), .B(x[2139]), .Z(n14066) );
  XOR U18419 ( .A(n14069), .B(n14068), .Z(n14067) );
  XOR U18420 ( .A(y[2141]), .B(x[2141]), .Z(n14068) );
  XOR U18421 ( .A(y[2140]), .B(x[2140]), .Z(n14069) );
  XOR U18422 ( .A(n14061), .B(n14060), .Z(n14070) );
  XOR U18423 ( .A(n14063), .B(n14062), .Z(n14060) );
  XOR U18424 ( .A(y[2138]), .B(x[2138]), .Z(n14062) );
  XOR U18425 ( .A(y[2137]), .B(x[2137]), .Z(n14063) );
  XOR U18426 ( .A(y[2136]), .B(x[2136]), .Z(n14061) );
  XNOR U18427 ( .A(n14054), .B(n14053), .Z(n14056) );
  XNOR U18428 ( .A(n14050), .B(n14049), .Z(n14053) );
  XOR U18429 ( .A(n14052), .B(n14051), .Z(n14049) );
  XOR U18430 ( .A(y[2135]), .B(x[2135]), .Z(n14051) );
  XOR U18431 ( .A(y[2134]), .B(x[2134]), .Z(n14052) );
  XOR U18432 ( .A(y[2133]), .B(x[2133]), .Z(n14050) );
  XOR U18433 ( .A(n14044), .B(n14043), .Z(n14054) );
  XOR U18434 ( .A(n14046), .B(n14045), .Z(n14043) );
  XOR U18435 ( .A(y[2132]), .B(x[2132]), .Z(n14045) );
  XOR U18436 ( .A(y[2131]), .B(x[2131]), .Z(n14046) );
  XOR U18437 ( .A(y[2130]), .B(x[2130]), .Z(n14044) );
  XNOR U18438 ( .A(n14021), .B(n14020), .Z(n14038) );
  XNOR U18439 ( .A(n14035), .B(n14036), .Z(n14020) );
  XOR U18440 ( .A(n14032), .B(n14031), .Z(n14036) );
  XOR U18441 ( .A(y[2127]), .B(x[2127]), .Z(n14031) );
  XOR U18442 ( .A(n14034), .B(n14033), .Z(n14032) );
  XOR U18443 ( .A(y[2129]), .B(x[2129]), .Z(n14033) );
  XOR U18444 ( .A(y[2128]), .B(x[2128]), .Z(n14034) );
  XOR U18445 ( .A(n14026), .B(n14025), .Z(n14035) );
  XOR U18446 ( .A(n14028), .B(n14027), .Z(n14025) );
  XOR U18447 ( .A(y[2126]), .B(x[2126]), .Z(n14027) );
  XOR U18448 ( .A(y[2125]), .B(x[2125]), .Z(n14028) );
  XOR U18449 ( .A(y[2124]), .B(x[2124]), .Z(n14026) );
  XNOR U18450 ( .A(n14019), .B(n14018), .Z(n14021) );
  XNOR U18451 ( .A(n14015), .B(n14014), .Z(n14018) );
  XOR U18452 ( .A(n14017), .B(n14016), .Z(n14014) );
  XOR U18453 ( .A(y[2123]), .B(x[2123]), .Z(n14016) );
  XOR U18454 ( .A(y[2122]), .B(x[2122]), .Z(n14017) );
  XOR U18455 ( .A(y[2121]), .B(x[2121]), .Z(n14015) );
  XOR U18456 ( .A(n14009), .B(n14008), .Z(n14019) );
  XOR U18457 ( .A(n14011), .B(n14010), .Z(n14008) );
  XOR U18458 ( .A(y[2120]), .B(x[2120]), .Z(n14010) );
  XOR U18459 ( .A(y[2119]), .B(x[2119]), .Z(n14011) );
  XOR U18460 ( .A(y[2118]), .B(x[2118]), .Z(n14009) );
  NAND U18461 ( .A(n14072), .B(n14073), .Z(N28989) );
  NAND U18462 ( .A(n14074), .B(n14075), .Z(n14073) );
  NANDN U18463 ( .A(n14076), .B(n14077), .Z(n14075) );
  NANDN U18464 ( .A(n14077), .B(n14076), .Z(n14072) );
  XOR U18465 ( .A(n14076), .B(n14078), .Z(N28988) );
  XNOR U18466 ( .A(n14074), .B(n14077), .Z(n14078) );
  NAND U18467 ( .A(n14079), .B(n14080), .Z(n14077) );
  NAND U18468 ( .A(n14081), .B(n14082), .Z(n14080) );
  NANDN U18469 ( .A(n14083), .B(n14084), .Z(n14082) );
  NANDN U18470 ( .A(n14084), .B(n14083), .Z(n14079) );
  AND U18471 ( .A(n14085), .B(n14086), .Z(n14074) );
  NAND U18472 ( .A(n14087), .B(n14088), .Z(n14086) );
  OR U18473 ( .A(n14089), .B(n14090), .Z(n14088) );
  NAND U18474 ( .A(n14090), .B(n14089), .Z(n14085) );
  IV U18475 ( .A(n14091), .Z(n14090) );
  AND U18476 ( .A(n14092), .B(n14093), .Z(n14076) );
  NAND U18477 ( .A(n14094), .B(n14095), .Z(n14093) );
  NANDN U18478 ( .A(n14096), .B(n14097), .Z(n14095) );
  NANDN U18479 ( .A(n14097), .B(n14096), .Z(n14092) );
  XOR U18480 ( .A(n14089), .B(n14098), .Z(N28987) );
  XOR U18481 ( .A(n14087), .B(n14091), .Z(n14098) );
  XNOR U18482 ( .A(n14084), .B(n14099), .Z(n14091) );
  XNOR U18483 ( .A(n14081), .B(n14083), .Z(n14099) );
  AND U18484 ( .A(n14100), .B(n14101), .Z(n14083) );
  NANDN U18485 ( .A(n14102), .B(n14103), .Z(n14101) );
  NANDN U18486 ( .A(n14104), .B(n14105), .Z(n14103) );
  IV U18487 ( .A(n14106), .Z(n14105) );
  NAND U18488 ( .A(n14106), .B(n14104), .Z(n14100) );
  AND U18489 ( .A(n14107), .B(n14108), .Z(n14081) );
  NAND U18490 ( .A(n14109), .B(n14110), .Z(n14108) );
  OR U18491 ( .A(n14111), .B(n14112), .Z(n14110) );
  NAND U18492 ( .A(n14112), .B(n14111), .Z(n14107) );
  IV U18493 ( .A(n14113), .Z(n14112) );
  NAND U18494 ( .A(n14114), .B(n14115), .Z(n14084) );
  NANDN U18495 ( .A(n14116), .B(n14117), .Z(n14115) );
  NAND U18496 ( .A(n14118), .B(n14119), .Z(n14117) );
  OR U18497 ( .A(n14119), .B(n14118), .Z(n14114) );
  IV U18498 ( .A(n14120), .Z(n14118) );
  AND U18499 ( .A(n14121), .B(n14122), .Z(n14087) );
  NAND U18500 ( .A(n14123), .B(n14124), .Z(n14122) );
  NANDN U18501 ( .A(n14125), .B(n14126), .Z(n14124) );
  NANDN U18502 ( .A(n14126), .B(n14125), .Z(n14121) );
  XOR U18503 ( .A(n14097), .B(n14127), .Z(n14089) );
  XNOR U18504 ( .A(n14094), .B(n14096), .Z(n14127) );
  AND U18505 ( .A(n14128), .B(n14129), .Z(n14096) );
  NANDN U18506 ( .A(n14130), .B(n14131), .Z(n14129) );
  NANDN U18507 ( .A(n14132), .B(n14133), .Z(n14131) );
  IV U18508 ( .A(n14134), .Z(n14133) );
  NAND U18509 ( .A(n14134), .B(n14132), .Z(n14128) );
  AND U18510 ( .A(n14135), .B(n14136), .Z(n14094) );
  NAND U18511 ( .A(n14137), .B(n14138), .Z(n14136) );
  OR U18512 ( .A(n14139), .B(n14140), .Z(n14138) );
  NAND U18513 ( .A(n14140), .B(n14139), .Z(n14135) );
  IV U18514 ( .A(n14141), .Z(n14140) );
  NAND U18515 ( .A(n14142), .B(n14143), .Z(n14097) );
  NANDN U18516 ( .A(n14144), .B(n14145), .Z(n14143) );
  NAND U18517 ( .A(n14146), .B(n14147), .Z(n14145) );
  OR U18518 ( .A(n14147), .B(n14146), .Z(n14142) );
  IV U18519 ( .A(n14148), .Z(n14146) );
  XOR U18520 ( .A(n14123), .B(n14149), .Z(N28986) );
  XNOR U18521 ( .A(n14126), .B(n14125), .Z(n14149) );
  XNOR U18522 ( .A(n14137), .B(n14150), .Z(n14125) );
  XOR U18523 ( .A(n14141), .B(n14139), .Z(n14150) );
  XOR U18524 ( .A(n14147), .B(n14151), .Z(n14139) );
  XOR U18525 ( .A(n14144), .B(n14148), .Z(n14151) );
  NAND U18526 ( .A(n14152), .B(n14153), .Z(n14148) );
  NAND U18527 ( .A(n14154), .B(n14155), .Z(n14153) );
  NAND U18528 ( .A(n14156), .B(n14157), .Z(n14152) );
  AND U18529 ( .A(n14158), .B(n14159), .Z(n14144) );
  NAND U18530 ( .A(n14160), .B(n14161), .Z(n14159) );
  NAND U18531 ( .A(n14162), .B(n14163), .Z(n14158) );
  NANDN U18532 ( .A(n14164), .B(n14165), .Z(n14147) );
  NANDN U18533 ( .A(n14166), .B(n14167), .Z(n14141) );
  XNOR U18534 ( .A(n14132), .B(n14168), .Z(n14137) );
  XOR U18535 ( .A(n14130), .B(n14134), .Z(n14168) );
  NAND U18536 ( .A(n14169), .B(n14170), .Z(n14134) );
  NAND U18537 ( .A(n14171), .B(n14172), .Z(n14170) );
  NAND U18538 ( .A(n14173), .B(n14174), .Z(n14169) );
  AND U18539 ( .A(n14175), .B(n14176), .Z(n14130) );
  NAND U18540 ( .A(n14177), .B(n14178), .Z(n14176) );
  NAND U18541 ( .A(n14179), .B(n14180), .Z(n14175) );
  AND U18542 ( .A(n14181), .B(n14182), .Z(n14132) );
  NAND U18543 ( .A(n14183), .B(n14184), .Z(n14126) );
  XNOR U18544 ( .A(n14109), .B(n14185), .Z(n14123) );
  XOR U18545 ( .A(n14113), .B(n14111), .Z(n14185) );
  XOR U18546 ( .A(n14119), .B(n14186), .Z(n14111) );
  XOR U18547 ( .A(n14116), .B(n14120), .Z(n14186) );
  NAND U18548 ( .A(n14187), .B(n14188), .Z(n14120) );
  NAND U18549 ( .A(n14189), .B(n14190), .Z(n14188) );
  NAND U18550 ( .A(n14191), .B(n14192), .Z(n14187) );
  AND U18551 ( .A(n14193), .B(n14194), .Z(n14116) );
  NAND U18552 ( .A(n14195), .B(n14196), .Z(n14194) );
  NAND U18553 ( .A(n14197), .B(n14198), .Z(n14193) );
  NANDN U18554 ( .A(n14199), .B(n14200), .Z(n14119) );
  NANDN U18555 ( .A(n14201), .B(n14202), .Z(n14113) );
  XNOR U18556 ( .A(n14104), .B(n14203), .Z(n14109) );
  XOR U18557 ( .A(n14102), .B(n14106), .Z(n14203) );
  NAND U18558 ( .A(n14204), .B(n14205), .Z(n14106) );
  NAND U18559 ( .A(n14206), .B(n14207), .Z(n14205) );
  NAND U18560 ( .A(n14208), .B(n14209), .Z(n14204) );
  AND U18561 ( .A(n14210), .B(n14211), .Z(n14102) );
  NAND U18562 ( .A(n14212), .B(n14213), .Z(n14211) );
  NAND U18563 ( .A(n14214), .B(n14215), .Z(n14210) );
  AND U18564 ( .A(n14216), .B(n14217), .Z(n14104) );
  XOR U18565 ( .A(n14184), .B(n14183), .Z(N28985) );
  XNOR U18566 ( .A(n14202), .B(n14201), .Z(n14183) );
  XNOR U18567 ( .A(n14216), .B(n14217), .Z(n14201) );
  XOR U18568 ( .A(n14213), .B(n14212), .Z(n14217) );
  XOR U18569 ( .A(y[2115]), .B(x[2115]), .Z(n14212) );
  XOR U18570 ( .A(n14215), .B(n14214), .Z(n14213) );
  XOR U18571 ( .A(y[2117]), .B(x[2117]), .Z(n14214) );
  XOR U18572 ( .A(y[2116]), .B(x[2116]), .Z(n14215) );
  XOR U18573 ( .A(n14207), .B(n14206), .Z(n14216) );
  XOR U18574 ( .A(n14209), .B(n14208), .Z(n14206) );
  XOR U18575 ( .A(y[2114]), .B(x[2114]), .Z(n14208) );
  XOR U18576 ( .A(y[2113]), .B(x[2113]), .Z(n14209) );
  XOR U18577 ( .A(y[2112]), .B(x[2112]), .Z(n14207) );
  XNOR U18578 ( .A(n14200), .B(n14199), .Z(n14202) );
  XNOR U18579 ( .A(n14196), .B(n14195), .Z(n14199) );
  XOR U18580 ( .A(n14198), .B(n14197), .Z(n14195) );
  XOR U18581 ( .A(y[2111]), .B(x[2111]), .Z(n14197) );
  XOR U18582 ( .A(y[2110]), .B(x[2110]), .Z(n14198) );
  XOR U18583 ( .A(y[2109]), .B(x[2109]), .Z(n14196) );
  XOR U18584 ( .A(n14190), .B(n14189), .Z(n14200) );
  XOR U18585 ( .A(n14192), .B(n14191), .Z(n14189) );
  XOR U18586 ( .A(y[2108]), .B(x[2108]), .Z(n14191) );
  XOR U18587 ( .A(y[2107]), .B(x[2107]), .Z(n14192) );
  XOR U18588 ( .A(y[2106]), .B(x[2106]), .Z(n14190) );
  XNOR U18589 ( .A(n14167), .B(n14166), .Z(n14184) );
  XNOR U18590 ( .A(n14181), .B(n14182), .Z(n14166) );
  XOR U18591 ( .A(n14178), .B(n14177), .Z(n14182) );
  XOR U18592 ( .A(y[2103]), .B(x[2103]), .Z(n14177) );
  XOR U18593 ( .A(n14180), .B(n14179), .Z(n14178) );
  XOR U18594 ( .A(y[2105]), .B(x[2105]), .Z(n14179) );
  XOR U18595 ( .A(y[2104]), .B(x[2104]), .Z(n14180) );
  XOR U18596 ( .A(n14172), .B(n14171), .Z(n14181) );
  XOR U18597 ( .A(n14174), .B(n14173), .Z(n14171) );
  XOR U18598 ( .A(y[2102]), .B(x[2102]), .Z(n14173) );
  XOR U18599 ( .A(y[2101]), .B(x[2101]), .Z(n14174) );
  XOR U18600 ( .A(y[2100]), .B(x[2100]), .Z(n14172) );
  XNOR U18601 ( .A(n14165), .B(n14164), .Z(n14167) );
  XNOR U18602 ( .A(n14161), .B(n14160), .Z(n14164) );
  XOR U18603 ( .A(n14163), .B(n14162), .Z(n14160) );
  XOR U18604 ( .A(y[2099]), .B(x[2099]), .Z(n14162) );
  XOR U18605 ( .A(y[2098]), .B(x[2098]), .Z(n14163) );
  XOR U18606 ( .A(y[2097]), .B(x[2097]), .Z(n14161) );
  XOR U18607 ( .A(n14155), .B(n14154), .Z(n14165) );
  XOR U18608 ( .A(n14157), .B(n14156), .Z(n14154) );
  XOR U18609 ( .A(y[2096]), .B(x[2096]), .Z(n14156) );
  XOR U18610 ( .A(y[2095]), .B(x[2095]), .Z(n14157) );
  XOR U18611 ( .A(y[2094]), .B(x[2094]), .Z(n14155) );
  NAND U18612 ( .A(n14218), .B(n14219), .Z(N28977) );
  NAND U18613 ( .A(n14220), .B(n14221), .Z(n14219) );
  NANDN U18614 ( .A(n14222), .B(n14223), .Z(n14221) );
  NANDN U18615 ( .A(n14223), .B(n14222), .Z(n14218) );
  XOR U18616 ( .A(n14222), .B(n14224), .Z(N28976) );
  XNOR U18617 ( .A(n14220), .B(n14223), .Z(n14224) );
  NAND U18618 ( .A(n14225), .B(n14226), .Z(n14223) );
  NAND U18619 ( .A(n14227), .B(n14228), .Z(n14226) );
  NANDN U18620 ( .A(n14229), .B(n14230), .Z(n14228) );
  NANDN U18621 ( .A(n14230), .B(n14229), .Z(n14225) );
  AND U18622 ( .A(n14231), .B(n14232), .Z(n14220) );
  NAND U18623 ( .A(n14233), .B(n14234), .Z(n14232) );
  OR U18624 ( .A(n14235), .B(n14236), .Z(n14234) );
  NAND U18625 ( .A(n14236), .B(n14235), .Z(n14231) );
  IV U18626 ( .A(n14237), .Z(n14236) );
  AND U18627 ( .A(n14238), .B(n14239), .Z(n14222) );
  NAND U18628 ( .A(n14240), .B(n14241), .Z(n14239) );
  NANDN U18629 ( .A(n14242), .B(n14243), .Z(n14241) );
  NANDN U18630 ( .A(n14243), .B(n14242), .Z(n14238) );
  XOR U18631 ( .A(n14235), .B(n14244), .Z(N28975) );
  XOR U18632 ( .A(n14233), .B(n14237), .Z(n14244) );
  XNOR U18633 ( .A(n14230), .B(n14245), .Z(n14237) );
  XNOR U18634 ( .A(n14227), .B(n14229), .Z(n14245) );
  AND U18635 ( .A(n14246), .B(n14247), .Z(n14229) );
  NANDN U18636 ( .A(n14248), .B(n14249), .Z(n14247) );
  NANDN U18637 ( .A(n14250), .B(n14251), .Z(n14249) );
  IV U18638 ( .A(n14252), .Z(n14251) );
  NAND U18639 ( .A(n14252), .B(n14250), .Z(n14246) );
  AND U18640 ( .A(n14253), .B(n14254), .Z(n14227) );
  NAND U18641 ( .A(n14255), .B(n14256), .Z(n14254) );
  OR U18642 ( .A(n14257), .B(n14258), .Z(n14256) );
  NAND U18643 ( .A(n14258), .B(n14257), .Z(n14253) );
  IV U18644 ( .A(n14259), .Z(n14258) );
  NAND U18645 ( .A(n14260), .B(n14261), .Z(n14230) );
  NANDN U18646 ( .A(n14262), .B(n14263), .Z(n14261) );
  NAND U18647 ( .A(n14264), .B(n14265), .Z(n14263) );
  OR U18648 ( .A(n14265), .B(n14264), .Z(n14260) );
  IV U18649 ( .A(n14266), .Z(n14264) );
  AND U18650 ( .A(n14267), .B(n14268), .Z(n14233) );
  NAND U18651 ( .A(n14269), .B(n14270), .Z(n14268) );
  NANDN U18652 ( .A(n14271), .B(n14272), .Z(n14270) );
  NANDN U18653 ( .A(n14272), .B(n14271), .Z(n14267) );
  XOR U18654 ( .A(n14243), .B(n14273), .Z(n14235) );
  XNOR U18655 ( .A(n14240), .B(n14242), .Z(n14273) );
  AND U18656 ( .A(n14274), .B(n14275), .Z(n14242) );
  NANDN U18657 ( .A(n14276), .B(n14277), .Z(n14275) );
  NANDN U18658 ( .A(n14278), .B(n14279), .Z(n14277) );
  IV U18659 ( .A(n14280), .Z(n14279) );
  NAND U18660 ( .A(n14280), .B(n14278), .Z(n14274) );
  AND U18661 ( .A(n14281), .B(n14282), .Z(n14240) );
  NAND U18662 ( .A(n14283), .B(n14284), .Z(n14282) );
  OR U18663 ( .A(n14285), .B(n14286), .Z(n14284) );
  NAND U18664 ( .A(n14286), .B(n14285), .Z(n14281) );
  IV U18665 ( .A(n14287), .Z(n14286) );
  NAND U18666 ( .A(n14288), .B(n14289), .Z(n14243) );
  NANDN U18667 ( .A(n14290), .B(n14291), .Z(n14289) );
  NAND U18668 ( .A(n14292), .B(n14293), .Z(n14291) );
  OR U18669 ( .A(n14293), .B(n14292), .Z(n14288) );
  IV U18670 ( .A(n14294), .Z(n14292) );
  XOR U18671 ( .A(n14269), .B(n14295), .Z(N28974) );
  XNOR U18672 ( .A(n14272), .B(n14271), .Z(n14295) );
  XNOR U18673 ( .A(n14283), .B(n14296), .Z(n14271) );
  XOR U18674 ( .A(n14287), .B(n14285), .Z(n14296) );
  XOR U18675 ( .A(n14293), .B(n14297), .Z(n14285) );
  XOR U18676 ( .A(n14290), .B(n14294), .Z(n14297) );
  NAND U18677 ( .A(n14298), .B(n14299), .Z(n14294) );
  NAND U18678 ( .A(n14300), .B(n14301), .Z(n14299) );
  NAND U18679 ( .A(n14302), .B(n14303), .Z(n14298) );
  AND U18680 ( .A(n14304), .B(n14305), .Z(n14290) );
  NAND U18681 ( .A(n14306), .B(n14307), .Z(n14305) );
  NAND U18682 ( .A(n14308), .B(n14309), .Z(n14304) );
  NANDN U18683 ( .A(n14310), .B(n14311), .Z(n14293) );
  NANDN U18684 ( .A(n14312), .B(n14313), .Z(n14287) );
  XNOR U18685 ( .A(n14278), .B(n14314), .Z(n14283) );
  XOR U18686 ( .A(n14276), .B(n14280), .Z(n14314) );
  NAND U18687 ( .A(n14315), .B(n14316), .Z(n14280) );
  NAND U18688 ( .A(n14317), .B(n14318), .Z(n14316) );
  NAND U18689 ( .A(n14319), .B(n14320), .Z(n14315) );
  AND U18690 ( .A(n14321), .B(n14322), .Z(n14276) );
  NAND U18691 ( .A(n14323), .B(n14324), .Z(n14322) );
  NAND U18692 ( .A(n14325), .B(n14326), .Z(n14321) );
  AND U18693 ( .A(n14327), .B(n14328), .Z(n14278) );
  NAND U18694 ( .A(n14329), .B(n14330), .Z(n14272) );
  XNOR U18695 ( .A(n14255), .B(n14331), .Z(n14269) );
  XOR U18696 ( .A(n14259), .B(n14257), .Z(n14331) );
  XOR U18697 ( .A(n14265), .B(n14332), .Z(n14257) );
  XOR U18698 ( .A(n14262), .B(n14266), .Z(n14332) );
  NAND U18699 ( .A(n14333), .B(n14334), .Z(n14266) );
  NAND U18700 ( .A(n14335), .B(n14336), .Z(n14334) );
  NAND U18701 ( .A(n14337), .B(n14338), .Z(n14333) );
  AND U18702 ( .A(n14339), .B(n14340), .Z(n14262) );
  NAND U18703 ( .A(n14341), .B(n14342), .Z(n14340) );
  NAND U18704 ( .A(n14343), .B(n14344), .Z(n14339) );
  NANDN U18705 ( .A(n14345), .B(n14346), .Z(n14265) );
  NANDN U18706 ( .A(n14347), .B(n14348), .Z(n14259) );
  XNOR U18707 ( .A(n14250), .B(n14349), .Z(n14255) );
  XOR U18708 ( .A(n14248), .B(n14252), .Z(n14349) );
  NAND U18709 ( .A(n14350), .B(n14351), .Z(n14252) );
  NAND U18710 ( .A(n14352), .B(n14353), .Z(n14351) );
  NAND U18711 ( .A(n14354), .B(n14355), .Z(n14350) );
  AND U18712 ( .A(n14356), .B(n14357), .Z(n14248) );
  NAND U18713 ( .A(n14358), .B(n14359), .Z(n14357) );
  NAND U18714 ( .A(n14360), .B(n14361), .Z(n14356) );
  AND U18715 ( .A(n14362), .B(n14363), .Z(n14250) );
  XOR U18716 ( .A(n14330), .B(n14329), .Z(N28973) );
  XNOR U18717 ( .A(n14348), .B(n14347), .Z(n14329) );
  XNOR U18718 ( .A(n14362), .B(n14363), .Z(n14347) );
  XOR U18719 ( .A(n14359), .B(n14358), .Z(n14363) );
  XOR U18720 ( .A(y[2091]), .B(x[2091]), .Z(n14358) );
  XOR U18721 ( .A(n14361), .B(n14360), .Z(n14359) );
  XOR U18722 ( .A(y[2093]), .B(x[2093]), .Z(n14360) );
  XOR U18723 ( .A(y[2092]), .B(x[2092]), .Z(n14361) );
  XOR U18724 ( .A(n14353), .B(n14352), .Z(n14362) );
  XOR U18725 ( .A(n14355), .B(n14354), .Z(n14352) );
  XOR U18726 ( .A(y[2090]), .B(x[2090]), .Z(n14354) );
  XOR U18727 ( .A(y[2089]), .B(x[2089]), .Z(n14355) );
  XOR U18728 ( .A(y[2088]), .B(x[2088]), .Z(n14353) );
  XNOR U18729 ( .A(n14346), .B(n14345), .Z(n14348) );
  XNOR U18730 ( .A(n14342), .B(n14341), .Z(n14345) );
  XOR U18731 ( .A(n14344), .B(n14343), .Z(n14341) );
  XOR U18732 ( .A(y[2087]), .B(x[2087]), .Z(n14343) );
  XOR U18733 ( .A(y[2086]), .B(x[2086]), .Z(n14344) );
  XOR U18734 ( .A(y[2085]), .B(x[2085]), .Z(n14342) );
  XOR U18735 ( .A(n14336), .B(n14335), .Z(n14346) );
  XOR U18736 ( .A(n14338), .B(n14337), .Z(n14335) );
  XOR U18737 ( .A(y[2084]), .B(x[2084]), .Z(n14337) );
  XOR U18738 ( .A(y[2083]), .B(x[2083]), .Z(n14338) );
  XOR U18739 ( .A(y[2082]), .B(x[2082]), .Z(n14336) );
  XNOR U18740 ( .A(n14313), .B(n14312), .Z(n14330) );
  XNOR U18741 ( .A(n14327), .B(n14328), .Z(n14312) );
  XOR U18742 ( .A(n14324), .B(n14323), .Z(n14328) );
  XOR U18743 ( .A(y[2079]), .B(x[2079]), .Z(n14323) );
  XOR U18744 ( .A(n14326), .B(n14325), .Z(n14324) );
  XOR U18745 ( .A(y[2081]), .B(x[2081]), .Z(n14325) );
  XOR U18746 ( .A(y[2080]), .B(x[2080]), .Z(n14326) );
  XOR U18747 ( .A(n14318), .B(n14317), .Z(n14327) );
  XOR U18748 ( .A(n14320), .B(n14319), .Z(n14317) );
  XOR U18749 ( .A(y[2078]), .B(x[2078]), .Z(n14319) );
  XOR U18750 ( .A(y[2077]), .B(x[2077]), .Z(n14320) );
  XOR U18751 ( .A(y[2076]), .B(x[2076]), .Z(n14318) );
  XNOR U18752 ( .A(n14311), .B(n14310), .Z(n14313) );
  XNOR U18753 ( .A(n14307), .B(n14306), .Z(n14310) );
  XOR U18754 ( .A(n14309), .B(n14308), .Z(n14306) );
  XOR U18755 ( .A(y[2075]), .B(x[2075]), .Z(n14308) );
  XOR U18756 ( .A(y[2074]), .B(x[2074]), .Z(n14309) );
  XOR U18757 ( .A(y[2073]), .B(x[2073]), .Z(n14307) );
  XOR U18758 ( .A(n14301), .B(n14300), .Z(n14311) );
  XOR U18759 ( .A(n14303), .B(n14302), .Z(n14300) );
  XOR U18760 ( .A(y[2072]), .B(x[2072]), .Z(n14302) );
  XOR U18761 ( .A(y[2071]), .B(x[2071]), .Z(n14303) );
  XOR U18762 ( .A(y[2070]), .B(x[2070]), .Z(n14301) );
  NAND U18763 ( .A(n14364), .B(n14365), .Z(N28965) );
  NAND U18764 ( .A(n14366), .B(n14367), .Z(n14365) );
  NANDN U18765 ( .A(n14368), .B(n14369), .Z(n14367) );
  NANDN U18766 ( .A(n14369), .B(n14368), .Z(n14364) );
  XOR U18767 ( .A(n14368), .B(n14370), .Z(N28964) );
  XNOR U18768 ( .A(n14366), .B(n14369), .Z(n14370) );
  NAND U18769 ( .A(n14371), .B(n14372), .Z(n14369) );
  NAND U18770 ( .A(n14373), .B(n14374), .Z(n14372) );
  NANDN U18771 ( .A(n14375), .B(n14376), .Z(n14374) );
  NANDN U18772 ( .A(n14376), .B(n14375), .Z(n14371) );
  AND U18773 ( .A(n14377), .B(n14378), .Z(n14366) );
  NAND U18774 ( .A(n14379), .B(n14380), .Z(n14378) );
  OR U18775 ( .A(n14381), .B(n14382), .Z(n14380) );
  NAND U18776 ( .A(n14382), .B(n14381), .Z(n14377) );
  IV U18777 ( .A(n14383), .Z(n14382) );
  AND U18778 ( .A(n14384), .B(n14385), .Z(n14368) );
  NAND U18779 ( .A(n14386), .B(n14387), .Z(n14385) );
  NANDN U18780 ( .A(n14388), .B(n14389), .Z(n14387) );
  NANDN U18781 ( .A(n14389), .B(n14388), .Z(n14384) );
  XOR U18782 ( .A(n14381), .B(n14390), .Z(N28963) );
  XOR U18783 ( .A(n14379), .B(n14383), .Z(n14390) );
  XNOR U18784 ( .A(n14376), .B(n14391), .Z(n14383) );
  XNOR U18785 ( .A(n14373), .B(n14375), .Z(n14391) );
  AND U18786 ( .A(n14392), .B(n14393), .Z(n14375) );
  NANDN U18787 ( .A(n14394), .B(n14395), .Z(n14393) );
  NANDN U18788 ( .A(n14396), .B(n14397), .Z(n14395) );
  IV U18789 ( .A(n14398), .Z(n14397) );
  NAND U18790 ( .A(n14398), .B(n14396), .Z(n14392) );
  AND U18791 ( .A(n14399), .B(n14400), .Z(n14373) );
  NAND U18792 ( .A(n14401), .B(n14402), .Z(n14400) );
  OR U18793 ( .A(n14403), .B(n14404), .Z(n14402) );
  NAND U18794 ( .A(n14404), .B(n14403), .Z(n14399) );
  IV U18795 ( .A(n14405), .Z(n14404) );
  NAND U18796 ( .A(n14406), .B(n14407), .Z(n14376) );
  NANDN U18797 ( .A(n14408), .B(n14409), .Z(n14407) );
  NAND U18798 ( .A(n14410), .B(n14411), .Z(n14409) );
  OR U18799 ( .A(n14411), .B(n14410), .Z(n14406) );
  IV U18800 ( .A(n14412), .Z(n14410) );
  AND U18801 ( .A(n14413), .B(n14414), .Z(n14379) );
  NAND U18802 ( .A(n14415), .B(n14416), .Z(n14414) );
  NANDN U18803 ( .A(n14417), .B(n14418), .Z(n14416) );
  NANDN U18804 ( .A(n14418), .B(n14417), .Z(n14413) );
  XOR U18805 ( .A(n14389), .B(n14419), .Z(n14381) );
  XNOR U18806 ( .A(n14386), .B(n14388), .Z(n14419) );
  AND U18807 ( .A(n14420), .B(n14421), .Z(n14388) );
  NANDN U18808 ( .A(n14422), .B(n14423), .Z(n14421) );
  NANDN U18809 ( .A(n14424), .B(n14425), .Z(n14423) );
  IV U18810 ( .A(n14426), .Z(n14425) );
  NAND U18811 ( .A(n14426), .B(n14424), .Z(n14420) );
  AND U18812 ( .A(n14427), .B(n14428), .Z(n14386) );
  NAND U18813 ( .A(n14429), .B(n14430), .Z(n14428) );
  OR U18814 ( .A(n14431), .B(n14432), .Z(n14430) );
  NAND U18815 ( .A(n14432), .B(n14431), .Z(n14427) );
  IV U18816 ( .A(n14433), .Z(n14432) );
  NAND U18817 ( .A(n14434), .B(n14435), .Z(n14389) );
  NANDN U18818 ( .A(n14436), .B(n14437), .Z(n14435) );
  NAND U18819 ( .A(n14438), .B(n14439), .Z(n14437) );
  OR U18820 ( .A(n14439), .B(n14438), .Z(n14434) );
  IV U18821 ( .A(n14440), .Z(n14438) );
  XOR U18822 ( .A(n14415), .B(n14441), .Z(N28962) );
  XNOR U18823 ( .A(n14418), .B(n14417), .Z(n14441) );
  XNOR U18824 ( .A(n14429), .B(n14442), .Z(n14417) );
  XOR U18825 ( .A(n14433), .B(n14431), .Z(n14442) );
  XOR U18826 ( .A(n14439), .B(n14443), .Z(n14431) );
  XOR U18827 ( .A(n14436), .B(n14440), .Z(n14443) );
  NAND U18828 ( .A(n14444), .B(n14445), .Z(n14440) );
  NAND U18829 ( .A(n14446), .B(n14447), .Z(n14445) );
  NAND U18830 ( .A(n14448), .B(n14449), .Z(n14444) );
  AND U18831 ( .A(n14450), .B(n14451), .Z(n14436) );
  NAND U18832 ( .A(n14452), .B(n14453), .Z(n14451) );
  NAND U18833 ( .A(n14454), .B(n14455), .Z(n14450) );
  NANDN U18834 ( .A(n14456), .B(n14457), .Z(n14439) );
  NANDN U18835 ( .A(n14458), .B(n14459), .Z(n14433) );
  XNOR U18836 ( .A(n14424), .B(n14460), .Z(n14429) );
  XOR U18837 ( .A(n14422), .B(n14426), .Z(n14460) );
  NAND U18838 ( .A(n14461), .B(n14462), .Z(n14426) );
  NAND U18839 ( .A(n14463), .B(n14464), .Z(n14462) );
  NAND U18840 ( .A(n14465), .B(n14466), .Z(n14461) );
  AND U18841 ( .A(n14467), .B(n14468), .Z(n14422) );
  NAND U18842 ( .A(n14469), .B(n14470), .Z(n14468) );
  NAND U18843 ( .A(n14471), .B(n14472), .Z(n14467) );
  AND U18844 ( .A(n14473), .B(n14474), .Z(n14424) );
  NAND U18845 ( .A(n14475), .B(n14476), .Z(n14418) );
  XNOR U18846 ( .A(n14401), .B(n14477), .Z(n14415) );
  XOR U18847 ( .A(n14405), .B(n14403), .Z(n14477) );
  XOR U18848 ( .A(n14411), .B(n14478), .Z(n14403) );
  XOR U18849 ( .A(n14408), .B(n14412), .Z(n14478) );
  NAND U18850 ( .A(n14479), .B(n14480), .Z(n14412) );
  NAND U18851 ( .A(n14481), .B(n14482), .Z(n14480) );
  NAND U18852 ( .A(n14483), .B(n14484), .Z(n14479) );
  AND U18853 ( .A(n14485), .B(n14486), .Z(n14408) );
  NAND U18854 ( .A(n14487), .B(n14488), .Z(n14486) );
  NAND U18855 ( .A(n14489), .B(n14490), .Z(n14485) );
  NANDN U18856 ( .A(n14491), .B(n14492), .Z(n14411) );
  NANDN U18857 ( .A(n14493), .B(n14494), .Z(n14405) );
  XNOR U18858 ( .A(n14396), .B(n14495), .Z(n14401) );
  XOR U18859 ( .A(n14394), .B(n14398), .Z(n14495) );
  NAND U18860 ( .A(n14496), .B(n14497), .Z(n14398) );
  NAND U18861 ( .A(n14498), .B(n14499), .Z(n14497) );
  NAND U18862 ( .A(n14500), .B(n14501), .Z(n14496) );
  AND U18863 ( .A(n14502), .B(n14503), .Z(n14394) );
  NAND U18864 ( .A(n14504), .B(n14505), .Z(n14503) );
  NAND U18865 ( .A(n14506), .B(n14507), .Z(n14502) );
  AND U18866 ( .A(n14508), .B(n14509), .Z(n14396) );
  XOR U18867 ( .A(n14476), .B(n14475), .Z(N28961) );
  XNOR U18868 ( .A(n14494), .B(n14493), .Z(n14475) );
  XNOR U18869 ( .A(n14508), .B(n14509), .Z(n14493) );
  XOR U18870 ( .A(n14505), .B(n14504), .Z(n14509) );
  XOR U18871 ( .A(y[2067]), .B(x[2067]), .Z(n14504) );
  XOR U18872 ( .A(n14507), .B(n14506), .Z(n14505) );
  XOR U18873 ( .A(y[2069]), .B(x[2069]), .Z(n14506) );
  XOR U18874 ( .A(y[2068]), .B(x[2068]), .Z(n14507) );
  XOR U18875 ( .A(n14499), .B(n14498), .Z(n14508) );
  XOR U18876 ( .A(n14501), .B(n14500), .Z(n14498) );
  XOR U18877 ( .A(y[2066]), .B(x[2066]), .Z(n14500) );
  XOR U18878 ( .A(y[2065]), .B(x[2065]), .Z(n14501) );
  XOR U18879 ( .A(y[2064]), .B(x[2064]), .Z(n14499) );
  XNOR U18880 ( .A(n14492), .B(n14491), .Z(n14494) );
  XNOR U18881 ( .A(n14488), .B(n14487), .Z(n14491) );
  XOR U18882 ( .A(n14490), .B(n14489), .Z(n14487) );
  XOR U18883 ( .A(y[2063]), .B(x[2063]), .Z(n14489) );
  XOR U18884 ( .A(y[2062]), .B(x[2062]), .Z(n14490) );
  XOR U18885 ( .A(y[2061]), .B(x[2061]), .Z(n14488) );
  XOR U18886 ( .A(n14482), .B(n14481), .Z(n14492) );
  XOR U18887 ( .A(n14484), .B(n14483), .Z(n14481) );
  XOR U18888 ( .A(y[2060]), .B(x[2060]), .Z(n14483) );
  XOR U18889 ( .A(y[2059]), .B(x[2059]), .Z(n14484) );
  XOR U18890 ( .A(y[2058]), .B(x[2058]), .Z(n14482) );
  XNOR U18891 ( .A(n14459), .B(n14458), .Z(n14476) );
  XNOR U18892 ( .A(n14473), .B(n14474), .Z(n14458) );
  XOR U18893 ( .A(n14470), .B(n14469), .Z(n14474) );
  XOR U18894 ( .A(y[2055]), .B(x[2055]), .Z(n14469) );
  XOR U18895 ( .A(n14472), .B(n14471), .Z(n14470) );
  XOR U18896 ( .A(y[2057]), .B(x[2057]), .Z(n14471) );
  XOR U18897 ( .A(y[2056]), .B(x[2056]), .Z(n14472) );
  XOR U18898 ( .A(n14464), .B(n14463), .Z(n14473) );
  XOR U18899 ( .A(n14466), .B(n14465), .Z(n14463) );
  XOR U18900 ( .A(y[2054]), .B(x[2054]), .Z(n14465) );
  XOR U18901 ( .A(y[2053]), .B(x[2053]), .Z(n14466) );
  XOR U18902 ( .A(y[2052]), .B(x[2052]), .Z(n14464) );
  XNOR U18903 ( .A(n14457), .B(n14456), .Z(n14459) );
  XNOR U18904 ( .A(n14453), .B(n14452), .Z(n14456) );
  XOR U18905 ( .A(n14455), .B(n14454), .Z(n14452) );
  XOR U18906 ( .A(y[2051]), .B(x[2051]), .Z(n14454) );
  XOR U18907 ( .A(y[2050]), .B(x[2050]), .Z(n14455) );
  XOR U18908 ( .A(y[2049]), .B(x[2049]), .Z(n14453) );
  XOR U18909 ( .A(n14447), .B(n14446), .Z(n14457) );
  XOR U18910 ( .A(n14449), .B(n14448), .Z(n14446) );
  XOR U18911 ( .A(y[2048]), .B(x[2048]), .Z(n14448) );
  XOR U18912 ( .A(y[2047]), .B(x[2047]), .Z(n14449) );
  XOR U18913 ( .A(y[2046]), .B(x[2046]), .Z(n14447) );
  NAND U18914 ( .A(n14510), .B(n14511), .Z(N28953) );
  NAND U18915 ( .A(n14512), .B(n14513), .Z(n14511) );
  NANDN U18916 ( .A(n14514), .B(n14515), .Z(n14513) );
  NANDN U18917 ( .A(n14515), .B(n14514), .Z(n14510) );
  XOR U18918 ( .A(n14514), .B(n14516), .Z(N28952) );
  XNOR U18919 ( .A(n14512), .B(n14515), .Z(n14516) );
  NAND U18920 ( .A(n14517), .B(n14518), .Z(n14515) );
  NAND U18921 ( .A(n14519), .B(n14520), .Z(n14518) );
  NANDN U18922 ( .A(n14521), .B(n14522), .Z(n14520) );
  NANDN U18923 ( .A(n14522), .B(n14521), .Z(n14517) );
  AND U18924 ( .A(n14523), .B(n14524), .Z(n14512) );
  NAND U18925 ( .A(n14525), .B(n14526), .Z(n14524) );
  OR U18926 ( .A(n14527), .B(n14528), .Z(n14526) );
  NAND U18927 ( .A(n14528), .B(n14527), .Z(n14523) );
  IV U18928 ( .A(n14529), .Z(n14528) );
  AND U18929 ( .A(n14530), .B(n14531), .Z(n14514) );
  NAND U18930 ( .A(n14532), .B(n14533), .Z(n14531) );
  NANDN U18931 ( .A(n14534), .B(n14535), .Z(n14533) );
  NANDN U18932 ( .A(n14535), .B(n14534), .Z(n14530) );
  XOR U18933 ( .A(n14527), .B(n14536), .Z(N28951) );
  XOR U18934 ( .A(n14525), .B(n14529), .Z(n14536) );
  XNOR U18935 ( .A(n14522), .B(n14537), .Z(n14529) );
  XNOR U18936 ( .A(n14519), .B(n14521), .Z(n14537) );
  AND U18937 ( .A(n14538), .B(n14539), .Z(n14521) );
  NANDN U18938 ( .A(n14540), .B(n14541), .Z(n14539) );
  NANDN U18939 ( .A(n14542), .B(n14543), .Z(n14541) );
  IV U18940 ( .A(n14544), .Z(n14543) );
  NAND U18941 ( .A(n14544), .B(n14542), .Z(n14538) );
  AND U18942 ( .A(n14545), .B(n14546), .Z(n14519) );
  NAND U18943 ( .A(n14547), .B(n14548), .Z(n14546) );
  OR U18944 ( .A(n14549), .B(n14550), .Z(n14548) );
  NAND U18945 ( .A(n14550), .B(n14549), .Z(n14545) );
  IV U18946 ( .A(n14551), .Z(n14550) );
  NAND U18947 ( .A(n14552), .B(n14553), .Z(n14522) );
  NANDN U18948 ( .A(n14554), .B(n14555), .Z(n14553) );
  NAND U18949 ( .A(n14556), .B(n14557), .Z(n14555) );
  OR U18950 ( .A(n14557), .B(n14556), .Z(n14552) );
  IV U18951 ( .A(n14558), .Z(n14556) );
  AND U18952 ( .A(n14559), .B(n14560), .Z(n14525) );
  NAND U18953 ( .A(n14561), .B(n14562), .Z(n14560) );
  NANDN U18954 ( .A(n14563), .B(n14564), .Z(n14562) );
  NANDN U18955 ( .A(n14564), .B(n14563), .Z(n14559) );
  XOR U18956 ( .A(n14535), .B(n14565), .Z(n14527) );
  XNOR U18957 ( .A(n14532), .B(n14534), .Z(n14565) );
  AND U18958 ( .A(n14566), .B(n14567), .Z(n14534) );
  NANDN U18959 ( .A(n14568), .B(n14569), .Z(n14567) );
  NANDN U18960 ( .A(n14570), .B(n14571), .Z(n14569) );
  IV U18961 ( .A(n14572), .Z(n14571) );
  NAND U18962 ( .A(n14572), .B(n14570), .Z(n14566) );
  AND U18963 ( .A(n14573), .B(n14574), .Z(n14532) );
  NAND U18964 ( .A(n14575), .B(n14576), .Z(n14574) );
  OR U18965 ( .A(n14577), .B(n14578), .Z(n14576) );
  NAND U18966 ( .A(n14578), .B(n14577), .Z(n14573) );
  IV U18967 ( .A(n14579), .Z(n14578) );
  NAND U18968 ( .A(n14580), .B(n14581), .Z(n14535) );
  NANDN U18969 ( .A(n14582), .B(n14583), .Z(n14581) );
  NAND U18970 ( .A(n14584), .B(n14585), .Z(n14583) );
  OR U18971 ( .A(n14585), .B(n14584), .Z(n14580) );
  IV U18972 ( .A(n14586), .Z(n14584) );
  XOR U18973 ( .A(n14561), .B(n14587), .Z(N28950) );
  XNOR U18974 ( .A(n14564), .B(n14563), .Z(n14587) );
  XNOR U18975 ( .A(n14575), .B(n14588), .Z(n14563) );
  XOR U18976 ( .A(n14579), .B(n14577), .Z(n14588) );
  XOR U18977 ( .A(n14585), .B(n14589), .Z(n14577) );
  XOR U18978 ( .A(n14582), .B(n14586), .Z(n14589) );
  NAND U18979 ( .A(n14590), .B(n14591), .Z(n14586) );
  NAND U18980 ( .A(n14592), .B(n14593), .Z(n14591) );
  NAND U18981 ( .A(n14594), .B(n14595), .Z(n14590) );
  AND U18982 ( .A(n14596), .B(n14597), .Z(n14582) );
  NAND U18983 ( .A(n14598), .B(n14599), .Z(n14597) );
  NAND U18984 ( .A(n14600), .B(n14601), .Z(n14596) );
  NANDN U18985 ( .A(n14602), .B(n14603), .Z(n14585) );
  NANDN U18986 ( .A(n14604), .B(n14605), .Z(n14579) );
  XNOR U18987 ( .A(n14570), .B(n14606), .Z(n14575) );
  XOR U18988 ( .A(n14568), .B(n14572), .Z(n14606) );
  NAND U18989 ( .A(n14607), .B(n14608), .Z(n14572) );
  NAND U18990 ( .A(n14609), .B(n14610), .Z(n14608) );
  NAND U18991 ( .A(n14611), .B(n14612), .Z(n14607) );
  AND U18992 ( .A(n14613), .B(n14614), .Z(n14568) );
  NAND U18993 ( .A(n14615), .B(n14616), .Z(n14614) );
  NAND U18994 ( .A(n14617), .B(n14618), .Z(n14613) );
  AND U18995 ( .A(n14619), .B(n14620), .Z(n14570) );
  NAND U18996 ( .A(n14621), .B(n14622), .Z(n14564) );
  XNOR U18997 ( .A(n14547), .B(n14623), .Z(n14561) );
  XOR U18998 ( .A(n14551), .B(n14549), .Z(n14623) );
  XOR U18999 ( .A(n14557), .B(n14624), .Z(n14549) );
  XOR U19000 ( .A(n14554), .B(n14558), .Z(n14624) );
  NAND U19001 ( .A(n14625), .B(n14626), .Z(n14558) );
  NAND U19002 ( .A(n14627), .B(n14628), .Z(n14626) );
  NAND U19003 ( .A(n14629), .B(n14630), .Z(n14625) );
  AND U19004 ( .A(n14631), .B(n14632), .Z(n14554) );
  NAND U19005 ( .A(n14633), .B(n14634), .Z(n14632) );
  NAND U19006 ( .A(n14635), .B(n14636), .Z(n14631) );
  NANDN U19007 ( .A(n14637), .B(n14638), .Z(n14557) );
  NANDN U19008 ( .A(n14639), .B(n14640), .Z(n14551) );
  XNOR U19009 ( .A(n14542), .B(n14641), .Z(n14547) );
  XOR U19010 ( .A(n14540), .B(n14544), .Z(n14641) );
  NAND U19011 ( .A(n14642), .B(n14643), .Z(n14544) );
  NAND U19012 ( .A(n14644), .B(n14645), .Z(n14643) );
  NAND U19013 ( .A(n14646), .B(n14647), .Z(n14642) );
  AND U19014 ( .A(n14648), .B(n14649), .Z(n14540) );
  NAND U19015 ( .A(n14650), .B(n14651), .Z(n14649) );
  NAND U19016 ( .A(n14652), .B(n14653), .Z(n14648) );
  AND U19017 ( .A(n14654), .B(n14655), .Z(n14542) );
  XOR U19018 ( .A(n14622), .B(n14621), .Z(N28949) );
  XNOR U19019 ( .A(n14640), .B(n14639), .Z(n14621) );
  XNOR U19020 ( .A(n14654), .B(n14655), .Z(n14639) );
  XOR U19021 ( .A(n14651), .B(n14650), .Z(n14655) );
  XOR U19022 ( .A(y[2043]), .B(x[2043]), .Z(n14650) );
  XOR U19023 ( .A(n14653), .B(n14652), .Z(n14651) );
  XOR U19024 ( .A(y[2045]), .B(x[2045]), .Z(n14652) );
  XOR U19025 ( .A(y[2044]), .B(x[2044]), .Z(n14653) );
  XOR U19026 ( .A(n14645), .B(n14644), .Z(n14654) );
  XOR U19027 ( .A(n14647), .B(n14646), .Z(n14644) );
  XOR U19028 ( .A(y[2042]), .B(x[2042]), .Z(n14646) );
  XOR U19029 ( .A(y[2041]), .B(x[2041]), .Z(n14647) );
  XOR U19030 ( .A(y[2040]), .B(x[2040]), .Z(n14645) );
  XNOR U19031 ( .A(n14638), .B(n14637), .Z(n14640) );
  XNOR U19032 ( .A(n14634), .B(n14633), .Z(n14637) );
  XOR U19033 ( .A(n14636), .B(n14635), .Z(n14633) );
  XOR U19034 ( .A(y[2039]), .B(x[2039]), .Z(n14635) );
  XOR U19035 ( .A(y[2038]), .B(x[2038]), .Z(n14636) );
  XOR U19036 ( .A(y[2037]), .B(x[2037]), .Z(n14634) );
  XOR U19037 ( .A(n14628), .B(n14627), .Z(n14638) );
  XOR U19038 ( .A(n14630), .B(n14629), .Z(n14627) );
  XOR U19039 ( .A(y[2036]), .B(x[2036]), .Z(n14629) );
  XOR U19040 ( .A(y[2035]), .B(x[2035]), .Z(n14630) );
  XOR U19041 ( .A(y[2034]), .B(x[2034]), .Z(n14628) );
  XNOR U19042 ( .A(n14605), .B(n14604), .Z(n14622) );
  XNOR U19043 ( .A(n14619), .B(n14620), .Z(n14604) );
  XOR U19044 ( .A(n14616), .B(n14615), .Z(n14620) );
  XOR U19045 ( .A(y[2031]), .B(x[2031]), .Z(n14615) );
  XOR U19046 ( .A(n14618), .B(n14617), .Z(n14616) );
  XOR U19047 ( .A(y[2033]), .B(x[2033]), .Z(n14617) );
  XOR U19048 ( .A(y[2032]), .B(x[2032]), .Z(n14618) );
  XOR U19049 ( .A(n14610), .B(n14609), .Z(n14619) );
  XOR U19050 ( .A(n14612), .B(n14611), .Z(n14609) );
  XOR U19051 ( .A(y[2030]), .B(x[2030]), .Z(n14611) );
  XOR U19052 ( .A(y[2029]), .B(x[2029]), .Z(n14612) );
  XOR U19053 ( .A(y[2028]), .B(x[2028]), .Z(n14610) );
  XNOR U19054 ( .A(n14603), .B(n14602), .Z(n14605) );
  XNOR U19055 ( .A(n14599), .B(n14598), .Z(n14602) );
  XOR U19056 ( .A(n14601), .B(n14600), .Z(n14598) );
  XOR U19057 ( .A(y[2027]), .B(x[2027]), .Z(n14600) );
  XOR U19058 ( .A(y[2026]), .B(x[2026]), .Z(n14601) );
  XOR U19059 ( .A(y[2025]), .B(x[2025]), .Z(n14599) );
  XOR U19060 ( .A(n14593), .B(n14592), .Z(n14603) );
  XOR U19061 ( .A(n14595), .B(n14594), .Z(n14592) );
  XOR U19062 ( .A(y[2024]), .B(x[2024]), .Z(n14594) );
  XOR U19063 ( .A(y[2023]), .B(x[2023]), .Z(n14595) );
  XOR U19064 ( .A(y[2022]), .B(x[2022]), .Z(n14593) );
  NAND U19065 ( .A(n14656), .B(n14657), .Z(N28941) );
  NAND U19066 ( .A(n14658), .B(n14659), .Z(n14657) );
  NANDN U19067 ( .A(n14660), .B(n14661), .Z(n14659) );
  NANDN U19068 ( .A(n14661), .B(n14660), .Z(n14656) );
  XOR U19069 ( .A(n14660), .B(n14662), .Z(N28940) );
  XNOR U19070 ( .A(n14658), .B(n14661), .Z(n14662) );
  NAND U19071 ( .A(n14663), .B(n14664), .Z(n14661) );
  NAND U19072 ( .A(n14665), .B(n14666), .Z(n14664) );
  NANDN U19073 ( .A(n14667), .B(n14668), .Z(n14666) );
  NANDN U19074 ( .A(n14668), .B(n14667), .Z(n14663) );
  AND U19075 ( .A(n14669), .B(n14670), .Z(n14658) );
  NAND U19076 ( .A(n14671), .B(n14672), .Z(n14670) );
  OR U19077 ( .A(n14673), .B(n14674), .Z(n14672) );
  NAND U19078 ( .A(n14674), .B(n14673), .Z(n14669) );
  IV U19079 ( .A(n14675), .Z(n14674) );
  AND U19080 ( .A(n14676), .B(n14677), .Z(n14660) );
  NAND U19081 ( .A(n14678), .B(n14679), .Z(n14677) );
  NANDN U19082 ( .A(n14680), .B(n14681), .Z(n14679) );
  NANDN U19083 ( .A(n14681), .B(n14680), .Z(n14676) );
  XOR U19084 ( .A(n14673), .B(n14682), .Z(N28939) );
  XOR U19085 ( .A(n14671), .B(n14675), .Z(n14682) );
  XNOR U19086 ( .A(n14668), .B(n14683), .Z(n14675) );
  XNOR U19087 ( .A(n14665), .B(n14667), .Z(n14683) );
  AND U19088 ( .A(n14684), .B(n14685), .Z(n14667) );
  NANDN U19089 ( .A(n14686), .B(n14687), .Z(n14685) );
  NANDN U19090 ( .A(n14688), .B(n14689), .Z(n14687) );
  IV U19091 ( .A(n14690), .Z(n14689) );
  NAND U19092 ( .A(n14690), .B(n14688), .Z(n14684) );
  AND U19093 ( .A(n14691), .B(n14692), .Z(n14665) );
  NAND U19094 ( .A(n14693), .B(n14694), .Z(n14692) );
  OR U19095 ( .A(n14695), .B(n14696), .Z(n14694) );
  NAND U19096 ( .A(n14696), .B(n14695), .Z(n14691) );
  IV U19097 ( .A(n14697), .Z(n14696) );
  NAND U19098 ( .A(n14698), .B(n14699), .Z(n14668) );
  NANDN U19099 ( .A(n14700), .B(n14701), .Z(n14699) );
  NAND U19100 ( .A(n14702), .B(n14703), .Z(n14701) );
  OR U19101 ( .A(n14703), .B(n14702), .Z(n14698) );
  IV U19102 ( .A(n14704), .Z(n14702) );
  AND U19103 ( .A(n14705), .B(n14706), .Z(n14671) );
  NAND U19104 ( .A(n14707), .B(n14708), .Z(n14706) );
  NANDN U19105 ( .A(n14709), .B(n14710), .Z(n14708) );
  NANDN U19106 ( .A(n14710), .B(n14709), .Z(n14705) );
  XOR U19107 ( .A(n14681), .B(n14711), .Z(n14673) );
  XNOR U19108 ( .A(n14678), .B(n14680), .Z(n14711) );
  AND U19109 ( .A(n14712), .B(n14713), .Z(n14680) );
  NANDN U19110 ( .A(n14714), .B(n14715), .Z(n14713) );
  NANDN U19111 ( .A(n14716), .B(n14717), .Z(n14715) );
  IV U19112 ( .A(n14718), .Z(n14717) );
  NAND U19113 ( .A(n14718), .B(n14716), .Z(n14712) );
  AND U19114 ( .A(n14719), .B(n14720), .Z(n14678) );
  NAND U19115 ( .A(n14721), .B(n14722), .Z(n14720) );
  OR U19116 ( .A(n14723), .B(n14724), .Z(n14722) );
  NAND U19117 ( .A(n14724), .B(n14723), .Z(n14719) );
  IV U19118 ( .A(n14725), .Z(n14724) );
  NAND U19119 ( .A(n14726), .B(n14727), .Z(n14681) );
  NANDN U19120 ( .A(n14728), .B(n14729), .Z(n14727) );
  NAND U19121 ( .A(n14730), .B(n14731), .Z(n14729) );
  OR U19122 ( .A(n14731), .B(n14730), .Z(n14726) );
  IV U19123 ( .A(n14732), .Z(n14730) );
  XOR U19124 ( .A(n14707), .B(n14733), .Z(N28938) );
  XNOR U19125 ( .A(n14710), .B(n14709), .Z(n14733) );
  XNOR U19126 ( .A(n14721), .B(n14734), .Z(n14709) );
  XOR U19127 ( .A(n14725), .B(n14723), .Z(n14734) );
  XOR U19128 ( .A(n14731), .B(n14735), .Z(n14723) );
  XOR U19129 ( .A(n14728), .B(n14732), .Z(n14735) );
  NAND U19130 ( .A(n14736), .B(n14737), .Z(n14732) );
  NAND U19131 ( .A(n14738), .B(n14739), .Z(n14737) );
  NAND U19132 ( .A(n14740), .B(n14741), .Z(n14736) );
  AND U19133 ( .A(n14742), .B(n14743), .Z(n14728) );
  NAND U19134 ( .A(n14744), .B(n14745), .Z(n14743) );
  NAND U19135 ( .A(n14746), .B(n14747), .Z(n14742) );
  NANDN U19136 ( .A(n14748), .B(n14749), .Z(n14731) );
  NANDN U19137 ( .A(n14750), .B(n14751), .Z(n14725) );
  XNOR U19138 ( .A(n14716), .B(n14752), .Z(n14721) );
  XOR U19139 ( .A(n14714), .B(n14718), .Z(n14752) );
  NAND U19140 ( .A(n14753), .B(n14754), .Z(n14718) );
  NAND U19141 ( .A(n14755), .B(n14756), .Z(n14754) );
  NAND U19142 ( .A(n14757), .B(n14758), .Z(n14753) );
  AND U19143 ( .A(n14759), .B(n14760), .Z(n14714) );
  NAND U19144 ( .A(n14761), .B(n14762), .Z(n14760) );
  NAND U19145 ( .A(n14763), .B(n14764), .Z(n14759) );
  AND U19146 ( .A(n14765), .B(n14766), .Z(n14716) );
  NAND U19147 ( .A(n14767), .B(n14768), .Z(n14710) );
  XNOR U19148 ( .A(n14693), .B(n14769), .Z(n14707) );
  XOR U19149 ( .A(n14697), .B(n14695), .Z(n14769) );
  XOR U19150 ( .A(n14703), .B(n14770), .Z(n14695) );
  XOR U19151 ( .A(n14700), .B(n14704), .Z(n14770) );
  NAND U19152 ( .A(n14771), .B(n14772), .Z(n14704) );
  NAND U19153 ( .A(n14773), .B(n14774), .Z(n14772) );
  NAND U19154 ( .A(n14775), .B(n14776), .Z(n14771) );
  AND U19155 ( .A(n14777), .B(n14778), .Z(n14700) );
  NAND U19156 ( .A(n14779), .B(n14780), .Z(n14778) );
  NAND U19157 ( .A(n14781), .B(n14782), .Z(n14777) );
  NANDN U19158 ( .A(n14783), .B(n14784), .Z(n14703) );
  NANDN U19159 ( .A(n14785), .B(n14786), .Z(n14697) );
  XNOR U19160 ( .A(n14688), .B(n14787), .Z(n14693) );
  XOR U19161 ( .A(n14686), .B(n14690), .Z(n14787) );
  NAND U19162 ( .A(n14788), .B(n14789), .Z(n14690) );
  NAND U19163 ( .A(n14790), .B(n14791), .Z(n14789) );
  NAND U19164 ( .A(n14792), .B(n14793), .Z(n14788) );
  AND U19165 ( .A(n14794), .B(n14795), .Z(n14686) );
  NAND U19166 ( .A(n14796), .B(n14797), .Z(n14795) );
  NAND U19167 ( .A(n14798), .B(n14799), .Z(n14794) );
  AND U19168 ( .A(n14800), .B(n14801), .Z(n14688) );
  XOR U19169 ( .A(n14768), .B(n14767), .Z(N28937) );
  XNOR U19170 ( .A(n14786), .B(n14785), .Z(n14767) );
  XNOR U19171 ( .A(n14800), .B(n14801), .Z(n14785) );
  XOR U19172 ( .A(n14797), .B(n14796), .Z(n14801) );
  XOR U19173 ( .A(y[2019]), .B(x[2019]), .Z(n14796) );
  XOR U19174 ( .A(n14799), .B(n14798), .Z(n14797) );
  XOR U19175 ( .A(y[2021]), .B(x[2021]), .Z(n14798) );
  XOR U19176 ( .A(y[2020]), .B(x[2020]), .Z(n14799) );
  XOR U19177 ( .A(n14791), .B(n14790), .Z(n14800) );
  XOR U19178 ( .A(n14793), .B(n14792), .Z(n14790) );
  XOR U19179 ( .A(y[2018]), .B(x[2018]), .Z(n14792) );
  XOR U19180 ( .A(y[2017]), .B(x[2017]), .Z(n14793) );
  XOR U19181 ( .A(y[2016]), .B(x[2016]), .Z(n14791) );
  XNOR U19182 ( .A(n14784), .B(n14783), .Z(n14786) );
  XNOR U19183 ( .A(n14780), .B(n14779), .Z(n14783) );
  XOR U19184 ( .A(n14782), .B(n14781), .Z(n14779) );
  XOR U19185 ( .A(y[2015]), .B(x[2015]), .Z(n14781) );
  XOR U19186 ( .A(y[2014]), .B(x[2014]), .Z(n14782) );
  XOR U19187 ( .A(y[2013]), .B(x[2013]), .Z(n14780) );
  XOR U19188 ( .A(n14774), .B(n14773), .Z(n14784) );
  XOR U19189 ( .A(n14776), .B(n14775), .Z(n14773) );
  XOR U19190 ( .A(y[2012]), .B(x[2012]), .Z(n14775) );
  XOR U19191 ( .A(y[2011]), .B(x[2011]), .Z(n14776) );
  XOR U19192 ( .A(y[2010]), .B(x[2010]), .Z(n14774) );
  XNOR U19193 ( .A(n14751), .B(n14750), .Z(n14768) );
  XNOR U19194 ( .A(n14765), .B(n14766), .Z(n14750) );
  XOR U19195 ( .A(n14762), .B(n14761), .Z(n14766) );
  XOR U19196 ( .A(y[2007]), .B(x[2007]), .Z(n14761) );
  XOR U19197 ( .A(n14764), .B(n14763), .Z(n14762) );
  XOR U19198 ( .A(y[2009]), .B(x[2009]), .Z(n14763) );
  XOR U19199 ( .A(y[2008]), .B(x[2008]), .Z(n14764) );
  XOR U19200 ( .A(n14756), .B(n14755), .Z(n14765) );
  XOR U19201 ( .A(n14758), .B(n14757), .Z(n14755) );
  XOR U19202 ( .A(y[2006]), .B(x[2006]), .Z(n14757) );
  XOR U19203 ( .A(y[2005]), .B(x[2005]), .Z(n14758) );
  XOR U19204 ( .A(y[2004]), .B(x[2004]), .Z(n14756) );
  XNOR U19205 ( .A(n14749), .B(n14748), .Z(n14751) );
  XNOR U19206 ( .A(n14745), .B(n14744), .Z(n14748) );
  XOR U19207 ( .A(n14747), .B(n14746), .Z(n14744) );
  XOR U19208 ( .A(y[2003]), .B(x[2003]), .Z(n14746) );
  XOR U19209 ( .A(y[2002]), .B(x[2002]), .Z(n14747) );
  XOR U19210 ( .A(y[2001]), .B(x[2001]), .Z(n14745) );
  XOR U19211 ( .A(n14739), .B(n14738), .Z(n14749) );
  XOR U19212 ( .A(n14741), .B(n14740), .Z(n14738) );
  XOR U19213 ( .A(y[2000]), .B(x[2000]), .Z(n14740) );
  XOR U19214 ( .A(y[1999]), .B(x[1999]), .Z(n14741) );
  XOR U19215 ( .A(y[1998]), .B(x[1998]), .Z(n14739) );
  NAND U19216 ( .A(n14802), .B(n14803), .Z(N28929) );
  NAND U19217 ( .A(n14804), .B(n14805), .Z(n14803) );
  NANDN U19218 ( .A(n14806), .B(n14807), .Z(n14805) );
  NANDN U19219 ( .A(n14807), .B(n14806), .Z(n14802) );
  XOR U19220 ( .A(n14806), .B(n14808), .Z(N28928) );
  XNOR U19221 ( .A(n14804), .B(n14807), .Z(n14808) );
  NAND U19222 ( .A(n14809), .B(n14810), .Z(n14807) );
  NAND U19223 ( .A(n14811), .B(n14812), .Z(n14810) );
  NANDN U19224 ( .A(n14813), .B(n14814), .Z(n14812) );
  NANDN U19225 ( .A(n14814), .B(n14813), .Z(n14809) );
  AND U19226 ( .A(n14815), .B(n14816), .Z(n14804) );
  NAND U19227 ( .A(n14817), .B(n14818), .Z(n14816) );
  OR U19228 ( .A(n14819), .B(n14820), .Z(n14818) );
  NAND U19229 ( .A(n14820), .B(n14819), .Z(n14815) );
  IV U19230 ( .A(n14821), .Z(n14820) );
  AND U19231 ( .A(n14822), .B(n14823), .Z(n14806) );
  NAND U19232 ( .A(n14824), .B(n14825), .Z(n14823) );
  NANDN U19233 ( .A(n14826), .B(n14827), .Z(n14825) );
  NANDN U19234 ( .A(n14827), .B(n14826), .Z(n14822) );
  XOR U19235 ( .A(n14819), .B(n14828), .Z(N28927) );
  XOR U19236 ( .A(n14817), .B(n14821), .Z(n14828) );
  XNOR U19237 ( .A(n14814), .B(n14829), .Z(n14821) );
  XNOR U19238 ( .A(n14811), .B(n14813), .Z(n14829) );
  AND U19239 ( .A(n14830), .B(n14831), .Z(n14813) );
  NANDN U19240 ( .A(n14832), .B(n14833), .Z(n14831) );
  NANDN U19241 ( .A(n14834), .B(n14835), .Z(n14833) );
  IV U19242 ( .A(n14836), .Z(n14835) );
  NAND U19243 ( .A(n14836), .B(n14834), .Z(n14830) );
  AND U19244 ( .A(n14837), .B(n14838), .Z(n14811) );
  NAND U19245 ( .A(n14839), .B(n14840), .Z(n14838) );
  OR U19246 ( .A(n14841), .B(n14842), .Z(n14840) );
  NAND U19247 ( .A(n14842), .B(n14841), .Z(n14837) );
  IV U19248 ( .A(n14843), .Z(n14842) );
  NAND U19249 ( .A(n14844), .B(n14845), .Z(n14814) );
  NANDN U19250 ( .A(n14846), .B(n14847), .Z(n14845) );
  NAND U19251 ( .A(n14848), .B(n14849), .Z(n14847) );
  OR U19252 ( .A(n14849), .B(n14848), .Z(n14844) );
  IV U19253 ( .A(n14850), .Z(n14848) );
  AND U19254 ( .A(n14851), .B(n14852), .Z(n14817) );
  NAND U19255 ( .A(n14853), .B(n14854), .Z(n14852) );
  NANDN U19256 ( .A(n14855), .B(n14856), .Z(n14854) );
  NANDN U19257 ( .A(n14856), .B(n14855), .Z(n14851) );
  XOR U19258 ( .A(n14827), .B(n14857), .Z(n14819) );
  XNOR U19259 ( .A(n14824), .B(n14826), .Z(n14857) );
  AND U19260 ( .A(n14858), .B(n14859), .Z(n14826) );
  NANDN U19261 ( .A(n14860), .B(n14861), .Z(n14859) );
  NANDN U19262 ( .A(n14862), .B(n14863), .Z(n14861) );
  IV U19263 ( .A(n14864), .Z(n14863) );
  NAND U19264 ( .A(n14864), .B(n14862), .Z(n14858) );
  AND U19265 ( .A(n14865), .B(n14866), .Z(n14824) );
  NAND U19266 ( .A(n14867), .B(n14868), .Z(n14866) );
  OR U19267 ( .A(n14869), .B(n14870), .Z(n14868) );
  NAND U19268 ( .A(n14870), .B(n14869), .Z(n14865) );
  IV U19269 ( .A(n14871), .Z(n14870) );
  NAND U19270 ( .A(n14872), .B(n14873), .Z(n14827) );
  NANDN U19271 ( .A(n14874), .B(n14875), .Z(n14873) );
  NAND U19272 ( .A(n14876), .B(n14877), .Z(n14875) );
  OR U19273 ( .A(n14877), .B(n14876), .Z(n14872) );
  IV U19274 ( .A(n14878), .Z(n14876) );
  XOR U19275 ( .A(n14853), .B(n14879), .Z(N28926) );
  XNOR U19276 ( .A(n14856), .B(n14855), .Z(n14879) );
  XNOR U19277 ( .A(n14867), .B(n14880), .Z(n14855) );
  XOR U19278 ( .A(n14871), .B(n14869), .Z(n14880) );
  XOR U19279 ( .A(n14877), .B(n14881), .Z(n14869) );
  XOR U19280 ( .A(n14874), .B(n14878), .Z(n14881) );
  NAND U19281 ( .A(n14882), .B(n14883), .Z(n14878) );
  NAND U19282 ( .A(n14884), .B(n14885), .Z(n14883) );
  NAND U19283 ( .A(n14886), .B(n14887), .Z(n14882) );
  AND U19284 ( .A(n14888), .B(n14889), .Z(n14874) );
  NAND U19285 ( .A(n14890), .B(n14891), .Z(n14889) );
  NAND U19286 ( .A(n14892), .B(n14893), .Z(n14888) );
  NANDN U19287 ( .A(n14894), .B(n14895), .Z(n14877) );
  NANDN U19288 ( .A(n14896), .B(n14897), .Z(n14871) );
  XNOR U19289 ( .A(n14862), .B(n14898), .Z(n14867) );
  XOR U19290 ( .A(n14860), .B(n14864), .Z(n14898) );
  NAND U19291 ( .A(n14899), .B(n14900), .Z(n14864) );
  NAND U19292 ( .A(n14901), .B(n14902), .Z(n14900) );
  NAND U19293 ( .A(n14903), .B(n14904), .Z(n14899) );
  AND U19294 ( .A(n14905), .B(n14906), .Z(n14860) );
  NAND U19295 ( .A(n14907), .B(n14908), .Z(n14906) );
  NAND U19296 ( .A(n14909), .B(n14910), .Z(n14905) );
  AND U19297 ( .A(n14911), .B(n14912), .Z(n14862) );
  NAND U19298 ( .A(n14913), .B(n14914), .Z(n14856) );
  XNOR U19299 ( .A(n14839), .B(n14915), .Z(n14853) );
  XOR U19300 ( .A(n14843), .B(n14841), .Z(n14915) );
  XOR U19301 ( .A(n14849), .B(n14916), .Z(n14841) );
  XOR U19302 ( .A(n14846), .B(n14850), .Z(n14916) );
  NAND U19303 ( .A(n14917), .B(n14918), .Z(n14850) );
  NAND U19304 ( .A(n14919), .B(n14920), .Z(n14918) );
  NAND U19305 ( .A(n14921), .B(n14922), .Z(n14917) );
  AND U19306 ( .A(n14923), .B(n14924), .Z(n14846) );
  NAND U19307 ( .A(n14925), .B(n14926), .Z(n14924) );
  NAND U19308 ( .A(n14927), .B(n14928), .Z(n14923) );
  NANDN U19309 ( .A(n14929), .B(n14930), .Z(n14849) );
  NANDN U19310 ( .A(n14931), .B(n14932), .Z(n14843) );
  XNOR U19311 ( .A(n14834), .B(n14933), .Z(n14839) );
  XOR U19312 ( .A(n14832), .B(n14836), .Z(n14933) );
  NAND U19313 ( .A(n14934), .B(n14935), .Z(n14836) );
  NAND U19314 ( .A(n14936), .B(n14937), .Z(n14935) );
  NAND U19315 ( .A(n14938), .B(n14939), .Z(n14934) );
  AND U19316 ( .A(n14940), .B(n14941), .Z(n14832) );
  NAND U19317 ( .A(n14942), .B(n14943), .Z(n14941) );
  NAND U19318 ( .A(n14944), .B(n14945), .Z(n14940) );
  AND U19319 ( .A(n14946), .B(n14947), .Z(n14834) );
  XOR U19320 ( .A(n14914), .B(n14913), .Z(N28925) );
  XNOR U19321 ( .A(n14932), .B(n14931), .Z(n14913) );
  XNOR U19322 ( .A(n14946), .B(n14947), .Z(n14931) );
  XOR U19323 ( .A(n14943), .B(n14942), .Z(n14947) );
  XOR U19324 ( .A(y[1995]), .B(x[1995]), .Z(n14942) );
  XOR U19325 ( .A(n14945), .B(n14944), .Z(n14943) );
  XOR U19326 ( .A(y[1997]), .B(x[1997]), .Z(n14944) );
  XOR U19327 ( .A(y[1996]), .B(x[1996]), .Z(n14945) );
  XOR U19328 ( .A(n14937), .B(n14936), .Z(n14946) );
  XOR U19329 ( .A(n14939), .B(n14938), .Z(n14936) );
  XOR U19330 ( .A(y[1994]), .B(x[1994]), .Z(n14938) );
  XOR U19331 ( .A(y[1993]), .B(x[1993]), .Z(n14939) );
  XOR U19332 ( .A(y[1992]), .B(x[1992]), .Z(n14937) );
  XNOR U19333 ( .A(n14930), .B(n14929), .Z(n14932) );
  XNOR U19334 ( .A(n14926), .B(n14925), .Z(n14929) );
  XOR U19335 ( .A(n14928), .B(n14927), .Z(n14925) );
  XOR U19336 ( .A(y[1991]), .B(x[1991]), .Z(n14927) );
  XOR U19337 ( .A(y[1990]), .B(x[1990]), .Z(n14928) );
  XOR U19338 ( .A(y[1989]), .B(x[1989]), .Z(n14926) );
  XOR U19339 ( .A(n14920), .B(n14919), .Z(n14930) );
  XOR U19340 ( .A(n14922), .B(n14921), .Z(n14919) );
  XOR U19341 ( .A(y[1988]), .B(x[1988]), .Z(n14921) );
  XOR U19342 ( .A(y[1987]), .B(x[1987]), .Z(n14922) );
  XOR U19343 ( .A(y[1986]), .B(x[1986]), .Z(n14920) );
  XNOR U19344 ( .A(n14897), .B(n14896), .Z(n14914) );
  XNOR U19345 ( .A(n14911), .B(n14912), .Z(n14896) );
  XOR U19346 ( .A(n14908), .B(n14907), .Z(n14912) );
  XOR U19347 ( .A(y[1983]), .B(x[1983]), .Z(n14907) );
  XOR U19348 ( .A(n14910), .B(n14909), .Z(n14908) );
  XOR U19349 ( .A(y[1985]), .B(x[1985]), .Z(n14909) );
  XOR U19350 ( .A(y[1984]), .B(x[1984]), .Z(n14910) );
  XOR U19351 ( .A(n14902), .B(n14901), .Z(n14911) );
  XOR U19352 ( .A(n14904), .B(n14903), .Z(n14901) );
  XOR U19353 ( .A(y[1982]), .B(x[1982]), .Z(n14903) );
  XOR U19354 ( .A(y[1981]), .B(x[1981]), .Z(n14904) );
  XOR U19355 ( .A(y[1980]), .B(x[1980]), .Z(n14902) );
  XNOR U19356 ( .A(n14895), .B(n14894), .Z(n14897) );
  XNOR U19357 ( .A(n14891), .B(n14890), .Z(n14894) );
  XOR U19358 ( .A(n14893), .B(n14892), .Z(n14890) );
  XOR U19359 ( .A(y[1979]), .B(x[1979]), .Z(n14892) );
  XOR U19360 ( .A(y[1978]), .B(x[1978]), .Z(n14893) );
  XOR U19361 ( .A(y[1977]), .B(x[1977]), .Z(n14891) );
  XOR U19362 ( .A(n14885), .B(n14884), .Z(n14895) );
  XOR U19363 ( .A(n14887), .B(n14886), .Z(n14884) );
  XOR U19364 ( .A(y[1976]), .B(x[1976]), .Z(n14886) );
  XOR U19365 ( .A(y[1975]), .B(x[1975]), .Z(n14887) );
  XOR U19366 ( .A(y[1974]), .B(x[1974]), .Z(n14885) );
  NAND U19367 ( .A(n14948), .B(n14949), .Z(N28917) );
  NAND U19368 ( .A(n14950), .B(n14951), .Z(n14949) );
  NANDN U19369 ( .A(n14952), .B(n14953), .Z(n14951) );
  NANDN U19370 ( .A(n14953), .B(n14952), .Z(n14948) );
  XOR U19371 ( .A(n14952), .B(n14954), .Z(N28916) );
  XNOR U19372 ( .A(n14950), .B(n14953), .Z(n14954) );
  NAND U19373 ( .A(n14955), .B(n14956), .Z(n14953) );
  NAND U19374 ( .A(n14957), .B(n14958), .Z(n14956) );
  NANDN U19375 ( .A(n14959), .B(n14960), .Z(n14958) );
  NANDN U19376 ( .A(n14960), .B(n14959), .Z(n14955) );
  AND U19377 ( .A(n14961), .B(n14962), .Z(n14950) );
  NAND U19378 ( .A(n14963), .B(n14964), .Z(n14962) );
  OR U19379 ( .A(n14965), .B(n14966), .Z(n14964) );
  NAND U19380 ( .A(n14966), .B(n14965), .Z(n14961) );
  IV U19381 ( .A(n14967), .Z(n14966) );
  AND U19382 ( .A(n14968), .B(n14969), .Z(n14952) );
  NAND U19383 ( .A(n14970), .B(n14971), .Z(n14969) );
  NANDN U19384 ( .A(n14972), .B(n14973), .Z(n14971) );
  NANDN U19385 ( .A(n14973), .B(n14972), .Z(n14968) );
  XOR U19386 ( .A(n14965), .B(n14974), .Z(N28915) );
  XOR U19387 ( .A(n14963), .B(n14967), .Z(n14974) );
  XNOR U19388 ( .A(n14960), .B(n14975), .Z(n14967) );
  XNOR U19389 ( .A(n14957), .B(n14959), .Z(n14975) );
  AND U19390 ( .A(n14976), .B(n14977), .Z(n14959) );
  NANDN U19391 ( .A(n14978), .B(n14979), .Z(n14977) );
  NANDN U19392 ( .A(n14980), .B(n14981), .Z(n14979) );
  IV U19393 ( .A(n14982), .Z(n14981) );
  NAND U19394 ( .A(n14982), .B(n14980), .Z(n14976) );
  AND U19395 ( .A(n14983), .B(n14984), .Z(n14957) );
  NAND U19396 ( .A(n14985), .B(n14986), .Z(n14984) );
  OR U19397 ( .A(n14987), .B(n14988), .Z(n14986) );
  NAND U19398 ( .A(n14988), .B(n14987), .Z(n14983) );
  IV U19399 ( .A(n14989), .Z(n14988) );
  NAND U19400 ( .A(n14990), .B(n14991), .Z(n14960) );
  NANDN U19401 ( .A(n14992), .B(n14993), .Z(n14991) );
  NAND U19402 ( .A(n14994), .B(n14995), .Z(n14993) );
  OR U19403 ( .A(n14995), .B(n14994), .Z(n14990) );
  IV U19404 ( .A(n14996), .Z(n14994) );
  AND U19405 ( .A(n14997), .B(n14998), .Z(n14963) );
  NAND U19406 ( .A(n14999), .B(n15000), .Z(n14998) );
  NANDN U19407 ( .A(n15001), .B(n15002), .Z(n15000) );
  NANDN U19408 ( .A(n15002), .B(n15001), .Z(n14997) );
  XOR U19409 ( .A(n14973), .B(n15003), .Z(n14965) );
  XNOR U19410 ( .A(n14970), .B(n14972), .Z(n15003) );
  AND U19411 ( .A(n15004), .B(n15005), .Z(n14972) );
  NANDN U19412 ( .A(n15006), .B(n15007), .Z(n15005) );
  NANDN U19413 ( .A(n15008), .B(n15009), .Z(n15007) );
  IV U19414 ( .A(n15010), .Z(n15009) );
  NAND U19415 ( .A(n15010), .B(n15008), .Z(n15004) );
  AND U19416 ( .A(n15011), .B(n15012), .Z(n14970) );
  NAND U19417 ( .A(n15013), .B(n15014), .Z(n15012) );
  OR U19418 ( .A(n15015), .B(n15016), .Z(n15014) );
  NAND U19419 ( .A(n15016), .B(n15015), .Z(n15011) );
  IV U19420 ( .A(n15017), .Z(n15016) );
  NAND U19421 ( .A(n15018), .B(n15019), .Z(n14973) );
  NANDN U19422 ( .A(n15020), .B(n15021), .Z(n15019) );
  NAND U19423 ( .A(n15022), .B(n15023), .Z(n15021) );
  OR U19424 ( .A(n15023), .B(n15022), .Z(n15018) );
  IV U19425 ( .A(n15024), .Z(n15022) );
  XOR U19426 ( .A(n14999), .B(n15025), .Z(N28914) );
  XNOR U19427 ( .A(n15002), .B(n15001), .Z(n15025) );
  XNOR U19428 ( .A(n15013), .B(n15026), .Z(n15001) );
  XOR U19429 ( .A(n15017), .B(n15015), .Z(n15026) );
  XOR U19430 ( .A(n15023), .B(n15027), .Z(n15015) );
  XOR U19431 ( .A(n15020), .B(n15024), .Z(n15027) );
  NAND U19432 ( .A(n15028), .B(n15029), .Z(n15024) );
  NAND U19433 ( .A(n15030), .B(n15031), .Z(n15029) );
  NAND U19434 ( .A(n15032), .B(n15033), .Z(n15028) );
  AND U19435 ( .A(n15034), .B(n15035), .Z(n15020) );
  NAND U19436 ( .A(n15036), .B(n15037), .Z(n15035) );
  NAND U19437 ( .A(n15038), .B(n15039), .Z(n15034) );
  NANDN U19438 ( .A(n15040), .B(n15041), .Z(n15023) );
  NANDN U19439 ( .A(n15042), .B(n15043), .Z(n15017) );
  XNOR U19440 ( .A(n15008), .B(n15044), .Z(n15013) );
  XOR U19441 ( .A(n15006), .B(n15010), .Z(n15044) );
  NAND U19442 ( .A(n15045), .B(n15046), .Z(n15010) );
  NAND U19443 ( .A(n15047), .B(n15048), .Z(n15046) );
  NAND U19444 ( .A(n15049), .B(n15050), .Z(n15045) );
  AND U19445 ( .A(n15051), .B(n15052), .Z(n15006) );
  NAND U19446 ( .A(n15053), .B(n15054), .Z(n15052) );
  NAND U19447 ( .A(n15055), .B(n15056), .Z(n15051) );
  AND U19448 ( .A(n15057), .B(n15058), .Z(n15008) );
  NAND U19449 ( .A(n15059), .B(n15060), .Z(n15002) );
  XNOR U19450 ( .A(n14985), .B(n15061), .Z(n14999) );
  XOR U19451 ( .A(n14989), .B(n14987), .Z(n15061) );
  XOR U19452 ( .A(n14995), .B(n15062), .Z(n14987) );
  XOR U19453 ( .A(n14992), .B(n14996), .Z(n15062) );
  NAND U19454 ( .A(n15063), .B(n15064), .Z(n14996) );
  NAND U19455 ( .A(n15065), .B(n15066), .Z(n15064) );
  NAND U19456 ( .A(n15067), .B(n15068), .Z(n15063) );
  AND U19457 ( .A(n15069), .B(n15070), .Z(n14992) );
  NAND U19458 ( .A(n15071), .B(n15072), .Z(n15070) );
  NAND U19459 ( .A(n15073), .B(n15074), .Z(n15069) );
  NANDN U19460 ( .A(n15075), .B(n15076), .Z(n14995) );
  NANDN U19461 ( .A(n15077), .B(n15078), .Z(n14989) );
  XNOR U19462 ( .A(n14980), .B(n15079), .Z(n14985) );
  XOR U19463 ( .A(n14978), .B(n14982), .Z(n15079) );
  NAND U19464 ( .A(n15080), .B(n15081), .Z(n14982) );
  NAND U19465 ( .A(n15082), .B(n15083), .Z(n15081) );
  NAND U19466 ( .A(n15084), .B(n15085), .Z(n15080) );
  AND U19467 ( .A(n15086), .B(n15087), .Z(n14978) );
  NAND U19468 ( .A(n15088), .B(n15089), .Z(n15087) );
  NAND U19469 ( .A(n15090), .B(n15091), .Z(n15086) );
  AND U19470 ( .A(n15092), .B(n15093), .Z(n14980) );
  XOR U19471 ( .A(n15060), .B(n15059), .Z(N28913) );
  XNOR U19472 ( .A(n15078), .B(n15077), .Z(n15059) );
  XNOR U19473 ( .A(n15092), .B(n15093), .Z(n15077) );
  XOR U19474 ( .A(n15089), .B(n15088), .Z(n15093) );
  XOR U19475 ( .A(y[1971]), .B(x[1971]), .Z(n15088) );
  XOR U19476 ( .A(n15091), .B(n15090), .Z(n15089) );
  XOR U19477 ( .A(y[1973]), .B(x[1973]), .Z(n15090) );
  XOR U19478 ( .A(y[1972]), .B(x[1972]), .Z(n15091) );
  XOR U19479 ( .A(n15083), .B(n15082), .Z(n15092) );
  XOR U19480 ( .A(n15085), .B(n15084), .Z(n15082) );
  XOR U19481 ( .A(y[1970]), .B(x[1970]), .Z(n15084) );
  XOR U19482 ( .A(y[1969]), .B(x[1969]), .Z(n15085) );
  XOR U19483 ( .A(y[1968]), .B(x[1968]), .Z(n15083) );
  XNOR U19484 ( .A(n15076), .B(n15075), .Z(n15078) );
  XNOR U19485 ( .A(n15072), .B(n15071), .Z(n15075) );
  XOR U19486 ( .A(n15074), .B(n15073), .Z(n15071) );
  XOR U19487 ( .A(y[1967]), .B(x[1967]), .Z(n15073) );
  XOR U19488 ( .A(y[1966]), .B(x[1966]), .Z(n15074) );
  XOR U19489 ( .A(y[1965]), .B(x[1965]), .Z(n15072) );
  XOR U19490 ( .A(n15066), .B(n15065), .Z(n15076) );
  XOR U19491 ( .A(n15068), .B(n15067), .Z(n15065) );
  XOR U19492 ( .A(y[1964]), .B(x[1964]), .Z(n15067) );
  XOR U19493 ( .A(y[1963]), .B(x[1963]), .Z(n15068) );
  XOR U19494 ( .A(y[1962]), .B(x[1962]), .Z(n15066) );
  XNOR U19495 ( .A(n15043), .B(n15042), .Z(n15060) );
  XNOR U19496 ( .A(n15057), .B(n15058), .Z(n15042) );
  XOR U19497 ( .A(n15054), .B(n15053), .Z(n15058) );
  XOR U19498 ( .A(y[1959]), .B(x[1959]), .Z(n15053) );
  XOR U19499 ( .A(n15056), .B(n15055), .Z(n15054) );
  XOR U19500 ( .A(y[1961]), .B(x[1961]), .Z(n15055) );
  XOR U19501 ( .A(y[1960]), .B(x[1960]), .Z(n15056) );
  XOR U19502 ( .A(n15048), .B(n15047), .Z(n15057) );
  XOR U19503 ( .A(n15050), .B(n15049), .Z(n15047) );
  XOR U19504 ( .A(y[1958]), .B(x[1958]), .Z(n15049) );
  XOR U19505 ( .A(y[1957]), .B(x[1957]), .Z(n15050) );
  XOR U19506 ( .A(y[1956]), .B(x[1956]), .Z(n15048) );
  XNOR U19507 ( .A(n15041), .B(n15040), .Z(n15043) );
  XNOR U19508 ( .A(n15037), .B(n15036), .Z(n15040) );
  XOR U19509 ( .A(n15039), .B(n15038), .Z(n15036) );
  XOR U19510 ( .A(y[1955]), .B(x[1955]), .Z(n15038) );
  XOR U19511 ( .A(y[1954]), .B(x[1954]), .Z(n15039) );
  XOR U19512 ( .A(y[1953]), .B(x[1953]), .Z(n15037) );
  XOR U19513 ( .A(n15031), .B(n15030), .Z(n15041) );
  XOR U19514 ( .A(n15033), .B(n15032), .Z(n15030) );
  XOR U19515 ( .A(y[1952]), .B(x[1952]), .Z(n15032) );
  XOR U19516 ( .A(y[1951]), .B(x[1951]), .Z(n15033) );
  XOR U19517 ( .A(y[1950]), .B(x[1950]), .Z(n15031) );
  NAND U19518 ( .A(n15094), .B(n15095), .Z(N28905) );
  NAND U19519 ( .A(n15096), .B(n15097), .Z(n15095) );
  NANDN U19520 ( .A(n15098), .B(n15099), .Z(n15097) );
  NANDN U19521 ( .A(n15099), .B(n15098), .Z(n15094) );
  XOR U19522 ( .A(n15098), .B(n15100), .Z(N28904) );
  XNOR U19523 ( .A(n15096), .B(n15099), .Z(n15100) );
  NAND U19524 ( .A(n15101), .B(n15102), .Z(n15099) );
  NAND U19525 ( .A(n15103), .B(n15104), .Z(n15102) );
  NANDN U19526 ( .A(n15105), .B(n15106), .Z(n15104) );
  NANDN U19527 ( .A(n15106), .B(n15105), .Z(n15101) );
  AND U19528 ( .A(n15107), .B(n15108), .Z(n15096) );
  NAND U19529 ( .A(n15109), .B(n15110), .Z(n15108) );
  OR U19530 ( .A(n15111), .B(n15112), .Z(n15110) );
  NAND U19531 ( .A(n15112), .B(n15111), .Z(n15107) );
  IV U19532 ( .A(n15113), .Z(n15112) );
  AND U19533 ( .A(n15114), .B(n15115), .Z(n15098) );
  NAND U19534 ( .A(n15116), .B(n15117), .Z(n15115) );
  NANDN U19535 ( .A(n15118), .B(n15119), .Z(n15117) );
  NANDN U19536 ( .A(n15119), .B(n15118), .Z(n15114) );
  XOR U19537 ( .A(n15111), .B(n15120), .Z(N28903) );
  XOR U19538 ( .A(n15109), .B(n15113), .Z(n15120) );
  XNOR U19539 ( .A(n15106), .B(n15121), .Z(n15113) );
  XNOR U19540 ( .A(n15103), .B(n15105), .Z(n15121) );
  AND U19541 ( .A(n15122), .B(n15123), .Z(n15105) );
  NANDN U19542 ( .A(n15124), .B(n15125), .Z(n15123) );
  NANDN U19543 ( .A(n15126), .B(n15127), .Z(n15125) );
  IV U19544 ( .A(n15128), .Z(n15127) );
  NAND U19545 ( .A(n15128), .B(n15126), .Z(n15122) );
  AND U19546 ( .A(n15129), .B(n15130), .Z(n15103) );
  NAND U19547 ( .A(n15131), .B(n15132), .Z(n15130) );
  OR U19548 ( .A(n15133), .B(n15134), .Z(n15132) );
  NAND U19549 ( .A(n15134), .B(n15133), .Z(n15129) );
  IV U19550 ( .A(n15135), .Z(n15134) );
  NAND U19551 ( .A(n15136), .B(n15137), .Z(n15106) );
  NANDN U19552 ( .A(n15138), .B(n15139), .Z(n15137) );
  NAND U19553 ( .A(n15140), .B(n15141), .Z(n15139) );
  OR U19554 ( .A(n15141), .B(n15140), .Z(n15136) );
  IV U19555 ( .A(n15142), .Z(n15140) );
  AND U19556 ( .A(n15143), .B(n15144), .Z(n15109) );
  NAND U19557 ( .A(n15145), .B(n15146), .Z(n15144) );
  NANDN U19558 ( .A(n15147), .B(n15148), .Z(n15146) );
  NANDN U19559 ( .A(n15148), .B(n15147), .Z(n15143) );
  XOR U19560 ( .A(n15119), .B(n15149), .Z(n15111) );
  XNOR U19561 ( .A(n15116), .B(n15118), .Z(n15149) );
  AND U19562 ( .A(n15150), .B(n15151), .Z(n15118) );
  NANDN U19563 ( .A(n15152), .B(n15153), .Z(n15151) );
  NANDN U19564 ( .A(n15154), .B(n15155), .Z(n15153) );
  IV U19565 ( .A(n15156), .Z(n15155) );
  NAND U19566 ( .A(n15156), .B(n15154), .Z(n15150) );
  AND U19567 ( .A(n15157), .B(n15158), .Z(n15116) );
  NAND U19568 ( .A(n15159), .B(n15160), .Z(n15158) );
  OR U19569 ( .A(n15161), .B(n15162), .Z(n15160) );
  NAND U19570 ( .A(n15162), .B(n15161), .Z(n15157) );
  IV U19571 ( .A(n15163), .Z(n15162) );
  NAND U19572 ( .A(n15164), .B(n15165), .Z(n15119) );
  NANDN U19573 ( .A(n15166), .B(n15167), .Z(n15165) );
  NAND U19574 ( .A(n15168), .B(n15169), .Z(n15167) );
  OR U19575 ( .A(n15169), .B(n15168), .Z(n15164) );
  IV U19576 ( .A(n15170), .Z(n15168) );
  XOR U19577 ( .A(n15145), .B(n15171), .Z(N28902) );
  XNOR U19578 ( .A(n15148), .B(n15147), .Z(n15171) );
  XNOR U19579 ( .A(n15159), .B(n15172), .Z(n15147) );
  XOR U19580 ( .A(n15163), .B(n15161), .Z(n15172) );
  XOR U19581 ( .A(n15169), .B(n15173), .Z(n15161) );
  XOR U19582 ( .A(n15166), .B(n15170), .Z(n15173) );
  NAND U19583 ( .A(n15174), .B(n15175), .Z(n15170) );
  NAND U19584 ( .A(n15176), .B(n15177), .Z(n15175) );
  NAND U19585 ( .A(n15178), .B(n15179), .Z(n15174) );
  AND U19586 ( .A(n15180), .B(n15181), .Z(n15166) );
  NAND U19587 ( .A(n15182), .B(n15183), .Z(n15181) );
  NAND U19588 ( .A(n15184), .B(n15185), .Z(n15180) );
  NANDN U19589 ( .A(n15186), .B(n15187), .Z(n15169) );
  NANDN U19590 ( .A(n15188), .B(n15189), .Z(n15163) );
  XNOR U19591 ( .A(n15154), .B(n15190), .Z(n15159) );
  XOR U19592 ( .A(n15152), .B(n15156), .Z(n15190) );
  NAND U19593 ( .A(n15191), .B(n15192), .Z(n15156) );
  NAND U19594 ( .A(n15193), .B(n15194), .Z(n15192) );
  NAND U19595 ( .A(n15195), .B(n15196), .Z(n15191) );
  AND U19596 ( .A(n15197), .B(n15198), .Z(n15152) );
  NAND U19597 ( .A(n15199), .B(n15200), .Z(n15198) );
  NAND U19598 ( .A(n15201), .B(n15202), .Z(n15197) );
  AND U19599 ( .A(n15203), .B(n15204), .Z(n15154) );
  NAND U19600 ( .A(n15205), .B(n15206), .Z(n15148) );
  XNOR U19601 ( .A(n15131), .B(n15207), .Z(n15145) );
  XOR U19602 ( .A(n15135), .B(n15133), .Z(n15207) );
  XOR U19603 ( .A(n15141), .B(n15208), .Z(n15133) );
  XOR U19604 ( .A(n15138), .B(n15142), .Z(n15208) );
  NAND U19605 ( .A(n15209), .B(n15210), .Z(n15142) );
  NAND U19606 ( .A(n15211), .B(n15212), .Z(n15210) );
  NAND U19607 ( .A(n15213), .B(n15214), .Z(n15209) );
  AND U19608 ( .A(n15215), .B(n15216), .Z(n15138) );
  NAND U19609 ( .A(n15217), .B(n15218), .Z(n15216) );
  NAND U19610 ( .A(n15219), .B(n15220), .Z(n15215) );
  NANDN U19611 ( .A(n15221), .B(n15222), .Z(n15141) );
  NANDN U19612 ( .A(n15223), .B(n15224), .Z(n15135) );
  XNOR U19613 ( .A(n15126), .B(n15225), .Z(n15131) );
  XOR U19614 ( .A(n15124), .B(n15128), .Z(n15225) );
  NAND U19615 ( .A(n15226), .B(n15227), .Z(n15128) );
  NAND U19616 ( .A(n15228), .B(n15229), .Z(n15227) );
  NAND U19617 ( .A(n15230), .B(n15231), .Z(n15226) );
  AND U19618 ( .A(n15232), .B(n15233), .Z(n15124) );
  NAND U19619 ( .A(n15234), .B(n15235), .Z(n15233) );
  NAND U19620 ( .A(n15236), .B(n15237), .Z(n15232) );
  AND U19621 ( .A(n15238), .B(n15239), .Z(n15126) );
  XOR U19622 ( .A(n15206), .B(n15205), .Z(N28901) );
  XNOR U19623 ( .A(n15224), .B(n15223), .Z(n15205) );
  XNOR U19624 ( .A(n15238), .B(n15239), .Z(n15223) );
  XOR U19625 ( .A(n15235), .B(n15234), .Z(n15239) );
  XOR U19626 ( .A(y[1947]), .B(x[1947]), .Z(n15234) );
  XOR U19627 ( .A(n15237), .B(n15236), .Z(n15235) );
  XOR U19628 ( .A(y[1949]), .B(x[1949]), .Z(n15236) );
  XOR U19629 ( .A(y[1948]), .B(x[1948]), .Z(n15237) );
  XOR U19630 ( .A(n15229), .B(n15228), .Z(n15238) );
  XOR U19631 ( .A(n15231), .B(n15230), .Z(n15228) );
  XOR U19632 ( .A(y[1946]), .B(x[1946]), .Z(n15230) );
  XOR U19633 ( .A(y[1945]), .B(x[1945]), .Z(n15231) );
  XOR U19634 ( .A(y[1944]), .B(x[1944]), .Z(n15229) );
  XNOR U19635 ( .A(n15222), .B(n15221), .Z(n15224) );
  XNOR U19636 ( .A(n15218), .B(n15217), .Z(n15221) );
  XOR U19637 ( .A(n15220), .B(n15219), .Z(n15217) );
  XOR U19638 ( .A(y[1943]), .B(x[1943]), .Z(n15219) );
  XOR U19639 ( .A(y[1942]), .B(x[1942]), .Z(n15220) );
  XOR U19640 ( .A(y[1941]), .B(x[1941]), .Z(n15218) );
  XOR U19641 ( .A(n15212), .B(n15211), .Z(n15222) );
  XOR U19642 ( .A(n15214), .B(n15213), .Z(n15211) );
  XOR U19643 ( .A(y[1940]), .B(x[1940]), .Z(n15213) );
  XOR U19644 ( .A(y[1939]), .B(x[1939]), .Z(n15214) );
  XOR U19645 ( .A(y[1938]), .B(x[1938]), .Z(n15212) );
  XNOR U19646 ( .A(n15189), .B(n15188), .Z(n15206) );
  XNOR U19647 ( .A(n15203), .B(n15204), .Z(n15188) );
  XOR U19648 ( .A(n15200), .B(n15199), .Z(n15204) );
  XOR U19649 ( .A(y[1935]), .B(x[1935]), .Z(n15199) );
  XOR U19650 ( .A(n15202), .B(n15201), .Z(n15200) );
  XOR U19651 ( .A(y[1937]), .B(x[1937]), .Z(n15201) );
  XOR U19652 ( .A(y[1936]), .B(x[1936]), .Z(n15202) );
  XOR U19653 ( .A(n15194), .B(n15193), .Z(n15203) );
  XOR U19654 ( .A(n15196), .B(n15195), .Z(n15193) );
  XOR U19655 ( .A(y[1934]), .B(x[1934]), .Z(n15195) );
  XOR U19656 ( .A(y[1933]), .B(x[1933]), .Z(n15196) );
  XOR U19657 ( .A(y[1932]), .B(x[1932]), .Z(n15194) );
  XNOR U19658 ( .A(n15187), .B(n15186), .Z(n15189) );
  XNOR U19659 ( .A(n15183), .B(n15182), .Z(n15186) );
  XOR U19660 ( .A(n15185), .B(n15184), .Z(n15182) );
  XOR U19661 ( .A(y[1931]), .B(x[1931]), .Z(n15184) );
  XOR U19662 ( .A(y[1930]), .B(x[1930]), .Z(n15185) );
  XOR U19663 ( .A(y[1929]), .B(x[1929]), .Z(n15183) );
  XOR U19664 ( .A(n15177), .B(n15176), .Z(n15187) );
  XOR U19665 ( .A(n15179), .B(n15178), .Z(n15176) );
  XOR U19666 ( .A(y[1928]), .B(x[1928]), .Z(n15178) );
  XOR U19667 ( .A(y[1927]), .B(x[1927]), .Z(n15179) );
  XOR U19668 ( .A(y[1926]), .B(x[1926]), .Z(n15177) );
  NAND U19669 ( .A(n15240), .B(n15241), .Z(N28893) );
  NAND U19670 ( .A(n15242), .B(n15243), .Z(n15241) );
  NANDN U19671 ( .A(n15244), .B(n15245), .Z(n15243) );
  NANDN U19672 ( .A(n15245), .B(n15244), .Z(n15240) );
  XOR U19673 ( .A(n15244), .B(n15246), .Z(N28892) );
  XNOR U19674 ( .A(n15242), .B(n15245), .Z(n15246) );
  NAND U19675 ( .A(n15247), .B(n15248), .Z(n15245) );
  NAND U19676 ( .A(n15249), .B(n15250), .Z(n15248) );
  NANDN U19677 ( .A(n15251), .B(n15252), .Z(n15250) );
  NANDN U19678 ( .A(n15252), .B(n15251), .Z(n15247) );
  AND U19679 ( .A(n15253), .B(n15254), .Z(n15242) );
  NAND U19680 ( .A(n15255), .B(n15256), .Z(n15254) );
  OR U19681 ( .A(n15257), .B(n15258), .Z(n15256) );
  NAND U19682 ( .A(n15258), .B(n15257), .Z(n15253) );
  IV U19683 ( .A(n15259), .Z(n15258) );
  AND U19684 ( .A(n15260), .B(n15261), .Z(n15244) );
  NAND U19685 ( .A(n15262), .B(n15263), .Z(n15261) );
  NANDN U19686 ( .A(n15264), .B(n15265), .Z(n15263) );
  NANDN U19687 ( .A(n15265), .B(n15264), .Z(n15260) );
  XOR U19688 ( .A(n15257), .B(n15266), .Z(N28891) );
  XOR U19689 ( .A(n15255), .B(n15259), .Z(n15266) );
  XNOR U19690 ( .A(n15252), .B(n15267), .Z(n15259) );
  XNOR U19691 ( .A(n15249), .B(n15251), .Z(n15267) );
  AND U19692 ( .A(n15268), .B(n15269), .Z(n15251) );
  NANDN U19693 ( .A(n15270), .B(n15271), .Z(n15269) );
  NANDN U19694 ( .A(n15272), .B(n15273), .Z(n15271) );
  IV U19695 ( .A(n15274), .Z(n15273) );
  NAND U19696 ( .A(n15274), .B(n15272), .Z(n15268) );
  AND U19697 ( .A(n15275), .B(n15276), .Z(n15249) );
  NAND U19698 ( .A(n15277), .B(n15278), .Z(n15276) );
  OR U19699 ( .A(n15279), .B(n15280), .Z(n15278) );
  NAND U19700 ( .A(n15280), .B(n15279), .Z(n15275) );
  IV U19701 ( .A(n15281), .Z(n15280) );
  NAND U19702 ( .A(n15282), .B(n15283), .Z(n15252) );
  NANDN U19703 ( .A(n15284), .B(n15285), .Z(n15283) );
  NAND U19704 ( .A(n15286), .B(n15287), .Z(n15285) );
  OR U19705 ( .A(n15287), .B(n15286), .Z(n15282) );
  IV U19706 ( .A(n15288), .Z(n15286) );
  AND U19707 ( .A(n15289), .B(n15290), .Z(n15255) );
  NAND U19708 ( .A(n15291), .B(n15292), .Z(n15290) );
  NANDN U19709 ( .A(n15293), .B(n15294), .Z(n15292) );
  NANDN U19710 ( .A(n15294), .B(n15293), .Z(n15289) );
  XOR U19711 ( .A(n15265), .B(n15295), .Z(n15257) );
  XNOR U19712 ( .A(n15262), .B(n15264), .Z(n15295) );
  AND U19713 ( .A(n15296), .B(n15297), .Z(n15264) );
  NANDN U19714 ( .A(n15298), .B(n15299), .Z(n15297) );
  NANDN U19715 ( .A(n15300), .B(n15301), .Z(n15299) );
  IV U19716 ( .A(n15302), .Z(n15301) );
  NAND U19717 ( .A(n15302), .B(n15300), .Z(n15296) );
  AND U19718 ( .A(n15303), .B(n15304), .Z(n15262) );
  NAND U19719 ( .A(n15305), .B(n15306), .Z(n15304) );
  OR U19720 ( .A(n15307), .B(n15308), .Z(n15306) );
  NAND U19721 ( .A(n15308), .B(n15307), .Z(n15303) );
  IV U19722 ( .A(n15309), .Z(n15308) );
  NAND U19723 ( .A(n15310), .B(n15311), .Z(n15265) );
  NANDN U19724 ( .A(n15312), .B(n15313), .Z(n15311) );
  NAND U19725 ( .A(n15314), .B(n15315), .Z(n15313) );
  OR U19726 ( .A(n15315), .B(n15314), .Z(n15310) );
  IV U19727 ( .A(n15316), .Z(n15314) );
  XOR U19728 ( .A(n15291), .B(n15317), .Z(N28890) );
  XNOR U19729 ( .A(n15294), .B(n15293), .Z(n15317) );
  XNOR U19730 ( .A(n15305), .B(n15318), .Z(n15293) );
  XOR U19731 ( .A(n15309), .B(n15307), .Z(n15318) );
  XOR U19732 ( .A(n15315), .B(n15319), .Z(n15307) );
  XOR U19733 ( .A(n15312), .B(n15316), .Z(n15319) );
  NAND U19734 ( .A(n15320), .B(n15321), .Z(n15316) );
  NAND U19735 ( .A(n15322), .B(n15323), .Z(n15321) );
  NAND U19736 ( .A(n15324), .B(n15325), .Z(n15320) );
  AND U19737 ( .A(n15326), .B(n15327), .Z(n15312) );
  NAND U19738 ( .A(n15328), .B(n15329), .Z(n15327) );
  NAND U19739 ( .A(n15330), .B(n15331), .Z(n15326) );
  NANDN U19740 ( .A(n15332), .B(n15333), .Z(n15315) );
  NANDN U19741 ( .A(n15334), .B(n15335), .Z(n15309) );
  XNOR U19742 ( .A(n15300), .B(n15336), .Z(n15305) );
  XOR U19743 ( .A(n15298), .B(n15302), .Z(n15336) );
  NAND U19744 ( .A(n15337), .B(n15338), .Z(n15302) );
  NAND U19745 ( .A(n15339), .B(n15340), .Z(n15338) );
  NAND U19746 ( .A(n15341), .B(n15342), .Z(n15337) );
  AND U19747 ( .A(n15343), .B(n15344), .Z(n15298) );
  NAND U19748 ( .A(n15345), .B(n15346), .Z(n15344) );
  NAND U19749 ( .A(n15347), .B(n15348), .Z(n15343) );
  AND U19750 ( .A(n15349), .B(n15350), .Z(n15300) );
  NAND U19751 ( .A(n15351), .B(n15352), .Z(n15294) );
  XNOR U19752 ( .A(n15277), .B(n15353), .Z(n15291) );
  XOR U19753 ( .A(n15281), .B(n15279), .Z(n15353) );
  XOR U19754 ( .A(n15287), .B(n15354), .Z(n15279) );
  XOR U19755 ( .A(n15284), .B(n15288), .Z(n15354) );
  NAND U19756 ( .A(n15355), .B(n15356), .Z(n15288) );
  NAND U19757 ( .A(n15357), .B(n15358), .Z(n15356) );
  NAND U19758 ( .A(n15359), .B(n15360), .Z(n15355) );
  AND U19759 ( .A(n15361), .B(n15362), .Z(n15284) );
  NAND U19760 ( .A(n15363), .B(n15364), .Z(n15362) );
  NAND U19761 ( .A(n15365), .B(n15366), .Z(n15361) );
  NANDN U19762 ( .A(n15367), .B(n15368), .Z(n15287) );
  NANDN U19763 ( .A(n15369), .B(n15370), .Z(n15281) );
  XNOR U19764 ( .A(n15272), .B(n15371), .Z(n15277) );
  XOR U19765 ( .A(n15270), .B(n15274), .Z(n15371) );
  NAND U19766 ( .A(n15372), .B(n15373), .Z(n15274) );
  NAND U19767 ( .A(n15374), .B(n15375), .Z(n15373) );
  NAND U19768 ( .A(n15376), .B(n15377), .Z(n15372) );
  AND U19769 ( .A(n15378), .B(n15379), .Z(n15270) );
  NAND U19770 ( .A(n15380), .B(n15381), .Z(n15379) );
  NAND U19771 ( .A(n15382), .B(n15383), .Z(n15378) );
  AND U19772 ( .A(n15384), .B(n15385), .Z(n15272) );
  XOR U19773 ( .A(n15352), .B(n15351), .Z(N28889) );
  XNOR U19774 ( .A(n15370), .B(n15369), .Z(n15351) );
  XNOR U19775 ( .A(n15384), .B(n15385), .Z(n15369) );
  XOR U19776 ( .A(n15381), .B(n15380), .Z(n15385) );
  XOR U19777 ( .A(y[1923]), .B(x[1923]), .Z(n15380) );
  XOR U19778 ( .A(n15383), .B(n15382), .Z(n15381) );
  XOR U19779 ( .A(y[1925]), .B(x[1925]), .Z(n15382) );
  XOR U19780 ( .A(y[1924]), .B(x[1924]), .Z(n15383) );
  XOR U19781 ( .A(n15375), .B(n15374), .Z(n15384) );
  XOR U19782 ( .A(n15377), .B(n15376), .Z(n15374) );
  XOR U19783 ( .A(y[1922]), .B(x[1922]), .Z(n15376) );
  XOR U19784 ( .A(y[1921]), .B(x[1921]), .Z(n15377) );
  XOR U19785 ( .A(y[1920]), .B(x[1920]), .Z(n15375) );
  XNOR U19786 ( .A(n15368), .B(n15367), .Z(n15370) );
  XNOR U19787 ( .A(n15364), .B(n15363), .Z(n15367) );
  XOR U19788 ( .A(n15366), .B(n15365), .Z(n15363) );
  XOR U19789 ( .A(y[1919]), .B(x[1919]), .Z(n15365) );
  XOR U19790 ( .A(y[1918]), .B(x[1918]), .Z(n15366) );
  XOR U19791 ( .A(y[1917]), .B(x[1917]), .Z(n15364) );
  XOR U19792 ( .A(n15358), .B(n15357), .Z(n15368) );
  XOR U19793 ( .A(n15360), .B(n15359), .Z(n15357) );
  XOR U19794 ( .A(y[1916]), .B(x[1916]), .Z(n15359) );
  XOR U19795 ( .A(y[1915]), .B(x[1915]), .Z(n15360) );
  XOR U19796 ( .A(y[1914]), .B(x[1914]), .Z(n15358) );
  XNOR U19797 ( .A(n15335), .B(n15334), .Z(n15352) );
  XNOR U19798 ( .A(n15349), .B(n15350), .Z(n15334) );
  XOR U19799 ( .A(n15346), .B(n15345), .Z(n15350) );
  XOR U19800 ( .A(y[1911]), .B(x[1911]), .Z(n15345) );
  XOR U19801 ( .A(n15348), .B(n15347), .Z(n15346) );
  XOR U19802 ( .A(y[1913]), .B(x[1913]), .Z(n15347) );
  XOR U19803 ( .A(y[1912]), .B(x[1912]), .Z(n15348) );
  XOR U19804 ( .A(n15340), .B(n15339), .Z(n15349) );
  XOR U19805 ( .A(n15342), .B(n15341), .Z(n15339) );
  XOR U19806 ( .A(y[1910]), .B(x[1910]), .Z(n15341) );
  XOR U19807 ( .A(y[1909]), .B(x[1909]), .Z(n15342) );
  XOR U19808 ( .A(y[1908]), .B(x[1908]), .Z(n15340) );
  XNOR U19809 ( .A(n15333), .B(n15332), .Z(n15335) );
  XNOR U19810 ( .A(n15329), .B(n15328), .Z(n15332) );
  XOR U19811 ( .A(n15331), .B(n15330), .Z(n15328) );
  XOR U19812 ( .A(y[1907]), .B(x[1907]), .Z(n15330) );
  XOR U19813 ( .A(y[1906]), .B(x[1906]), .Z(n15331) );
  XOR U19814 ( .A(y[1905]), .B(x[1905]), .Z(n15329) );
  XOR U19815 ( .A(n15323), .B(n15322), .Z(n15333) );
  XOR U19816 ( .A(n15325), .B(n15324), .Z(n15322) );
  XOR U19817 ( .A(y[1904]), .B(x[1904]), .Z(n15324) );
  XOR U19818 ( .A(y[1903]), .B(x[1903]), .Z(n15325) );
  XOR U19819 ( .A(y[1902]), .B(x[1902]), .Z(n15323) );
  NAND U19820 ( .A(n15386), .B(n15387), .Z(N28881) );
  NAND U19821 ( .A(n15388), .B(n15389), .Z(n15387) );
  NANDN U19822 ( .A(n15390), .B(n15391), .Z(n15389) );
  NANDN U19823 ( .A(n15391), .B(n15390), .Z(n15386) );
  XOR U19824 ( .A(n15390), .B(n15392), .Z(N28880) );
  XNOR U19825 ( .A(n15388), .B(n15391), .Z(n15392) );
  NAND U19826 ( .A(n15393), .B(n15394), .Z(n15391) );
  NAND U19827 ( .A(n15395), .B(n15396), .Z(n15394) );
  NANDN U19828 ( .A(n15397), .B(n15398), .Z(n15396) );
  NANDN U19829 ( .A(n15398), .B(n15397), .Z(n15393) );
  AND U19830 ( .A(n15399), .B(n15400), .Z(n15388) );
  NAND U19831 ( .A(n15401), .B(n15402), .Z(n15400) );
  OR U19832 ( .A(n15403), .B(n15404), .Z(n15402) );
  NAND U19833 ( .A(n15404), .B(n15403), .Z(n15399) );
  IV U19834 ( .A(n15405), .Z(n15404) );
  AND U19835 ( .A(n15406), .B(n15407), .Z(n15390) );
  NAND U19836 ( .A(n15408), .B(n15409), .Z(n15407) );
  NANDN U19837 ( .A(n15410), .B(n15411), .Z(n15409) );
  NANDN U19838 ( .A(n15411), .B(n15410), .Z(n15406) );
  XOR U19839 ( .A(n15403), .B(n15412), .Z(N28879) );
  XOR U19840 ( .A(n15401), .B(n15405), .Z(n15412) );
  XNOR U19841 ( .A(n15398), .B(n15413), .Z(n15405) );
  XNOR U19842 ( .A(n15395), .B(n15397), .Z(n15413) );
  AND U19843 ( .A(n15414), .B(n15415), .Z(n15397) );
  NANDN U19844 ( .A(n15416), .B(n15417), .Z(n15415) );
  NANDN U19845 ( .A(n15418), .B(n15419), .Z(n15417) );
  IV U19846 ( .A(n15420), .Z(n15419) );
  NAND U19847 ( .A(n15420), .B(n15418), .Z(n15414) );
  AND U19848 ( .A(n15421), .B(n15422), .Z(n15395) );
  NAND U19849 ( .A(n15423), .B(n15424), .Z(n15422) );
  OR U19850 ( .A(n15425), .B(n15426), .Z(n15424) );
  NAND U19851 ( .A(n15426), .B(n15425), .Z(n15421) );
  IV U19852 ( .A(n15427), .Z(n15426) );
  NAND U19853 ( .A(n15428), .B(n15429), .Z(n15398) );
  NANDN U19854 ( .A(n15430), .B(n15431), .Z(n15429) );
  NAND U19855 ( .A(n15432), .B(n15433), .Z(n15431) );
  OR U19856 ( .A(n15433), .B(n15432), .Z(n15428) );
  IV U19857 ( .A(n15434), .Z(n15432) );
  AND U19858 ( .A(n15435), .B(n15436), .Z(n15401) );
  NAND U19859 ( .A(n15437), .B(n15438), .Z(n15436) );
  NANDN U19860 ( .A(n15439), .B(n15440), .Z(n15438) );
  NANDN U19861 ( .A(n15440), .B(n15439), .Z(n15435) );
  XOR U19862 ( .A(n15411), .B(n15441), .Z(n15403) );
  XNOR U19863 ( .A(n15408), .B(n15410), .Z(n15441) );
  AND U19864 ( .A(n15442), .B(n15443), .Z(n15410) );
  NANDN U19865 ( .A(n15444), .B(n15445), .Z(n15443) );
  NANDN U19866 ( .A(n15446), .B(n15447), .Z(n15445) );
  IV U19867 ( .A(n15448), .Z(n15447) );
  NAND U19868 ( .A(n15448), .B(n15446), .Z(n15442) );
  AND U19869 ( .A(n15449), .B(n15450), .Z(n15408) );
  NAND U19870 ( .A(n15451), .B(n15452), .Z(n15450) );
  OR U19871 ( .A(n15453), .B(n15454), .Z(n15452) );
  NAND U19872 ( .A(n15454), .B(n15453), .Z(n15449) );
  IV U19873 ( .A(n15455), .Z(n15454) );
  NAND U19874 ( .A(n15456), .B(n15457), .Z(n15411) );
  NANDN U19875 ( .A(n15458), .B(n15459), .Z(n15457) );
  NAND U19876 ( .A(n15460), .B(n15461), .Z(n15459) );
  OR U19877 ( .A(n15461), .B(n15460), .Z(n15456) );
  IV U19878 ( .A(n15462), .Z(n15460) );
  XOR U19879 ( .A(n15437), .B(n15463), .Z(N28878) );
  XNOR U19880 ( .A(n15440), .B(n15439), .Z(n15463) );
  XNOR U19881 ( .A(n15451), .B(n15464), .Z(n15439) );
  XOR U19882 ( .A(n15455), .B(n15453), .Z(n15464) );
  XOR U19883 ( .A(n15461), .B(n15465), .Z(n15453) );
  XOR U19884 ( .A(n15458), .B(n15462), .Z(n15465) );
  NAND U19885 ( .A(n15466), .B(n15467), .Z(n15462) );
  NAND U19886 ( .A(n15468), .B(n15469), .Z(n15467) );
  NAND U19887 ( .A(n15470), .B(n15471), .Z(n15466) );
  AND U19888 ( .A(n15472), .B(n15473), .Z(n15458) );
  NAND U19889 ( .A(n15474), .B(n15475), .Z(n15473) );
  NAND U19890 ( .A(n15476), .B(n15477), .Z(n15472) );
  NANDN U19891 ( .A(n15478), .B(n15479), .Z(n15461) );
  NANDN U19892 ( .A(n15480), .B(n15481), .Z(n15455) );
  XNOR U19893 ( .A(n15446), .B(n15482), .Z(n15451) );
  XOR U19894 ( .A(n15444), .B(n15448), .Z(n15482) );
  NAND U19895 ( .A(n15483), .B(n15484), .Z(n15448) );
  NAND U19896 ( .A(n15485), .B(n15486), .Z(n15484) );
  NAND U19897 ( .A(n15487), .B(n15488), .Z(n15483) );
  AND U19898 ( .A(n15489), .B(n15490), .Z(n15444) );
  NAND U19899 ( .A(n15491), .B(n15492), .Z(n15490) );
  NAND U19900 ( .A(n15493), .B(n15494), .Z(n15489) );
  AND U19901 ( .A(n15495), .B(n15496), .Z(n15446) );
  NAND U19902 ( .A(n15497), .B(n15498), .Z(n15440) );
  XNOR U19903 ( .A(n15423), .B(n15499), .Z(n15437) );
  XOR U19904 ( .A(n15427), .B(n15425), .Z(n15499) );
  XOR U19905 ( .A(n15433), .B(n15500), .Z(n15425) );
  XOR U19906 ( .A(n15430), .B(n15434), .Z(n15500) );
  NAND U19907 ( .A(n15501), .B(n15502), .Z(n15434) );
  NAND U19908 ( .A(n15503), .B(n15504), .Z(n15502) );
  NAND U19909 ( .A(n15505), .B(n15506), .Z(n15501) );
  AND U19910 ( .A(n15507), .B(n15508), .Z(n15430) );
  NAND U19911 ( .A(n15509), .B(n15510), .Z(n15508) );
  NAND U19912 ( .A(n15511), .B(n15512), .Z(n15507) );
  NANDN U19913 ( .A(n15513), .B(n15514), .Z(n15433) );
  NANDN U19914 ( .A(n15515), .B(n15516), .Z(n15427) );
  XNOR U19915 ( .A(n15418), .B(n15517), .Z(n15423) );
  XOR U19916 ( .A(n15416), .B(n15420), .Z(n15517) );
  NAND U19917 ( .A(n15518), .B(n15519), .Z(n15420) );
  NAND U19918 ( .A(n15520), .B(n15521), .Z(n15519) );
  NAND U19919 ( .A(n15522), .B(n15523), .Z(n15518) );
  AND U19920 ( .A(n15524), .B(n15525), .Z(n15416) );
  NAND U19921 ( .A(n15526), .B(n15527), .Z(n15525) );
  NAND U19922 ( .A(n15528), .B(n15529), .Z(n15524) );
  AND U19923 ( .A(n15530), .B(n15531), .Z(n15418) );
  XOR U19924 ( .A(n15498), .B(n15497), .Z(N28877) );
  XNOR U19925 ( .A(n15516), .B(n15515), .Z(n15497) );
  XNOR U19926 ( .A(n15530), .B(n15531), .Z(n15515) );
  XOR U19927 ( .A(n15527), .B(n15526), .Z(n15531) );
  XOR U19928 ( .A(y[1899]), .B(x[1899]), .Z(n15526) );
  XOR U19929 ( .A(n15529), .B(n15528), .Z(n15527) );
  XOR U19930 ( .A(y[1901]), .B(x[1901]), .Z(n15528) );
  XOR U19931 ( .A(y[1900]), .B(x[1900]), .Z(n15529) );
  XOR U19932 ( .A(n15521), .B(n15520), .Z(n15530) );
  XOR U19933 ( .A(n15523), .B(n15522), .Z(n15520) );
  XOR U19934 ( .A(y[1898]), .B(x[1898]), .Z(n15522) );
  XOR U19935 ( .A(y[1897]), .B(x[1897]), .Z(n15523) );
  XOR U19936 ( .A(y[1896]), .B(x[1896]), .Z(n15521) );
  XNOR U19937 ( .A(n15514), .B(n15513), .Z(n15516) );
  XNOR U19938 ( .A(n15510), .B(n15509), .Z(n15513) );
  XOR U19939 ( .A(n15512), .B(n15511), .Z(n15509) );
  XOR U19940 ( .A(y[1895]), .B(x[1895]), .Z(n15511) );
  XOR U19941 ( .A(y[1894]), .B(x[1894]), .Z(n15512) );
  XOR U19942 ( .A(y[1893]), .B(x[1893]), .Z(n15510) );
  XOR U19943 ( .A(n15504), .B(n15503), .Z(n15514) );
  XOR U19944 ( .A(n15506), .B(n15505), .Z(n15503) );
  XOR U19945 ( .A(y[1892]), .B(x[1892]), .Z(n15505) );
  XOR U19946 ( .A(y[1891]), .B(x[1891]), .Z(n15506) );
  XOR U19947 ( .A(y[1890]), .B(x[1890]), .Z(n15504) );
  XNOR U19948 ( .A(n15481), .B(n15480), .Z(n15498) );
  XNOR U19949 ( .A(n15495), .B(n15496), .Z(n15480) );
  XOR U19950 ( .A(n15492), .B(n15491), .Z(n15496) );
  XOR U19951 ( .A(y[1887]), .B(x[1887]), .Z(n15491) );
  XOR U19952 ( .A(n15494), .B(n15493), .Z(n15492) );
  XOR U19953 ( .A(y[1889]), .B(x[1889]), .Z(n15493) );
  XOR U19954 ( .A(y[1888]), .B(x[1888]), .Z(n15494) );
  XOR U19955 ( .A(n15486), .B(n15485), .Z(n15495) );
  XOR U19956 ( .A(n15488), .B(n15487), .Z(n15485) );
  XOR U19957 ( .A(y[1886]), .B(x[1886]), .Z(n15487) );
  XOR U19958 ( .A(y[1885]), .B(x[1885]), .Z(n15488) );
  XOR U19959 ( .A(y[1884]), .B(x[1884]), .Z(n15486) );
  XNOR U19960 ( .A(n15479), .B(n15478), .Z(n15481) );
  XNOR U19961 ( .A(n15475), .B(n15474), .Z(n15478) );
  XOR U19962 ( .A(n15477), .B(n15476), .Z(n15474) );
  XOR U19963 ( .A(y[1883]), .B(x[1883]), .Z(n15476) );
  XOR U19964 ( .A(y[1882]), .B(x[1882]), .Z(n15477) );
  XOR U19965 ( .A(y[1881]), .B(x[1881]), .Z(n15475) );
  XOR U19966 ( .A(n15469), .B(n15468), .Z(n15479) );
  XOR U19967 ( .A(n15471), .B(n15470), .Z(n15468) );
  XOR U19968 ( .A(y[1880]), .B(x[1880]), .Z(n15470) );
  XOR U19969 ( .A(y[1879]), .B(x[1879]), .Z(n15471) );
  XOR U19970 ( .A(y[1878]), .B(x[1878]), .Z(n15469) );
  NAND U19971 ( .A(n15532), .B(n15533), .Z(N28869) );
  NAND U19972 ( .A(n15534), .B(n15535), .Z(n15533) );
  NANDN U19973 ( .A(n15536), .B(n15537), .Z(n15535) );
  NANDN U19974 ( .A(n15537), .B(n15536), .Z(n15532) );
  XOR U19975 ( .A(n15536), .B(n15538), .Z(N28868) );
  XNOR U19976 ( .A(n15534), .B(n15537), .Z(n15538) );
  NAND U19977 ( .A(n15539), .B(n15540), .Z(n15537) );
  NAND U19978 ( .A(n15541), .B(n15542), .Z(n15540) );
  NANDN U19979 ( .A(n15543), .B(n15544), .Z(n15542) );
  NANDN U19980 ( .A(n15544), .B(n15543), .Z(n15539) );
  AND U19981 ( .A(n15545), .B(n15546), .Z(n15534) );
  NAND U19982 ( .A(n15547), .B(n15548), .Z(n15546) );
  OR U19983 ( .A(n15549), .B(n15550), .Z(n15548) );
  NAND U19984 ( .A(n15550), .B(n15549), .Z(n15545) );
  IV U19985 ( .A(n15551), .Z(n15550) );
  AND U19986 ( .A(n15552), .B(n15553), .Z(n15536) );
  NAND U19987 ( .A(n15554), .B(n15555), .Z(n15553) );
  NANDN U19988 ( .A(n15556), .B(n15557), .Z(n15555) );
  NANDN U19989 ( .A(n15557), .B(n15556), .Z(n15552) );
  XOR U19990 ( .A(n15549), .B(n15558), .Z(N28867) );
  XOR U19991 ( .A(n15547), .B(n15551), .Z(n15558) );
  XNOR U19992 ( .A(n15544), .B(n15559), .Z(n15551) );
  XNOR U19993 ( .A(n15541), .B(n15543), .Z(n15559) );
  AND U19994 ( .A(n15560), .B(n15561), .Z(n15543) );
  NANDN U19995 ( .A(n15562), .B(n15563), .Z(n15561) );
  NANDN U19996 ( .A(n15564), .B(n15565), .Z(n15563) );
  IV U19997 ( .A(n15566), .Z(n15565) );
  NAND U19998 ( .A(n15566), .B(n15564), .Z(n15560) );
  AND U19999 ( .A(n15567), .B(n15568), .Z(n15541) );
  NAND U20000 ( .A(n15569), .B(n15570), .Z(n15568) );
  OR U20001 ( .A(n15571), .B(n15572), .Z(n15570) );
  NAND U20002 ( .A(n15572), .B(n15571), .Z(n15567) );
  IV U20003 ( .A(n15573), .Z(n15572) );
  NAND U20004 ( .A(n15574), .B(n15575), .Z(n15544) );
  NANDN U20005 ( .A(n15576), .B(n15577), .Z(n15575) );
  NAND U20006 ( .A(n15578), .B(n15579), .Z(n15577) );
  OR U20007 ( .A(n15579), .B(n15578), .Z(n15574) );
  IV U20008 ( .A(n15580), .Z(n15578) );
  AND U20009 ( .A(n15581), .B(n15582), .Z(n15547) );
  NAND U20010 ( .A(n15583), .B(n15584), .Z(n15582) );
  NANDN U20011 ( .A(n15585), .B(n15586), .Z(n15584) );
  NANDN U20012 ( .A(n15586), .B(n15585), .Z(n15581) );
  XOR U20013 ( .A(n15557), .B(n15587), .Z(n15549) );
  XNOR U20014 ( .A(n15554), .B(n15556), .Z(n15587) );
  AND U20015 ( .A(n15588), .B(n15589), .Z(n15556) );
  NANDN U20016 ( .A(n15590), .B(n15591), .Z(n15589) );
  NANDN U20017 ( .A(n15592), .B(n15593), .Z(n15591) );
  IV U20018 ( .A(n15594), .Z(n15593) );
  NAND U20019 ( .A(n15594), .B(n15592), .Z(n15588) );
  AND U20020 ( .A(n15595), .B(n15596), .Z(n15554) );
  NAND U20021 ( .A(n15597), .B(n15598), .Z(n15596) );
  OR U20022 ( .A(n15599), .B(n15600), .Z(n15598) );
  NAND U20023 ( .A(n15600), .B(n15599), .Z(n15595) );
  IV U20024 ( .A(n15601), .Z(n15600) );
  NAND U20025 ( .A(n15602), .B(n15603), .Z(n15557) );
  NANDN U20026 ( .A(n15604), .B(n15605), .Z(n15603) );
  NAND U20027 ( .A(n15606), .B(n15607), .Z(n15605) );
  OR U20028 ( .A(n15607), .B(n15606), .Z(n15602) );
  IV U20029 ( .A(n15608), .Z(n15606) );
  XOR U20030 ( .A(n15583), .B(n15609), .Z(N28866) );
  XNOR U20031 ( .A(n15586), .B(n15585), .Z(n15609) );
  XNOR U20032 ( .A(n15597), .B(n15610), .Z(n15585) );
  XOR U20033 ( .A(n15601), .B(n15599), .Z(n15610) );
  XOR U20034 ( .A(n15607), .B(n15611), .Z(n15599) );
  XOR U20035 ( .A(n15604), .B(n15608), .Z(n15611) );
  NAND U20036 ( .A(n15612), .B(n15613), .Z(n15608) );
  NAND U20037 ( .A(n15614), .B(n15615), .Z(n15613) );
  NAND U20038 ( .A(n15616), .B(n15617), .Z(n15612) );
  AND U20039 ( .A(n15618), .B(n15619), .Z(n15604) );
  NAND U20040 ( .A(n15620), .B(n15621), .Z(n15619) );
  NAND U20041 ( .A(n15622), .B(n15623), .Z(n15618) );
  NANDN U20042 ( .A(n15624), .B(n15625), .Z(n15607) );
  NANDN U20043 ( .A(n15626), .B(n15627), .Z(n15601) );
  XNOR U20044 ( .A(n15592), .B(n15628), .Z(n15597) );
  XOR U20045 ( .A(n15590), .B(n15594), .Z(n15628) );
  NAND U20046 ( .A(n15629), .B(n15630), .Z(n15594) );
  NAND U20047 ( .A(n15631), .B(n15632), .Z(n15630) );
  NAND U20048 ( .A(n15633), .B(n15634), .Z(n15629) );
  AND U20049 ( .A(n15635), .B(n15636), .Z(n15590) );
  NAND U20050 ( .A(n15637), .B(n15638), .Z(n15636) );
  NAND U20051 ( .A(n15639), .B(n15640), .Z(n15635) );
  AND U20052 ( .A(n15641), .B(n15642), .Z(n15592) );
  NAND U20053 ( .A(n15643), .B(n15644), .Z(n15586) );
  XNOR U20054 ( .A(n15569), .B(n15645), .Z(n15583) );
  XOR U20055 ( .A(n15573), .B(n15571), .Z(n15645) );
  XOR U20056 ( .A(n15579), .B(n15646), .Z(n15571) );
  XOR U20057 ( .A(n15576), .B(n15580), .Z(n15646) );
  NAND U20058 ( .A(n15647), .B(n15648), .Z(n15580) );
  NAND U20059 ( .A(n15649), .B(n15650), .Z(n15648) );
  NAND U20060 ( .A(n15651), .B(n15652), .Z(n15647) );
  AND U20061 ( .A(n15653), .B(n15654), .Z(n15576) );
  NAND U20062 ( .A(n15655), .B(n15656), .Z(n15654) );
  NAND U20063 ( .A(n15657), .B(n15658), .Z(n15653) );
  NANDN U20064 ( .A(n15659), .B(n15660), .Z(n15579) );
  NANDN U20065 ( .A(n15661), .B(n15662), .Z(n15573) );
  XNOR U20066 ( .A(n15564), .B(n15663), .Z(n15569) );
  XOR U20067 ( .A(n15562), .B(n15566), .Z(n15663) );
  NAND U20068 ( .A(n15664), .B(n15665), .Z(n15566) );
  NAND U20069 ( .A(n15666), .B(n15667), .Z(n15665) );
  NAND U20070 ( .A(n15668), .B(n15669), .Z(n15664) );
  AND U20071 ( .A(n15670), .B(n15671), .Z(n15562) );
  NAND U20072 ( .A(n15672), .B(n15673), .Z(n15671) );
  NAND U20073 ( .A(n15674), .B(n15675), .Z(n15670) );
  AND U20074 ( .A(n15676), .B(n15677), .Z(n15564) );
  XOR U20075 ( .A(n15644), .B(n15643), .Z(N28865) );
  XNOR U20076 ( .A(n15662), .B(n15661), .Z(n15643) );
  XNOR U20077 ( .A(n15676), .B(n15677), .Z(n15661) );
  XOR U20078 ( .A(n15673), .B(n15672), .Z(n15677) );
  XOR U20079 ( .A(y[1875]), .B(x[1875]), .Z(n15672) );
  XOR U20080 ( .A(n15675), .B(n15674), .Z(n15673) );
  XOR U20081 ( .A(y[1877]), .B(x[1877]), .Z(n15674) );
  XOR U20082 ( .A(y[1876]), .B(x[1876]), .Z(n15675) );
  XOR U20083 ( .A(n15667), .B(n15666), .Z(n15676) );
  XOR U20084 ( .A(n15669), .B(n15668), .Z(n15666) );
  XOR U20085 ( .A(y[1874]), .B(x[1874]), .Z(n15668) );
  XOR U20086 ( .A(y[1873]), .B(x[1873]), .Z(n15669) );
  XOR U20087 ( .A(y[1872]), .B(x[1872]), .Z(n15667) );
  XNOR U20088 ( .A(n15660), .B(n15659), .Z(n15662) );
  XNOR U20089 ( .A(n15656), .B(n15655), .Z(n15659) );
  XOR U20090 ( .A(n15658), .B(n15657), .Z(n15655) );
  XOR U20091 ( .A(y[1871]), .B(x[1871]), .Z(n15657) );
  XOR U20092 ( .A(y[1870]), .B(x[1870]), .Z(n15658) );
  XOR U20093 ( .A(y[1869]), .B(x[1869]), .Z(n15656) );
  XOR U20094 ( .A(n15650), .B(n15649), .Z(n15660) );
  XOR U20095 ( .A(n15652), .B(n15651), .Z(n15649) );
  XOR U20096 ( .A(y[1868]), .B(x[1868]), .Z(n15651) );
  XOR U20097 ( .A(y[1867]), .B(x[1867]), .Z(n15652) );
  XOR U20098 ( .A(y[1866]), .B(x[1866]), .Z(n15650) );
  XNOR U20099 ( .A(n15627), .B(n15626), .Z(n15644) );
  XNOR U20100 ( .A(n15641), .B(n15642), .Z(n15626) );
  XOR U20101 ( .A(n15638), .B(n15637), .Z(n15642) );
  XOR U20102 ( .A(y[1863]), .B(x[1863]), .Z(n15637) );
  XOR U20103 ( .A(n15640), .B(n15639), .Z(n15638) );
  XOR U20104 ( .A(y[1865]), .B(x[1865]), .Z(n15639) );
  XOR U20105 ( .A(y[1864]), .B(x[1864]), .Z(n15640) );
  XOR U20106 ( .A(n15632), .B(n15631), .Z(n15641) );
  XOR U20107 ( .A(n15634), .B(n15633), .Z(n15631) );
  XOR U20108 ( .A(y[1862]), .B(x[1862]), .Z(n15633) );
  XOR U20109 ( .A(y[1861]), .B(x[1861]), .Z(n15634) );
  XOR U20110 ( .A(y[1860]), .B(x[1860]), .Z(n15632) );
  XNOR U20111 ( .A(n15625), .B(n15624), .Z(n15627) );
  XNOR U20112 ( .A(n15621), .B(n15620), .Z(n15624) );
  XOR U20113 ( .A(n15623), .B(n15622), .Z(n15620) );
  XOR U20114 ( .A(y[1859]), .B(x[1859]), .Z(n15622) );
  XOR U20115 ( .A(y[1858]), .B(x[1858]), .Z(n15623) );
  XOR U20116 ( .A(y[1857]), .B(x[1857]), .Z(n15621) );
  XOR U20117 ( .A(n15615), .B(n15614), .Z(n15625) );
  XOR U20118 ( .A(n15617), .B(n15616), .Z(n15614) );
  XOR U20119 ( .A(y[1856]), .B(x[1856]), .Z(n15616) );
  XOR U20120 ( .A(y[1855]), .B(x[1855]), .Z(n15617) );
  XOR U20121 ( .A(y[1854]), .B(x[1854]), .Z(n15615) );
  NAND U20122 ( .A(n15678), .B(n15679), .Z(N28857) );
  NAND U20123 ( .A(n15680), .B(n15681), .Z(n15679) );
  NANDN U20124 ( .A(n15682), .B(n15683), .Z(n15681) );
  NANDN U20125 ( .A(n15683), .B(n15682), .Z(n15678) );
  XOR U20126 ( .A(n15682), .B(n15684), .Z(N28856) );
  XNOR U20127 ( .A(n15680), .B(n15683), .Z(n15684) );
  NAND U20128 ( .A(n15685), .B(n15686), .Z(n15683) );
  NAND U20129 ( .A(n15687), .B(n15688), .Z(n15686) );
  NANDN U20130 ( .A(n15689), .B(n15690), .Z(n15688) );
  NANDN U20131 ( .A(n15690), .B(n15689), .Z(n15685) );
  AND U20132 ( .A(n15691), .B(n15692), .Z(n15680) );
  NAND U20133 ( .A(n15693), .B(n15694), .Z(n15692) );
  OR U20134 ( .A(n15695), .B(n15696), .Z(n15694) );
  NAND U20135 ( .A(n15696), .B(n15695), .Z(n15691) );
  IV U20136 ( .A(n15697), .Z(n15696) );
  AND U20137 ( .A(n15698), .B(n15699), .Z(n15682) );
  NAND U20138 ( .A(n15700), .B(n15701), .Z(n15699) );
  NANDN U20139 ( .A(n15702), .B(n15703), .Z(n15701) );
  NANDN U20140 ( .A(n15703), .B(n15702), .Z(n15698) );
  XOR U20141 ( .A(n15695), .B(n15704), .Z(N28855) );
  XOR U20142 ( .A(n15693), .B(n15697), .Z(n15704) );
  XNOR U20143 ( .A(n15690), .B(n15705), .Z(n15697) );
  XNOR U20144 ( .A(n15687), .B(n15689), .Z(n15705) );
  AND U20145 ( .A(n15706), .B(n15707), .Z(n15689) );
  NANDN U20146 ( .A(n15708), .B(n15709), .Z(n15707) );
  NANDN U20147 ( .A(n15710), .B(n15711), .Z(n15709) );
  IV U20148 ( .A(n15712), .Z(n15711) );
  NAND U20149 ( .A(n15712), .B(n15710), .Z(n15706) );
  AND U20150 ( .A(n15713), .B(n15714), .Z(n15687) );
  NAND U20151 ( .A(n15715), .B(n15716), .Z(n15714) );
  OR U20152 ( .A(n15717), .B(n15718), .Z(n15716) );
  NAND U20153 ( .A(n15718), .B(n15717), .Z(n15713) );
  IV U20154 ( .A(n15719), .Z(n15718) );
  NAND U20155 ( .A(n15720), .B(n15721), .Z(n15690) );
  NANDN U20156 ( .A(n15722), .B(n15723), .Z(n15721) );
  NAND U20157 ( .A(n15724), .B(n15725), .Z(n15723) );
  OR U20158 ( .A(n15725), .B(n15724), .Z(n15720) );
  IV U20159 ( .A(n15726), .Z(n15724) );
  AND U20160 ( .A(n15727), .B(n15728), .Z(n15693) );
  NAND U20161 ( .A(n15729), .B(n15730), .Z(n15728) );
  NANDN U20162 ( .A(n15731), .B(n15732), .Z(n15730) );
  NANDN U20163 ( .A(n15732), .B(n15731), .Z(n15727) );
  XOR U20164 ( .A(n15703), .B(n15733), .Z(n15695) );
  XNOR U20165 ( .A(n15700), .B(n15702), .Z(n15733) );
  AND U20166 ( .A(n15734), .B(n15735), .Z(n15702) );
  NANDN U20167 ( .A(n15736), .B(n15737), .Z(n15735) );
  NANDN U20168 ( .A(n15738), .B(n15739), .Z(n15737) );
  IV U20169 ( .A(n15740), .Z(n15739) );
  NAND U20170 ( .A(n15740), .B(n15738), .Z(n15734) );
  AND U20171 ( .A(n15741), .B(n15742), .Z(n15700) );
  NAND U20172 ( .A(n15743), .B(n15744), .Z(n15742) );
  OR U20173 ( .A(n15745), .B(n15746), .Z(n15744) );
  NAND U20174 ( .A(n15746), .B(n15745), .Z(n15741) );
  IV U20175 ( .A(n15747), .Z(n15746) );
  NAND U20176 ( .A(n15748), .B(n15749), .Z(n15703) );
  NANDN U20177 ( .A(n15750), .B(n15751), .Z(n15749) );
  NAND U20178 ( .A(n15752), .B(n15753), .Z(n15751) );
  OR U20179 ( .A(n15753), .B(n15752), .Z(n15748) );
  IV U20180 ( .A(n15754), .Z(n15752) );
  XOR U20181 ( .A(n15729), .B(n15755), .Z(N28854) );
  XNOR U20182 ( .A(n15732), .B(n15731), .Z(n15755) );
  XNOR U20183 ( .A(n15743), .B(n15756), .Z(n15731) );
  XOR U20184 ( .A(n15747), .B(n15745), .Z(n15756) );
  XOR U20185 ( .A(n15753), .B(n15757), .Z(n15745) );
  XOR U20186 ( .A(n15750), .B(n15754), .Z(n15757) );
  NAND U20187 ( .A(n15758), .B(n15759), .Z(n15754) );
  NAND U20188 ( .A(n15760), .B(n15761), .Z(n15759) );
  NAND U20189 ( .A(n15762), .B(n15763), .Z(n15758) );
  AND U20190 ( .A(n15764), .B(n15765), .Z(n15750) );
  NAND U20191 ( .A(n15766), .B(n15767), .Z(n15765) );
  NAND U20192 ( .A(n15768), .B(n15769), .Z(n15764) );
  NANDN U20193 ( .A(n15770), .B(n15771), .Z(n15753) );
  NANDN U20194 ( .A(n15772), .B(n15773), .Z(n15747) );
  XNOR U20195 ( .A(n15738), .B(n15774), .Z(n15743) );
  XOR U20196 ( .A(n15736), .B(n15740), .Z(n15774) );
  NAND U20197 ( .A(n15775), .B(n15776), .Z(n15740) );
  NAND U20198 ( .A(n15777), .B(n15778), .Z(n15776) );
  NAND U20199 ( .A(n15779), .B(n15780), .Z(n15775) );
  AND U20200 ( .A(n15781), .B(n15782), .Z(n15736) );
  NAND U20201 ( .A(n15783), .B(n15784), .Z(n15782) );
  NAND U20202 ( .A(n15785), .B(n15786), .Z(n15781) );
  AND U20203 ( .A(n15787), .B(n15788), .Z(n15738) );
  NAND U20204 ( .A(n15789), .B(n15790), .Z(n15732) );
  XNOR U20205 ( .A(n15715), .B(n15791), .Z(n15729) );
  XOR U20206 ( .A(n15719), .B(n15717), .Z(n15791) );
  XOR U20207 ( .A(n15725), .B(n15792), .Z(n15717) );
  XOR U20208 ( .A(n15722), .B(n15726), .Z(n15792) );
  NAND U20209 ( .A(n15793), .B(n15794), .Z(n15726) );
  NAND U20210 ( .A(n15795), .B(n15796), .Z(n15794) );
  NAND U20211 ( .A(n15797), .B(n15798), .Z(n15793) );
  AND U20212 ( .A(n15799), .B(n15800), .Z(n15722) );
  NAND U20213 ( .A(n15801), .B(n15802), .Z(n15800) );
  NAND U20214 ( .A(n15803), .B(n15804), .Z(n15799) );
  NANDN U20215 ( .A(n15805), .B(n15806), .Z(n15725) );
  NANDN U20216 ( .A(n15807), .B(n15808), .Z(n15719) );
  XNOR U20217 ( .A(n15710), .B(n15809), .Z(n15715) );
  XOR U20218 ( .A(n15708), .B(n15712), .Z(n15809) );
  NAND U20219 ( .A(n15810), .B(n15811), .Z(n15712) );
  NAND U20220 ( .A(n15812), .B(n15813), .Z(n15811) );
  NAND U20221 ( .A(n15814), .B(n15815), .Z(n15810) );
  AND U20222 ( .A(n15816), .B(n15817), .Z(n15708) );
  NAND U20223 ( .A(n15818), .B(n15819), .Z(n15817) );
  NAND U20224 ( .A(n15820), .B(n15821), .Z(n15816) );
  AND U20225 ( .A(n15822), .B(n15823), .Z(n15710) );
  XOR U20226 ( .A(n15790), .B(n15789), .Z(N28853) );
  XNOR U20227 ( .A(n15808), .B(n15807), .Z(n15789) );
  XNOR U20228 ( .A(n15822), .B(n15823), .Z(n15807) );
  XOR U20229 ( .A(n15819), .B(n15818), .Z(n15823) );
  XOR U20230 ( .A(y[1851]), .B(x[1851]), .Z(n15818) );
  XOR U20231 ( .A(n15821), .B(n15820), .Z(n15819) );
  XOR U20232 ( .A(y[1853]), .B(x[1853]), .Z(n15820) );
  XOR U20233 ( .A(y[1852]), .B(x[1852]), .Z(n15821) );
  XOR U20234 ( .A(n15813), .B(n15812), .Z(n15822) );
  XOR U20235 ( .A(n15815), .B(n15814), .Z(n15812) );
  XOR U20236 ( .A(y[1850]), .B(x[1850]), .Z(n15814) );
  XOR U20237 ( .A(y[1849]), .B(x[1849]), .Z(n15815) );
  XOR U20238 ( .A(y[1848]), .B(x[1848]), .Z(n15813) );
  XNOR U20239 ( .A(n15806), .B(n15805), .Z(n15808) );
  XNOR U20240 ( .A(n15802), .B(n15801), .Z(n15805) );
  XOR U20241 ( .A(n15804), .B(n15803), .Z(n15801) );
  XOR U20242 ( .A(y[1847]), .B(x[1847]), .Z(n15803) );
  XOR U20243 ( .A(y[1846]), .B(x[1846]), .Z(n15804) );
  XOR U20244 ( .A(y[1845]), .B(x[1845]), .Z(n15802) );
  XOR U20245 ( .A(n15796), .B(n15795), .Z(n15806) );
  XOR U20246 ( .A(n15798), .B(n15797), .Z(n15795) );
  XOR U20247 ( .A(y[1844]), .B(x[1844]), .Z(n15797) );
  XOR U20248 ( .A(y[1843]), .B(x[1843]), .Z(n15798) );
  XOR U20249 ( .A(y[1842]), .B(x[1842]), .Z(n15796) );
  XNOR U20250 ( .A(n15773), .B(n15772), .Z(n15790) );
  XNOR U20251 ( .A(n15787), .B(n15788), .Z(n15772) );
  XOR U20252 ( .A(n15784), .B(n15783), .Z(n15788) );
  XOR U20253 ( .A(y[1839]), .B(x[1839]), .Z(n15783) );
  XOR U20254 ( .A(n15786), .B(n15785), .Z(n15784) );
  XOR U20255 ( .A(y[1841]), .B(x[1841]), .Z(n15785) );
  XOR U20256 ( .A(y[1840]), .B(x[1840]), .Z(n15786) );
  XOR U20257 ( .A(n15778), .B(n15777), .Z(n15787) );
  XOR U20258 ( .A(n15780), .B(n15779), .Z(n15777) );
  XOR U20259 ( .A(y[1838]), .B(x[1838]), .Z(n15779) );
  XOR U20260 ( .A(y[1837]), .B(x[1837]), .Z(n15780) );
  XOR U20261 ( .A(y[1836]), .B(x[1836]), .Z(n15778) );
  XNOR U20262 ( .A(n15771), .B(n15770), .Z(n15773) );
  XNOR U20263 ( .A(n15767), .B(n15766), .Z(n15770) );
  XOR U20264 ( .A(n15769), .B(n15768), .Z(n15766) );
  XOR U20265 ( .A(y[1835]), .B(x[1835]), .Z(n15768) );
  XOR U20266 ( .A(y[1834]), .B(x[1834]), .Z(n15769) );
  XOR U20267 ( .A(y[1833]), .B(x[1833]), .Z(n15767) );
  XOR U20268 ( .A(n15761), .B(n15760), .Z(n15771) );
  XOR U20269 ( .A(n15763), .B(n15762), .Z(n15760) );
  XOR U20270 ( .A(y[1832]), .B(x[1832]), .Z(n15762) );
  XOR U20271 ( .A(y[1831]), .B(x[1831]), .Z(n15763) );
  XOR U20272 ( .A(y[1830]), .B(x[1830]), .Z(n15761) );
  NAND U20273 ( .A(n15824), .B(n15825), .Z(N28845) );
  NAND U20274 ( .A(n15826), .B(n15827), .Z(n15825) );
  NANDN U20275 ( .A(n15828), .B(n15829), .Z(n15827) );
  NANDN U20276 ( .A(n15829), .B(n15828), .Z(n15824) );
  XOR U20277 ( .A(n15828), .B(n15830), .Z(N28844) );
  XNOR U20278 ( .A(n15826), .B(n15829), .Z(n15830) );
  NAND U20279 ( .A(n15831), .B(n15832), .Z(n15829) );
  NAND U20280 ( .A(n15833), .B(n15834), .Z(n15832) );
  NANDN U20281 ( .A(n15835), .B(n15836), .Z(n15834) );
  NANDN U20282 ( .A(n15836), .B(n15835), .Z(n15831) );
  AND U20283 ( .A(n15837), .B(n15838), .Z(n15826) );
  NAND U20284 ( .A(n15839), .B(n15840), .Z(n15838) );
  OR U20285 ( .A(n15841), .B(n15842), .Z(n15840) );
  NAND U20286 ( .A(n15842), .B(n15841), .Z(n15837) );
  IV U20287 ( .A(n15843), .Z(n15842) );
  AND U20288 ( .A(n15844), .B(n15845), .Z(n15828) );
  NAND U20289 ( .A(n15846), .B(n15847), .Z(n15845) );
  NANDN U20290 ( .A(n15848), .B(n15849), .Z(n15847) );
  NANDN U20291 ( .A(n15849), .B(n15848), .Z(n15844) );
  XOR U20292 ( .A(n15841), .B(n15850), .Z(N28843) );
  XOR U20293 ( .A(n15839), .B(n15843), .Z(n15850) );
  XNOR U20294 ( .A(n15836), .B(n15851), .Z(n15843) );
  XNOR U20295 ( .A(n15833), .B(n15835), .Z(n15851) );
  AND U20296 ( .A(n15852), .B(n15853), .Z(n15835) );
  NANDN U20297 ( .A(n15854), .B(n15855), .Z(n15853) );
  NANDN U20298 ( .A(n15856), .B(n15857), .Z(n15855) );
  IV U20299 ( .A(n15858), .Z(n15857) );
  NAND U20300 ( .A(n15858), .B(n15856), .Z(n15852) );
  AND U20301 ( .A(n15859), .B(n15860), .Z(n15833) );
  NAND U20302 ( .A(n15861), .B(n15862), .Z(n15860) );
  OR U20303 ( .A(n15863), .B(n15864), .Z(n15862) );
  NAND U20304 ( .A(n15864), .B(n15863), .Z(n15859) );
  IV U20305 ( .A(n15865), .Z(n15864) );
  NAND U20306 ( .A(n15866), .B(n15867), .Z(n15836) );
  NANDN U20307 ( .A(n15868), .B(n15869), .Z(n15867) );
  NAND U20308 ( .A(n15870), .B(n15871), .Z(n15869) );
  OR U20309 ( .A(n15871), .B(n15870), .Z(n15866) );
  IV U20310 ( .A(n15872), .Z(n15870) );
  AND U20311 ( .A(n15873), .B(n15874), .Z(n15839) );
  NAND U20312 ( .A(n15875), .B(n15876), .Z(n15874) );
  NANDN U20313 ( .A(n15877), .B(n15878), .Z(n15876) );
  NANDN U20314 ( .A(n15878), .B(n15877), .Z(n15873) );
  XOR U20315 ( .A(n15849), .B(n15879), .Z(n15841) );
  XNOR U20316 ( .A(n15846), .B(n15848), .Z(n15879) );
  AND U20317 ( .A(n15880), .B(n15881), .Z(n15848) );
  NANDN U20318 ( .A(n15882), .B(n15883), .Z(n15881) );
  NANDN U20319 ( .A(n15884), .B(n15885), .Z(n15883) );
  IV U20320 ( .A(n15886), .Z(n15885) );
  NAND U20321 ( .A(n15886), .B(n15884), .Z(n15880) );
  AND U20322 ( .A(n15887), .B(n15888), .Z(n15846) );
  NAND U20323 ( .A(n15889), .B(n15890), .Z(n15888) );
  OR U20324 ( .A(n15891), .B(n15892), .Z(n15890) );
  NAND U20325 ( .A(n15892), .B(n15891), .Z(n15887) );
  IV U20326 ( .A(n15893), .Z(n15892) );
  NAND U20327 ( .A(n15894), .B(n15895), .Z(n15849) );
  NANDN U20328 ( .A(n15896), .B(n15897), .Z(n15895) );
  NAND U20329 ( .A(n15898), .B(n15899), .Z(n15897) );
  OR U20330 ( .A(n15899), .B(n15898), .Z(n15894) );
  IV U20331 ( .A(n15900), .Z(n15898) );
  XOR U20332 ( .A(n15875), .B(n15901), .Z(N28842) );
  XNOR U20333 ( .A(n15878), .B(n15877), .Z(n15901) );
  XNOR U20334 ( .A(n15889), .B(n15902), .Z(n15877) );
  XOR U20335 ( .A(n15893), .B(n15891), .Z(n15902) );
  XOR U20336 ( .A(n15899), .B(n15903), .Z(n15891) );
  XOR U20337 ( .A(n15896), .B(n15900), .Z(n15903) );
  NAND U20338 ( .A(n15904), .B(n15905), .Z(n15900) );
  NAND U20339 ( .A(n15906), .B(n15907), .Z(n15905) );
  NAND U20340 ( .A(n15908), .B(n15909), .Z(n15904) );
  AND U20341 ( .A(n15910), .B(n15911), .Z(n15896) );
  NAND U20342 ( .A(n15912), .B(n15913), .Z(n15911) );
  NAND U20343 ( .A(n15914), .B(n15915), .Z(n15910) );
  NANDN U20344 ( .A(n15916), .B(n15917), .Z(n15899) );
  NANDN U20345 ( .A(n15918), .B(n15919), .Z(n15893) );
  XNOR U20346 ( .A(n15884), .B(n15920), .Z(n15889) );
  XOR U20347 ( .A(n15882), .B(n15886), .Z(n15920) );
  NAND U20348 ( .A(n15921), .B(n15922), .Z(n15886) );
  NAND U20349 ( .A(n15923), .B(n15924), .Z(n15922) );
  NAND U20350 ( .A(n15925), .B(n15926), .Z(n15921) );
  AND U20351 ( .A(n15927), .B(n15928), .Z(n15882) );
  NAND U20352 ( .A(n15929), .B(n15930), .Z(n15928) );
  NAND U20353 ( .A(n15931), .B(n15932), .Z(n15927) );
  AND U20354 ( .A(n15933), .B(n15934), .Z(n15884) );
  NAND U20355 ( .A(n15935), .B(n15936), .Z(n15878) );
  XNOR U20356 ( .A(n15861), .B(n15937), .Z(n15875) );
  XOR U20357 ( .A(n15865), .B(n15863), .Z(n15937) );
  XOR U20358 ( .A(n15871), .B(n15938), .Z(n15863) );
  XOR U20359 ( .A(n15868), .B(n15872), .Z(n15938) );
  NAND U20360 ( .A(n15939), .B(n15940), .Z(n15872) );
  NAND U20361 ( .A(n15941), .B(n15942), .Z(n15940) );
  NAND U20362 ( .A(n15943), .B(n15944), .Z(n15939) );
  AND U20363 ( .A(n15945), .B(n15946), .Z(n15868) );
  NAND U20364 ( .A(n15947), .B(n15948), .Z(n15946) );
  NAND U20365 ( .A(n15949), .B(n15950), .Z(n15945) );
  NANDN U20366 ( .A(n15951), .B(n15952), .Z(n15871) );
  NANDN U20367 ( .A(n15953), .B(n15954), .Z(n15865) );
  XNOR U20368 ( .A(n15856), .B(n15955), .Z(n15861) );
  XOR U20369 ( .A(n15854), .B(n15858), .Z(n15955) );
  NAND U20370 ( .A(n15956), .B(n15957), .Z(n15858) );
  NAND U20371 ( .A(n15958), .B(n15959), .Z(n15957) );
  NAND U20372 ( .A(n15960), .B(n15961), .Z(n15956) );
  AND U20373 ( .A(n15962), .B(n15963), .Z(n15854) );
  NAND U20374 ( .A(n15964), .B(n15965), .Z(n15963) );
  NAND U20375 ( .A(n15966), .B(n15967), .Z(n15962) );
  AND U20376 ( .A(n15968), .B(n15969), .Z(n15856) );
  XOR U20377 ( .A(n15936), .B(n15935), .Z(N28841) );
  XNOR U20378 ( .A(n15954), .B(n15953), .Z(n15935) );
  XNOR U20379 ( .A(n15968), .B(n15969), .Z(n15953) );
  XOR U20380 ( .A(n15965), .B(n15964), .Z(n15969) );
  XOR U20381 ( .A(y[1827]), .B(x[1827]), .Z(n15964) );
  XOR U20382 ( .A(n15967), .B(n15966), .Z(n15965) );
  XOR U20383 ( .A(y[1829]), .B(x[1829]), .Z(n15966) );
  XOR U20384 ( .A(y[1828]), .B(x[1828]), .Z(n15967) );
  XOR U20385 ( .A(n15959), .B(n15958), .Z(n15968) );
  XOR U20386 ( .A(n15961), .B(n15960), .Z(n15958) );
  XOR U20387 ( .A(y[1826]), .B(x[1826]), .Z(n15960) );
  XOR U20388 ( .A(y[1825]), .B(x[1825]), .Z(n15961) );
  XOR U20389 ( .A(y[1824]), .B(x[1824]), .Z(n15959) );
  XNOR U20390 ( .A(n15952), .B(n15951), .Z(n15954) );
  XNOR U20391 ( .A(n15948), .B(n15947), .Z(n15951) );
  XOR U20392 ( .A(n15950), .B(n15949), .Z(n15947) );
  XOR U20393 ( .A(y[1823]), .B(x[1823]), .Z(n15949) );
  XOR U20394 ( .A(y[1822]), .B(x[1822]), .Z(n15950) );
  XOR U20395 ( .A(y[1821]), .B(x[1821]), .Z(n15948) );
  XOR U20396 ( .A(n15942), .B(n15941), .Z(n15952) );
  XOR U20397 ( .A(n15944), .B(n15943), .Z(n15941) );
  XOR U20398 ( .A(y[1820]), .B(x[1820]), .Z(n15943) );
  XOR U20399 ( .A(y[1819]), .B(x[1819]), .Z(n15944) );
  XOR U20400 ( .A(y[1818]), .B(x[1818]), .Z(n15942) );
  XNOR U20401 ( .A(n15919), .B(n15918), .Z(n15936) );
  XNOR U20402 ( .A(n15933), .B(n15934), .Z(n15918) );
  XOR U20403 ( .A(n15930), .B(n15929), .Z(n15934) );
  XOR U20404 ( .A(y[1815]), .B(x[1815]), .Z(n15929) );
  XOR U20405 ( .A(n15932), .B(n15931), .Z(n15930) );
  XOR U20406 ( .A(y[1817]), .B(x[1817]), .Z(n15931) );
  XOR U20407 ( .A(y[1816]), .B(x[1816]), .Z(n15932) );
  XOR U20408 ( .A(n15924), .B(n15923), .Z(n15933) );
  XOR U20409 ( .A(n15926), .B(n15925), .Z(n15923) );
  XOR U20410 ( .A(y[1814]), .B(x[1814]), .Z(n15925) );
  XOR U20411 ( .A(y[1813]), .B(x[1813]), .Z(n15926) );
  XOR U20412 ( .A(y[1812]), .B(x[1812]), .Z(n15924) );
  XNOR U20413 ( .A(n15917), .B(n15916), .Z(n15919) );
  XNOR U20414 ( .A(n15913), .B(n15912), .Z(n15916) );
  XOR U20415 ( .A(n15915), .B(n15914), .Z(n15912) );
  XOR U20416 ( .A(y[1811]), .B(x[1811]), .Z(n15914) );
  XOR U20417 ( .A(y[1810]), .B(x[1810]), .Z(n15915) );
  XOR U20418 ( .A(y[1809]), .B(x[1809]), .Z(n15913) );
  XOR U20419 ( .A(n15907), .B(n15906), .Z(n15917) );
  XOR U20420 ( .A(n15909), .B(n15908), .Z(n15906) );
  XOR U20421 ( .A(y[1808]), .B(x[1808]), .Z(n15908) );
  XOR U20422 ( .A(y[1807]), .B(x[1807]), .Z(n15909) );
  XOR U20423 ( .A(y[1806]), .B(x[1806]), .Z(n15907) );
  NAND U20424 ( .A(n15970), .B(n15971), .Z(N28833) );
  NAND U20425 ( .A(n15972), .B(n15973), .Z(n15971) );
  NANDN U20426 ( .A(n15974), .B(n15975), .Z(n15973) );
  NANDN U20427 ( .A(n15975), .B(n15974), .Z(n15970) );
  XOR U20428 ( .A(n15974), .B(n15976), .Z(N28832) );
  XNOR U20429 ( .A(n15972), .B(n15975), .Z(n15976) );
  NAND U20430 ( .A(n15977), .B(n15978), .Z(n15975) );
  NAND U20431 ( .A(n15979), .B(n15980), .Z(n15978) );
  NANDN U20432 ( .A(n15981), .B(n15982), .Z(n15980) );
  NANDN U20433 ( .A(n15982), .B(n15981), .Z(n15977) );
  AND U20434 ( .A(n15983), .B(n15984), .Z(n15972) );
  NAND U20435 ( .A(n15985), .B(n15986), .Z(n15984) );
  OR U20436 ( .A(n15987), .B(n15988), .Z(n15986) );
  NAND U20437 ( .A(n15988), .B(n15987), .Z(n15983) );
  IV U20438 ( .A(n15989), .Z(n15988) );
  AND U20439 ( .A(n15990), .B(n15991), .Z(n15974) );
  NAND U20440 ( .A(n15992), .B(n15993), .Z(n15991) );
  NANDN U20441 ( .A(n15994), .B(n15995), .Z(n15993) );
  NANDN U20442 ( .A(n15995), .B(n15994), .Z(n15990) );
  XOR U20443 ( .A(n15987), .B(n15996), .Z(N28831) );
  XOR U20444 ( .A(n15985), .B(n15989), .Z(n15996) );
  XNOR U20445 ( .A(n15982), .B(n15997), .Z(n15989) );
  XNOR U20446 ( .A(n15979), .B(n15981), .Z(n15997) );
  AND U20447 ( .A(n15998), .B(n15999), .Z(n15981) );
  NANDN U20448 ( .A(n16000), .B(n16001), .Z(n15999) );
  NANDN U20449 ( .A(n16002), .B(n16003), .Z(n16001) );
  IV U20450 ( .A(n16004), .Z(n16003) );
  NAND U20451 ( .A(n16004), .B(n16002), .Z(n15998) );
  AND U20452 ( .A(n16005), .B(n16006), .Z(n15979) );
  NAND U20453 ( .A(n16007), .B(n16008), .Z(n16006) );
  OR U20454 ( .A(n16009), .B(n16010), .Z(n16008) );
  NAND U20455 ( .A(n16010), .B(n16009), .Z(n16005) );
  IV U20456 ( .A(n16011), .Z(n16010) );
  NAND U20457 ( .A(n16012), .B(n16013), .Z(n15982) );
  NANDN U20458 ( .A(n16014), .B(n16015), .Z(n16013) );
  NAND U20459 ( .A(n16016), .B(n16017), .Z(n16015) );
  OR U20460 ( .A(n16017), .B(n16016), .Z(n16012) );
  IV U20461 ( .A(n16018), .Z(n16016) );
  AND U20462 ( .A(n16019), .B(n16020), .Z(n15985) );
  NAND U20463 ( .A(n16021), .B(n16022), .Z(n16020) );
  NANDN U20464 ( .A(n16023), .B(n16024), .Z(n16022) );
  NANDN U20465 ( .A(n16024), .B(n16023), .Z(n16019) );
  XOR U20466 ( .A(n15995), .B(n16025), .Z(n15987) );
  XNOR U20467 ( .A(n15992), .B(n15994), .Z(n16025) );
  AND U20468 ( .A(n16026), .B(n16027), .Z(n15994) );
  NANDN U20469 ( .A(n16028), .B(n16029), .Z(n16027) );
  NANDN U20470 ( .A(n16030), .B(n16031), .Z(n16029) );
  IV U20471 ( .A(n16032), .Z(n16031) );
  NAND U20472 ( .A(n16032), .B(n16030), .Z(n16026) );
  AND U20473 ( .A(n16033), .B(n16034), .Z(n15992) );
  NAND U20474 ( .A(n16035), .B(n16036), .Z(n16034) );
  OR U20475 ( .A(n16037), .B(n16038), .Z(n16036) );
  NAND U20476 ( .A(n16038), .B(n16037), .Z(n16033) );
  IV U20477 ( .A(n16039), .Z(n16038) );
  NAND U20478 ( .A(n16040), .B(n16041), .Z(n15995) );
  NANDN U20479 ( .A(n16042), .B(n16043), .Z(n16041) );
  NAND U20480 ( .A(n16044), .B(n16045), .Z(n16043) );
  OR U20481 ( .A(n16045), .B(n16044), .Z(n16040) );
  IV U20482 ( .A(n16046), .Z(n16044) );
  XOR U20483 ( .A(n16021), .B(n16047), .Z(N28830) );
  XNOR U20484 ( .A(n16024), .B(n16023), .Z(n16047) );
  XNOR U20485 ( .A(n16035), .B(n16048), .Z(n16023) );
  XOR U20486 ( .A(n16039), .B(n16037), .Z(n16048) );
  XOR U20487 ( .A(n16045), .B(n16049), .Z(n16037) );
  XOR U20488 ( .A(n16042), .B(n16046), .Z(n16049) );
  NAND U20489 ( .A(n16050), .B(n16051), .Z(n16046) );
  NAND U20490 ( .A(n16052), .B(n16053), .Z(n16051) );
  NAND U20491 ( .A(n16054), .B(n16055), .Z(n16050) );
  AND U20492 ( .A(n16056), .B(n16057), .Z(n16042) );
  NAND U20493 ( .A(n16058), .B(n16059), .Z(n16057) );
  NAND U20494 ( .A(n16060), .B(n16061), .Z(n16056) );
  NANDN U20495 ( .A(n16062), .B(n16063), .Z(n16045) );
  NANDN U20496 ( .A(n16064), .B(n16065), .Z(n16039) );
  XNOR U20497 ( .A(n16030), .B(n16066), .Z(n16035) );
  XOR U20498 ( .A(n16028), .B(n16032), .Z(n16066) );
  NAND U20499 ( .A(n16067), .B(n16068), .Z(n16032) );
  NAND U20500 ( .A(n16069), .B(n16070), .Z(n16068) );
  NAND U20501 ( .A(n16071), .B(n16072), .Z(n16067) );
  AND U20502 ( .A(n16073), .B(n16074), .Z(n16028) );
  NAND U20503 ( .A(n16075), .B(n16076), .Z(n16074) );
  NAND U20504 ( .A(n16077), .B(n16078), .Z(n16073) );
  AND U20505 ( .A(n16079), .B(n16080), .Z(n16030) );
  NAND U20506 ( .A(n16081), .B(n16082), .Z(n16024) );
  XNOR U20507 ( .A(n16007), .B(n16083), .Z(n16021) );
  XOR U20508 ( .A(n16011), .B(n16009), .Z(n16083) );
  XOR U20509 ( .A(n16017), .B(n16084), .Z(n16009) );
  XOR U20510 ( .A(n16014), .B(n16018), .Z(n16084) );
  NAND U20511 ( .A(n16085), .B(n16086), .Z(n16018) );
  NAND U20512 ( .A(n16087), .B(n16088), .Z(n16086) );
  NAND U20513 ( .A(n16089), .B(n16090), .Z(n16085) );
  AND U20514 ( .A(n16091), .B(n16092), .Z(n16014) );
  NAND U20515 ( .A(n16093), .B(n16094), .Z(n16092) );
  NAND U20516 ( .A(n16095), .B(n16096), .Z(n16091) );
  NANDN U20517 ( .A(n16097), .B(n16098), .Z(n16017) );
  NANDN U20518 ( .A(n16099), .B(n16100), .Z(n16011) );
  XNOR U20519 ( .A(n16002), .B(n16101), .Z(n16007) );
  XOR U20520 ( .A(n16000), .B(n16004), .Z(n16101) );
  NAND U20521 ( .A(n16102), .B(n16103), .Z(n16004) );
  NAND U20522 ( .A(n16104), .B(n16105), .Z(n16103) );
  NAND U20523 ( .A(n16106), .B(n16107), .Z(n16102) );
  AND U20524 ( .A(n16108), .B(n16109), .Z(n16000) );
  NAND U20525 ( .A(n16110), .B(n16111), .Z(n16109) );
  NAND U20526 ( .A(n16112), .B(n16113), .Z(n16108) );
  AND U20527 ( .A(n16114), .B(n16115), .Z(n16002) );
  XOR U20528 ( .A(n16082), .B(n16081), .Z(N28829) );
  XNOR U20529 ( .A(n16100), .B(n16099), .Z(n16081) );
  XNOR U20530 ( .A(n16114), .B(n16115), .Z(n16099) );
  XOR U20531 ( .A(n16111), .B(n16110), .Z(n16115) );
  XOR U20532 ( .A(y[1803]), .B(x[1803]), .Z(n16110) );
  XOR U20533 ( .A(n16113), .B(n16112), .Z(n16111) );
  XOR U20534 ( .A(y[1805]), .B(x[1805]), .Z(n16112) );
  XOR U20535 ( .A(y[1804]), .B(x[1804]), .Z(n16113) );
  XOR U20536 ( .A(n16105), .B(n16104), .Z(n16114) );
  XOR U20537 ( .A(n16107), .B(n16106), .Z(n16104) );
  XOR U20538 ( .A(y[1802]), .B(x[1802]), .Z(n16106) );
  XOR U20539 ( .A(y[1801]), .B(x[1801]), .Z(n16107) );
  XOR U20540 ( .A(y[1800]), .B(x[1800]), .Z(n16105) );
  XNOR U20541 ( .A(n16098), .B(n16097), .Z(n16100) );
  XNOR U20542 ( .A(n16094), .B(n16093), .Z(n16097) );
  XOR U20543 ( .A(n16096), .B(n16095), .Z(n16093) );
  XOR U20544 ( .A(y[1799]), .B(x[1799]), .Z(n16095) );
  XOR U20545 ( .A(y[1798]), .B(x[1798]), .Z(n16096) );
  XOR U20546 ( .A(y[1797]), .B(x[1797]), .Z(n16094) );
  XOR U20547 ( .A(n16088), .B(n16087), .Z(n16098) );
  XOR U20548 ( .A(n16090), .B(n16089), .Z(n16087) );
  XOR U20549 ( .A(y[1796]), .B(x[1796]), .Z(n16089) );
  XOR U20550 ( .A(y[1795]), .B(x[1795]), .Z(n16090) );
  XOR U20551 ( .A(y[1794]), .B(x[1794]), .Z(n16088) );
  XNOR U20552 ( .A(n16065), .B(n16064), .Z(n16082) );
  XNOR U20553 ( .A(n16079), .B(n16080), .Z(n16064) );
  XOR U20554 ( .A(n16076), .B(n16075), .Z(n16080) );
  XOR U20555 ( .A(y[1791]), .B(x[1791]), .Z(n16075) );
  XOR U20556 ( .A(n16078), .B(n16077), .Z(n16076) );
  XOR U20557 ( .A(y[1793]), .B(x[1793]), .Z(n16077) );
  XOR U20558 ( .A(y[1792]), .B(x[1792]), .Z(n16078) );
  XOR U20559 ( .A(n16070), .B(n16069), .Z(n16079) );
  XOR U20560 ( .A(n16072), .B(n16071), .Z(n16069) );
  XOR U20561 ( .A(y[1790]), .B(x[1790]), .Z(n16071) );
  XOR U20562 ( .A(y[1789]), .B(x[1789]), .Z(n16072) );
  XOR U20563 ( .A(y[1788]), .B(x[1788]), .Z(n16070) );
  XNOR U20564 ( .A(n16063), .B(n16062), .Z(n16065) );
  XNOR U20565 ( .A(n16059), .B(n16058), .Z(n16062) );
  XOR U20566 ( .A(n16061), .B(n16060), .Z(n16058) );
  XOR U20567 ( .A(y[1787]), .B(x[1787]), .Z(n16060) );
  XOR U20568 ( .A(y[1786]), .B(x[1786]), .Z(n16061) );
  XOR U20569 ( .A(y[1785]), .B(x[1785]), .Z(n16059) );
  XOR U20570 ( .A(n16053), .B(n16052), .Z(n16063) );
  XOR U20571 ( .A(n16055), .B(n16054), .Z(n16052) );
  XOR U20572 ( .A(y[1784]), .B(x[1784]), .Z(n16054) );
  XOR U20573 ( .A(y[1783]), .B(x[1783]), .Z(n16055) );
  XOR U20574 ( .A(y[1782]), .B(x[1782]), .Z(n16053) );
  NAND U20575 ( .A(n16116), .B(n16117), .Z(N28821) );
  NAND U20576 ( .A(n16118), .B(n16119), .Z(n16117) );
  NANDN U20577 ( .A(n16120), .B(n16121), .Z(n16119) );
  NANDN U20578 ( .A(n16121), .B(n16120), .Z(n16116) );
  XOR U20579 ( .A(n16120), .B(n16122), .Z(N28820) );
  XNOR U20580 ( .A(n16118), .B(n16121), .Z(n16122) );
  NAND U20581 ( .A(n16123), .B(n16124), .Z(n16121) );
  NAND U20582 ( .A(n16125), .B(n16126), .Z(n16124) );
  NANDN U20583 ( .A(n16127), .B(n16128), .Z(n16126) );
  NANDN U20584 ( .A(n16128), .B(n16127), .Z(n16123) );
  AND U20585 ( .A(n16129), .B(n16130), .Z(n16118) );
  NAND U20586 ( .A(n16131), .B(n16132), .Z(n16130) );
  OR U20587 ( .A(n16133), .B(n16134), .Z(n16132) );
  NAND U20588 ( .A(n16134), .B(n16133), .Z(n16129) );
  IV U20589 ( .A(n16135), .Z(n16134) );
  AND U20590 ( .A(n16136), .B(n16137), .Z(n16120) );
  NAND U20591 ( .A(n16138), .B(n16139), .Z(n16137) );
  NANDN U20592 ( .A(n16140), .B(n16141), .Z(n16139) );
  NANDN U20593 ( .A(n16141), .B(n16140), .Z(n16136) );
  XOR U20594 ( .A(n16133), .B(n16142), .Z(N28819) );
  XOR U20595 ( .A(n16131), .B(n16135), .Z(n16142) );
  XNOR U20596 ( .A(n16128), .B(n16143), .Z(n16135) );
  XNOR U20597 ( .A(n16125), .B(n16127), .Z(n16143) );
  AND U20598 ( .A(n16144), .B(n16145), .Z(n16127) );
  NANDN U20599 ( .A(n16146), .B(n16147), .Z(n16145) );
  NANDN U20600 ( .A(n16148), .B(n16149), .Z(n16147) );
  IV U20601 ( .A(n16150), .Z(n16149) );
  NAND U20602 ( .A(n16150), .B(n16148), .Z(n16144) );
  AND U20603 ( .A(n16151), .B(n16152), .Z(n16125) );
  NAND U20604 ( .A(n16153), .B(n16154), .Z(n16152) );
  OR U20605 ( .A(n16155), .B(n16156), .Z(n16154) );
  NAND U20606 ( .A(n16156), .B(n16155), .Z(n16151) );
  IV U20607 ( .A(n16157), .Z(n16156) );
  NAND U20608 ( .A(n16158), .B(n16159), .Z(n16128) );
  NANDN U20609 ( .A(n16160), .B(n16161), .Z(n16159) );
  NAND U20610 ( .A(n16162), .B(n16163), .Z(n16161) );
  OR U20611 ( .A(n16163), .B(n16162), .Z(n16158) );
  IV U20612 ( .A(n16164), .Z(n16162) );
  AND U20613 ( .A(n16165), .B(n16166), .Z(n16131) );
  NAND U20614 ( .A(n16167), .B(n16168), .Z(n16166) );
  NANDN U20615 ( .A(n16169), .B(n16170), .Z(n16168) );
  NANDN U20616 ( .A(n16170), .B(n16169), .Z(n16165) );
  XOR U20617 ( .A(n16141), .B(n16171), .Z(n16133) );
  XNOR U20618 ( .A(n16138), .B(n16140), .Z(n16171) );
  AND U20619 ( .A(n16172), .B(n16173), .Z(n16140) );
  NANDN U20620 ( .A(n16174), .B(n16175), .Z(n16173) );
  NANDN U20621 ( .A(n16176), .B(n16177), .Z(n16175) );
  IV U20622 ( .A(n16178), .Z(n16177) );
  NAND U20623 ( .A(n16178), .B(n16176), .Z(n16172) );
  AND U20624 ( .A(n16179), .B(n16180), .Z(n16138) );
  NAND U20625 ( .A(n16181), .B(n16182), .Z(n16180) );
  OR U20626 ( .A(n16183), .B(n16184), .Z(n16182) );
  NAND U20627 ( .A(n16184), .B(n16183), .Z(n16179) );
  IV U20628 ( .A(n16185), .Z(n16184) );
  NAND U20629 ( .A(n16186), .B(n16187), .Z(n16141) );
  NANDN U20630 ( .A(n16188), .B(n16189), .Z(n16187) );
  NAND U20631 ( .A(n16190), .B(n16191), .Z(n16189) );
  OR U20632 ( .A(n16191), .B(n16190), .Z(n16186) );
  IV U20633 ( .A(n16192), .Z(n16190) );
  XOR U20634 ( .A(n16167), .B(n16193), .Z(N28818) );
  XNOR U20635 ( .A(n16170), .B(n16169), .Z(n16193) );
  XNOR U20636 ( .A(n16181), .B(n16194), .Z(n16169) );
  XOR U20637 ( .A(n16185), .B(n16183), .Z(n16194) );
  XOR U20638 ( .A(n16191), .B(n16195), .Z(n16183) );
  XOR U20639 ( .A(n16188), .B(n16192), .Z(n16195) );
  NAND U20640 ( .A(n16196), .B(n16197), .Z(n16192) );
  NAND U20641 ( .A(n16198), .B(n16199), .Z(n16197) );
  NAND U20642 ( .A(n16200), .B(n16201), .Z(n16196) );
  AND U20643 ( .A(n16202), .B(n16203), .Z(n16188) );
  NAND U20644 ( .A(n16204), .B(n16205), .Z(n16203) );
  NAND U20645 ( .A(n16206), .B(n16207), .Z(n16202) );
  NANDN U20646 ( .A(n16208), .B(n16209), .Z(n16191) );
  NANDN U20647 ( .A(n16210), .B(n16211), .Z(n16185) );
  XNOR U20648 ( .A(n16176), .B(n16212), .Z(n16181) );
  XOR U20649 ( .A(n16174), .B(n16178), .Z(n16212) );
  NAND U20650 ( .A(n16213), .B(n16214), .Z(n16178) );
  NAND U20651 ( .A(n16215), .B(n16216), .Z(n16214) );
  NAND U20652 ( .A(n16217), .B(n16218), .Z(n16213) );
  AND U20653 ( .A(n16219), .B(n16220), .Z(n16174) );
  NAND U20654 ( .A(n16221), .B(n16222), .Z(n16220) );
  NAND U20655 ( .A(n16223), .B(n16224), .Z(n16219) );
  AND U20656 ( .A(n16225), .B(n16226), .Z(n16176) );
  NAND U20657 ( .A(n16227), .B(n16228), .Z(n16170) );
  XNOR U20658 ( .A(n16153), .B(n16229), .Z(n16167) );
  XOR U20659 ( .A(n16157), .B(n16155), .Z(n16229) );
  XOR U20660 ( .A(n16163), .B(n16230), .Z(n16155) );
  XOR U20661 ( .A(n16160), .B(n16164), .Z(n16230) );
  NAND U20662 ( .A(n16231), .B(n16232), .Z(n16164) );
  NAND U20663 ( .A(n16233), .B(n16234), .Z(n16232) );
  NAND U20664 ( .A(n16235), .B(n16236), .Z(n16231) );
  AND U20665 ( .A(n16237), .B(n16238), .Z(n16160) );
  NAND U20666 ( .A(n16239), .B(n16240), .Z(n16238) );
  NAND U20667 ( .A(n16241), .B(n16242), .Z(n16237) );
  NANDN U20668 ( .A(n16243), .B(n16244), .Z(n16163) );
  NANDN U20669 ( .A(n16245), .B(n16246), .Z(n16157) );
  XNOR U20670 ( .A(n16148), .B(n16247), .Z(n16153) );
  XOR U20671 ( .A(n16146), .B(n16150), .Z(n16247) );
  NAND U20672 ( .A(n16248), .B(n16249), .Z(n16150) );
  NAND U20673 ( .A(n16250), .B(n16251), .Z(n16249) );
  NAND U20674 ( .A(n16252), .B(n16253), .Z(n16248) );
  AND U20675 ( .A(n16254), .B(n16255), .Z(n16146) );
  NAND U20676 ( .A(n16256), .B(n16257), .Z(n16255) );
  NAND U20677 ( .A(n16258), .B(n16259), .Z(n16254) );
  AND U20678 ( .A(n16260), .B(n16261), .Z(n16148) );
  XOR U20679 ( .A(n16228), .B(n16227), .Z(N28817) );
  XNOR U20680 ( .A(n16246), .B(n16245), .Z(n16227) );
  XNOR U20681 ( .A(n16260), .B(n16261), .Z(n16245) );
  XOR U20682 ( .A(n16257), .B(n16256), .Z(n16261) );
  XOR U20683 ( .A(y[1779]), .B(x[1779]), .Z(n16256) );
  XOR U20684 ( .A(n16259), .B(n16258), .Z(n16257) );
  XOR U20685 ( .A(y[1781]), .B(x[1781]), .Z(n16258) );
  XOR U20686 ( .A(y[1780]), .B(x[1780]), .Z(n16259) );
  XOR U20687 ( .A(n16251), .B(n16250), .Z(n16260) );
  XOR U20688 ( .A(n16253), .B(n16252), .Z(n16250) );
  XOR U20689 ( .A(y[1778]), .B(x[1778]), .Z(n16252) );
  XOR U20690 ( .A(y[1777]), .B(x[1777]), .Z(n16253) );
  XOR U20691 ( .A(y[1776]), .B(x[1776]), .Z(n16251) );
  XNOR U20692 ( .A(n16244), .B(n16243), .Z(n16246) );
  XNOR U20693 ( .A(n16240), .B(n16239), .Z(n16243) );
  XOR U20694 ( .A(n16242), .B(n16241), .Z(n16239) );
  XOR U20695 ( .A(y[1775]), .B(x[1775]), .Z(n16241) );
  XOR U20696 ( .A(y[1774]), .B(x[1774]), .Z(n16242) );
  XOR U20697 ( .A(y[1773]), .B(x[1773]), .Z(n16240) );
  XOR U20698 ( .A(n16234), .B(n16233), .Z(n16244) );
  XOR U20699 ( .A(n16236), .B(n16235), .Z(n16233) );
  XOR U20700 ( .A(y[1772]), .B(x[1772]), .Z(n16235) );
  XOR U20701 ( .A(y[1771]), .B(x[1771]), .Z(n16236) );
  XOR U20702 ( .A(y[1770]), .B(x[1770]), .Z(n16234) );
  XNOR U20703 ( .A(n16211), .B(n16210), .Z(n16228) );
  XNOR U20704 ( .A(n16225), .B(n16226), .Z(n16210) );
  XOR U20705 ( .A(n16222), .B(n16221), .Z(n16226) );
  XOR U20706 ( .A(y[1767]), .B(x[1767]), .Z(n16221) );
  XOR U20707 ( .A(n16224), .B(n16223), .Z(n16222) );
  XOR U20708 ( .A(y[1769]), .B(x[1769]), .Z(n16223) );
  XOR U20709 ( .A(y[1768]), .B(x[1768]), .Z(n16224) );
  XOR U20710 ( .A(n16216), .B(n16215), .Z(n16225) );
  XOR U20711 ( .A(n16218), .B(n16217), .Z(n16215) );
  XOR U20712 ( .A(y[1766]), .B(x[1766]), .Z(n16217) );
  XOR U20713 ( .A(y[1765]), .B(x[1765]), .Z(n16218) );
  XOR U20714 ( .A(y[1764]), .B(x[1764]), .Z(n16216) );
  XNOR U20715 ( .A(n16209), .B(n16208), .Z(n16211) );
  XNOR U20716 ( .A(n16205), .B(n16204), .Z(n16208) );
  XOR U20717 ( .A(n16207), .B(n16206), .Z(n16204) );
  XOR U20718 ( .A(y[1763]), .B(x[1763]), .Z(n16206) );
  XOR U20719 ( .A(y[1762]), .B(x[1762]), .Z(n16207) );
  XOR U20720 ( .A(y[1761]), .B(x[1761]), .Z(n16205) );
  XOR U20721 ( .A(n16199), .B(n16198), .Z(n16209) );
  XOR U20722 ( .A(n16201), .B(n16200), .Z(n16198) );
  XOR U20723 ( .A(y[1760]), .B(x[1760]), .Z(n16200) );
  XOR U20724 ( .A(y[1759]), .B(x[1759]), .Z(n16201) );
  XOR U20725 ( .A(y[1758]), .B(x[1758]), .Z(n16199) );
  NAND U20726 ( .A(n16262), .B(n16263), .Z(N28809) );
  NAND U20727 ( .A(n16264), .B(n16265), .Z(n16263) );
  NANDN U20728 ( .A(n16266), .B(n16267), .Z(n16265) );
  NANDN U20729 ( .A(n16267), .B(n16266), .Z(n16262) );
  XOR U20730 ( .A(n16266), .B(n16268), .Z(N28808) );
  XNOR U20731 ( .A(n16264), .B(n16267), .Z(n16268) );
  NAND U20732 ( .A(n16269), .B(n16270), .Z(n16267) );
  NAND U20733 ( .A(n16271), .B(n16272), .Z(n16270) );
  NANDN U20734 ( .A(n16273), .B(n16274), .Z(n16272) );
  NANDN U20735 ( .A(n16274), .B(n16273), .Z(n16269) );
  AND U20736 ( .A(n16275), .B(n16276), .Z(n16264) );
  NAND U20737 ( .A(n16277), .B(n16278), .Z(n16276) );
  OR U20738 ( .A(n16279), .B(n16280), .Z(n16278) );
  NAND U20739 ( .A(n16280), .B(n16279), .Z(n16275) );
  IV U20740 ( .A(n16281), .Z(n16280) );
  AND U20741 ( .A(n16282), .B(n16283), .Z(n16266) );
  NAND U20742 ( .A(n16284), .B(n16285), .Z(n16283) );
  NANDN U20743 ( .A(n16286), .B(n16287), .Z(n16285) );
  NANDN U20744 ( .A(n16287), .B(n16286), .Z(n16282) );
  XOR U20745 ( .A(n16279), .B(n16288), .Z(N28807) );
  XOR U20746 ( .A(n16277), .B(n16281), .Z(n16288) );
  XNOR U20747 ( .A(n16274), .B(n16289), .Z(n16281) );
  XNOR U20748 ( .A(n16271), .B(n16273), .Z(n16289) );
  AND U20749 ( .A(n16290), .B(n16291), .Z(n16273) );
  NANDN U20750 ( .A(n16292), .B(n16293), .Z(n16291) );
  NANDN U20751 ( .A(n16294), .B(n16295), .Z(n16293) );
  IV U20752 ( .A(n16296), .Z(n16295) );
  NAND U20753 ( .A(n16296), .B(n16294), .Z(n16290) );
  AND U20754 ( .A(n16297), .B(n16298), .Z(n16271) );
  NAND U20755 ( .A(n16299), .B(n16300), .Z(n16298) );
  OR U20756 ( .A(n16301), .B(n16302), .Z(n16300) );
  NAND U20757 ( .A(n16302), .B(n16301), .Z(n16297) );
  IV U20758 ( .A(n16303), .Z(n16302) );
  NAND U20759 ( .A(n16304), .B(n16305), .Z(n16274) );
  NANDN U20760 ( .A(n16306), .B(n16307), .Z(n16305) );
  NAND U20761 ( .A(n16308), .B(n16309), .Z(n16307) );
  OR U20762 ( .A(n16309), .B(n16308), .Z(n16304) );
  IV U20763 ( .A(n16310), .Z(n16308) );
  AND U20764 ( .A(n16311), .B(n16312), .Z(n16277) );
  NAND U20765 ( .A(n16313), .B(n16314), .Z(n16312) );
  NANDN U20766 ( .A(n16315), .B(n16316), .Z(n16314) );
  NANDN U20767 ( .A(n16316), .B(n16315), .Z(n16311) );
  XOR U20768 ( .A(n16287), .B(n16317), .Z(n16279) );
  XNOR U20769 ( .A(n16284), .B(n16286), .Z(n16317) );
  AND U20770 ( .A(n16318), .B(n16319), .Z(n16286) );
  NANDN U20771 ( .A(n16320), .B(n16321), .Z(n16319) );
  NANDN U20772 ( .A(n16322), .B(n16323), .Z(n16321) );
  IV U20773 ( .A(n16324), .Z(n16323) );
  NAND U20774 ( .A(n16324), .B(n16322), .Z(n16318) );
  AND U20775 ( .A(n16325), .B(n16326), .Z(n16284) );
  NAND U20776 ( .A(n16327), .B(n16328), .Z(n16326) );
  OR U20777 ( .A(n16329), .B(n16330), .Z(n16328) );
  NAND U20778 ( .A(n16330), .B(n16329), .Z(n16325) );
  IV U20779 ( .A(n16331), .Z(n16330) );
  NAND U20780 ( .A(n16332), .B(n16333), .Z(n16287) );
  NANDN U20781 ( .A(n16334), .B(n16335), .Z(n16333) );
  NAND U20782 ( .A(n16336), .B(n16337), .Z(n16335) );
  OR U20783 ( .A(n16337), .B(n16336), .Z(n16332) );
  IV U20784 ( .A(n16338), .Z(n16336) );
  XOR U20785 ( .A(n16313), .B(n16339), .Z(N28806) );
  XNOR U20786 ( .A(n16316), .B(n16315), .Z(n16339) );
  XNOR U20787 ( .A(n16327), .B(n16340), .Z(n16315) );
  XOR U20788 ( .A(n16331), .B(n16329), .Z(n16340) );
  XOR U20789 ( .A(n16337), .B(n16341), .Z(n16329) );
  XOR U20790 ( .A(n16334), .B(n16338), .Z(n16341) );
  NAND U20791 ( .A(n16342), .B(n16343), .Z(n16338) );
  NAND U20792 ( .A(n16344), .B(n16345), .Z(n16343) );
  NAND U20793 ( .A(n16346), .B(n16347), .Z(n16342) );
  AND U20794 ( .A(n16348), .B(n16349), .Z(n16334) );
  NAND U20795 ( .A(n16350), .B(n16351), .Z(n16349) );
  NAND U20796 ( .A(n16352), .B(n16353), .Z(n16348) );
  NANDN U20797 ( .A(n16354), .B(n16355), .Z(n16337) );
  NANDN U20798 ( .A(n16356), .B(n16357), .Z(n16331) );
  XNOR U20799 ( .A(n16322), .B(n16358), .Z(n16327) );
  XOR U20800 ( .A(n16320), .B(n16324), .Z(n16358) );
  NAND U20801 ( .A(n16359), .B(n16360), .Z(n16324) );
  NAND U20802 ( .A(n16361), .B(n16362), .Z(n16360) );
  NAND U20803 ( .A(n16363), .B(n16364), .Z(n16359) );
  AND U20804 ( .A(n16365), .B(n16366), .Z(n16320) );
  NAND U20805 ( .A(n16367), .B(n16368), .Z(n16366) );
  NAND U20806 ( .A(n16369), .B(n16370), .Z(n16365) );
  AND U20807 ( .A(n16371), .B(n16372), .Z(n16322) );
  NAND U20808 ( .A(n16373), .B(n16374), .Z(n16316) );
  XNOR U20809 ( .A(n16299), .B(n16375), .Z(n16313) );
  XOR U20810 ( .A(n16303), .B(n16301), .Z(n16375) );
  XOR U20811 ( .A(n16309), .B(n16376), .Z(n16301) );
  XOR U20812 ( .A(n16306), .B(n16310), .Z(n16376) );
  NAND U20813 ( .A(n16377), .B(n16378), .Z(n16310) );
  NAND U20814 ( .A(n16379), .B(n16380), .Z(n16378) );
  NAND U20815 ( .A(n16381), .B(n16382), .Z(n16377) );
  AND U20816 ( .A(n16383), .B(n16384), .Z(n16306) );
  NAND U20817 ( .A(n16385), .B(n16386), .Z(n16384) );
  NAND U20818 ( .A(n16387), .B(n16388), .Z(n16383) );
  NANDN U20819 ( .A(n16389), .B(n16390), .Z(n16309) );
  NANDN U20820 ( .A(n16391), .B(n16392), .Z(n16303) );
  XNOR U20821 ( .A(n16294), .B(n16393), .Z(n16299) );
  XOR U20822 ( .A(n16292), .B(n16296), .Z(n16393) );
  NAND U20823 ( .A(n16394), .B(n16395), .Z(n16296) );
  NAND U20824 ( .A(n16396), .B(n16397), .Z(n16395) );
  NAND U20825 ( .A(n16398), .B(n16399), .Z(n16394) );
  AND U20826 ( .A(n16400), .B(n16401), .Z(n16292) );
  NAND U20827 ( .A(n16402), .B(n16403), .Z(n16401) );
  NAND U20828 ( .A(n16404), .B(n16405), .Z(n16400) );
  AND U20829 ( .A(n16406), .B(n16407), .Z(n16294) );
  XOR U20830 ( .A(n16374), .B(n16373), .Z(N28805) );
  XNOR U20831 ( .A(n16392), .B(n16391), .Z(n16373) );
  XNOR U20832 ( .A(n16406), .B(n16407), .Z(n16391) );
  XOR U20833 ( .A(n16403), .B(n16402), .Z(n16407) );
  XOR U20834 ( .A(y[1755]), .B(x[1755]), .Z(n16402) );
  XOR U20835 ( .A(n16405), .B(n16404), .Z(n16403) );
  XOR U20836 ( .A(y[1757]), .B(x[1757]), .Z(n16404) );
  XOR U20837 ( .A(y[1756]), .B(x[1756]), .Z(n16405) );
  XOR U20838 ( .A(n16397), .B(n16396), .Z(n16406) );
  XOR U20839 ( .A(n16399), .B(n16398), .Z(n16396) );
  XOR U20840 ( .A(y[1754]), .B(x[1754]), .Z(n16398) );
  XOR U20841 ( .A(y[1753]), .B(x[1753]), .Z(n16399) );
  XOR U20842 ( .A(y[1752]), .B(x[1752]), .Z(n16397) );
  XNOR U20843 ( .A(n16390), .B(n16389), .Z(n16392) );
  XNOR U20844 ( .A(n16386), .B(n16385), .Z(n16389) );
  XOR U20845 ( .A(n16388), .B(n16387), .Z(n16385) );
  XOR U20846 ( .A(y[1751]), .B(x[1751]), .Z(n16387) );
  XOR U20847 ( .A(y[1750]), .B(x[1750]), .Z(n16388) );
  XOR U20848 ( .A(y[1749]), .B(x[1749]), .Z(n16386) );
  XOR U20849 ( .A(n16380), .B(n16379), .Z(n16390) );
  XOR U20850 ( .A(n16382), .B(n16381), .Z(n16379) );
  XOR U20851 ( .A(y[1748]), .B(x[1748]), .Z(n16381) );
  XOR U20852 ( .A(y[1747]), .B(x[1747]), .Z(n16382) );
  XOR U20853 ( .A(y[1746]), .B(x[1746]), .Z(n16380) );
  XNOR U20854 ( .A(n16357), .B(n16356), .Z(n16374) );
  XNOR U20855 ( .A(n16371), .B(n16372), .Z(n16356) );
  XOR U20856 ( .A(n16368), .B(n16367), .Z(n16372) );
  XOR U20857 ( .A(y[1743]), .B(x[1743]), .Z(n16367) );
  XOR U20858 ( .A(n16370), .B(n16369), .Z(n16368) );
  XOR U20859 ( .A(y[1745]), .B(x[1745]), .Z(n16369) );
  XOR U20860 ( .A(y[1744]), .B(x[1744]), .Z(n16370) );
  XOR U20861 ( .A(n16362), .B(n16361), .Z(n16371) );
  XOR U20862 ( .A(n16364), .B(n16363), .Z(n16361) );
  XOR U20863 ( .A(y[1742]), .B(x[1742]), .Z(n16363) );
  XOR U20864 ( .A(y[1741]), .B(x[1741]), .Z(n16364) );
  XOR U20865 ( .A(y[1740]), .B(x[1740]), .Z(n16362) );
  XNOR U20866 ( .A(n16355), .B(n16354), .Z(n16357) );
  XNOR U20867 ( .A(n16351), .B(n16350), .Z(n16354) );
  XOR U20868 ( .A(n16353), .B(n16352), .Z(n16350) );
  XOR U20869 ( .A(y[1739]), .B(x[1739]), .Z(n16352) );
  XOR U20870 ( .A(y[1738]), .B(x[1738]), .Z(n16353) );
  XOR U20871 ( .A(y[1737]), .B(x[1737]), .Z(n16351) );
  XOR U20872 ( .A(n16345), .B(n16344), .Z(n16355) );
  XOR U20873 ( .A(n16347), .B(n16346), .Z(n16344) );
  XOR U20874 ( .A(y[1736]), .B(x[1736]), .Z(n16346) );
  XOR U20875 ( .A(y[1735]), .B(x[1735]), .Z(n16347) );
  XOR U20876 ( .A(y[1734]), .B(x[1734]), .Z(n16345) );
  NAND U20877 ( .A(n16408), .B(n16409), .Z(N28797) );
  NAND U20878 ( .A(n16410), .B(n16411), .Z(n16409) );
  NANDN U20879 ( .A(n16412), .B(n16413), .Z(n16411) );
  NANDN U20880 ( .A(n16413), .B(n16412), .Z(n16408) );
  XOR U20881 ( .A(n16412), .B(n16414), .Z(N28796) );
  XNOR U20882 ( .A(n16410), .B(n16413), .Z(n16414) );
  NAND U20883 ( .A(n16415), .B(n16416), .Z(n16413) );
  NAND U20884 ( .A(n16417), .B(n16418), .Z(n16416) );
  NANDN U20885 ( .A(n16419), .B(n16420), .Z(n16418) );
  NANDN U20886 ( .A(n16420), .B(n16419), .Z(n16415) );
  AND U20887 ( .A(n16421), .B(n16422), .Z(n16410) );
  NAND U20888 ( .A(n16423), .B(n16424), .Z(n16422) );
  OR U20889 ( .A(n16425), .B(n16426), .Z(n16424) );
  NAND U20890 ( .A(n16426), .B(n16425), .Z(n16421) );
  IV U20891 ( .A(n16427), .Z(n16426) );
  AND U20892 ( .A(n16428), .B(n16429), .Z(n16412) );
  NAND U20893 ( .A(n16430), .B(n16431), .Z(n16429) );
  NANDN U20894 ( .A(n16432), .B(n16433), .Z(n16431) );
  NANDN U20895 ( .A(n16433), .B(n16432), .Z(n16428) );
  XOR U20896 ( .A(n16425), .B(n16434), .Z(N28795) );
  XOR U20897 ( .A(n16423), .B(n16427), .Z(n16434) );
  XNOR U20898 ( .A(n16420), .B(n16435), .Z(n16427) );
  XNOR U20899 ( .A(n16417), .B(n16419), .Z(n16435) );
  AND U20900 ( .A(n16436), .B(n16437), .Z(n16419) );
  NANDN U20901 ( .A(n16438), .B(n16439), .Z(n16437) );
  NANDN U20902 ( .A(n16440), .B(n16441), .Z(n16439) );
  IV U20903 ( .A(n16442), .Z(n16441) );
  NAND U20904 ( .A(n16442), .B(n16440), .Z(n16436) );
  AND U20905 ( .A(n16443), .B(n16444), .Z(n16417) );
  NAND U20906 ( .A(n16445), .B(n16446), .Z(n16444) );
  OR U20907 ( .A(n16447), .B(n16448), .Z(n16446) );
  NAND U20908 ( .A(n16448), .B(n16447), .Z(n16443) );
  IV U20909 ( .A(n16449), .Z(n16448) );
  NAND U20910 ( .A(n16450), .B(n16451), .Z(n16420) );
  NANDN U20911 ( .A(n16452), .B(n16453), .Z(n16451) );
  NAND U20912 ( .A(n16454), .B(n16455), .Z(n16453) );
  OR U20913 ( .A(n16455), .B(n16454), .Z(n16450) );
  IV U20914 ( .A(n16456), .Z(n16454) );
  AND U20915 ( .A(n16457), .B(n16458), .Z(n16423) );
  NAND U20916 ( .A(n16459), .B(n16460), .Z(n16458) );
  NANDN U20917 ( .A(n16461), .B(n16462), .Z(n16460) );
  NANDN U20918 ( .A(n16462), .B(n16461), .Z(n16457) );
  XOR U20919 ( .A(n16433), .B(n16463), .Z(n16425) );
  XNOR U20920 ( .A(n16430), .B(n16432), .Z(n16463) );
  AND U20921 ( .A(n16464), .B(n16465), .Z(n16432) );
  NANDN U20922 ( .A(n16466), .B(n16467), .Z(n16465) );
  NANDN U20923 ( .A(n16468), .B(n16469), .Z(n16467) );
  IV U20924 ( .A(n16470), .Z(n16469) );
  NAND U20925 ( .A(n16470), .B(n16468), .Z(n16464) );
  AND U20926 ( .A(n16471), .B(n16472), .Z(n16430) );
  NAND U20927 ( .A(n16473), .B(n16474), .Z(n16472) );
  OR U20928 ( .A(n16475), .B(n16476), .Z(n16474) );
  NAND U20929 ( .A(n16476), .B(n16475), .Z(n16471) );
  IV U20930 ( .A(n16477), .Z(n16476) );
  NAND U20931 ( .A(n16478), .B(n16479), .Z(n16433) );
  NANDN U20932 ( .A(n16480), .B(n16481), .Z(n16479) );
  NAND U20933 ( .A(n16482), .B(n16483), .Z(n16481) );
  OR U20934 ( .A(n16483), .B(n16482), .Z(n16478) );
  IV U20935 ( .A(n16484), .Z(n16482) );
  XOR U20936 ( .A(n16459), .B(n16485), .Z(N28794) );
  XNOR U20937 ( .A(n16462), .B(n16461), .Z(n16485) );
  XNOR U20938 ( .A(n16473), .B(n16486), .Z(n16461) );
  XOR U20939 ( .A(n16477), .B(n16475), .Z(n16486) );
  XOR U20940 ( .A(n16483), .B(n16487), .Z(n16475) );
  XOR U20941 ( .A(n16480), .B(n16484), .Z(n16487) );
  NAND U20942 ( .A(n16488), .B(n16489), .Z(n16484) );
  NAND U20943 ( .A(n16490), .B(n16491), .Z(n16489) );
  NAND U20944 ( .A(n16492), .B(n16493), .Z(n16488) );
  AND U20945 ( .A(n16494), .B(n16495), .Z(n16480) );
  NAND U20946 ( .A(n16496), .B(n16497), .Z(n16495) );
  NAND U20947 ( .A(n16498), .B(n16499), .Z(n16494) );
  NANDN U20948 ( .A(n16500), .B(n16501), .Z(n16483) );
  NANDN U20949 ( .A(n16502), .B(n16503), .Z(n16477) );
  XNOR U20950 ( .A(n16468), .B(n16504), .Z(n16473) );
  XOR U20951 ( .A(n16466), .B(n16470), .Z(n16504) );
  NAND U20952 ( .A(n16505), .B(n16506), .Z(n16470) );
  NAND U20953 ( .A(n16507), .B(n16508), .Z(n16506) );
  NAND U20954 ( .A(n16509), .B(n16510), .Z(n16505) );
  AND U20955 ( .A(n16511), .B(n16512), .Z(n16466) );
  NAND U20956 ( .A(n16513), .B(n16514), .Z(n16512) );
  NAND U20957 ( .A(n16515), .B(n16516), .Z(n16511) );
  AND U20958 ( .A(n16517), .B(n16518), .Z(n16468) );
  NAND U20959 ( .A(n16519), .B(n16520), .Z(n16462) );
  XNOR U20960 ( .A(n16445), .B(n16521), .Z(n16459) );
  XOR U20961 ( .A(n16449), .B(n16447), .Z(n16521) );
  XOR U20962 ( .A(n16455), .B(n16522), .Z(n16447) );
  XOR U20963 ( .A(n16452), .B(n16456), .Z(n16522) );
  NAND U20964 ( .A(n16523), .B(n16524), .Z(n16456) );
  NAND U20965 ( .A(n16525), .B(n16526), .Z(n16524) );
  NAND U20966 ( .A(n16527), .B(n16528), .Z(n16523) );
  AND U20967 ( .A(n16529), .B(n16530), .Z(n16452) );
  NAND U20968 ( .A(n16531), .B(n16532), .Z(n16530) );
  NAND U20969 ( .A(n16533), .B(n16534), .Z(n16529) );
  NANDN U20970 ( .A(n16535), .B(n16536), .Z(n16455) );
  NANDN U20971 ( .A(n16537), .B(n16538), .Z(n16449) );
  XNOR U20972 ( .A(n16440), .B(n16539), .Z(n16445) );
  XOR U20973 ( .A(n16438), .B(n16442), .Z(n16539) );
  NAND U20974 ( .A(n16540), .B(n16541), .Z(n16442) );
  NAND U20975 ( .A(n16542), .B(n16543), .Z(n16541) );
  NAND U20976 ( .A(n16544), .B(n16545), .Z(n16540) );
  AND U20977 ( .A(n16546), .B(n16547), .Z(n16438) );
  NAND U20978 ( .A(n16548), .B(n16549), .Z(n16547) );
  NAND U20979 ( .A(n16550), .B(n16551), .Z(n16546) );
  AND U20980 ( .A(n16552), .B(n16553), .Z(n16440) );
  XOR U20981 ( .A(n16520), .B(n16519), .Z(N28793) );
  XNOR U20982 ( .A(n16538), .B(n16537), .Z(n16519) );
  XNOR U20983 ( .A(n16552), .B(n16553), .Z(n16537) );
  XOR U20984 ( .A(n16549), .B(n16548), .Z(n16553) );
  XOR U20985 ( .A(y[1731]), .B(x[1731]), .Z(n16548) );
  XOR U20986 ( .A(n16551), .B(n16550), .Z(n16549) );
  XOR U20987 ( .A(y[1733]), .B(x[1733]), .Z(n16550) );
  XOR U20988 ( .A(y[1732]), .B(x[1732]), .Z(n16551) );
  XOR U20989 ( .A(n16543), .B(n16542), .Z(n16552) );
  XOR U20990 ( .A(n16545), .B(n16544), .Z(n16542) );
  XOR U20991 ( .A(y[1730]), .B(x[1730]), .Z(n16544) );
  XOR U20992 ( .A(y[1729]), .B(x[1729]), .Z(n16545) );
  XOR U20993 ( .A(y[1728]), .B(x[1728]), .Z(n16543) );
  XNOR U20994 ( .A(n16536), .B(n16535), .Z(n16538) );
  XNOR U20995 ( .A(n16532), .B(n16531), .Z(n16535) );
  XOR U20996 ( .A(n16534), .B(n16533), .Z(n16531) );
  XOR U20997 ( .A(y[1727]), .B(x[1727]), .Z(n16533) );
  XOR U20998 ( .A(y[1726]), .B(x[1726]), .Z(n16534) );
  XOR U20999 ( .A(y[1725]), .B(x[1725]), .Z(n16532) );
  XOR U21000 ( .A(n16526), .B(n16525), .Z(n16536) );
  XOR U21001 ( .A(n16528), .B(n16527), .Z(n16525) );
  XOR U21002 ( .A(y[1724]), .B(x[1724]), .Z(n16527) );
  XOR U21003 ( .A(y[1723]), .B(x[1723]), .Z(n16528) );
  XOR U21004 ( .A(y[1722]), .B(x[1722]), .Z(n16526) );
  XNOR U21005 ( .A(n16503), .B(n16502), .Z(n16520) );
  XNOR U21006 ( .A(n16517), .B(n16518), .Z(n16502) );
  XOR U21007 ( .A(n16514), .B(n16513), .Z(n16518) );
  XOR U21008 ( .A(y[1719]), .B(x[1719]), .Z(n16513) );
  XOR U21009 ( .A(n16516), .B(n16515), .Z(n16514) );
  XOR U21010 ( .A(y[1721]), .B(x[1721]), .Z(n16515) );
  XOR U21011 ( .A(y[1720]), .B(x[1720]), .Z(n16516) );
  XOR U21012 ( .A(n16508), .B(n16507), .Z(n16517) );
  XOR U21013 ( .A(n16510), .B(n16509), .Z(n16507) );
  XOR U21014 ( .A(y[1718]), .B(x[1718]), .Z(n16509) );
  XOR U21015 ( .A(y[1717]), .B(x[1717]), .Z(n16510) );
  XOR U21016 ( .A(y[1716]), .B(x[1716]), .Z(n16508) );
  XNOR U21017 ( .A(n16501), .B(n16500), .Z(n16503) );
  XNOR U21018 ( .A(n16497), .B(n16496), .Z(n16500) );
  XOR U21019 ( .A(n16499), .B(n16498), .Z(n16496) );
  XOR U21020 ( .A(y[1715]), .B(x[1715]), .Z(n16498) );
  XOR U21021 ( .A(y[1714]), .B(x[1714]), .Z(n16499) );
  XOR U21022 ( .A(y[1713]), .B(x[1713]), .Z(n16497) );
  XOR U21023 ( .A(n16491), .B(n16490), .Z(n16501) );
  XOR U21024 ( .A(n16493), .B(n16492), .Z(n16490) );
  XOR U21025 ( .A(y[1712]), .B(x[1712]), .Z(n16492) );
  XOR U21026 ( .A(y[1711]), .B(x[1711]), .Z(n16493) );
  XOR U21027 ( .A(y[1710]), .B(x[1710]), .Z(n16491) );
  NAND U21028 ( .A(n16554), .B(n16555), .Z(N28785) );
  NAND U21029 ( .A(n16556), .B(n16557), .Z(n16555) );
  NANDN U21030 ( .A(n16558), .B(n16559), .Z(n16557) );
  NANDN U21031 ( .A(n16559), .B(n16558), .Z(n16554) );
  XOR U21032 ( .A(n16558), .B(n16560), .Z(N28784) );
  XNOR U21033 ( .A(n16556), .B(n16559), .Z(n16560) );
  NAND U21034 ( .A(n16561), .B(n16562), .Z(n16559) );
  NAND U21035 ( .A(n16563), .B(n16564), .Z(n16562) );
  NANDN U21036 ( .A(n16565), .B(n16566), .Z(n16564) );
  NANDN U21037 ( .A(n16566), .B(n16565), .Z(n16561) );
  AND U21038 ( .A(n16567), .B(n16568), .Z(n16556) );
  NAND U21039 ( .A(n16569), .B(n16570), .Z(n16568) );
  OR U21040 ( .A(n16571), .B(n16572), .Z(n16570) );
  NAND U21041 ( .A(n16572), .B(n16571), .Z(n16567) );
  IV U21042 ( .A(n16573), .Z(n16572) );
  AND U21043 ( .A(n16574), .B(n16575), .Z(n16558) );
  NAND U21044 ( .A(n16576), .B(n16577), .Z(n16575) );
  NANDN U21045 ( .A(n16578), .B(n16579), .Z(n16577) );
  NANDN U21046 ( .A(n16579), .B(n16578), .Z(n16574) );
  XOR U21047 ( .A(n16571), .B(n16580), .Z(N28783) );
  XOR U21048 ( .A(n16569), .B(n16573), .Z(n16580) );
  XNOR U21049 ( .A(n16566), .B(n16581), .Z(n16573) );
  XNOR U21050 ( .A(n16563), .B(n16565), .Z(n16581) );
  AND U21051 ( .A(n16582), .B(n16583), .Z(n16565) );
  NANDN U21052 ( .A(n16584), .B(n16585), .Z(n16583) );
  NANDN U21053 ( .A(n16586), .B(n16587), .Z(n16585) );
  IV U21054 ( .A(n16588), .Z(n16587) );
  NAND U21055 ( .A(n16588), .B(n16586), .Z(n16582) );
  AND U21056 ( .A(n16589), .B(n16590), .Z(n16563) );
  NAND U21057 ( .A(n16591), .B(n16592), .Z(n16590) );
  OR U21058 ( .A(n16593), .B(n16594), .Z(n16592) );
  NAND U21059 ( .A(n16594), .B(n16593), .Z(n16589) );
  IV U21060 ( .A(n16595), .Z(n16594) );
  NAND U21061 ( .A(n16596), .B(n16597), .Z(n16566) );
  NANDN U21062 ( .A(n16598), .B(n16599), .Z(n16597) );
  NAND U21063 ( .A(n16600), .B(n16601), .Z(n16599) );
  OR U21064 ( .A(n16601), .B(n16600), .Z(n16596) );
  IV U21065 ( .A(n16602), .Z(n16600) );
  AND U21066 ( .A(n16603), .B(n16604), .Z(n16569) );
  NAND U21067 ( .A(n16605), .B(n16606), .Z(n16604) );
  NANDN U21068 ( .A(n16607), .B(n16608), .Z(n16606) );
  NANDN U21069 ( .A(n16608), .B(n16607), .Z(n16603) );
  XOR U21070 ( .A(n16579), .B(n16609), .Z(n16571) );
  XNOR U21071 ( .A(n16576), .B(n16578), .Z(n16609) );
  AND U21072 ( .A(n16610), .B(n16611), .Z(n16578) );
  NANDN U21073 ( .A(n16612), .B(n16613), .Z(n16611) );
  NANDN U21074 ( .A(n16614), .B(n16615), .Z(n16613) );
  IV U21075 ( .A(n16616), .Z(n16615) );
  NAND U21076 ( .A(n16616), .B(n16614), .Z(n16610) );
  AND U21077 ( .A(n16617), .B(n16618), .Z(n16576) );
  NAND U21078 ( .A(n16619), .B(n16620), .Z(n16618) );
  OR U21079 ( .A(n16621), .B(n16622), .Z(n16620) );
  NAND U21080 ( .A(n16622), .B(n16621), .Z(n16617) );
  IV U21081 ( .A(n16623), .Z(n16622) );
  NAND U21082 ( .A(n16624), .B(n16625), .Z(n16579) );
  NANDN U21083 ( .A(n16626), .B(n16627), .Z(n16625) );
  NAND U21084 ( .A(n16628), .B(n16629), .Z(n16627) );
  OR U21085 ( .A(n16629), .B(n16628), .Z(n16624) );
  IV U21086 ( .A(n16630), .Z(n16628) );
  XOR U21087 ( .A(n16605), .B(n16631), .Z(N28782) );
  XNOR U21088 ( .A(n16608), .B(n16607), .Z(n16631) );
  XNOR U21089 ( .A(n16619), .B(n16632), .Z(n16607) );
  XOR U21090 ( .A(n16623), .B(n16621), .Z(n16632) );
  XOR U21091 ( .A(n16629), .B(n16633), .Z(n16621) );
  XOR U21092 ( .A(n16626), .B(n16630), .Z(n16633) );
  NAND U21093 ( .A(n16634), .B(n16635), .Z(n16630) );
  NAND U21094 ( .A(n16636), .B(n16637), .Z(n16635) );
  NAND U21095 ( .A(n16638), .B(n16639), .Z(n16634) );
  AND U21096 ( .A(n16640), .B(n16641), .Z(n16626) );
  NAND U21097 ( .A(n16642), .B(n16643), .Z(n16641) );
  NAND U21098 ( .A(n16644), .B(n16645), .Z(n16640) );
  NANDN U21099 ( .A(n16646), .B(n16647), .Z(n16629) );
  NANDN U21100 ( .A(n16648), .B(n16649), .Z(n16623) );
  XNOR U21101 ( .A(n16614), .B(n16650), .Z(n16619) );
  XOR U21102 ( .A(n16612), .B(n16616), .Z(n16650) );
  NAND U21103 ( .A(n16651), .B(n16652), .Z(n16616) );
  NAND U21104 ( .A(n16653), .B(n16654), .Z(n16652) );
  NAND U21105 ( .A(n16655), .B(n16656), .Z(n16651) );
  AND U21106 ( .A(n16657), .B(n16658), .Z(n16612) );
  NAND U21107 ( .A(n16659), .B(n16660), .Z(n16658) );
  NAND U21108 ( .A(n16661), .B(n16662), .Z(n16657) );
  AND U21109 ( .A(n16663), .B(n16664), .Z(n16614) );
  NAND U21110 ( .A(n16665), .B(n16666), .Z(n16608) );
  XNOR U21111 ( .A(n16591), .B(n16667), .Z(n16605) );
  XOR U21112 ( .A(n16595), .B(n16593), .Z(n16667) );
  XOR U21113 ( .A(n16601), .B(n16668), .Z(n16593) );
  XOR U21114 ( .A(n16598), .B(n16602), .Z(n16668) );
  NAND U21115 ( .A(n16669), .B(n16670), .Z(n16602) );
  NAND U21116 ( .A(n16671), .B(n16672), .Z(n16670) );
  NAND U21117 ( .A(n16673), .B(n16674), .Z(n16669) );
  AND U21118 ( .A(n16675), .B(n16676), .Z(n16598) );
  NAND U21119 ( .A(n16677), .B(n16678), .Z(n16676) );
  NAND U21120 ( .A(n16679), .B(n16680), .Z(n16675) );
  NANDN U21121 ( .A(n16681), .B(n16682), .Z(n16601) );
  NANDN U21122 ( .A(n16683), .B(n16684), .Z(n16595) );
  XNOR U21123 ( .A(n16586), .B(n16685), .Z(n16591) );
  XOR U21124 ( .A(n16584), .B(n16588), .Z(n16685) );
  NAND U21125 ( .A(n16686), .B(n16687), .Z(n16588) );
  NAND U21126 ( .A(n16688), .B(n16689), .Z(n16687) );
  NAND U21127 ( .A(n16690), .B(n16691), .Z(n16686) );
  AND U21128 ( .A(n16692), .B(n16693), .Z(n16584) );
  NAND U21129 ( .A(n16694), .B(n16695), .Z(n16693) );
  NAND U21130 ( .A(n16696), .B(n16697), .Z(n16692) );
  AND U21131 ( .A(n16698), .B(n16699), .Z(n16586) );
  XOR U21132 ( .A(n16666), .B(n16665), .Z(N28781) );
  XNOR U21133 ( .A(n16684), .B(n16683), .Z(n16665) );
  XNOR U21134 ( .A(n16698), .B(n16699), .Z(n16683) );
  XOR U21135 ( .A(n16695), .B(n16694), .Z(n16699) );
  XOR U21136 ( .A(y[1707]), .B(x[1707]), .Z(n16694) );
  XOR U21137 ( .A(n16697), .B(n16696), .Z(n16695) );
  XOR U21138 ( .A(y[1709]), .B(x[1709]), .Z(n16696) );
  XOR U21139 ( .A(y[1708]), .B(x[1708]), .Z(n16697) );
  XOR U21140 ( .A(n16689), .B(n16688), .Z(n16698) );
  XOR U21141 ( .A(n16691), .B(n16690), .Z(n16688) );
  XOR U21142 ( .A(y[1706]), .B(x[1706]), .Z(n16690) );
  XOR U21143 ( .A(y[1705]), .B(x[1705]), .Z(n16691) );
  XOR U21144 ( .A(y[1704]), .B(x[1704]), .Z(n16689) );
  XNOR U21145 ( .A(n16682), .B(n16681), .Z(n16684) );
  XNOR U21146 ( .A(n16678), .B(n16677), .Z(n16681) );
  XOR U21147 ( .A(n16680), .B(n16679), .Z(n16677) );
  XOR U21148 ( .A(y[1703]), .B(x[1703]), .Z(n16679) );
  XOR U21149 ( .A(y[1702]), .B(x[1702]), .Z(n16680) );
  XOR U21150 ( .A(y[1701]), .B(x[1701]), .Z(n16678) );
  XOR U21151 ( .A(n16672), .B(n16671), .Z(n16682) );
  XOR U21152 ( .A(n16674), .B(n16673), .Z(n16671) );
  XOR U21153 ( .A(y[1700]), .B(x[1700]), .Z(n16673) );
  XOR U21154 ( .A(y[1699]), .B(x[1699]), .Z(n16674) );
  XOR U21155 ( .A(y[1698]), .B(x[1698]), .Z(n16672) );
  XNOR U21156 ( .A(n16649), .B(n16648), .Z(n16666) );
  XNOR U21157 ( .A(n16663), .B(n16664), .Z(n16648) );
  XOR U21158 ( .A(n16660), .B(n16659), .Z(n16664) );
  XOR U21159 ( .A(y[1695]), .B(x[1695]), .Z(n16659) );
  XOR U21160 ( .A(n16662), .B(n16661), .Z(n16660) );
  XOR U21161 ( .A(y[1697]), .B(x[1697]), .Z(n16661) );
  XOR U21162 ( .A(y[1696]), .B(x[1696]), .Z(n16662) );
  XOR U21163 ( .A(n16654), .B(n16653), .Z(n16663) );
  XOR U21164 ( .A(n16656), .B(n16655), .Z(n16653) );
  XOR U21165 ( .A(y[1694]), .B(x[1694]), .Z(n16655) );
  XOR U21166 ( .A(y[1693]), .B(x[1693]), .Z(n16656) );
  XOR U21167 ( .A(y[1692]), .B(x[1692]), .Z(n16654) );
  XNOR U21168 ( .A(n16647), .B(n16646), .Z(n16649) );
  XNOR U21169 ( .A(n16643), .B(n16642), .Z(n16646) );
  XOR U21170 ( .A(n16645), .B(n16644), .Z(n16642) );
  XOR U21171 ( .A(y[1691]), .B(x[1691]), .Z(n16644) );
  XOR U21172 ( .A(y[1690]), .B(x[1690]), .Z(n16645) );
  XOR U21173 ( .A(y[1689]), .B(x[1689]), .Z(n16643) );
  XOR U21174 ( .A(n16637), .B(n16636), .Z(n16647) );
  XOR U21175 ( .A(n16639), .B(n16638), .Z(n16636) );
  XOR U21176 ( .A(y[1688]), .B(x[1688]), .Z(n16638) );
  XOR U21177 ( .A(y[1687]), .B(x[1687]), .Z(n16639) );
  XOR U21178 ( .A(y[1686]), .B(x[1686]), .Z(n16637) );
  NAND U21179 ( .A(n16700), .B(n16701), .Z(N28773) );
  NAND U21180 ( .A(n16702), .B(n16703), .Z(n16701) );
  NANDN U21181 ( .A(n16704), .B(n16705), .Z(n16703) );
  NANDN U21182 ( .A(n16705), .B(n16704), .Z(n16700) );
  XOR U21183 ( .A(n16704), .B(n16706), .Z(N28772) );
  XNOR U21184 ( .A(n16702), .B(n16705), .Z(n16706) );
  NAND U21185 ( .A(n16707), .B(n16708), .Z(n16705) );
  NAND U21186 ( .A(n16709), .B(n16710), .Z(n16708) );
  NANDN U21187 ( .A(n16711), .B(n16712), .Z(n16710) );
  NANDN U21188 ( .A(n16712), .B(n16711), .Z(n16707) );
  AND U21189 ( .A(n16713), .B(n16714), .Z(n16702) );
  NAND U21190 ( .A(n16715), .B(n16716), .Z(n16714) );
  OR U21191 ( .A(n16717), .B(n16718), .Z(n16716) );
  NAND U21192 ( .A(n16718), .B(n16717), .Z(n16713) );
  IV U21193 ( .A(n16719), .Z(n16718) );
  AND U21194 ( .A(n16720), .B(n16721), .Z(n16704) );
  NAND U21195 ( .A(n16722), .B(n16723), .Z(n16721) );
  NANDN U21196 ( .A(n16724), .B(n16725), .Z(n16723) );
  NANDN U21197 ( .A(n16725), .B(n16724), .Z(n16720) );
  XOR U21198 ( .A(n16717), .B(n16726), .Z(N28771) );
  XOR U21199 ( .A(n16715), .B(n16719), .Z(n16726) );
  XNOR U21200 ( .A(n16712), .B(n16727), .Z(n16719) );
  XNOR U21201 ( .A(n16709), .B(n16711), .Z(n16727) );
  AND U21202 ( .A(n16728), .B(n16729), .Z(n16711) );
  NANDN U21203 ( .A(n16730), .B(n16731), .Z(n16729) );
  NANDN U21204 ( .A(n16732), .B(n16733), .Z(n16731) );
  IV U21205 ( .A(n16734), .Z(n16733) );
  NAND U21206 ( .A(n16734), .B(n16732), .Z(n16728) );
  AND U21207 ( .A(n16735), .B(n16736), .Z(n16709) );
  NAND U21208 ( .A(n16737), .B(n16738), .Z(n16736) );
  OR U21209 ( .A(n16739), .B(n16740), .Z(n16738) );
  NAND U21210 ( .A(n16740), .B(n16739), .Z(n16735) );
  IV U21211 ( .A(n16741), .Z(n16740) );
  NAND U21212 ( .A(n16742), .B(n16743), .Z(n16712) );
  NANDN U21213 ( .A(n16744), .B(n16745), .Z(n16743) );
  NAND U21214 ( .A(n16746), .B(n16747), .Z(n16745) );
  OR U21215 ( .A(n16747), .B(n16746), .Z(n16742) );
  IV U21216 ( .A(n16748), .Z(n16746) );
  AND U21217 ( .A(n16749), .B(n16750), .Z(n16715) );
  NAND U21218 ( .A(n16751), .B(n16752), .Z(n16750) );
  NANDN U21219 ( .A(n16753), .B(n16754), .Z(n16752) );
  NANDN U21220 ( .A(n16754), .B(n16753), .Z(n16749) );
  XOR U21221 ( .A(n16725), .B(n16755), .Z(n16717) );
  XNOR U21222 ( .A(n16722), .B(n16724), .Z(n16755) );
  AND U21223 ( .A(n16756), .B(n16757), .Z(n16724) );
  NANDN U21224 ( .A(n16758), .B(n16759), .Z(n16757) );
  NANDN U21225 ( .A(n16760), .B(n16761), .Z(n16759) );
  IV U21226 ( .A(n16762), .Z(n16761) );
  NAND U21227 ( .A(n16762), .B(n16760), .Z(n16756) );
  AND U21228 ( .A(n16763), .B(n16764), .Z(n16722) );
  NAND U21229 ( .A(n16765), .B(n16766), .Z(n16764) );
  OR U21230 ( .A(n16767), .B(n16768), .Z(n16766) );
  NAND U21231 ( .A(n16768), .B(n16767), .Z(n16763) );
  IV U21232 ( .A(n16769), .Z(n16768) );
  NAND U21233 ( .A(n16770), .B(n16771), .Z(n16725) );
  NANDN U21234 ( .A(n16772), .B(n16773), .Z(n16771) );
  NAND U21235 ( .A(n16774), .B(n16775), .Z(n16773) );
  OR U21236 ( .A(n16775), .B(n16774), .Z(n16770) );
  IV U21237 ( .A(n16776), .Z(n16774) );
  XOR U21238 ( .A(n16751), .B(n16777), .Z(N28770) );
  XNOR U21239 ( .A(n16754), .B(n16753), .Z(n16777) );
  XNOR U21240 ( .A(n16765), .B(n16778), .Z(n16753) );
  XOR U21241 ( .A(n16769), .B(n16767), .Z(n16778) );
  XOR U21242 ( .A(n16775), .B(n16779), .Z(n16767) );
  XOR U21243 ( .A(n16772), .B(n16776), .Z(n16779) );
  NAND U21244 ( .A(n16780), .B(n16781), .Z(n16776) );
  NAND U21245 ( .A(n16782), .B(n16783), .Z(n16781) );
  NAND U21246 ( .A(n16784), .B(n16785), .Z(n16780) );
  AND U21247 ( .A(n16786), .B(n16787), .Z(n16772) );
  NAND U21248 ( .A(n16788), .B(n16789), .Z(n16787) );
  NAND U21249 ( .A(n16790), .B(n16791), .Z(n16786) );
  NANDN U21250 ( .A(n16792), .B(n16793), .Z(n16775) );
  NANDN U21251 ( .A(n16794), .B(n16795), .Z(n16769) );
  XNOR U21252 ( .A(n16760), .B(n16796), .Z(n16765) );
  XOR U21253 ( .A(n16758), .B(n16762), .Z(n16796) );
  NAND U21254 ( .A(n16797), .B(n16798), .Z(n16762) );
  NAND U21255 ( .A(n16799), .B(n16800), .Z(n16798) );
  NAND U21256 ( .A(n16801), .B(n16802), .Z(n16797) );
  AND U21257 ( .A(n16803), .B(n16804), .Z(n16758) );
  NAND U21258 ( .A(n16805), .B(n16806), .Z(n16804) );
  NAND U21259 ( .A(n16807), .B(n16808), .Z(n16803) );
  AND U21260 ( .A(n16809), .B(n16810), .Z(n16760) );
  NAND U21261 ( .A(n16811), .B(n16812), .Z(n16754) );
  XNOR U21262 ( .A(n16737), .B(n16813), .Z(n16751) );
  XOR U21263 ( .A(n16741), .B(n16739), .Z(n16813) );
  XOR U21264 ( .A(n16747), .B(n16814), .Z(n16739) );
  XOR U21265 ( .A(n16744), .B(n16748), .Z(n16814) );
  NAND U21266 ( .A(n16815), .B(n16816), .Z(n16748) );
  NAND U21267 ( .A(n16817), .B(n16818), .Z(n16816) );
  NAND U21268 ( .A(n16819), .B(n16820), .Z(n16815) );
  AND U21269 ( .A(n16821), .B(n16822), .Z(n16744) );
  NAND U21270 ( .A(n16823), .B(n16824), .Z(n16822) );
  NAND U21271 ( .A(n16825), .B(n16826), .Z(n16821) );
  NANDN U21272 ( .A(n16827), .B(n16828), .Z(n16747) );
  NANDN U21273 ( .A(n16829), .B(n16830), .Z(n16741) );
  XNOR U21274 ( .A(n16732), .B(n16831), .Z(n16737) );
  XOR U21275 ( .A(n16730), .B(n16734), .Z(n16831) );
  NAND U21276 ( .A(n16832), .B(n16833), .Z(n16734) );
  NAND U21277 ( .A(n16834), .B(n16835), .Z(n16833) );
  NAND U21278 ( .A(n16836), .B(n16837), .Z(n16832) );
  AND U21279 ( .A(n16838), .B(n16839), .Z(n16730) );
  NAND U21280 ( .A(n16840), .B(n16841), .Z(n16839) );
  NAND U21281 ( .A(n16842), .B(n16843), .Z(n16838) );
  AND U21282 ( .A(n16844), .B(n16845), .Z(n16732) );
  XOR U21283 ( .A(n16812), .B(n16811), .Z(N28769) );
  XNOR U21284 ( .A(n16830), .B(n16829), .Z(n16811) );
  XNOR U21285 ( .A(n16844), .B(n16845), .Z(n16829) );
  XOR U21286 ( .A(n16841), .B(n16840), .Z(n16845) );
  XOR U21287 ( .A(y[1683]), .B(x[1683]), .Z(n16840) );
  XOR U21288 ( .A(n16843), .B(n16842), .Z(n16841) );
  XOR U21289 ( .A(y[1685]), .B(x[1685]), .Z(n16842) );
  XOR U21290 ( .A(y[1684]), .B(x[1684]), .Z(n16843) );
  XOR U21291 ( .A(n16835), .B(n16834), .Z(n16844) );
  XOR U21292 ( .A(n16837), .B(n16836), .Z(n16834) );
  XOR U21293 ( .A(y[1682]), .B(x[1682]), .Z(n16836) );
  XOR U21294 ( .A(y[1681]), .B(x[1681]), .Z(n16837) );
  XOR U21295 ( .A(y[1680]), .B(x[1680]), .Z(n16835) );
  XNOR U21296 ( .A(n16828), .B(n16827), .Z(n16830) );
  XNOR U21297 ( .A(n16824), .B(n16823), .Z(n16827) );
  XOR U21298 ( .A(n16826), .B(n16825), .Z(n16823) );
  XOR U21299 ( .A(y[1679]), .B(x[1679]), .Z(n16825) );
  XOR U21300 ( .A(y[1678]), .B(x[1678]), .Z(n16826) );
  XOR U21301 ( .A(y[1677]), .B(x[1677]), .Z(n16824) );
  XOR U21302 ( .A(n16818), .B(n16817), .Z(n16828) );
  XOR U21303 ( .A(n16820), .B(n16819), .Z(n16817) );
  XOR U21304 ( .A(y[1676]), .B(x[1676]), .Z(n16819) );
  XOR U21305 ( .A(y[1675]), .B(x[1675]), .Z(n16820) );
  XOR U21306 ( .A(y[1674]), .B(x[1674]), .Z(n16818) );
  XNOR U21307 ( .A(n16795), .B(n16794), .Z(n16812) );
  XNOR U21308 ( .A(n16809), .B(n16810), .Z(n16794) );
  XOR U21309 ( .A(n16806), .B(n16805), .Z(n16810) );
  XOR U21310 ( .A(y[1671]), .B(x[1671]), .Z(n16805) );
  XOR U21311 ( .A(n16808), .B(n16807), .Z(n16806) );
  XOR U21312 ( .A(y[1673]), .B(x[1673]), .Z(n16807) );
  XOR U21313 ( .A(y[1672]), .B(x[1672]), .Z(n16808) );
  XOR U21314 ( .A(n16800), .B(n16799), .Z(n16809) );
  XOR U21315 ( .A(n16802), .B(n16801), .Z(n16799) );
  XOR U21316 ( .A(y[1670]), .B(x[1670]), .Z(n16801) );
  XOR U21317 ( .A(y[1669]), .B(x[1669]), .Z(n16802) );
  XOR U21318 ( .A(y[1668]), .B(x[1668]), .Z(n16800) );
  XNOR U21319 ( .A(n16793), .B(n16792), .Z(n16795) );
  XNOR U21320 ( .A(n16789), .B(n16788), .Z(n16792) );
  XOR U21321 ( .A(n16791), .B(n16790), .Z(n16788) );
  XOR U21322 ( .A(y[1667]), .B(x[1667]), .Z(n16790) );
  XOR U21323 ( .A(y[1666]), .B(x[1666]), .Z(n16791) );
  XOR U21324 ( .A(y[1665]), .B(x[1665]), .Z(n16789) );
  XOR U21325 ( .A(n16783), .B(n16782), .Z(n16793) );
  XOR U21326 ( .A(n16785), .B(n16784), .Z(n16782) );
  XOR U21327 ( .A(y[1664]), .B(x[1664]), .Z(n16784) );
  XOR U21328 ( .A(y[1663]), .B(x[1663]), .Z(n16785) );
  XOR U21329 ( .A(y[1662]), .B(x[1662]), .Z(n16783) );
  NAND U21330 ( .A(n16846), .B(n16847), .Z(N28761) );
  NAND U21331 ( .A(n16848), .B(n16849), .Z(n16847) );
  NANDN U21332 ( .A(n16850), .B(n16851), .Z(n16849) );
  NANDN U21333 ( .A(n16851), .B(n16850), .Z(n16846) );
  XOR U21334 ( .A(n16850), .B(n16852), .Z(N28760) );
  XNOR U21335 ( .A(n16848), .B(n16851), .Z(n16852) );
  NAND U21336 ( .A(n16853), .B(n16854), .Z(n16851) );
  NAND U21337 ( .A(n16855), .B(n16856), .Z(n16854) );
  NANDN U21338 ( .A(n16857), .B(n16858), .Z(n16856) );
  NANDN U21339 ( .A(n16858), .B(n16857), .Z(n16853) );
  AND U21340 ( .A(n16859), .B(n16860), .Z(n16848) );
  NAND U21341 ( .A(n16861), .B(n16862), .Z(n16860) );
  OR U21342 ( .A(n16863), .B(n16864), .Z(n16862) );
  NAND U21343 ( .A(n16864), .B(n16863), .Z(n16859) );
  IV U21344 ( .A(n16865), .Z(n16864) );
  AND U21345 ( .A(n16866), .B(n16867), .Z(n16850) );
  NAND U21346 ( .A(n16868), .B(n16869), .Z(n16867) );
  NANDN U21347 ( .A(n16870), .B(n16871), .Z(n16869) );
  NANDN U21348 ( .A(n16871), .B(n16870), .Z(n16866) );
  XOR U21349 ( .A(n16863), .B(n16872), .Z(N28759) );
  XOR U21350 ( .A(n16861), .B(n16865), .Z(n16872) );
  XNOR U21351 ( .A(n16858), .B(n16873), .Z(n16865) );
  XNOR U21352 ( .A(n16855), .B(n16857), .Z(n16873) );
  AND U21353 ( .A(n16874), .B(n16875), .Z(n16857) );
  NANDN U21354 ( .A(n16876), .B(n16877), .Z(n16875) );
  NANDN U21355 ( .A(n16878), .B(n16879), .Z(n16877) );
  IV U21356 ( .A(n16880), .Z(n16879) );
  NAND U21357 ( .A(n16880), .B(n16878), .Z(n16874) );
  AND U21358 ( .A(n16881), .B(n16882), .Z(n16855) );
  NAND U21359 ( .A(n16883), .B(n16884), .Z(n16882) );
  OR U21360 ( .A(n16885), .B(n16886), .Z(n16884) );
  NAND U21361 ( .A(n16886), .B(n16885), .Z(n16881) );
  IV U21362 ( .A(n16887), .Z(n16886) );
  NAND U21363 ( .A(n16888), .B(n16889), .Z(n16858) );
  NANDN U21364 ( .A(n16890), .B(n16891), .Z(n16889) );
  NAND U21365 ( .A(n16892), .B(n16893), .Z(n16891) );
  OR U21366 ( .A(n16893), .B(n16892), .Z(n16888) );
  IV U21367 ( .A(n16894), .Z(n16892) );
  AND U21368 ( .A(n16895), .B(n16896), .Z(n16861) );
  NAND U21369 ( .A(n16897), .B(n16898), .Z(n16896) );
  NANDN U21370 ( .A(n16899), .B(n16900), .Z(n16898) );
  NANDN U21371 ( .A(n16900), .B(n16899), .Z(n16895) );
  XOR U21372 ( .A(n16871), .B(n16901), .Z(n16863) );
  XNOR U21373 ( .A(n16868), .B(n16870), .Z(n16901) );
  AND U21374 ( .A(n16902), .B(n16903), .Z(n16870) );
  NANDN U21375 ( .A(n16904), .B(n16905), .Z(n16903) );
  NANDN U21376 ( .A(n16906), .B(n16907), .Z(n16905) );
  IV U21377 ( .A(n16908), .Z(n16907) );
  NAND U21378 ( .A(n16908), .B(n16906), .Z(n16902) );
  AND U21379 ( .A(n16909), .B(n16910), .Z(n16868) );
  NAND U21380 ( .A(n16911), .B(n16912), .Z(n16910) );
  OR U21381 ( .A(n16913), .B(n16914), .Z(n16912) );
  NAND U21382 ( .A(n16914), .B(n16913), .Z(n16909) );
  IV U21383 ( .A(n16915), .Z(n16914) );
  NAND U21384 ( .A(n16916), .B(n16917), .Z(n16871) );
  NANDN U21385 ( .A(n16918), .B(n16919), .Z(n16917) );
  NAND U21386 ( .A(n16920), .B(n16921), .Z(n16919) );
  OR U21387 ( .A(n16921), .B(n16920), .Z(n16916) );
  IV U21388 ( .A(n16922), .Z(n16920) );
  XOR U21389 ( .A(n16897), .B(n16923), .Z(N28758) );
  XNOR U21390 ( .A(n16900), .B(n16899), .Z(n16923) );
  XNOR U21391 ( .A(n16911), .B(n16924), .Z(n16899) );
  XOR U21392 ( .A(n16915), .B(n16913), .Z(n16924) );
  XOR U21393 ( .A(n16921), .B(n16925), .Z(n16913) );
  XOR U21394 ( .A(n16918), .B(n16922), .Z(n16925) );
  NAND U21395 ( .A(n16926), .B(n16927), .Z(n16922) );
  NAND U21396 ( .A(n16928), .B(n16929), .Z(n16927) );
  NAND U21397 ( .A(n16930), .B(n16931), .Z(n16926) );
  AND U21398 ( .A(n16932), .B(n16933), .Z(n16918) );
  NAND U21399 ( .A(n16934), .B(n16935), .Z(n16933) );
  NAND U21400 ( .A(n16936), .B(n16937), .Z(n16932) );
  NANDN U21401 ( .A(n16938), .B(n16939), .Z(n16921) );
  NANDN U21402 ( .A(n16940), .B(n16941), .Z(n16915) );
  XNOR U21403 ( .A(n16906), .B(n16942), .Z(n16911) );
  XOR U21404 ( .A(n16904), .B(n16908), .Z(n16942) );
  NAND U21405 ( .A(n16943), .B(n16944), .Z(n16908) );
  NAND U21406 ( .A(n16945), .B(n16946), .Z(n16944) );
  NAND U21407 ( .A(n16947), .B(n16948), .Z(n16943) );
  AND U21408 ( .A(n16949), .B(n16950), .Z(n16904) );
  NAND U21409 ( .A(n16951), .B(n16952), .Z(n16950) );
  NAND U21410 ( .A(n16953), .B(n16954), .Z(n16949) );
  AND U21411 ( .A(n16955), .B(n16956), .Z(n16906) );
  NAND U21412 ( .A(n16957), .B(n16958), .Z(n16900) );
  XNOR U21413 ( .A(n16883), .B(n16959), .Z(n16897) );
  XOR U21414 ( .A(n16887), .B(n16885), .Z(n16959) );
  XOR U21415 ( .A(n16893), .B(n16960), .Z(n16885) );
  XOR U21416 ( .A(n16890), .B(n16894), .Z(n16960) );
  NAND U21417 ( .A(n16961), .B(n16962), .Z(n16894) );
  NAND U21418 ( .A(n16963), .B(n16964), .Z(n16962) );
  NAND U21419 ( .A(n16965), .B(n16966), .Z(n16961) );
  AND U21420 ( .A(n16967), .B(n16968), .Z(n16890) );
  NAND U21421 ( .A(n16969), .B(n16970), .Z(n16968) );
  NAND U21422 ( .A(n16971), .B(n16972), .Z(n16967) );
  NANDN U21423 ( .A(n16973), .B(n16974), .Z(n16893) );
  NANDN U21424 ( .A(n16975), .B(n16976), .Z(n16887) );
  XNOR U21425 ( .A(n16878), .B(n16977), .Z(n16883) );
  XOR U21426 ( .A(n16876), .B(n16880), .Z(n16977) );
  NAND U21427 ( .A(n16978), .B(n16979), .Z(n16880) );
  NAND U21428 ( .A(n16980), .B(n16981), .Z(n16979) );
  NAND U21429 ( .A(n16982), .B(n16983), .Z(n16978) );
  AND U21430 ( .A(n16984), .B(n16985), .Z(n16876) );
  NAND U21431 ( .A(n16986), .B(n16987), .Z(n16985) );
  NAND U21432 ( .A(n16988), .B(n16989), .Z(n16984) );
  AND U21433 ( .A(n16990), .B(n16991), .Z(n16878) );
  XOR U21434 ( .A(n16958), .B(n16957), .Z(N28757) );
  XNOR U21435 ( .A(n16976), .B(n16975), .Z(n16957) );
  XNOR U21436 ( .A(n16990), .B(n16991), .Z(n16975) );
  XOR U21437 ( .A(n16987), .B(n16986), .Z(n16991) );
  XOR U21438 ( .A(y[1659]), .B(x[1659]), .Z(n16986) );
  XOR U21439 ( .A(n16989), .B(n16988), .Z(n16987) );
  XOR U21440 ( .A(y[1661]), .B(x[1661]), .Z(n16988) );
  XOR U21441 ( .A(y[1660]), .B(x[1660]), .Z(n16989) );
  XOR U21442 ( .A(n16981), .B(n16980), .Z(n16990) );
  XOR U21443 ( .A(n16983), .B(n16982), .Z(n16980) );
  XOR U21444 ( .A(y[1658]), .B(x[1658]), .Z(n16982) );
  XOR U21445 ( .A(y[1657]), .B(x[1657]), .Z(n16983) );
  XOR U21446 ( .A(y[1656]), .B(x[1656]), .Z(n16981) );
  XNOR U21447 ( .A(n16974), .B(n16973), .Z(n16976) );
  XNOR U21448 ( .A(n16970), .B(n16969), .Z(n16973) );
  XOR U21449 ( .A(n16972), .B(n16971), .Z(n16969) );
  XOR U21450 ( .A(y[1655]), .B(x[1655]), .Z(n16971) );
  XOR U21451 ( .A(y[1654]), .B(x[1654]), .Z(n16972) );
  XOR U21452 ( .A(y[1653]), .B(x[1653]), .Z(n16970) );
  XOR U21453 ( .A(n16964), .B(n16963), .Z(n16974) );
  XOR U21454 ( .A(n16966), .B(n16965), .Z(n16963) );
  XOR U21455 ( .A(y[1652]), .B(x[1652]), .Z(n16965) );
  XOR U21456 ( .A(y[1651]), .B(x[1651]), .Z(n16966) );
  XOR U21457 ( .A(y[1650]), .B(x[1650]), .Z(n16964) );
  XNOR U21458 ( .A(n16941), .B(n16940), .Z(n16958) );
  XNOR U21459 ( .A(n16955), .B(n16956), .Z(n16940) );
  XOR U21460 ( .A(n16952), .B(n16951), .Z(n16956) );
  XOR U21461 ( .A(y[1647]), .B(x[1647]), .Z(n16951) );
  XOR U21462 ( .A(n16954), .B(n16953), .Z(n16952) );
  XOR U21463 ( .A(y[1649]), .B(x[1649]), .Z(n16953) );
  XOR U21464 ( .A(y[1648]), .B(x[1648]), .Z(n16954) );
  XOR U21465 ( .A(n16946), .B(n16945), .Z(n16955) );
  XOR U21466 ( .A(n16948), .B(n16947), .Z(n16945) );
  XOR U21467 ( .A(y[1646]), .B(x[1646]), .Z(n16947) );
  XOR U21468 ( .A(y[1645]), .B(x[1645]), .Z(n16948) );
  XOR U21469 ( .A(y[1644]), .B(x[1644]), .Z(n16946) );
  XNOR U21470 ( .A(n16939), .B(n16938), .Z(n16941) );
  XNOR U21471 ( .A(n16935), .B(n16934), .Z(n16938) );
  XOR U21472 ( .A(n16937), .B(n16936), .Z(n16934) );
  XOR U21473 ( .A(y[1643]), .B(x[1643]), .Z(n16936) );
  XOR U21474 ( .A(y[1642]), .B(x[1642]), .Z(n16937) );
  XOR U21475 ( .A(y[1641]), .B(x[1641]), .Z(n16935) );
  XOR U21476 ( .A(n16929), .B(n16928), .Z(n16939) );
  XOR U21477 ( .A(n16931), .B(n16930), .Z(n16928) );
  XOR U21478 ( .A(y[1640]), .B(x[1640]), .Z(n16930) );
  XOR U21479 ( .A(y[1639]), .B(x[1639]), .Z(n16931) );
  XOR U21480 ( .A(y[1638]), .B(x[1638]), .Z(n16929) );
  NAND U21481 ( .A(n16992), .B(n16993), .Z(N28749) );
  NAND U21482 ( .A(n16994), .B(n16995), .Z(n16993) );
  NANDN U21483 ( .A(n16996), .B(n16997), .Z(n16995) );
  NANDN U21484 ( .A(n16997), .B(n16996), .Z(n16992) );
  XOR U21485 ( .A(n16996), .B(n16998), .Z(N28748) );
  XNOR U21486 ( .A(n16994), .B(n16997), .Z(n16998) );
  NAND U21487 ( .A(n16999), .B(n17000), .Z(n16997) );
  NAND U21488 ( .A(n17001), .B(n17002), .Z(n17000) );
  NANDN U21489 ( .A(n17003), .B(n17004), .Z(n17002) );
  NANDN U21490 ( .A(n17004), .B(n17003), .Z(n16999) );
  AND U21491 ( .A(n17005), .B(n17006), .Z(n16994) );
  NAND U21492 ( .A(n17007), .B(n17008), .Z(n17006) );
  OR U21493 ( .A(n17009), .B(n17010), .Z(n17008) );
  NAND U21494 ( .A(n17010), .B(n17009), .Z(n17005) );
  IV U21495 ( .A(n17011), .Z(n17010) );
  AND U21496 ( .A(n17012), .B(n17013), .Z(n16996) );
  NAND U21497 ( .A(n17014), .B(n17015), .Z(n17013) );
  NANDN U21498 ( .A(n17016), .B(n17017), .Z(n17015) );
  NANDN U21499 ( .A(n17017), .B(n17016), .Z(n17012) );
  XOR U21500 ( .A(n17009), .B(n17018), .Z(N28747) );
  XOR U21501 ( .A(n17007), .B(n17011), .Z(n17018) );
  XNOR U21502 ( .A(n17004), .B(n17019), .Z(n17011) );
  XNOR U21503 ( .A(n17001), .B(n17003), .Z(n17019) );
  AND U21504 ( .A(n17020), .B(n17021), .Z(n17003) );
  NANDN U21505 ( .A(n17022), .B(n17023), .Z(n17021) );
  NANDN U21506 ( .A(n17024), .B(n17025), .Z(n17023) );
  IV U21507 ( .A(n17026), .Z(n17025) );
  NAND U21508 ( .A(n17026), .B(n17024), .Z(n17020) );
  AND U21509 ( .A(n17027), .B(n17028), .Z(n17001) );
  NAND U21510 ( .A(n17029), .B(n17030), .Z(n17028) );
  OR U21511 ( .A(n17031), .B(n17032), .Z(n17030) );
  NAND U21512 ( .A(n17032), .B(n17031), .Z(n17027) );
  IV U21513 ( .A(n17033), .Z(n17032) );
  NAND U21514 ( .A(n17034), .B(n17035), .Z(n17004) );
  NANDN U21515 ( .A(n17036), .B(n17037), .Z(n17035) );
  NAND U21516 ( .A(n17038), .B(n17039), .Z(n17037) );
  OR U21517 ( .A(n17039), .B(n17038), .Z(n17034) );
  IV U21518 ( .A(n17040), .Z(n17038) );
  AND U21519 ( .A(n17041), .B(n17042), .Z(n17007) );
  NAND U21520 ( .A(n17043), .B(n17044), .Z(n17042) );
  NANDN U21521 ( .A(n17045), .B(n17046), .Z(n17044) );
  NANDN U21522 ( .A(n17046), .B(n17045), .Z(n17041) );
  XOR U21523 ( .A(n17017), .B(n17047), .Z(n17009) );
  XNOR U21524 ( .A(n17014), .B(n17016), .Z(n17047) );
  AND U21525 ( .A(n17048), .B(n17049), .Z(n17016) );
  NANDN U21526 ( .A(n17050), .B(n17051), .Z(n17049) );
  NANDN U21527 ( .A(n17052), .B(n17053), .Z(n17051) );
  IV U21528 ( .A(n17054), .Z(n17053) );
  NAND U21529 ( .A(n17054), .B(n17052), .Z(n17048) );
  AND U21530 ( .A(n17055), .B(n17056), .Z(n17014) );
  NAND U21531 ( .A(n17057), .B(n17058), .Z(n17056) );
  OR U21532 ( .A(n17059), .B(n17060), .Z(n17058) );
  NAND U21533 ( .A(n17060), .B(n17059), .Z(n17055) );
  IV U21534 ( .A(n17061), .Z(n17060) );
  NAND U21535 ( .A(n17062), .B(n17063), .Z(n17017) );
  NANDN U21536 ( .A(n17064), .B(n17065), .Z(n17063) );
  NAND U21537 ( .A(n17066), .B(n17067), .Z(n17065) );
  OR U21538 ( .A(n17067), .B(n17066), .Z(n17062) );
  IV U21539 ( .A(n17068), .Z(n17066) );
  XOR U21540 ( .A(n17043), .B(n17069), .Z(N28746) );
  XNOR U21541 ( .A(n17046), .B(n17045), .Z(n17069) );
  XNOR U21542 ( .A(n17057), .B(n17070), .Z(n17045) );
  XOR U21543 ( .A(n17061), .B(n17059), .Z(n17070) );
  XOR U21544 ( .A(n17067), .B(n17071), .Z(n17059) );
  XOR U21545 ( .A(n17064), .B(n17068), .Z(n17071) );
  NAND U21546 ( .A(n17072), .B(n17073), .Z(n17068) );
  NAND U21547 ( .A(n17074), .B(n17075), .Z(n17073) );
  NAND U21548 ( .A(n17076), .B(n17077), .Z(n17072) );
  AND U21549 ( .A(n17078), .B(n17079), .Z(n17064) );
  NAND U21550 ( .A(n17080), .B(n17081), .Z(n17079) );
  NAND U21551 ( .A(n17082), .B(n17083), .Z(n17078) );
  NANDN U21552 ( .A(n17084), .B(n17085), .Z(n17067) );
  NANDN U21553 ( .A(n17086), .B(n17087), .Z(n17061) );
  XNOR U21554 ( .A(n17052), .B(n17088), .Z(n17057) );
  XOR U21555 ( .A(n17050), .B(n17054), .Z(n17088) );
  NAND U21556 ( .A(n17089), .B(n17090), .Z(n17054) );
  NAND U21557 ( .A(n17091), .B(n17092), .Z(n17090) );
  NAND U21558 ( .A(n17093), .B(n17094), .Z(n17089) );
  AND U21559 ( .A(n17095), .B(n17096), .Z(n17050) );
  NAND U21560 ( .A(n17097), .B(n17098), .Z(n17096) );
  NAND U21561 ( .A(n17099), .B(n17100), .Z(n17095) );
  AND U21562 ( .A(n17101), .B(n17102), .Z(n17052) );
  NAND U21563 ( .A(n17103), .B(n17104), .Z(n17046) );
  XNOR U21564 ( .A(n17029), .B(n17105), .Z(n17043) );
  XOR U21565 ( .A(n17033), .B(n17031), .Z(n17105) );
  XOR U21566 ( .A(n17039), .B(n17106), .Z(n17031) );
  XOR U21567 ( .A(n17036), .B(n17040), .Z(n17106) );
  NAND U21568 ( .A(n17107), .B(n17108), .Z(n17040) );
  NAND U21569 ( .A(n17109), .B(n17110), .Z(n17108) );
  NAND U21570 ( .A(n17111), .B(n17112), .Z(n17107) );
  AND U21571 ( .A(n17113), .B(n17114), .Z(n17036) );
  NAND U21572 ( .A(n17115), .B(n17116), .Z(n17114) );
  NAND U21573 ( .A(n17117), .B(n17118), .Z(n17113) );
  NANDN U21574 ( .A(n17119), .B(n17120), .Z(n17039) );
  NANDN U21575 ( .A(n17121), .B(n17122), .Z(n17033) );
  XNOR U21576 ( .A(n17024), .B(n17123), .Z(n17029) );
  XOR U21577 ( .A(n17022), .B(n17026), .Z(n17123) );
  NAND U21578 ( .A(n17124), .B(n17125), .Z(n17026) );
  NAND U21579 ( .A(n17126), .B(n17127), .Z(n17125) );
  NAND U21580 ( .A(n17128), .B(n17129), .Z(n17124) );
  AND U21581 ( .A(n17130), .B(n17131), .Z(n17022) );
  NAND U21582 ( .A(n17132), .B(n17133), .Z(n17131) );
  NAND U21583 ( .A(n17134), .B(n17135), .Z(n17130) );
  AND U21584 ( .A(n17136), .B(n17137), .Z(n17024) );
  XOR U21585 ( .A(n17104), .B(n17103), .Z(N28745) );
  XNOR U21586 ( .A(n17122), .B(n17121), .Z(n17103) );
  XNOR U21587 ( .A(n17136), .B(n17137), .Z(n17121) );
  XOR U21588 ( .A(n17133), .B(n17132), .Z(n17137) );
  XOR U21589 ( .A(y[1635]), .B(x[1635]), .Z(n17132) );
  XOR U21590 ( .A(n17135), .B(n17134), .Z(n17133) );
  XOR U21591 ( .A(y[1637]), .B(x[1637]), .Z(n17134) );
  XOR U21592 ( .A(y[1636]), .B(x[1636]), .Z(n17135) );
  XOR U21593 ( .A(n17127), .B(n17126), .Z(n17136) );
  XOR U21594 ( .A(n17129), .B(n17128), .Z(n17126) );
  XOR U21595 ( .A(y[1634]), .B(x[1634]), .Z(n17128) );
  XOR U21596 ( .A(y[1633]), .B(x[1633]), .Z(n17129) );
  XOR U21597 ( .A(y[1632]), .B(x[1632]), .Z(n17127) );
  XNOR U21598 ( .A(n17120), .B(n17119), .Z(n17122) );
  XNOR U21599 ( .A(n17116), .B(n17115), .Z(n17119) );
  XOR U21600 ( .A(n17118), .B(n17117), .Z(n17115) );
  XOR U21601 ( .A(y[1631]), .B(x[1631]), .Z(n17117) );
  XOR U21602 ( .A(y[1630]), .B(x[1630]), .Z(n17118) );
  XOR U21603 ( .A(y[1629]), .B(x[1629]), .Z(n17116) );
  XOR U21604 ( .A(n17110), .B(n17109), .Z(n17120) );
  XOR U21605 ( .A(n17112), .B(n17111), .Z(n17109) );
  XOR U21606 ( .A(y[1628]), .B(x[1628]), .Z(n17111) );
  XOR U21607 ( .A(y[1627]), .B(x[1627]), .Z(n17112) );
  XOR U21608 ( .A(y[1626]), .B(x[1626]), .Z(n17110) );
  XNOR U21609 ( .A(n17087), .B(n17086), .Z(n17104) );
  XNOR U21610 ( .A(n17101), .B(n17102), .Z(n17086) );
  XOR U21611 ( .A(n17098), .B(n17097), .Z(n17102) );
  XOR U21612 ( .A(y[1623]), .B(x[1623]), .Z(n17097) );
  XOR U21613 ( .A(n17100), .B(n17099), .Z(n17098) );
  XOR U21614 ( .A(y[1625]), .B(x[1625]), .Z(n17099) );
  XOR U21615 ( .A(y[1624]), .B(x[1624]), .Z(n17100) );
  XOR U21616 ( .A(n17092), .B(n17091), .Z(n17101) );
  XOR U21617 ( .A(n17094), .B(n17093), .Z(n17091) );
  XOR U21618 ( .A(y[1622]), .B(x[1622]), .Z(n17093) );
  XOR U21619 ( .A(y[1621]), .B(x[1621]), .Z(n17094) );
  XOR U21620 ( .A(y[1620]), .B(x[1620]), .Z(n17092) );
  XNOR U21621 ( .A(n17085), .B(n17084), .Z(n17087) );
  XNOR U21622 ( .A(n17081), .B(n17080), .Z(n17084) );
  XOR U21623 ( .A(n17083), .B(n17082), .Z(n17080) );
  XOR U21624 ( .A(y[1619]), .B(x[1619]), .Z(n17082) );
  XOR U21625 ( .A(y[1618]), .B(x[1618]), .Z(n17083) );
  XOR U21626 ( .A(y[1617]), .B(x[1617]), .Z(n17081) );
  XOR U21627 ( .A(n17075), .B(n17074), .Z(n17085) );
  XOR U21628 ( .A(n17077), .B(n17076), .Z(n17074) );
  XOR U21629 ( .A(y[1616]), .B(x[1616]), .Z(n17076) );
  XOR U21630 ( .A(y[1615]), .B(x[1615]), .Z(n17077) );
  XOR U21631 ( .A(y[1614]), .B(x[1614]), .Z(n17075) );
  NAND U21632 ( .A(n17138), .B(n17139), .Z(N28737) );
  NAND U21633 ( .A(n17140), .B(n17141), .Z(n17139) );
  NANDN U21634 ( .A(n17142), .B(n17143), .Z(n17141) );
  NANDN U21635 ( .A(n17143), .B(n17142), .Z(n17138) );
  XOR U21636 ( .A(n17142), .B(n17144), .Z(N28736) );
  XNOR U21637 ( .A(n17140), .B(n17143), .Z(n17144) );
  NAND U21638 ( .A(n17145), .B(n17146), .Z(n17143) );
  NAND U21639 ( .A(n17147), .B(n17148), .Z(n17146) );
  NANDN U21640 ( .A(n17149), .B(n17150), .Z(n17148) );
  NANDN U21641 ( .A(n17150), .B(n17149), .Z(n17145) );
  AND U21642 ( .A(n17151), .B(n17152), .Z(n17140) );
  NAND U21643 ( .A(n17153), .B(n17154), .Z(n17152) );
  OR U21644 ( .A(n17155), .B(n17156), .Z(n17154) );
  NAND U21645 ( .A(n17156), .B(n17155), .Z(n17151) );
  IV U21646 ( .A(n17157), .Z(n17156) );
  AND U21647 ( .A(n17158), .B(n17159), .Z(n17142) );
  NAND U21648 ( .A(n17160), .B(n17161), .Z(n17159) );
  NANDN U21649 ( .A(n17162), .B(n17163), .Z(n17161) );
  NANDN U21650 ( .A(n17163), .B(n17162), .Z(n17158) );
  XOR U21651 ( .A(n17155), .B(n17164), .Z(N28735) );
  XOR U21652 ( .A(n17153), .B(n17157), .Z(n17164) );
  XNOR U21653 ( .A(n17150), .B(n17165), .Z(n17157) );
  XNOR U21654 ( .A(n17147), .B(n17149), .Z(n17165) );
  AND U21655 ( .A(n17166), .B(n17167), .Z(n17149) );
  NANDN U21656 ( .A(n17168), .B(n17169), .Z(n17167) );
  NANDN U21657 ( .A(n17170), .B(n17171), .Z(n17169) );
  IV U21658 ( .A(n17172), .Z(n17171) );
  NAND U21659 ( .A(n17172), .B(n17170), .Z(n17166) );
  AND U21660 ( .A(n17173), .B(n17174), .Z(n17147) );
  NAND U21661 ( .A(n17175), .B(n17176), .Z(n17174) );
  OR U21662 ( .A(n17177), .B(n17178), .Z(n17176) );
  NAND U21663 ( .A(n17178), .B(n17177), .Z(n17173) );
  IV U21664 ( .A(n17179), .Z(n17178) );
  NAND U21665 ( .A(n17180), .B(n17181), .Z(n17150) );
  NANDN U21666 ( .A(n17182), .B(n17183), .Z(n17181) );
  NAND U21667 ( .A(n17184), .B(n17185), .Z(n17183) );
  OR U21668 ( .A(n17185), .B(n17184), .Z(n17180) );
  IV U21669 ( .A(n17186), .Z(n17184) );
  AND U21670 ( .A(n17187), .B(n17188), .Z(n17153) );
  NAND U21671 ( .A(n17189), .B(n17190), .Z(n17188) );
  NANDN U21672 ( .A(n17191), .B(n17192), .Z(n17190) );
  NANDN U21673 ( .A(n17192), .B(n17191), .Z(n17187) );
  XOR U21674 ( .A(n17163), .B(n17193), .Z(n17155) );
  XNOR U21675 ( .A(n17160), .B(n17162), .Z(n17193) );
  AND U21676 ( .A(n17194), .B(n17195), .Z(n17162) );
  NANDN U21677 ( .A(n17196), .B(n17197), .Z(n17195) );
  NANDN U21678 ( .A(n17198), .B(n17199), .Z(n17197) );
  IV U21679 ( .A(n17200), .Z(n17199) );
  NAND U21680 ( .A(n17200), .B(n17198), .Z(n17194) );
  AND U21681 ( .A(n17201), .B(n17202), .Z(n17160) );
  NAND U21682 ( .A(n17203), .B(n17204), .Z(n17202) );
  OR U21683 ( .A(n17205), .B(n17206), .Z(n17204) );
  NAND U21684 ( .A(n17206), .B(n17205), .Z(n17201) );
  IV U21685 ( .A(n17207), .Z(n17206) );
  NAND U21686 ( .A(n17208), .B(n17209), .Z(n17163) );
  NANDN U21687 ( .A(n17210), .B(n17211), .Z(n17209) );
  NAND U21688 ( .A(n17212), .B(n17213), .Z(n17211) );
  OR U21689 ( .A(n17213), .B(n17212), .Z(n17208) );
  IV U21690 ( .A(n17214), .Z(n17212) );
  XOR U21691 ( .A(n17189), .B(n17215), .Z(N28734) );
  XNOR U21692 ( .A(n17192), .B(n17191), .Z(n17215) );
  XNOR U21693 ( .A(n17203), .B(n17216), .Z(n17191) );
  XOR U21694 ( .A(n17207), .B(n17205), .Z(n17216) );
  XOR U21695 ( .A(n17213), .B(n17217), .Z(n17205) );
  XOR U21696 ( .A(n17210), .B(n17214), .Z(n17217) );
  NAND U21697 ( .A(n17218), .B(n17219), .Z(n17214) );
  NAND U21698 ( .A(n17220), .B(n17221), .Z(n17219) );
  NAND U21699 ( .A(n17222), .B(n17223), .Z(n17218) );
  AND U21700 ( .A(n17224), .B(n17225), .Z(n17210) );
  NAND U21701 ( .A(n17226), .B(n17227), .Z(n17225) );
  NAND U21702 ( .A(n17228), .B(n17229), .Z(n17224) );
  NANDN U21703 ( .A(n17230), .B(n17231), .Z(n17213) );
  NANDN U21704 ( .A(n17232), .B(n17233), .Z(n17207) );
  XNOR U21705 ( .A(n17198), .B(n17234), .Z(n17203) );
  XOR U21706 ( .A(n17196), .B(n17200), .Z(n17234) );
  NAND U21707 ( .A(n17235), .B(n17236), .Z(n17200) );
  NAND U21708 ( .A(n17237), .B(n17238), .Z(n17236) );
  NAND U21709 ( .A(n17239), .B(n17240), .Z(n17235) );
  AND U21710 ( .A(n17241), .B(n17242), .Z(n17196) );
  NAND U21711 ( .A(n17243), .B(n17244), .Z(n17242) );
  NAND U21712 ( .A(n17245), .B(n17246), .Z(n17241) );
  AND U21713 ( .A(n17247), .B(n17248), .Z(n17198) );
  NAND U21714 ( .A(n17249), .B(n17250), .Z(n17192) );
  XNOR U21715 ( .A(n17175), .B(n17251), .Z(n17189) );
  XOR U21716 ( .A(n17179), .B(n17177), .Z(n17251) );
  XOR U21717 ( .A(n17185), .B(n17252), .Z(n17177) );
  XOR U21718 ( .A(n17182), .B(n17186), .Z(n17252) );
  NAND U21719 ( .A(n17253), .B(n17254), .Z(n17186) );
  NAND U21720 ( .A(n17255), .B(n17256), .Z(n17254) );
  NAND U21721 ( .A(n17257), .B(n17258), .Z(n17253) );
  AND U21722 ( .A(n17259), .B(n17260), .Z(n17182) );
  NAND U21723 ( .A(n17261), .B(n17262), .Z(n17260) );
  NAND U21724 ( .A(n17263), .B(n17264), .Z(n17259) );
  NANDN U21725 ( .A(n17265), .B(n17266), .Z(n17185) );
  NANDN U21726 ( .A(n17267), .B(n17268), .Z(n17179) );
  XNOR U21727 ( .A(n17170), .B(n17269), .Z(n17175) );
  XOR U21728 ( .A(n17168), .B(n17172), .Z(n17269) );
  NAND U21729 ( .A(n17270), .B(n17271), .Z(n17172) );
  NAND U21730 ( .A(n17272), .B(n17273), .Z(n17271) );
  NAND U21731 ( .A(n17274), .B(n17275), .Z(n17270) );
  AND U21732 ( .A(n17276), .B(n17277), .Z(n17168) );
  NAND U21733 ( .A(n17278), .B(n17279), .Z(n17277) );
  NAND U21734 ( .A(n17280), .B(n17281), .Z(n17276) );
  AND U21735 ( .A(n17282), .B(n17283), .Z(n17170) );
  XOR U21736 ( .A(n17250), .B(n17249), .Z(N28733) );
  XNOR U21737 ( .A(n17268), .B(n17267), .Z(n17249) );
  XNOR U21738 ( .A(n17282), .B(n17283), .Z(n17267) );
  XOR U21739 ( .A(n17279), .B(n17278), .Z(n17283) );
  XOR U21740 ( .A(y[1611]), .B(x[1611]), .Z(n17278) );
  XOR U21741 ( .A(n17281), .B(n17280), .Z(n17279) );
  XOR U21742 ( .A(y[1613]), .B(x[1613]), .Z(n17280) );
  XOR U21743 ( .A(y[1612]), .B(x[1612]), .Z(n17281) );
  XOR U21744 ( .A(n17273), .B(n17272), .Z(n17282) );
  XOR U21745 ( .A(n17275), .B(n17274), .Z(n17272) );
  XOR U21746 ( .A(y[1610]), .B(x[1610]), .Z(n17274) );
  XOR U21747 ( .A(y[1609]), .B(x[1609]), .Z(n17275) );
  XOR U21748 ( .A(y[1608]), .B(x[1608]), .Z(n17273) );
  XNOR U21749 ( .A(n17266), .B(n17265), .Z(n17268) );
  XNOR U21750 ( .A(n17262), .B(n17261), .Z(n17265) );
  XOR U21751 ( .A(n17264), .B(n17263), .Z(n17261) );
  XOR U21752 ( .A(y[1607]), .B(x[1607]), .Z(n17263) );
  XOR U21753 ( .A(y[1606]), .B(x[1606]), .Z(n17264) );
  XOR U21754 ( .A(y[1605]), .B(x[1605]), .Z(n17262) );
  XOR U21755 ( .A(n17256), .B(n17255), .Z(n17266) );
  XOR U21756 ( .A(n17258), .B(n17257), .Z(n17255) );
  XOR U21757 ( .A(y[1604]), .B(x[1604]), .Z(n17257) );
  XOR U21758 ( .A(y[1603]), .B(x[1603]), .Z(n17258) );
  XOR U21759 ( .A(y[1602]), .B(x[1602]), .Z(n17256) );
  XNOR U21760 ( .A(n17233), .B(n17232), .Z(n17250) );
  XNOR U21761 ( .A(n17247), .B(n17248), .Z(n17232) );
  XOR U21762 ( .A(n17244), .B(n17243), .Z(n17248) );
  XOR U21763 ( .A(y[1599]), .B(x[1599]), .Z(n17243) );
  XOR U21764 ( .A(n17246), .B(n17245), .Z(n17244) );
  XOR U21765 ( .A(y[1601]), .B(x[1601]), .Z(n17245) );
  XOR U21766 ( .A(y[1600]), .B(x[1600]), .Z(n17246) );
  XOR U21767 ( .A(n17238), .B(n17237), .Z(n17247) );
  XOR U21768 ( .A(n17240), .B(n17239), .Z(n17237) );
  XOR U21769 ( .A(y[1598]), .B(x[1598]), .Z(n17239) );
  XOR U21770 ( .A(y[1597]), .B(x[1597]), .Z(n17240) );
  XOR U21771 ( .A(y[1596]), .B(x[1596]), .Z(n17238) );
  XNOR U21772 ( .A(n17231), .B(n17230), .Z(n17233) );
  XNOR U21773 ( .A(n17227), .B(n17226), .Z(n17230) );
  XOR U21774 ( .A(n17229), .B(n17228), .Z(n17226) );
  XOR U21775 ( .A(y[1595]), .B(x[1595]), .Z(n17228) );
  XOR U21776 ( .A(y[1594]), .B(x[1594]), .Z(n17229) );
  XOR U21777 ( .A(y[1593]), .B(x[1593]), .Z(n17227) );
  XOR U21778 ( .A(n17221), .B(n17220), .Z(n17231) );
  XOR U21779 ( .A(n17223), .B(n17222), .Z(n17220) );
  XOR U21780 ( .A(y[1592]), .B(x[1592]), .Z(n17222) );
  XOR U21781 ( .A(y[1591]), .B(x[1591]), .Z(n17223) );
  XOR U21782 ( .A(y[1590]), .B(x[1590]), .Z(n17221) );
  NAND U21783 ( .A(n17284), .B(n17285), .Z(N28725) );
  NAND U21784 ( .A(n17286), .B(n17287), .Z(n17285) );
  NANDN U21785 ( .A(n17288), .B(n17289), .Z(n17287) );
  NANDN U21786 ( .A(n17289), .B(n17288), .Z(n17284) );
  XOR U21787 ( .A(n17288), .B(n17290), .Z(N28724) );
  XNOR U21788 ( .A(n17286), .B(n17289), .Z(n17290) );
  NAND U21789 ( .A(n17291), .B(n17292), .Z(n17289) );
  NAND U21790 ( .A(n17293), .B(n17294), .Z(n17292) );
  NANDN U21791 ( .A(n17295), .B(n17296), .Z(n17294) );
  NANDN U21792 ( .A(n17296), .B(n17295), .Z(n17291) );
  AND U21793 ( .A(n17297), .B(n17298), .Z(n17286) );
  NAND U21794 ( .A(n17299), .B(n17300), .Z(n17298) );
  OR U21795 ( .A(n17301), .B(n17302), .Z(n17300) );
  NAND U21796 ( .A(n17302), .B(n17301), .Z(n17297) );
  IV U21797 ( .A(n17303), .Z(n17302) );
  AND U21798 ( .A(n17304), .B(n17305), .Z(n17288) );
  NAND U21799 ( .A(n17306), .B(n17307), .Z(n17305) );
  NANDN U21800 ( .A(n17308), .B(n17309), .Z(n17307) );
  NANDN U21801 ( .A(n17309), .B(n17308), .Z(n17304) );
  XOR U21802 ( .A(n17301), .B(n17310), .Z(N28723) );
  XOR U21803 ( .A(n17299), .B(n17303), .Z(n17310) );
  XNOR U21804 ( .A(n17296), .B(n17311), .Z(n17303) );
  XNOR U21805 ( .A(n17293), .B(n17295), .Z(n17311) );
  AND U21806 ( .A(n17312), .B(n17313), .Z(n17295) );
  NANDN U21807 ( .A(n17314), .B(n17315), .Z(n17313) );
  NANDN U21808 ( .A(n17316), .B(n17317), .Z(n17315) );
  IV U21809 ( .A(n17318), .Z(n17317) );
  NAND U21810 ( .A(n17318), .B(n17316), .Z(n17312) );
  AND U21811 ( .A(n17319), .B(n17320), .Z(n17293) );
  NAND U21812 ( .A(n17321), .B(n17322), .Z(n17320) );
  OR U21813 ( .A(n17323), .B(n17324), .Z(n17322) );
  NAND U21814 ( .A(n17324), .B(n17323), .Z(n17319) );
  IV U21815 ( .A(n17325), .Z(n17324) );
  NAND U21816 ( .A(n17326), .B(n17327), .Z(n17296) );
  NANDN U21817 ( .A(n17328), .B(n17329), .Z(n17327) );
  NAND U21818 ( .A(n17330), .B(n17331), .Z(n17329) );
  OR U21819 ( .A(n17331), .B(n17330), .Z(n17326) );
  IV U21820 ( .A(n17332), .Z(n17330) );
  AND U21821 ( .A(n17333), .B(n17334), .Z(n17299) );
  NAND U21822 ( .A(n17335), .B(n17336), .Z(n17334) );
  NANDN U21823 ( .A(n17337), .B(n17338), .Z(n17336) );
  NANDN U21824 ( .A(n17338), .B(n17337), .Z(n17333) );
  XOR U21825 ( .A(n17309), .B(n17339), .Z(n17301) );
  XNOR U21826 ( .A(n17306), .B(n17308), .Z(n17339) );
  AND U21827 ( .A(n17340), .B(n17341), .Z(n17308) );
  NANDN U21828 ( .A(n17342), .B(n17343), .Z(n17341) );
  NANDN U21829 ( .A(n17344), .B(n17345), .Z(n17343) );
  IV U21830 ( .A(n17346), .Z(n17345) );
  NAND U21831 ( .A(n17346), .B(n17344), .Z(n17340) );
  AND U21832 ( .A(n17347), .B(n17348), .Z(n17306) );
  NAND U21833 ( .A(n17349), .B(n17350), .Z(n17348) );
  OR U21834 ( .A(n17351), .B(n17352), .Z(n17350) );
  NAND U21835 ( .A(n17352), .B(n17351), .Z(n17347) );
  IV U21836 ( .A(n17353), .Z(n17352) );
  NAND U21837 ( .A(n17354), .B(n17355), .Z(n17309) );
  NANDN U21838 ( .A(n17356), .B(n17357), .Z(n17355) );
  NAND U21839 ( .A(n17358), .B(n17359), .Z(n17357) );
  OR U21840 ( .A(n17359), .B(n17358), .Z(n17354) );
  IV U21841 ( .A(n17360), .Z(n17358) );
  XOR U21842 ( .A(n17335), .B(n17361), .Z(N28722) );
  XNOR U21843 ( .A(n17338), .B(n17337), .Z(n17361) );
  XNOR U21844 ( .A(n17349), .B(n17362), .Z(n17337) );
  XOR U21845 ( .A(n17353), .B(n17351), .Z(n17362) );
  XOR U21846 ( .A(n17359), .B(n17363), .Z(n17351) );
  XOR U21847 ( .A(n17356), .B(n17360), .Z(n17363) );
  NAND U21848 ( .A(n17364), .B(n17365), .Z(n17360) );
  NAND U21849 ( .A(n17366), .B(n17367), .Z(n17365) );
  NAND U21850 ( .A(n17368), .B(n17369), .Z(n17364) );
  AND U21851 ( .A(n17370), .B(n17371), .Z(n17356) );
  NAND U21852 ( .A(n17372), .B(n17373), .Z(n17371) );
  NAND U21853 ( .A(n17374), .B(n17375), .Z(n17370) );
  NANDN U21854 ( .A(n17376), .B(n17377), .Z(n17359) );
  NANDN U21855 ( .A(n17378), .B(n17379), .Z(n17353) );
  XNOR U21856 ( .A(n17344), .B(n17380), .Z(n17349) );
  XOR U21857 ( .A(n17342), .B(n17346), .Z(n17380) );
  NAND U21858 ( .A(n17381), .B(n17382), .Z(n17346) );
  NAND U21859 ( .A(n17383), .B(n17384), .Z(n17382) );
  NAND U21860 ( .A(n17385), .B(n17386), .Z(n17381) );
  AND U21861 ( .A(n17387), .B(n17388), .Z(n17342) );
  NAND U21862 ( .A(n17389), .B(n17390), .Z(n17388) );
  NAND U21863 ( .A(n17391), .B(n17392), .Z(n17387) );
  AND U21864 ( .A(n17393), .B(n17394), .Z(n17344) );
  NAND U21865 ( .A(n17395), .B(n17396), .Z(n17338) );
  XNOR U21866 ( .A(n17321), .B(n17397), .Z(n17335) );
  XOR U21867 ( .A(n17325), .B(n17323), .Z(n17397) );
  XOR U21868 ( .A(n17331), .B(n17398), .Z(n17323) );
  XOR U21869 ( .A(n17328), .B(n17332), .Z(n17398) );
  NAND U21870 ( .A(n17399), .B(n17400), .Z(n17332) );
  NAND U21871 ( .A(n17401), .B(n17402), .Z(n17400) );
  NAND U21872 ( .A(n17403), .B(n17404), .Z(n17399) );
  AND U21873 ( .A(n17405), .B(n17406), .Z(n17328) );
  NAND U21874 ( .A(n17407), .B(n17408), .Z(n17406) );
  NAND U21875 ( .A(n17409), .B(n17410), .Z(n17405) );
  NANDN U21876 ( .A(n17411), .B(n17412), .Z(n17331) );
  NANDN U21877 ( .A(n17413), .B(n17414), .Z(n17325) );
  XNOR U21878 ( .A(n17316), .B(n17415), .Z(n17321) );
  XOR U21879 ( .A(n17314), .B(n17318), .Z(n17415) );
  NAND U21880 ( .A(n17416), .B(n17417), .Z(n17318) );
  NAND U21881 ( .A(n17418), .B(n17419), .Z(n17417) );
  NAND U21882 ( .A(n17420), .B(n17421), .Z(n17416) );
  AND U21883 ( .A(n17422), .B(n17423), .Z(n17314) );
  NAND U21884 ( .A(n17424), .B(n17425), .Z(n17423) );
  NAND U21885 ( .A(n17426), .B(n17427), .Z(n17422) );
  AND U21886 ( .A(n17428), .B(n17429), .Z(n17316) );
  XOR U21887 ( .A(n17396), .B(n17395), .Z(N28721) );
  XNOR U21888 ( .A(n17414), .B(n17413), .Z(n17395) );
  XNOR U21889 ( .A(n17428), .B(n17429), .Z(n17413) );
  XOR U21890 ( .A(n17425), .B(n17424), .Z(n17429) );
  XOR U21891 ( .A(y[1587]), .B(x[1587]), .Z(n17424) );
  XOR U21892 ( .A(n17427), .B(n17426), .Z(n17425) );
  XOR U21893 ( .A(y[1589]), .B(x[1589]), .Z(n17426) );
  XOR U21894 ( .A(y[1588]), .B(x[1588]), .Z(n17427) );
  XOR U21895 ( .A(n17419), .B(n17418), .Z(n17428) );
  XOR U21896 ( .A(n17421), .B(n17420), .Z(n17418) );
  XOR U21897 ( .A(y[1586]), .B(x[1586]), .Z(n17420) );
  XOR U21898 ( .A(y[1585]), .B(x[1585]), .Z(n17421) );
  XOR U21899 ( .A(y[1584]), .B(x[1584]), .Z(n17419) );
  XNOR U21900 ( .A(n17412), .B(n17411), .Z(n17414) );
  XNOR U21901 ( .A(n17408), .B(n17407), .Z(n17411) );
  XOR U21902 ( .A(n17410), .B(n17409), .Z(n17407) );
  XOR U21903 ( .A(y[1583]), .B(x[1583]), .Z(n17409) );
  XOR U21904 ( .A(y[1582]), .B(x[1582]), .Z(n17410) );
  XOR U21905 ( .A(y[1581]), .B(x[1581]), .Z(n17408) );
  XOR U21906 ( .A(n17402), .B(n17401), .Z(n17412) );
  XOR U21907 ( .A(n17404), .B(n17403), .Z(n17401) );
  XOR U21908 ( .A(y[1580]), .B(x[1580]), .Z(n17403) );
  XOR U21909 ( .A(y[1579]), .B(x[1579]), .Z(n17404) );
  XOR U21910 ( .A(y[1578]), .B(x[1578]), .Z(n17402) );
  XNOR U21911 ( .A(n17379), .B(n17378), .Z(n17396) );
  XNOR U21912 ( .A(n17393), .B(n17394), .Z(n17378) );
  XOR U21913 ( .A(n17390), .B(n17389), .Z(n17394) );
  XOR U21914 ( .A(y[1575]), .B(x[1575]), .Z(n17389) );
  XOR U21915 ( .A(n17392), .B(n17391), .Z(n17390) );
  XOR U21916 ( .A(y[1577]), .B(x[1577]), .Z(n17391) );
  XOR U21917 ( .A(y[1576]), .B(x[1576]), .Z(n17392) );
  XOR U21918 ( .A(n17384), .B(n17383), .Z(n17393) );
  XOR U21919 ( .A(n17386), .B(n17385), .Z(n17383) );
  XOR U21920 ( .A(y[1574]), .B(x[1574]), .Z(n17385) );
  XOR U21921 ( .A(y[1573]), .B(x[1573]), .Z(n17386) );
  XOR U21922 ( .A(y[1572]), .B(x[1572]), .Z(n17384) );
  XNOR U21923 ( .A(n17377), .B(n17376), .Z(n17379) );
  XNOR U21924 ( .A(n17373), .B(n17372), .Z(n17376) );
  XOR U21925 ( .A(n17375), .B(n17374), .Z(n17372) );
  XOR U21926 ( .A(y[1571]), .B(x[1571]), .Z(n17374) );
  XOR U21927 ( .A(y[1570]), .B(x[1570]), .Z(n17375) );
  XOR U21928 ( .A(y[1569]), .B(x[1569]), .Z(n17373) );
  XOR U21929 ( .A(n17367), .B(n17366), .Z(n17377) );
  XOR U21930 ( .A(n17369), .B(n17368), .Z(n17366) );
  XOR U21931 ( .A(y[1568]), .B(x[1568]), .Z(n17368) );
  XOR U21932 ( .A(y[1567]), .B(x[1567]), .Z(n17369) );
  XOR U21933 ( .A(y[1566]), .B(x[1566]), .Z(n17367) );
  NAND U21934 ( .A(n17430), .B(n17431), .Z(N28713) );
  NAND U21935 ( .A(n17432), .B(n17433), .Z(n17431) );
  NANDN U21936 ( .A(n17434), .B(n17435), .Z(n17433) );
  NANDN U21937 ( .A(n17435), .B(n17434), .Z(n17430) );
  XOR U21938 ( .A(n17434), .B(n17436), .Z(N28712) );
  XNOR U21939 ( .A(n17432), .B(n17435), .Z(n17436) );
  NAND U21940 ( .A(n17437), .B(n17438), .Z(n17435) );
  NAND U21941 ( .A(n17439), .B(n17440), .Z(n17438) );
  NANDN U21942 ( .A(n17441), .B(n17442), .Z(n17440) );
  NANDN U21943 ( .A(n17442), .B(n17441), .Z(n17437) );
  AND U21944 ( .A(n17443), .B(n17444), .Z(n17432) );
  NAND U21945 ( .A(n17445), .B(n17446), .Z(n17444) );
  OR U21946 ( .A(n17447), .B(n17448), .Z(n17446) );
  NAND U21947 ( .A(n17448), .B(n17447), .Z(n17443) );
  IV U21948 ( .A(n17449), .Z(n17448) );
  AND U21949 ( .A(n17450), .B(n17451), .Z(n17434) );
  NAND U21950 ( .A(n17452), .B(n17453), .Z(n17451) );
  NANDN U21951 ( .A(n17454), .B(n17455), .Z(n17453) );
  NANDN U21952 ( .A(n17455), .B(n17454), .Z(n17450) );
  XOR U21953 ( .A(n17447), .B(n17456), .Z(N28711) );
  XOR U21954 ( .A(n17445), .B(n17449), .Z(n17456) );
  XNOR U21955 ( .A(n17442), .B(n17457), .Z(n17449) );
  XNOR U21956 ( .A(n17439), .B(n17441), .Z(n17457) );
  AND U21957 ( .A(n17458), .B(n17459), .Z(n17441) );
  NANDN U21958 ( .A(n17460), .B(n17461), .Z(n17459) );
  NANDN U21959 ( .A(n17462), .B(n17463), .Z(n17461) );
  IV U21960 ( .A(n17464), .Z(n17463) );
  NAND U21961 ( .A(n17464), .B(n17462), .Z(n17458) );
  AND U21962 ( .A(n17465), .B(n17466), .Z(n17439) );
  NAND U21963 ( .A(n17467), .B(n17468), .Z(n17466) );
  OR U21964 ( .A(n17469), .B(n17470), .Z(n17468) );
  NAND U21965 ( .A(n17470), .B(n17469), .Z(n17465) );
  IV U21966 ( .A(n17471), .Z(n17470) );
  NAND U21967 ( .A(n17472), .B(n17473), .Z(n17442) );
  NANDN U21968 ( .A(n17474), .B(n17475), .Z(n17473) );
  NAND U21969 ( .A(n17476), .B(n17477), .Z(n17475) );
  OR U21970 ( .A(n17477), .B(n17476), .Z(n17472) );
  IV U21971 ( .A(n17478), .Z(n17476) );
  AND U21972 ( .A(n17479), .B(n17480), .Z(n17445) );
  NAND U21973 ( .A(n17481), .B(n17482), .Z(n17480) );
  NANDN U21974 ( .A(n17483), .B(n17484), .Z(n17482) );
  NANDN U21975 ( .A(n17484), .B(n17483), .Z(n17479) );
  XOR U21976 ( .A(n17455), .B(n17485), .Z(n17447) );
  XNOR U21977 ( .A(n17452), .B(n17454), .Z(n17485) );
  AND U21978 ( .A(n17486), .B(n17487), .Z(n17454) );
  NANDN U21979 ( .A(n17488), .B(n17489), .Z(n17487) );
  NANDN U21980 ( .A(n17490), .B(n17491), .Z(n17489) );
  IV U21981 ( .A(n17492), .Z(n17491) );
  NAND U21982 ( .A(n17492), .B(n17490), .Z(n17486) );
  AND U21983 ( .A(n17493), .B(n17494), .Z(n17452) );
  NAND U21984 ( .A(n17495), .B(n17496), .Z(n17494) );
  OR U21985 ( .A(n17497), .B(n17498), .Z(n17496) );
  NAND U21986 ( .A(n17498), .B(n17497), .Z(n17493) );
  IV U21987 ( .A(n17499), .Z(n17498) );
  NAND U21988 ( .A(n17500), .B(n17501), .Z(n17455) );
  NANDN U21989 ( .A(n17502), .B(n17503), .Z(n17501) );
  NAND U21990 ( .A(n17504), .B(n17505), .Z(n17503) );
  OR U21991 ( .A(n17505), .B(n17504), .Z(n17500) );
  IV U21992 ( .A(n17506), .Z(n17504) );
  XOR U21993 ( .A(n17481), .B(n17507), .Z(N28710) );
  XNOR U21994 ( .A(n17484), .B(n17483), .Z(n17507) );
  XNOR U21995 ( .A(n17495), .B(n17508), .Z(n17483) );
  XOR U21996 ( .A(n17499), .B(n17497), .Z(n17508) );
  XOR U21997 ( .A(n17505), .B(n17509), .Z(n17497) );
  XOR U21998 ( .A(n17502), .B(n17506), .Z(n17509) );
  NAND U21999 ( .A(n17510), .B(n17511), .Z(n17506) );
  NAND U22000 ( .A(n17512), .B(n17513), .Z(n17511) );
  NAND U22001 ( .A(n17514), .B(n17515), .Z(n17510) );
  AND U22002 ( .A(n17516), .B(n17517), .Z(n17502) );
  NAND U22003 ( .A(n17518), .B(n17519), .Z(n17517) );
  NAND U22004 ( .A(n17520), .B(n17521), .Z(n17516) );
  NANDN U22005 ( .A(n17522), .B(n17523), .Z(n17505) );
  NANDN U22006 ( .A(n17524), .B(n17525), .Z(n17499) );
  XNOR U22007 ( .A(n17490), .B(n17526), .Z(n17495) );
  XOR U22008 ( .A(n17488), .B(n17492), .Z(n17526) );
  NAND U22009 ( .A(n17527), .B(n17528), .Z(n17492) );
  NAND U22010 ( .A(n17529), .B(n17530), .Z(n17528) );
  NAND U22011 ( .A(n17531), .B(n17532), .Z(n17527) );
  AND U22012 ( .A(n17533), .B(n17534), .Z(n17488) );
  NAND U22013 ( .A(n17535), .B(n17536), .Z(n17534) );
  NAND U22014 ( .A(n17537), .B(n17538), .Z(n17533) );
  AND U22015 ( .A(n17539), .B(n17540), .Z(n17490) );
  NAND U22016 ( .A(n17541), .B(n17542), .Z(n17484) );
  XNOR U22017 ( .A(n17467), .B(n17543), .Z(n17481) );
  XOR U22018 ( .A(n17471), .B(n17469), .Z(n17543) );
  XOR U22019 ( .A(n17477), .B(n17544), .Z(n17469) );
  XOR U22020 ( .A(n17474), .B(n17478), .Z(n17544) );
  NAND U22021 ( .A(n17545), .B(n17546), .Z(n17478) );
  NAND U22022 ( .A(n17547), .B(n17548), .Z(n17546) );
  NAND U22023 ( .A(n17549), .B(n17550), .Z(n17545) );
  AND U22024 ( .A(n17551), .B(n17552), .Z(n17474) );
  NAND U22025 ( .A(n17553), .B(n17554), .Z(n17552) );
  NAND U22026 ( .A(n17555), .B(n17556), .Z(n17551) );
  NANDN U22027 ( .A(n17557), .B(n17558), .Z(n17477) );
  NANDN U22028 ( .A(n17559), .B(n17560), .Z(n17471) );
  XNOR U22029 ( .A(n17462), .B(n17561), .Z(n17467) );
  XOR U22030 ( .A(n17460), .B(n17464), .Z(n17561) );
  NAND U22031 ( .A(n17562), .B(n17563), .Z(n17464) );
  NAND U22032 ( .A(n17564), .B(n17565), .Z(n17563) );
  NAND U22033 ( .A(n17566), .B(n17567), .Z(n17562) );
  AND U22034 ( .A(n17568), .B(n17569), .Z(n17460) );
  NAND U22035 ( .A(n17570), .B(n17571), .Z(n17569) );
  NAND U22036 ( .A(n17572), .B(n17573), .Z(n17568) );
  AND U22037 ( .A(n17574), .B(n17575), .Z(n17462) );
  XOR U22038 ( .A(n17542), .B(n17541), .Z(N28709) );
  XNOR U22039 ( .A(n17560), .B(n17559), .Z(n17541) );
  XNOR U22040 ( .A(n17574), .B(n17575), .Z(n17559) );
  XOR U22041 ( .A(n17571), .B(n17570), .Z(n17575) );
  XOR U22042 ( .A(y[1563]), .B(x[1563]), .Z(n17570) );
  XOR U22043 ( .A(n17573), .B(n17572), .Z(n17571) );
  XOR U22044 ( .A(y[1565]), .B(x[1565]), .Z(n17572) );
  XOR U22045 ( .A(y[1564]), .B(x[1564]), .Z(n17573) );
  XOR U22046 ( .A(n17565), .B(n17564), .Z(n17574) );
  XOR U22047 ( .A(n17567), .B(n17566), .Z(n17564) );
  XOR U22048 ( .A(y[1562]), .B(x[1562]), .Z(n17566) );
  XOR U22049 ( .A(y[1561]), .B(x[1561]), .Z(n17567) );
  XOR U22050 ( .A(y[1560]), .B(x[1560]), .Z(n17565) );
  XNOR U22051 ( .A(n17558), .B(n17557), .Z(n17560) );
  XNOR U22052 ( .A(n17554), .B(n17553), .Z(n17557) );
  XOR U22053 ( .A(n17556), .B(n17555), .Z(n17553) );
  XOR U22054 ( .A(y[1559]), .B(x[1559]), .Z(n17555) );
  XOR U22055 ( .A(y[1558]), .B(x[1558]), .Z(n17556) );
  XOR U22056 ( .A(y[1557]), .B(x[1557]), .Z(n17554) );
  XOR U22057 ( .A(n17548), .B(n17547), .Z(n17558) );
  XOR U22058 ( .A(n17550), .B(n17549), .Z(n17547) );
  XOR U22059 ( .A(y[1556]), .B(x[1556]), .Z(n17549) );
  XOR U22060 ( .A(y[1555]), .B(x[1555]), .Z(n17550) );
  XOR U22061 ( .A(y[1554]), .B(x[1554]), .Z(n17548) );
  XNOR U22062 ( .A(n17525), .B(n17524), .Z(n17542) );
  XNOR U22063 ( .A(n17539), .B(n17540), .Z(n17524) );
  XOR U22064 ( .A(n17536), .B(n17535), .Z(n17540) );
  XOR U22065 ( .A(y[1551]), .B(x[1551]), .Z(n17535) );
  XOR U22066 ( .A(n17538), .B(n17537), .Z(n17536) );
  XOR U22067 ( .A(y[1553]), .B(x[1553]), .Z(n17537) );
  XOR U22068 ( .A(y[1552]), .B(x[1552]), .Z(n17538) );
  XOR U22069 ( .A(n17530), .B(n17529), .Z(n17539) );
  XOR U22070 ( .A(n17532), .B(n17531), .Z(n17529) );
  XOR U22071 ( .A(y[1550]), .B(x[1550]), .Z(n17531) );
  XOR U22072 ( .A(y[1549]), .B(x[1549]), .Z(n17532) );
  XOR U22073 ( .A(y[1548]), .B(x[1548]), .Z(n17530) );
  XNOR U22074 ( .A(n17523), .B(n17522), .Z(n17525) );
  XNOR U22075 ( .A(n17519), .B(n17518), .Z(n17522) );
  XOR U22076 ( .A(n17521), .B(n17520), .Z(n17518) );
  XOR U22077 ( .A(y[1547]), .B(x[1547]), .Z(n17520) );
  XOR U22078 ( .A(y[1546]), .B(x[1546]), .Z(n17521) );
  XOR U22079 ( .A(y[1545]), .B(x[1545]), .Z(n17519) );
  XOR U22080 ( .A(n17513), .B(n17512), .Z(n17523) );
  XOR U22081 ( .A(n17515), .B(n17514), .Z(n17512) );
  XOR U22082 ( .A(y[1544]), .B(x[1544]), .Z(n17514) );
  XOR U22083 ( .A(y[1543]), .B(x[1543]), .Z(n17515) );
  XOR U22084 ( .A(y[1542]), .B(x[1542]), .Z(n17513) );
  NAND U22085 ( .A(n17576), .B(n17577), .Z(N28701) );
  NAND U22086 ( .A(n17578), .B(n17579), .Z(n17577) );
  NANDN U22087 ( .A(n17580), .B(n17581), .Z(n17579) );
  NANDN U22088 ( .A(n17581), .B(n17580), .Z(n17576) );
  XOR U22089 ( .A(n17580), .B(n17582), .Z(N28700) );
  XNOR U22090 ( .A(n17578), .B(n17581), .Z(n17582) );
  NAND U22091 ( .A(n17583), .B(n17584), .Z(n17581) );
  NAND U22092 ( .A(n17585), .B(n17586), .Z(n17584) );
  NANDN U22093 ( .A(n17587), .B(n17588), .Z(n17586) );
  NANDN U22094 ( .A(n17588), .B(n17587), .Z(n17583) );
  AND U22095 ( .A(n17589), .B(n17590), .Z(n17578) );
  NAND U22096 ( .A(n17591), .B(n17592), .Z(n17590) );
  OR U22097 ( .A(n17593), .B(n17594), .Z(n17592) );
  NAND U22098 ( .A(n17594), .B(n17593), .Z(n17589) );
  IV U22099 ( .A(n17595), .Z(n17594) );
  AND U22100 ( .A(n17596), .B(n17597), .Z(n17580) );
  NAND U22101 ( .A(n17598), .B(n17599), .Z(n17597) );
  NANDN U22102 ( .A(n17600), .B(n17601), .Z(n17599) );
  NANDN U22103 ( .A(n17601), .B(n17600), .Z(n17596) );
  XOR U22104 ( .A(n17593), .B(n17602), .Z(N28699) );
  XOR U22105 ( .A(n17591), .B(n17595), .Z(n17602) );
  XNOR U22106 ( .A(n17588), .B(n17603), .Z(n17595) );
  XNOR U22107 ( .A(n17585), .B(n17587), .Z(n17603) );
  AND U22108 ( .A(n17604), .B(n17605), .Z(n17587) );
  NANDN U22109 ( .A(n17606), .B(n17607), .Z(n17605) );
  NANDN U22110 ( .A(n17608), .B(n17609), .Z(n17607) );
  IV U22111 ( .A(n17610), .Z(n17609) );
  NAND U22112 ( .A(n17610), .B(n17608), .Z(n17604) );
  AND U22113 ( .A(n17611), .B(n17612), .Z(n17585) );
  NAND U22114 ( .A(n17613), .B(n17614), .Z(n17612) );
  OR U22115 ( .A(n17615), .B(n17616), .Z(n17614) );
  NAND U22116 ( .A(n17616), .B(n17615), .Z(n17611) );
  IV U22117 ( .A(n17617), .Z(n17616) );
  NAND U22118 ( .A(n17618), .B(n17619), .Z(n17588) );
  NANDN U22119 ( .A(n17620), .B(n17621), .Z(n17619) );
  NAND U22120 ( .A(n17622), .B(n17623), .Z(n17621) );
  OR U22121 ( .A(n17623), .B(n17622), .Z(n17618) );
  IV U22122 ( .A(n17624), .Z(n17622) );
  AND U22123 ( .A(n17625), .B(n17626), .Z(n17591) );
  NAND U22124 ( .A(n17627), .B(n17628), .Z(n17626) );
  NANDN U22125 ( .A(n17629), .B(n17630), .Z(n17628) );
  NANDN U22126 ( .A(n17630), .B(n17629), .Z(n17625) );
  XOR U22127 ( .A(n17601), .B(n17631), .Z(n17593) );
  XNOR U22128 ( .A(n17598), .B(n17600), .Z(n17631) );
  AND U22129 ( .A(n17632), .B(n17633), .Z(n17600) );
  NANDN U22130 ( .A(n17634), .B(n17635), .Z(n17633) );
  NANDN U22131 ( .A(n17636), .B(n17637), .Z(n17635) );
  IV U22132 ( .A(n17638), .Z(n17637) );
  NAND U22133 ( .A(n17638), .B(n17636), .Z(n17632) );
  AND U22134 ( .A(n17639), .B(n17640), .Z(n17598) );
  NAND U22135 ( .A(n17641), .B(n17642), .Z(n17640) );
  OR U22136 ( .A(n17643), .B(n17644), .Z(n17642) );
  NAND U22137 ( .A(n17644), .B(n17643), .Z(n17639) );
  IV U22138 ( .A(n17645), .Z(n17644) );
  NAND U22139 ( .A(n17646), .B(n17647), .Z(n17601) );
  NANDN U22140 ( .A(n17648), .B(n17649), .Z(n17647) );
  NAND U22141 ( .A(n17650), .B(n17651), .Z(n17649) );
  OR U22142 ( .A(n17651), .B(n17650), .Z(n17646) );
  IV U22143 ( .A(n17652), .Z(n17650) );
  XOR U22144 ( .A(n17627), .B(n17653), .Z(N28698) );
  XNOR U22145 ( .A(n17630), .B(n17629), .Z(n17653) );
  XNOR U22146 ( .A(n17641), .B(n17654), .Z(n17629) );
  XOR U22147 ( .A(n17645), .B(n17643), .Z(n17654) );
  XOR U22148 ( .A(n17651), .B(n17655), .Z(n17643) );
  XOR U22149 ( .A(n17648), .B(n17652), .Z(n17655) );
  NAND U22150 ( .A(n17656), .B(n17657), .Z(n17652) );
  NAND U22151 ( .A(n17658), .B(n17659), .Z(n17657) );
  NAND U22152 ( .A(n17660), .B(n17661), .Z(n17656) );
  AND U22153 ( .A(n17662), .B(n17663), .Z(n17648) );
  NAND U22154 ( .A(n17664), .B(n17665), .Z(n17663) );
  NAND U22155 ( .A(n17666), .B(n17667), .Z(n17662) );
  NANDN U22156 ( .A(n17668), .B(n17669), .Z(n17651) );
  NANDN U22157 ( .A(n17670), .B(n17671), .Z(n17645) );
  XNOR U22158 ( .A(n17636), .B(n17672), .Z(n17641) );
  XOR U22159 ( .A(n17634), .B(n17638), .Z(n17672) );
  NAND U22160 ( .A(n17673), .B(n17674), .Z(n17638) );
  NAND U22161 ( .A(n17675), .B(n17676), .Z(n17674) );
  NAND U22162 ( .A(n17677), .B(n17678), .Z(n17673) );
  AND U22163 ( .A(n17679), .B(n17680), .Z(n17634) );
  NAND U22164 ( .A(n17681), .B(n17682), .Z(n17680) );
  NAND U22165 ( .A(n17683), .B(n17684), .Z(n17679) );
  AND U22166 ( .A(n17685), .B(n17686), .Z(n17636) );
  NAND U22167 ( .A(n17687), .B(n17688), .Z(n17630) );
  XNOR U22168 ( .A(n17613), .B(n17689), .Z(n17627) );
  XOR U22169 ( .A(n17617), .B(n17615), .Z(n17689) );
  XOR U22170 ( .A(n17623), .B(n17690), .Z(n17615) );
  XOR U22171 ( .A(n17620), .B(n17624), .Z(n17690) );
  NAND U22172 ( .A(n17691), .B(n17692), .Z(n17624) );
  NAND U22173 ( .A(n17693), .B(n17694), .Z(n17692) );
  NAND U22174 ( .A(n17695), .B(n17696), .Z(n17691) );
  AND U22175 ( .A(n17697), .B(n17698), .Z(n17620) );
  NAND U22176 ( .A(n17699), .B(n17700), .Z(n17698) );
  NAND U22177 ( .A(n17701), .B(n17702), .Z(n17697) );
  NANDN U22178 ( .A(n17703), .B(n17704), .Z(n17623) );
  NANDN U22179 ( .A(n17705), .B(n17706), .Z(n17617) );
  XNOR U22180 ( .A(n17608), .B(n17707), .Z(n17613) );
  XOR U22181 ( .A(n17606), .B(n17610), .Z(n17707) );
  NAND U22182 ( .A(n17708), .B(n17709), .Z(n17610) );
  NAND U22183 ( .A(n17710), .B(n17711), .Z(n17709) );
  NAND U22184 ( .A(n17712), .B(n17713), .Z(n17708) );
  AND U22185 ( .A(n17714), .B(n17715), .Z(n17606) );
  NAND U22186 ( .A(n17716), .B(n17717), .Z(n17715) );
  NAND U22187 ( .A(n17718), .B(n17719), .Z(n17714) );
  AND U22188 ( .A(n17720), .B(n17721), .Z(n17608) );
  XOR U22189 ( .A(n17688), .B(n17687), .Z(N28697) );
  XNOR U22190 ( .A(n17706), .B(n17705), .Z(n17687) );
  XNOR U22191 ( .A(n17720), .B(n17721), .Z(n17705) );
  XOR U22192 ( .A(n17717), .B(n17716), .Z(n17721) );
  XOR U22193 ( .A(y[1539]), .B(x[1539]), .Z(n17716) );
  XOR U22194 ( .A(n17719), .B(n17718), .Z(n17717) );
  XOR U22195 ( .A(y[1541]), .B(x[1541]), .Z(n17718) );
  XOR U22196 ( .A(y[1540]), .B(x[1540]), .Z(n17719) );
  XOR U22197 ( .A(n17711), .B(n17710), .Z(n17720) );
  XOR U22198 ( .A(n17713), .B(n17712), .Z(n17710) );
  XOR U22199 ( .A(y[1538]), .B(x[1538]), .Z(n17712) );
  XOR U22200 ( .A(y[1537]), .B(x[1537]), .Z(n17713) );
  XOR U22201 ( .A(y[1536]), .B(x[1536]), .Z(n17711) );
  XNOR U22202 ( .A(n17704), .B(n17703), .Z(n17706) );
  XNOR U22203 ( .A(n17700), .B(n17699), .Z(n17703) );
  XOR U22204 ( .A(n17702), .B(n17701), .Z(n17699) );
  XOR U22205 ( .A(y[1535]), .B(x[1535]), .Z(n17701) );
  XOR U22206 ( .A(y[1534]), .B(x[1534]), .Z(n17702) );
  XOR U22207 ( .A(y[1533]), .B(x[1533]), .Z(n17700) );
  XOR U22208 ( .A(n17694), .B(n17693), .Z(n17704) );
  XOR U22209 ( .A(n17696), .B(n17695), .Z(n17693) );
  XOR U22210 ( .A(y[1532]), .B(x[1532]), .Z(n17695) );
  XOR U22211 ( .A(y[1531]), .B(x[1531]), .Z(n17696) );
  XOR U22212 ( .A(y[1530]), .B(x[1530]), .Z(n17694) );
  XNOR U22213 ( .A(n17671), .B(n17670), .Z(n17688) );
  XNOR U22214 ( .A(n17685), .B(n17686), .Z(n17670) );
  XOR U22215 ( .A(n17682), .B(n17681), .Z(n17686) );
  XOR U22216 ( .A(y[1527]), .B(x[1527]), .Z(n17681) );
  XOR U22217 ( .A(n17684), .B(n17683), .Z(n17682) );
  XOR U22218 ( .A(y[1529]), .B(x[1529]), .Z(n17683) );
  XOR U22219 ( .A(y[1528]), .B(x[1528]), .Z(n17684) );
  XOR U22220 ( .A(n17676), .B(n17675), .Z(n17685) );
  XOR U22221 ( .A(n17678), .B(n17677), .Z(n17675) );
  XOR U22222 ( .A(y[1526]), .B(x[1526]), .Z(n17677) );
  XOR U22223 ( .A(y[1525]), .B(x[1525]), .Z(n17678) );
  XOR U22224 ( .A(y[1524]), .B(x[1524]), .Z(n17676) );
  XNOR U22225 ( .A(n17669), .B(n17668), .Z(n17671) );
  XNOR U22226 ( .A(n17665), .B(n17664), .Z(n17668) );
  XOR U22227 ( .A(n17667), .B(n17666), .Z(n17664) );
  XOR U22228 ( .A(y[1523]), .B(x[1523]), .Z(n17666) );
  XOR U22229 ( .A(y[1522]), .B(x[1522]), .Z(n17667) );
  XOR U22230 ( .A(y[1521]), .B(x[1521]), .Z(n17665) );
  XOR U22231 ( .A(n17659), .B(n17658), .Z(n17669) );
  XOR U22232 ( .A(n17661), .B(n17660), .Z(n17658) );
  XOR U22233 ( .A(y[1520]), .B(x[1520]), .Z(n17660) );
  XOR U22234 ( .A(y[1519]), .B(x[1519]), .Z(n17661) );
  XOR U22235 ( .A(y[1518]), .B(x[1518]), .Z(n17659) );
  NAND U22236 ( .A(n17722), .B(n17723), .Z(N28689) );
  NAND U22237 ( .A(n17724), .B(n17725), .Z(n17723) );
  NANDN U22238 ( .A(n17726), .B(n17727), .Z(n17725) );
  NANDN U22239 ( .A(n17727), .B(n17726), .Z(n17722) );
  XOR U22240 ( .A(n17726), .B(n17728), .Z(N28688) );
  XNOR U22241 ( .A(n17724), .B(n17727), .Z(n17728) );
  NAND U22242 ( .A(n17729), .B(n17730), .Z(n17727) );
  NAND U22243 ( .A(n17731), .B(n17732), .Z(n17730) );
  NANDN U22244 ( .A(n17733), .B(n17734), .Z(n17732) );
  NANDN U22245 ( .A(n17734), .B(n17733), .Z(n17729) );
  AND U22246 ( .A(n17735), .B(n17736), .Z(n17724) );
  NAND U22247 ( .A(n17737), .B(n17738), .Z(n17736) );
  OR U22248 ( .A(n17739), .B(n17740), .Z(n17738) );
  NAND U22249 ( .A(n17740), .B(n17739), .Z(n17735) );
  IV U22250 ( .A(n17741), .Z(n17740) );
  AND U22251 ( .A(n17742), .B(n17743), .Z(n17726) );
  NAND U22252 ( .A(n17744), .B(n17745), .Z(n17743) );
  NANDN U22253 ( .A(n17746), .B(n17747), .Z(n17745) );
  NANDN U22254 ( .A(n17747), .B(n17746), .Z(n17742) );
  XOR U22255 ( .A(n17739), .B(n17748), .Z(N28687) );
  XOR U22256 ( .A(n17737), .B(n17741), .Z(n17748) );
  XNOR U22257 ( .A(n17734), .B(n17749), .Z(n17741) );
  XNOR U22258 ( .A(n17731), .B(n17733), .Z(n17749) );
  AND U22259 ( .A(n17750), .B(n17751), .Z(n17733) );
  NANDN U22260 ( .A(n17752), .B(n17753), .Z(n17751) );
  NANDN U22261 ( .A(n17754), .B(n17755), .Z(n17753) );
  IV U22262 ( .A(n17756), .Z(n17755) );
  NAND U22263 ( .A(n17756), .B(n17754), .Z(n17750) );
  AND U22264 ( .A(n17757), .B(n17758), .Z(n17731) );
  NAND U22265 ( .A(n17759), .B(n17760), .Z(n17758) );
  OR U22266 ( .A(n17761), .B(n17762), .Z(n17760) );
  NAND U22267 ( .A(n17762), .B(n17761), .Z(n17757) );
  IV U22268 ( .A(n17763), .Z(n17762) );
  NAND U22269 ( .A(n17764), .B(n17765), .Z(n17734) );
  NANDN U22270 ( .A(n17766), .B(n17767), .Z(n17765) );
  NAND U22271 ( .A(n17768), .B(n17769), .Z(n17767) );
  OR U22272 ( .A(n17769), .B(n17768), .Z(n17764) );
  IV U22273 ( .A(n17770), .Z(n17768) );
  AND U22274 ( .A(n17771), .B(n17772), .Z(n17737) );
  NAND U22275 ( .A(n17773), .B(n17774), .Z(n17772) );
  NANDN U22276 ( .A(n17775), .B(n17776), .Z(n17774) );
  NANDN U22277 ( .A(n17776), .B(n17775), .Z(n17771) );
  XOR U22278 ( .A(n17747), .B(n17777), .Z(n17739) );
  XNOR U22279 ( .A(n17744), .B(n17746), .Z(n17777) );
  AND U22280 ( .A(n17778), .B(n17779), .Z(n17746) );
  NANDN U22281 ( .A(n17780), .B(n17781), .Z(n17779) );
  NANDN U22282 ( .A(n17782), .B(n17783), .Z(n17781) );
  IV U22283 ( .A(n17784), .Z(n17783) );
  NAND U22284 ( .A(n17784), .B(n17782), .Z(n17778) );
  AND U22285 ( .A(n17785), .B(n17786), .Z(n17744) );
  NAND U22286 ( .A(n17787), .B(n17788), .Z(n17786) );
  OR U22287 ( .A(n17789), .B(n17790), .Z(n17788) );
  NAND U22288 ( .A(n17790), .B(n17789), .Z(n17785) );
  IV U22289 ( .A(n17791), .Z(n17790) );
  NAND U22290 ( .A(n17792), .B(n17793), .Z(n17747) );
  NANDN U22291 ( .A(n17794), .B(n17795), .Z(n17793) );
  NAND U22292 ( .A(n17796), .B(n17797), .Z(n17795) );
  OR U22293 ( .A(n17797), .B(n17796), .Z(n17792) );
  IV U22294 ( .A(n17798), .Z(n17796) );
  XOR U22295 ( .A(n17773), .B(n17799), .Z(N28686) );
  XNOR U22296 ( .A(n17776), .B(n17775), .Z(n17799) );
  XNOR U22297 ( .A(n17787), .B(n17800), .Z(n17775) );
  XOR U22298 ( .A(n17791), .B(n17789), .Z(n17800) );
  XOR U22299 ( .A(n17797), .B(n17801), .Z(n17789) );
  XOR U22300 ( .A(n17794), .B(n17798), .Z(n17801) );
  NAND U22301 ( .A(n17802), .B(n17803), .Z(n17798) );
  NAND U22302 ( .A(n17804), .B(n17805), .Z(n17803) );
  NAND U22303 ( .A(n17806), .B(n17807), .Z(n17802) );
  AND U22304 ( .A(n17808), .B(n17809), .Z(n17794) );
  NAND U22305 ( .A(n17810), .B(n17811), .Z(n17809) );
  NAND U22306 ( .A(n17812), .B(n17813), .Z(n17808) );
  NANDN U22307 ( .A(n17814), .B(n17815), .Z(n17797) );
  NANDN U22308 ( .A(n17816), .B(n17817), .Z(n17791) );
  XNOR U22309 ( .A(n17782), .B(n17818), .Z(n17787) );
  XOR U22310 ( .A(n17780), .B(n17784), .Z(n17818) );
  NAND U22311 ( .A(n17819), .B(n17820), .Z(n17784) );
  NAND U22312 ( .A(n17821), .B(n17822), .Z(n17820) );
  NAND U22313 ( .A(n17823), .B(n17824), .Z(n17819) );
  AND U22314 ( .A(n17825), .B(n17826), .Z(n17780) );
  NAND U22315 ( .A(n17827), .B(n17828), .Z(n17826) );
  NAND U22316 ( .A(n17829), .B(n17830), .Z(n17825) );
  AND U22317 ( .A(n17831), .B(n17832), .Z(n17782) );
  NAND U22318 ( .A(n17833), .B(n17834), .Z(n17776) );
  XNOR U22319 ( .A(n17759), .B(n17835), .Z(n17773) );
  XOR U22320 ( .A(n17763), .B(n17761), .Z(n17835) );
  XOR U22321 ( .A(n17769), .B(n17836), .Z(n17761) );
  XOR U22322 ( .A(n17766), .B(n17770), .Z(n17836) );
  NAND U22323 ( .A(n17837), .B(n17838), .Z(n17770) );
  NAND U22324 ( .A(n17839), .B(n17840), .Z(n17838) );
  NAND U22325 ( .A(n17841), .B(n17842), .Z(n17837) );
  AND U22326 ( .A(n17843), .B(n17844), .Z(n17766) );
  NAND U22327 ( .A(n17845), .B(n17846), .Z(n17844) );
  NAND U22328 ( .A(n17847), .B(n17848), .Z(n17843) );
  NANDN U22329 ( .A(n17849), .B(n17850), .Z(n17769) );
  NANDN U22330 ( .A(n17851), .B(n17852), .Z(n17763) );
  XNOR U22331 ( .A(n17754), .B(n17853), .Z(n17759) );
  XOR U22332 ( .A(n17752), .B(n17756), .Z(n17853) );
  NAND U22333 ( .A(n17854), .B(n17855), .Z(n17756) );
  NAND U22334 ( .A(n17856), .B(n17857), .Z(n17855) );
  NAND U22335 ( .A(n17858), .B(n17859), .Z(n17854) );
  AND U22336 ( .A(n17860), .B(n17861), .Z(n17752) );
  NAND U22337 ( .A(n17862), .B(n17863), .Z(n17861) );
  NAND U22338 ( .A(n17864), .B(n17865), .Z(n17860) );
  AND U22339 ( .A(n17866), .B(n17867), .Z(n17754) );
  XOR U22340 ( .A(n17834), .B(n17833), .Z(N28685) );
  XNOR U22341 ( .A(n17852), .B(n17851), .Z(n17833) );
  XNOR U22342 ( .A(n17866), .B(n17867), .Z(n17851) );
  XOR U22343 ( .A(n17863), .B(n17862), .Z(n17867) );
  XOR U22344 ( .A(y[1515]), .B(x[1515]), .Z(n17862) );
  XOR U22345 ( .A(n17865), .B(n17864), .Z(n17863) );
  XOR U22346 ( .A(y[1517]), .B(x[1517]), .Z(n17864) );
  XOR U22347 ( .A(y[1516]), .B(x[1516]), .Z(n17865) );
  XOR U22348 ( .A(n17857), .B(n17856), .Z(n17866) );
  XOR U22349 ( .A(n17859), .B(n17858), .Z(n17856) );
  XOR U22350 ( .A(y[1514]), .B(x[1514]), .Z(n17858) );
  XOR U22351 ( .A(y[1513]), .B(x[1513]), .Z(n17859) );
  XOR U22352 ( .A(y[1512]), .B(x[1512]), .Z(n17857) );
  XNOR U22353 ( .A(n17850), .B(n17849), .Z(n17852) );
  XNOR U22354 ( .A(n17846), .B(n17845), .Z(n17849) );
  XOR U22355 ( .A(n17848), .B(n17847), .Z(n17845) );
  XOR U22356 ( .A(y[1511]), .B(x[1511]), .Z(n17847) );
  XOR U22357 ( .A(y[1510]), .B(x[1510]), .Z(n17848) );
  XOR U22358 ( .A(y[1509]), .B(x[1509]), .Z(n17846) );
  XOR U22359 ( .A(n17840), .B(n17839), .Z(n17850) );
  XOR U22360 ( .A(n17842), .B(n17841), .Z(n17839) );
  XOR U22361 ( .A(y[1508]), .B(x[1508]), .Z(n17841) );
  XOR U22362 ( .A(y[1507]), .B(x[1507]), .Z(n17842) );
  XOR U22363 ( .A(y[1506]), .B(x[1506]), .Z(n17840) );
  XNOR U22364 ( .A(n17817), .B(n17816), .Z(n17834) );
  XNOR U22365 ( .A(n17831), .B(n17832), .Z(n17816) );
  XOR U22366 ( .A(n17828), .B(n17827), .Z(n17832) );
  XOR U22367 ( .A(y[1503]), .B(x[1503]), .Z(n17827) );
  XOR U22368 ( .A(n17830), .B(n17829), .Z(n17828) );
  XOR U22369 ( .A(y[1505]), .B(x[1505]), .Z(n17829) );
  XOR U22370 ( .A(y[1504]), .B(x[1504]), .Z(n17830) );
  XOR U22371 ( .A(n17822), .B(n17821), .Z(n17831) );
  XOR U22372 ( .A(n17824), .B(n17823), .Z(n17821) );
  XOR U22373 ( .A(y[1502]), .B(x[1502]), .Z(n17823) );
  XOR U22374 ( .A(y[1501]), .B(x[1501]), .Z(n17824) );
  XOR U22375 ( .A(y[1500]), .B(x[1500]), .Z(n17822) );
  XNOR U22376 ( .A(n17815), .B(n17814), .Z(n17817) );
  XNOR U22377 ( .A(n17811), .B(n17810), .Z(n17814) );
  XOR U22378 ( .A(n17813), .B(n17812), .Z(n17810) );
  XOR U22379 ( .A(y[1499]), .B(x[1499]), .Z(n17812) );
  XOR U22380 ( .A(y[1498]), .B(x[1498]), .Z(n17813) );
  XOR U22381 ( .A(y[1497]), .B(x[1497]), .Z(n17811) );
  XOR U22382 ( .A(n17805), .B(n17804), .Z(n17815) );
  XOR U22383 ( .A(n17807), .B(n17806), .Z(n17804) );
  XOR U22384 ( .A(y[1496]), .B(x[1496]), .Z(n17806) );
  XOR U22385 ( .A(y[1495]), .B(x[1495]), .Z(n17807) );
  XOR U22386 ( .A(y[1494]), .B(x[1494]), .Z(n17805) );
  NAND U22387 ( .A(n17868), .B(n17869), .Z(N28677) );
  NAND U22388 ( .A(n17870), .B(n17871), .Z(n17869) );
  NANDN U22389 ( .A(n17872), .B(n17873), .Z(n17871) );
  NANDN U22390 ( .A(n17873), .B(n17872), .Z(n17868) );
  XOR U22391 ( .A(n17872), .B(n17874), .Z(N28676) );
  XNOR U22392 ( .A(n17870), .B(n17873), .Z(n17874) );
  NAND U22393 ( .A(n17875), .B(n17876), .Z(n17873) );
  NAND U22394 ( .A(n17877), .B(n17878), .Z(n17876) );
  NANDN U22395 ( .A(n17879), .B(n17880), .Z(n17878) );
  NANDN U22396 ( .A(n17880), .B(n17879), .Z(n17875) );
  AND U22397 ( .A(n17881), .B(n17882), .Z(n17870) );
  NAND U22398 ( .A(n17883), .B(n17884), .Z(n17882) );
  OR U22399 ( .A(n17885), .B(n17886), .Z(n17884) );
  NAND U22400 ( .A(n17886), .B(n17885), .Z(n17881) );
  IV U22401 ( .A(n17887), .Z(n17886) );
  AND U22402 ( .A(n17888), .B(n17889), .Z(n17872) );
  NAND U22403 ( .A(n17890), .B(n17891), .Z(n17889) );
  NANDN U22404 ( .A(n17892), .B(n17893), .Z(n17891) );
  NANDN U22405 ( .A(n17893), .B(n17892), .Z(n17888) );
  XOR U22406 ( .A(n17885), .B(n17894), .Z(N28675) );
  XOR U22407 ( .A(n17883), .B(n17887), .Z(n17894) );
  XNOR U22408 ( .A(n17880), .B(n17895), .Z(n17887) );
  XNOR U22409 ( .A(n17877), .B(n17879), .Z(n17895) );
  AND U22410 ( .A(n17896), .B(n17897), .Z(n17879) );
  NANDN U22411 ( .A(n17898), .B(n17899), .Z(n17897) );
  NANDN U22412 ( .A(n17900), .B(n17901), .Z(n17899) );
  IV U22413 ( .A(n17902), .Z(n17901) );
  NAND U22414 ( .A(n17902), .B(n17900), .Z(n17896) );
  AND U22415 ( .A(n17903), .B(n17904), .Z(n17877) );
  NAND U22416 ( .A(n17905), .B(n17906), .Z(n17904) );
  OR U22417 ( .A(n17907), .B(n17908), .Z(n17906) );
  NAND U22418 ( .A(n17908), .B(n17907), .Z(n17903) );
  IV U22419 ( .A(n17909), .Z(n17908) );
  NAND U22420 ( .A(n17910), .B(n17911), .Z(n17880) );
  NANDN U22421 ( .A(n17912), .B(n17913), .Z(n17911) );
  NAND U22422 ( .A(n17914), .B(n17915), .Z(n17913) );
  OR U22423 ( .A(n17915), .B(n17914), .Z(n17910) );
  IV U22424 ( .A(n17916), .Z(n17914) );
  AND U22425 ( .A(n17917), .B(n17918), .Z(n17883) );
  NAND U22426 ( .A(n17919), .B(n17920), .Z(n17918) );
  NANDN U22427 ( .A(n17921), .B(n17922), .Z(n17920) );
  NANDN U22428 ( .A(n17922), .B(n17921), .Z(n17917) );
  XOR U22429 ( .A(n17893), .B(n17923), .Z(n17885) );
  XNOR U22430 ( .A(n17890), .B(n17892), .Z(n17923) );
  AND U22431 ( .A(n17924), .B(n17925), .Z(n17892) );
  NANDN U22432 ( .A(n17926), .B(n17927), .Z(n17925) );
  NANDN U22433 ( .A(n17928), .B(n17929), .Z(n17927) );
  IV U22434 ( .A(n17930), .Z(n17929) );
  NAND U22435 ( .A(n17930), .B(n17928), .Z(n17924) );
  AND U22436 ( .A(n17931), .B(n17932), .Z(n17890) );
  NAND U22437 ( .A(n17933), .B(n17934), .Z(n17932) );
  OR U22438 ( .A(n17935), .B(n17936), .Z(n17934) );
  NAND U22439 ( .A(n17936), .B(n17935), .Z(n17931) );
  IV U22440 ( .A(n17937), .Z(n17936) );
  NAND U22441 ( .A(n17938), .B(n17939), .Z(n17893) );
  NANDN U22442 ( .A(n17940), .B(n17941), .Z(n17939) );
  NAND U22443 ( .A(n17942), .B(n17943), .Z(n17941) );
  OR U22444 ( .A(n17943), .B(n17942), .Z(n17938) );
  IV U22445 ( .A(n17944), .Z(n17942) );
  XOR U22446 ( .A(n17919), .B(n17945), .Z(N28674) );
  XNOR U22447 ( .A(n17922), .B(n17921), .Z(n17945) );
  XNOR U22448 ( .A(n17933), .B(n17946), .Z(n17921) );
  XOR U22449 ( .A(n17937), .B(n17935), .Z(n17946) );
  XOR U22450 ( .A(n17943), .B(n17947), .Z(n17935) );
  XOR U22451 ( .A(n17940), .B(n17944), .Z(n17947) );
  NAND U22452 ( .A(n17948), .B(n17949), .Z(n17944) );
  NAND U22453 ( .A(n17950), .B(n17951), .Z(n17949) );
  NAND U22454 ( .A(n17952), .B(n17953), .Z(n17948) );
  AND U22455 ( .A(n17954), .B(n17955), .Z(n17940) );
  NAND U22456 ( .A(n17956), .B(n17957), .Z(n17955) );
  NAND U22457 ( .A(n17958), .B(n17959), .Z(n17954) );
  NANDN U22458 ( .A(n17960), .B(n17961), .Z(n17943) );
  NANDN U22459 ( .A(n17962), .B(n17963), .Z(n17937) );
  XNOR U22460 ( .A(n17928), .B(n17964), .Z(n17933) );
  XOR U22461 ( .A(n17926), .B(n17930), .Z(n17964) );
  NAND U22462 ( .A(n17965), .B(n17966), .Z(n17930) );
  NAND U22463 ( .A(n17967), .B(n17968), .Z(n17966) );
  NAND U22464 ( .A(n17969), .B(n17970), .Z(n17965) );
  AND U22465 ( .A(n17971), .B(n17972), .Z(n17926) );
  NAND U22466 ( .A(n17973), .B(n17974), .Z(n17972) );
  NAND U22467 ( .A(n17975), .B(n17976), .Z(n17971) );
  AND U22468 ( .A(n17977), .B(n17978), .Z(n17928) );
  NAND U22469 ( .A(n17979), .B(n17980), .Z(n17922) );
  XNOR U22470 ( .A(n17905), .B(n17981), .Z(n17919) );
  XOR U22471 ( .A(n17909), .B(n17907), .Z(n17981) );
  XOR U22472 ( .A(n17915), .B(n17982), .Z(n17907) );
  XOR U22473 ( .A(n17912), .B(n17916), .Z(n17982) );
  NAND U22474 ( .A(n17983), .B(n17984), .Z(n17916) );
  NAND U22475 ( .A(n17985), .B(n17986), .Z(n17984) );
  NAND U22476 ( .A(n17987), .B(n17988), .Z(n17983) );
  AND U22477 ( .A(n17989), .B(n17990), .Z(n17912) );
  NAND U22478 ( .A(n17991), .B(n17992), .Z(n17990) );
  NAND U22479 ( .A(n17993), .B(n17994), .Z(n17989) );
  NANDN U22480 ( .A(n17995), .B(n17996), .Z(n17915) );
  NANDN U22481 ( .A(n17997), .B(n17998), .Z(n17909) );
  XNOR U22482 ( .A(n17900), .B(n17999), .Z(n17905) );
  XOR U22483 ( .A(n17898), .B(n17902), .Z(n17999) );
  NAND U22484 ( .A(n18000), .B(n18001), .Z(n17902) );
  NAND U22485 ( .A(n18002), .B(n18003), .Z(n18001) );
  NAND U22486 ( .A(n18004), .B(n18005), .Z(n18000) );
  AND U22487 ( .A(n18006), .B(n18007), .Z(n17898) );
  NAND U22488 ( .A(n18008), .B(n18009), .Z(n18007) );
  NAND U22489 ( .A(n18010), .B(n18011), .Z(n18006) );
  AND U22490 ( .A(n18012), .B(n18013), .Z(n17900) );
  XOR U22491 ( .A(n17980), .B(n17979), .Z(N28673) );
  XNOR U22492 ( .A(n17998), .B(n17997), .Z(n17979) );
  XNOR U22493 ( .A(n18012), .B(n18013), .Z(n17997) );
  XOR U22494 ( .A(n18009), .B(n18008), .Z(n18013) );
  XOR U22495 ( .A(y[1491]), .B(x[1491]), .Z(n18008) );
  XOR U22496 ( .A(n18011), .B(n18010), .Z(n18009) );
  XOR U22497 ( .A(y[1493]), .B(x[1493]), .Z(n18010) );
  XOR U22498 ( .A(y[1492]), .B(x[1492]), .Z(n18011) );
  XOR U22499 ( .A(n18003), .B(n18002), .Z(n18012) );
  XOR U22500 ( .A(n18005), .B(n18004), .Z(n18002) );
  XOR U22501 ( .A(y[1490]), .B(x[1490]), .Z(n18004) );
  XOR U22502 ( .A(y[1489]), .B(x[1489]), .Z(n18005) );
  XOR U22503 ( .A(y[1488]), .B(x[1488]), .Z(n18003) );
  XNOR U22504 ( .A(n17996), .B(n17995), .Z(n17998) );
  XNOR U22505 ( .A(n17992), .B(n17991), .Z(n17995) );
  XOR U22506 ( .A(n17994), .B(n17993), .Z(n17991) );
  XOR U22507 ( .A(y[1487]), .B(x[1487]), .Z(n17993) );
  XOR U22508 ( .A(y[1486]), .B(x[1486]), .Z(n17994) );
  XOR U22509 ( .A(y[1485]), .B(x[1485]), .Z(n17992) );
  XOR U22510 ( .A(n17986), .B(n17985), .Z(n17996) );
  XOR U22511 ( .A(n17988), .B(n17987), .Z(n17985) );
  XOR U22512 ( .A(y[1484]), .B(x[1484]), .Z(n17987) );
  XOR U22513 ( .A(y[1483]), .B(x[1483]), .Z(n17988) );
  XOR U22514 ( .A(y[1482]), .B(x[1482]), .Z(n17986) );
  XNOR U22515 ( .A(n17963), .B(n17962), .Z(n17980) );
  XNOR U22516 ( .A(n17977), .B(n17978), .Z(n17962) );
  XOR U22517 ( .A(n17974), .B(n17973), .Z(n17978) );
  XOR U22518 ( .A(y[1479]), .B(x[1479]), .Z(n17973) );
  XOR U22519 ( .A(n17976), .B(n17975), .Z(n17974) );
  XOR U22520 ( .A(y[1481]), .B(x[1481]), .Z(n17975) );
  XOR U22521 ( .A(y[1480]), .B(x[1480]), .Z(n17976) );
  XOR U22522 ( .A(n17968), .B(n17967), .Z(n17977) );
  XOR U22523 ( .A(n17970), .B(n17969), .Z(n17967) );
  XOR U22524 ( .A(y[1478]), .B(x[1478]), .Z(n17969) );
  XOR U22525 ( .A(y[1477]), .B(x[1477]), .Z(n17970) );
  XOR U22526 ( .A(y[1476]), .B(x[1476]), .Z(n17968) );
  XNOR U22527 ( .A(n17961), .B(n17960), .Z(n17963) );
  XNOR U22528 ( .A(n17957), .B(n17956), .Z(n17960) );
  XOR U22529 ( .A(n17959), .B(n17958), .Z(n17956) );
  XOR U22530 ( .A(y[1475]), .B(x[1475]), .Z(n17958) );
  XOR U22531 ( .A(y[1474]), .B(x[1474]), .Z(n17959) );
  XOR U22532 ( .A(y[1473]), .B(x[1473]), .Z(n17957) );
  XOR U22533 ( .A(n17951), .B(n17950), .Z(n17961) );
  XOR U22534 ( .A(n17953), .B(n17952), .Z(n17950) );
  XOR U22535 ( .A(y[1472]), .B(x[1472]), .Z(n17952) );
  XOR U22536 ( .A(y[1471]), .B(x[1471]), .Z(n17953) );
  XOR U22537 ( .A(y[1470]), .B(x[1470]), .Z(n17951) );
  NAND U22538 ( .A(n18014), .B(n18015), .Z(N28665) );
  NAND U22539 ( .A(n18016), .B(n18017), .Z(n18015) );
  NANDN U22540 ( .A(n18018), .B(n18019), .Z(n18017) );
  NANDN U22541 ( .A(n18019), .B(n18018), .Z(n18014) );
  XOR U22542 ( .A(n18018), .B(n18020), .Z(N28664) );
  XNOR U22543 ( .A(n18016), .B(n18019), .Z(n18020) );
  NAND U22544 ( .A(n18021), .B(n18022), .Z(n18019) );
  NAND U22545 ( .A(n18023), .B(n18024), .Z(n18022) );
  NANDN U22546 ( .A(n18025), .B(n18026), .Z(n18024) );
  NANDN U22547 ( .A(n18026), .B(n18025), .Z(n18021) );
  AND U22548 ( .A(n18027), .B(n18028), .Z(n18016) );
  NAND U22549 ( .A(n18029), .B(n18030), .Z(n18028) );
  OR U22550 ( .A(n18031), .B(n18032), .Z(n18030) );
  NAND U22551 ( .A(n18032), .B(n18031), .Z(n18027) );
  IV U22552 ( .A(n18033), .Z(n18032) );
  AND U22553 ( .A(n18034), .B(n18035), .Z(n18018) );
  NAND U22554 ( .A(n18036), .B(n18037), .Z(n18035) );
  NANDN U22555 ( .A(n18038), .B(n18039), .Z(n18037) );
  NANDN U22556 ( .A(n18039), .B(n18038), .Z(n18034) );
  XOR U22557 ( .A(n18031), .B(n18040), .Z(N28663) );
  XOR U22558 ( .A(n18029), .B(n18033), .Z(n18040) );
  XNOR U22559 ( .A(n18026), .B(n18041), .Z(n18033) );
  XNOR U22560 ( .A(n18023), .B(n18025), .Z(n18041) );
  AND U22561 ( .A(n18042), .B(n18043), .Z(n18025) );
  NANDN U22562 ( .A(n18044), .B(n18045), .Z(n18043) );
  NANDN U22563 ( .A(n18046), .B(n18047), .Z(n18045) );
  IV U22564 ( .A(n18048), .Z(n18047) );
  NAND U22565 ( .A(n18048), .B(n18046), .Z(n18042) );
  AND U22566 ( .A(n18049), .B(n18050), .Z(n18023) );
  NAND U22567 ( .A(n18051), .B(n18052), .Z(n18050) );
  OR U22568 ( .A(n18053), .B(n18054), .Z(n18052) );
  NAND U22569 ( .A(n18054), .B(n18053), .Z(n18049) );
  IV U22570 ( .A(n18055), .Z(n18054) );
  NAND U22571 ( .A(n18056), .B(n18057), .Z(n18026) );
  NANDN U22572 ( .A(n18058), .B(n18059), .Z(n18057) );
  NAND U22573 ( .A(n18060), .B(n18061), .Z(n18059) );
  OR U22574 ( .A(n18061), .B(n18060), .Z(n18056) );
  IV U22575 ( .A(n18062), .Z(n18060) );
  AND U22576 ( .A(n18063), .B(n18064), .Z(n18029) );
  NAND U22577 ( .A(n18065), .B(n18066), .Z(n18064) );
  NANDN U22578 ( .A(n18067), .B(n18068), .Z(n18066) );
  NANDN U22579 ( .A(n18068), .B(n18067), .Z(n18063) );
  XOR U22580 ( .A(n18039), .B(n18069), .Z(n18031) );
  XNOR U22581 ( .A(n18036), .B(n18038), .Z(n18069) );
  AND U22582 ( .A(n18070), .B(n18071), .Z(n18038) );
  NANDN U22583 ( .A(n18072), .B(n18073), .Z(n18071) );
  NANDN U22584 ( .A(n18074), .B(n18075), .Z(n18073) );
  IV U22585 ( .A(n18076), .Z(n18075) );
  NAND U22586 ( .A(n18076), .B(n18074), .Z(n18070) );
  AND U22587 ( .A(n18077), .B(n18078), .Z(n18036) );
  NAND U22588 ( .A(n18079), .B(n18080), .Z(n18078) );
  OR U22589 ( .A(n18081), .B(n18082), .Z(n18080) );
  NAND U22590 ( .A(n18082), .B(n18081), .Z(n18077) );
  IV U22591 ( .A(n18083), .Z(n18082) );
  NAND U22592 ( .A(n18084), .B(n18085), .Z(n18039) );
  NANDN U22593 ( .A(n18086), .B(n18087), .Z(n18085) );
  NAND U22594 ( .A(n18088), .B(n18089), .Z(n18087) );
  OR U22595 ( .A(n18089), .B(n18088), .Z(n18084) );
  IV U22596 ( .A(n18090), .Z(n18088) );
  XOR U22597 ( .A(n18065), .B(n18091), .Z(N28662) );
  XNOR U22598 ( .A(n18068), .B(n18067), .Z(n18091) );
  XNOR U22599 ( .A(n18079), .B(n18092), .Z(n18067) );
  XOR U22600 ( .A(n18083), .B(n18081), .Z(n18092) );
  XOR U22601 ( .A(n18089), .B(n18093), .Z(n18081) );
  XOR U22602 ( .A(n18086), .B(n18090), .Z(n18093) );
  NAND U22603 ( .A(n18094), .B(n18095), .Z(n18090) );
  NAND U22604 ( .A(n18096), .B(n18097), .Z(n18095) );
  NAND U22605 ( .A(n18098), .B(n18099), .Z(n18094) );
  AND U22606 ( .A(n18100), .B(n18101), .Z(n18086) );
  NAND U22607 ( .A(n18102), .B(n18103), .Z(n18101) );
  NAND U22608 ( .A(n18104), .B(n18105), .Z(n18100) );
  NANDN U22609 ( .A(n18106), .B(n18107), .Z(n18089) );
  NANDN U22610 ( .A(n18108), .B(n18109), .Z(n18083) );
  XNOR U22611 ( .A(n18074), .B(n18110), .Z(n18079) );
  XOR U22612 ( .A(n18072), .B(n18076), .Z(n18110) );
  NAND U22613 ( .A(n18111), .B(n18112), .Z(n18076) );
  NAND U22614 ( .A(n18113), .B(n18114), .Z(n18112) );
  NAND U22615 ( .A(n18115), .B(n18116), .Z(n18111) );
  AND U22616 ( .A(n18117), .B(n18118), .Z(n18072) );
  NAND U22617 ( .A(n18119), .B(n18120), .Z(n18118) );
  NAND U22618 ( .A(n18121), .B(n18122), .Z(n18117) );
  AND U22619 ( .A(n18123), .B(n18124), .Z(n18074) );
  NAND U22620 ( .A(n18125), .B(n18126), .Z(n18068) );
  XNOR U22621 ( .A(n18051), .B(n18127), .Z(n18065) );
  XOR U22622 ( .A(n18055), .B(n18053), .Z(n18127) );
  XOR U22623 ( .A(n18061), .B(n18128), .Z(n18053) );
  XOR U22624 ( .A(n18058), .B(n18062), .Z(n18128) );
  NAND U22625 ( .A(n18129), .B(n18130), .Z(n18062) );
  NAND U22626 ( .A(n18131), .B(n18132), .Z(n18130) );
  NAND U22627 ( .A(n18133), .B(n18134), .Z(n18129) );
  AND U22628 ( .A(n18135), .B(n18136), .Z(n18058) );
  NAND U22629 ( .A(n18137), .B(n18138), .Z(n18136) );
  NAND U22630 ( .A(n18139), .B(n18140), .Z(n18135) );
  NANDN U22631 ( .A(n18141), .B(n18142), .Z(n18061) );
  NANDN U22632 ( .A(n18143), .B(n18144), .Z(n18055) );
  XNOR U22633 ( .A(n18046), .B(n18145), .Z(n18051) );
  XOR U22634 ( .A(n18044), .B(n18048), .Z(n18145) );
  NAND U22635 ( .A(n18146), .B(n18147), .Z(n18048) );
  NAND U22636 ( .A(n18148), .B(n18149), .Z(n18147) );
  NAND U22637 ( .A(n18150), .B(n18151), .Z(n18146) );
  AND U22638 ( .A(n18152), .B(n18153), .Z(n18044) );
  NAND U22639 ( .A(n18154), .B(n18155), .Z(n18153) );
  NAND U22640 ( .A(n18156), .B(n18157), .Z(n18152) );
  AND U22641 ( .A(n18158), .B(n18159), .Z(n18046) );
  XOR U22642 ( .A(n18126), .B(n18125), .Z(N28661) );
  XNOR U22643 ( .A(n18144), .B(n18143), .Z(n18125) );
  XNOR U22644 ( .A(n18158), .B(n18159), .Z(n18143) );
  XOR U22645 ( .A(n18155), .B(n18154), .Z(n18159) );
  XOR U22646 ( .A(y[1467]), .B(x[1467]), .Z(n18154) );
  XOR U22647 ( .A(n18157), .B(n18156), .Z(n18155) );
  XOR U22648 ( .A(y[1469]), .B(x[1469]), .Z(n18156) );
  XOR U22649 ( .A(y[1468]), .B(x[1468]), .Z(n18157) );
  XOR U22650 ( .A(n18149), .B(n18148), .Z(n18158) );
  XOR U22651 ( .A(n18151), .B(n18150), .Z(n18148) );
  XOR U22652 ( .A(y[1466]), .B(x[1466]), .Z(n18150) );
  XOR U22653 ( .A(y[1465]), .B(x[1465]), .Z(n18151) );
  XOR U22654 ( .A(y[1464]), .B(x[1464]), .Z(n18149) );
  XNOR U22655 ( .A(n18142), .B(n18141), .Z(n18144) );
  XNOR U22656 ( .A(n18138), .B(n18137), .Z(n18141) );
  XOR U22657 ( .A(n18140), .B(n18139), .Z(n18137) );
  XOR U22658 ( .A(y[1463]), .B(x[1463]), .Z(n18139) );
  XOR U22659 ( .A(y[1462]), .B(x[1462]), .Z(n18140) );
  XOR U22660 ( .A(y[1461]), .B(x[1461]), .Z(n18138) );
  XOR U22661 ( .A(n18132), .B(n18131), .Z(n18142) );
  XOR U22662 ( .A(n18134), .B(n18133), .Z(n18131) );
  XOR U22663 ( .A(y[1460]), .B(x[1460]), .Z(n18133) );
  XOR U22664 ( .A(y[1459]), .B(x[1459]), .Z(n18134) );
  XOR U22665 ( .A(y[1458]), .B(x[1458]), .Z(n18132) );
  XNOR U22666 ( .A(n18109), .B(n18108), .Z(n18126) );
  XNOR U22667 ( .A(n18123), .B(n18124), .Z(n18108) );
  XOR U22668 ( .A(n18120), .B(n18119), .Z(n18124) );
  XOR U22669 ( .A(y[1455]), .B(x[1455]), .Z(n18119) );
  XOR U22670 ( .A(n18122), .B(n18121), .Z(n18120) );
  XOR U22671 ( .A(y[1457]), .B(x[1457]), .Z(n18121) );
  XOR U22672 ( .A(y[1456]), .B(x[1456]), .Z(n18122) );
  XOR U22673 ( .A(n18114), .B(n18113), .Z(n18123) );
  XOR U22674 ( .A(n18116), .B(n18115), .Z(n18113) );
  XOR U22675 ( .A(y[1454]), .B(x[1454]), .Z(n18115) );
  XOR U22676 ( .A(y[1453]), .B(x[1453]), .Z(n18116) );
  XOR U22677 ( .A(y[1452]), .B(x[1452]), .Z(n18114) );
  XNOR U22678 ( .A(n18107), .B(n18106), .Z(n18109) );
  XNOR U22679 ( .A(n18103), .B(n18102), .Z(n18106) );
  XOR U22680 ( .A(n18105), .B(n18104), .Z(n18102) );
  XOR U22681 ( .A(y[1451]), .B(x[1451]), .Z(n18104) );
  XOR U22682 ( .A(y[1450]), .B(x[1450]), .Z(n18105) );
  XOR U22683 ( .A(y[1449]), .B(x[1449]), .Z(n18103) );
  XOR U22684 ( .A(n18097), .B(n18096), .Z(n18107) );
  XOR U22685 ( .A(n18099), .B(n18098), .Z(n18096) );
  XOR U22686 ( .A(y[1448]), .B(x[1448]), .Z(n18098) );
  XOR U22687 ( .A(y[1447]), .B(x[1447]), .Z(n18099) );
  XOR U22688 ( .A(y[1446]), .B(x[1446]), .Z(n18097) );
  NAND U22689 ( .A(n18160), .B(n18161), .Z(N28653) );
  NAND U22690 ( .A(n18162), .B(n18163), .Z(n18161) );
  NANDN U22691 ( .A(n18164), .B(n18165), .Z(n18163) );
  NANDN U22692 ( .A(n18165), .B(n18164), .Z(n18160) );
  XOR U22693 ( .A(n18164), .B(n18166), .Z(N28652) );
  XNOR U22694 ( .A(n18162), .B(n18165), .Z(n18166) );
  NAND U22695 ( .A(n18167), .B(n18168), .Z(n18165) );
  NAND U22696 ( .A(n18169), .B(n18170), .Z(n18168) );
  NANDN U22697 ( .A(n18171), .B(n18172), .Z(n18170) );
  NANDN U22698 ( .A(n18172), .B(n18171), .Z(n18167) );
  AND U22699 ( .A(n18173), .B(n18174), .Z(n18162) );
  NAND U22700 ( .A(n18175), .B(n18176), .Z(n18174) );
  OR U22701 ( .A(n18177), .B(n18178), .Z(n18176) );
  NAND U22702 ( .A(n18178), .B(n18177), .Z(n18173) );
  IV U22703 ( .A(n18179), .Z(n18178) );
  AND U22704 ( .A(n18180), .B(n18181), .Z(n18164) );
  NAND U22705 ( .A(n18182), .B(n18183), .Z(n18181) );
  NANDN U22706 ( .A(n18184), .B(n18185), .Z(n18183) );
  NANDN U22707 ( .A(n18185), .B(n18184), .Z(n18180) );
  XOR U22708 ( .A(n18177), .B(n18186), .Z(N28651) );
  XOR U22709 ( .A(n18175), .B(n18179), .Z(n18186) );
  XNOR U22710 ( .A(n18172), .B(n18187), .Z(n18179) );
  XNOR U22711 ( .A(n18169), .B(n18171), .Z(n18187) );
  AND U22712 ( .A(n18188), .B(n18189), .Z(n18171) );
  NANDN U22713 ( .A(n18190), .B(n18191), .Z(n18189) );
  NANDN U22714 ( .A(n18192), .B(n18193), .Z(n18191) );
  IV U22715 ( .A(n18194), .Z(n18193) );
  NAND U22716 ( .A(n18194), .B(n18192), .Z(n18188) );
  AND U22717 ( .A(n18195), .B(n18196), .Z(n18169) );
  NAND U22718 ( .A(n18197), .B(n18198), .Z(n18196) );
  OR U22719 ( .A(n18199), .B(n18200), .Z(n18198) );
  NAND U22720 ( .A(n18200), .B(n18199), .Z(n18195) );
  IV U22721 ( .A(n18201), .Z(n18200) );
  NAND U22722 ( .A(n18202), .B(n18203), .Z(n18172) );
  NANDN U22723 ( .A(n18204), .B(n18205), .Z(n18203) );
  NAND U22724 ( .A(n18206), .B(n18207), .Z(n18205) );
  OR U22725 ( .A(n18207), .B(n18206), .Z(n18202) );
  IV U22726 ( .A(n18208), .Z(n18206) );
  AND U22727 ( .A(n18209), .B(n18210), .Z(n18175) );
  NAND U22728 ( .A(n18211), .B(n18212), .Z(n18210) );
  NANDN U22729 ( .A(n18213), .B(n18214), .Z(n18212) );
  NANDN U22730 ( .A(n18214), .B(n18213), .Z(n18209) );
  XOR U22731 ( .A(n18185), .B(n18215), .Z(n18177) );
  XNOR U22732 ( .A(n18182), .B(n18184), .Z(n18215) );
  AND U22733 ( .A(n18216), .B(n18217), .Z(n18184) );
  NANDN U22734 ( .A(n18218), .B(n18219), .Z(n18217) );
  NANDN U22735 ( .A(n18220), .B(n18221), .Z(n18219) );
  IV U22736 ( .A(n18222), .Z(n18221) );
  NAND U22737 ( .A(n18222), .B(n18220), .Z(n18216) );
  AND U22738 ( .A(n18223), .B(n18224), .Z(n18182) );
  NAND U22739 ( .A(n18225), .B(n18226), .Z(n18224) );
  OR U22740 ( .A(n18227), .B(n18228), .Z(n18226) );
  NAND U22741 ( .A(n18228), .B(n18227), .Z(n18223) );
  IV U22742 ( .A(n18229), .Z(n18228) );
  NAND U22743 ( .A(n18230), .B(n18231), .Z(n18185) );
  NANDN U22744 ( .A(n18232), .B(n18233), .Z(n18231) );
  NAND U22745 ( .A(n18234), .B(n18235), .Z(n18233) );
  OR U22746 ( .A(n18235), .B(n18234), .Z(n18230) );
  IV U22747 ( .A(n18236), .Z(n18234) );
  XOR U22748 ( .A(n18211), .B(n18237), .Z(N28650) );
  XNOR U22749 ( .A(n18214), .B(n18213), .Z(n18237) );
  XNOR U22750 ( .A(n18225), .B(n18238), .Z(n18213) );
  XOR U22751 ( .A(n18229), .B(n18227), .Z(n18238) );
  XOR U22752 ( .A(n18235), .B(n18239), .Z(n18227) );
  XOR U22753 ( .A(n18232), .B(n18236), .Z(n18239) );
  NAND U22754 ( .A(n18240), .B(n18241), .Z(n18236) );
  NAND U22755 ( .A(n18242), .B(n18243), .Z(n18241) );
  NAND U22756 ( .A(n18244), .B(n18245), .Z(n18240) );
  AND U22757 ( .A(n18246), .B(n18247), .Z(n18232) );
  NAND U22758 ( .A(n18248), .B(n18249), .Z(n18247) );
  NAND U22759 ( .A(n18250), .B(n18251), .Z(n18246) );
  NANDN U22760 ( .A(n18252), .B(n18253), .Z(n18235) );
  NANDN U22761 ( .A(n18254), .B(n18255), .Z(n18229) );
  XNOR U22762 ( .A(n18220), .B(n18256), .Z(n18225) );
  XOR U22763 ( .A(n18218), .B(n18222), .Z(n18256) );
  NAND U22764 ( .A(n18257), .B(n18258), .Z(n18222) );
  NAND U22765 ( .A(n18259), .B(n18260), .Z(n18258) );
  NAND U22766 ( .A(n18261), .B(n18262), .Z(n18257) );
  AND U22767 ( .A(n18263), .B(n18264), .Z(n18218) );
  NAND U22768 ( .A(n18265), .B(n18266), .Z(n18264) );
  NAND U22769 ( .A(n18267), .B(n18268), .Z(n18263) );
  AND U22770 ( .A(n18269), .B(n18270), .Z(n18220) );
  NAND U22771 ( .A(n18271), .B(n18272), .Z(n18214) );
  XNOR U22772 ( .A(n18197), .B(n18273), .Z(n18211) );
  XOR U22773 ( .A(n18201), .B(n18199), .Z(n18273) );
  XOR U22774 ( .A(n18207), .B(n18274), .Z(n18199) );
  XOR U22775 ( .A(n18204), .B(n18208), .Z(n18274) );
  NAND U22776 ( .A(n18275), .B(n18276), .Z(n18208) );
  NAND U22777 ( .A(n18277), .B(n18278), .Z(n18276) );
  NAND U22778 ( .A(n18279), .B(n18280), .Z(n18275) );
  AND U22779 ( .A(n18281), .B(n18282), .Z(n18204) );
  NAND U22780 ( .A(n18283), .B(n18284), .Z(n18282) );
  NAND U22781 ( .A(n18285), .B(n18286), .Z(n18281) );
  NANDN U22782 ( .A(n18287), .B(n18288), .Z(n18207) );
  NANDN U22783 ( .A(n18289), .B(n18290), .Z(n18201) );
  XNOR U22784 ( .A(n18192), .B(n18291), .Z(n18197) );
  XOR U22785 ( .A(n18190), .B(n18194), .Z(n18291) );
  NAND U22786 ( .A(n18292), .B(n18293), .Z(n18194) );
  NAND U22787 ( .A(n18294), .B(n18295), .Z(n18293) );
  NAND U22788 ( .A(n18296), .B(n18297), .Z(n18292) );
  AND U22789 ( .A(n18298), .B(n18299), .Z(n18190) );
  NAND U22790 ( .A(n18300), .B(n18301), .Z(n18299) );
  NAND U22791 ( .A(n18302), .B(n18303), .Z(n18298) );
  AND U22792 ( .A(n18304), .B(n18305), .Z(n18192) );
  XOR U22793 ( .A(n18272), .B(n18271), .Z(N28649) );
  XNOR U22794 ( .A(n18290), .B(n18289), .Z(n18271) );
  XNOR U22795 ( .A(n18304), .B(n18305), .Z(n18289) );
  XOR U22796 ( .A(n18301), .B(n18300), .Z(n18305) );
  XOR U22797 ( .A(y[1443]), .B(x[1443]), .Z(n18300) );
  XOR U22798 ( .A(n18303), .B(n18302), .Z(n18301) );
  XOR U22799 ( .A(y[1445]), .B(x[1445]), .Z(n18302) );
  XOR U22800 ( .A(y[1444]), .B(x[1444]), .Z(n18303) );
  XOR U22801 ( .A(n18295), .B(n18294), .Z(n18304) );
  XOR U22802 ( .A(n18297), .B(n18296), .Z(n18294) );
  XOR U22803 ( .A(y[1442]), .B(x[1442]), .Z(n18296) );
  XOR U22804 ( .A(y[1441]), .B(x[1441]), .Z(n18297) );
  XOR U22805 ( .A(y[1440]), .B(x[1440]), .Z(n18295) );
  XNOR U22806 ( .A(n18288), .B(n18287), .Z(n18290) );
  XNOR U22807 ( .A(n18284), .B(n18283), .Z(n18287) );
  XOR U22808 ( .A(n18286), .B(n18285), .Z(n18283) );
  XOR U22809 ( .A(y[1439]), .B(x[1439]), .Z(n18285) );
  XOR U22810 ( .A(y[1438]), .B(x[1438]), .Z(n18286) );
  XOR U22811 ( .A(y[1437]), .B(x[1437]), .Z(n18284) );
  XOR U22812 ( .A(n18278), .B(n18277), .Z(n18288) );
  XOR U22813 ( .A(n18280), .B(n18279), .Z(n18277) );
  XOR U22814 ( .A(y[1436]), .B(x[1436]), .Z(n18279) );
  XOR U22815 ( .A(y[1435]), .B(x[1435]), .Z(n18280) );
  XOR U22816 ( .A(y[1434]), .B(x[1434]), .Z(n18278) );
  XNOR U22817 ( .A(n18255), .B(n18254), .Z(n18272) );
  XNOR U22818 ( .A(n18269), .B(n18270), .Z(n18254) );
  XOR U22819 ( .A(n18266), .B(n18265), .Z(n18270) );
  XOR U22820 ( .A(y[1431]), .B(x[1431]), .Z(n18265) );
  XOR U22821 ( .A(n18268), .B(n18267), .Z(n18266) );
  XOR U22822 ( .A(y[1433]), .B(x[1433]), .Z(n18267) );
  XOR U22823 ( .A(y[1432]), .B(x[1432]), .Z(n18268) );
  XOR U22824 ( .A(n18260), .B(n18259), .Z(n18269) );
  XOR U22825 ( .A(n18262), .B(n18261), .Z(n18259) );
  XOR U22826 ( .A(y[1430]), .B(x[1430]), .Z(n18261) );
  XOR U22827 ( .A(y[1429]), .B(x[1429]), .Z(n18262) );
  XOR U22828 ( .A(y[1428]), .B(x[1428]), .Z(n18260) );
  XNOR U22829 ( .A(n18253), .B(n18252), .Z(n18255) );
  XNOR U22830 ( .A(n18249), .B(n18248), .Z(n18252) );
  XOR U22831 ( .A(n18251), .B(n18250), .Z(n18248) );
  XOR U22832 ( .A(y[1427]), .B(x[1427]), .Z(n18250) );
  XOR U22833 ( .A(y[1426]), .B(x[1426]), .Z(n18251) );
  XOR U22834 ( .A(y[1425]), .B(x[1425]), .Z(n18249) );
  XOR U22835 ( .A(n18243), .B(n18242), .Z(n18253) );
  XOR U22836 ( .A(n18245), .B(n18244), .Z(n18242) );
  XOR U22837 ( .A(y[1424]), .B(x[1424]), .Z(n18244) );
  XOR U22838 ( .A(y[1423]), .B(x[1423]), .Z(n18245) );
  XOR U22839 ( .A(y[1422]), .B(x[1422]), .Z(n18243) );
  NAND U22840 ( .A(n18306), .B(n18307), .Z(N28641) );
  NAND U22841 ( .A(n18308), .B(n18309), .Z(n18307) );
  NANDN U22842 ( .A(n18310), .B(n18311), .Z(n18309) );
  NANDN U22843 ( .A(n18311), .B(n18310), .Z(n18306) );
  XOR U22844 ( .A(n18310), .B(n18312), .Z(N28640) );
  XNOR U22845 ( .A(n18308), .B(n18311), .Z(n18312) );
  NAND U22846 ( .A(n18313), .B(n18314), .Z(n18311) );
  NAND U22847 ( .A(n18315), .B(n18316), .Z(n18314) );
  NANDN U22848 ( .A(n18317), .B(n18318), .Z(n18316) );
  NANDN U22849 ( .A(n18318), .B(n18317), .Z(n18313) );
  AND U22850 ( .A(n18319), .B(n18320), .Z(n18308) );
  NAND U22851 ( .A(n18321), .B(n18322), .Z(n18320) );
  OR U22852 ( .A(n18323), .B(n18324), .Z(n18322) );
  NAND U22853 ( .A(n18324), .B(n18323), .Z(n18319) );
  IV U22854 ( .A(n18325), .Z(n18324) );
  AND U22855 ( .A(n18326), .B(n18327), .Z(n18310) );
  NAND U22856 ( .A(n18328), .B(n18329), .Z(n18327) );
  NANDN U22857 ( .A(n18330), .B(n18331), .Z(n18329) );
  NANDN U22858 ( .A(n18331), .B(n18330), .Z(n18326) );
  XOR U22859 ( .A(n18323), .B(n18332), .Z(N28639) );
  XOR U22860 ( .A(n18321), .B(n18325), .Z(n18332) );
  XNOR U22861 ( .A(n18318), .B(n18333), .Z(n18325) );
  XNOR U22862 ( .A(n18315), .B(n18317), .Z(n18333) );
  AND U22863 ( .A(n18334), .B(n18335), .Z(n18317) );
  NANDN U22864 ( .A(n18336), .B(n18337), .Z(n18335) );
  NANDN U22865 ( .A(n18338), .B(n18339), .Z(n18337) );
  IV U22866 ( .A(n18340), .Z(n18339) );
  NAND U22867 ( .A(n18340), .B(n18338), .Z(n18334) );
  AND U22868 ( .A(n18341), .B(n18342), .Z(n18315) );
  NAND U22869 ( .A(n18343), .B(n18344), .Z(n18342) );
  OR U22870 ( .A(n18345), .B(n18346), .Z(n18344) );
  NAND U22871 ( .A(n18346), .B(n18345), .Z(n18341) );
  IV U22872 ( .A(n18347), .Z(n18346) );
  NAND U22873 ( .A(n18348), .B(n18349), .Z(n18318) );
  NANDN U22874 ( .A(n18350), .B(n18351), .Z(n18349) );
  NAND U22875 ( .A(n18352), .B(n18353), .Z(n18351) );
  OR U22876 ( .A(n18353), .B(n18352), .Z(n18348) );
  IV U22877 ( .A(n18354), .Z(n18352) );
  AND U22878 ( .A(n18355), .B(n18356), .Z(n18321) );
  NAND U22879 ( .A(n18357), .B(n18358), .Z(n18356) );
  NANDN U22880 ( .A(n18359), .B(n18360), .Z(n18358) );
  NANDN U22881 ( .A(n18360), .B(n18359), .Z(n18355) );
  XOR U22882 ( .A(n18331), .B(n18361), .Z(n18323) );
  XNOR U22883 ( .A(n18328), .B(n18330), .Z(n18361) );
  AND U22884 ( .A(n18362), .B(n18363), .Z(n18330) );
  NANDN U22885 ( .A(n18364), .B(n18365), .Z(n18363) );
  NANDN U22886 ( .A(n18366), .B(n18367), .Z(n18365) );
  IV U22887 ( .A(n18368), .Z(n18367) );
  NAND U22888 ( .A(n18368), .B(n18366), .Z(n18362) );
  AND U22889 ( .A(n18369), .B(n18370), .Z(n18328) );
  NAND U22890 ( .A(n18371), .B(n18372), .Z(n18370) );
  OR U22891 ( .A(n18373), .B(n18374), .Z(n18372) );
  NAND U22892 ( .A(n18374), .B(n18373), .Z(n18369) );
  IV U22893 ( .A(n18375), .Z(n18374) );
  NAND U22894 ( .A(n18376), .B(n18377), .Z(n18331) );
  NANDN U22895 ( .A(n18378), .B(n18379), .Z(n18377) );
  NAND U22896 ( .A(n18380), .B(n18381), .Z(n18379) );
  OR U22897 ( .A(n18381), .B(n18380), .Z(n18376) );
  IV U22898 ( .A(n18382), .Z(n18380) );
  XOR U22899 ( .A(n18357), .B(n18383), .Z(N28638) );
  XNOR U22900 ( .A(n18360), .B(n18359), .Z(n18383) );
  XNOR U22901 ( .A(n18371), .B(n18384), .Z(n18359) );
  XOR U22902 ( .A(n18375), .B(n18373), .Z(n18384) );
  XOR U22903 ( .A(n18381), .B(n18385), .Z(n18373) );
  XOR U22904 ( .A(n18378), .B(n18382), .Z(n18385) );
  NAND U22905 ( .A(n18386), .B(n18387), .Z(n18382) );
  NAND U22906 ( .A(n18388), .B(n18389), .Z(n18387) );
  NAND U22907 ( .A(n18390), .B(n18391), .Z(n18386) );
  AND U22908 ( .A(n18392), .B(n18393), .Z(n18378) );
  NAND U22909 ( .A(n18394), .B(n18395), .Z(n18393) );
  NAND U22910 ( .A(n18396), .B(n18397), .Z(n18392) );
  NANDN U22911 ( .A(n18398), .B(n18399), .Z(n18381) );
  NANDN U22912 ( .A(n18400), .B(n18401), .Z(n18375) );
  XNOR U22913 ( .A(n18366), .B(n18402), .Z(n18371) );
  XOR U22914 ( .A(n18364), .B(n18368), .Z(n18402) );
  NAND U22915 ( .A(n18403), .B(n18404), .Z(n18368) );
  NAND U22916 ( .A(n18405), .B(n18406), .Z(n18404) );
  NAND U22917 ( .A(n18407), .B(n18408), .Z(n18403) );
  AND U22918 ( .A(n18409), .B(n18410), .Z(n18364) );
  NAND U22919 ( .A(n18411), .B(n18412), .Z(n18410) );
  NAND U22920 ( .A(n18413), .B(n18414), .Z(n18409) );
  AND U22921 ( .A(n18415), .B(n18416), .Z(n18366) );
  NAND U22922 ( .A(n18417), .B(n18418), .Z(n18360) );
  XNOR U22923 ( .A(n18343), .B(n18419), .Z(n18357) );
  XOR U22924 ( .A(n18347), .B(n18345), .Z(n18419) );
  XOR U22925 ( .A(n18353), .B(n18420), .Z(n18345) );
  XOR U22926 ( .A(n18350), .B(n18354), .Z(n18420) );
  NAND U22927 ( .A(n18421), .B(n18422), .Z(n18354) );
  NAND U22928 ( .A(n18423), .B(n18424), .Z(n18422) );
  NAND U22929 ( .A(n18425), .B(n18426), .Z(n18421) );
  AND U22930 ( .A(n18427), .B(n18428), .Z(n18350) );
  NAND U22931 ( .A(n18429), .B(n18430), .Z(n18428) );
  NAND U22932 ( .A(n18431), .B(n18432), .Z(n18427) );
  NANDN U22933 ( .A(n18433), .B(n18434), .Z(n18353) );
  NANDN U22934 ( .A(n18435), .B(n18436), .Z(n18347) );
  XNOR U22935 ( .A(n18338), .B(n18437), .Z(n18343) );
  XOR U22936 ( .A(n18336), .B(n18340), .Z(n18437) );
  NAND U22937 ( .A(n18438), .B(n18439), .Z(n18340) );
  NAND U22938 ( .A(n18440), .B(n18441), .Z(n18439) );
  NAND U22939 ( .A(n18442), .B(n18443), .Z(n18438) );
  AND U22940 ( .A(n18444), .B(n18445), .Z(n18336) );
  NAND U22941 ( .A(n18446), .B(n18447), .Z(n18445) );
  NAND U22942 ( .A(n18448), .B(n18449), .Z(n18444) );
  AND U22943 ( .A(n18450), .B(n18451), .Z(n18338) );
  XOR U22944 ( .A(n18418), .B(n18417), .Z(N28637) );
  XNOR U22945 ( .A(n18436), .B(n18435), .Z(n18417) );
  XNOR U22946 ( .A(n18450), .B(n18451), .Z(n18435) );
  XOR U22947 ( .A(n18447), .B(n18446), .Z(n18451) );
  XOR U22948 ( .A(y[1419]), .B(x[1419]), .Z(n18446) );
  XOR U22949 ( .A(n18449), .B(n18448), .Z(n18447) );
  XOR U22950 ( .A(y[1421]), .B(x[1421]), .Z(n18448) );
  XOR U22951 ( .A(y[1420]), .B(x[1420]), .Z(n18449) );
  XOR U22952 ( .A(n18441), .B(n18440), .Z(n18450) );
  XOR U22953 ( .A(n18443), .B(n18442), .Z(n18440) );
  XOR U22954 ( .A(y[1418]), .B(x[1418]), .Z(n18442) );
  XOR U22955 ( .A(y[1417]), .B(x[1417]), .Z(n18443) );
  XOR U22956 ( .A(y[1416]), .B(x[1416]), .Z(n18441) );
  XNOR U22957 ( .A(n18434), .B(n18433), .Z(n18436) );
  XNOR U22958 ( .A(n18430), .B(n18429), .Z(n18433) );
  XOR U22959 ( .A(n18432), .B(n18431), .Z(n18429) );
  XOR U22960 ( .A(y[1415]), .B(x[1415]), .Z(n18431) );
  XOR U22961 ( .A(y[1414]), .B(x[1414]), .Z(n18432) );
  XOR U22962 ( .A(y[1413]), .B(x[1413]), .Z(n18430) );
  XOR U22963 ( .A(n18424), .B(n18423), .Z(n18434) );
  XOR U22964 ( .A(n18426), .B(n18425), .Z(n18423) );
  XOR U22965 ( .A(y[1412]), .B(x[1412]), .Z(n18425) );
  XOR U22966 ( .A(y[1411]), .B(x[1411]), .Z(n18426) );
  XOR U22967 ( .A(y[1410]), .B(x[1410]), .Z(n18424) );
  XNOR U22968 ( .A(n18401), .B(n18400), .Z(n18418) );
  XNOR U22969 ( .A(n18415), .B(n18416), .Z(n18400) );
  XOR U22970 ( .A(n18412), .B(n18411), .Z(n18416) );
  XOR U22971 ( .A(y[1407]), .B(x[1407]), .Z(n18411) );
  XOR U22972 ( .A(n18414), .B(n18413), .Z(n18412) );
  XOR U22973 ( .A(y[1409]), .B(x[1409]), .Z(n18413) );
  XOR U22974 ( .A(y[1408]), .B(x[1408]), .Z(n18414) );
  XOR U22975 ( .A(n18406), .B(n18405), .Z(n18415) );
  XOR U22976 ( .A(n18408), .B(n18407), .Z(n18405) );
  XOR U22977 ( .A(y[1406]), .B(x[1406]), .Z(n18407) );
  XOR U22978 ( .A(y[1405]), .B(x[1405]), .Z(n18408) );
  XOR U22979 ( .A(y[1404]), .B(x[1404]), .Z(n18406) );
  XNOR U22980 ( .A(n18399), .B(n18398), .Z(n18401) );
  XNOR U22981 ( .A(n18395), .B(n18394), .Z(n18398) );
  XOR U22982 ( .A(n18397), .B(n18396), .Z(n18394) );
  XOR U22983 ( .A(y[1403]), .B(x[1403]), .Z(n18396) );
  XOR U22984 ( .A(y[1402]), .B(x[1402]), .Z(n18397) );
  XOR U22985 ( .A(y[1401]), .B(x[1401]), .Z(n18395) );
  XOR U22986 ( .A(n18389), .B(n18388), .Z(n18399) );
  XOR U22987 ( .A(n18391), .B(n18390), .Z(n18388) );
  XOR U22988 ( .A(y[1400]), .B(x[1400]), .Z(n18390) );
  XOR U22989 ( .A(y[1399]), .B(x[1399]), .Z(n18391) );
  XOR U22990 ( .A(y[1398]), .B(x[1398]), .Z(n18389) );
  NAND U22991 ( .A(n18452), .B(n18453), .Z(N28629) );
  NAND U22992 ( .A(n18454), .B(n18455), .Z(n18453) );
  NANDN U22993 ( .A(n18456), .B(n18457), .Z(n18455) );
  NANDN U22994 ( .A(n18457), .B(n18456), .Z(n18452) );
  XOR U22995 ( .A(n18456), .B(n18458), .Z(N28628) );
  XNOR U22996 ( .A(n18454), .B(n18457), .Z(n18458) );
  NAND U22997 ( .A(n18459), .B(n18460), .Z(n18457) );
  NAND U22998 ( .A(n18461), .B(n18462), .Z(n18460) );
  NANDN U22999 ( .A(n18463), .B(n18464), .Z(n18462) );
  NANDN U23000 ( .A(n18464), .B(n18463), .Z(n18459) );
  AND U23001 ( .A(n18465), .B(n18466), .Z(n18454) );
  NAND U23002 ( .A(n18467), .B(n18468), .Z(n18466) );
  OR U23003 ( .A(n18469), .B(n18470), .Z(n18468) );
  NAND U23004 ( .A(n18470), .B(n18469), .Z(n18465) );
  IV U23005 ( .A(n18471), .Z(n18470) );
  AND U23006 ( .A(n18472), .B(n18473), .Z(n18456) );
  NAND U23007 ( .A(n18474), .B(n18475), .Z(n18473) );
  NANDN U23008 ( .A(n18476), .B(n18477), .Z(n18475) );
  NANDN U23009 ( .A(n18477), .B(n18476), .Z(n18472) );
  XOR U23010 ( .A(n18469), .B(n18478), .Z(N28627) );
  XOR U23011 ( .A(n18467), .B(n18471), .Z(n18478) );
  XNOR U23012 ( .A(n18464), .B(n18479), .Z(n18471) );
  XNOR U23013 ( .A(n18461), .B(n18463), .Z(n18479) );
  AND U23014 ( .A(n18480), .B(n18481), .Z(n18463) );
  NANDN U23015 ( .A(n18482), .B(n18483), .Z(n18481) );
  NANDN U23016 ( .A(n18484), .B(n18485), .Z(n18483) );
  IV U23017 ( .A(n18486), .Z(n18485) );
  NAND U23018 ( .A(n18486), .B(n18484), .Z(n18480) );
  AND U23019 ( .A(n18487), .B(n18488), .Z(n18461) );
  NAND U23020 ( .A(n18489), .B(n18490), .Z(n18488) );
  OR U23021 ( .A(n18491), .B(n18492), .Z(n18490) );
  NAND U23022 ( .A(n18492), .B(n18491), .Z(n18487) );
  IV U23023 ( .A(n18493), .Z(n18492) );
  NAND U23024 ( .A(n18494), .B(n18495), .Z(n18464) );
  NANDN U23025 ( .A(n18496), .B(n18497), .Z(n18495) );
  NAND U23026 ( .A(n18498), .B(n18499), .Z(n18497) );
  OR U23027 ( .A(n18499), .B(n18498), .Z(n18494) );
  IV U23028 ( .A(n18500), .Z(n18498) );
  AND U23029 ( .A(n18501), .B(n18502), .Z(n18467) );
  NAND U23030 ( .A(n18503), .B(n18504), .Z(n18502) );
  NANDN U23031 ( .A(n18505), .B(n18506), .Z(n18504) );
  NANDN U23032 ( .A(n18506), .B(n18505), .Z(n18501) );
  XOR U23033 ( .A(n18477), .B(n18507), .Z(n18469) );
  XNOR U23034 ( .A(n18474), .B(n18476), .Z(n18507) );
  AND U23035 ( .A(n18508), .B(n18509), .Z(n18476) );
  NANDN U23036 ( .A(n18510), .B(n18511), .Z(n18509) );
  NANDN U23037 ( .A(n18512), .B(n18513), .Z(n18511) );
  IV U23038 ( .A(n18514), .Z(n18513) );
  NAND U23039 ( .A(n18514), .B(n18512), .Z(n18508) );
  AND U23040 ( .A(n18515), .B(n18516), .Z(n18474) );
  NAND U23041 ( .A(n18517), .B(n18518), .Z(n18516) );
  OR U23042 ( .A(n18519), .B(n18520), .Z(n18518) );
  NAND U23043 ( .A(n18520), .B(n18519), .Z(n18515) );
  IV U23044 ( .A(n18521), .Z(n18520) );
  NAND U23045 ( .A(n18522), .B(n18523), .Z(n18477) );
  NANDN U23046 ( .A(n18524), .B(n18525), .Z(n18523) );
  NAND U23047 ( .A(n18526), .B(n18527), .Z(n18525) );
  OR U23048 ( .A(n18527), .B(n18526), .Z(n18522) );
  IV U23049 ( .A(n18528), .Z(n18526) );
  XOR U23050 ( .A(n18503), .B(n18529), .Z(N28626) );
  XNOR U23051 ( .A(n18506), .B(n18505), .Z(n18529) );
  XNOR U23052 ( .A(n18517), .B(n18530), .Z(n18505) );
  XOR U23053 ( .A(n18521), .B(n18519), .Z(n18530) );
  XOR U23054 ( .A(n18527), .B(n18531), .Z(n18519) );
  XOR U23055 ( .A(n18524), .B(n18528), .Z(n18531) );
  NAND U23056 ( .A(n18532), .B(n18533), .Z(n18528) );
  NAND U23057 ( .A(n18534), .B(n18535), .Z(n18533) );
  NAND U23058 ( .A(n18536), .B(n18537), .Z(n18532) );
  AND U23059 ( .A(n18538), .B(n18539), .Z(n18524) );
  NAND U23060 ( .A(n18540), .B(n18541), .Z(n18539) );
  NAND U23061 ( .A(n18542), .B(n18543), .Z(n18538) );
  NANDN U23062 ( .A(n18544), .B(n18545), .Z(n18527) );
  NANDN U23063 ( .A(n18546), .B(n18547), .Z(n18521) );
  XNOR U23064 ( .A(n18512), .B(n18548), .Z(n18517) );
  XOR U23065 ( .A(n18510), .B(n18514), .Z(n18548) );
  NAND U23066 ( .A(n18549), .B(n18550), .Z(n18514) );
  NAND U23067 ( .A(n18551), .B(n18552), .Z(n18550) );
  NAND U23068 ( .A(n18553), .B(n18554), .Z(n18549) );
  AND U23069 ( .A(n18555), .B(n18556), .Z(n18510) );
  NAND U23070 ( .A(n18557), .B(n18558), .Z(n18556) );
  NAND U23071 ( .A(n18559), .B(n18560), .Z(n18555) );
  AND U23072 ( .A(n18561), .B(n18562), .Z(n18512) );
  NAND U23073 ( .A(n18563), .B(n18564), .Z(n18506) );
  XNOR U23074 ( .A(n18489), .B(n18565), .Z(n18503) );
  XOR U23075 ( .A(n18493), .B(n18491), .Z(n18565) );
  XOR U23076 ( .A(n18499), .B(n18566), .Z(n18491) );
  XOR U23077 ( .A(n18496), .B(n18500), .Z(n18566) );
  NAND U23078 ( .A(n18567), .B(n18568), .Z(n18500) );
  NAND U23079 ( .A(n18569), .B(n18570), .Z(n18568) );
  NAND U23080 ( .A(n18571), .B(n18572), .Z(n18567) );
  AND U23081 ( .A(n18573), .B(n18574), .Z(n18496) );
  NAND U23082 ( .A(n18575), .B(n18576), .Z(n18574) );
  NAND U23083 ( .A(n18577), .B(n18578), .Z(n18573) );
  NANDN U23084 ( .A(n18579), .B(n18580), .Z(n18499) );
  NANDN U23085 ( .A(n18581), .B(n18582), .Z(n18493) );
  XNOR U23086 ( .A(n18484), .B(n18583), .Z(n18489) );
  XOR U23087 ( .A(n18482), .B(n18486), .Z(n18583) );
  NAND U23088 ( .A(n18584), .B(n18585), .Z(n18486) );
  NAND U23089 ( .A(n18586), .B(n18587), .Z(n18585) );
  NAND U23090 ( .A(n18588), .B(n18589), .Z(n18584) );
  AND U23091 ( .A(n18590), .B(n18591), .Z(n18482) );
  NAND U23092 ( .A(n18592), .B(n18593), .Z(n18591) );
  NAND U23093 ( .A(n18594), .B(n18595), .Z(n18590) );
  AND U23094 ( .A(n18596), .B(n18597), .Z(n18484) );
  XOR U23095 ( .A(n18564), .B(n18563), .Z(N28625) );
  XNOR U23096 ( .A(n18582), .B(n18581), .Z(n18563) );
  XNOR U23097 ( .A(n18596), .B(n18597), .Z(n18581) );
  XOR U23098 ( .A(n18593), .B(n18592), .Z(n18597) );
  XOR U23099 ( .A(y[1395]), .B(x[1395]), .Z(n18592) );
  XOR U23100 ( .A(n18595), .B(n18594), .Z(n18593) );
  XOR U23101 ( .A(y[1397]), .B(x[1397]), .Z(n18594) );
  XOR U23102 ( .A(y[1396]), .B(x[1396]), .Z(n18595) );
  XOR U23103 ( .A(n18587), .B(n18586), .Z(n18596) );
  XOR U23104 ( .A(n18589), .B(n18588), .Z(n18586) );
  XOR U23105 ( .A(y[1394]), .B(x[1394]), .Z(n18588) );
  XOR U23106 ( .A(y[1393]), .B(x[1393]), .Z(n18589) );
  XOR U23107 ( .A(y[1392]), .B(x[1392]), .Z(n18587) );
  XNOR U23108 ( .A(n18580), .B(n18579), .Z(n18582) );
  XNOR U23109 ( .A(n18576), .B(n18575), .Z(n18579) );
  XOR U23110 ( .A(n18578), .B(n18577), .Z(n18575) );
  XOR U23111 ( .A(y[1391]), .B(x[1391]), .Z(n18577) );
  XOR U23112 ( .A(y[1390]), .B(x[1390]), .Z(n18578) );
  XOR U23113 ( .A(y[1389]), .B(x[1389]), .Z(n18576) );
  XOR U23114 ( .A(n18570), .B(n18569), .Z(n18580) );
  XOR U23115 ( .A(n18572), .B(n18571), .Z(n18569) );
  XOR U23116 ( .A(y[1388]), .B(x[1388]), .Z(n18571) );
  XOR U23117 ( .A(y[1387]), .B(x[1387]), .Z(n18572) );
  XOR U23118 ( .A(y[1386]), .B(x[1386]), .Z(n18570) );
  XNOR U23119 ( .A(n18547), .B(n18546), .Z(n18564) );
  XNOR U23120 ( .A(n18561), .B(n18562), .Z(n18546) );
  XOR U23121 ( .A(n18558), .B(n18557), .Z(n18562) );
  XOR U23122 ( .A(y[1383]), .B(x[1383]), .Z(n18557) );
  XOR U23123 ( .A(n18560), .B(n18559), .Z(n18558) );
  XOR U23124 ( .A(y[1385]), .B(x[1385]), .Z(n18559) );
  XOR U23125 ( .A(y[1384]), .B(x[1384]), .Z(n18560) );
  XOR U23126 ( .A(n18552), .B(n18551), .Z(n18561) );
  XOR U23127 ( .A(n18554), .B(n18553), .Z(n18551) );
  XOR U23128 ( .A(y[1382]), .B(x[1382]), .Z(n18553) );
  XOR U23129 ( .A(y[1381]), .B(x[1381]), .Z(n18554) );
  XOR U23130 ( .A(y[1380]), .B(x[1380]), .Z(n18552) );
  XNOR U23131 ( .A(n18545), .B(n18544), .Z(n18547) );
  XNOR U23132 ( .A(n18541), .B(n18540), .Z(n18544) );
  XOR U23133 ( .A(n18543), .B(n18542), .Z(n18540) );
  XOR U23134 ( .A(y[1379]), .B(x[1379]), .Z(n18542) );
  XOR U23135 ( .A(y[1378]), .B(x[1378]), .Z(n18543) );
  XOR U23136 ( .A(y[1377]), .B(x[1377]), .Z(n18541) );
  XOR U23137 ( .A(n18535), .B(n18534), .Z(n18545) );
  XOR U23138 ( .A(n18537), .B(n18536), .Z(n18534) );
  XOR U23139 ( .A(y[1376]), .B(x[1376]), .Z(n18536) );
  XOR U23140 ( .A(y[1375]), .B(x[1375]), .Z(n18537) );
  XOR U23141 ( .A(y[1374]), .B(x[1374]), .Z(n18535) );
  NAND U23142 ( .A(n18598), .B(n18599), .Z(N28617) );
  NAND U23143 ( .A(n18600), .B(n18601), .Z(n18599) );
  NANDN U23144 ( .A(n18602), .B(n18603), .Z(n18601) );
  NANDN U23145 ( .A(n18603), .B(n18602), .Z(n18598) );
  XOR U23146 ( .A(n18602), .B(n18604), .Z(N28616) );
  XNOR U23147 ( .A(n18600), .B(n18603), .Z(n18604) );
  NAND U23148 ( .A(n18605), .B(n18606), .Z(n18603) );
  NAND U23149 ( .A(n18607), .B(n18608), .Z(n18606) );
  NANDN U23150 ( .A(n18609), .B(n18610), .Z(n18608) );
  NANDN U23151 ( .A(n18610), .B(n18609), .Z(n18605) );
  AND U23152 ( .A(n18611), .B(n18612), .Z(n18600) );
  NAND U23153 ( .A(n18613), .B(n18614), .Z(n18612) );
  OR U23154 ( .A(n18615), .B(n18616), .Z(n18614) );
  NAND U23155 ( .A(n18616), .B(n18615), .Z(n18611) );
  IV U23156 ( .A(n18617), .Z(n18616) );
  AND U23157 ( .A(n18618), .B(n18619), .Z(n18602) );
  NAND U23158 ( .A(n18620), .B(n18621), .Z(n18619) );
  NANDN U23159 ( .A(n18622), .B(n18623), .Z(n18621) );
  NANDN U23160 ( .A(n18623), .B(n18622), .Z(n18618) );
  XOR U23161 ( .A(n18615), .B(n18624), .Z(N28615) );
  XOR U23162 ( .A(n18613), .B(n18617), .Z(n18624) );
  XNOR U23163 ( .A(n18610), .B(n18625), .Z(n18617) );
  XNOR U23164 ( .A(n18607), .B(n18609), .Z(n18625) );
  AND U23165 ( .A(n18626), .B(n18627), .Z(n18609) );
  NANDN U23166 ( .A(n18628), .B(n18629), .Z(n18627) );
  NANDN U23167 ( .A(n18630), .B(n18631), .Z(n18629) );
  IV U23168 ( .A(n18632), .Z(n18631) );
  NAND U23169 ( .A(n18632), .B(n18630), .Z(n18626) );
  AND U23170 ( .A(n18633), .B(n18634), .Z(n18607) );
  NAND U23171 ( .A(n18635), .B(n18636), .Z(n18634) );
  OR U23172 ( .A(n18637), .B(n18638), .Z(n18636) );
  NAND U23173 ( .A(n18638), .B(n18637), .Z(n18633) );
  IV U23174 ( .A(n18639), .Z(n18638) );
  NAND U23175 ( .A(n18640), .B(n18641), .Z(n18610) );
  NANDN U23176 ( .A(n18642), .B(n18643), .Z(n18641) );
  NAND U23177 ( .A(n18644), .B(n18645), .Z(n18643) );
  OR U23178 ( .A(n18645), .B(n18644), .Z(n18640) );
  IV U23179 ( .A(n18646), .Z(n18644) );
  AND U23180 ( .A(n18647), .B(n18648), .Z(n18613) );
  NAND U23181 ( .A(n18649), .B(n18650), .Z(n18648) );
  NANDN U23182 ( .A(n18651), .B(n18652), .Z(n18650) );
  NANDN U23183 ( .A(n18652), .B(n18651), .Z(n18647) );
  XOR U23184 ( .A(n18623), .B(n18653), .Z(n18615) );
  XNOR U23185 ( .A(n18620), .B(n18622), .Z(n18653) );
  AND U23186 ( .A(n18654), .B(n18655), .Z(n18622) );
  NANDN U23187 ( .A(n18656), .B(n18657), .Z(n18655) );
  NANDN U23188 ( .A(n18658), .B(n18659), .Z(n18657) );
  IV U23189 ( .A(n18660), .Z(n18659) );
  NAND U23190 ( .A(n18660), .B(n18658), .Z(n18654) );
  AND U23191 ( .A(n18661), .B(n18662), .Z(n18620) );
  NAND U23192 ( .A(n18663), .B(n18664), .Z(n18662) );
  OR U23193 ( .A(n18665), .B(n18666), .Z(n18664) );
  NAND U23194 ( .A(n18666), .B(n18665), .Z(n18661) );
  IV U23195 ( .A(n18667), .Z(n18666) );
  NAND U23196 ( .A(n18668), .B(n18669), .Z(n18623) );
  NANDN U23197 ( .A(n18670), .B(n18671), .Z(n18669) );
  NAND U23198 ( .A(n18672), .B(n18673), .Z(n18671) );
  OR U23199 ( .A(n18673), .B(n18672), .Z(n18668) );
  IV U23200 ( .A(n18674), .Z(n18672) );
  XOR U23201 ( .A(n18649), .B(n18675), .Z(N28614) );
  XNOR U23202 ( .A(n18652), .B(n18651), .Z(n18675) );
  XNOR U23203 ( .A(n18663), .B(n18676), .Z(n18651) );
  XOR U23204 ( .A(n18667), .B(n18665), .Z(n18676) );
  XOR U23205 ( .A(n18673), .B(n18677), .Z(n18665) );
  XOR U23206 ( .A(n18670), .B(n18674), .Z(n18677) );
  NAND U23207 ( .A(n18678), .B(n18679), .Z(n18674) );
  NAND U23208 ( .A(n18680), .B(n18681), .Z(n18679) );
  NAND U23209 ( .A(n18682), .B(n18683), .Z(n18678) );
  AND U23210 ( .A(n18684), .B(n18685), .Z(n18670) );
  NAND U23211 ( .A(n18686), .B(n18687), .Z(n18685) );
  NAND U23212 ( .A(n18688), .B(n18689), .Z(n18684) );
  NANDN U23213 ( .A(n18690), .B(n18691), .Z(n18673) );
  NANDN U23214 ( .A(n18692), .B(n18693), .Z(n18667) );
  XNOR U23215 ( .A(n18658), .B(n18694), .Z(n18663) );
  XOR U23216 ( .A(n18656), .B(n18660), .Z(n18694) );
  NAND U23217 ( .A(n18695), .B(n18696), .Z(n18660) );
  NAND U23218 ( .A(n18697), .B(n18698), .Z(n18696) );
  NAND U23219 ( .A(n18699), .B(n18700), .Z(n18695) );
  AND U23220 ( .A(n18701), .B(n18702), .Z(n18656) );
  NAND U23221 ( .A(n18703), .B(n18704), .Z(n18702) );
  NAND U23222 ( .A(n18705), .B(n18706), .Z(n18701) );
  AND U23223 ( .A(n18707), .B(n18708), .Z(n18658) );
  NAND U23224 ( .A(n18709), .B(n18710), .Z(n18652) );
  XNOR U23225 ( .A(n18635), .B(n18711), .Z(n18649) );
  XOR U23226 ( .A(n18639), .B(n18637), .Z(n18711) );
  XOR U23227 ( .A(n18645), .B(n18712), .Z(n18637) );
  XOR U23228 ( .A(n18642), .B(n18646), .Z(n18712) );
  NAND U23229 ( .A(n18713), .B(n18714), .Z(n18646) );
  NAND U23230 ( .A(n18715), .B(n18716), .Z(n18714) );
  NAND U23231 ( .A(n18717), .B(n18718), .Z(n18713) );
  AND U23232 ( .A(n18719), .B(n18720), .Z(n18642) );
  NAND U23233 ( .A(n18721), .B(n18722), .Z(n18720) );
  NAND U23234 ( .A(n18723), .B(n18724), .Z(n18719) );
  NANDN U23235 ( .A(n18725), .B(n18726), .Z(n18645) );
  NANDN U23236 ( .A(n18727), .B(n18728), .Z(n18639) );
  XNOR U23237 ( .A(n18630), .B(n18729), .Z(n18635) );
  XOR U23238 ( .A(n18628), .B(n18632), .Z(n18729) );
  NAND U23239 ( .A(n18730), .B(n18731), .Z(n18632) );
  NAND U23240 ( .A(n18732), .B(n18733), .Z(n18731) );
  NAND U23241 ( .A(n18734), .B(n18735), .Z(n18730) );
  AND U23242 ( .A(n18736), .B(n18737), .Z(n18628) );
  NAND U23243 ( .A(n18738), .B(n18739), .Z(n18737) );
  NAND U23244 ( .A(n18740), .B(n18741), .Z(n18736) );
  AND U23245 ( .A(n18742), .B(n18743), .Z(n18630) );
  XOR U23246 ( .A(n18710), .B(n18709), .Z(N28613) );
  XNOR U23247 ( .A(n18728), .B(n18727), .Z(n18709) );
  XNOR U23248 ( .A(n18742), .B(n18743), .Z(n18727) );
  XOR U23249 ( .A(n18739), .B(n18738), .Z(n18743) );
  XOR U23250 ( .A(y[1371]), .B(x[1371]), .Z(n18738) );
  XOR U23251 ( .A(n18741), .B(n18740), .Z(n18739) );
  XOR U23252 ( .A(y[1373]), .B(x[1373]), .Z(n18740) );
  XOR U23253 ( .A(y[1372]), .B(x[1372]), .Z(n18741) );
  XOR U23254 ( .A(n18733), .B(n18732), .Z(n18742) );
  XOR U23255 ( .A(n18735), .B(n18734), .Z(n18732) );
  XOR U23256 ( .A(y[1370]), .B(x[1370]), .Z(n18734) );
  XOR U23257 ( .A(y[1369]), .B(x[1369]), .Z(n18735) );
  XOR U23258 ( .A(y[1368]), .B(x[1368]), .Z(n18733) );
  XNOR U23259 ( .A(n18726), .B(n18725), .Z(n18728) );
  XNOR U23260 ( .A(n18722), .B(n18721), .Z(n18725) );
  XOR U23261 ( .A(n18724), .B(n18723), .Z(n18721) );
  XOR U23262 ( .A(y[1367]), .B(x[1367]), .Z(n18723) );
  XOR U23263 ( .A(y[1366]), .B(x[1366]), .Z(n18724) );
  XOR U23264 ( .A(y[1365]), .B(x[1365]), .Z(n18722) );
  XOR U23265 ( .A(n18716), .B(n18715), .Z(n18726) );
  XOR U23266 ( .A(n18718), .B(n18717), .Z(n18715) );
  XOR U23267 ( .A(y[1364]), .B(x[1364]), .Z(n18717) );
  XOR U23268 ( .A(y[1363]), .B(x[1363]), .Z(n18718) );
  XOR U23269 ( .A(y[1362]), .B(x[1362]), .Z(n18716) );
  XNOR U23270 ( .A(n18693), .B(n18692), .Z(n18710) );
  XNOR U23271 ( .A(n18707), .B(n18708), .Z(n18692) );
  XOR U23272 ( .A(n18704), .B(n18703), .Z(n18708) );
  XOR U23273 ( .A(y[1359]), .B(x[1359]), .Z(n18703) );
  XOR U23274 ( .A(n18706), .B(n18705), .Z(n18704) );
  XOR U23275 ( .A(y[1361]), .B(x[1361]), .Z(n18705) );
  XOR U23276 ( .A(y[1360]), .B(x[1360]), .Z(n18706) );
  XOR U23277 ( .A(n18698), .B(n18697), .Z(n18707) );
  XOR U23278 ( .A(n18700), .B(n18699), .Z(n18697) );
  XOR U23279 ( .A(y[1358]), .B(x[1358]), .Z(n18699) );
  XOR U23280 ( .A(y[1357]), .B(x[1357]), .Z(n18700) );
  XOR U23281 ( .A(y[1356]), .B(x[1356]), .Z(n18698) );
  XNOR U23282 ( .A(n18691), .B(n18690), .Z(n18693) );
  XNOR U23283 ( .A(n18687), .B(n18686), .Z(n18690) );
  XOR U23284 ( .A(n18689), .B(n18688), .Z(n18686) );
  XOR U23285 ( .A(y[1355]), .B(x[1355]), .Z(n18688) );
  XOR U23286 ( .A(y[1354]), .B(x[1354]), .Z(n18689) );
  XOR U23287 ( .A(y[1353]), .B(x[1353]), .Z(n18687) );
  XOR U23288 ( .A(n18681), .B(n18680), .Z(n18691) );
  XOR U23289 ( .A(n18683), .B(n18682), .Z(n18680) );
  XOR U23290 ( .A(y[1352]), .B(x[1352]), .Z(n18682) );
  XOR U23291 ( .A(y[1351]), .B(x[1351]), .Z(n18683) );
  XOR U23292 ( .A(y[1350]), .B(x[1350]), .Z(n18681) );
  NAND U23293 ( .A(n18744), .B(n18745), .Z(N28605) );
  NAND U23294 ( .A(n18746), .B(n18747), .Z(n18745) );
  NANDN U23295 ( .A(n18748), .B(n18749), .Z(n18747) );
  NANDN U23296 ( .A(n18749), .B(n18748), .Z(n18744) );
  XOR U23297 ( .A(n18748), .B(n18750), .Z(N28604) );
  XNOR U23298 ( .A(n18746), .B(n18749), .Z(n18750) );
  NAND U23299 ( .A(n18751), .B(n18752), .Z(n18749) );
  NAND U23300 ( .A(n18753), .B(n18754), .Z(n18752) );
  NANDN U23301 ( .A(n18755), .B(n18756), .Z(n18754) );
  NANDN U23302 ( .A(n18756), .B(n18755), .Z(n18751) );
  AND U23303 ( .A(n18757), .B(n18758), .Z(n18746) );
  NAND U23304 ( .A(n18759), .B(n18760), .Z(n18758) );
  OR U23305 ( .A(n18761), .B(n18762), .Z(n18760) );
  NAND U23306 ( .A(n18762), .B(n18761), .Z(n18757) );
  IV U23307 ( .A(n18763), .Z(n18762) );
  AND U23308 ( .A(n18764), .B(n18765), .Z(n18748) );
  NAND U23309 ( .A(n18766), .B(n18767), .Z(n18765) );
  NANDN U23310 ( .A(n18768), .B(n18769), .Z(n18767) );
  NANDN U23311 ( .A(n18769), .B(n18768), .Z(n18764) );
  XOR U23312 ( .A(n18761), .B(n18770), .Z(N28603) );
  XOR U23313 ( .A(n18759), .B(n18763), .Z(n18770) );
  XNOR U23314 ( .A(n18756), .B(n18771), .Z(n18763) );
  XNOR U23315 ( .A(n18753), .B(n18755), .Z(n18771) );
  AND U23316 ( .A(n18772), .B(n18773), .Z(n18755) );
  NANDN U23317 ( .A(n18774), .B(n18775), .Z(n18773) );
  NANDN U23318 ( .A(n18776), .B(n18777), .Z(n18775) );
  IV U23319 ( .A(n18778), .Z(n18777) );
  NAND U23320 ( .A(n18778), .B(n18776), .Z(n18772) );
  AND U23321 ( .A(n18779), .B(n18780), .Z(n18753) );
  NAND U23322 ( .A(n18781), .B(n18782), .Z(n18780) );
  OR U23323 ( .A(n18783), .B(n18784), .Z(n18782) );
  NAND U23324 ( .A(n18784), .B(n18783), .Z(n18779) );
  IV U23325 ( .A(n18785), .Z(n18784) );
  NAND U23326 ( .A(n18786), .B(n18787), .Z(n18756) );
  NANDN U23327 ( .A(n18788), .B(n18789), .Z(n18787) );
  NAND U23328 ( .A(n18790), .B(n18791), .Z(n18789) );
  OR U23329 ( .A(n18791), .B(n18790), .Z(n18786) );
  IV U23330 ( .A(n18792), .Z(n18790) );
  AND U23331 ( .A(n18793), .B(n18794), .Z(n18759) );
  NAND U23332 ( .A(n18795), .B(n18796), .Z(n18794) );
  NANDN U23333 ( .A(n18797), .B(n18798), .Z(n18796) );
  NANDN U23334 ( .A(n18798), .B(n18797), .Z(n18793) );
  XOR U23335 ( .A(n18769), .B(n18799), .Z(n18761) );
  XNOR U23336 ( .A(n18766), .B(n18768), .Z(n18799) );
  AND U23337 ( .A(n18800), .B(n18801), .Z(n18768) );
  NANDN U23338 ( .A(n18802), .B(n18803), .Z(n18801) );
  NANDN U23339 ( .A(n18804), .B(n18805), .Z(n18803) );
  IV U23340 ( .A(n18806), .Z(n18805) );
  NAND U23341 ( .A(n18806), .B(n18804), .Z(n18800) );
  AND U23342 ( .A(n18807), .B(n18808), .Z(n18766) );
  NAND U23343 ( .A(n18809), .B(n18810), .Z(n18808) );
  OR U23344 ( .A(n18811), .B(n18812), .Z(n18810) );
  NAND U23345 ( .A(n18812), .B(n18811), .Z(n18807) );
  IV U23346 ( .A(n18813), .Z(n18812) );
  NAND U23347 ( .A(n18814), .B(n18815), .Z(n18769) );
  NANDN U23348 ( .A(n18816), .B(n18817), .Z(n18815) );
  NAND U23349 ( .A(n18818), .B(n18819), .Z(n18817) );
  OR U23350 ( .A(n18819), .B(n18818), .Z(n18814) );
  IV U23351 ( .A(n18820), .Z(n18818) );
  XOR U23352 ( .A(n18795), .B(n18821), .Z(N28602) );
  XNOR U23353 ( .A(n18798), .B(n18797), .Z(n18821) );
  XNOR U23354 ( .A(n18809), .B(n18822), .Z(n18797) );
  XOR U23355 ( .A(n18813), .B(n18811), .Z(n18822) );
  XOR U23356 ( .A(n18819), .B(n18823), .Z(n18811) );
  XOR U23357 ( .A(n18816), .B(n18820), .Z(n18823) );
  NAND U23358 ( .A(n18824), .B(n18825), .Z(n18820) );
  NAND U23359 ( .A(n18826), .B(n18827), .Z(n18825) );
  NAND U23360 ( .A(n18828), .B(n18829), .Z(n18824) );
  AND U23361 ( .A(n18830), .B(n18831), .Z(n18816) );
  NAND U23362 ( .A(n18832), .B(n18833), .Z(n18831) );
  NAND U23363 ( .A(n18834), .B(n18835), .Z(n18830) );
  NANDN U23364 ( .A(n18836), .B(n18837), .Z(n18819) );
  NANDN U23365 ( .A(n18838), .B(n18839), .Z(n18813) );
  XNOR U23366 ( .A(n18804), .B(n18840), .Z(n18809) );
  XOR U23367 ( .A(n18802), .B(n18806), .Z(n18840) );
  NAND U23368 ( .A(n18841), .B(n18842), .Z(n18806) );
  NAND U23369 ( .A(n18843), .B(n18844), .Z(n18842) );
  NAND U23370 ( .A(n18845), .B(n18846), .Z(n18841) );
  AND U23371 ( .A(n18847), .B(n18848), .Z(n18802) );
  NAND U23372 ( .A(n18849), .B(n18850), .Z(n18848) );
  NAND U23373 ( .A(n18851), .B(n18852), .Z(n18847) );
  AND U23374 ( .A(n18853), .B(n18854), .Z(n18804) );
  NAND U23375 ( .A(n18855), .B(n18856), .Z(n18798) );
  XNOR U23376 ( .A(n18781), .B(n18857), .Z(n18795) );
  XOR U23377 ( .A(n18785), .B(n18783), .Z(n18857) );
  XOR U23378 ( .A(n18791), .B(n18858), .Z(n18783) );
  XOR U23379 ( .A(n18788), .B(n18792), .Z(n18858) );
  NAND U23380 ( .A(n18859), .B(n18860), .Z(n18792) );
  NAND U23381 ( .A(n18861), .B(n18862), .Z(n18860) );
  NAND U23382 ( .A(n18863), .B(n18864), .Z(n18859) );
  AND U23383 ( .A(n18865), .B(n18866), .Z(n18788) );
  NAND U23384 ( .A(n18867), .B(n18868), .Z(n18866) );
  NAND U23385 ( .A(n18869), .B(n18870), .Z(n18865) );
  NANDN U23386 ( .A(n18871), .B(n18872), .Z(n18791) );
  NANDN U23387 ( .A(n18873), .B(n18874), .Z(n18785) );
  XNOR U23388 ( .A(n18776), .B(n18875), .Z(n18781) );
  XOR U23389 ( .A(n18774), .B(n18778), .Z(n18875) );
  NAND U23390 ( .A(n18876), .B(n18877), .Z(n18778) );
  NAND U23391 ( .A(n18878), .B(n18879), .Z(n18877) );
  NAND U23392 ( .A(n18880), .B(n18881), .Z(n18876) );
  AND U23393 ( .A(n18882), .B(n18883), .Z(n18774) );
  NAND U23394 ( .A(n18884), .B(n18885), .Z(n18883) );
  NAND U23395 ( .A(n18886), .B(n18887), .Z(n18882) );
  AND U23396 ( .A(n18888), .B(n18889), .Z(n18776) );
  XOR U23397 ( .A(n18856), .B(n18855), .Z(N28601) );
  XNOR U23398 ( .A(n18874), .B(n18873), .Z(n18855) );
  XNOR U23399 ( .A(n18888), .B(n18889), .Z(n18873) );
  XOR U23400 ( .A(n18885), .B(n18884), .Z(n18889) );
  XOR U23401 ( .A(y[1347]), .B(x[1347]), .Z(n18884) );
  XOR U23402 ( .A(n18887), .B(n18886), .Z(n18885) );
  XOR U23403 ( .A(y[1349]), .B(x[1349]), .Z(n18886) );
  XOR U23404 ( .A(y[1348]), .B(x[1348]), .Z(n18887) );
  XOR U23405 ( .A(n18879), .B(n18878), .Z(n18888) );
  XOR U23406 ( .A(n18881), .B(n18880), .Z(n18878) );
  XOR U23407 ( .A(y[1346]), .B(x[1346]), .Z(n18880) );
  XOR U23408 ( .A(y[1345]), .B(x[1345]), .Z(n18881) );
  XOR U23409 ( .A(y[1344]), .B(x[1344]), .Z(n18879) );
  XNOR U23410 ( .A(n18872), .B(n18871), .Z(n18874) );
  XNOR U23411 ( .A(n18868), .B(n18867), .Z(n18871) );
  XOR U23412 ( .A(n18870), .B(n18869), .Z(n18867) );
  XOR U23413 ( .A(y[1343]), .B(x[1343]), .Z(n18869) );
  XOR U23414 ( .A(y[1342]), .B(x[1342]), .Z(n18870) );
  XOR U23415 ( .A(y[1341]), .B(x[1341]), .Z(n18868) );
  XOR U23416 ( .A(n18862), .B(n18861), .Z(n18872) );
  XOR U23417 ( .A(n18864), .B(n18863), .Z(n18861) );
  XOR U23418 ( .A(y[1340]), .B(x[1340]), .Z(n18863) );
  XOR U23419 ( .A(y[1339]), .B(x[1339]), .Z(n18864) );
  XOR U23420 ( .A(y[1338]), .B(x[1338]), .Z(n18862) );
  XNOR U23421 ( .A(n18839), .B(n18838), .Z(n18856) );
  XNOR U23422 ( .A(n18853), .B(n18854), .Z(n18838) );
  XOR U23423 ( .A(n18850), .B(n18849), .Z(n18854) );
  XOR U23424 ( .A(y[1335]), .B(x[1335]), .Z(n18849) );
  XOR U23425 ( .A(n18852), .B(n18851), .Z(n18850) );
  XOR U23426 ( .A(y[1337]), .B(x[1337]), .Z(n18851) );
  XOR U23427 ( .A(y[1336]), .B(x[1336]), .Z(n18852) );
  XOR U23428 ( .A(n18844), .B(n18843), .Z(n18853) );
  XOR U23429 ( .A(n18846), .B(n18845), .Z(n18843) );
  XOR U23430 ( .A(y[1334]), .B(x[1334]), .Z(n18845) );
  XOR U23431 ( .A(y[1333]), .B(x[1333]), .Z(n18846) );
  XOR U23432 ( .A(y[1332]), .B(x[1332]), .Z(n18844) );
  XNOR U23433 ( .A(n18837), .B(n18836), .Z(n18839) );
  XNOR U23434 ( .A(n18833), .B(n18832), .Z(n18836) );
  XOR U23435 ( .A(n18835), .B(n18834), .Z(n18832) );
  XOR U23436 ( .A(y[1331]), .B(x[1331]), .Z(n18834) );
  XOR U23437 ( .A(y[1330]), .B(x[1330]), .Z(n18835) );
  XOR U23438 ( .A(y[1329]), .B(x[1329]), .Z(n18833) );
  XOR U23439 ( .A(n18827), .B(n18826), .Z(n18837) );
  XOR U23440 ( .A(n18829), .B(n18828), .Z(n18826) );
  XOR U23441 ( .A(y[1328]), .B(x[1328]), .Z(n18828) );
  XOR U23442 ( .A(y[1327]), .B(x[1327]), .Z(n18829) );
  XOR U23443 ( .A(y[1326]), .B(x[1326]), .Z(n18827) );
  NAND U23444 ( .A(n18890), .B(n18891), .Z(N28593) );
  NAND U23445 ( .A(n18892), .B(n18893), .Z(n18891) );
  NANDN U23446 ( .A(n18894), .B(n18895), .Z(n18893) );
  NANDN U23447 ( .A(n18895), .B(n18894), .Z(n18890) );
  XOR U23448 ( .A(n18894), .B(n18896), .Z(N28592) );
  XNOR U23449 ( .A(n18892), .B(n18895), .Z(n18896) );
  NAND U23450 ( .A(n18897), .B(n18898), .Z(n18895) );
  NAND U23451 ( .A(n18899), .B(n18900), .Z(n18898) );
  NANDN U23452 ( .A(n18901), .B(n18902), .Z(n18900) );
  NANDN U23453 ( .A(n18902), .B(n18901), .Z(n18897) );
  AND U23454 ( .A(n18903), .B(n18904), .Z(n18892) );
  NAND U23455 ( .A(n18905), .B(n18906), .Z(n18904) );
  OR U23456 ( .A(n18907), .B(n18908), .Z(n18906) );
  NAND U23457 ( .A(n18908), .B(n18907), .Z(n18903) );
  IV U23458 ( .A(n18909), .Z(n18908) );
  AND U23459 ( .A(n18910), .B(n18911), .Z(n18894) );
  NAND U23460 ( .A(n18912), .B(n18913), .Z(n18911) );
  NANDN U23461 ( .A(n18914), .B(n18915), .Z(n18913) );
  NANDN U23462 ( .A(n18915), .B(n18914), .Z(n18910) );
  XOR U23463 ( .A(n18907), .B(n18916), .Z(N28591) );
  XOR U23464 ( .A(n18905), .B(n18909), .Z(n18916) );
  XNOR U23465 ( .A(n18902), .B(n18917), .Z(n18909) );
  XNOR U23466 ( .A(n18899), .B(n18901), .Z(n18917) );
  AND U23467 ( .A(n18918), .B(n18919), .Z(n18901) );
  NANDN U23468 ( .A(n18920), .B(n18921), .Z(n18919) );
  NANDN U23469 ( .A(n18922), .B(n18923), .Z(n18921) );
  IV U23470 ( .A(n18924), .Z(n18923) );
  NAND U23471 ( .A(n18924), .B(n18922), .Z(n18918) );
  AND U23472 ( .A(n18925), .B(n18926), .Z(n18899) );
  NAND U23473 ( .A(n18927), .B(n18928), .Z(n18926) );
  OR U23474 ( .A(n18929), .B(n18930), .Z(n18928) );
  NAND U23475 ( .A(n18930), .B(n18929), .Z(n18925) );
  IV U23476 ( .A(n18931), .Z(n18930) );
  NAND U23477 ( .A(n18932), .B(n18933), .Z(n18902) );
  NANDN U23478 ( .A(n18934), .B(n18935), .Z(n18933) );
  NAND U23479 ( .A(n18936), .B(n18937), .Z(n18935) );
  OR U23480 ( .A(n18937), .B(n18936), .Z(n18932) );
  IV U23481 ( .A(n18938), .Z(n18936) );
  AND U23482 ( .A(n18939), .B(n18940), .Z(n18905) );
  NAND U23483 ( .A(n18941), .B(n18942), .Z(n18940) );
  NANDN U23484 ( .A(n18943), .B(n18944), .Z(n18942) );
  NANDN U23485 ( .A(n18944), .B(n18943), .Z(n18939) );
  XOR U23486 ( .A(n18915), .B(n18945), .Z(n18907) );
  XNOR U23487 ( .A(n18912), .B(n18914), .Z(n18945) );
  AND U23488 ( .A(n18946), .B(n18947), .Z(n18914) );
  NANDN U23489 ( .A(n18948), .B(n18949), .Z(n18947) );
  NANDN U23490 ( .A(n18950), .B(n18951), .Z(n18949) );
  IV U23491 ( .A(n18952), .Z(n18951) );
  NAND U23492 ( .A(n18952), .B(n18950), .Z(n18946) );
  AND U23493 ( .A(n18953), .B(n18954), .Z(n18912) );
  NAND U23494 ( .A(n18955), .B(n18956), .Z(n18954) );
  OR U23495 ( .A(n18957), .B(n18958), .Z(n18956) );
  NAND U23496 ( .A(n18958), .B(n18957), .Z(n18953) );
  IV U23497 ( .A(n18959), .Z(n18958) );
  NAND U23498 ( .A(n18960), .B(n18961), .Z(n18915) );
  NANDN U23499 ( .A(n18962), .B(n18963), .Z(n18961) );
  NAND U23500 ( .A(n18964), .B(n18965), .Z(n18963) );
  OR U23501 ( .A(n18965), .B(n18964), .Z(n18960) );
  IV U23502 ( .A(n18966), .Z(n18964) );
  XOR U23503 ( .A(n18941), .B(n18967), .Z(N28590) );
  XNOR U23504 ( .A(n18944), .B(n18943), .Z(n18967) );
  XNOR U23505 ( .A(n18955), .B(n18968), .Z(n18943) );
  XOR U23506 ( .A(n18959), .B(n18957), .Z(n18968) );
  XOR U23507 ( .A(n18965), .B(n18969), .Z(n18957) );
  XOR U23508 ( .A(n18962), .B(n18966), .Z(n18969) );
  NAND U23509 ( .A(n18970), .B(n18971), .Z(n18966) );
  NAND U23510 ( .A(n18972), .B(n18973), .Z(n18971) );
  NAND U23511 ( .A(n18974), .B(n18975), .Z(n18970) );
  AND U23512 ( .A(n18976), .B(n18977), .Z(n18962) );
  NAND U23513 ( .A(n18978), .B(n18979), .Z(n18977) );
  NAND U23514 ( .A(n18980), .B(n18981), .Z(n18976) );
  NANDN U23515 ( .A(n18982), .B(n18983), .Z(n18965) );
  NANDN U23516 ( .A(n18984), .B(n18985), .Z(n18959) );
  XNOR U23517 ( .A(n18950), .B(n18986), .Z(n18955) );
  XOR U23518 ( .A(n18948), .B(n18952), .Z(n18986) );
  NAND U23519 ( .A(n18987), .B(n18988), .Z(n18952) );
  NAND U23520 ( .A(n18989), .B(n18990), .Z(n18988) );
  NAND U23521 ( .A(n18991), .B(n18992), .Z(n18987) );
  AND U23522 ( .A(n18993), .B(n18994), .Z(n18948) );
  NAND U23523 ( .A(n18995), .B(n18996), .Z(n18994) );
  NAND U23524 ( .A(n18997), .B(n18998), .Z(n18993) );
  AND U23525 ( .A(n18999), .B(n19000), .Z(n18950) );
  NAND U23526 ( .A(n19001), .B(n19002), .Z(n18944) );
  XNOR U23527 ( .A(n18927), .B(n19003), .Z(n18941) );
  XOR U23528 ( .A(n18931), .B(n18929), .Z(n19003) );
  XOR U23529 ( .A(n18937), .B(n19004), .Z(n18929) );
  XOR U23530 ( .A(n18934), .B(n18938), .Z(n19004) );
  NAND U23531 ( .A(n19005), .B(n19006), .Z(n18938) );
  NAND U23532 ( .A(n19007), .B(n19008), .Z(n19006) );
  NAND U23533 ( .A(n19009), .B(n19010), .Z(n19005) );
  AND U23534 ( .A(n19011), .B(n19012), .Z(n18934) );
  NAND U23535 ( .A(n19013), .B(n19014), .Z(n19012) );
  NAND U23536 ( .A(n19015), .B(n19016), .Z(n19011) );
  NANDN U23537 ( .A(n19017), .B(n19018), .Z(n18937) );
  NANDN U23538 ( .A(n19019), .B(n19020), .Z(n18931) );
  XNOR U23539 ( .A(n18922), .B(n19021), .Z(n18927) );
  XOR U23540 ( .A(n18920), .B(n18924), .Z(n19021) );
  NAND U23541 ( .A(n19022), .B(n19023), .Z(n18924) );
  NAND U23542 ( .A(n19024), .B(n19025), .Z(n19023) );
  NAND U23543 ( .A(n19026), .B(n19027), .Z(n19022) );
  AND U23544 ( .A(n19028), .B(n19029), .Z(n18920) );
  NAND U23545 ( .A(n19030), .B(n19031), .Z(n19029) );
  NAND U23546 ( .A(n19032), .B(n19033), .Z(n19028) );
  AND U23547 ( .A(n19034), .B(n19035), .Z(n18922) );
  XOR U23548 ( .A(n19002), .B(n19001), .Z(N28589) );
  XNOR U23549 ( .A(n19020), .B(n19019), .Z(n19001) );
  XNOR U23550 ( .A(n19034), .B(n19035), .Z(n19019) );
  XOR U23551 ( .A(n19031), .B(n19030), .Z(n19035) );
  XOR U23552 ( .A(y[1323]), .B(x[1323]), .Z(n19030) );
  XOR U23553 ( .A(n19033), .B(n19032), .Z(n19031) );
  XOR U23554 ( .A(y[1325]), .B(x[1325]), .Z(n19032) );
  XOR U23555 ( .A(y[1324]), .B(x[1324]), .Z(n19033) );
  XOR U23556 ( .A(n19025), .B(n19024), .Z(n19034) );
  XOR U23557 ( .A(n19027), .B(n19026), .Z(n19024) );
  XOR U23558 ( .A(y[1322]), .B(x[1322]), .Z(n19026) );
  XOR U23559 ( .A(y[1321]), .B(x[1321]), .Z(n19027) );
  XOR U23560 ( .A(y[1320]), .B(x[1320]), .Z(n19025) );
  XNOR U23561 ( .A(n19018), .B(n19017), .Z(n19020) );
  XNOR U23562 ( .A(n19014), .B(n19013), .Z(n19017) );
  XOR U23563 ( .A(n19016), .B(n19015), .Z(n19013) );
  XOR U23564 ( .A(y[1319]), .B(x[1319]), .Z(n19015) );
  XOR U23565 ( .A(y[1318]), .B(x[1318]), .Z(n19016) );
  XOR U23566 ( .A(y[1317]), .B(x[1317]), .Z(n19014) );
  XOR U23567 ( .A(n19008), .B(n19007), .Z(n19018) );
  XOR U23568 ( .A(n19010), .B(n19009), .Z(n19007) );
  XOR U23569 ( .A(y[1316]), .B(x[1316]), .Z(n19009) );
  XOR U23570 ( .A(y[1315]), .B(x[1315]), .Z(n19010) );
  XOR U23571 ( .A(y[1314]), .B(x[1314]), .Z(n19008) );
  XNOR U23572 ( .A(n18985), .B(n18984), .Z(n19002) );
  XNOR U23573 ( .A(n18999), .B(n19000), .Z(n18984) );
  XOR U23574 ( .A(n18996), .B(n18995), .Z(n19000) );
  XOR U23575 ( .A(y[1311]), .B(x[1311]), .Z(n18995) );
  XOR U23576 ( .A(n18998), .B(n18997), .Z(n18996) );
  XOR U23577 ( .A(y[1313]), .B(x[1313]), .Z(n18997) );
  XOR U23578 ( .A(y[1312]), .B(x[1312]), .Z(n18998) );
  XOR U23579 ( .A(n18990), .B(n18989), .Z(n18999) );
  XOR U23580 ( .A(n18992), .B(n18991), .Z(n18989) );
  XOR U23581 ( .A(y[1310]), .B(x[1310]), .Z(n18991) );
  XOR U23582 ( .A(y[1309]), .B(x[1309]), .Z(n18992) );
  XOR U23583 ( .A(y[1308]), .B(x[1308]), .Z(n18990) );
  XNOR U23584 ( .A(n18983), .B(n18982), .Z(n18985) );
  XNOR U23585 ( .A(n18979), .B(n18978), .Z(n18982) );
  XOR U23586 ( .A(n18981), .B(n18980), .Z(n18978) );
  XOR U23587 ( .A(y[1307]), .B(x[1307]), .Z(n18980) );
  XOR U23588 ( .A(y[1306]), .B(x[1306]), .Z(n18981) );
  XOR U23589 ( .A(y[1305]), .B(x[1305]), .Z(n18979) );
  XOR U23590 ( .A(n18973), .B(n18972), .Z(n18983) );
  XOR U23591 ( .A(n18975), .B(n18974), .Z(n18972) );
  XOR U23592 ( .A(y[1304]), .B(x[1304]), .Z(n18974) );
  XOR U23593 ( .A(y[1303]), .B(x[1303]), .Z(n18975) );
  XOR U23594 ( .A(y[1302]), .B(x[1302]), .Z(n18973) );
  NAND U23595 ( .A(n19036), .B(n19037), .Z(N28581) );
  NAND U23596 ( .A(n19038), .B(n19039), .Z(n19037) );
  NANDN U23597 ( .A(n19040), .B(n19041), .Z(n19039) );
  NANDN U23598 ( .A(n19041), .B(n19040), .Z(n19036) );
  XOR U23599 ( .A(n19040), .B(n19042), .Z(N28580) );
  XNOR U23600 ( .A(n19038), .B(n19041), .Z(n19042) );
  NAND U23601 ( .A(n19043), .B(n19044), .Z(n19041) );
  NAND U23602 ( .A(n19045), .B(n19046), .Z(n19044) );
  NANDN U23603 ( .A(n19047), .B(n19048), .Z(n19046) );
  NANDN U23604 ( .A(n19048), .B(n19047), .Z(n19043) );
  AND U23605 ( .A(n19049), .B(n19050), .Z(n19038) );
  NAND U23606 ( .A(n19051), .B(n19052), .Z(n19050) );
  OR U23607 ( .A(n19053), .B(n19054), .Z(n19052) );
  NAND U23608 ( .A(n19054), .B(n19053), .Z(n19049) );
  IV U23609 ( .A(n19055), .Z(n19054) );
  AND U23610 ( .A(n19056), .B(n19057), .Z(n19040) );
  NAND U23611 ( .A(n19058), .B(n19059), .Z(n19057) );
  NANDN U23612 ( .A(n19060), .B(n19061), .Z(n19059) );
  NANDN U23613 ( .A(n19061), .B(n19060), .Z(n19056) );
  XOR U23614 ( .A(n19053), .B(n19062), .Z(N28579) );
  XOR U23615 ( .A(n19051), .B(n19055), .Z(n19062) );
  XNOR U23616 ( .A(n19048), .B(n19063), .Z(n19055) );
  XNOR U23617 ( .A(n19045), .B(n19047), .Z(n19063) );
  AND U23618 ( .A(n19064), .B(n19065), .Z(n19047) );
  NANDN U23619 ( .A(n19066), .B(n19067), .Z(n19065) );
  NANDN U23620 ( .A(n19068), .B(n19069), .Z(n19067) );
  IV U23621 ( .A(n19070), .Z(n19069) );
  NAND U23622 ( .A(n19070), .B(n19068), .Z(n19064) );
  AND U23623 ( .A(n19071), .B(n19072), .Z(n19045) );
  NAND U23624 ( .A(n19073), .B(n19074), .Z(n19072) );
  OR U23625 ( .A(n19075), .B(n19076), .Z(n19074) );
  NAND U23626 ( .A(n19076), .B(n19075), .Z(n19071) );
  IV U23627 ( .A(n19077), .Z(n19076) );
  NAND U23628 ( .A(n19078), .B(n19079), .Z(n19048) );
  NANDN U23629 ( .A(n19080), .B(n19081), .Z(n19079) );
  NAND U23630 ( .A(n19082), .B(n19083), .Z(n19081) );
  OR U23631 ( .A(n19083), .B(n19082), .Z(n19078) );
  IV U23632 ( .A(n19084), .Z(n19082) );
  AND U23633 ( .A(n19085), .B(n19086), .Z(n19051) );
  NAND U23634 ( .A(n19087), .B(n19088), .Z(n19086) );
  NANDN U23635 ( .A(n19089), .B(n19090), .Z(n19088) );
  NANDN U23636 ( .A(n19090), .B(n19089), .Z(n19085) );
  XOR U23637 ( .A(n19061), .B(n19091), .Z(n19053) );
  XNOR U23638 ( .A(n19058), .B(n19060), .Z(n19091) );
  AND U23639 ( .A(n19092), .B(n19093), .Z(n19060) );
  NANDN U23640 ( .A(n19094), .B(n19095), .Z(n19093) );
  NANDN U23641 ( .A(n19096), .B(n19097), .Z(n19095) );
  IV U23642 ( .A(n19098), .Z(n19097) );
  NAND U23643 ( .A(n19098), .B(n19096), .Z(n19092) );
  AND U23644 ( .A(n19099), .B(n19100), .Z(n19058) );
  NAND U23645 ( .A(n19101), .B(n19102), .Z(n19100) );
  OR U23646 ( .A(n19103), .B(n19104), .Z(n19102) );
  NAND U23647 ( .A(n19104), .B(n19103), .Z(n19099) );
  IV U23648 ( .A(n19105), .Z(n19104) );
  NAND U23649 ( .A(n19106), .B(n19107), .Z(n19061) );
  NANDN U23650 ( .A(n19108), .B(n19109), .Z(n19107) );
  NAND U23651 ( .A(n19110), .B(n19111), .Z(n19109) );
  OR U23652 ( .A(n19111), .B(n19110), .Z(n19106) );
  IV U23653 ( .A(n19112), .Z(n19110) );
  XOR U23654 ( .A(n19087), .B(n19113), .Z(N28578) );
  XNOR U23655 ( .A(n19090), .B(n19089), .Z(n19113) );
  XNOR U23656 ( .A(n19101), .B(n19114), .Z(n19089) );
  XOR U23657 ( .A(n19105), .B(n19103), .Z(n19114) );
  XOR U23658 ( .A(n19111), .B(n19115), .Z(n19103) );
  XOR U23659 ( .A(n19108), .B(n19112), .Z(n19115) );
  NAND U23660 ( .A(n19116), .B(n19117), .Z(n19112) );
  NAND U23661 ( .A(n19118), .B(n19119), .Z(n19117) );
  NAND U23662 ( .A(n19120), .B(n19121), .Z(n19116) );
  AND U23663 ( .A(n19122), .B(n19123), .Z(n19108) );
  NAND U23664 ( .A(n19124), .B(n19125), .Z(n19123) );
  NAND U23665 ( .A(n19126), .B(n19127), .Z(n19122) );
  NANDN U23666 ( .A(n19128), .B(n19129), .Z(n19111) );
  NANDN U23667 ( .A(n19130), .B(n19131), .Z(n19105) );
  XNOR U23668 ( .A(n19096), .B(n19132), .Z(n19101) );
  XOR U23669 ( .A(n19094), .B(n19098), .Z(n19132) );
  NAND U23670 ( .A(n19133), .B(n19134), .Z(n19098) );
  NAND U23671 ( .A(n19135), .B(n19136), .Z(n19134) );
  NAND U23672 ( .A(n19137), .B(n19138), .Z(n19133) );
  AND U23673 ( .A(n19139), .B(n19140), .Z(n19094) );
  NAND U23674 ( .A(n19141), .B(n19142), .Z(n19140) );
  NAND U23675 ( .A(n19143), .B(n19144), .Z(n19139) );
  AND U23676 ( .A(n19145), .B(n19146), .Z(n19096) );
  NAND U23677 ( .A(n19147), .B(n19148), .Z(n19090) );
  XNOR U23678 ( .A(n19073), .B(n19149), .Z(n19087) );
  XOR U23679 ( .A(n19077), .B(n19075), .Z(n19149) );
  XOR U23680 ( .A(n19083), .B(n19150), .Z(n19075) );
  XOR U23681 ( .A(n19080), .B(n19084), .Z(n19150) );
  NAND U23682 ( .A(n19151), .B(n19152), .Z(n19084) );
  NAND U23683 ( .A(n19153), .B(n19154), .Z(n19152) );
  NAND U23684 ( .A(n19155), .B(n19156), .Z(n19151) );
  AND U23685 ( .A(n19157), .B(n19158), .Z(n19080) );
  NAND U23686 ( .A(n19159), .B(n19160), .Z(n19158) );
  NAND U23687 ( .A(n19161), .B(n19162), .Z(n19157) );
  NANDN U23688 ( .A(n19163), .B(n19164), .Z(n19083) );
  NANDN U23689 ( .A(n19165), .B(n19166), .Z(n19077) );
  XNOR U23690 ( .A(n19068), .B(n19167), .Z(n19073) );
  XOR U23691 ( .A(n19066), .B(n19070), .Z(n19167) );
  NAND U23692 ( .A(n19168), .B(n19169), .Z(n19070) );
  NAND U23693 ( .A(n19170), .B(n19171), .Z(n19169) );
  NAND U23694 ( .A(n19172), .B(n19173), .Z(n19168) );
  AND U23695 ( .A(n19174), .B(n19175), .Z(n19066) );
  NAND U23696 ( .A(n19176), .B(n19177), .Z(n19175) );
  NAND U23697 ( .A(n19178), .B(n19179), .Z(n19174) );
  AND U23698 ( .A(n19180), .B(n19181), .Z(n19068) );
  XOR U23699 ( .A(n19148), .B(n19147), .Z(N28577) );
  XNOR U23700 ( .A(n19166), .B(n19165), .Z(n19147) );
  XNOR U23701 ( .A(n19180), .B(n19181), .Z(n19165) );
  XOR U23702 ( .A(n19177), .B(n19176), .Z(n19181) );
  XOR U23703 ( .A(y[1299]), .B(x[1299]), .Z(n19176) );
  XOR U23704 ( .A(n19179), .B(n19178), .Z(n19177) );
  XOR U23705 ( .A(y[1301]), .B(x[1301]), .Z(n19178) );
  XOR U23706 ( .A(y[1300]), .B(x[1300]), .Z(n19179) );
  XOR U23707 ( .A(n19171), .B(n19170), .Z(n19180) );
  XOR U23708 ( .A(n19173), .B(n19172), .Z(n19170) );
  XOR U23709 ( .A(y[1298]), .B(x[1298]), .Z(n19172) );
  XOR U23710 ( .A(y[1297]), .B(x[1297]), .Z(n19173) );
  XOR U23711 ( .A(y[1296]), .B(x[1296]), .Z(n19171) );
  XNOR U23712 ( .A(n19164), .B(n19163), .Z(n19166) );
  XNOR U23713 ( .A(n19160), .B(n19159), .Z(n19163) );
  XOR U23714 ( .A(n19162), .B(n19161), .Z(n19159) );
  XOR U23715 ( .A(y[1295]), .B(x[1295]), .Z(n19161) );
  XOR U23716 ( .A(y[1294]), .B(x[1294]), .Z(n19162) );
  XOR U23717 ( .A(y[1293]), .B(x[1293]), .Z(n19160) );
  XOR U23718 ( .A(n19154), .B(n19153), .Z(n19164) );
  XOR U23719 ( .A(n19156), .B(n19155), .Z(n19153) );
  XOR U23720 ( .A(y[1292]), .B(x[1292]), .Z(n19155) );
  XOR U23721 ( .A(y[1291]), .B(x[1291]), .Z(n19156) );
  XOR U23722 ( .A(y[1290]), .B(x[1290]), .Z(n19154) );
  XNOR U23723 ( .A(n19131), .B(n19130), .Z(n19148) );
  XNOR U23724 ( .A(n19145), .B(n19146), .Z(n19130) );
  XOR U23725 ( .A(n19142), .B(n19141), .Z(n19146) );
  XOR U23726 ( .A(y[1287]), .B(x[1287]), .Z(n19141) );
  XOR U23727 ( .A(n19144), .B(n19143), .Z(n19142) );
  XOR U23728 ( .A(y[1289]), .B(x[1289]), .Z(n19143) );
  XOR U23729 ( .A(y[1288]), .B(x[1288]), .Z(n19144) );
  XOR U23730 ( .A(n19136), .B(n19135), .Z(n19145) );
  XOR U23731 ( .A(n19138), .B(n19137), .Z(n19135) );
  XOR U23732 ( .A(y[1286]), .B(x[1286]), .Z(n19137) );
  XOR U23733 ( .A(y[1285]), .B(x[1285]), .Z(n19138) );
  XOR U23734 ( .A(y[1284]), .B(x[1284]), .Z(n19136) );
  XNOR U23735 ( .A(n19129), .B(n19128), .Z(n19131) );
  XNOR U23736 ( .A(n19125), .B(n19124), .Z(n19128) );
  XOR U23737 ( .A(n19127), .B(n19126), .Z(n19124) );
  XOR U23738 ( .A(y[1283]), .B(x[1283]), .Z(n19126) );
  XOR U23739 ( .A(y[1282]), .B(x[1282]), .Z(n19127) );
  XOR U23740 ( .A(y[1281]), .B(x[1281]), .Z(n19125) );
  XOR U23741 ( .A(n19119), .B(n19118), .Z(n19129) );
  XOR U23742 ( .A(n19121), .B(n19120), .Z(n19118) );
  XOR U23743 ( .A(y[1280]), .B(x[1280]), .Z(n19120) );
  XOR U23744 ( .A(y[1279]), .B(x[1279]), .Z(n19121) );
  XOR U23745 ( .A(y[1278]), .B(x[1278]), .Z(n19119) );
  NAND U23746 ( .A(n19182), .B(n19183), .Z(N28569) );
  NAND U23747 ( .A(n19184), .B(n19185), .Z(n19183) );
  NANDN U23748 ( .A(n19186), .B(n19187), .Z(n19185) );
  NANDN U23749 ( .A(n19187), .B(n19186), .Z(n19182) );
  XOR U23750 ( .A(n19186), .B(n19188), .Z(N28568) );
  XNOR U23751 ( .A(n19184), .B(n19187), .Z(n19188) );
  NAND U23752 ( .A(n19189), .B(n19190), .Z(n19187) );
  NAND U23753 ( .A(n19191), .B(n19192), .Z(n19190) );
  NANDN U23754 ( .A(n19193), .B(n19194), .Z(n19192) );
  NANDN U23755 ( .A(n19194), .B(n19193), .Z(n19189) );
  AND U23756 ( .A(n19195), .B(n19196), .Z(n19184) );
  NAND U23757 ( .A(n19197), .B(n19198), .Z(n19196) );
  OR U23758 ( .A(n19199), .B(n19200), .Z(n19198) );
  NAND U23759 ( .A(n19200), .B(n19199), .Z(n19195) );
  IV U23760 ( .A(n19201), .Z(n19200) );
  AND U23761 ( .A(n19202), .B(n19203), .Z(n19186) );
  NAND U23762 ( .A(n19204), .B(n19205), .Z(n19203) );
  NANDN U23763 ( .A(n19206), .B(n19207), .Z(n19205) );
  NANDN U23764 ( .A(n19207), .B(n19206), .Z(n19202) );
  XOR U23765 ( .A(n19199), .B(n19208), .Z(N28567) );
  XOR U23766 ( .A(n19197), .B(n19201), .Z(n19208) );
  XNOR U23767 ( .A(n19194), .B(n19209), .Z(n19201) );
  XNOR U23768 ( .A(n19191), .B(n19193), .Z(n19209) );
  AND U23769 ( .A(n19210), .B(n19211), .Z(n19193) );
  NANDN U23770 ( .A(n19212), .B(n19213), .Z(n19211) );
  NANDN U23771 ( .A(n19214), .B(n19215), .Z(n19213) );
  IV U23772 ( .A(n19216), .Z(n19215) );
  NAND U23773 ( .A(n19216), .B(n19214), .Z(n19210) );
  AND U23774 ( .A(n19217), .B(n19218), .Z(n19191) );
  NAND U23775 ( .A(n19219), .B(n19220), .Z(n19218) );
  OR U23776 ( .A(n19221), .B(n19222), .Z(n19220) );
  NAND U23777 ( .A(n19222), .B(n19221), .Z(n19217) );
  IV U23778 ( .A(n19223), .Z(n19222) );
  NAND U23779 ( .A(n19224), .B(n19225), .Z(n19194) );
  NANDN U23780 ( .A(n19226), .B(n19227), .Z(n19225) );
  NAND U23781 ( .A(n19228), .B(n19229), .Z(n19227) );
  OR U23782 ( .A(n19229), .B(n19228), .Z(n19224) );
  IV U23783 ( .A(n19230), .Z(n19228) );
  AND U23784 ( .A(n19231), .B(n19232), .Z(n19197) );
  NAND U23785 ( .A(n19233), .B(n19234), .Z(n19232) );
  NANDN U23786 ( .A(n19235), .B(n19236), .Z(n19234) );
  NANDN U23787 ( .A(n19236), .B(n19235), .Z(n19231) );
  XOR U23788 ( .A(n19207), .B(n19237), .Z(n19199) );
  XNOR U23789 ( .A(n19204), .B(n19206), .Z(n19237) );
  AND U23790 ( .A(n19238), .B(n19239), .Z(n19206) );
  NANDN U23791 ( .A(n19240), .B(n19241), .Z(n19239) );
  NANDN U23792 ( .A(n19242), .B(n19243), .Z(n19241) );
  IV U23793 ( .A(n19244), .Z(n19243) );
  NAND U23794 ( .A(n19244), .B(n19242), .Z(n19238) );
  AND U23795 ( .A(n19245), .B(n19246), .Z(n19204) );
  NAND U23796 ( .A(n19247), .B(n19248), .Z(n19246) );
  OR U23797 ( .A(n19249), .B(n19250), .Z(n19248) );
  NAND U23798 ( .A(n19250), .B(n19249), .Z(n19245) );
  IV U23799 ( .A(n19251), .Z(n19250) );
  NAND U23800 ( .A(n19252), .B(n19253), .Z(n19207) );
  NANDN U23801 ( .A(n19254), .B(n19255), .Z(n19253) );
  NAND U23802 ( .A(n19256), .B(n19257), .Z(n19255) );
  OR U23803 ( .A(n19257), .B(n19256), .Z(n19252) );
  IV U23804 ( .A(n19258), .Z(n19256) );
  XOR U23805 ( .A(n19233), .B(n19259), .Z(N28566) );
  XNOR U23806 ( .A(n19236), .B(n19235), .Z(n19259) );
  XNOR U23807 ( .A(n19247), .B(n19260), .Z(n19235) );
  XOR U23808 ( .A(n19251), .B(n19249), .Z(n19260) );
  XOR U23809 ( .A(n19257), .B(n19261), .Z(n19249) );
  XOR U23810 ( .A(n19254), .B(n19258), .Z(n19261) );
  NAND U23811 ( .A(n19262), .B(n19263), .Z(n19258) );
  NAND U23812 ( .A(n19264), .B(n19265), .Z(n19263) );
  NAND U23813 ( .A(n19266), .B(n19267), .Z(n19262) );
  AND U23814 ( .A(n19268), .B(n19269), .Z(n19254) );
  NAND U23815 ( .A(n19270), .B(n19271), .Z(n19269) );
  NAND U23816 ( .A(n19272), .B(n19273), .Z(n19268) );
  NANDN U23817 ( .A(n19274), .B(n19275), .Z(n19257) );
  NANDN U23818 ( .A(n19276), .B(n19277), .Z(n19251) );
  XNOR U23819 ( .A(n19242), .B(n19278), .Z(n19247) );
  XOR U23820 ( .A(n19240), .B(n19244), .Z(n19278) );
  NAND U23821 ( .A(n19279), .B(n19280), .Z(n19244) );
  NAND U23822 ( .A(n19281), .B(n19282), .Z(n19280) );
  NAND U23823 ( .A(n19283), .B(n19284), .Z(n19279) );
  AND U23824 ( .A(n19285), .B(n19286), .Z(n19240) );
  NAND U23825 ( .A(n19287), .B(n19288), .Z(n19286) );
  NAND U23826 ( .A(n19289), .B(n19290), .Z(n19285) );
  AND U23827 ( .A(n19291), .B(n19292), .Z(n19242) );
  NAND U23828 ( .A(n19293), .B(n19294), .Z(n19236) );
  XNOR U23829 ( .A(n19219), .B(n19295), .Z(n19233) );
  XOR U23830 ( .A(n19223), .B(n19221), .Z(n19295) );
  XOR U23831 ( .A(n19229), .B(n19296), .Z(n19221) );
  XOR U23832 ( .A(n19226), .B(n19230), .Z(n19296) );
  NAND U23833 ( .A(n19297), .B(n19298), .Z(n19230) );
  NAND U23834 ( .A(n19299), .B(n19300), .Z(n19298) );
  NAND U23835 ( .A(n19301), .B(n19302), .Z(n19297) );
  AND U23836 ( .A(n19303), .B(n19304), .Z(n19226) );
  NAND U23837 ( .A(n19305), .B(n19306), .Z(n19304) );
  NAND U23838 ( .A(n19307), .B(n19308), .Z(n19303) );
  NANDN U23839 ( .A(n19309), .B(n19310), .Z(n19229) );
  NANDN U23840 ( .A(n19311), .B(n19312), .Z(n19223) );
  XNOR U23841 ( .A(n19214), .B(n19313), .Z(n19219) );
  XOR U23842 ( .A(n19212), .B(n19216), .Z(n19313) );
  NAND U23843 ( .A(n19314), .B(n19315), .Z(n19216) );
  NAND U23844 ( .A(n19316), .B(n19317), .Z(n19315) );
  NAND U23845 ( .A(n19318), .B(n19319), .Z(n19314) );
  AND U23846 ( .A(n19320), .B(n19321), .Z(n19212) );
  NAND U23847 ( .A(n19322), .B(n19323), .Z(n19321) );
  NAND U23848 ( .A(n19324), .B(n19325), .Z(n19320) );
  AND U23849 ( .A(n19326), .B(n19327), .Z(n19214) );
  XOR U23850 ( .A(n19294), .B(n19293), .Z(N28565) );
  XNOR U23851 ( .A(n19312), .B(n19311), .Z(n19293) );
  XNOR U23852 ( .A(n19326), .B(n19327), .Z(n19311) );
  XOR U23853 ( .A(n19323), .B(n19322), .Z(n19327) );
  XOR U23854 ( .A(y[1275]), .B(x[1275]), .Z(n19322) );
  XOR U23855 ( .A(n19325), .B(n19324), .Z(n19323) );
  XOR U23856 ( .A(y[1277]), .B(x[1277]), .Z(n19324) );
  XOR U23857 ( .A(y[1276]), .B(x[1276]), .Z(n19325) );
  XOR U23858 ( .A(n19317), .B(n19316), .Z(n19326) );
  XOR U23859 ( .A(n19319), .B(n19318), .Z(n19316) );
  XOR U23860 ( .A(y[1274]), .B(x[1274]), .Z(n19318) );
  XOR U23861 ( .A(y[1273]), .B(x[1273]), .Z(n19319) );
  XOR U23862 ( .A(y[1272]), .B(x[1272]), .Z(n19317) );
  XNOR U23863 ( .A(n19310), .B(n19309), .Z(n19312) );
  XNOR U23864 ( .A(n19306), .B(n19305), .Z(n19309) );
  XOR U23865 ( .A(n19308), .B(n19307), .Z(n19305) );
  XOR U23866 ( .A(y[1271]), .B(x[1271]), .Z(n19307) );
  XOR U23867 ( .A(y[1270]), .B(x[1270]), .Z(n19308) );
  XOR U23868 ( .A(y[1269]), .B(x[1269]), .Z(n19306) );
  XOR U23869 ( .A(n19300), .B(n19299), .Z(n19310) );
  XOR U23870 ( .A(n19302), .B(n19301), .Z(n19299) );
  XOR U23871 ( .A(y[1268]), .B(x[1268]), .Z(n19301) );
  XOR U23872 ( .A(y[1267]), .B(x[1267]), .Z(n19302) );
  XOR U23873 ( .A(y[1266]), .B(x[1266]), .Z(n19300) );
  XNOR U23874 ( .A(n19277), .B(n19276), .Z(n19294) );
  XNOR U23875 ( .A(n19291), .B(n19292), .Z(n19276) );
  XOR U23876 ( .A(n19288), .B(n19287), .Z(n19292) );
  XOR U23877 ( .A(y[1263]), .B(x[1263]), .Z(n19287) );
  XOR U23878 ( .A(n19290), .B(n19289), .Z(n19288) );
  XOR U23879 ( .A(y[1265]), .B(x[1265]), .Z(n19289) );
  XOR U23880 ( .A(y[1264]), .B(x[1264]), .Z(n19290) );
  XOR U23881 ( .A(n19282), .B(n19281), .Z(n19291) );
  XOR U23882 ( .A(n19284), .B(n19283), .Z(n19281) );
  XOR U23883 ( .A(y[1262]), .B(x[1262]), .Z(n19283) );
  XOR U23884 ( .A(y[1261]), .B(x[1261]), .Z(n19284) );
  XOR U23885 ( .A(y[1260]), .B(x[1260]), .Z(n19282) );
  XNOR U23886 ( .A(n19275), .B(n19274), .Z(n19277) );
  XNOR U23887 ( .A(n19271), .B(n19270), .Z(n19274) );
  XOR U23888 ( .A(n19273), .B(n19272), .Z(n19270) );
  XOR U23889 ( .A(y[1259]), .B(x[1259]), .Z(n19272) );
  XOR U23890 ( .A(y[1258]), .B(x[1258]), .Z(n19273) );
  XOR U23891 ( .A(y[1257]), .B(x[1257]), .Z(n19271) );
  XOR U23892 ( .A(n19265), .B(n19264), .Z(n19275) );
  XOR U23893 ( .A(n19267), .B(n19266), .Z(n19264) );
  XOR U23894 ( .A(y[1256]), .B(x[1256]), .Z(n19266) );
  XOR U23895 ( .A(y[1255]), .B(x[1255]), .Z(n19267) );
  XOR U23896 ( .A(y[1254]), .B(x[1254]), .Z(n19265) );
  NAND U23897 ( .A(n19328), .B(n19329), .Z(N28557) );
  NAND U23898 ( .A(n19330), .B(n19331), .Z(n19329) );
  NANDN U23899 ( .A(n19332), .B(n19333), .Z(n19331) );
  NANDN U23900 ( .A(n19333), .B(n19332), .Z(n19328) );
  XOR U23901 ( .A(n19332), .B(n19334), .Z(N28556) );
  XNOR U23902 ( .A(n19330), .B(n19333), .Z(n19334) );
  NAND U23903 ( .A(n19335), .B(n19336), .Z(n19333) );
  NAND U23904 ( .A(n19337), .B(n19338), .Z(n19336) );
  NANDN U23905 ( .A(n19339), .B(n19340), .Z(n19338) );
  NANDN U23906 ( .A(n19340), .B(n19339), .Z(n19335) );
  AND U23907 ( .A(n19341), .B(n19342), .Z(n19330) );
  NAND U23908 ( .A(n19343), .B(n19344), .Z(n19342) );
  OR U23909 ( .A(n19345), .B(n19346), .Z(n19344) );
  NAND U23910 ( .A(n19346), .B(n19345), .Z(n19341) );
  IV U23911 ( .A(n19347), .Z(n19346) );
  AND U23912 ( .A(n19348), .B(n19349), .Z(n19332) );
  NAND U23913 ( .A(n19350), .B(n19351), .Z(n19349) );
  NANDN U23914 ( .A(n19352), .B(n19353), .Z(n19351) );
  NANDN U23915 ( .A(n19353), .B(n19352), .Z(n19348) );
  XOR U23916 ( .A(n19345), .B(n19354), .Z(N28555) );
  XOR U23917 ( .A(n19343), .B(n19347), .Z(n19354) );
  XNOR U23918 ( .A(n19340), .B(n19355), .Z(n19347) );
  XNOR U23919 ( .A(n19337), .B(n19339), .Z(n19355) );
  AND U23920 ( .A(n19356), .B(n19357), .Z(n19339) );
  NANDN U23921 ( .A(n19358), .B(n19359), .Z(n19357) );
  NANDN U23922 ( .A(n19360), .B(n19361), .Z(n19359) );
  IV U23923 ( .A(n19362), .Z(n19361) );
  NAND U23924 ( .A(n19362), .B(n19360), .Z(n19356) );
  AND U23925 ( .A(n19363), .B(n19364), .Z(n19337) );
  NAND U23926 ( .A(n19365), .B(n19366), .Z(n19364) );
  OR U23927 ( .A(n19367), .B(n19368), .Z(n19366) );
  NAND U23928 ( .A(n19368), .B(n19367), .Z(n19363) );
  IV U23929 ( .A(n19369), .Z(n19368) );
  NAND U23930 ( .A(n19370), .B(n19371), .Z(n19340) );
  NANDN U23931 ( .A(n19372), .B(n19373), .Z(n19371) );
  NAND U23932 ( .A(n19374), .B(n19375), .Z(n19373) );
  OR U23933 ( .A(n19375), .B(n19374), .Z(n19370) );
  IV U23934 ( .A(n19376), .Z(n19374) );
  AND U23935 ( .A(n19377), .B(n19378), .Z(n19343) );
  NAND U23936 ( .A(n19379), .B(n19380), .Z(n19378) );
  NANDN U23937 ( .A(n19381), .B(n19382), .Z(n19380) );
  NANDN U23938 ( .A(n19382), .B(n19381), .Z(n19377) );
  XOR U23939 ( .A(n19353), .B(n19383), .Z(n19345) );
  XNOR U23940 ( .A(n19350), .B(n19352), .Z(n19383) );
  AND U23941 ( .A(n19384), .B(n19385), .Z(n19352) );
  NANDN U23942 ( .A(n19386), .B(n19387), .Z(n19385) );
  NANDN U23943 ( .A(n19388), .B(n19389), .Z(n19387) );
  IV U23944 ( .A(n19390), .Z(n19389) );
  NAND U23945 ( .A(n19390), .B(n19388), .Z(n19384) );
  AND U23946 ( .A(n19391), .B(n19392), .Z(n19350) );
  NAND U23947 ( .A(n19393), .B(n19394), .Z(n19392) );
  OR U23948 ( .A(n19395), .B(n19396), .Z(n19394) );
  NAND U23949 ( .A(n19396), .B(n19395), .Z(n19391) );
  IV U23950 ( .A(n19397), .Z(n19396) );
  NAND U23951 ( .A(n19398), .B(n19399), .Z(n19353) );
  NANDN U23952 ( .A(n19400), .B(n19401), .Z(n19399) );
  NAND U23953 ( .A(n19402), .B(n19403), .Z(n19401) );
  OR U23954 ( .A(n19403), .B(n19402), .Z(n19398) );
  IV U23955 ( .A(n19404), .Z(n19402) );
  XOR U23956 ( .A(n19379), .B(n19405), .Z(N28554) );
  XNOR U23957 ( .A(n19382), .B(n19381), .Z(n19405) );
  XNOR U23958 ( .A(n19393), .B(n19406), .Z(n19381) );
  XOR U23959 ( .A(n19397), .B(n19395), .Z(n19406) );
  XOR U23960 ( .A(n19403), .B(n19407), .Z(n19395) );
  XOR U23961 ( .A(n19400), .B(n19404), .Z(n19407) );
  NAND U23962 ( .A(n19408), .B(n19409), .Z(n19404) );
  NAND U23963 ( .A(n19410), .B(n19411), .Z(n19409) );
  NAND U23964 ( .A(n19412), .B(n19413), .Z(n19408) );
  AND U23965 ( .A(n19414), .B(n19415), .Z(n19400) );
  NAND U23966 ( .A(n19416), .B(n19417), .Z(n19415) );
  NAND U23967 ( .A(n19418), .B(n19419), .Z(n19414) );
  NANDN U23968 ( .A(n19420), .B(n19421), .Z(n19403) );
  NANDN U23969 ( .A(n19422), .B(n19423), .Z(n19397) );
  XNOR U23970 ( .A(n19388), .B(n19424), .Z(n19393) );
  XOR U23971 ( .A(n19386), .B(n19390), .Z(n19424) );
  NAND U23972 ( .A(n19425), .B(n19426), .Z(n19390) );
  NAND U23973 ( .A(n19427), .B(n19428), .Z(n19426) );
  NAND U23974 ( .A(n19429), .B(n19430), .Z(n19425) );
  AND U23975 ( .A(n19431), .B(n19432), .Z(n19386) );
  NAND U23976 ( .A(n19433), .B(n19434), .Z(n19432) );
  NAND U23977 ( .A(n19435), .B(n19436), .Z(n19431) );
  AND U23978 ( .A(n19437), .B(n19438), .Z(n19388) );
  NAND U23979 ( .A(n19439), .B(n19440), .Z(n19382) );
  XNOR U23980 ( .A(n19365), .B(n19441), .Z(n19379) );
  XOR U23981 ( .A(n19369), .B(n19367), .Z(n19441) );
  XOR U23982 ( .A(n19375), .B(n19442), .Z(n19367) );
  XOR U23983 ( .A(n19372), .B(n19376), .Z(n19442) );
  NAND U23984 ( .A(n19443), .B(n19444), .Z(n19376) );
  NAND U23985 ( .A(n19445), .B(n19446), .Z(n19444) );
  NAND U23986 ( .A(n19447), .B(n19448), .Z(n19443) );
  AND U23987 ( .A(n19449), .B(n19450), .Z(n19372) );
  NAND U23988 ( .A(n19451), .B(n19452), .Z(n19450) );
  NAND U23989 ( .A(n19453), .B(n19454), .Z(n19449) );
  NANDN U23990 ( .A(n19455), .B(n19456), .Z(n19375) );
  NANDN U23991 ( .A(n19457), .B(n19458), .Z(n19369) );
  XNOR U23992 ( .A(n19360), .B(n19459), .Z(n19365) );
  XOR U23993 ( .A(n19358), .B(n19362), .Z(n19459) );
  NAND U23994 ( .A(n19460), .B(n19461), .Z(n19362) );
  NAND U23995 ( .A(n19462), .B(n19463), .Z(n19461) );
  NAND U23996 ( .A(n19464), .B(n19465), .Z(n19460) );
  AND U23997 ( .A(n19466), .B(n19467), .Z(n19358) );
  NAND U23998 ( .A(n19468), .B(n19469), .Z(n19467) );
  NAND U23999 ( .A(n19470), .B(n19471), .Z(n19466) );
  AND U24000 ( .A(n19472), .B(n19473), .Z(n19360) );
  XOR U24001 ( .A(n19440), .B(n19439), .Z(N28553) );
  XNOR U24002 ( .A(n19458), .B(n19457), .Z(n19439) );
  XNOR U24003 ( .A(n19472), .B(n19473), .Z(n19457) );
  XOR U24004 ( .A(n19469), .B(n19468), .Z(n19473) );
  XOR U24005 ( .A(y[1251]), .B(x[1251]), .Z(n19468) );
  XOR U24006 ( .A(n19471), .B(n19470), .Z(n19469) );
  XOR U24007 ( .A(y[1253]), .B(x[1253]), .Z(n19470) );
  XOR U24008 ( .A(y[1252]), .B(x[1252]), .Z(n19471) );
  XOR U24009 ( .A(n19463), .B(n19462), .Z(n19472) );
  XOR U24010 ( .A(n19465), .B(n19464), .Z(n19462) );
  XOR U24011 ( .A(y[1250]), .B(x[1250]), .Z(n19464) );
  XOR U24012 ( .A(y[1249]), .B(x[1249]), .Z(n19465) );
  XOR U24013 ( .A(y[1248]), .B(x[1248]), .Z(n19463) );
  XNOR U24014 ( .A(n19456), .B(n19455), .Z(n19458) );
  XNOR U24015 ( .A(n19452), .B(n19451), .Z(n19455) );
  XOR U24016 ( .A(n19454), .B(n19453), .Z(n19451) );
  XOR U24017 ( .A(y[1247]), .B(x[1247]), .Z(n19453) );
  XOR U24018 ( .A(y[1246]), .B(x[1246]), .Z(n19454) );
  XOR U24019 ( .A(y[1245]), .B(x[1245]), .Z(n19452) );
  XOR U24020 ( .A(n19446), .B(n19445), .Z(n19456) );
  XOR U24021 ( .A(n19448), .B(n19447), .Z(n19445) );
  XOR U24022 ( .A(y[1244]), .B(x[1244]), .Z(n19447) );
  XOR U24023 ( .A(y[1243]), .B(x[1243]), .Z(n19448) );
  XOR U24024 ( .A(y[1242]), .B(x[1242]), .Z(n19446) );
  XNOR U24025 ( .A(n19423), .B(n19422), .Z(n19440) );
  XNOR U24026 ( .A(n19437), .B(n19438), .Z(n19422) );
  XOR U24027 ( .A(n19434), .B(n19433), .Z(n19438) );
  XOR U24028 ( .A(y[1239]), .B(x[1239]), .Z(n19433) );
  XOR U24029 ( .A(n19436), .B(n19435), .Z(n19434) );
  XOR U24030 ( .A(y[1241]), .B(x[1241]), .Z(n19435) );
  XOR U24031 ( .A(y[1240]), .B(x[1240]), .Z(n19436) );
  XOR U24032 ( .A(n19428), .B(n19427), .Z(n19437) );
  XOR U24033 ( .A(n19430), .B(n19429), .Z(n19427) );
  XOR U24034 ( .A(y[1238]), .B(x[1238]), .Z(n19429) );
  XOR U24035 ( .A(y[1237]), .B(x[1237]), .Z(n19430) );
  XOR U24036 ( .A(y[1236]), .B(x[1236]), .Z(n19428) );
  XNOR U24037 ( .A(n19421), .B(n19420), .Z(n19423) );
  XNOR U24038 ( .A(n19417), .B(n19416), .Z(n19420) );
  XOR U24039 ( .A(n19419), .B(n19418), .Z(n19416) );
  XOR U24040 ( .A(y[1235]), .B(x[1235]), .Z(n19418) );
  XOR U24041 ( .A(y[1234]), .B(x[1234]), .Z(n19419) );
  XOR U24042 ( .A(y[1233]), .B(x[1233]), .Z(n19417) );
  XOR U24043 ( .A(n19411), .B(n19410), .Z(n19421) );
  XOR U24044 ( .A(n19413), .B(n19412), .Z(n19410) );
  XOR U24045 ( .A(y[1232]), .B(x[1232]), .Z(n19412) );
  XOR U24046 ( .A(y[1231]), .B(x[1231]), .Z(n19413) );
  XOR U24047 ( .A(y[1230]), .B(x[1230]), .Z(n19411) );
  NAND U24048 ( .A(n19474), .B(n19475), .Z(N28545) );
  NAND U24049 ( .A(n19476), .B(n19477), .Z(n19475) );
  NANDN U24050 ( .A(n19478), .B(n19479), .Z(n19477) );
  NANDN U24051 ( .A(n19479), .B(n19478), .Z(n19474) );
  XOR U24052 ( .A(n19478), .B(n19480), .Z(N28544) );
  XNOR U24053 ( .A(n19476), .B(n19479), .Z(n19480) );
  NAND U24054 ( .A(n19481), .B(n19482), .Z(n19479) );
  NAND U24055 ( .A(n19483), .B(n19484), .Z(n19482) );
  NANDN U24056 ( .A(n19485), .B(n19486), .Z(n19484) );
  NANDN U24057 ( .A(n19486), .B(n19485), .Z(n19481) );
  AND U24058 ( .A(n19487), .B(n19488), .Z(n19476) );
  NAND U24059 ( .A(n19489), .B(n19490), .Z(n19488) );
  OR U24060 ( .A(n19491), .B(n19492), .Z(n19490) );
  NAND U24061 ( .A(n19492), .B(n19491), .Z(n19487) );
  IV U24062 ( .A(n19493), .Z(n19492) );
  AND U24063 ( .A(n19494), .B(n19495), .Z(n19478) );
  NAND U24064 ( .A(n19496), .B(n19497), .Z(n19495) );
  NANDN U24065 ( .A(n19498), .B(n19499), .Z(n19497) );
  NANDN U24066 ( .A(n19499), .B(n19498), .Z(n19494) );
  XOR U24067 ( .A(n19491), .B(n19500), .Z(N28543) );
  XOR U24068 ( .A(n19489), .B(n19493), .Z(n19500) );
  XNOR U24069 ( .A(n19486), .B(n19501), .Z(n19493) );
  XNOR U24070 ( .A(n19483), .B(n19485), .Z(n19501) );
  AND U24071 ( .A(n19502), .B(n19503), .Z(n19485) );
  NANDN U24072 ( .A(n19504), .B(n19505), .Z(n19503) );
  NANDN U24073 ( .A(n19506), .B(n19507), .Z(n19505) );
  IV U24074 ( .A(n19508), .Z(n19507) );
  NAND U24075 ( .A(n19508), .B(n19506), .Z(n19502) );
  AND U24076 ( .A(n19509), .B(n19510), .Z(n19483) );
  NAND U24077 ( .A(n19511), .B(n19512), .Z(n19510) );
  OR U24078 ( .A(n19513), .B(n19514), .Z(n19512) );
  NAND U24079 ( .A(n19514), .B(n19513), .Z(n19509) );
  IV U24080 ( .A(n19515), .Z(n19514) );
  NAND U24081 ( .A(n19516), .B(n19517), .Z(n19486) );
  NANDN U24082 ( .A(n19518), .B(n19519), .Z(n19517) );
  NAND U24083 ( .A(n19520), .B(n19521), .Z(n19519) );
  OR U24084 ( .A(n19521), .B(n19520), .Z(n19516) );
  IV U24085 ( .A(n19522), .Z(n19520) );
  AND U24086 ( .A(n19523), .B(n19524), .Z(n19489) );
  NAND U24087 ( .A(n19525), .B(n19526), .Z(n19524) );
  NANDN U24088 ( .A(n19527), .B(n19528), .Z(n19526) );
  NANDN U24089 ( .A(n19528), .B(n19527), .Z(n19523) );
  XOR U24090 ( .A(n19499), .B(n19529), .Z(n19491) );
  XNOR U24091 ( .A(n19496), .B(n19498), .Z(n19529) );
  AND U24092 ( .A(n19530), .B(n19531), .Z(n19498) );
  NANDN U24093 ( .A(n19532), .B(n19533), .Z(n19531) );
  NANDN U24094 ( .A(n19534), .B(n19535), .Z(n19533) );
  IV U24095 ( .A(n19536), .Z(n19535) );
  NAND U24096 ( .A(n19536), .B(n19534), .Z(n19530) );
  AND U24097 ( .A(n19537), .B(n19538), .Z(n19496) );
  NAND U24098 ( .A(n19539), .B(n19540), .Z(n19538) );
  OR U24099 ( .A(n19541), .B(n19542), .Z(n19540) );
  NAND U24100 ( .A(n19542), .B(n19541), .Z(n19537) );
  IV U24101 ( .A(n19543), .Z(n19542) );
  NAND U24102 ( .A(n19544), .B(n19545), .Z(n19499) );
  NANDN U24103 ( .A(n19546), .B(n19547), .Z(n19545) );
  NAND U24104 ( .A(n19548), .B(n19549), .Z(n19547) );
  OR U24105 ( .A(n19549), .B(n19548), .Z(n19544) );
  IV U24106 ( .A(n19550), .Z(n19548) );
  XOR U24107 ( .A(n19525), .B(n19551), .Z(N28542) );
  XNOR U24108 ( .A(n19528), .B(n19527), .Z(n19551) );
  XNOR U24109 ( .A(n19539), .B(n19552), .Z(n19527) );
  XOR U24110 ( .A(n19543), .B(n19541), .Z(n19552) );
  XOR U24111 ( .A(n19549), .B(n19553), .Z(n19541) );
  XOR U24112 ( .A(n19546), .B(n19550), .Z(n19553) );
  NAND U24113 ( .A(n19554), .B(n19555), .Z(n19550) );
  NAND U24114 ( .A(n19556), .B(n19557), .Z(n19555) );
  NAND U24115 ( .A(n19558), .B(n19559), .Z(n19554) );
  AND U24116 ( .A(n19560), .B(n19561), .Z(n19546) );
  NAND U24117 ( .A(n19562), .B(n19563), .Z(n19561) );
  NAND U24118 ( .A(n19564), .B(n19565), .Z(n19560) );
  NANDN U24119 ( .A(n19566), .B(n19567), .Z(n19549) );
  NANDN U24120 ( .A(n19568), .B(n19569), .Z(n19543) );
  XNOR U24121 ( .A(n19534), .B(n19570), .Z(n19539) );
  XOR U24122 ( .A(n19532), .B(n19536), .Z(n19570) );
  NAND U24123 ( .A(n19571), .B(n19572), .Z(n19536) );
  NAND U24124 ( .A(n19573), .B(n19574), .Z(n19572) );
  NAND U24125 ( .A(n19575), .B(n19576), .Z(n19571) );
  AND U24126 ( .A(n19577), .B(n19578), .Z(n19532) );
  NAND U24127 ( .A(n19579), .B(n19580), .Z(n19578) );
  NAND U24128 ( .A(n19581), .B(n19582), .Z(n19577) );
  AND U24129 ( .A(n19583), .B(n19584), .Z(n19534) );
  NAND U24130 ( .A(n19585), .B(n19586), .Z(n19528) );
  XNOR U24131 ( .A(n19511), .B(n19587), .Z(n19525) );
  XOR U24132 ( .A(n19515), .B(n19513), .Z(n19587) );
  XOR U24133 ( .A(n19521), .B(n19588), .Z(n19513) );
  XOR U24134 ( .A(n19518), .B(n19522), .Z(n19588) );
  NAND U24135 ( .A(n19589), .B(n19590), .Z(n19522) );
  NAND U24136 ( .A(n19591), .B(n19592), .Z(n19590) );
  NAND U24137 ( .A(n19593), .B(n19594), .Z(n19589) );
  AND U24138 ( .A(n19595), .B(n19596), .Z(n19518) );
  NAND U24139 ( .A(n19597), .B(n19598), .Z(n19596) );
  NAND U24140 ( .A(n19599), .B(n19600), .Z(n19595) );
  NANDN U24141 ( .A(n19601), .B(n19602), .Z(n19521) );
  NANDN U24142 ( .A(n19603), .B(n19604), .Z(n19515) );
  XNOR U24143 ( .A(n19506), .B(n19605), .Z(n19511) );
  XOR U24144 ( .A(n19504), .B(n19508), .Z(n19605) );
  NAND U24145 ( .A(n19606), .B(n19607), .Z(n19508) );
  NAND U24146 ( .A(n19608), .B(n19609), .Z(n19607) );
  NAND U24147 ( .A(n19610), .B(n19611), .Z(n19606) );
  AND U24148 ( .A(n19612), .B(n19613), .Z(n19504) );
  NAND U24149 ( .A(n19614), .B(n19615), .Z(n19613) );
  NAND U24150 ( .A(n19616), .B(n19617), .Z(n19612) );
  AND U24151 ( .A(n19618), .B(n19619), .Z(n19506) );
  XOR U24152 ( .A(n19586), .B(n19585), .Z(N28541) );
  XNOR U24153 ( .A(n19604), .B(n19603), .Z(n19585) );
  XNOR U24154 ( .A(n19618), .B(n19619), .Z(n19603) );
  XOR U24155 ( .A(n19615), .B(n19614), .Z(n19619) );
  XOR U24156 ( .A(y[1227]), .B(x[1227]), .Z(n19614) );
  XOR U24157 ( .A(n19617), .B(n19616), .Z(n19615) );
  XOR U24158 ( .A(y[1229]), .B(x[1229]), .Z(n19616) );
  XOR U24159 ( .A(y[1228]), .B(x[1228]), .Z(n19617) );
  XOR U24160 ( .A(n19609), .B(n19608), .Z(n19618) );
  XOR U24161 ( .A(n19611), .B(n19610), .Z(n19608) );
  XOR U24162 ( .A(y[1226]), .B(x[1226]), .Z(n19610) );
  XOR U24163 ( .A(y[1225]), .B(x[1225]), .Z(n19611) );
  XOR U24164 ( .A(y[1224]), .B(x[1224]), .Z(n19609) );
  XNOR U24165 ( .A(n19602), .B(n19601), .Z(n19604) );
  XNOR U24166 ( .A(n19598), .B(n19597), .Z(n19601) );
  XOR U24167 ( .A(n19600), .B(n19599), .Z(n19597) );
  XOR U24168 ( .A(y[1223]), .B(x[1223]), .Z(n19599) );
  XOR U24169 ( .A(y[1222]), .B(x[1222]), .Z(n19600) );
  XOR U24170 ( .A(y[1221]), .B(x[1221]), .Z(n19598) );
  XOR U24171 ( .A(n19592), .B(n19591), .Z(n19602) );
  XOR U24172 ( .A(n19594), .B(n19593), .Z(n19591) );
  XOR U24173 ( .A(y[1220]), .B(x[1220]), .Z(n19593) );
  XOR U24174 ( .A(y[1219]), .B(x[1219]), .Z(n19594) );
  XOR U24175 ( .A(y[1218]), .B(x[1218]), .Z(n19592) );
  XNOR U24176 ( .A(n19569), .B(n19568), .Z(n19586) );
  XNOR U24177 ( .A(n19583), .B(n19584), .Z(n19568) );
  XOR U24178 ( .A(n19580), .B(n19579), .Z(n19584) );
  XOR U24179 ( .A(y[1215]), .B(x[1215]), .Z(n19579) );
  XOR U24180 ( .A(n19582), .B(n19581), .Z(n19580) );
  XOR U24181 ( .A(y[1217]), .B(x[1217]), .Z(n19581) );
  XOR U24182 ( .A(y[1216]), .B(x[1216]), .Z(n19582) );
  XOR U24183 ( .A(n19574), .B(n19573), .Z(n19583) );
  XOR U24184 ( .A(n19576), .B(n19575), .Z(n19573) );
  XOR U24185 ( .A(y[1214]), .B(x[1214]), .Z(n19575) );
  XOR U24186 ( .A(y[1213]), .B(x[1213]), .Z(n19576) );
  XOR U24187 ( .A(y[1212]), .B(x[1212]), .Z(n19574) );
  XNOR U24188 ( .A(n19567), .B(n19566), .Z(n19569) );
  XNOR U24189 ( .A(n19563), .B(n19562), .Z(n19566) );
  XOR U24190 ( .A(n19565), .B(n19564), .Z(n19562) );
  XOR U24191 ( .A(y[1211]), .B(x[1211]), .Z(n19564) );
  XOR U24192 ( .A(y[1210]), .B(x[1210]), .Z(n19565) );
  XOR U24193 ( .A(y[1209]), .B(x[1209]), .Z(n19563) );
  XOR U24194 ( .A(n19557), .B(n19556), .Z(n19567) );
  XOR U24195 ( .A(n19559), .B(n19558), .Z(n19556) );
  XOR U24196 ( .A(y[1208]), .B(x[1208]), .Z(n19558) );
  XOR U24197 ( .A(y[1207]), .B(x[1207]), .Z(n19559) );
  XOR U24198 ( .A(y[1206]), .B(x[1206]), .Z(n19557) );
  NAND U24199 ( .A(n19620), .B(n19621), .Z(N28533) );
  NAND U24200 ( .A(n19622), .B(n19623), .Z(n19621) );
  NANDN U24201 ( .A(n19624), .B(n19625), .Z(n19623) );
  NANDN U24202 ( .A(n19625), .B(n19624), .Z(n19620) );
  XOR U24203 ( .A(n19624), .B(n19626), .Z(N28532) );
  XNOR U24204 ( .A(n19622), .B(n19625), .Z(n19626) );
  NAND U24205 ( .A(n19627), .B(n19628), .Z(n19625) );
  NAND U24206 ( .A(n19629), .B(n19630), .Z(n19628) );
  NANDN U24207 ( .A(n19631), .B(n19632), .Z(n19630) );
  NANDN U24208 ( .A(n19632), .B(n19631), .Z(n19627) );
  AND U24209 ( .A(n19633), .B(n19634), .Z(n19622) );
  NAND U24210 ( .A(n19635), .B(n19636), .Z(n19634) );
  OR U24211 ( .A(n19637), .B(n19638), .Z(n19636) );
  NAND U24212 ( .A(n19638), .B(n19637), .Z(n19633) );
  IV U24213 ( .A(n19639), .Z(n19638) );
  AND U24214 ( .A(n19640), .B(n19641), .Z(n19624) );
  NAND U24215 ( .A(n19642), .B(n19643), .Z(n19641) );
  NANDN U24216 ( .A(n19644), .B(n19645), .Z(n19643) );
  NANDN U24217 ( .A(n19645), .B(n19644), .Z(n19640) );
  XOR U24218 ( .A(n19637), .B(n19646), .Z(N28531) );
  XOR U24219 ( .A(n19635), .B(n19639), .Z(n19646) );
  XNOR U24220 ( .A(n19632), .B(n19647), .Z(n19639) );
  XNOR U24221 ( .A(n19629), .B(n19631), .Z(n19647) );
  AND U24222 ( .A(n19648), .B(n19649), .Z(n19631) );
  NANDN U24223 ( .A(n19650), .B(n19651), .Z(n19649) );
  NANDN U24224 ( .A(n19652), .B(n19653), .Z(n19651) );
  IV U24225 ( .A(n19654), .Z(n19653) );
  NAND U24226 ( .A(n19654), .B(n19652), .Z(n19648) );
  AND U24227 ( .A(n19655), .B(n19656), .Z(n19629) );
  NAND U24228 ( .A(n19657), .B(n19658), .Z(n19656) );
  OR U24229 ( .A(n19659), .B(n19660), .Z(n19658) );
  NAND U24230 ( .A(n19660), .B(n19659), .Z(n19655) );
  IV U24231 ( .A(n19661), .Z(n19660) );
  NAND U24232 ( .A(n19662), .B(n19663), .Z(n19632) );
  NANDN U24233 ( .A(n19664), .B(n19665), .Z(n19663) );
  NAND U24234 ( .A(n19666), .B(n19667), .Z(n19665) );
  OR U24235 ( .A(n19667), .B(n19666), .Z(n19662) );
  IV U24236 ( .A(n19668), .Z(n19666) );
  AND U24237 ( .A(n19669), .B(n19670), .Z(n19635) );
  NAND U24238 ( .A(n19671), .B(n19672), .Z(n19670) );
  NANDN U24239 ( .A(n19673), .B(n19674), .Z(n19672) );
  NANDN U24240 ( .A(n19674), .B(n19673), .Z(n19669) );
  XOR U24241 ( .A(n19645), .B(n19675), .Z(n19637) );
  XNOR U24242 ( .A(n19642), .B(n19644), .Z(n19675) );
  AND U24243 ( .A(n19676), .B(n19677), .Z(n19644) );
  NANDN U24244 ( .A(n19678), .B(n19679), .Z(n19677) );
  NANDN U24245 ( .A(n19680), .B(n19681), .Z(n19679) );
  IV U24246 ( .A(n19682), .Z(n19681) );
  NAND U24247 ( .A(n19682), .B(n19680), .Z(n19676) );
  AND U24248 ( .A(n19683), .B(n19684), .Z(n19642) );
  NAND U24249 ( .A(n19685), .B(n19686), .Z(n19684) );
  OR U24250 ( .A(n19687), .B(n19688), .Z(n19686) );
  NAND U24251 ( .A(n19688), .B(n19687), .Z(n19683) );
  IV U24252 ( .A(n19689), .Z(n19688) );
  NAND U24253 ( .A(n19690), .B(n19691), .Z(n19645) );
  NANDN U24254 ( .A(n19692), .B(n19693), .Z(n19691) );
  NAND U24255 ( .A(n19694), .B(n19695), .Z(n19693) );
  OR U24256 ( .A(n19695), .B(n19694), .Z(n19690) );
  IV U24257 ( .A(n19696), .Z(n19694) );
  XOR U24258 ( .A(n19671), .B(n19697), .Z(N28530) );
  XNOR U24259 ( .A(n19674), .B(n19673), .Z(n19697) );
  XNOR U24260 ( .A(n19685), .B(n19698), .Z(n19673) );
  XOR U24261 ( .A(n19689), .B(n19687), .Z(n19698) );
  XOR U24262 ( .A(n19695), .B(n19699), .Z(n19687) );
  XOR U24263 ( .A(n19692), .B(n19696), .Z(n19699) );
  NAND U24264 ( .A(n19700), .B(n19701), .Z(n19696) );
  NAND U24265 ( .A(n19702), .B(n19703), .Z(n19701) );
  NAND U24266 ( .A(n19704), .B(n19705), .Z(n19700) );
  AND U24267 ( .A(n19706), .B(n19707), .Z(n19692) );
  NAND U24268 ( .A(n19708), .B(n19709), .Z(n19707) );
  NAND U24269 ( .A(n19710), .B(n19711), .Z(n19706) );
  NANDN U24270 ( .A(n19712), .B(n19713), .Z(n19695) );
  NANDN U24271 ( .A(n19714), .B(n19715), .Z(n19689) );
  XNOR U24272 ( .A(n19680), .B(n19716), .Z(n19685) );
  XOR U24273 ( .A(n19678), .B(n19682), .Z(n19716) );
  NAND U24274 ( .A(n19717), .B(n19718), .Z(n19682) );
  NAND U24275 ( .A(n19719), .B(n19720), .Z(n19718) );
  NAND U24276 ( .A(n19721), .B(n19722), .Z(n19717) );
  AND U24277 ( .A(n19723), .B(n19724), .Z(n19678) );
  NAND U24278 ( .A(n19725), .B(n19726), .Z(n19724) );
  NAND U24279 ( .A(n19727), .B(n19728), .Z(n19723) );
  AND U24280 ( .A(n19729), .B(n19730), .Z(n19680) );
  NAND U24281 ( .A(n19731), .B(n19732), .Z(n19674) );
  XNOR U24282 ( .A(n19657), .B(n19733), .Z(n19671) );
  XOR U24283 ( .A(n19661), .B(n19659), .Z(n19733) );
  XOR U24284 ( .A(n19667), .B(n19734), .Z(n19659) );
  XOR U24285 ( .A(n19664), .B(n19668), .Z(n19734) );
  NAND U24286 ( .A(n19735), .B(n19736), .Z(n19668) );
  NAND U24287 ( .A(n19737), .B(n19738), .Z(n19736) );
  NAND U24288 ( .A(n19739), .B(n19740), .Z(n19735) );
  AND U24289 ( .A(n19741), .B(n19742), .Z(n19664) );
  NAND U24290 ( .A(n19743), .B(n19744), .Z(n19742) );
  NAND U24291 ( .A(n19745), .B(n19746), .Z(n19741) );
  NANDN U24292 ( .A(n19747), .B(n19748), .Z(n19667) );
  NANDN U24293 ( .A(n19749), .B(n19750), .Z(n19661) );
  XNOR U24294 ( .A(n19652), .B(n19751), .Z(n19657) );
  XOR U24295 ( .A(n19650), .B(n19654), .Z(n19751) );
  NAND U24296 ( .A(n19752), .B(n19753), .Z(n19654) );
  NAND U24297 ( .A(n19754), .B(n19755), .Z(n19753) );
  NAND U24298 ( .A(n19756), .B(n19757), .Z(n19752) );
  AND U24299 ( .A(n19758), .B(n19759), .Z(n19650) );
  NAND U24300 ( .A(n19760), .B(n19761), .Z(n19759) );
  NAND U24301 ( .A(n19762), .B(n19763), .Z(n19758) );
  AND U24302 ( .A(n19764), .B(n19765), .Z(n19652) );
  XOR U24303 ( .A(n19732), .B(n19731), .Z(N28529) );
  XNOR U24304 ( .A(n19750), .B(n19749), .Z(n19731) );
  XNOR U24305 ( .A(n19764), .B(n19765), .Z(n19749) );
  XOR U24306 ( .A(n19761), .B(n19760), .Z(n19765) );
  XOR U24307 ( .A(y[1203]), .B(x[1203]), .Z(n19760) );
  XOR U24308 ( .A(n19763), .B(n19762), .Z(n19761) );
  XOR U24309 ( .A(y[1205]), .B(x[1205]), .Z(n19762) );
  XOR U24310 ( .A(y[1204]), .B(x[1204]), .Z(n19763) );
  XOR U24311 ( .A(n19755), .B(n19754), .Z(n19764) );
  XOR U24312 ( .A(n19757), .B(n19756), .Z(n19754) );
  XOR U24313 ( .A(y[1202]), .B(x[1202]), .Z(n19756) );
  XOR U24314 ( .A(y[1201]), .B(x[1201]), .Z(n19757) );
  XOR U24315 ( .A(y[1200]), .B(x[1200]), .Z(n19755) );
  XNOR U24316 ( .A(n19748), .B(n19747), .Z(n19750) );
  XNOR U24317 ( .A(n19744), .B(n19743), .Z(n19747) );
  XOR U24318 ( .A(n19746), .B(n19745), .Z(n19743) );
  XOR U24319 ( .A(y[1199]), .B(x[1199]), .Z(n19745) );
  XOR U24320 ( .A(y[1198]), .B(x[1198]), .Z(n19746) );
  XOR U24321 ( .A(y[1197]), .B(x[1197]), .Z(n19744) );
  XOR U24322 ( .A(n19738), .B(n19737), .Z(n19748) );
  XOR U24323 ( .A(n19740), .B(n19739), .Z(n19737) );
  XOR U24324 ( .A(y[1196]), .B(x[1196]), .Z(n19739) );
  XOR U24325 ( .A(y[1195]), .B(x[1195]), .Z(n19740) );
  XOR U24326 ( .A(y[1194]), .B(x[1194]), .Z(n19738) );
  XNOR U24327 ( .A(n19715), .B(n19714), .Z(n19732) );
  XNOR U24328 ( .A(n19729), .B(n19730), .Z(n19714) );
  XOR U24329 ( .A(n19726), .B(n19725), .Z(n19730) );
  XOR U24330 ( .A(y[1191]), .B(x[1191]), .Z(n19725) );
  XOR U24331 ( .A(n19728), .B(n19727), .Z(n19726) );
  XOR U24332 ( .A(y[1193]), .B(x[1193]), .Z(n19727) );
  XOR U24333 ( .A(y[1192]), .B(x[1192]), .Z(n19728) );
  XOR U24334 ( .A(n19720), .B(n19719), .Z(n19729) );
  XOR U24335 ( .A(n19722), .B(n19721), .Z(n19719) );
  XOR U24336 ( .A(y[1190]), .B(x[1190]), .Z(n19721) );
  XOR U24337 ( .A(y[1189]), .B(x[1189]), .Z(n19722) );
  XOR U24338 ( .A(y[1188]), .B(x[1188]), .Z(n19720) );
  XNOR U24339 ( .A(n19713), .B(n19712), .Z(n19715) );
  XNOR U24340 ( .A(n19709), .B(n19708), .Z(n19712) );
  XOR U24341 ( .A(n19711), .B(n19710), .Z(n19708) );
  XOR U24342 ( .A(y[1187]), .B(x[1187]), .Z(n19710) );
  XOR U24343 ( .A(y[1186]), .B(x[1186]), .Z(n19711) );
  XOR U24344 ( .A(y[1185]), .B(x[1185]), .Z(n19709) );
  XOR U24345 ( .A(n19703), .B(n19702), .Z(n19713) );
  XOR U24346 ( .A(n19705), .B(n19704), .Z(n19702) );
  XOR U24347 ( .A(y[1184]), .B(x[1184]), .Z(n19704) );
  XOR U24348 ( .A(y[1183]), .B(x[1183]), .Z(n19705) );
  XOR U24349 ( .A(y[1182]), .B(x[1182]), .Z(n19703) );
  NAND U24350 ( .A(n19766), .B(n19767), .Z(N28521) );
  NAND U24351 ( .A(n19768), .B(n19769), .Z(n19767) );
  NANDN U24352 ( .A(n19770), .B(n19771), .Z(n19769) );
  NANDN U24353 ( .A(n19771), .B(n19770), .Z(n19766) );
  XOR U24354 ( .A(n19770), .B(n19772), .Z(N28520) );
  XNOR U24355 ( .A(n19768), .B(n19771), .Z(n19772) );
  NAND U24356 ( .A(n19773), .B(n19774), .Z(n19771) );
  NAND U24357 ( .A(n19775), .B(n19776), .Z(n19774) );
  NANDN U24358 ( .A(n19777), .B(n19778), .Z(n19776) );
  NANDN U24359 ( .A(n19778), .B(n19777), .Z(n19773) );
  AND U24360 ( .A(n19779), .B(n19780), .Z(n19768) );
  NAND U24361 ( .A(n19781), .B(n19782), .Z(n19780) );
  OR U24362 ( .A(n19783), .B(n19784), .Z(n19782) );
  NAND U24363 ( .A(n19784), .B(n19783), .Z(n19779) );
  IV U24364 ( .A(n19785), .Z(n19784) );
  AND U24365 ( .A(n19786), .B(n19787), .Z(n19770) );
  NAND U24366 ( .A(n19788), .B(n19789), .Z(n19787) );
  NANDN U24367 ( .A(n19790), .B(n19791), .Z(n19789) );
  NANDN U24368 ( .A(n19791), .B(n19790), .Z(n19786) );
  XOR U24369 ( .A(n19783), .B(n19792), .Z(N28519) );
  XOR U24370 ( .A(n19781), .B(n19785), .Z(n19792) );
  XNOR U24371 ( .A(n19778), .B(n19793), .Z(n19785) );
  XNOR U24372 ( .A(n19775), .B(n19777), .Z(n19793) );
  AND U24373 ( .A(n19794), .B(n19795), .Z(n19777) );
  NANDN U24374 ( .A(n19796), .B(n19797), .Z(n19795) );
  NANDN U24375 ( .A(n19798), .B(n19799), .Z(n19797) );
  IV U24376 ( .A(n19800), .Z(n19799) );
  NAND U24377 ( .A(n19800), .B(n19798), .Z(n19794) );
  AND U24378 ( .A(n19801), .B(n19802), .Z(n19775) );
  NAND U24379 ( .A(n19803), .B(n19804), .Z(n19802) );
  OR U24380 ( .A(n19805), .B(n19806), .Z(n19804) );
  NAND U24381 ( .A(n19806), .B(n19805), .Z(n19801) );
  IV U24382 ( .A(n19807), .Z(n19806) );
  NAND U24383 ( .A(n19808), .B(n19809), .Z(n19778) );
  NANDN U24384 ( .A(n19810), .B(n19811), .Z(n19809) );
  NAND U24385 ( .A(n19812), .B(n19813), .Z(n19811) );
  OR U24386 ( .A(n19813), .B(n19812), .Z(n19808) );
  IV U24387 ( .A(n19814), .Z(n19812) );
  AND U24388 ( .A(n19815), .B(n19816), .Z(n19781) );
  NAND U24389 ( .A(n19817), .B(n19818), .Z(n19816) );
  NANDN U24390 ( .A(n19819), .B(n19820), .Z(n19818) );
  NANDN U24391 ( .A(n19820), .B(n19819), .Z(n19815) );
  XOR U24392 ( .A(n19791), .B(n19821), .Z(n19783) );
  XNOR U24393 ( .A(n19788), .B(n19790), .Z(n19821) );
  AND U24394 ( .A(n19822), .B(n19823), .Z(n19790) );
  NANDN U24395 ( .A(n19824), .B(n19825), .Z(n19823) );
  NANDN U24396 ( .A(n19826), .B(n19827), .Z(n19825) );
  IV U24397 ( .A(n19828), .Z(n19827) );
  NAND U24398 ( .A(n19828), .B(n19826), .Z(n19822) );
  AND U24399 ( .A(n19829), .B(n19830), .Z(n19788) );
  NAND U24400 ( .A(n19831), .B(n19832), .Z(n19830) );
  OR U24401 ( .A(n19833), .B(n19834), .Z(n19832) );
  NAND U24402 ( .A(n19834), .B(n19833), .Z(n19829) );
  IV U24403 ( .A(n19835), .Z(n19834) );
  NAND U24404 ( .A(n19836), .B(n19837), .Z(n19791) );
  NANDN U24405 ( .A(n19838), .B(n19839), .Z(n19837) );
  NAND U24406 ( .A(n19840), .B(n19841), .Z(n19839) );
  OR U24407 ( .A(n19841), .B(n19840), .Z(n19836) );
  IV U24408 ( .A(n19842), .Z(n19840) );
  XOR U24409 ( .A(n19817), .B(n19843), .Z(N28518) );
  XNOR U24410 ( .A(n19820), .B(n19819), .Z(n19843) );
  XNOR U24411 ( .A(n19831), .B(n19844), .Z(n19819) );
  XOR U24412 ( .A(n19835), .B(n19833), .Z(n19844) );
  XOR U24413 ( .A(n19841), .B(n19845), .Z(n19833) );
  XOR U24414 ( .A(n19838), .B(n19842), .Z(n19845) );
  NAND U24415 ( .A(n19846), .B(n19847), .Z(n19842) );
  NAND U24416 ( .A(n19848), .B(n19849), .Z(n19847) );
  NAND U24417 ( .A(n19850), .B(n19851), .Z(n19846) );
  AND U24418 ( .A(n19852), .B(n19853), .Z(n19838) );
  NAND U24419 ( .A(n19854), .B(n19855), .Z(n19853) );
  NAND U24420 ( .A(n19856), .B(n19857), .Z(n19852) );
  NANDN U24421 ( .A(n19858), .B(n19859), .Z(n19841) );
  NANDN U24422 ( .A(n19860), .B(n19861), .Z(n19835) );
  XNOR U24423 ( .A(n19826), .B(n19862), .Z(n19831) );
  XOR U24424 ( .A(n19824), .B(n19828), .Z(n19862) );
  NAND U24425 ( .A(n19863), .B(n19864), .Z(n19828) );
  NAND U24426 ( .A(n19865), .B(n19866), .Z(n19864) );
  NAND U24427 ( .A(n19867), .B(n19868), .Z(n19863) );
  AND U24428 ( .A(n19869), .B(n19870), .Z(n19824) );
  NAND U24429 ( .A(n19871), .B(n19872), .Z(n19870) );
  NAND U24430 ( .A(n19873), .B(n19874), .Z(n19869) );
  AND U24431 ( .A(n19875), .B(n19876), .Z(n19826) );
  NAND U24432 ( .A(n19877), .B(n19878), .Z(n19820) );
  XNOR U24433 ( .A(n19803), .B(n19879), .Z(n19817) );
  XOR U24434 ( .A(n19807), .B(n19805), .Z(n19879) );
  XOR U24435 ( .A(n19813), .B(n19880), .Z(n19805) );
  XOR U24436 ( .A(n19810), .B(n19814), .Z(n19880) );
  NAND U24437 ( .A(n19881), .B(n19882), .Z(n19814) );
  NAND U24438 ( .A(n19883), .B(n19884), .Z(n19882) );
  NAND U24439 ( .A(n19885), .B(n19886), .Z(n19881) );
  AND U24440 ( .A(n19887), .B(n19888), .Z(n19810) );
  NAND U24441 ( .A(n19889), .B(n19890), .Z(n19888) );
  NAND U24442 ( .A(n19891), .B(n19892), .Z(n19887) );
  NANDN U24443 ( .A(n19893), .B(n19894), .Z(n19813) );
  NANDN U24444 ( .A(n19895), .B(n19896), .Z(n19807) );
  XNOR U24445 ( .A(n19798), .B(n19897), .Z(n19803) );
  XOR U24446 ( .A(n19796), .B(n19800), .Z(n19897) );
  NAND U24447 ( .A(n19898), .B(n19899), .Z(n19800) );
  NAND U24448 ( .A(n19900), .B(n19901), .Z(n19899) );
  NAND U24449 ( .A(n19902), .B(n19903), .Z(n19898) );
  AND U24450 ( .A(n19904), .B(n19905), .Z(n19796) );
  NAND U24451 ( .A(n19906), .B(n19907), .Z(n19905) );
  NAND U24452 ( .A(n19908), .B(n19909), .Z(n19904) );
  AND U24453 ( .A(n19910), .B(n19911), .Z(n19798) );
  XOR U24454 ( .A(n19878), .B(n19877), .Z(N28517) );
  XNOR U24455 ( .A(n19896), .B(n19895), .Z(n19877) );
  XNOR U24456 ( .A(n19910), .B(n19911), .Z(n19895) );
  XOR U24457 ( .A(n19907), .B(n19906), .Z(n19911) );
  XOR U24458 ( .A(y[1179]), .B(x[1179]), .Z(n19906) );
  XOR U24459 ( .A(n19909), .B(n19908), .Z(n19907) );
  XOR U24460 ( .A(y[1181]), .B(x[1181]), .Z(n19908) );
  XOR U24461 ( .A(y[1180]), .B(x[1180]), .Z(n19909) );
  XOR U24462 ( .A(n19901), .B(n19900), .Z(n19910) );
  XOR U24463 ( .A(n19903), .B(n19902), .Z(n19900) );
  XOR U24464 ( .A(y[1178]), .B(x[1178]), .Z(n19902) );
  XOR U24465 ( .A(y[1177]), .B(x[1177]), .Z(n19903) );
  XOR U24466 ( .A(y[1176]), .B(x[1176]), .Z(n19901) );
  XNOR U24467 ( .A(n19894), .B(n19893), .Z(n19896) );
  XNOR U24468 ( .A(n19890), .B(n19889), .Z(n19893) );
  XOR U24469 ( .A(n19892), .B(n19891), .Z(n19889) );
  XOR U24470 ( .A(y[1175]), .B(x[1175]), .Z(n19891) );
  XOR U24471 ( .A(y[1174]), .B(x[1174]), .Z(n19892) );
  XOR U24472 ( .A(y[1173]), .B(x[1173]), .Z(n19890) );
  XOR U24473 ( .A(n19884), .B(n19883), .Z(n19894) );
  XOR U24474 ( .A(n19886), .B(n19885), .Z(n19883) );
  XOR U24475 ( .A(y[1172]), .B(x[1172]), .Z(n19885) );
  XOR U24476 ( .A(y[1171]), .B(x[1171]), .Z(n19886) );
  XOR U24477 ( .A(y[1170]), .B(x[1170]), .Z(n19884) );
  XNOR U24478 ( .A(n19861), .B(n19860), .Z(n19878) );
  XNOR U24479 ( .A(n19875), .B(n19876), .Z(n19860) );
  XOR U24480 ( .A(n19872), .B(n19871), .Z(n19876) );
  XOR U24481 ( .A(y[1167]), .B(x[1167]), .Z(n19871) );
  XOR U24482 ( .A(n19874), .B(n19873), .Z(n19872) );
  XOR U24483 ( .A(y[1169]), .B(x[1169]), .Z(n19873) );
  XOR U24484 ( .A(y[1168]), .B(x[1168]), .Z(n19874) );
  XOR U24485 ( .A(n19866), .B(n19865), .Z(n19875) );
  XOR U24486 ( .A(n19868), .B(n19867), .Z(n19865) );
  XOR U24487 ( .A(y[1166]), .B(x[1166]), .Z(n19867) );
  XOR U24488 ( .A(y[1165]), .B(x[1165]), .Z(n19868) );
  XOR U24489 ( .A(y[1164]), .B(x[1164]), .Z(n19866) );
  XNOR U24490 ( .A(n19859), .B(n19858), .Z(n19861) );
  XNOR U24491 ( .A(n19855), .B(n19854), .Z(n19858) );
  XOR U24492 ( .A(n19857), .B(n19856), .Z(n19854) );
  XOR U24493 ( .A(y[1163]), .B(x[1163]), .Z(n19856) );
  XOR U24494 ( .A(y[1162]), .B(x[1162]), .Z(n19857) );
  XOR U24495 ( .A(y[1161]), .B(x[1161]), .Z(n19855) );
  XOR U24496 ( .A(n19849), .B(n19848), .Z(n19859) );
  XOR U24497 ( .A(n19851), .B(n19850), .Z(n19848) );
  XOR U24498 ( .A(y[1160]), .B(x[1160]), .Z(n19850) );
  XOR U24499 ( .A(y[1159]), .B(x[1159]), .Z(n19851) );
  XOR U24500 ( .A(y[1158]), .B(x[1158]), .Z(n19849) );
  NAND U24501 ( .A(n19912), .B(n19913), .Z(N28509) );
  NAND U24502 ( .A(n19914), .B(n19915), .Z(n19913) );
  NANDN U24503 ( .A(n19916), .B(n19917), .Z(n19915) );
  NANDN U24504 ( .A(n19917), .B(n19916), .Z(n19912) );
  XOR U24505 ( .A(n19916), .B(n19918), .Z(N28508) );
  XNOR U24506 ( .A(n19914), .B(n19917), .Z(n19918) );
  NAND U24507 ( .A(n19919), .B(n19920), .Z(n19917) );
  NAND U24508 ( .A(n19921), .B(n19922), .Z(n19920) );
  NANDN U24509 ( .A(n19923), .B(n19924), .Z(n19922) );
  NANDN U24510 ( .A(n19924), .B(n19923), .Z(n19919) );
  AND U24511 ( .A(n19925), .B(n19926), .Z(n19914) );
  NAND U24512 ( .A(n19927), .B(n19928), .Z(n19926) );
  OR U24513 ( .A(n19929), .B(n19930), .Z(n19928) );
  NAND U24514 ( .A(n19930), .B(n19929), .Z(n19925) );
  IV U24515 ( .A(n19931), .Z(n19930) );
  AND U24516 ( .A(n19932), .B(n19933), .Z(n19916) );
  NAND U24517 ( .A(n19934), .B(n19935), .Z(n19933) );
  NANDN U24518 ( .A(n19936), .B(n19937), .Z(n19935) );
  NANDN U24519 ( .A(n19937), .B(n19936), .Z(n19932) );
  XOR U24520 ( .A(n19929), .B(n19938), .Z(N28507) );
  XOR U24521 ( .A(n19927), .B(n19931), .Z(n19938) );
  XNOR U24522 ( .A(n19924), .B(n19939), .Z(n19931) );
  XNOR U24523 ( .A(n19921), .B(n19923), .Z(n19939) );
  AND U24524 ( .A(n19940), .B(n19941), .Z(n19923) );
  NANDN U24525 ( .A(n19942), .B(n19943), .Z(n19941) );
  NANDN U24526 ( .A(n19944), .B(n19945), .Z(n19943) );
  IV U24527 ( .A(n19946), .Z(n19945) );
  NAND U24528 ( .A(n19946), .B(n19944), .Z(n19940) );
  AND U24529 ( .A(n19947), .B(n19948), .Z(n19921) );
  NAND U24530 ( .A(n19949), .B(n19950), .Z(n19948) );
  OR U24531 ( .A(n19951), .B(n19952), .Z(n19950) );
  NAND U24532 ( .A(n19952), .B(n19951), .Z(n19947) );
  IV U24533 ( .A(n19953), .Z(n19952) );
  NAND U24534 ( .A(n19954), .B(n19955), .Z(n19924) );
  NANDN U24535 ( .A(n19956), .B(n19957), .Z(n19955) );
  NAND U24536 ( .A(n19958), .B(n19959), .Z(n19957) );
  OR U24537 ( .A(n19959), .B(n19958), .Z(n19954) );
  IV U24538 ( .A(n19960), .Z(n19958) );
  AND U24539 ( .A(n19961), .B(n19962), .Z(n19927) );
  NAND U24540 ( .A(n19963), .B(n19964), .Z(n19962) );
  NANDN U24541 ( .A(n19965), .B(n19966), .Z(n19964) );
  NANDN U24542 ( .A(n19966), .B(n19965), .Z(n19961) );
  XOR U24543 ( .A(n19937), .B(n19967), .Z(n19929) );
  XNOR U24544 ( .A(n19934), .B(n19936), .Z(n19967) );
  AND U24545 ( .A(n19968), .B(n19969), .Z(n19936) );
  NANDN U24546 ( .A(n19970), .B(n19971), .Z(n19969) );
  NANDN U24547 ( .A(n19972), .B(n19973), .Z(n19971) );
  IV U24548 ( .A(n19974), .Z(n19973) );
  NAND U24549 ( .A(n19974), .B(n19972), .Z(n19968) );
  AND U24550 ( .A(n19975), .B(n19976), .Z(n19934) );
  NAND U24551 ( .A(n19977), .B(n19978), .Z(n19976) );
  OR U24552 ( .A(n19979), .B(n19980), .Z(n19978) );
  NAND U24553 ( .A(n19980), .B(n19979), .Z(n19975) );
  IV U24554 ( .A(n19981), .Z(n19980) );
  NAND U24555 ( .A(n19982), .B(n19983), .Z(n19937) );
  NANDN U24556 ( .A(n19984), .B(n19985), .Z(n19983) );
  NAND U24557 ( .A(n19986), .B(n19987), .Z(n19985) );
  OR U24558 ( .A(n19987), .B(n19986), .Z(n19982) );
  IV U24559 ( .A(n19988), .Z(n19986) );
  XOR U24560 ( .A(n19963), .B(n19989), .Z(N28506) );
  XNOR U24561 ( .A(n19966), .B(n19965), .Z(n19989) );
  XNOR U24562 ( .A(n19977), .B(n19990), .Z(n19965) );
  XOR U24563 ( .A(n19981), .B(n19979), .Z(n19990) );
  XOR U24564 ( .A(n19987), .B(n19991), .Z(n19979) );
  XOR U24565 ( .A(n19984), .B(n19988), .Z(n19991) );
  NAND U24566 ( .A(n19992), .B(n19993), .Z(n19988) );
  NAND U24567 ( .A(n19994), .B(n19995), .Z(n19993) );
  NAND U24568 ( .A(n19996), .B(n19997), .Z(n19992) );
  AND U24569 ( .A(n19998), .B(n19999), .Z(n19984) );
  NAND U24570 ( .A(n20000), .B(n20001), .Z(n19999) );
  NAND U24571 ( .A(n20002), .B(n20003), .Z(n19998) );
  NANDN U24572 ( .A(n20004), .B(n20005), .Z(n19987) );
  NANDN U24573 ( .A(n20006), .B(n20007), .Z(n19981) );
  XNOR U24574 ( .A(n19972), .B(n20008), .Z(n19977) );
  XOR U24575 ( .A(n19970), .B(n19974), .Z(n20008) );
  NAND U24576 ( .A(n20009), .B(n20010), .Z(n19974) );
  NAND U24577 ( .A(n20011), .B(n20012), .Z(n20010) );
  NAND U24578 ( .A(n20013), .B(n20014), .Z(n20009) );
  AND U24579 ( .A(n20015), .B(n20016), .Z(n19970) );
  NAND U24580 ( .A(n20017), .B(n20018), .Z(n20016) );
  NAND U24581 ( .A(n20019), .B(n20020), .Z(n20015) );
  AND U24582 ( .A(n20021), .B(n20022), .Z(n19972) );
  NAND U24583 ( .A(n20023), .B(n20024), .Z(n19966) );
  XNOR U24584 ( .A(n19949), .B(n20025), .Z(n19963) );
  XOR U24585 ( .A(n19953), .B(n19951), .Z(n20025) );
  XOR U24586 ( .A(n19959), .B(n20026), .Z(n19951) );
  XOR U24587 ( .A(n19956), .B(n19960), .Z(n20026) );
  NAND U24588 ( .A(n20027), .B(n20028), .Z(n19960) );
  NAND U24589 ( .A(n20029), .B(n20030), .Z(n20028) );
  NAND U24590 ( .A(n20031), .B(n20032), .Z(n20027) );
  AND U24591 ( .A(n20033), .B(n20034), .Z(n19956) );
  NAND U24592 ( .A(n20035), .B(n20036), .Z(n20034) );
  NAND U24593 ( .A(n20037), .B(n20038), .Z(n20033) );
  NANDN U24594 ( .A(n20039), .B(n20040), .Z(n19959) );
  NANDN U24595 ( .A(n20041), .B(n20042), .Z(n19953) );
  XNOR U24596 ( .A(n19944), .B(n20043), .Z(n19949) );
  XOR U24597 ( .A(n19942), .B(n19946), .Z(n20043) );
  NAND U24598 ( .A(n20044), .B(n20045), .Z(n19946) );
  NAND U24599 ( .A(n20046), .B(n20047), .Z(n20045) );
  NAND U24600 ( .A(n20048), .B(n20049), .Z(n20044) );
  AND U24601 ( .A(n20050), .B(n20051), .Z(n19942) );
  NAND U24602 ( .A(n20052), .B(n20053), .Z(n20051) );
  NAND U24603 ( .A(n20054), .B(n20055), .Z(n20050) );
  AND U24604 ( .A(n20056), .B(n20057), .Z(n19944) );
  XOR U24605 ( .A(n20024), .B(n20023), .Z(N28505) );
  XNOR U24606 ( .A(n20042), .B(n20041), .Z(n20023) );
  XNOR U24607 ( .A(n20056), .B(n20057), .Z(n20041) );
  XOR U24608 ( .A(n20053), .B(n20052), .Z(n20057) );
  XOR U24609 ( .A(y[1155]), .B(x[1155]), .Z(n20052) );
  XOR U24610 ( .A(n20055), .B(n20054), .Z(n20053) );
  XOR U24611 ( .A(y[1157]), .B(x[1157]), .Z(n20054) );
  XOR U24612 ( .A(y[1156]), .B(x[1156]), .Z(n20055) );
  XOR U24613 ( .A(n20047), .B(n20046), .Z(n20056) );
  XOR U24614 ( .A(n20049), .B(n20048), .Z(n20046) );
  XOR U24615 ( .A(y[1154]), .B(x[1154]), .Z(n20048) );
  XOR U24616 ( .A(y[1153]), .B(x[1153]), .Z(n20049) );
  XOR U24617 ( .A(y[1152]), .B(x[1152]), .Z(n20047) );
  XNOR U24618 ( .A(n20040), .B(n20039), .Z(n20042) );
  XNOR U24619 ( .A(n20036), .B(n20035), .Z(n20039) );
  XOR U24620 ( .A(n20038), .B(n20037), .Z(n20035) );
  XOR U24621 ( .A(y[1151]), .B(x[1151]), .Z(n20037) );
  XOR U24622 ( .A(y[1150]), .B(x[1150]), .Z(n20038) );
  XOR U24623 ( .A(y[1149]), .B(x[1149]), .Z(n20036) );
  XOR U24624 ( .A(n20030), .B(n20029), .Z(n20040) );
  XOR U24625 ( .A(n20032), .B(n20031), .Z(n20029) );
  XOR U24626 ( .A(y[1148]), .B(x[1148]), .Z(n20031) );
  XOR U24627 ( .A(y[1147]), .B(x[1147]), .Z(n20032) );
  XOR U24628 ( .A(y[1146]), .B(x[1146]), .Z(n20030) );
  XNOR U24629 ( .A(n20007), .B(n20006), .Z(n20024) );
  XNOR U24630 ( .A(n20021), .B(n20022), .Z(n20006) );
  XOR U24631 ( .A(n20018), .B(n20017), .Z(n20022) );
  XOR U24632 ( .A(y[1143]), .B(x[1143]), .Z(n20017) );
  XOR U24633 ( .A(n20020), .B(n20019), .Z(n20018) );
  XOR U24634 ( .A(y[1145]), .B(x[1145]), .Z(n20019) );
  XOR U24635 ( .A(y[1144]), .B(x[1144]), .Z(n20020) );
  XOR U24636 ( .A(n20012), .B(n20011), .Z(n20021) );
  XOR U24637 ( .A(n20014), .B(n20013), .Z(n20011) );
  XOR U24638 ( .A(y[1142]), .B(x[1142]), .Z(n20013) );
  XOR U24639 ( .A(y[1141]), .B(x[1141]), .Z(n20014) );
  XOR U24640 ( .A(y[1140]), .B(x[1140]), .Z(n20012) );
  XNOR U24641 ( .A(n20005), .B(n20004), .Z(n20007) );
  XNOR U24642 ( .A(n20001), .B(n20000), .Z(n20004) );
  XOR U24643 ( .A(n20003), .B(n20002), .Z(n20000) );
  XOR U24644 ( .A(y[1139]), .B(x[1139]), .Z(n20002) );
  XOR U24645 ( .A(y[1138]), .B(x[1138]), .Z(n20003) );
  XOR U24646 ( .A(y[1137]), .B(x[1137]), .Z(n20001) );
  XOR U24647 ( .A(n19995), .B(n19994), .Z(n20005) );
  XOR U24648 ( .A(n19997), .B(n19996), .Z(n19994) );
  XOR U24649 ( .A(y[1136]), .B(x[1136]), .Z(n19996) );
  XOR U24650 ( .A(y[1135]), .B(x[1135]), .Z(n19997) );
  XOR U24651 ( .A(y[1134]), .B(x[1134]), .Z(n19995) );
  NAND U24652 ( .A(n20058), .B(n20059), .Z(N28497) );
  NAND U24653 ( .A(n20060), .B(n20061), .Z(n20059) );
  NANDN U24654 ( .A(n20062), .B(n20063), .Z(n20061) );
  NANDN U24655 ( .A(n20063), .B(n20062), .Z(n20058) );
  XOR U24656 ( .A(n20062), .B(n20064), .Z(N28496) );
  XNOR U24657 ( .A(n20060), .B(n20063), .Z(n20064) );
  NAND U24658 ( .A(n20065), .B(n20066), .Z(n20063) );
  NAND U24659 ( .A(n20067), .B(n20068), .Z(n20066) );
  NANDN U24660 ( .A(n20069), .B(n20070), .Z(n20068) );
  NANDN U24661 ( .A(n20070), .B(n20069), .Z(n20065) );
  AND U24662 ( .A(n20071), .B(n20072), .Z(n20060) );
  NAND U24663 ( .A(n20073), .B(n20074), .Z(n20072) );
  OR U24664 ( .A(n20075), .B(n20076), .Z(n20074) );
  NAND U24665 ( .A(n20076), .B(n20075), .Z(n20071) );
  IV U24666 ( .A(n20077), .Z(n20076) );
  AND U24667 ( .A(n20078), .B(n20079), .Z(n20062) );
  NAND U24668 ( .A(n20080), .B(n20081), .Z(n20079) );
  NANDN U24669 ( .A(n20082), .B(n20083), .Z(n20081) );
  NANDN U24670 ( .A(n20083), .B(n20082), .Z(n20078) );
  XOR U24671 ( .A(n20075), .B(n20084), .Z(N28495) );
  XOR U24672 ( .A(n20073), .B(n20077), .Z(n20084) );
  XNOR U24673 ( .A(n20070), .B(n20085), .Z(n20077) );
  XNOR U24674 ( .A(n20067), .B(n20069), .Z(n20085) );
  AND U24675 ( .A(n20086), .B(n20087), .Z(n20069) );
  NANDN U24676 ( .A(n20088), .B(n20089), .Z(n20087) );
  NANDN U24677 ( .A(n20090), .B(n20091), .Z(n20089) );
  IV U24678 ( .A(n20092), .Z(n20091) );
  NAND U24679 ( .A(n20092), .B(n20090), .Z(n20086) );
  AND U24680 ( .A(n20093), .B(n20094), .Z(n20067) );
  NAND U24681 ( .A(n20095), .B(n20096), .Z(n20094) );
  OR U24682 ( .A(n20097), .B(n20098), .Z(n20096) );
  NAND U24683 ( .A(n20098), .B(n20097), .Z(n20093) );
  IV U24684 ( .A(n20099), .Z(n20098) );
  NAND U24685 ( .A(n20100), .B(n20101), .Z(n20070) );
  NANDN U24686 ( .A(n20102), .B(n20103), .Z(n20101) );
  NAND U24687 ( .A(n20104), .B(n20105), .Z(n20103) );
  OR U24688 ( .A(n20105), .B(n20104), .Z(n20100) );
  IV U24689 ( .A(n20106), .Z(n20104) );
  AND U24690 ( .A(n20107), .B(n20108), .Z(n20073) );
  NAND U24691 ( .A(n20109), .B(n20110), .Z(n20108) );
  NANDN U24692 ( .A(n20111), .B(n20112), .Z(n20110) );
  NANDN U24693 ( .A(n20112), .B(n20111), .Z(n20107) );
  XOR U24694 ( .A(n20083), .B(n20113), .Z(n20075) );
  XNOR U24695 ( .A(n20080), .B(n20082), .Z(n20113) );
  AND U24696 ( .A(n20114), .B(n20115), .Z(n20082) );
  NANDN U24697 ( .A(n20116), .B(n20117), .Z(n20115) );
  NANDN U24698 ( .A(n20118), .B(n20119), .Z(n20117) );
  IV U24699 ( .A(n20120), .Z(n20119) );
  NAND U24700 ( .A(n20120), .B(n20118), .Z(n20114) );
  AND U24701 ( .A(n20121), .B(n20122), .Z(n20080) );
  NAND U24702 ( .A(n20123), .B(n20124), .Z(n20122) );
  OR U24703 ( .A(n20125), .B(n20126), .Z(n20124) );
  NAND U24704 ( .A(n20126), .B(n20125), .Z(n20121) );
  IV U24705 ( .A(n20127), .Z(n20126) );
  NAND U24706 ( .A(n20128), .B(n20129), .Z(n20083) );
  NANDN U24707 ( .A(n20130), .B(n20131), .Z(n20129) );
  NAND U24708 ( .A(n20132), .B(n20133), .Z(n20131) );
  OR U24709 ( .A(n20133), .B(n20132), .Z(n20128) );
  IV U24710 ( .A(n20134), .Z(n20132) );
  XOR U24711 ( .A(n20109), .B(n20135), .Z(N28494) );
  XNOR U24712 ( .A(n20112), .B(n20111), .Z(n20135) );
  XNOR U24713 ( .A(n20123), .B(n20136), .Z(n20111) );
  XOR U24714 ( .A(n20127), .B(n20125), .Z(n20136) );
  XOR U24715 ( .A(n20133), .B(n20137), .Z(n20125) );
  XOR U24716 ( .A(n20130), .B(n20134), .Z(n20137) );
  NAND U24717 ( .A(n20138), .B(n20139), .Z(n20134) );
  NAND U24718 ( .A(n20140), .B(n20141), .Z(n20139) );
  NAND U24719 ( .A(n20142), .B(n20143), .Z(n20138) );
  AND U24720 ( .A(n20144), .B(n20145), .Z(n20130) );
  NAND U24721 ( .A(n20146), .B(n20147), .Z(n20145) );
  NAND U24722 ( .A(n20148), .B(n20149), .Z(n20144) );
  NANDN U24723 ( .A(n20150), .B(n20151), .Z(n20133) );
  NANDN U24724 ( .A(n20152), .B(n20153), .Z(n20127) );
  XNOR U24725 ( .A(n20118), .B(n20154), .Z(n20123) );
  XOR U24726 ( .A(n20116), .B(n20120), .Z(n20154) );
  NAND U24727 ( .A(n20155), .B(n20156), .Z(n20120) );
  NAND U24728 ( .A(n20157), .B(n20158), .Z(n20156) );
  NAND U24729 ( .A(n20159), .B(n20160), .Z(n20155) );
  AND U24730 ( .A(n20161), .B(n20162), .Z(n20116) );
  NAND U24731 ( .A(n20163), .B(n20164), .Z(n20162) );
  NAND U24732 ( .A(n20165), .B(n20166), .Z(n20161) );
  AND U24733 ( .A(n20167), .B(n20168), .Z(n20118) );
  NAND U24734 ( .A(n20169), .B(n20170), .Z(n20112) );
  XNOR U24735 ( .A(n20095), .B(n20171), .Z(n20109) );
  XOR U24736 ( .A(n20099), .B(n20097), .Z(n20171) );
  XOR U24737 ( .A(n20105), .B(n20172), .Z(n20097) );
  XOR U24738 ( .A(n20102), .B(n20106), .Z(n20172) );
  NAND U24739 ( .A(n20173), .B(n20174), .Z(n20106) );
  NAND U24740 ( .A(n20175), .B(n20176), .Z(n20174) );
  NAND U24741 ( .A(n20177), .B(n20178), .Z(n20173) );
  AND U24742 ( .A(n20179), .B(n20180), .Z(n20102) );
  NAND U24743 ( .A(n20181), .B(n20182), .Z(n20180) );
  NAND U24744 ( .A(n20183), .B(n20184), .Z(n20179) );
  NANDN U24745 ( .A(n20185), .B(n20186), .Z(n20105) );
  NANDN U24746 ( .A(n20187), .B(n20188), .Z(n20099) );
  XNOR U24747 ( .A(n20090), .B(n20189), .Z(n20095) );
  XOR U24748 ( .A(n20088), .B(n20092), .Z(n20189) );
  NAND U24749 ( .A(n20190), .B(n20191), .Z(n20092) );
  NAND U24750 ( .A(n20192), .B(n20193), .Z(n20191) );
  NAND U24751 ( .A(n20194), .B(n20195), .Z(n20190) );
  AND U24752 ( .A(n20196), .B(n20197), .Z(n20088) );
  NAND U24753 ( .A(n20198), .B(n20199), .Z(n20197) );
  NAND U24754 ( .A(n20200), .B(n20201), .Z(n20196) );
  AND U24755 ( .A(n20202), .B(n20203), .Z(n20090) );
  XOR U24756 ( .A(n20170), .B(n20169), .Z(N28493) );
  XNOR U24757 ( .A(n20188), .B(n20187), .Z(n20169) );
  XNOR U24758 ( .A(n20202), .B(n20203), .Z(n20187) );
  XOR U24759 ( .A(n20199), .B(n20198), .Z(n20203) );
  XOR U24760 ( .A(y[1131]), .B(x[1131]), .Z(n20198) );
  XOR U24761 ( .A(n20201), .B(n20200), .Z(n20199) );
  XOR U24762 ( .A(y[1133]), .B(x[1133]), .Z(n20200) );
  XOR U24763 ( .A(y[1132]), .B(x[1132]), .Z(n20201) );
  XOR U24764 ( .A(n20193), .B(n20192), .Z(n20202) );
  XOR U24765 ( .A(n20195), .B(n20194), .Z(n20192) );
  XOR U24766 ( .A(y[1130]), .B(x[1130]), .Z(n20194) );
  XOR U24767 ( .A(y[1129]), .B(x[1129]), .Z(n20195) );
  XOR U24768 ( .A(y[1128]), .B(x[1128]), .Z(n20193) );
  XNOR U24769 ( .A(n20186), .B(n20185), .Z(n20188) );
  XNOR U24770 ( .A(n20182), .B(n20181), .Z(n20185) );
  XOR U24771 ( .A(n20184), .B(n20183), .Z(n20181) );
  XOR U24772 ( .A(y[1127]), .B(x[1127]), .Z(n20183) );
  XOR U24773 ( .A(y[1126]), .B(x[1126]), .Z(n20184) );
  XOR U24774 ( .A(y[1125]), .B(x[1125]), .Z(n20182) );
  XOR U24775 ( .A(n20176), .B(n20175), .Z(n20186) );
  XOR U24776 ( .A(n20178), .B(n20177), .Z(n20175) );
  XOR U24777 ( .A(y[1124]), .B(x[1124]), .Z(n20177) );
  XOR U24778 ( .A(y[1123]), .B(x[1123]), .Z(n20178) );
  XOR U24779 ( .A(y[1122]), .B(x[1122]), .Z(n20176) );
  XNOR U24780 ( .A(n20153), .B(n20152), .Z(n20170) );
  XNOR U24781 ( .A(n20167), .B(n20168), .Z(n20152) );
  XOR U24782 ( .A(n20164), .B(n20163), .Z(n20168) );
  XOR U24783 ( .A(y[1119]), .B(x[1119]), .Z(n20163) );
  XOR U24784 ( .A(n20166), .B(n20165), .Z(n20164) );
  XOR U24785 ( .A(y[1121]), .B(x[1121]), .Z(n20165) );
  XOR U24786 ( .A(y[1120]), .B(x[1120]), .Z(n20166) );
  XOR U24787 ( .A(n20158), .B(n20157), .Z(n20167) );
  XOR U24788 ( .A(n20160), .B(n20159), .Z(n20157) );
  XOR U24789 ( .A(y[1118]), .B(x[1118]), .Z(n20159) );
  XOR U24790 ( .A(y[1117]), .B(x[1117]), .Z(n20160) );
  XOR U24791 ( .A(y[1116]), .B(x[1116]), .Z(n20158) );
  XNOR U24792 ( .A(n20151), .B(n20150), .Z(n20153) );
  XNOR U24793 ( .A(n20147), .B(n20146), .Z(n20150) );
  XOR U24794 ( .A(n20149), .B(n20148), .Z(n20146) );
  XOR U24795 ( .A(y[1115]), .B(x[1115]), .Z(n20148) );
  XOR U24796 ( .A(y[1114]), .B(x[1114]), .Z(n20149) );
  XOR U24797 ( .A(y[1113]), .B(x[1113]), .Z(n20147) );
  XOR U24798 ( .A(n20141), .B(n20140), .Z(n20151) );
  XOR U24799 ( .A(n20143), .B(n20142), .Z(n20140) );
  XOR U24800 ( .A(y[1112]), .B(x[1112]), .Z(n20142) );
  XOR U24801 ( .A(y[1111]), .B(x[1111]), .Z(n20143) );
  XOR U24802 ( .A(y[1110]), .B(x[1110]), .Z(n20141) );
  NAND U24803 ( .A(n20204), .B(n20205), .Z(N28485) );
  NAND U24804 ( .A(n20206), .B(n20207), .Z(n20205) );
  NANDN U24805 ( .A(n20208), .B(n20209), .Z(n20207) );
  NANDN U24806 ( .A(n20209), .B(n20208), .Z(n20204) );
  XOR U24807 ( .A(n20208), .B(n20210), .Z(N28484) );
  XNOR U24808 ( .A(n20206), .B(n20209), .Z(n20210) );
  NAND U24809 ( .A(n20211), .B(n20212), .Z(n20209) );
  NAND U24810 ( .A(n20213), .B(n20214), .Z(n20212) );
  NANDN U24811 ( .A(n20215), .B(n20216), .Z(n20214) );
  NANDN U24812 ( .A(n20216), .B(n20215), .Z(n20211) );
  AND U24813 ( .A(n20217), .B(n20218), .Z(n20206) );
  NAND U24814 ( .A(n20219), .B(n20220), .Z(n20218) );
  OR U24815 ( .A(n20221), .B(n20222), .Z(n20220) );
  NAND U24816 ( .A(n20222), .B(n20221), .Z(n20217) );
  IV U24817 ( .A(n20223), .Z(n20222) );
  AND U24818 ( .A(n20224), .B(n20225), .Z(n20208) );
  NAND U24819 ( .A(n20226), .B(n20227), .Z(n20225) );
  NANDN U24820 ( .A(n20228), .B(n20229), .Z(n20227) );
  NANDN U24821 ( .A(n20229), .B(n20228), .Z(n20224) );
  XOR U24822 ( .A(n20221), .B(n20230), .Z(N28483) );
  XOR U24823 ( .A(n20219), .B(n20223), .Z(n20230) );
  XNOR U24824 ( .A(n20216), .B(n20231), .Z(n20223) );
  XNOR U24825 ( .A(n20213), .B(n20215), .Z(n20231) );
  AND U24826 ( .A(n20232), .B(n20233), .Z(n20215) );
  NANDN U24827 ( .A(n20234), .B(n20235), .Z(n20233) );
  NANDN U24828 ( .A(n20236), .B(n20237), .Z(n20235) );
  IV U24829 ( .A(n20238), .Z(n20237) );
  NAND U24830 ( .A(n20238), .B(n20236), .Z(n20232) );
  AND U24831 ( .A(n20239), .B(n20240), .Z(n20213) );
  NAND U24832 ( .A(n20241), .B(n20242), .Z(n20240) );
  OR U24833 ( .A(n20243), .B(n20244), .Z(n20242) );
  NAND U24834 ( .A(n20244), .B(n20243), .Z(n20239) );
  IV U24835 ( .A(n20245), .Z(n20244) );
  NAND U24836 ( .A(n20246), .B(n20247), .Z(n20216) );
  NANDN U24837 ( .A(n20248), .B(n20249), .Z(n20247) );
  NAND U24838 ( .A(n20250), .B(n20251), .Z(n20249) );
  OR U24839 ( .A(n20251), .B(n20250), .Z(n20246) );
  IV U24840 ( .A(n20252), .Z(n20250) );
  AND U24841 ( .A(n20253), .B(n20254), .Z(n20219) );
  NAND U24842 ( .A(n20255), .B(n20256), .Z(n20254) );
  NANDN U24843 ( .A(n20257), .B(n20258), .Z(n20256) );
  NANDN U24844 ( .A(n20258), .B(n20257), .Z(n20253) );
  XOR U24845 ( .A(n20229), .B(n20259), .Z(n20221) );
  XNOR U24846 ( .A(n20226), .B(n20228), .Z(n20259) );
  AND U24847 ( .A(n20260), .B(n20261), .Z(n20228) );
  NANDN U24848 ( .A(n20262), .B(n20263), .Z(n20261) );
  NANDN U24849 ( .A(n20264), .B(n20265), .Z(n20263) );
  IV U24850 ( .A(n20266), .Z(n20265) );
  NAND U24851 ( .A(n20266), .B(n20264), .Z(n20260) );
  AND U24852 ( .A(n20267), .B(n20268), .Z(n20226) );
  NAND U24853 ( .A(n20269), .B(n20270), .Z(n20268) );
  OR U24854 ( .A(n20271), .B(n20272), .Z(n20270) );
  NAND U24855 ( .A(n20272), .B(n20271), .Z(n20267) );
  IV U24856 ( .A(n20273), .Z(n20272) );
  NAND U24857 ( .A(n20274), .B(n20275), .Z(n20229) );
  NANDN U24858 ( .A(n20276), .B(n20277), .Z(n20275) );
  NAND U24859 ( .A(n20278), .B(n20279), .Z(n20277) );
  OR U24860 ( .A(n20279), .B(n20278), .Z(n20274) );
  IV U24861 ( .A(n20280), .Z(n20278) );
  XOR U24862 ( .A(n20255), .B(n20281), .Z(N28482) );
  XNOR U24863 ( .A(n20258), .B(n20257), .Z(n20281) );
  XNOR U24864 ( .A(n20269), .B(n20282), .Z(n20257) );
  XOR U24865 ( .A(n20273), .B(n20271), .Z(n20282) );
  XOR U24866 ( .A(n20279), .B(n20283), .Z(n20271) );
  XOR U24867 ( .A(n20276), .B(n20280), .Z(n20283) );
  NAND U24868 ( .A(n20284), .B(n20285), .Z(n20280) );
  NAND U24869 ( .A(n20286), .B(n20287), .Z(n20285) );
  NAND U24870 ( .A(n20288), .B(n20289), .Z(n20284) );
  AND U24871 ( .A(n20290), .B(n20291), .Z(n20276) );
  NAND U24872 ( .A(n20292), .B(n20293), .Z(n20291) );
  NAND U24873 ( .A(n20294), .B(n20295), .Z(n20290) );
  NANDN U24874 ( .A(n20296), .B(n20297), .Z(n20279) );
  NANDN U24875 ( .A(n20298), .B(n20299), .Z(n20273) );
  XNOR U24876 ( .A(n20264), .B(n20300), .Z(n20269) );
  XOR U24877 ( .A(n20262), .B(n20266), .Z(n20300) );
  NAND U24878 ( .A(n20301), .B(n20302), .Z(n20266) );
  NAND U24879 ( .A(n20303), .B(n20304), .Z(n20302) );
  NAND U24880 ( .A(n20305), .B(n20306), .Z(n20301) );
  AND U24881 ( .A(n20307), .B(n20308), .Z(n20262) );
  NAND U24882 ( .A(n20309), .B(n20310), .Z(n20308) );
  NAND U24883 ( .A(n20311), .B(n20312), .Z(n20307) );
  AND U24884 ( .A(n20313), .B(n20314), .Z(n20264) );
  NAND U24885 ( .A(n20315), .B(n20316), .Z(n20258) );
  XNOR U24886 ( .A(n20241), .B(n20317), .Z(n20255) );
  XOR U24887 ( .A(n20245), .B(n20243), .Z(n20317) );
  XOR U24888 ( .A(n20251), .B(n20318), .Z(n20243) );
  XOR U24889 ( .A(n20248), .B(n20252), .Z(n20318) );
  NAND U24890 ( .A(n20319), .B(n20320), .Z(n20252) );
  NAND U24891 ( .A(n20321), .B(n20322), .Z(n20320) );
  NAND U24892 ( .A(n20323), .B(n20324), .Z(n20319) );
  AND U24893 ( .A(n20325), .B(n20326), .Z(n20248) );
  NAND U24894 ( .A(n20327), .B(n20328), .Z(n20326) );
  NAND U24895 ( .A(n20329), .B(n20330), .Z(n20325) );
  NANDN U24896 ( .A(n20331), .B(n20332), .Z(n20251) );
  NANDN U24897 ( .A(n20333), .B(n20334), .Z(n20245) );
  XNOR U24898 ( .A(n20236), .B(n20335), .Z(n20241) );
  XOR U24899 ( .A(n20234), .B(n20238), .Z(n20335) );
  NAND U24900 ( .A(n20336), .B(n20337), .Z(n20238) );
  NAND U24901 ( .A(n20338), .B(n20339), .Z(n20337) );
  NAND U24902 ( .A(n20340), .B(n20341), .Z(n20336) );
  AND U24903 ( .A(n20342), .B(n20343), .Z(n20234) );
  NAND U24904 ( .A(n20344), .B(n20345), .Z(n20343) );
  NAND U24905 ( .A(n20346), .B(n20347), .Z(n20342) );
  AND U24906 ( .A(n20348), .B(n20349), .Z(n20236) );
  XOR U24907 ( .A(n20316), .B(n20315), .Z(N28481) );
  XNOR U24908 ( .A(n20334), .B(n20333), .Z(n20315) );
  XNOR U24909 ( .A(n20348), .B(n20349), .Z(n20333) );
  XOR U24910 ( .A(n20345), .B(n20344), .Z(n20349) );
  XOR U24911 ( .A(y[1107]), .B(x[1107]), .Z(n20344) );
  XOR U24912 ( .A(n20347), .B(n20346), .Z(n20345) );
  XOR U24913 ( .A(y[1109]), .B(x[1109]), .Z(n20346) );
  XOR U24914 ( .A(y[1108]), .B(x[1108]), .Z(n20347) );
  XOR U24915 ( .A(n20339), .B(n20338), .Z(n20348) );
  XOR U24916 ( .A(n20341), .B(n20340), .Z(n20338) );
  XOR U24917 ( .A(y[1106]), .B(x[1106]), .Z(n20340) );
  XOR U24918 ( .A(y[1105]), .B(x[1105]), .Z(n20341) );
  XOR U24919 ( .A(y[1104]), .B(x[1104]), .Z(n20339) );
  XNOR U24920 ( .A(n20332), .B(n20331), .Z(n20334) );
  XNOR U24921 ( .A(n20328), .B(n20327), .Z(n20331) );
  XOR U24922 ( .A(n20330), .B(n20329), .Z(n20327) );
  XOR U24923 ( .A(y[1103]), .B(x[1103]), .Z(n20329) );
  XOR U24924 ( .A(y[1102]), .B(x[1102]), .Z(n20330) );
  XOR U24925 ( .A(y[1101]), .B(x[1101]), .Z(n20328) );
  XOR U24926 ( .A(n20322), .B(n20321), .Z(n20332) );
  XOR U24927 ( .A(n20324), .B(n20323), .Z(n20321) );
  XOR U24928 ( .A(y[1100]), .B(x[1100]), .Z(n20323) );
  XOR U24929 ( .A(y[1099]), .B(x[1099]), .Z(n20324) );
  XOR U24930 ( .A(y[1098]), .B(x[1098]), .Z(n20322) );
  XNOR U24931 ( .A(n20299), .B(n20298), .Z(n20316) );
  XNOR U24932 ( .A(n20313), .B(n20314), .Z(n20298) );
  XOR U24933 ( .A(n20310), .B(n20309), .Z(n20314) );
  XOR U24934 ( .A(y[1095]), .B(x[1095]), .Z(n20309) );
  XOR U24935 ( .A(n20312), .B(n20311), .Z(n20310) );
  XOR U24936 ( .A(y[1097]), .B(x[1097]), .Z(n20311) );
  XOR U24937 ( .A(y[1096]), .B(x[1096]), .Z(n20312) );
  XOR U24938 ( .A(n20304), .B(n20303), .Z(n20313) );
  XOR U24939 ( .A(n20306), .B(n20305), .Z(n20303) );
  XOR U24940 ( .A(y[1094]), .B(x[1094]), .Z(n20305) );
  XOR U24941 ( .A(y[1093]), .B(x[1093]), .Z(n20306) );
  XOR U24942 ( .A(y[1092]), .B(x[1092]), .Z(n20304) );
  XNOR U24943 ( .A(n20297), .B(n20296), .Z(n20299) );
  XNOR U24944 ( .A(n20293), .B(n20292), .Z(n20296) );
  XOR U24945 ( .A(n20295), .B(n20294), .Z(n20292) );
  XOR U24946 ( .A(y[1091]), .B(x[1091]), .Z(n20294) );
  XOR U24947 ( .A(y[1090]), .B(x[1090]), .Z(n20295) );
  XOR U24948 ( .A(y[1089]), .B(x[1089]), .Z(n20293) );
  XOR U24949 ( .A(n20287), .B(n20286), .Z(n20297) );
  XOR U24950 ( .A(n20289), .B(n20288), .Z(n20286) );
  XOR U24951 ( .A(y[1088]), .B(x[1088]), .Z(n20288) );
  XOR U24952 ( .A(y[1087]), .B(x[1087]), .Z(n20289) );
  XOR U24953 ( .A(y[1086]), .B(x[1086]), .Z(n20287) );
  NAND U24954 ( .A(n20350), .B(n20351), .Z(N28473) );
  NAND U24955 ( .A(n20352), .B(n20353), .Z(n20351) );
  NANDN U24956 ( .A(n20354), .B(n20355), .Z(n20353) );
  NANDN U24957 ( .A(n20355), .B(n20354), .Z(n20350) );
  XOR U24958 ( .A(n20354), .B(n20356), .Z(N28472) );
  XNOR U24959 ( .A(n20352), .B(n20355), .Z(n20356) );
  NAND U24960 ( .A(n20357), .B(n20358), .Z(n20355) );
  NAND U24961 ( .A(n20359), .B(n20360), .Z(n20358) );
  NANDN U24962 ( .A(n20361), .B(n20362), .Z(n20360) );
  NANDN U24963 ( .A(n20362), .B(n20361), .Z(n20357) );
  AND U24964 ( .A(n20363), .B(n20364), .Z(n20352) );
  NAND U24965 ( .A(n20365), .B(n20366), .Z(n20364) );
  OR U24966 ( .A(n20367), .B(n20368), .Z(n20366) );
  NAND U24967 ( .A(n20368), .B(n20367), .Z(n20363) );
  IV U24968 ( .A(n20369), .Z(n20368) );
  AND U24969 ( .A(n20370), .B(n20371), .Z(n20354) );
  NAND U24970 ( .A(n20372), .B(n20373), .Z(n20371) );
  NANDN U24971 ( .A(n20374), .B(n20375), .Z(n20373) );
  NANDN U24972 ( .A(n20375), .B(n20374), .Z(n20370) );
  XOR U24973 ( .A(n20367), .B(n20376), .Z(N28471) );
  XOR U24974 ( .A(n20365), .B(n20369), .Z(n20376) );
  XNOR U24975 ( .A(n20362), .B(n20377), .Z(n20369) );
  XNOR U24976 ( .A(n20359), .B(n20361), .Z(n20377) );
  AND U24977 ( .A(n20378), .B(n20379), .Z(n20361) );
  NANDN U24978 ( .A(n20380), .B(n20381), .Z(n20379) );
  NANDN U24979 ( .A(n20382), .B(n20383), .Z(n20381) );
  IV U24980 ( .A(n20384), .Z(n20383) );
  NAND U24981 ( .A(n20384), .B(n20382), .Z(n20378) );
  AND U24982 ( .A(n20385), .B(n20386), .Z(n20359) );
  NAND U24983 ( .A(n20387), .B(n20388), .Z(n20386) );
  OR U24984 ( .A(n20389), .B(n20390), .Z(n20388) );
  NAND U24985 ( .A(n20390), .B(n20389), .Z(n20385) );
  IV U24986 ( .A(n20391), .Z(n20390) );
  NAND U24987 ( .A(n20392), .B(n20393), .Z(n20362) );
  NANDN U24988 ( .A(n20394), .B(n20395), .Z(n20393) );
  NAND U24989 ( .A(n20396), .B(n20397), .Z(n20395) );
  OR U24990 ( .A(n20397), .B(n20396), .Z(n20392) );
  IV U24991 ( .A(n20398), .Z(n20396) );
  AND U24992 ( .A(n20399), .B(n20400), .Z(n20365) );
  NAND U24993 ( .A(n20401), .B(n20402), .Z(n20400) );
  NANDN U24994 ( .A(n20403), .B(n20404), .Z(n20402) );
  NANDN U24995 ( .A(n20404), .B(n20403), .Z(n20399) );
  XOR U24996 ( .A(n20375), .B(n20405), .Z(n20367) );
  XNOR U24997 ( .A(n20372), .B(n20374), .Z(n20405) );
  AND U24998 ( .A(n20406), .B(n20407), .Z(n20374) );
  NANDN U24999 ( .A(n20408), .B(n20409), .Z(n20407) );
  NANDN U25000 ( .A(n20410), .B(n20411), .Z(n20409) );
  IV U25001 ( .A(n20412), .Z(n20411) );
  NAND U25002 ( .A(n20412), .B(n20410), .Z(n20406) );
  AND U25003 ( .A(n20413), .B(n20414), .Z(n20372) );
  NAND U25004 ( .A(n20415), .B(n20416), .Z(n20414) );
  OR U25005 ( .A(n20417), .B(n20418), .Z(n20416) );
  NAND U25006 ( .A(n20418), .B(n20417), .Z(n20413) );
  IV U25007 ( .A(n20419), .Z(n20418) );
  NAND U25008 ( .A(n20420), .B(n20421), .Z(n20375) );
  NANDN U25009 ( .A(n20422), .B(n20423), .Z(n20421) );
  NAND U25010 ( .A(n20424), .B(n20425), .Z(n20423) );
  OR U25011 ( .A(n20425), .B(n20424), .Z(n20420) );
  IV U25012 ( .A(n20426), .Z(n20424) );
  XOR U25013 ( .A(n20401), .B(n20427), .Z(N28470) );
  XNOR U25014 ( .A(n20404), .B(n20403), .Z(n20427) );
  XNOR U25015 ( .A(n20415), .B(n20428), .Z(n20403) );
  XOR U25016 ( .A(n20419), .B(n20417), .Z(n20428) );
  XOR U25017 ( .A(n20425), .B(n20429), .Z(n20417) );
  XOR U25018 ( .A(n20422), .B(n20426), .Z(n20429) );
  NAND U25019 ( .A(n20430), .B(n20431), .Z(n20426) );
  NAND U25020 ( .A(n20432), .B(n20433), .Z(n20431) );
  NAND U25021 ( .A(n20434), .B(n20435), .Z(n20430) );
  AND U25022 ( .A(n20436), .B(n20437), .Z(n20422) );
  NAND U25023 ( .A(n20438), .B(n20439), .Z(n20437) );
  NAND U25024 ( .A(n20440), .B(n20441), .Z(n20436) );
  NANDN U25025 ( .A(n20442), .B(n20443), .Z(n20425) );
  NANDN U25026 ( .A(n20444), .B(n20445), .Z(n20419) );
  XNOR U25027 ( .A(n20410), .B(n20446), .Z(n20415) );
  XOR U25028 ( .A(n20408), .B(n20412), .Z(n20446) );
  NAND U25029 ( .A(n20447), .B(n20448), .Z(n20412) );
  NAND U25030 ( .A(n20449), .B(n20450), .Z(n20448) );
  NAND U25031 ( .A(n20451), .B(n20452), .Z(n20447) );
  AND U25032 ( .A(n20453), .B(n20454), .Z(n20408) );
  NAND U25033 ( .A(n20455), .B(n20456), .Z(n20454) );
  NAND U25034 ( .A(n20457), .B(n20458), .Z(n20453) );
  AND U25035 ( .A(n20459), .B(n20460), .Z(n20410) );
  NAND U25036 ( .A(n20461), .B(n20462), .Z(n20404) );
  XNOR U25037 ( .A(n20387), .B(n20463), .Z(n20401) );
  XOR U25038 ( .A(n20391), .B(n20389), .Z(n20463) );
  XOR U25039 ( .A(n20397), .B(n20464), .Z(n20389) );
  XOR U25040 ( .A(n20394), .B(n20398), .Z(n20464) );
  NAND U25041 ( .A(n20465), .B(n20466), .Z(n20398) );
  NAND U25042 ( .A(n20467), .B(n20468), .Z(n20466) );
  NAND U25043 ( .A(n20469), .B(n20470), .Z(n20465) );
  AND U25044 ( .A(n20471), .B(n20472), .Z(n20394) );
  NAND U25045 ( .A(n20473), .B(n20474), .Z(n20472) );
  NAND U25046 ( .A(n20475), .B(n20476), .Z(n20471) );
  NANDN U25047 ( .A(n20477), .B(n20478), .Z(n20397) );
  NANDN U25048 ( .A(n20479), .B(n20480), .Z(n20391) );
  XNOR U25049 ( .A(n20382), .B(n20481), .Z(n20387) );
  XOR U25050 ( .A(n20380), .B(n20384), .Z(n20481) );
  NAND U25051 ( .A(n20482), .B(n20483), .Z(n20384) );
  NAND U25052 ( .A(n20484), .B(n20485), .Z(n20483) );
  NAND U25053 ( .A(n20486), .B(n20487), .Z(n20482) );
  AND U25054 ( .A(n20488), .B(n20489), .Z(n20380) );
  NAND U25055 ( .A(n20490), .B(n20491), .Z(n20489) );
  NAND U25056 ( .A(n20492), .B(n20493), .Z(n20488) );
  AND U25057 ( .A(n20494), .B(n20495), .Z(n20382) );
  XOR U25058 ( .A(n20462), .B(n20461), .Z(N28469) );
  XNOR U25059 ( .A(n20480), .B(n20479), .Z(n20461) );
  XNOR U25060 ( .A(n20494), .B(n20495), .Z(n20479) );
  XOR U25061 ( .A(n20491), .B(n20490), .Z(n20495) );
  XOR U25062 ( .A(y[1083]), .B(x[1083]), .Z(n20490) );
  XOR U25063 ( .A(n20493), .B(n20492), .Z(n20491) );
  XOR U25064 ( .A(y[1085]), .B(x[1085]), .Z(n20492) );
  XOR U25065 ( .A(y[1084]), .B(x[1084]), .Z(n20493) );
  XOR U25066 ( .A(n20485), .B(n20484), .Z(n20494) );
  XOR U25067 ( .A(n20487), .B(n20486), .Z(n20484) );
  XOR U25068 ( .A(y[1082]), .B(x[1082]), .Z(n20486) );
  XOR U25069 ( .A(y[1081]), .B(x[1081]), .Z(n20487) );
  XOR U25070 ( .A(y[1080]), .B(x[1080]), .Z(n20485) );
  XNOR U25071 ( .A(n20478), .B(n20477), .Z(n20480) );
  XNOR U25072 ( .A(n20474), .B(n20473), .Z(n20477) );
  XOR U25073 ( .A(n20476), .B(n20475), .Z(n20473) );
  XOR U25074 ( .A(y[1079]), .B(x[1079]), .Z(n20475) );
  XOR U25075 ( .A(y[1078]), .B(x[1078]), .Z(n20476) );
  XOR U25076 ( .A(y[1077]), .B(x[1077]), .Z(n20474) );
  XOR U25077 ( .A(n20468), .B(n20467), .Z(n20478) );
  XOR U25078 ( .A(n20470), .B(n20469), .Z(n20467) );
  XOR U25079 ( .A(y[1076]), .B(x[1076]), .Z(n20469) );
  XOR U25080 ( .A(y[1075]), .B(x[1075]), .Z(n20470) );
  XOR U25081 ( .A(y[1074]), .B(x[1074]), .Z(n20468) );
  XNOR U25082 ( .A(n20445), .B(n20444), .Z(n20462) );
  XNOR U25083 ( .A(n20459), .B(n20460), .Z(n20444) );
  XOR U25084 ( .A(n20456), .B(n20455), .Z(n20460) );
  XOR U25085 ( .A(y[1071]), .B(x[1071]), .Z(n20455) );
  XOR U25086 ( .A(n20458), .B(n20457), .Z(n20456) );
  XOR U25087 ( .A(y[1073]), .B(x[1073]), .Z(n20457) );
  XOR U25088 ( .A(y[1072]), .B(x[1072]), .Z(n20458) );
  XOR U25089 ( .A(n20450), .B(n20449), .Z(n20459) );
  XOR U25090 ( .A(n20452), .B(n20451), .Z(n20449) );
  XOR U25091 ( .A(y[1070]), .B(x[1070]), .Z(n20451) );
  XOR U25092 ( .A(y[1069]), .B(x[1069]), .Z(n20452) );
  XOR U25093 ( .A(y[1068]), .B(x[1068]), .Z(n20450) );
  XNOR U25094 ( .A(n20443), .B(n20442), .Z(n20445) );
  XNOR U25095 ( .A(n20439), .B(n20438), .Z(n20442) );
  XOR U25096 ( .A(n20441), .B(n20440), .Z(n20438) );
  XOR U25097 ( .A(y[1067]), .B(x[1067]), .Z(n20440) );
  XOR U25098 ( .A(y[1066]), .B(x[1066]), .Z(n20441) );
  XOR U25099 ( .A(y[1065]), .B(x[1065]), .Z(n20439) );
  XOR U25100 ( .A(n20433), .B(n20432), .Z(n20443) );
  XOR U25101 ( .A(n20435), .B(n20434), .Z(n20432) );
  XOR U25102 ( .A(y[1064]), .B(x[1064]), .Z(n20434) );
  XOR U25103 ( .A(y[1063]), .B(x[1063]), .Z(n20435) );
  XOR U25104 ( .A(y[1062]), .B(x[1062]), .Z(n20433) );
  NAND U25105 ( .A(n20496), .B(n20497), .Z(N28461) );
  NAND U25106 ( .A(n20498), .B(n20499), .Z(n20497) );
  NANDN U25107 ( .A(n20500), .B(n20501), .Z(n20499) );
  NANDN U25108 ( .A(n20501), .B(n20500), .Z(n20496) );
  XOR U25109 ( .A(n20500), .B(n20502), .Z(N28460) );
  XNOR U25110 ( .A(n20498), .B(n20501), .Z(n20502) );
  NAND U25111 ( .A(n20503), .B(n20504), .Z(n20501) );
  NAND U25112 ( .A(n20505), .B(n20506), .Z(n20504) );
  NANDN U25113 ( .A(n20507), .B(n20508), .Z(n20506) );
  NANDN U25114 ( .A(n20508), .B(n20507), .Z(n20503) );
  AND U25115 ( .A(n20509), .B(n20510), .Z(n20498) );
  NAND U25116 ( .A(n20511), .B(n20512), .Z(n20510) );
  OR U25117 ( .A(n20513), .B(n20514), .Z(n20512) );
  NAND U25118 ( .A(n20514), .B(n20513), .Z(n20509) );
  IV U25119 ( .A(n20515), .Z(n20514) );
  AND U25120 ( .A(n20516), .B(n20517), .Z(n20500) );
  NAND U25121 ( .A(n20518), .B(n20519), .Z(n20517) );
  NANDN U25122 ( .A(n20520), .B(n20521), .Z(n20519) );
  NANDN U25123 ( .A(n20521), .B(n20520), .Z(n20516) );
  XOR U25124 ( .A(n20513), .B(n20522), .Z(N28459) );
  XOR U25125 ( .A(n20511), .B(n20515), .Z(n20522) );
  XNOR U25126 ( .A(n20508), .B(n20523), .Z(n20515) );
  XNOR U25127 ( .A(n20505), .B(n20507), .Z(n20523) );
  AND U25128 ( .A(n20524), .B(n20525), .Z(n20507) );
  NANDN U25129 ( .A(n20526), .B(n20527), .Z(n20525) );
  NANDN U25130 ( .A(n20528), .B(n20529), .Z(n20527) );
  IV U25131 ( .A(n20530), .Z(n20529) );
  NAND U25132 ( .A(n20530), .B(n20528), .Z(n20524) );
  AND U25133 ( .A(n20531), .B(n20532), .Z(n20505) );
  NAND U25134 ( .A(n20533), .B(n20534), .Z(n20532) );
  OR U25135 ( .A(n20535), .B(n20536), .Z(n20534) );
  NAND U25136 ( .A(n20536), .B(n20535), .Z(n20531) );
  IV U25137 ( .A(n20537), .Z(n20536) );
  NAND U25138 ( .A(n20538), .B(n20539), .Z(n20508) );
  NANDN U25139 ( .A(n20540), .B(n20541), .Z(n20539) );
  NAND U25140 ( .A(n20542), .B(n20543), .Z(n20541) );
  OR U25141 ( .A(n20543), .B(n20542), .Z(n20538) );
  IV U25142 ( .A(n20544), .Z(n20542) );
  AND U25143 ( .A(n20545), .B(n20546), .Z(n20511) );
  NAND U25144 ( .A(n20547), .B(n20548), .Z(n20546) );
  NANDN U25145 ( .A(n20549), .B(n20550), .Z(n20548) );
  NANDN U25146 ( .A(n20550), .B(n20549), .Z(n20545) );
  XOR U25147 ( .A(n20521), .B(n20551), .Z(n20513) );
  XNOR U25148 ( .A(n20518), .B(n20520), .Z(n20551) );
  AND U25149 ( .A(n20552), .B(n20553), .Z(n20520) );
  NANDN U25150 ( .A(n20554), .B(n20555), .Z(n20553) );
  NANDN U25151 ( .A(n20556), .B(n20557), .Z(n20555) );
  IV U25152 ( .A(n20558), .Z(n20557) );
  NAND U25153 ( .A(n20558), .B(n20556), .Z(n20552) );
  AND U25154 ( .A(n20559), .B(n20560), .Z(n20518) );
  NAND U25155 ( .A(n20561), .B(n20562), .Z(n20560) );
  OR U25156 ( .A(n20563), .B(n20564), .Z(n20562) );
  NAND U25157 ( .A(n20564), .B(n20563), .Z(n20559) );
  IV U25158 ( .A(n20565), .Z(n20564) );
  NAND U25159 ( .A(n20566), .B(n20567), .Z(n20521) );
  NANDN U25160 ( .A(n20568), .B(n20569), .Z(n20567) );
  NAND U25161 ( .A(n20570), .B(n20571), .Z(n20569) );
  OR U25162 ( .A(n20571), .B(n20570), .Z(n20566) );
  IV U25163 ( .A(n20572), .Z(n20570) );
  XOR U25164 ( .A(n20547), .B(n20573), .Z(N28458) );
  XNOR U25165 ( .A(n20550), .B(n20549), .Z(n20573) );
  XNOR U25166 ( .A(n20561), .B(n20574), .Z(n20549) );
  XOR U25167 ( .A(n20565), .B(n20563), .Z(n20574) );
  XOR U25168 ( .A(n20571), .B(n20575), .Z(n20563) );
  XOR U25169 ( .A(n20568), .B(n20572), .Z(n20575) );
  NAND U25170 ( .A(n20576), .B(n20577), .Z(n20572) );
  NAND U25171 ( .A(n20578), .B(n20579), .Z(n20577) );
  NAND U25172 ( .A(n20580), .B(n20581), .Z(n20576) );
  AND U25173 ( .A(n20582), .B(n20583), .Z(n20568) );
  NAND U25174 ( .A(n20584), .B(n20585), .Z(n20583) );
  NAND U25175 ( .A(n20586), .B(n20587), .Z(n20582) );
  NANDN U25176 ( .A(n20588), .B(n20589), .Z(n20571) );
  NANDN U25177 ( .A(n20590), .B(n20591), .Z(n20565) );
  XNOR U25178 ( .A(n20556), .B(n20592), .Z(n20561) );
  XOR U25179 ( .A(n20554), .B(n20558), .Z(n20592) );
  NAND U25180 ( .A(n20593), .B(n20594), .Z(n20558) );
  NAND U25181 ( .A(n20595), .B(n20596), .Z(n20594) );
  NAND U25182 ( .A(n20597), .B(n20598), .Z(n20593) );
  AND U25183 ( .A(n20599), .B(n20600), .Z(n20554) );
  NAND U25184 ( .A(n20601), .B(n20602), .Z(n20600) );
  NAND U25185 ( .A(n20603), .B(n20604), .Z(n20599) );
  AND U25186 ( .A(n20605), .B(n20606), .Z(n20556) );
  NAND U25187 ( .A(n20607), .B(n20608), .Z(n20550) );
  XNOR U25188 ( .A(n20533), .B(n20609), .Z(n20547) );
  XOR U25189 ( .A(n20537), .B(n20535), .Z(n20609) );
  XOR U25190 ( .A(n20543), .B(n20610), .Z(n20535) );
  XOR U25191 ( .A(n20540), .B(n20544), .Z(n20610) );
  NAND U25192 ( .A(n20611), .B(n20612), .Z(n20544) );
  NAND U25193 ( .A(n20613), .B(n20614), .Z(n20612) );
  NAND U25194 ( .A(n20615), .B(n20616), .Z(n20611) );
  AND U25195 ( .A(n20617), .B(n20618), .Z(n20540) );
  NAND U25196 ( .A(n20619), .B(n20620), .Z(n20618) );
  NAND U25197 ( .A(n20621), .B(n20622), .Z(n20617) );
  NANDN U25198 ( .A(n20623), .B(n20624), .Z(n20543) );
  NANDN U25199 ( .A(n20625), .B(n20626), .Z(n20537) );
  XNOR U25200 ( .A(n20528), .B(n20627), .Z(n20533) );
  XOR U25201 ( .A(n20526), .B(n20530), .Z(n20627) );
  NAND U25202 ( .A(n20628), .B(n20629), .Z(n20530) );
  NAND U25203 ( .A(n20630), .B(n20631), .Z(n20629) );
  NAND U25204 ( .A(n20632), .B(n20633), .Z(n20628) );
  AND U25205 ( .A(n20634), .B(n20635), .Z(n20526) );
  NAND U25206 ( .A(n20636), .B(n20637), .Z(n20635) );
  NAND U25207 ( .A(n20638), .B(n20639), .Z(n20634) );
  AND U25208 ( .A(n20640), .B(n20641), .Z(n20528) );
  XOR U25209 ( .A(n20608), .B(n20607), .Z(N28457) );
  XNOR U25210 ( .A(n20626), .B(n20625), .Z(n20607) );
  XNOR U25211 ( .A(n20640), .B(n20641), .Z(n20625) );
  XOR U25212 ( .A(n20637), .B(n20636), .Z(n20641) );
  XOR U25213 ( .A(y[1059]), .B(x[1059]), .Z(n20636) );
  XOR U25214 ( .A(n20639), .B(n20638), .Z(n20637) );
  XOR U25215 ( .A(y[1061]), .B(x[1061]), .Z(n20638) );
  XOR U25216 ( .A(y[1060]), .B(x[1060]), .Z(n20639) );
  XOR U25217 ( .A(n20631), .B(n20630), .Z(n20640) );
  XOR U25218 ( .A(n20633), .B(n20632), .Z(n20630) );
  XOR U25219 ( .A(y[1058]), .B(x[1058]), .Z(n20632) );
  XOR U25220 ( .A(y[1057]), .B(x[1057]), .Z(n20633) );
  XOR U25221 ( .A(y[1056]), .B(x[1056]), .Z(n20631) );
  XNOR U25222 ( .A(n20624), .B(n20623), .Z(n20626) );
  XNOR U25223 ( .A(n20620), .B(n20619), .Z(n20623) );
  XOR U25224 ( .A(n20622), .B(n20621), .Z(n20619) );
  XOR U25225 ( .A(y[1055]), .B(x[1055]), .Z(n20621) );
  XOR U25226 ( .A(y[1054]), .B(x[1054]), .Z(n20622) );
  XOR U25227 ( .A(y[1053]), .B(x[1053]), .Z(n20620) );
  XOR U25228 ( .A(n20614), .B(n20613), .Z(n20624) );
  XOR U25229 ( .A(n20616), .B(n20615), .Z(n20613) );
  XOR U25230 ( .A(y[1052]), .B(x[1052]), .Z(n20615) );
  XOR U25231 ( .A(y[1051]), .B(x[1051]), .Z(n20616) );
  XOR U25232 ( .A(y[1050]), .B(x[1050]), .Z(n20614) );
  XNOR U25233 ( .A(n20591), .B(n20590), .Z(n20608) );
  XNOR U25234 ( .A(n20605), .B(n20606), .Z(n20590) );
  XOR U25235 ( .A(n20602), .B(n20601), .Z(n20606) );
  XOR U25236 ( .A(y[1047]), .B(x[1047]), .Z(n20601) );
  XOR U25237 ( .A(n20604), .B(n20603), .Z(n20602) );
  XOR U25238 ( .A(y[1049]), .B(x[1049]), .Z(n20603) );
  XOR U25239 ( .A(y[1048]), .B(x[1048]), .Z(n20604) );
  XOR U25240 ( .A(n20596), .B(n20595), .Z(n20605) );
  XOR U25241 ( .A(n20598), .B(n20597), .Z(n20595) );
  XOR U25242 ( .A(y[1046]), .B(x[1046]), .Z(n20597) );
  XOR U25243 ( .A(y[1045]), .B(x[1045]), .Z(n20598) );
  XOR U25244 ( .A(y[1044]), .B(x[1044]), .Z(n20596) );
  XNOR U25245 ( .A(n20589), .B(n20588), .Z(n20591) );
  XNOR U25246 ( .A(n20585), .B(n20584), .Z(n20588) );
  XOR U25247 ( .A(n20587), .B(n20586), .Z(n20584) );
  XOR U25248 ( .A(y[1043]), .B(x[1043]), .Z(n20586) );
  XOR U25249 ( .A(y[1042]), .B(x[1042]), .Z(n20587) );
  XOR U25250 ( .A(y[1041]), .B(x[1041]), .Z(n20585) );
  XOR U25251 ( .A(n20579), .B(n20578), .Z(n20589) );
  XOR U25252 ( .A(n20581), .B(n20580), .Z(n20578) );
  XOR U25253 ( .A(y[1040]), .B(x[1040]), .Z(n20580) );
  XOR U25254 ( .A(y[1039]), .B(x[1039]), .Z(n20581) );
  XOR U25255 ( .A(y[1038]), .B(x[1038]), .Z(n20579) );
  NAND U25256 ( .A(n20642), .B(n20643), .Z(N28449) );
  NAND U25257 ( .A(n20644), .B(n20645), .Z(n20643) );
  NANDN U25258 ( .A(n20646), .B(n20647), .Z(n20645) );
  NANDN U25259 ( .A(n20647), .B(n20646), .Z(n20642) );
  XOR U25260 ( .A(n20646), .B(n20648), .Z(N28448) );
  XNOR U25261 ( .A(n20644), .B(n20647), .Z(n20648) );
  NAND U25262 ( .A(n20649), .B(n20650), .Z(n20647) );
  NAND U25263 ( .A(n20651), .B(n20652), .Z(n20650) );
  NANDN U25264 ( .A(n20653), .B(n20654), .Z(n20652) );
  NANDN U25265 ( .A(n20654), .B(n20653), .Z(n20649) );
  AND U25266 ( .A(n20655), .B(n20656), .Z(n20644) );
  NAND U25267 ( .A(n20657), .B(n20658), .Z(n20656) );
  OR U25268 ( .A(n20659), .B(n20660), .Z(n20658) );
  NAND U25269 ( .A(n20660), .B(n20659), .Z(n20655) );
  IV U25270 ( .A(n20661), .Z(n20660) );
  AND U25271 ( .A(n20662), .B(n20663), .Z(n20646) );
  NAND U25272 ( .A(n20664), .B(n20665), .Z(n20663) );
  NANDN U25273 ( .A(n20666), .B(n20667), .Z(n20665) );
  NANDN U25274 ( .A(n20667), .B(n20666), .Z(n20662) );
  XOR U25275 ( .A(n20659), .B(n20668), .Z(N28447) );
  XOR U25276 ( .A(n20657), .B(n20661), .Z(n20668) );
  XNOR U25277 ( .A(n20654), .B(n20669), .Z(n20661) );
  XNOR U25278 ( .A(n20651), .B(n20653), .Z(n20669) );
  AND U25279 ( .A(n20670), .B(n20671), .Z(n20653) );
  NANDN U25280 ( .A(n20672), .B(n20673), .Z(n20671) );
  NANDN U25281 ( .A(n20674), .B(n20675), .Z(n20673) );
  IV U25282 ( .A(n20676), .Z(n20675) );
  NAND U25283 ( .A(n20676), .B(n20674), .Z(n20670) );
  AND U25284 ( .A(n20677), .B(n20678), .Z(n20651) );
  NAND U25285 ( .A(n20679), .B(n20680), .Z(n20678) );
  OR U25286 ( .A(n20681), .B(n20682), .Z(n20680) );
  NAND U25287 ( .A(n20682), .B(n20681), .Z(n20677) );
  IV U25288 ( .A(n20683), .Z(n20682) );
  NAND U25289 ( .A(n20684), .B(n20685), .Z(n20654) );
  NANDN U25290 ( .A(n20686), .B(n20687), .Z(n20685) );
  NAND U25291 ( .A(n20688), .B(n20689), .Z(n20687) );
  OR U25292 ( .A(n20689), .B(n20688), .Z(n20684) );
  IV U25293 ( .A(n20690), .Z(n20688) );
  AND U25294 ( .A(n20691), .B(n20692), .Z(n20657) );
  NAND U25295 ( .A(n20693), .B(n20694), .Z(n20692) );
  NANDN U25296 ( .A(n20695), .B(n20696), .Z(n20694) );
  NANDN U25297 ( .A(n20696), .B(n20695), .Z(n20691) );
  XOR U25298 ( .A(n20667), .B(n20697), .Z(n20659) );
  XNOR U25299 ( .A(n20664), .B(n20666), .Z(n20697) );
  AND U25300 ( .A(n20698), .B(n20699), .Z(n20666) );
  NANDN U25301 ( .A(n20700), .B(n20701), .Z(n20699) );
  NANDN U25302 ( .A(n20702), .B(n20703), .Z(n20701) );
  IV U25303 ( .A(n20704), .Z(n20703) );
  NAND U25304 ( .A(n20704), .B(n20702), .Z(n20698) );
  AND U25305 ( .A(n20705), .B(n20706), .Z(n20664) );
  NAND U25306 ( .A(n20707), .B(n20708), .Z(n20706) );
  OR U25307 ( .A(n20709), .B(n20710), .Z(n20708) );
  NAND U25308 ( .A(n20710), .B(n20709), .Z(n20705) );
  IV U25309 ( .A(n20711), .Z(n20710) );
  NAND U25310 ( .A(n20712), .B(n20713), .Z(n20667) );
  NANDN U25311 ( .A(n20714), .B(n20715), .Z(n20713) );
  NAND U25312 ( .A(n20716), .B(n20717), .Z(n20715) );
  OR U25313 ( .A(n20717), .B(n20716), .Z(n20712) );
  IV U25314 ( .A(n20718), .Z(n20716) );
  XOR U25315 ( .A(n20693), .B(n20719), .Z(N28446) );
  XNOR U25316 ( .A(n20696), .B(n20695), .Z(n20719) );
  XNOR U25317 ( .A(n20707), .B(n20720), .Z(n20695) );
  XOR U25318 ( .A(n20711), .B(n20709), .Z(n20720) );
  XOR U25319 ( .A(n20717), .B(n20721), .Z(n20709) );
  XOR U25320 ( .A(n20714), .B(n20718), .Z(n20721) );
  NAND U25321 ( .A(n20722), .B(n20723), .Z(n20718) );
  NAND U25322 ( .A(n20724), .B(n20725), .Z(n20723) );
  NAND U25323 ( .A(n20726), .B(n20727), .Z(n20722) );
  AND U25324 ( .A(n20728), .B(n20729), .Z(n20714) );
  NAND U25325 ( .A(n20730), .B(n20731), .Z(n20729) );
  NAND U25326 ( .A(n20732), .B(n20733), .Z(n20728) );
  NANDN U25327 ( .A(n20734), .B(n20735), .Z(n20717) );
  NANDN U25328 ( .A(n20736), .B(n20737), .Z(n20711) );
  XNOR U25329 ( .A(n20702), .B(n20738), .Z(n20707) );
  XOR U25330 ( .A(n20700), .B(n20704), .Z(n20738) );
  NAND U25331 ( .A(n20739), .B(n20740), .Z(n20704) );
  NAND U25332 ( .A(n20741), .B(n20742), .Z(n20740) );
  NAND U25333 ( .A(n20743), .B(n20744), .Z(n20739) );
  AND U25334 ( .A(n20745), .B(n20746), .Z(n20700) );
  NAND U25335 ( .A(n20747), .B(n20748), .Z(n20746) );
  NAND U25336 ( .A(n20749), .B(n20750), .Z(n20745) );
  AND U25337 ( .A(n20751), .B(n20752), .Z(n20702) );
  NAND U25338 ( .A(n20753), .B(n20754), .Z(n20696) );
  XNOR U25339 ( .A(n20679), .B(n20755), .Z(n20693) );
  XOR U25340 ( .A(n20683), .B(n20681), .Z(n20755) );
  XOR U25341 ( .A(n20689), .B(n20756), .Z(n20681) );
  XOR U25342 ( .A(n20686), .B(n20690), .Z(n20756) );
  NAND U25343 ( .A(n20757), .B(n20758), .Z(n20690) );
  NAND U25344 ( .A(n20759), .B(n20760), .Z(n20758) );
  NAND U25345 ( .A(n20761), .B(n20762), .Z(n20757) );
  AND U25346 ( .A(n20763), .B(n20764), .Z(n20686) );
  NAND U25347 ( .A(n20765), .B(n20766), .Z(n20764) );
  NAND U25348 ( .A(n20767), .B(n20768), .Z(n20763) );
  NANDN U25349 ( .A(n20769), .B(n20770), .Z(n20689) );
  NANDN U25350 ( .A(n20771), .B(n20772), .Z(n20683) );
  XNOR U25351 ( .A(n20674), .B(n20773), .Z(n20679) );
  XOR U25352 ( .A(n20672), .B(n20676), .Z(n20773) );
  NAND U25353 ( .A(n20774), .B(n20775), .Z(n20676) );
  NAND U25354 ( .A(n20776), .B(n20777), .Z(n20775) );
  NAND U25355 ( .A(n20778), .B(n20779), .Z(n20774) );
  AND U25356 ( .A(n20780), .B(n20781), .Z(n20672) );
  NAND U25357 ( .A(n20782), .B(n20783), .Z(n20781) );
  NAND U25358 ( .A(n20784), .B(n20785), .Z(n20780) );
  AND U25359 ( .A(n20786), .B(n20787), .Z(n20674) );
  XOR U25360 ( .A(n20754), .B(n20753), .Z(N28445) );
  XNOR U25361 ( .A(n20772), .B(n20771), .Z(n20753) );
  XNOR U25362 ( .A(n20786), .B(n20787), .Z(n20771) );
  XOR U25363 ( .A(n20783), .B(n20782), .Z(n20787) );
  XOR U25364 ( .A(y[1035]), .B(x[1035]), .Z(n20782) );
  XOR U25365 ( .A(n20785), .B(n20784), .Z(n20783) );
  XOR U25366 ( .A(y[1037]), .B(x[1037]), .Z(n20784) );
  XOR U25367 ( .A(y[1036]), .B(x[1036]), .Z(n20785) );
  XOR U25368 ( .A(n20777), .B(n20776), .Z(n20786) );
  XOR U25369 ( .A(n20779), .B(n20778), .Z(n20776) );
  XOR U25370 ( .A(y[1034]), .B(x[1034]), .Z(n20778) );
  XOR U25371 ( .A(y[1033]), .B(x[1033]), .Z(n20779) );
  XOR U25372 ( .A(y[1032]), .B(x[1032]), .Z(n20777) );
  XNOR U25373 ( .A(n20770), .B(n20769), .Z(n20772) );
  XNOR U25374 ( .A(n20766), .B(n20765), .Z(n20769) );
  XOR U25375 ( .A(n20768), .B(n20767), .Z(n20765) );
  XOR U25376 ( .A(y[1031]), .B(x[1031]), .Z(n20767) );
  XOR U25377 ( .A(y[1030]), .B(x[1030]), .Z(n20768) );
  XOR U25378 ( .A(y[1029]), .B(x[1029]), .Z(n20766) );
  XOR U25379 ( .A(n20760), .B(n20759), .Z(n20770) );
  XOR U25380 ( .A(n20762), .B(n20761), .Z(n20759) );
  XOR U25381 ( .A(y[1028]), .B(x[1028]), .Z(n20761) );
  XOR U25382 ( .A(y[1027]), .B(x[1027]), .Z(n20762) );
  XOR U25383 ( .A(y[1026]), .B(x[1026]), .Z(n20760) );
  XNOR U25384 ( .A(n20737), .B(n20736), .Z(n20754) );
  XNOR U25385 ( .A(n20751), .B(n20752), .Z(n20736) );
  XOR U25386 ( .A(n20748), .B(n20747), .Z(n20752) );
  XOR U25387 ( .A(y[1023]), .B(x[1023]), .Z(n20747) );
  XOR U25388 ( .A(n20750), .B(n20749), .Z(n20748) );
  XOR U25389 ( .A(y[1025]), .B(x[1025]), .Z(n20749) );
  XOR U25390 ( .A(y[1024]), .B(x[1024]), .Z(n20750) );
  XOR U25391 ( .A(n20742), .B(n20741), .Z(n20751) );
  XOR U25392 ( .A(n20744), .B(n20743), .Z(n20741) );
  XOR U25393 ( .A(y[1022]), .B(x[1022]), .Z(n20743) );
  XOR U25394 ( .A(y[1021]), .B(x[1021]), .Z(n20744) );
  XOR U25395 ( .A(y[1020]), .B(x[1020]), .Z(n20742) );
  XNOR U25396 ( .A(n20735), .B(n20734), .Z(n20737) );
  XNOR U25397 ( .A(n20731), .B(n20730), .Z(n20734) );
  XOR U25398 ( .A(n20733), .B(n20732), .Z(n20730) );
  XOR U25399 ( .A(y[1019]), .B(x[1019]), .Z(n20732) );
  XOR U25400 ( .A(y[1018]), .B(x[1018]), .Z(n20733) );
  XOR U25401 ( .A(y[1017]), .B(x[1017]), .Z(n20731) );
  XOR U25402 ( .A(n20725), .B(n20724), .Z(n20735) );
  XOR U25403 ( .A(n20727), .B(n20726), .Z(n20724) );
  XOR U25404 ( .A(y[1016]), .B(x[1016]), .Z(n20726) );
  XOR U25405 ( .A(y[1015]), .B(x[1015]), .Z(n20727) );
  XOR U25406 ( .A(y[1014]), .B(x[1014]), .Z(n20725) );
  NAND U25407 ( .A(n20788), .B(n20789), .Z(N28437) );
  NAND U25408 ( .A(n20790), .B(n20791), .Z(n20789) );
  NANDN U25409 ( .A(n20792), .B(n20793), .Z(n20791) );
  NANDN U25410 ( .A(n20793), .B(n20792), .Z(n20788) );
  XOR U25411 ( .A(n20792), .B(n20794), .Z(N28436) );
  XNOR U25412 ( .A(n20790), .B(n20793), .Z(n20794) );
  NAND U25413 ( .A(n20795), .B(n20796), .Z(n20793) );
  NAND U25414 ( .A(n20797), .B(n20798), .Z(n20796) );
  NANDN U25415 ( .A(n20799), .B(n20800), .Z(n20798) );
  NANDN U25416 ( .A(n20800), .B(n20799), .Z(n20795) );
  AND U25417 ( .A(n20801), .B(n20802), .Z(n20790) );
  NAND U25418 ( .A(n20803), .B(n20804), .Z(n20802) );
  OR U25419 ( .A(n20805), .B(n20806), .Z(n20804) );
  NAND U25420 ( .A(n20806), .B(n20805), .Z(n20801) );
  IV U25421 ( .A(n20807), .Z(n20806) );
  AND U25422 ( .A(n20808), .B(n20809), .Z(n20792) );
  NAND U25423 ( .A(n20810), .B(n20811), .Z(n20809) );
  NANDN U25424 ( .A(n20812), .B(n20813), .Z(n20811) );
  NANDN U25425 ( .A(n20813), .B(n20812), .Z(n20808) );
  XOR U25426 ( .A(n20805), .B(n20814), .Z(N28435) );
  XOR U25427 ( .A(n20803), .B(n20807), .Z(n20814) );
  XNOR U25428 ( .A(n20800), .B(n20815), .Z(n20807) );
  XNOR U25429 ( .A(n20797), .B(n20799), .Z(n20815) );
  AND U25430 ( .A(n20816), .B(n20817), .Z(n20799) );
  NANDN U25431 ( .A(n20818), .B(n20819), .Z(n20817) );
  NANDN U25432 ( .A(n20820), .B(n20821), .Z(n20819) );
  IV U25433 ( .A(n20822), .Z(n20821) );
  NAND U25434 ( .A(n20822), .B(n20820), .Z(n20816) );
  AND U25435 ( .A(n20823), .B(n20824), .Z(n20797) );
  NAND U25436 ( .A(n20825), .B(n20826), .Z(n20824) );
  OR U25437 ( .A(n20827), .B(n20828), .Z(n20826) );
  NAND U25438 ( .A(n20828), .B(n20827), .Z(n20823) );
  IV U25439 ( .A(n20829), .Z(n20828) );
  NAND U25440 ( .A(n20830), .B(n20831), .Z(n20800) );
  NANDN U25441 ( .A(n20832), .B(n20833), .Z(n20831) );
  NAND U25442 ( .A(n20834), .B(n20835), .Z(n20833) );
  OR U25443 ( .A(n20835), .B(n20834), .Z(n20830) );
  IV U25444 ( .A(n20836), .Z(n20834) );
  AND U25445 ( .A(n20837), .B(n20838), .Z(n20803) );
  NAND U25446 ( .A(n20839), .B(n20840), .Z(n20838) );
  NANDN U25447 ( .A(n20841), .B(n20842), .Z(n20840) );
  NANDN U25448 ( .A(n20842), .B(n20841), .Z(n20837) );
  XOR U25449 ( .A(n20813), .B(n20843), .Z(n20805) );
  XNOR U25450 ( .A(n20810), .B(n20812), .Z(n20843) );
  AND U25451 ( .A(n20844), .B(n20845), .Z(n20812) );
  NANDN U25452 ( .A(n20846), .B(n20847), .Z(n20845) );
  NANDN U25453 ( .A(n20848), .B(n20849), .Z(n20847) );
  IV U25454 ( .A(n20850), .Z(n20849) );
  NAND U25455 ( .A(n20850), .B(n20848), .Z(n20844) );
  AND U25456 ( .A(n20851), .B(n20852), .Z(n20810) );
  NAND U25457 ( .A(n20853), .B(n20854), .Z(n20852) );
  OR U25458 ( .A(n20855), .B(n20856), .Z(n20854) );
  NAND U25459 ( .A(n20856), .B(n20855), .Z(n20851) );
  IV U25460 ( .A(n20857), .Z(n20856) );
  NAND U25461 ( .A(n20858), .B(n20859), .Z(n20813) );
  NANDN U25462 ( .A(n20860), .B(n20861), .Z(n20859) );
  NAND U25463 ( .A(n20862), .B(n20863), .Z(n20861) );
  OR U25464 ( .A(n20863), .B(n20862), .Z(n20858) );
  IV U25465 ( .A(n20864), .Z(n20862) );
  XOR U25466 ( .A(n20839), .B(n20865), .Z(N28434) );
  XNOR U25467 ( .A(n20842), .B(n20841), .Z(n20865) );
  XNOR U25468 ( .A(n20853), .B(n20866), .Z(n20841) );
  XOR U25469 ( .A(n20857), .B(n20855), .Z(n20866) );
  XOR U25470 ( .A(n20863), .B(n20867), .Z(n20855) );
  XOR U25471 ( .A(n20860), .B(n20864), .Z(n20867) );
  NAND U25472 ( .A(n20868), .B(n20869), .Z(n20864) );
  NAND U25473 ( .A(n20870), .B(n20871), .Z(n20869) );
  NAND U25474 ( .A(n20872), .B(n20873), .Z(n20868) );
  AND U25475 ( .A(n20874), .B(n20875), .Z(n20860) );
  NAND U25476 ( .A(n20876), .B(n20877), .Z(n20875) );
  NAND U25477 ( .A(n20878), .B(n20879), .Z(n20874) );
  NANDN U25478 ( .A(n20880), .B(n20881), .Z(n20863) );
  NANDN U25479 ( .A(n20882), .B(n20883), .Z(n20857) );
  XNOR U25480 ( .A(n20848), .B(n20884), .Z(n20853) );
  XOR U25481 ( .A(n20846), .B(n20850), .Z(n20884) );
  NAND U25482 ( .A(n20885), .B(n20886), .Z(n20850) );
  NAND U25483 ( .A(n20887), .B(n20888), .Z(n20886) );
  NAND U25484 ( .A(n20889), .B(n20890), .Z(n20885) );
  AND U25485 ( .A(n20891), .B(n20892), .Z(n20846) );
  NAND U25486 ( .A(n20893), .B(n20894), .Z(n20892) );
  NAND U25487 ( .A(n20895), .B(n20896), .Z(n20891) );
  AND U25488 ( .A(n20897), .B(n20898), .Z(n20848) );
  NAND U25489 ( .A(n20899), .B(n20900), .Z(n20842) );
  XNOR U25490 ( .A(n20825), .B(n20901), .Z(n20839) );
  XOR U25491 ( .A(n20829), .B(n20827), .Z(n20901) );
  XOR U25492 ( .A(n20835), .B(n20902), .Z(n20827) );
  XOR U25493 ( .A(n20832), .B(n20836), .Z(n20902) );
  NAND U25494 ( .A(n20903), .B(n20904), .Z(n20836) );
  NAND U25495 ( .A(n20905), .B(n20906), .Z(n20904) );
  NAND U25496 ( .A(n20907), .B(n20908), .Z(n20903) );
  AND U25497 ( .A(n20909), .B(n20910), .Z(n20832) );
  NAND U25498 ( .A(n20911), .B(n20912), .Z(n20910) );
  NAND U25499 ( .A(n20913), .B(n20914), .Z(n20909) );
  NANDN U25500 ( .A(n20915), .B(n20916), .Z(n20835) );
  NANDN U25501 ( .A(n20917), .B(n20918), .Z(n20829) );
  XNOR U25502 ( .A(n20820), .B(n20919), .Z(n20825) );
  XOR U25503 ( .A(n20818), .B(n20822), .Z(n20919) );
  NAND U25504 ( .A(n20920), .B(n20921), .Z(n20822) );
  NAND U25505 ( .A(n20922), .B(n20923), .Z(n20921) );
  NAND U25506 ( .A(n20924), .B(n20925), .Z(n20920) );
  AND U25507 ( .A(n20926), .B(n20927), .Z(n20818) );
  NAND U25508 ( .A(n20928), .B(n20929), .Z(n20927) );
  NAND U25509 ( .A(n20930), .B(n20931), .Z(n20926) );
  AND U25510 ( .A(n20932), .B(n20933), .Z(n20820) );
  XOR U25511 ( .A(n20900), .B(n20899), .Z(N28433) );
  XNOR U25512 ( .A(n20918), .B(n20917), .Z(n20899) );
  XNOR U25513 ( .A(n20932), .B(n20933), .Z(n20917) );
  XOR U25514 ( .A(n20929), .B(n20928), .Z(n20933) );
  XOR U25515 ( .A(y[1011]), .B(x[1011]), .Z(n20928) );
  XOR U25516 ( .A(n20931), .B(n20930), .Z(n20929) );
  XOR U25517 ( .A(y[1013]), .B(x[1013]), .Z(n20930) );
  XOR U25518 ( .A(y[1012]), .B(x[1012]), .Z(n20931) );
  XOR U25519 ( .A(n20923), .B(n20922), .Z(n20932) );
  XOR U25520 ( .A(n20925), .B(n20924), .Z(n20922) );
  XOR U25521 ( .A(y[1010]), .B(x[1010]), .Z(n20924) );
  XOR U25522 ( .A(y[1009]), .B(x[1009]), .Z(n20925) );
  XOR U25523 ( .A(y[1008]), .B(x[1008]), .Z(n20923) );
  XNOR U25524 ( .A(n20916), .B(n20915), .Z(n20918) );
  XNOR U25525 ( .A(n20912), .B(n20911), .Z(n20915) );
  XOR U25526 ( .A(n20914), .B(n20913), .Z(n20911) );
  XOR U25527 ( .A(y[1007]), .B(x[1007]), .Z(n20913) );
  XOR U25528 ( .A(y[1006]), .B(x[1006]), .Z(n20914) );
  XOR U25529 ( .A(y[1005]), .B(x[1005]), .Z(n20912) );
  XOR U25530 ( .A(n20906), .B(n20905), .Z(n20916) );
  XOR U25531 ( .A(n20908), .B(n20907), .Z(n20905) );
  XOR U25532 ( .A(y[1004]), .B(x[1004]), .Z(n20907) );
  XOR U25533 ( .A(y[1003]), .B(x[1003]), .Z(n20908) );
  XOR U25534 ( .A(y[1002]), .B(x[1002]), .Z(n20906) );
  XNOR U25535 ( .A(n20883), .B(n20882), .Z(n20900) );
  XNOR U25536 ( .A(n20897), .B(n20898), .Z(n20882) );
  XOR U25537 ( .A(n20894), .B(n20893), .Z(n20898) );
  XOR U25538 ( .A(y[999]), .B(x[999]), .Z(n20893) );
  XOR U25539 ( .A(n20896), .B(n20895), .Z(n20894) );
  XOR U25540 ( .A(y[1001]), .B(x[1001]), .Z(n20895) );
  XOR U25541 ( .A(y[1000]), .B(x[1000]), .Z(n20896) );
  XOR U25542 ( .A(n20888), .B(n20887), .Z(n20897) );
  XOR U25543 ( .A(n20890), .B(n20889), .Z(n20887) );
  XOR U25544 ( .A(y[998]), .B(x[998]), .Z(n20889) );
  XOR U25545 ( .A(y[997]), .B(x[997]), .Z(n20890) );
  XOR U25546 ( .A(y[996]), .B(x[996]), .Z(n20888) );
  XNOR U25547 ( .A(n20881), .B(n20880), .Z(n20883) );
  XNOR U25548 ( .A(n20877), .B(n20876), .Z(n20880) );
  XOR U25549 ( .A(n20879), .B(n20878), .Z(n20876) );
  XOR U25550 ( .A(y[995]), .B(x[995]), .Z(n20878) );
  XOR U25551 ( .A(y[994]), .B(x[994]), .Z(n20879) );
  XOR U25552 ( .A(y[993]), .B(x[993]), .Z(n20877) );
  XOR U25553 ( .A(n20871), .B(n20870), .Z(n20881) );
  XOR U25554 ( .A(n20873), .B(n20872), .Z(n20870) );
  XOR U25555 ( .A(y[992]), .B(x[992]), .Z(n20872) );
  XOR U25556 ( .A(y[991]), .B(x[991]), .Z(n20873) );
  XOR U25557 ( .A(y[990]), .B(x[990]), .Z(n20871) );
  NAND U25558 ( .A(n20934), .B(n20935), .Z(N28425) );
  NAND U25559 ( .A(n20936), .B(n20937), .Z(n20935) );
  NANDN U25560 ( .A(n20938), .B(n20939), .Z(n20937) );
  NANDN U25561 ( .A(n20939), .B(n20938), .Z(n20934) );
  XOR U25562 ( .A(n20938), .B(n20940), .Z(N28424) );
  XNOR U25563 ( .A(n20936), .B(n20939), .Z(n20940) );
  NAND U25564 ( .A(n20941), .B(n20942), .Z(n20939) );
  NAND U25565 ( .A(n20943), .B(n20944), .Z(n20942) );
  NANDN U25566 ( .A(n20945), .B(n20946), .Z(n20944) );
  NANDN U25567 ( .A(n20946), .B(n20945), .Z(n20941) );
  AND U25568 ( .A(n20947), .B(n20948), .Z(n20936) );
  NAND U25569 ( .A(n20949), .B(n20950), .Z(n20948) );
  OR U25570 ( .A(n20951), .B(n20952), .Z(n20950) );
  NAND U25571 ( .A(n20952), .B(n20951), .Z(n20947) );
  IV U25572 ( .A(n20953), .Z(n20952) );
  AND U25573 ( .A(n20954), .B(n20955), .Z(n20938) );
  NAND U25574 ( .A(n20956), .B(n20957), .Z(n20955) );
  NANDN U25575 ( .A(n20958), .B(n20959), .Z(n20957) );
  NANDN U25576 ( .A(n20959), .B(n20958), .Z(n20954) );
  XOR U25577 ( .A(n20951), .B(n20960), .Z(N28423) );
  XOR U25578 ( .A(n20949), .B(n20953), .Z(n20960) );
  XNOR U25579 ( .A(n20946), .B(n20961), .Z(n20953) );
  XNOR U25580 ( .A(n20943), .B(n20945), .Z(n20961) );
  AND U25581 ( .A(n20962), .B(n20963), .Z(n20945) );
  NANDN U25582 ( .A(n20964), .B(n20965), .Z(n20963) );
  NANDN U25583 ( .A(n20966), .B(n20967), .Z(n20965) );
  IV U25584 ( .A(n20968), .Z(n20967) );
  NAND U25585 ( .A(n20968), .B(n20966), .Z(n20962) );
  AND U25586 ( .A(n20969), .B(n20970), .Z(n20943) );
  NAND U25587 ( .A(n20971), .B(n20972), .Z(n20970) );
  OR U25588 ( .A(n20973), .B(n20974), .Z(n20972) );
  NAND U25589 ( .A(n20974), .B(n20973), .Z(n20969) );
  IV U25590 ( .A(n20975), .Z(n20974) );
  NAND U25591 ( .A(n20976), .B(n20977), .Z(n20946) );
  NANDN U25592 ( .A(n20978), .B(n20979), .Z(n20977) );
  NAND U25593 ( .A(n20980), .B(n20981), .Z(n20979) );
  OR U25594 ( .A(n20981), .B(n20980), .Z(n20976) );
  IV U25595 ( .A(n20982), .Z(n20980) );
  AND U25596 ( .A(n20983), .B(n20984), .Z(n20949) );
  NAND U25597 ( .A(n20985), .B(n20986), .Z(n20984) );
  NANDN U25598 ( .A(n20987), .B(n20988), .Z(n20986) );
  NANDN U25599 ( .A(n20988), .B(n20987), .Z(n20983) );
  XOR U25600 ( .A(n20959), .B(n20989), .Z(n20951) );
  XNOR U25601 ( .A(n20956), .B(n20958), .Z(n20989) );
  AND U25602 ( .A(n20990), .B(n20991), .Z(n20958) );
  NANDN U25603 ( .A(n20992), .B(n20993), .Z(n20991) );
  NANDN U25604 ( .A(n20994), .B(n20995), .Z(n20993) );
  IV U25605 ( .A(n20996), .Z(n20995) );
  NAND U25606 ( .A(n20996), .B(n20994), .Z(n20990) );
  AND U25607 ( .A(n20997), .B(n20998), .Z(n20956) );
  NAND U25608 ( .A(n20999), .B(n21000), .Z(n20998) );
  OR U25609 ( .A(n21001), .B(n21002), .Z(n21000) );
  NAND U25610 ( .A(n21002), .B(n21001), .Z(n20997) );
  IV U25611 ( .A(n21003), .Z(n21002) );
  NAND U25612 ( .A(n21004), .B(n21005), .Z(n20959) );
  NANDN U25613 ( .A(n21006), .B(n21007), .Z(n21005) );
  NAND U25614 ( .A(n21008), .B(n21009), .Z(n21007) );
  OR U25615 ( .A(n21009), .B(n21008), .Z(n21004) );
  IV U25616 ( .A(n21010), .Z(n21008) );
  XOR U25617 ( .A(n20985), .B(n21011), .Z(N28422) );
  XNOR U25618 ( .A(n20988), .B(n20987), .Z(n21011) );
  XNOR U25619 ( .A(n20999), .B(n21012), .Z(n20987) );
  XOR U25620 ( .A(n21003), .B(n21001), .Z(n21012) );
  XOR U25621 ( .A(n21009), .B(n21013), .Z(n21001) );
  XOR U25622 ( .A(n21006), .B(n21010), .Z(n21013) );
  NAND U25623 ( .A(n21014), .B(n21015), .Z(n21010) );
  NAND U25624 ( .A(n21016), .B(n21017), .Z(n21015) );
  NAND U25625 ( .A(n21018), .B(n21019), .Z(n21014) );
  AND U25626 ( .A(n21020), .B(n21021), .Z(n21006) );
  NAND U25627 ( .A(n21022), .B(n21023), .Z(n21021) );
  NAND U25628 ( .A(n21024), .B(n21025), .Z(n21020) );
  NANDN U25629 ( .A(n21026), .B(n21027), .Z(n21009) );
  NANDN U25630 ( .A(n21028), .B(n21029), .Z(n21003) );
  XNOR U25631 ( .A(n20994), .B(n21030), .Z(n20999) );
  XOR U25632 ( .A(n20992), .B(n20996), .Z(n21030) );
  NAND U25633 ( .A(n21031), .B(n21032), .Z(n20996) );
  NAND U25634 ( .A(n21033), .B(n21034), .Z(n21032) );
  NAND U25635 ( .A(n21035), .B(n21036), .Z(n21031) );
  AND U25636 ( .A(n21037), .B(n21038), .Z(n20992) );
  NAND U25637 ( .A(n21039), .B(n21040), .Z(n21038) );
  NAND U25638 ( .A(n21041), .B(n21042), .Z(n21037) );
  AND U25639 ( .A(n21043), .B(n21044), .Z(n20994) );
  NAND U25640 ( .A(n21045), .B(n21046), .Z(n20988) );
  XNOR U25641 ( .A(n20971), .B(n21047), .Z(n20985) );
  XOR U25642 ( .A(n20975), .B(n20973), .Z(n21047) );
  XOR U25643 ( .A(n20981), .B(n21048), .Z(n20973) );
  XOR U25644 ( .A(n20978), .B(n20982), .Z(n21048) );
  NAND U25645 ( .A(n21049), .B(n21050), .Z(n20982) );
  NAND U25646 ( .A(n21051), .B(n21052), .Z(n21050) );
  NAND U25647 ( .A(n21053), .B(n21054), .Z(n21049) );
  AND U25648 ( .A(n21055), .B(n21056), .Z(n20978) );
  NAND U25649 ( .A(n21057), .B(n21058), .Z(n21056) );
  NAND U25650 ( .A(n21059), .B(n21060), .Z(n21055) );
  NANDN U25651 ( .A(n21061), .B(n21062), .Z(n20981) );
  NANDN U25652 ( .A(n21063), .B(n21064), .Z(n20975) );
  XNOR U25653 ( .A(n20966), .B(n21065), .Z(n20971) );
  XOR U25654 ( .A(n20964), .B(n20968), .Z(n21065) );
  NAND U25655 ( .A(n21066), .B(n21067), .Z(n20968) );
  NAND U25656 ( .A(n21068), .B(n21069), .Z(n21067) );
  NAND U25657 ( .A(n21070), .B(n21071), .Z(n21066) );
  AND U25658 ( .A(n21072), .B(n21073), .Z(n20964) );
  NAND U25659 ( .A(n21074), .B(n21075), .Z(n21073) );
  NAND U25660 ( .A(n21076), .B(n21077), .Z(n21072) );
  AND U25661 ( .A(n21078), .B(n21079), .Z(n20966) );
  XOR U25662 ( .A(n21046), .B(n21045), .Z(N28421) );
  XNOR U25663 ( .A(n21064), .B(n21063), .Z(n21045) );
  XNOR U25664 ( .A(n21078), .B(n21079), .Z(n21063) );
  XOR U25665 ( .A(n21075), .B(n21074), .Z(n21079) );
  XOR U25666 ( .A(y[987]), .B(x[987]), .Z(n21074) );
  XOR U25667 ( .A(n21077), .B(n21076), .Z(n21075) );
  XOR U25668 ( .A(y[989]), .B(x[989]), .Z(n21076) );
  XOR U25669 ( .A(y[988]), .B(x[988]), .Z(n21077) );
  XOR U25670 ( .A(n21069), .B(n21068), .Z(n21078) );
  XOR U25671 ( .A(n21071), .B(n21070), .Z(n21068) );
  XOR U25672 ( .A(y[986]), .B(x[986]), .Z(n21070) );
  XOR U25673 ( .A(y[985]), .B(x[985]), .Z(n21071) );
  XOR U25674 ( .A(y[984]), .B(x[984]), .Z(n21069) );
  XNOR U25675 ( .A(n21062), .B(n21061), .Z(n21064) );
  XNOR U25676 ( .A(n21058), .B(n21057), .Z(n21061) );
  XOR U25677 ( .A(n21060), .B(n21059), .Z(n21057) );
  XOR U25678 ( .A(y[983]), .B(x[983]), .Z(n21059) );
  XOR U25679 ( .A(y[982]), .B(x[982]), .Z(n21060) );
  XOR U25680 ( .A(y[981]), .B(x[981]), .Z(n21058) );
  XOR U25681 ( .A(n21052), .B(n21051), .Z(n21062) );
  XOR U25682 ( .A(n21054), .B(n21053), .Z(n21051) );
  XOR U25683 ( .A(y[980]), .B(x[980]), .Z(n21053) );
  XOR U25684 ( .A(y[979]), .B(x[979]), .Z(n21054) );
  XOR U25685 ( .A(y[978]), .B(x[978]), .Z(n21052) );
  XNOR U25686 ( .A(n21029), .B(n21028), .Z(n21046) );
  XNOR U25687 ( .A(n21043), .B(n21044), .Z(n21028) );
  XOR U25688 ( .A(n21040), .B(n21039), .Z(n21044) );
  XOR U25689 ( .A(y[975]), .B(x[975]), .Z(n21039) );
  XOR U25690 ( .A(n21042), .B(n21041), .Z(n21040) );
  XOR U25691 ( .A(y[977]), .B(x[977]), .Z(n21041) );
  XOR U25692 ( .A(y[976]), .B(x[976]), .Z(n21042) );
  XOR U25693 ( .A(n21034), .B(n21033), .Z(n21043) );
  XOR U25694 ( .A(n21036), .B(n21035), .Z(n21033) );
  XOR U25695 ( .A(y[974]), .B(x[974]), .Z(n21035) );
  XOR U25696 ( .A(y[973]), .B(x[973]), .Z(n21036) );
  XOR U25697 ( .A(y[972]), .B(x[972]), .Z(n21034) );
  XNOR U25698 ( .A(n21027), .B(n21026), .Z(n21029) );
  XNOR U25699 ( .A(n21023), .B(n21022), .Z(n21026) );
  XOR U25700 ( .A(n21025), .B(n21024), .Z(n21022) );
  XOR U25701 ( .A(y[971]), .B(x[971]), .Z(n21024) );
  XOR U25702 ( .A(y[970]), .B(x[970]), .Z(n21025) );
  XOR U25703 ( .A(y[969]), .B(x[969]), .Z(n21023) );
  XOR U25704 ( .A(n21017), .B(n21016), .Z(n21027) );
  XOR U25705 ( .A(n21019), .B(n21018), .Z(n21016) );
  XOR U25706 ( .A(y[968]), .B(x[968]), .Z(n21018) );
  XOR U25707 ( .A(y[967]), .B(x[967]), .Z(n21019) );
  XOR U25708 ( .A(y[966]), .B(x[966]), .Z(n21017) );
  NAND U25709 ( .A(n21080), .B(n21081), .Z(N28413) );
  NAND U25710 ( .A(n21082), .B(n21083), .Z(n21081) );
  NANDN U25711 ( .A(n21084), .B(n21085), .Z(n21083) );
  NANDN U25712 ( .A(n21085), .B(n21084), .Z(n21080) );
  XOR U25713 ( .A(n21084), .B(n21086), .Z(N28412) );
  XNOR U25714 ( .A(n21082), .B(n21085), .Z(n21086) );
  NAND U25715 ( .A(n21087), .B(n21088), .Z(n21085) );
  NAND U25716 ( .A(n21089), .B(n21090), .Z(n21088) );
  NANDN U25717 ( .A(n21091), .B(n21092), .Z(n21090) );
  NANDN U25718 ( .A(n21092), .B(n21091), .Z(n21087) );
  AND U25719 ( .A(n21093), .B(n21094), .Z(n21082) );
  NAND U25720 ( .A(n21095), .B(n21096), .Z(n21094) );
  OR U25721 ( .A(n21097), .B(n21098), .Z(n21096) );
  NAND U25722 ( .A(n21098), .B(n21097), .Z(n21093) );
  IV U25723 ( .A(n21099), .Z(n21098) );
  AND U25724 ( .A(n21100), .B(n21101), .Z(n21084) );
  NAND U25725 ( .A(n21102), .B(n21103), .Z(n21101) );
  NANDN U25726 ( .A(n21104), .B(n21105), .Z(n21103) );
  NANDN U25727 ( .A(n21105), .B(n21104), .Z(n21100) );
  XOR U25728 ( .A(n21097), .B(n21106), .Z(N28411) );
  XOR U25729 ( .A(n21095), .B(n21099), .Z(n21106) );
  XNOR U25730 ( .A(n21092), .B(n21107), .Z(n21099) );
  XNOR U25731 ( .A(n21089), .B(n21091), .Z(n21107) );
  AND U25732 ( .A(n21108), .B(n21109), .Z(n21091) );
  NANDN U25733 ( .A(n21110), .B(n21111), .Z(n21109) );
  NANDN U25734 ( .A(n21112), .B(n21113), .Z(n21111) );
  IV U25735 ( .A(n21114), .Z(n21113) );
  NAND U25736 ( .A(n21114), .B(n21112), .Z(n21108) );
  AND U25737 ( .A(n21115), .B(n21116), .Z(n21089) );
  NAND U25738 ( .A(n21117), .B(n21118), .Z(n21116) );
  OR U25739 ( .A(n21119), .B(n21120), .Z(n21118) );
  NAND U25740 ( .A(n21120), .B(n21119), .Z(n21115) );
  IV U25741 ( .A(n21121), .Z(n21120) );
  NAND U25742 ( .A(n21122), .B(n21123), .Z(n21092) );
  NANDN U25743 ( .A(n21124), .B(n21125), .Z(n21123) );
  NAND U25744 ( .A(n21126), .B(n21127), .Z(n21125) );
  OR U25745 ( .A(n21127), .B(n21126), .Z(n21122) );
  IV U25746 ( .A(n21128), .Z(n21126) );
  AND U25747 ( .A(n21129), .B(n21130), .Z(n21095) );
  NAND U25748 ( .A(n21131), .B(n21132), .Z(n21130) );
  NANDN U25749 ( .A(n21133), .B(n21134), .Z(n21132) );
  NANDN U25750 ( .A(n21134), .B(n21133), .Z(n21129) );
  XOR U25751 ( .A(n21105), .B(n21135), .Z(n21097) );
  XNOR U25752 ( .A(n21102), .B(n21104), .Z(n21135) );
  AND U25753 ( .A(n21136), .B(n21137), .Z(n21104) );
  NANDN U25754 ( .A(n21138), .B(n21139), .Z(n21137) );
  NANDN U25755 ( .A(n21140), .B(n21141), .Z(n21139) );
  IV U25756 ( .A(n21142), .Z(n21141) );
  NAND U25757 ( .A(n21142), .B(n21140), .Z(n21136) );
  AND U25758 ( .A(n21143), .B(n21144), .Z(n21102) );
  NAND U25759 ( .A(n21145), .B(n21146), .Z(n21144) );
  OR U25760 ( .A(n21147), .B(n21148), .Z(n21146) );
  NAND U25761 ( .A(n21148), .B(n21147), .Z(n21143) );
  IV U25762 ( .A(n21149), .Z(n21148) );
  NAND U25763 ( .A(n21150), .B(n21151), .Z(n21105) );
  NANDN U25764 ( .A(n21152), .B(n21153), .Z(n21151) );
  NAND U25765 ( .A(n21154), .B(n21155), .Z(n21153) );
  OR U25766 ( .A(n21155), .B(n21154), .Z(n21150) );
  IV U25767 ( .A(n21156), .Z(n21154) );
  XOR U25768 ( .A(n21131), .B(n21157), .Z(N28410) );
  XNOR U25769 ( .A(n21134), .B(n21133), .Z(n21157) );
  XNOR U25770 ( .A(n21145), .B(n21158), .Z(n21133) );
  XOR U25771 ( .A(n21149), .B(n21147), .Z(n21158) );
  XOR U25772 ( .A(n21155), .B(n21159), .Z(n21147) );
  XOR U25773 ( .A(n21152), .B(n21156), .Z(n21159) );
  NAND U25774 ( .A(n21160), .B(n21161), .Z(n21156) );
  NAND U25775 ( .A(n21162), .B(n21163), .Z(n21161) );
  NAND U25776 ( .A(n21164), .B(n21165), .Z(n21160) );
  AND U25777 ( .A(n21166), .B(n21167), .Z(n21152) );
  NAND U25778 ( .A(n21168), .B(n21169), .Z(n21167) );
  NAND U25779 ( .A(n21170), .B(n21171), .Z(n21166) );
  NANDN U25780 ( .A(n21172), .B(n21173), .Z(n21155) );
  NANDN U25781 ( .A(n21174), .B(n21175), .Z(n21149) );
  XNOR U25782 ( .A(n21140), .B(n21176), .Z(n21145) );
  XOR U25783 ( .A(n21138), .B(n21142), .Z(n21176) );
  NAND U25784 ( .A(n21177), .B(n21178), .Z(n21142) );
  NAND U25785 ( .A(n21179), .B(n21180), .Z(n21178) );
  NAND U25786 ( .A(n21181), .B(n21182), .Z(n21177) );
  AND U25787 ( .A(n21183), .B(n21184), .Z(n21138) );
  NAND U25788 ( .A(n21185), .B(n21186), .Z(n21184) );
  NAND U25789 ( .A(n21187), .B(n21188), .Z(n21183) );
  AND U25790 ( .A(n21189), .B(n21190), .Z(n21140) );
  NAND U25791 ( .A(n21191), .B(n21192), .Z(n21134) );
  XNOR U25792 ( .A(n21117), .B(n21193), .Z(n21131) );
  XOR U25793 ( .A(n21121), .B(n21119), .Z(n21193) );
  XOR U25794 ( .A(n21127), .B(n21194), .Z(n21119) );
  XOR U25795 ( .A(n21124), .B(n21128), .Z(n21194) );
  NAND U25796 ( .A(n21195), .B(n21196), .Z(n21128) );
  NAND U25797 ( .A(n21197), .B(n21198), .Z(n21196) );
  NAND U25798 ( .A(n21199), .B(n21200), .Z(n21195) );
  AND U25799 ( .A(n21201), .B(n21202), .Z(n21124) );
  NAND U25800 ( .A(n21203), .B(n21204), .Z(n21202) );
  NAND U25801 ( .A(n21205), .B(n21206), .Z(n21201) );
  NANDN U25802 ( .A(n21207), .B(n21208), .Z(n21127) );
  NANDN U25803 ( .A(n21209), .B(n21210), .Z(n21121) );
  XNOR U25804 ( .A(n21112), .B(n21211), .Z(n21117) );
  XOR U25805 ( .A(n21110), .B(n21114), .Z(n21211) );
  NAND U25806 ( .A(n21212), .B(n21213), .Z(n21114) );
  NAND U25807 ( .A(n21214), .B(n21215), .Z(n21213) );
  NAND U25808 ( .A(n21216), .B(n21217), .Z(n21212) );
  AND U25809 ( .A(n21218), .B(n21219), .Z(n21110) );
  NAND U25810 ( .A(n21220), .B(n21221), .Z(n21219) );
  NAND U25811 ( .A(n21222), .B(n21223), .Z(n21218) );
  AND U25812 ( .A(n21224), .B(n21225), .Z(n21112) );
  XOR U25813 ( .A(n21192), .B(n21191), .Z(N28409) );
  XNOR U25814 ( .A(n21210), .B(n21209), .Z(n21191) );
  XNOR U25815 ( .A(n21224), .B(n21225), .Z(n21209) );
  XOR U25816 ( .A(n21221), .B(n21220), .Z(n21225) );
  XOR U25817 ( .A(y[963]), .B(x[963]), .Z(n21220) );
  XOR U25818 ( .A(n21223), .B(n21222), .Z(n21221) );
  XOR U25819 ( .A(y[965]), .B(x[965]), .Z(n21222) );
  XOR U25820 ( .A(y[964]), .B(x[964]), .Z(n21223) );
  XOR U25821 ( .A(n21215), .B(n21214), .Z(n21224) );
  XOR U25822 ( .A(n21217), .B(n21216), .Z(n21214) );
  XOR U25823 ( .A(y[962]), .B(x[962]), .Z(n21216) );
  XOR U25824 ( .A(y[961]), .B(x[961]), .Z(n21217) );
  XOR U25825 ( .A(y[960]), .B(x[960]), .Z(n21215) );
  XNOR U25826 ( .A(n21208), .B(n21207), .Z(n21210) );
  XNOR U25827 ( .A(n21204), .B(n21203), .Z(n21207) );
  XOR U25828 ( .A(n21206), .B(n21205), .Z(n21203) );
  XOR U25829 ( .A(y[959]), .B(x[959]), .Z(n21205) );
  XOR U25830 ( .A(y[958]), .B(x[958]), .Z(n21206) );
  XOR U25831 ( .A(y[957]), .B(x[957]), .Z(n21204) );
  XOR U25832 ( .A(n21198), .B(n21197), .Z(n21208) );
  XOR U25833 ( .A(n21200), .B(n21199), .Z(n21197) );
  XOR U25834 ( .A(y[956]), .B(x[956]), .Z(n21199) );
  XOR U25835 ( .A(y[955]), .B(x[955]), .Z(n21200) );
  XOR U25836 ( .A(y[954]), .B(x[954]), .Z(n21198) );
  XNOR U25837 ( .A(n21175), .B(n21174), .Z(n21192) );
  XNOR U25838 ( .A(n21189), .B(n21190), .Z(n21174) );
  XOR U25839 ( .A(n21186), .B(n21185), .Z(n21190) );
  XOR U25840 ( .A(y[951]), .B(x[951]), .Z(n21185) );
  XOR U25841 ( .A(n21188), .B(n21187), .Z(n21186) );
  XOR U25842 ( .A(y[953]), .B(x[953]), .Z(n21187) );
  XOR U25843 ( .A(y[952]), .B(x[952]), .Z(n21188) );
  XOR U25844 ( .A(n21180), .B(n21179), .Z(n21189) );
  XOR U25845 ( .A(n21182), .B(n21181), .Z(n21179) );
  XOR U25846 ( .A(y[950]), .B(x[950]), .Z(n21181) );
  XOR U25847 ( .A(y[949]), .B(x[949]), .Z(n21182) );
  XOR U25848 ( .A(y[948]), .B(x[948]), .Z(n21180) );
  XNOR U25849 ( .A(n21173), .B(n21172), .Z(n21175) );
  XNOR U25850 ( .A(n21169), .B(n21168), .Z(n21172) );
  XOR U25851 ( .A(n21171), .B(n21170), .Z(n21168) );
  XOR U25852 ( .A(y[947]), .B(x[947]), .Z(n21170) );
  XOR U25853 ( .A(y[946]), .B(x[946]), .Z(n21171) );
  XOR U25854 ( .A(y[945]), .B(x[945]), .Z(n21169) );
  XOR U25855 ( .A(n21163), .B(n21162), .Z(n21173) );
  XOR U25856 ( .A(n21165), .B(n21164), .Z(n21162) );
  XOR U25857 ( .A(y[944]), .B(x[944]), .Z(n21164) );
  XOR U25858 ( .A(y[943]), .B(x[943]), .Z(n21165) );
  XOR U25859 ( .A(y[942]), .B(x[942]), .Z(n21163) );
  NAND U25860 ( .A(n21226), .B(n21227), .Z(N28401) );
  NAND U25861 ( .A(n21228), .B(n21229), .Z(n21227) );
  NANDN U25862 ( .A(n21230), .B(n21231), .Z(n21229) );
  NANDN U25863 ( .A(n21231), .B(n21230), .Z(n21226) );
  XOR U25864 ( .A(n21230), .B(n21232), .Z(N28400) );
  XNOR U25865 ( .A(n21228), .B(n21231), .Z(n21232) );
  NAND U25866 ( .A(n21233), .B(n21234), .Z(n21231) );
  NAND U25867 ( .A(n21235), .B(n21236), .Z(n21234) );
  NANDN U25868 ( .A(n21237), .B(n21238), .Z(n21236) );
  NANDN U25869 ( .A(n21238), .B(n21237), .Z(n21233) );
  AND U25870 ( .A(n21239), .B(n21240), .Z(n21228) );
  NAND U25871 ( .A(n21241), .B(n21242), .Z(n21240) );
  OR U25872 ( .A(n21243), .B(n21244), .Z(n21242) );
  NAND U25873 ( .A(n21244), .B(n21243), .Z(n21239) );
  IV U25874 ( .A(n21245), .Z(n21244) );
  AND U25875 ( .A(n21246), .B(n21247), .Z(n21230) );
  NAND U25876 ( .A(n21248), .B(n21249), .Z(n21247) );
  NANDN U25877 ( .A(n21250), .B(n21251), .Z(n21249) );
  NANDN U25878 ( .A(n21251), .B(n21250), .Z(n21246) );
  XOR U25879 ( .A(n21243), .B(n21252), .Z(N28399) );
  XOR U25880 ( .A(n21241), .B(n21245), .Z(n21252) );
  XNOR U25881 ( .A(n21238), .B(n21253), .Z(n21245) );
  XNOR U25882 ( .A(n21235), .B(n21237), .Z(n21253) );
  AND U25883 ( .A(n21254), .B(n21255), .Z(n21237) );
  NANDN U25884 ( .A(n21256), .B(n21257), .Z(n21255) );
  NANDN U25885 ( .A(n21258), .B(n21259), .Z(n21257) );
  IV U25886 ( .A(n21260), .Z(n21259) );
  NAND U25887 ( .A(n21260), .B(n21258), .Z(n21254) );
  AND U25888 ( .A(n21261), .B(n21262), .Z(n21235) );
  NAND U25889 ( .A(n21263), .B(n21264), .Z(n21262) );
  OR U25890 ( .A(n21265), .B(n21266), .Z(n21264) );
  NAND U25891 ( .A(n21266), .B(n21265), .Z(n21261) );
  IV U25892 ( .A(n21267), .Z(n21266) );
  NAND U25893 ( .A(n21268), .B(n21269), .Z(n21238) );
  NANDN U25894 ( .A(n21270), .B(n21271), .Z(n21269) );
  NAND U25895 ( .A(n21272), .B(n21273), .Z(n21271) );
  OR U25896 ( .A(n21273), .B(n21272), .Z(n21268) );
  IV U25897 ( .A(n21274), .Z(n21272) );
  AND U25898 ( .A(n21275), .B(n21276), .Z(n21241) );
  NAND U25899 ( .A(n21277), .B(n21278), .Z(n21276) );
  NANDN U25900 ( .A(n21279), .B(n21280), .Z(n21278) );
  NANDN U25901 ( .A(n21280), .B(n21279), .Z(n21275) );
  XOR U25902 ( .A(n21251), .B(n21281), .Z(n21243) );
  XNOR U25903 ( .A(n21248), .B(n21250), .Z(n21281) );
  AND U25904 ( .A(n21282), .B(n21283), .Z(n21250) );
  NANDN U25905 ( .A(n21284), .B(n21285), .Z(n21283) );
  NANDN U25906 ( .A(n21286), .B(n21287), .Z(n21285) );
  IV U25907 ( .A(n21288), .Z(n21287) );
  NAND U25908 ( .A(n21288), .B(n21286), .Z(n21282) );
  AND U25909 ( .A(n21289), .B(n21290), .Z(n21248) );
  NAND U25910 ( .A(n21291), .B(n21292), .Z(n21290) );
  OR U25911 ( .A(n21293), .B(n21294), .Z(n21292) );
  NAND U25912 ( .A(n21294), .B(n21293), .Z(n21289) );
  IV U25913 ( .A(n21295), .Z(n21294) );
  NAND U25914 ( .A(n21296), .B(n21297), .Z(n21251) );
  NANDN U25915 ( .A(n21298), .B(n21299), .Z(n21297) );
  NAND U25916 ( .A(n21300), .B(n21301), .Z(n21299) );
  OR U25917 ( .A(n21301), .B(n21300), .Z(n21296) );
  IV U25918 ( .A(n21302), .Z(n21300) );
  XOR U25919 ( .A(n21277), .B(n21303), .Z(N28398) );
  XNOR U25920 ( .A(n21280), .B(n21279), .Z(n21303) );
  XNOR U25921 ( .A(n21291), .B(n21304), .Z(n21279) );
  XOR U25922 ( .A(n21295), .B(n21293), .Z(n21304) );
  XOR U25923 ( .A(n21301), .B(n21305), .Z(n21293) );
  XOR U25924 ( .A(n21298), .B(n21302), .Z(n21305) );
  NAND U25925 ( .A(n21306), .B(n21307), .Z(n21302) );
  NAND U25926 ( .A(n21308), .B(n21309), .Z(n21307) );
  NAND U25927 ( .A(n21310), .B(n21311), .Z(n21306) );
  AND U25928 ( .A(n21312), .B(n21313), .Z(n21298) );
  NAND U25929 ( .A(n21314), .B(n21315), .Z(n21313) );
  NAND U25930 ( .A(n21316), .B(n21317), .Z(n21312) );
  NANDN U25931 ( .A(n21318), .B(n21319), .Z(n21301) );
  NANDN U25932 ( .A(n21320), .B(n21321), .Z(n21295) );
  XNOR U25933 ( .A(n21286), .B(n21322), .Z(n21291) );
  XOR U25934 ( .A(n21284), .B(n21288), .Z(n21322) );
  NAND U25935 ( .A(n21323), .B(n21324), .Z(n21288) );
  NAND U25936 ( .A(n21325), .B(n21326), .Z(n21324) );
  NAND U25937 ( .A(n21327), .B(n21328), .Z(n21323) );
  AND U25938 ( .A(n21329), .B(n21330), .Z(n21284) );
  NAND U25939 ( .A(n21331), .B(n21332), .Z(n21330) );
  NAND U25940 ( .A(n21333), .B(n21334), .Z(n21329) );
  AND U25941 ( .A(n21335), .B(n21336), .Z(n21286) );
  NAND U25942 ( .A(n21337), .B(n21338), .Z(n21280) );
  XNOR U25943 ( .A(n21263), .B(n21339), .Z(n21277) );
  XOR U25944 ( .A(n21267), .B(n21265), .Z(n21339) );
  XOR U25945 ( .A(n21273), .B(n21340), .Z(n21265) );
  XOR U25946 ( .A(n21270), .B(n21274), .Z(n21340) );
  NAND U25947 ( .A(n21341), .B(n21342), .Z(n21274) );
  NAND U25948 ( .A(n21343), .B(n21344), .Z(n21342) );
  NAND U25949 ( .A(n21345), .B(n21346), .Z(n21341) );
  AND U25950 ( .A(n21347), .B(n21348), .Z(n21270) );
  NAND U25951 ( .A(n21349), .B(n21350), .Z(n21348) );
  NAND U25952 ( .A(n21351), .B(n21352), .Z(n21347) );
  NANDN U25953 ( .A(n21353), .B(n21354), .Z(n21273) );
  NANDN U25954 ( .A(n21355), .B(n21356), .Z(n21267) );
  XNOR U25955 ( .A(n21258), .B(n21357), .Z(n21263) );
  XOR U25956 ( .A(n21256), .B(n21260), .Z(n21357) );
  NAND U25957 ( .A(n21358), .B(n21359), .Z(n21260) );
  NAND U25958 ( .A(n21360), .B(n21361), .Z(n21359) );
  NAND U25959 ( .A(n21362), .B(n21363), .Z(n21358) );
  AND U25960 ( .A(n21364), .B(n21365), .Z(n21256) );
  NAND U25961 ( .A(n21366), .B(n21367), .Z(n21365) );
  NAND U25962 ( .A(n21368), .B(n21369), .Z(n21364) );
  AND U25963 ( .A(n21370), .B(n21371), .Z(n21258) );
  XOR U25964 ( .A(n21338), .B(n21337), .Z(N28397) );
  XNOR U25965 ( .A(n21356), .B(n21355), .Z(n21337) );
  XNOR U25966 ( .A(n21370), .B(n21371), .Z(n21355) );
  XOR U25967 ( .A(n21367), .B(n21366), .Z(n21371) );
  XOR U25968 ( .A(y[939]), .B(x[939]), .Z(n21366) );
  XOR U25969 ( .A(n21369), .B(n21368), .Z(n21367) );
  XOR U25970 ( .A(y[941]), .B(x[941]), .Z(n21368) );
  XOR U25971 ( .A(y[940]), .B(x[940]), .Z(n21369) );
  XOR U25972 ( .A(n21361), .B(n21360), .Z(n21370) );
  XOR U25973 ( .A(n21363), .B(n21362), .Z(n21360) );
  XOR U25974 ( .A(y[938]), .B(x[938]), .Z(n21362) );
  XOR U25975 ( .A(y[937]), .B(x[937]), .Z(n21363) );
  XOR U25976 ( .A(y[936]), .B(x[936]), .Z(n21361) );
  XNOR U25977 ( .A(n21354), .B(n21353), .Z(n21356) );
  XNOR U25978 ( .A(n21350), .B(n21349), .Z(n21353) );
  XOR U25979 ( .A(n21352), .B(n21351), .Z(n21349) );
  XOR U25980 ( .A(y[935]), .B(x[935]), .Z(n21351) );
  XOR U25981 ( .A(y[934]), .B(x[934]), .Z(n21352) );
  XOR U25982 ( .A(y[933]), .B(x[933]), .Z(n21350) );
  XOR U25983 ( .A(n21344), .B(n21343), .Z(n21354) );
  XOR U25984 ( .A(n21346), .B(n21345), .Z(n21343) );
  XOR U25985 ( .A(y[932]), .B(x[932]), .Z(n21345) );
  XOR U25986 ( .A(y[931]), .B(x[931]), .Z(n21346) );
  XOR U25987 ( .A(y[930]), .B(x[930]), .Z(n21344) );
  XNOR U25988 ( .A(n21321), .B(n21320), .Z(n21338) );
  XNOR U25989 ( .A(n21335), .B(n21336), .Z(n21320) );
  XOR U25990 ( .A(n21332), .B(n21331), .Z(n21336) );
  XOR U25991 ( .A(y[927]), .B(x[927]), .Z(n21331) );
  XOR U25992 ( .A(n21334), .B(n21333), .Z(n21332) );
  XOR U25993 ( .A(y[929]), .B(x[929]), .Z(n21333) );
  XOR U25994 ( .A(y[928]), .B(x[928]), .Z(n21334) );
  XOR U25995 ( .A(n21326), .B(n21325), .Z(n21335) );
  XOR U25996 ( .A(n21328), .B(n21327), .Z(n21325) );
  XOR U25997 ( .A(y[926]), .B(x[926]), .Z(n21327) );
  XOR U25998 ( .A(y[925]), .B(x[925]), .Z(n21328) );
  XOR U25999 ( .A(y[924]), .B(x[924]), .Z(n21326) );
  XNOR U26000 ( .A(n21319), .B(n21318), .Z(n21321) );
  XNOR U26001 ( .A(n21315), .B(n21314), .Z(n21318) );
  XOR U26002 ( .A(n21317), .B(n21316), .Z(n21314) );
  XOR U26003 ( .A(y[923]), .B(x[923]), .Z(n21316) );
  XOR U26004 ( .A(y[922]), .B(x[922]), .Z(n21317) );
  XOR U26005 ( .A(y[921]), .B(x[921]), .Z(n21315) );
  XOR U26006 ( .A(n21309), .B(n21308), .Z(n21319) );
  XOR U26007 ( .A(n21311), .B(n21310), .Z(n21308) );
  XOR U26008 ( .A(y[920]), .B(x[920]), .Z(n21310) );
  XOR U26009 ( .A(y[919]), .B(x[919]), .Z(n21311) );
  XOR U26010 ( .A(y[918]), .B(x[918]), .Z(n21309) );
  NAND U26011 ( .A(n21372), .B(n21373), .Z(N28389) );
  NAND U26012 ( .A(n21374), .B(n21375), .Z(n21373) );
  NANDN U26013 ( .A(n21376), .B(n21377), .Z(n21375) );
  NANDN U26014 ( .A(n21377), .B(n21376), .Z(n21372) );
  XOR U26015 ( .A(n21376), .B(n21378), .Z(N28388) );
  XNOR U26016 ( .A(n21374), .B(n21377), .Z(n21378) );
  NAND U26017 ( .A(n21379), .B(n21380), .Z(n21377) );
  NAND U26018 ( .A(n21381), .B(n21382), .Z(n21380) );
  NANDN U26019 ( .A(n21383), .B(n21384), .Z(n21382) );
  NANDN U26020 ( .A(n21384), .B(n21383), .Z(n21379) );
  AND U26021 ( .A(n21385), .B(n21386), .Z(n21374) );
  NAND U26022 ( .A(n21387), .B(n21388), .Z(n21386) );
  OR U26023 ( .A(n21389), .B(n21390), .Z(n21388) );
  NAND U26024 ( .A(n21390), .B(n21389), .Z(n21385) );
  IV U26025 ( .A(n21391), .Z(n21390) );
  AND U26026 ( .A(n21392), .B(n21393), .Z(n21376) );
  NAND U26027 ( .A(n21394), .B(n21395), .Z(n21393) );
  NANDN U26028 ( .A(n21396), .B(n21397), .Z(n21395) );
  NANDN U26029 ( .A(n21397), .B(n21396), .Z(n21392) );
  XOR U26030 ( .A(n21389), .B(n21398), .Z(N28387) );
  XOR U26031 ( .A(n21387), .B(n21391), .Z(n21398) );
  XNOR U26032 ( .A(n21384), .B(n21399), .Z(n21391) );
  XNOR U26033 ( .A(n21381), .B(n21383), .Z(n21399) );
  AND U26034 ( .A(n21400), .B(n21401), .Z(n21383) );
  NANDN U26035 ( .A(n21402), .B(n21403), .Z(n21401) );
  NANDN U26036 ( .A(n21404), .B(n21405), .Z(n21403) );
  IV U26037 ( .A(n21406), .Z(n21405) );
  NAND U26038 ( .A(n21406), .B(n21404), .Z(n21400) );
  AND U26039 ( .A(n21407), .B(n21408), .Z(n21381) );
  NAND U26040 ( .A(n21409), .B(n21410), .Z(n21408) );
  OR U26041 ( .A(n21411), .B(n21412), .Z(n21410) );
  NAND U26042 ( .A(n21412), .B(n21411), .Z(n21407) );
  IV U26043 ( .A(n21413), .Z(n21412) );
  NAND U26044 ( .A(n21414), .B(n21415), .Z(n21384) );
  NANDN U26045 ( .A(n21416), .B(n21417), .Z(n21415) );
  NAND U26046 ( .A(n21418), .B(n21419), .Z(n21417) );
  OR U26047 ( .A(n21419), .B(n21418), .Z(n21414) );
  IV U26048 ( .A(n21420), .Z(n21418) );
  AND U26049 ( .A(n21421), .B(n21422), .Z(n21387) );
  NAND U26050 ( .A(n21423), .B(n21424), .Z(n21422) );
  NANDN U26051 ( .A(n21425), .B(n21426), .Z(n21424) );
  NANDN U26052 ( .A(n21426), .B(n21425), .Z(n21421) );
  XOR U26053 ( .A(n21397), .B(n21427), .Z(n21389) );
  XNOR U26054 ( .A(n21394), .B(n21396), .Z(n21427) );
  AND U26055 ( .A(n21428), .B(n21429), .Z(n21396) );
  NANDN U26056 ( .A(n21430), .B(n21431), .Z(n21429) );
  NANDN U26057 ( .A(n21432), .B(n21433), .Z(n21431) );
  IV U26058 ( .A(n21434), .Z(n21433) );
  NAND U26059 ( .A(n21434), .B(n21432), .Z(n21428) );
  AND U26060 ( .A(n21435), .B(n21436), .Z(n21394) );
  NAND U26061 ( .A(n21437), .B(n21438), .Z(n21436) );
  OR U26062 ( .A(n21439), .B(n21440), .Z(n21438) );
  NAND U26063 ( .A(n21440), .B(n21439), .Z(n21435) );
  IV U26064 ( .A(n21441), .Z(n21440) );
  NAND U26065 ( .A(n21442), .B(n21443), .Z(n21397) );
  NANDN U26066 ( .A(n21444), .B(n21445), .Z(n21443) );
  NAND U26067 ( .A(n21446), .B(n21447), .Z(n21445) );
  OR U26068 ( .A(n21447), .B(n21446), .Z(n21442) );
  IV U26069 ( .A(n21448), .Z(n21446) );
  XOR U26070 ( .A(n21423), .B(n21449), .Z(N28386) );
  XNOR U26071 ( .A(n21426), .B(n21425), .Z(n21449) );
  XNOR U26072 ( .A(n21437), .B(n21450), .Z(n21425) );
  XOR U26073 ( .A(n21441), .B(n21439), .Z(n21450) );
  XOR U26074 ( .A(n21447), .B(n21451), .Z(n21439) );
  XOR U26075 ( .A(n21444), .B(n21448), .Z(n21451) );
  NAND U26076 ( .A(n21452), .B(n21453), .Z(n21448) );
  NAND U26077 ( .A(n21454), .B(n21455), .Z(n21453) );
  NAND U26078 ( .A(n21456), .B(n21457), .Z(n21452) );
  AND U26079 ( .A(n21458), .B(n21459), .Z(n21444) );
  NAND U26080 ( .A(n21460), .B(n21461), .Z(n21459) );
  NAND U26081 ( .A(n21462), .B(n21463), .Z(n21458) );
  NANDN U26082 ( .A(n21464), .B(n21465), .Z(n21447) );
  NANDN U26083 ( .A(n21466), .B(n21467), .Z(n21441) );
  XNOR U26084 ( .A(n21432), .B(n21468), .Z(n21437) );
  XOR U26085 ( .A(n21430), .B(n21434), .Z(n21468) );
  NAND U26086 ( .A(n21469), .B(n21470), .Z(n21434) );
  NAND U26087 ( .A(n21471), .B(n21472), .Z(n21470) );
  NAND U26088 ( .A(n21473), .B(n21474), .Z(n21469) );
  AND U26089 ( .A(n21475), .B(n21476), .Z(n21430) );
  NAND U26090 ( .A(n21477), .B(n21478), .Z(n21476) );
  NAND U26091 ( .A(n21479), .B(n21480), .Z(n21475) );
  AND U26092 ( .A(n21481), .B(n21482), .Z(n21432) );
  NAND U26093 ( .A(n21483), .B(n21484), .Z(n21426) );
  XNOR U26094 ( .A(n21409), .B(n21485), .Z(n21423) );
  XOR U26095 ( .A(n21413), .B(n21411), .Z(n21485) );
  XOR U26096 ( .A(n21419), .B(n21486), .Z(n21411) );
  XOR U26097 ( .A(n21416), .B(n21420), .Z(n21486) );
  NAND U26098 ( .A(n21487), .B(n21488), .Z(n21420) );
  NAND U26099 ( .A(n21489), .B(n21490), .Z(n21488) );
  NAND U26100 ( .A(n21491), .B(n21492), .Z(n21487) );
  AND U26101 ( .A(n21493), .B(n21494), .Z(n21416) );
  NAND U26102 ( .A(n21495), .B(n21496), .Z(n21494) );
  NAND U26103 ( .A(n21497), .B(n21498), .Z(n21493) );
  NANDN U26104 ( .A(n21499), .B(n21500), .Z(n21419) );
  NANDN U26105 ( .A(n21501), .B(n21502), .Z(n21413) );
  XNOR U26106 ( .A(n21404), .B(n21503), .Z(n21409) );
  XOR U26107 ( .A(n21402), .B(n21406), .Z(n21503) );
  NAND U26108 ( .A(n21504), .B(n21505), .Z(n21406) );
  NAND U26109 ( .A(n21506), .B(n21507), .Z(n21505) );
  NAND U26110 ( .A(n21508), .B(n21509), .Z(n21504) );
  AND U26111 ( .A(n21510), .B(n21511), .Z(n21402) );
  NAND U26112 ( .A(n21512), .B(n21513), .Z(n21511) );
  NAND U26113 ( .A(n21514), .B(n21515), .Z(n21510) );
  AND U26114 ( .A(n21516), .B(n21517), .Z(n21404) );
  XOR U26115 ( .A(n21484), .B(n21483), .Z(N28385) );
  XNOR U26116 ( .A(n21502), .B(n21501), .Z(n21483) );
  XNOR U26117 ( .A(n21516), .B(n21517), .Z(n21501) );
  XOR U26118 ( .A(n21513), .B(n21512), .Z(n21517) );
  XOR U26119 ( .A(y[915]), .B(x[915]), .Z(n21512) );
  XOR U26120 ( .A(n21515), .B(n21514), .Z(n21513) );
  XOR U26121 ( .A(y[917]), .B(x[917]), .Z(n21514) );
  XOR U26122 ( .A(y[916]), .B(x[916]), .Z(n21515) );
  XOR U26123 ( .A(n21507), .B(n21506), .Z(n21516) );
  XOR U26124 ( .A(n21509), .B(n21508), .Z(n21506) );
  XOR U26125 ( .A(y[914]), .B(x[914]), .Z(n21508) );
  XOR U26126 ( .A(y[913]), .B(x[913]), .Z(n21509) );
  XOR U26127 ( .A(y[912]), .B(x[912]), .Z(n21507) );
  XNOR U26128 ( .A(n21500), .B(n21499), .Z(n21502) );
  XNOR U26129 ( .A(n21496), .B(n21495), .Z(n21499) );
  XOR U26130 ( .A(n21498), .B(n21497), .Z(n21495) );
  XOR U26131 ( .A(y[911]), .B(x[911]), .Z(n21497) );
  XOR U26132 ( .A(y[910]), .B(x[910]), .Z(n21498) );
  XOR U26133 ( .A(y[909]), .B(x[909]), .Z(n21496) );
  XOR U26134 ( .A(n21490), .B(n21489), .Z(n21500) );
  XOR U26135 ( .A(n21492), .B(n21491), .Z(n21489) );
  XOR U26136 ( .A(y[908]), .B(x[908]), .Z(n21491) );
  XOR U26137 ( .A(y[907]), .B(x[907]), .Z(n21492) );
  XOR U26138 ( .A(y[906]), .B(x[906]), .Z(n21490) );
  XNOR U26139 ( .A(n21467), .B(n21466), .Z(n21484) );
  XNOR U26140 ( .A(n21481), .B(n21482), .Z(n21466) );
  XOR U26141 ( .A(n21478), .B(n21477), .Z(n21482) );
  XOR U26142 ( .A(y[903]), .B(x[903]), .Z(n21477) );
  XOR U26143 ( .A(n21480), .B(n21479), .Z(n21478) );
  XOR U26144 ( .A(y[905]), .B(x[905]), .Z(n21479) );
  XOR U26145 ( .A(y[904]), .B(x[904]), .Z(n21480) );
  XOR U26146 ( .A(n21472), .B(n21471), .Z(n21481) );
  XOR U26147 ( .A(n21474), .B(n21473), .Z(n21471) );
  XOR U26148 ( .A(y[902]), .B(x[902]), .Z(n21473) );
  XOR U26149 ( .A(y[901]), .B(x[901]), .Z(n21474) );
  XOR U26150 ( .A(y[900]), .B(x[900]), .Z(n21472) );
  XNOR U26151 ( .A(n21465), .B(n21464), .Z(n21467) );
  XNOR U26152 ( .A(n21461), .B(n21460), .Z(n21464) );
  XOR U26153 ( .A(n21463), .B(n21462), .Z(n21460) );
  XOR U26154 ( .A(y[899]), .B(x[899]), .Z(n21462) );
  XOR U26155 ( .A(y[898]), .B(x[898]), .Z(n21463) );
  XOR U26156 ( .A(y[897]), .B(x[897]), .Z(n21461) );
  XOR U26157 ( .A(n21455), .B(n21454), .Z(n21465) );
  XOR U26158 ( .A(n21457), .B(n21456), .Z(n21454) );
  XOR U26159 ( .A(y[896]), .B(x[896]), .Z(n21456) );
  XOR U26160 ( .A(y[895]), .B(x[895]), .Z(n21457) );
  XOR U26161 ( .A(y[894]), .B(x[894]), .Z(n21455) );
  NAND U26162 ( .A(n21518), .B(n21519), .Z(N28377) );
  NAND U26163 ( .A(n21520), .B(n21521), .Z(n21519) );
  NANDN U26164 ( .A(n21522), .B(n21523), .Z(n21521) );
  NANDN U26165 ( .A(n21523), .B(n21522), .Z(n21518) );
  XOR U26166 ( .A(n21522), .B(n21524), .Z(N28376) );
  XNOR U26167 ( .A(n21520), .B(n21523), .Z(n21524) );
  NAND U26168 ( .A(n21525), .B(n21526), .Z(n21523) );
  NAND U26169 ( .A(n21527), .B(n21528), .Z(n21526) );
  NANDN U26170 ( .A(n21529), .B(n21530), .Z(n21528) );
  NANDN U26171 ( .A(n21530), .B(n21529), .Z(n21525) );
  AND U26172 ( .A(n21531), .B(n21532), .Z(n21520) );
  NAND U26173 ( .A(n21533), .B(n21534), .Z(n21532) );
  OR U26174 ( .A(n21535), .B(n21536), .Z(n21534) );
  NAND U26175 ( .A(n21536), .B(n21535), .Z(n21531) );
  IV U26176 ( .A(n21537), .Z(n21536) );
  AND U26177 ( .A(n21538), .B(n21539), .Z(n21522) );
  NAND U26178 ( .A(n21540), .B(n21541), .Z(n21539) );
  NANDN U26179 ( .A(n21542), .B(n21543), .Z(n21541) );
  NANDN U26180 ( .A(n21543), .B(n21542), .Z(n21538) );
  XOR U26181 ( .A(n21535), .B(n21544), .Z(N28375) );
  XOR U26182 ( .A(n21533), .B(n21537), .Z(n21544) );
  XNOR U26183 ( .A(n21530), .B(n21545), .Z(n21537) );
  XNOR U26184 ( .A(n21527), .B(n21529), .Z(n21545) );
  AND U26185 ( .A(n21546), .B(n21547), .Z(n21529) );
  NANDN U26186 ( .A(n21548), .B(n21549), .Z(n21547) );
  NANDN U26187 ( .A(n21550), .B(n21551), .Z(n21549) );
  IV U26188 ( .A(n21552), .Z(n21551) );
  NAND U26189 ( .A(n21552), .B(n21550), .Z(n21546) );
  AND U26190 ( .A(n21553), .B(n21554), .Z(n21527) );
  NAND U26191 ( .A(n21555), .B(n21556), .Z(n21554) );
  OR U26192 ( .A(n21557), .B(n21558), .Z(n21556) );
  NAND U26193 ( .A(n21558), .B(n21557), .Z(n21553) );
  IV U26194 ( .A(n21559), .Z(n21558) );
  NAND U26195 ( .A(n21560), .B(n21561), .Z(n21530) );
  NANDN U26196 ( .A(n21562), .B(n21563), .Z(n21561) );
  NAND U26197 ( .A(n21564), .B(n21565), .Z(n21563) );
  OR U26198 ( .A(n21565), .B(n21564), .Z(n21560) );
  IV U26199 ( .A(n21566), .Z(n21564) );
  AND U26200 ( .A(n21567), .B(n21568), .Z(n21533) );
  NAND U26201 ( .A(n21569), .B(n21570), .Z(n21568) );
  NANDN U26202 ( .A(n21571), .B(n21572), .Z(n21570) );
  NANDN U26203 ( .A(n21572), .B(n21571), .Z(n21567) );
  XOR U26204 ( .A(n21543), .B(n21573), .Z(n21535) );
  XNOR U26205 ( .A(n21540), .B(n21542), .Z(n21573) );
  AND U26206 ( .A(n21574), .B(n21575), .Z(n21542) );
  NANDN U26207 ( .A(n21576), .B(n21577), .Z(n21575) );
  NANDN U26208 ( .A(n21578), .B(n21579), .Z(n21577) );
  IV U26209 ( .A(n21580), .Z(n21579) );
  NAND U26210 ( .A(n21580), .B(n21578), .Z(n21574) );
  AND U26211 ( .A(n21581), .B(n21582), .Z(n21540) );
  NAND U26212 ( .A(n21583), .B(n21584), .Z(n21582) );
  OR U26213 ( .A(n21585), .B(n21586), .Z(n21584) );
  NAND U26214 ( .A(n21586), .B(n21585), .Z(n21581) );
  IV U26215 ( .A(n21587), .Z(n21586) );
  NAND U26216 ( .A(n21588), .B(n21589), .Z(n21543) );
  NANDN U26217 ( .A(n21590), .B(n21591), .Z(n21589) );
  NAND U26218 ( .A(n21592), .B(n21593), .Z(n21591) );
  OR U26219 ( .A(n21593), .B(n21592), .Z(n21588) );
  IV U26220 ( .A(n21594), .Z(n21592) );
  XOR U26221 ( .A(n21569), .B(n21595), .Z(N28374) );
  XNOR U26222 ( .A(n21572), .B(n21571), .Z(n21595) );
  XNOR U26223 ( .A(n21583), .B(n21596), .Z(n21571) );
  XOR U26224 ( .A(n21587), .B(n21585), .Z(n21596) );
  XOR U26225 ( .A(n21593), .B(n21597), .Z(n21585) );
  XOR U26226 ( .A(n21590), .B(n21594), .Z(n21597) );
  NAND U26227 ( .A(n21598), .B(n21599), .Z(n21594) );
  NAND U26228 ( .A(n21600), .B(n21601), .Z(n21599) );
  NAND U26229 ( .A(n21602), .B(n21603), .Z(n21598) );
  AND U26230 ( .A(n21604), .B(n21605), .Z(n21590) );
  NAND U26231 ( .A(n21606), .B(n21607), .Z(n21605) );
  NAND U26232 ( .A(n21608), .B(n21609), .Z(n21604) );
  NANDN U26233 ( .A(n21610), .B(n21611), .Z(n21593) );
  NANDN U26234 ( .A(n21612), .B(n21613), .Z(n21587) );
  XNOR U26235 ( .A(n21578), .B(n21614), .Z(n21583) );
  XOR U26236 ( .A(n21576), .B(n21580), .Z(n21614) );
  NAND U26237 ( .A(n21615), .B(n21616), .Z(n21580) );
  NAND U26238 ( .A(n21617), .B(n21618), .Z(n21616) );
  NAND U26239 ( .A(n21619), .B(n21620), .Z(n21615) );
  AND U26240 ( .A(n21621), .B(n21622), .Z(n21576) );
  NAND U26241 ( .A(n21623), .B(n21624), .Z(n21622) );
  NAND U26242 ( .A(n21625), .B(n21626), .Z(n21621) );
  AND U26243 ( .A(n21627), .B(n21628), .Z(n21578) );
  NAND U26244 ( .A(n21629), .B(n21630), .Z(n21572) );
  XNOR U26245 ( .A(n21555), .B(n21631), .Z(n21569) );
  XOR U26246 ( .A(n21559), .B(n21557), .Z(n21631) );
  XOR U26247 ( .A(n21565), .B(n21632), .Z(n21557) );
  XOR U26248 ( .A(n21562), .B(n21566), .Z(n21632) );
  NAND U26249 ( .A(n21633), .B(n21634), .Z(n21566) );
  NAND U26250 ( .A(n21635), .B(n21636), .Z(n21634) );
  NAND U26251 ( .A(n21637), .B(n21638), .Z(n21633) );
  AND U26252 ( .A(n21639), .B(n21640), .Z(n21562) );
  NAND U26253 ( .A(n21641), .B(n21642), .Z(n21640) );
  NAND U26254 ( .A(n21643), .B(n21644), .Z(n21639) );
  NANDN U26255 ( .A(n21645), .B(n21646), .Z(n21565) );
  NANDN U26256 ( .A(n21647), .B(n21648), .Z(n21559) );
  XNOR U26257 ( .A(n21550), .B(n21649), .Z(n21555) );
  XOR U26258 ( .A(n21548), .B(n21552), .Z(n21649) );
  NAND U26259 ( .A(n21650), .B(n21651), .Z(n21552) );
  NAND U26260 ( .A(n21652), .B(n21653), .Z(n21651) );
  NAND U26261 ( .A(n21654), .B(n21655), .Z(n21650) );
  AND U26262 ( .A(n21656), .B(n21657), .Z(n21548) );
  NAND U26263 ( .A(n21658), .B(n21659), .Z(n21657) );
  NAND U26264 ( .A(n21660), .B(n21661), .Z(n21656) );
  AND U26265 ( .A(n21662), .B(n21663), .Z(n21550) );
  XOR U26266 ( .A(n21630), .B(n21629), .Z(N28373) );
  XNOR U26267 ( .A(n21648), .B(n21647), .Z(n21629) );
  XNOR U26268 ( .A(n21662), .B(n21663), .Z(n21647) );
  XOR U26269 ( .A(n21659), .B(n21658), .Z(n21663) );
  XOR U26270 ( .A(y[891]), .B(x[891]), .Z(n21658) );
  XOR U26271 ( .A(n21661), .B(n21660), .Z(n21659) );
  XOR U26272 ( .A(y[893]), .B(x[893]), .Z(n21660) );
  XOR U26273 ( .A(y[892]), .B(x[892]), .Z(n21661) );
  XOR U26274 ( .A(n21653), .B(n21652), .Z(n21662) );
  XOR U26275 ( .A(n21655), .B(n21654), .Z(n21652) );
  XOR U26276 ( .A(y[890]), .B(x[890]), .Z(n21654) );
  XOR U26277 ( .A(y[889]), .B(x[889]), .Z(n21655) );
  XOR U26278 ( .A(y[888]), .B(x[888]), .Z(n21653) );
  XNOR U26279 ( .A(n21646), .B(n21645), .Z(n21648) );
  XNOR U26280 ( .A(n21642), .B(n21641), .Z(n21645) );
  XOR U26281 ( .A(n21644), .B(n21643), .Z(n21641) );
  XOR U26282 ( .A(y[887]), .B(x[887]), .Z(n21643) );
  XOR U26283 ( .A(y[886]), .B(x[886]), .Z(n21644) );
  XOR U26284 ( .A(y[885]), .B(x[885]), .Z(n21642) );
  XOR U26285 ( .A(n21636), .B(n21635), .Z(n21646) );
  XOR U26286 ( .A(n21638), .B(n21637), .Z(n21635) );
  XOR U26287 ( .A(y[884]), .B(x[884]), .Z(n21637) );
  XOR U26288 ( .A(y[883]), .B(x[883]), .Z(n21638) );
  XOR U26289 ( .A(y[882]), .B(x[882]), .Z(n21636) );
  XNOR U26290 ( .A(n21613), .B(n21612), .Z(n21630) );
  XNOR U26291 ( .A(n21627), .B(n21628), .Z(n21612) );
  XOR U26292 ( .A(n21624), .B(n21623), .Z(n21628) );
  XOR U26293 ( .A(y[879]), .B(x[879]), .Z(n21623) );
  XOR U26294 ( .A(n21626), .B(n21625), .Z(n21624) );
  XOR U26295 ( .A(y[881]), .B(x[881]), .Z(n21625) );
  XOR U26296 ( .A(y[880]), .B(x[880]), .Z(n21626) );
  XOR U26297 ( .A(n21618), .B(n21617), .Z(n21627) );
  XOR U26298 ( .A(n21620), .B(n21619), .Z(n21617) );
  XOR U26299 ( .A(y[878]), .B(x[878]), .Z(n21619) );
  XOR U26300 ( .A(y[877]), .B(x[877]), .Z(n21620) );
  XOR U26301 ( .A(y[876]), .B(x[876]), .Z(n21618) );
  XNOR U26302 ( .A(n21611), .B(n21610), .Z(n21613) );
  XNOR U26303 ( .A(n21607), .B(n21606), .Z(n21610) );
  XOR U26304 ( .A(n21609), .B(n21608), .Z(n21606) );
  XOR U26305 ( .A(y[875]), .B(x[875]), .Z(n21608) );
  XOR U26306 ( .A(y[874]), .B(x[874]), .Z(n21609) );
  XOR U26307 ( .A(y[873]), .B(x[873]), .Z(n21607) );
  XOR U26308 ( .A(n21601), .B(n21600), .Z(n21611) );
  XOR U26309 ( .A(n21603), .B(n21602), .Z(n21600) );
  XOR U26310 ( .A(y[872]), .B(x[872]), .Z(n21602) );
  XOR U26311 ( .A(y[871]), .B(x[871]), .Z(n21603) );
  XOR U26312 ( .A(y[870]), .B(x[870]), .Z(n21601) );
  NAND U26313 ( .A(n21664), .B(n21665), .Z(N28365) );
  NAND U26314 ( .A(n21666), .B(n21667), .Z(n21665) );
  NANDN U26315 ( .A(n21668), .B(n21669), .Z(n21667) );
  NANDN U26316 ( .A(n21669), .B(n21668), .Z(n21664) );
  XOR U26317 ( .A(n21668), .B(n21670), .Z(N28364) );
  XNOR U26318 ( .A(n21666), .B(n21669), .Z(n21670) );
  NAND U26319 ( .A(n21671), .B(n21672), .Z(n21669) );
  NAND U26320 ( .A(n21673), .B(n21674), .Z(n21672) );
  NANDN U26321 ( .A(n21675), .B(n21676), .Z(n21674) );
  NANDN U26322 ( .A(n21676), .B(n21675), .Z(n21671) );
  AND U26323 ( .A(n21677), .B(n21678), .Z(n21666) );
  NAND U26324 ( .A(n21679), .B(n21680), .Z(n21678) );
  OR U26325 ( .A(n21681), .B(n21682), .Z(n21680) );
  NAND U26326 ( .A(n21682), .B(n21681), .Z(n21677) );
  IV U26327 ( .A(n21683), .Z(n21682) );
  AND U26328 ( .A(n21684), .B(n21685), .Z(n21668) );
  NAND U26329 ( .A(n21686), .B(n21687), .Z(n21685) );
  NANDN U26330 ( .A(n21688), .B(n21689), .Z(n21687) );
  NANDN U26331 ( .A(n21689), .B(n21688), .Z(n21684) );
  XOR U26332 ( .A(n21681), .B(n21690), .Z(N28363) );
  XOR U26333 ( .A(n21679), .B(n21683), .Z(n21690) );
  XNOR U26334 ( .A(n21676), .B(n21691), .Z(n21683) );
  XNOR U26335 ( .A(n21673), .B(n21675), .Z(n21691) );
  AND U26336 ( .A(n21692), .B(n21693), .Z(n21675) );
  NANDN U26337 ( .A(n21694), .B(n21695), .Z(n21693) );
  NANDN U26338 ( .A(n21696), .B(n21697), .Z(n21695) );
  IV U26339 ( .A(n21698), .Z(n21697) );
  NAND U26340 ( .A(n21698), .B(n21696), .Z(n21692) );
  AND U26341 ( .A(n21699), .B(n21700), .Z(n21673) );
  NAND U26342 ( .A(n21701), .B(n21702), .Z(n21700) );
  OR U26343 ( .A(n21703), .B(n21704), .Z(n21702) );
  NAND U26344 ( .A(n21704), .B(n21703), .Z(n21699) );
  IV U26345 ( .A(n21705), .Z(n21704) );
  NAND U26346 ( .A(n21706), .B(n21707), .Z(n21676) );
  NANDN U26347 ( .A(n21708), .B(n21709), .Z(n21707) );
  NAND U26348 ( .A(n21710), .B(n21711), .Z(n21709) );
  OR U26349 ( .A(n21711), .B(n21710), .Z(n21706) );
  IV U26350 ( .A(n21712), .Z(n21710) );
  AND U26351 ( .A(n21713), .B(n21714), .Z(n21679) );
  NAND U26352 ( .A(n21715), .B(n21716), .Z(n21714) );
  NANDN U26353 ( .A(n21717), .B(n21718), .Z(n21716) );
  NANDN U26354 ( .A(n21718), .B(n21717), .Z(n21713) );
  XOR U26355 ( .A(n21689), .B(n21719), .Z(n21681) );
  XNOR U26356 ( .A(n21686), .B(n21688), .Z(n21719) );
  AND U26357 ( .A(n21720), .B(n21721), .Z(n21688) );
  NANDN U26358 ( .A(n21722), .B(n21723), .Z(n21721) );
  NANDN U26359 ( .A(n21724), .B(n21725), .Z(n21723) );
  IV U26360 ( .A(n21726), .Z(n21725) );
  NAND U26361 ( .A(n21726), .B(n21724), .Z(n21720) );
  AND U26362 ( .A(n21727), .B(n21728), .Z(n21686) );
  NAND U26363 ( .A(n21729), .B(n21730), .Z(n21728) );
  OR U26364 ( .A(n21731), .B(n21732), .Z(n21730) );
  NAND U26365 ( .A(n21732), .B(n21731), .Z(n21727) );
  IV U26366 ( .A(n21733), .Z(n21732) );
  NAND U26367 ( .A(n21734), .B(n21735), .Z(n21689) );
  NANDN U26368 ( .A(n21736), .B(n21737), .Z(n21735) );
  NAND U26369 ( .A(n21738), .B(n21739), .Z(n21737) );
  OR U26370 ( .A(n21739), .B(n21738), .Z(n21734) );
  IV U26371 ( .A(n21740), .Z(n21738) );
  XOR U26372 ( .A(n21715), .B(n21741), .Z(N28362) );
  XNOR U26373 ( .A(n21718), .B(n21717), .Z(n21741) );
  XNOR U26374 ( .A(n21729), .B(n21742), .Z(n21717) );
  XOR U26375 ( .A(n21733), .B(n21731), .Z(n21742) );
  XOR U26376 ( .A(n21739), .B(n21743), .Z(n21731) );
  XOR U26377 ( .A(n21736), .B(n21740), .Z(n21743) );
  NAND U26378 ( .A(n21744), .B(n21745), .Z(n21740) );
  NAND U26379 ( .A(n21746), .B(n21747), .Z(n21745) );
  NAND U26380 ( .A(n21748), .B(n21749), .Z(n21744) );
  AND U26381 ( .A(n21750), .B(n21751), .Z(n21736) );
  NAND U26382 ( .A(n21752), .B(n21753), .Z(n21751) );
  NAND U26383 ( .A(n21754), .B(n21755), .Z(n21750) );
  NANDN U26384 ( .A(n21756), .B(n21757), .Z(n21739) );
  NANDN U26385 ( .A(n21758), .B(n21759), .Z(n21733) );
  XNOR U26386 ( .A(n21724), .B(n21760), .Z(n21729) );
  XOR U26387 ( .A(n21722), .B(n21726), .Z(n21760) );
  NAND U26388 ( .A(n21761), .B(n21762), .Z(n21726) );
  NAND U26389 ( .A(n21763), .B(n21764), .Z(n21762) );
  NAND U26390 ( .A(n21765), .B(n21766), .Z(n21761) );
  AND U26391 ( .A(n21767), .B(n21768), .Z(n21722) );
  NAND U26392 ( .A(n21769), .B(n21770), .Z(n21768) );
  NAND U26393 ( .A(n21771), .B(n21772), .Z(n21767) );
  AND U26394 ( .A(n21773), .B(n21774), .Z(n21724) );
  NAND U26395 ( .A(n21775), .B(n21776), .Z(n21718) );
  XNOR U26396 ( .A(n21701), .B(n21777), .Z(n21715) );
  XOR U26397 ( .A(n21705), .B(n21703), .Z(n21777) );
  XOR U26398 ( .A(n21711), .B(n21778), .Z(n21703) );
  XOR U26399 ( .A(n21708), .B(n21712), .Z(n21778) );
  NAND U26400 ( .A(n21779), .B(n21780), .Z(n21712) );
  NAND U26401 ( .A(n21781), .B(n21782), .Z(n21780) );
  NAND U26402 ( .A(n21783), .B(n21784), .Z(n21779) );
  AND U26403 ( .A(n21785), .B(n21786), .Z(n21708) );
  NAND U26404 ( .A(n21787), .B(n21788), .Z(n21786) );
  NAND U26405 ( .A(n21789), .B(n21790), .Z(n21785) );
  NANDN U26406 ( .A(n21791), .B(n21792), .Z(n21711) );
  NANDN U26407 ( .A(n21793), .B(n21794), .Z(n21705) );
  XNOR U26408 ( .A(n21696), .B(n21795), .Z(n21701) );
  XOR U26409 ( .A(n21694), .B(n21698), .Z(n21795) );
  NAND U26410 ( .A(n21796), .B(n21797), .Z(n21698) );
  NAND U26411 ( .A(n21798), .B(n21799), .Z(n21797) );
  NAND U26412 ( .A(n21800), .B(n21801), .Z(n21796) );
  AND U26413 ( .A(n21802), .B(n21803), .Z(n21694) );
  NAND U26414 ( .A(n21804), .B(n21805), .Z(n21803) );
  NAND U26415 ( .A(n21806), .B(n21807), .Z(n21802) );
  AND U26416 ( .A(n21808), .B(n21809), .Z(n21696) );
  XOR U26417 ( .A(n21776), .B(n21775), .Z(N28361) );
  XNOR U26418 ( .A(n21794), .B(n21793), .Z(n21775) );
  XNOR U26419 ( .A(n21808), .B(n21809), .Z(n21793) );
  XOR U26420 ( .A(n21805), .B(n21804), .Z(n21809) );
  XOR U26421 ( .A(y[867]), .B(x[867]), .Z(n21804) );
  XOR U26422 ( .A(n21807), .B(n21806), .Z(n21805) );
  XOR U26423 ( .A(y[869]), .B(x[869]), .Z(n21806) );
  XOR U26424 ( .A(y[868]), .B(x[868]), .Z(n21807) );
  XOR U26425 ( .A(n21799), .B(n21798), .Z(n21808) );
  XOR U26426 ( .A(n21801), .B(n21800), .Z(n21798) );
  XOR U26427 ( .A(y[866]), .B(x[866]), .Z(n21800) );
  XOR U26428 ( .A(y[865]), .B(x[865]), .Z(n21801) );
  XOR U26429 ( .A(y[864]), .B(x[864]), .Z(n21799) );
  XNOR U26430 ( .A(n21792), .B(n21791), .Z(n21794) );
  XNOR U26431 ( .A(n21788), .B(n21787), .Z(n21791) );
  XOR U26432 ( .A(n21790), .B(n21789), .Z(n21787) );
  XOR U26433 ( .A(y[863]), .B(x[863]), .Z(n21789) );
  XOR U26434 ( .A(y[862]), .B(x[862]), .Z(n21790) );
  XOR U26435 ( .A(y[861]), .B(x[861]), .Z(n21788) );
  XOR U26436 ( .A(n21782), .B(n21781), .Z(n21792) );
  XOR U26437 ( .A(n21784), .B(n21783), .Z(n21781) );
  XOR U26438 ( .A(y[860]), .B(x[860]), .Z(n21783) );
  XOR U26439 ( .A(y[859]), .B(x[859]), .Z(n21784) );
  XOR U26440 ( .A(y[858]), .B(x[858]), .Z(n21782) );
  XNOR U26441 ( .A(n21759), .B(n21758), .Z(n21776) );
  XNOR U26442 ( .A(n21773), .B(n21774), .Z(n21758) );
  XOR U26443 ( .A(n21770), .B(n21769), .Z(n21774) );
  XOR U26444 ( .A(y[855]), .B(x[855]), .Z(n21769) );
  XOR U26445 ( .A(n21772), .B(n21771), .Z(n21770) );
  XOR U26446 ( .A(y[857]), .B(x[857]), .Z(n21771) );
  XOR U26447 ( .A(y[856]), .B(x[856]), .Z(n21772) );
  XOR U26448 ( .A(n21764), .B(n21763), .Z(n21773) );
  XOR U26449 ( .A(n21766), .B(n21765), .Z(n21763) );
  XOR U26450 ( .A(y[854]), .B(x[854]), .Z(n21765) );
  XOR U26451 ( .A(y[853]), .B(x[853]), .Z(n21766) );
  XOR U26452 ( .A(y[852]), .B(x[852]), .Z(n21764) );
  XNOR U26453 ( .A(n21757), .B(n21756), .Z(n21759) );
  XNOR U26454 ( .A(n21753), .B(n21752), .Z(n21756) );
  XOR U26455 ( .A(n21755), .B(n21754), .Z(n21752) );
  XOR U26456 ( .A(y[851]), .B(x[851]), .Z(n21754) );
  XOR U26457 ( .A(y[850]), .B(x[850]), .Z(n21755) );
  XOR U26458 ( .A(y[849]), .B(x[849]), .Z(n21753) );
  XOR U26459 ( .A(n21747), .B(n21746), .Z(n21757) );
  XOR U26460 ( .A(n21749), .B(n21748), .Z(n21746) );
  XOR U26461 ( .A(y[848]), .B(x[848]), .Z(n21748) );
  XOR U26462 ( .A(y[847]), .B(x[847]), .Z(n21749) );
  XOR U26463 ( .A(y[846]), .B(x[846]), .Z(n21747) );
  NAND U26464 ( .A(n21810), .B(n21811), .Z(N28353) );
  NAND U26465 ( .A(n21812), .B(n21813), .Z(n21811) );
  NANDN U26466 ( .A(n21814), .B(n21815), .Z(n21813) );
  NANDN U26467 ( .A(n21815), .B(n21814), .Z(n21810) );
  XOR U26468 ( .A(n21814), .B(n21816), .Z(N28352) );
  XNOR U26469 ( .A(n21812), .B(n21815), .Z(n21816) );
  NAND U26470 ( .A(n21817), .B(n21818), .Z(n21815) );
  NAND U26471 ( .A(n21819), .B(n21820), .Z(n21818) );
  NANDN U26472 ( .A(n21821), .B(n21822), .Z(n21820) );
  NANDN U26473 ( .A(n21822), .B(n21821), .Z(n21817) );
  AND U26474 ( .A(n21823), .B(n21824), .Z(n21812) );
  NAND U26475 ( .A(n21825), .B(n21826), .Z(n21824) );
  OR U26476 ( .A(n21827), .B(n21828), .Z(n21826) );
  NAND U26477 ( .A(n21828), .B(n21827), .Z(n21823) );
  IV U26478 ( .A(n21829), .Z(n21828) );
  AND U26479 ( .A(n21830), .B(n21831), .Z(n21814) );
  NAND U26480 ( .A(n21832), .B(n21833), .Z(n21831) );
  NANDN U26481 ( .A(n21834), .B(n21835), .Z(n21833) );
  NANDN U26482 ( .A(n21835), .B(n21834), .Z(n21830) );
  XOR U26483 ( .A(n21827), .B(n21836), .Z(N28351) );
  XOR U26484 ( .A(n21825), .B(n21829), .Z(n21836) );
  XNOR U26485 ( .A(n21822), .B(n21837), .Z(n21829) );
  XNOR U26486 ( .A(n21819), .B(n21821), .Z(n21837) );
  AND U26487 ( .A(n21838), .B(n21839), .Z(n21821) );
  NANDN U26488 ( .A(n21840), .B(n21841), .Z(n21839) );
  NANDN U26489 ( .A(n21842), .B(n21843), .Z(n21841) );
  IV U26490 ( .A(n21844), .Z(n21843) );
  NAND U26491 ( .A(n21844), .B(n21842), .Z(n21838) );
  AND U26492 ( .A(n21845), .B(n21846), .Z(n21819) );
  NAND U26493 ( .A(n21847), .B(n21848), .Z(n21846) );
  OR U26494 ( .A(n21849), .B(n21850), .Z(n21848) );
  NAND U26495 ( .A(n21850), .B(n21849), .Z(n21845) );
  IV U26496 ( .A(n21851), .Z(n21850) );
  NAND U26497 ( .A(n21852), .B(n21853), .Z(n21822) );
  NANDN U26498 ( .A(n21854), .B(n21855), .Z(n21853) );
  NAND U26499 ( .A(n21856), .B(n21857), .Z(n21855) );
  OR U26500 ( .A(n21857), .B(n21856), .Z(n21852) );
  IV U26501 ( .A(n21858), .Z(n21856) );
  AND U26502 ( .A(n21859), .B(n21860), .Z(n21825) );
  NAND U26503 ( .A(n21861), .B(n21862), .Z(n21860) );
  NANDN U26504 ( .A(n21863), .B(n21864), .Z(n21862) );
  NANDN U26505 ( .A(n21864), .B(n21863), .Z(n21859) );
  XOR U26506 ( .A(n21835), .B(n21865), .Z(n21827) );
  XNOR U26507 ( .A(n21832), .B(n21834), .Z(n21865) );
  AND U26508 ( .A(n21866), .B(n21867), .Z(n21834) );
  NANDN U26509 ( .A(n21868), .B(n21869), .Z(n21867) );
  NANDN U26510 ( .A(n21870), .B(n21871), .Z(n21869) );
  IV U26511 ( .A(n21872), .Z(n21871) );
  NAND U26512 ( .A(n21872), .B(n21870), .Z(n21866) );
  AND U26513 ( .A(n21873), .B(n21874), .Z(n21832) );
  NAND U26514 ( .A(n21875), .B(n21876), .Z(n21874) );
  OR U26515 ( .A(n21877), .B(n21878), .Z(n21876) );
  NAND U26516 ( .A(n21878), .B(n21877), .Z(n21873) );
  IV U26517 ( .A(n21879), .Z(n21878) );
  NAND U26518 ( .A(n21880), .B(n21881), .Z(n21835) );
  NANDN U26519 ( .A(n21882), .B(n21883), .Z(n21881) );
  NAND U26520 ( .A(n21884), .B(n21885), .Z(n21883) );
  OR U26521 ( .A(n21885), .B(n21884), .Z(n21880) );
  IV U26522 ( .A(n21886), .Z(n21884) );
  XOR U26523 ( .A(n21861), .B(n21887), .Z(N28350) );
  XNOR U26524 ( .A(n21864), .B(n21863), .Z(n21887) );
  XNOR U26525 ( .A(n21875), .B(n21888), .Z(n21863) );
  XOR U26526 ( .A(n21879), .B(n21877), .Z(n21888) );
  XOR U26527 ( .A(n21885), .B(n21889), .Z(n21877) );
  XOR U26528 ( .A(n21882), .B(n21886), .Z(n21889) );
  NAND U26529 ( .A(n21890), .B(n21891), .Z(n21886) );
  NAND U26530 ( .A(n21892), .B(n21893), .Z(n21891) );
  NAND U26531 ( .A(n21894), .B(n21895), .Z(n21890) );
  AND U26532 ( .A(n21896), .B(n21897), .Z(n21882) );
  NAND U26533 ( .A(n21898), .B(n21899), .Z(n21897) );
  NAND U26534 ( .A(n21900), .B(n21901), .Z(n21896) );
  NANDN U26535 ( .A(n21902), .B(n21903), .Z(n21885) );
  NANDN U26536 ( .A(n21904), .B(n21905), .Z(n21879) );
  XNOR U26537 ( .A(n21870), .B(n21906), .Z(n21875) );
  XOR U26538 ( .A(n21868), .B(n21872), .Z(n21906) );
  NAND U26539 ( .A(n21907), .B(n21908), .Z(n21872) );
  NAND U26540 ( .A(n21909), .B(n21910), .Z(n21908) );
  NAND U26541 ( .A(n21911), .B(n21912), .Z(n21907) );
  AND U26542 ( .A(n21913), .B(n21914), .Z(n21868) );
  NAND U26543 ( .A(n21915), .B(n21916), .Z(n21914) );
  NAND U26544 ( .A(n21917), .B(n21918), .Z(n21913) );
  AND U26545 ( .A(n21919), .B(n21920), .Z(n21870) );
  NAND U26546 ( .A(n21921), .B(n21922), .Z(n21864) );
  XNOR U26547 ( .A(n21847), .B(n21923), .Z(n21861) );
  XOR U26548 ( .A(n21851), .B(n21849), .Z(n21923) );
  XOR U26549 ( .A(n21857), .B(n21924), .Z(n21849) );
  XOR U26550 ( .A(n21854), .B(n21858), .Z(n21924) );
  NAND U26551 ( .A(n21925), .B(n21926), .Z(n21858) );
  NAND U26552 ( .A(n21927), .B(n21928), .Z(n21926) );
  NAND U26553 ( .A(n21929), .B(n21930), .Z(n21925) );
  AND U26554 ( .A(n21931), .B(n21932), .Z(n21854) );
  NAND U26555 ( .A(n21933), .B(n21934), .Z(n21932) );
  NAND U26556 ( .A(n21935), .B(n21936), .Z(n21931) );
  NANDN U26557 ( .A(n21937), .B(n21938), .Z(n21857) );
  NANDN U26558 ( .A(n21939), .B(n21940), .Z(n21851) );
  XNOR U26559 ( .A(n21842), .B(n21941), .Z(n21847) );
  XOR U26560 ( .A(n21840), .B(n21844), .Z(n21941) );
  NAND U26561 ( .A(n21942), .B(n21943), .Z(n21844) );
  NAND U26562 ( .A(n21944), .B(n21945), .Z(n21943) );
  NAND U26563 ( .A(n21946), .B(n21947), .Z(n21942) );
  AND U26564 ( .A(n21948), .B(n21949), .Z(n21840) );
  NAND U26565 ( .A(n21950), .B(n21951), .Z(n21949) );
  NAND U26566 ( .A(n21952), .B(n21953), .Z(n21948) );
  AND U26567 ( .A(n21954), .B(n21955), .Z(n21842) );
  XOR U26568 ( .A(n21922), .B(n21921), .Z(N28349) );
  XNOR U26569 ( .A(n21940), .B(n21939), .Z(n21921) );
  XNOR U26570 ( .A(n21954), .B(n21955), .Z(n21939) );
  XOR U26571 ( .A(n21951), .B(n21950), .Z(n21955) );
  XOR U26572 ( .A(y[843]), .B(x[843]), .Z(n21950) );
  XOR U26573 ( .A(n21953), .B(n21952), .Z(n21951) );
  XOR U26574 ( .A(y[845]), .B(x[845]), .Z(n21952) );
  XOR U26575 ( .A(y[844]), .B(x[844]), .Z(n21953) );
  XOR U26576 ( .A(n21945), .B(n21944), .Z(n21954) );
  XOR U26577 ( .A(n21947), .B(n21946), .Z(n21944) );
  XOR U26578 ( .A(y[842]), .B(x[842]), .Z(n21946) );
  XOR U26579 ( .A(y[841]), .B(x[841]), .Z(n21947) );
  XOR U26580 ( .A(y[840]), .B(x[840]), .Z(n21945) );
  XNOR U26581 ( .A(n21938), .B(n21937), .Z(n21940) );
  XNOR U26582 ( .A(n21934), .B(n21933), .Z(n21937) );
  XOR U26583 ( .A(n21936), .B(n21935), .Z(n21933) );
  XOR U26584 ( .A(y[839]), .B(x[839]), .Z(n21935) );
  XOR U26585 ( .A(y[838]), .B(x[838]), .Z(n21936) );
  XOR U26586 ( .A(y[837]), .B(x[837]), .Z(n21934) );
  XOR U26587 ( .A(n21928), .B(n21927), .Z(n21938) );
  XOR U26588 ( .A(n21930), .B(n21929), .Z(n21927) );
  XOR U26589 ( .A(y[836]), .B(x[836]), .Z(n21929) );
  XOR U26590 ( .A(y[835]), .B(x[835]), .Z(n21930) );
  XOR U26591 ( .A(y[834]), .B(x[834]), .Z(n21928) );
  XNOR U26592 ( .A(n21905), .B(n21904), .Z(n21922) );
  XNOR U26593 ( .A(n21919), .B(n21920), .Z(n21904) );
  XOR U26594 ( .A(n21916), .B(n21915), .Z(n21920) );
  XOR U26595 ( .A(y[831]), .B(x[831]), .Z(n21915) );
  XOR U26596 ( .A(n21918), .B(n21917), .Z(n21916) );
  XOR U26597 ( .A(y[833]), .B(x[833]), .Z(n21917) );
  XOR U26598 ( .A(y[832]), .B(x[832]), .Z(n21918) );
  XOR U26599 ( .A(n21910), .B(n21909), .Z(n21919) );
  XOR U26600 ( .A(n21912), .B(n21911), .Z(n21909) );
  XOR U26601 ( .A(y[830]), .B(x[830]), .Z(n21911) );
  XOR U26602 ( .A(y[829]), .B(x[829]), .Z(n21912) );
  XOR U26603 ( .A(y[828]), .B(x[828]), .Z(n21910) );
  XNOR U26604 ( .A(n21903), .B(n21902), .Z(n21905) );
  XNOR U26605 ( .A(n21899), .B(n21898), .Z(n21902) );
  XOR U26606 ( .A(n21901), .B(n21900), .Z(n21898) );
  XOR U26607 ( .A(y[827]), .B(x[827]), .Z(n21900) );
  XOR U26608 ( .A(y[826]), .B(x[826]), .Z(n21901) );
  XOR U26609 ( .A(y[825]), .B(x[825]), .Z(n21899) );
  XOR U26610 ( .A(n21893), .B(n21892), .Z(n21903) );
  XOR U26611 ( .A(n21895), .B(n21894), .Z(n21892) );
  XOR U26612 ( .A(y[824]), .B(x[824]), .Z(n21894) );
  XOR U26613 ( .A(y[823]), .B(x[823]), .Z(n21895) );
  XOR U26614 ( .A(y[822]), .B(x[822]), .Z(n21893) );
  NAND U26615 ( .A(n21956), .B(n21957), .Z(N28341) );
  NAND U26616 ( .A(n21958), .B(n21959), .Z(n21957) );
  NANDN U26617 ( .A(n21960), .B(n21961), .Z(n21959) );
  NANDN U26618 ( .A(n21961), .B(n21960), .Z(n21956) );
  XOR U26619 ( .A(n21960), .B(n21962), .Z(N28340) );
  XNOR U26620 ( .A(n21958), .B(n21961), .Z(n21962) );
  NAND U26621 ( .A(n21963), .B(n21964), .Z(n21961) );
  NAND U26622 ( .A(n21965), .B(n21966), .Z(n21964) );
  NANDN U26623 ( .A(n21967), .B(n21968), .Z(n21966) );
  NANDN U26624 ( .A(n21968), .B(n21967), .Z(n21963) );
  AND U26625 ( .A(n21969), .B(n21970), .Z(n21958) );
  NAND U26626 ( .A(n21971), .B(n21972), .Z(n21970) );
  OR U26627 ( .A(n21973), .B(n21974), .Z(n21972) );
  NAND U26628 ( .A(n21974), .B(n21973), .Z(n21969) );
  IV U26629 ( .A(n21975), .Z(n21974) );
  AND U26630 ( .A(n21976), .B(n21977), .Z(n21960) );
  NAND U26631 ( .A(n21978), .B(n21979), .Z(n21977) );
  NANDN U26632 ( .A(n21980), .B(n21981), .Z(n21979) );
  NANDN U26633 ( .A(n21981), .B(n21980), .Z(n21976) );
  XOR U26634 ( .A(n21973), .B(n21982), .Z(N28339) );
  XOR U26635 ( .A(n21971), .B(n21975), .Z(n21982) );
  XNOR U26636 ( .A(n21968), .B(n21983), .Z(n21975) );
  XNOR U26637 ( .A(n21965), .B(n21967), .Z(n21983) );
  AND U26638 ( .A(n21984), .B(n21985), .Z(n21967) );
  NANDN U26639 ( .A(n21986), .B(n21987), .Z(n21985) );
  NANDN U26640 ( .A(n21988), .B(n21989), .Z(n21987) );
  IV U26641 ( .A(n21990), .Z(n21989) );
  NAND U26642 ( .A(n21990), .B(n21988), .Z(n21984) );
  AND U26643 ( .A(n21991), .B(n21992), .Z(n21965) );
  NAND U26644 ( .A(n21993), .B(n21994), .Z(n21992) );
  OR U26645 ( .A(n21995), .B(n21996), .Z(n21994) );
  NAND U26646 ( .A(n21996), .B(n21995), .Z(n21991) );
  IV U26647 ( .A(n21997), .Z(n21996) );
  NAND U26648 ( .A(n21998), .B(n21999), .Z(n21968) );
  NANDN U26649 ( .A(n22000), .B(n22001), .Z(n21999) );
  NAND U26650 ( .A(n22002), .B(n22003), .Z(n22001) );
  OR U26651 ( .A(n22003), .B(n22002), .Z(n21998) );
  IV U26652 ( .A(n22004), .Z(n22002) );
  AND U26653 ( .A(n22005), .B(n22006), .Z(n21971) );
  NAND U26654 ( .A(n22007), .B(n22008), .Z(n22006) );
  NANDN U26655 ( .A(n22009), .B(n22010), .Z(n22008) );
  NANDN U26656 ( .A(n22010), .B(n22009), .Z(n22005) );
  XOR U26657 ( .A(n21981), .B(n22011), .Z(n21973) );
  XNOR U26658 ( .A(n21978), .B(n21980), .Z(n22011) );
  AND U26659 ( .A(n22012), .B(n22013), .Z(n21980) );
  NANDN U26660 ( .A(n22014), .B(n22015), .Z(n22013) );
  NANDN U26661 ( .A(n22016), .B(n22017), .Z(n22015) );
  IV U26662 ( .A(n22018), .Z(n22017) );
  NAND U26663 ( .A(n22018), .B(n22016), .Z(n22012) );
  AND U26664 ( .A(n22019), .B(n22020), .Z(n21978) );
  NAND U26665 ( .A(n22021), .B(n22022), .Z(n22020) );
  OR U26666 ( .A(n22023), .B(n22024), .Z(n22022) );
  NAND U26667 ( .A(n22024), .B(n22023), .Z(n22019) );
  IV U26668 ( .A(n22025), .Z(n22024) );
  NAND U26669 ( .A(n22026), .B(n22027), .Z(n21981) );
  NANDN U26670 ( .A(n22028), .B(n22029), .Z(n22027) );
  NAND U26671 ( .A(n22030), .B(n22031), .Z(n22029) );
  OR U26672 ( .A(n22031), .B(n22030), .Z(n22026) );
  IV U26673 ( .A(n22032), .Z(n22030) );
  XOR U26674 ( .A(n22007), .B(n22033), .Z(N28338) );
  XNOR U26675 ( .A(n22010), .B(n22009), .Z(n22033) );
  XNOR U26676 ( .A(n22021), .B(n22034), .Z(n22009) );
  XOR U26677 ( .A(n22025), .B(n22023), .Z(n22034) );
  XOR U26678 ( .A(n22031), .B(n22035), .Z(n22023) );
  XOR U26679 ( .A(n22028), .B(n22032), .Z(n22035) );
  NAND U26680 ( .A(n22036), .B(n22037), .Z(n22032) );
  NAND U26681 ( .A(n22038), .B(n22039), .Z(n22037) );
  NAND U26682 ( .A(n22040), .B(n22041), .Z(n22036) );
  AND U26683 ( .A(n22042), .B(n22043), .Z(n22028) );
  NAND U26684 ( .A(n22044), .B(n22045), .Z(n22043) );
  NAND U26685 ( .A(n22046), .B(n22047), .Z(n22042) );
  NANDN U26686 ( .A(n22048), .B(n22049), .Z(n22031) );
  NANDN U26687 ( .A(n22050), .B(n22051), .Z(n22025) );
  XNOR U26688 ( .A(n22016), .B(n22052), .Z(n22021) );
  XOR U26689 ( .A(n22014), .B(n22018), .Z(n22052) );
  NAND U26690 ( .A(n22053), .B(n22054), .Z(n22018) );
  NAND U26691 ( .A(n22055), .B(n22056), .Z(n22054) );
  NAND U26692 ( .A(n22057), .B(n22058), .Z(n22053) );
  AND U26693 ( .A(n22059), .B(n22060), .Z(n22014) );
  NAND U26694 ( .A(n22061), .B(n22062), .Z(n22060) );
  NAND U26695 ( .A(n22063), .B(n22064), .Z(n22059) );
  AND U26696 ( .A(n22065), .B(n22066), .Z(n22016) );
  NAND U26697 ( .A(n22067), .B(n22068), .Z(n22010) );
  XNOR U26698 ( .A(n21993), .B(n22069), .Z(n22007) );
  XOR U26699 ( .A(n21997), .B(n21995), .Z(n22069) );
  XOR U26700 ( .A(n22003), .B(n22070), .Z(n21995) );
  XOR U26701 ( .A(n22000), .B(n22004), .Z(n22070) );
  NAND U26702 ( .A(n22071), .B(n22072), .Z(n22004) );
  NAND U26703 ( .A(n22073), .B(n22074), .Z(n22072) );
  NAND U26704 ( .A(n22075), .B(n22076), .Z(n22071) );
  AND U26705 ( .A(n22077), .B(n22078), .Z(n22000) );
  NAND U26706 ( .A(n22079), .B(n22080), .Z(n22078) );
  NAND U26707 ( .A(n22081), .B(n22082), .Z(n22077) );
  NANDN U26708 ( .A(n22083), .B(n22084), .Z(n22003) );
  NANDN U26709 ( .A(n22085), .B(n22086), .Z(n21997) );
  XNOR U26710 ( .A(n21988), .B(n22087), .Z(n21993) );
  XOR U26711 ( .A(n21986), .B(n21990), .Z(n22087) );
  NAND U26712 ( .A(n22088), .B(n22089), .Z(n21990) );
  NAND U26713 ( .A(n22090), .B(n22091), .Z(n22089) );
  NAND U26714 ( .A(n22092), .B(n22093), .Z(n22088) );
  AND U26715 ( .A(n22094), .B(n22095), .Z(n21986) );
  NAND U26716 ( .A(n22096), .B(n22097), .Z(n22095) );
  NAND U26717 ( .A(n22098), .B(n22099), .Z(n22094) );
  AND U26718 ( .A(n22100), .B(n22101), .Z(n21988) );
  XOR U26719 ( .A(n22068), .B(n22067), .Z(N28337) );
  XNOR U26720 ( .A(n22086), .B(n22085), .Z(n22067) );
  XNOR U26721 ( .A(n22100), .B(n22101), .Z(n22085) );
  XOR U26722 ( .A(n22097), .B(n22096), .Z(n22101) );
  XOR U26723 ( .A(y[819]), .B(x[819]), .Z(n22096) );
  XOR U26724 ( .A(n22099), .B(n22098), .Z(n22097) );
  XOR U26725 ( .A(y[821]), .B(x[821]), .Z(n22098) );
  XOR U26726 ( .A(y[820]), .B(x[820]), .Z(n22099) );
  XOR U26727 ( .A(n22091), .B(n22090), .Z(n22100) );
  XOR U26728 ( .A(n22093), .B(n22092), .Z(n22090) );
  XOR U26729 ( .A(y[818]), .B(x[818]), .Z(n22092) );
  XOR U26730 ( .A(y[817]), .B(x[817]), .Z(n22093) );
  XOR U26731 ( .A(y[816]), .B(x[816]), .Z(n22091) );
  XNOR U26732 ( .A(n22084), .B(n22083), .Z(n22086) );
  XNOR U26733 ( .A(n22080), .B(n22079), .Z(n22083) );
  XOR U26734 ( .A(n22082), .B(n22081), .Z(n22079) );
  XOR U26735 ( .A(y[815]), .B(x[815]), .Z(n22081) );
  XOR U26736 ( .A(y[814]), .B(x[814]), .Z(n22082) );
  XOR U26737 ( .A(y[813]), .B(x[813]), .Z(n22080) );
  XOR U26738 ( .A(n22074), .B(n22073), .Z(n22084) );
  XOR U26739 ( .A(n22076), .B(n22075), .Z(n22073) );
  XOR U26740 ( .A(y[812]), .B(x[812]), .Z(n22075) );
  XOR U26741 ( .A(y[811]), .B(x[811]), .Z(n22076) );
  XOR U26742 ( .A(y[810]), .B(x[810]), .Z(n22074) );
  XNOR U26743 ( .A(n22051), .B(n22050), .Z(n22068) );
  XNOR U26744 ( .A(n22065), .B(n22066), .Z(n22050) );
  XOR U26745 ( .A(n22062), .B(n22061), .Z(n22066) );
  XOR U26746 ( .A(y[807]), .B(x[807]), .Z(n22061) );
  XOR U26747 ( .A(n22064), .B(n22063), .Z(n22062) );
  XOR U26748 ( .A(y[809]), .B(x[809]), .Z(n22063) );
  XOR U26749 ( .A(y[808]), .B(x[808]), .Z(n22064) );
  XOR U26750 ( .A(n22056), .B(n22055), .Z(n22065) );
  XOR U26751 ( .A(n22058), .B(n22057), .Z(n22055) );
  XOR U26752 ( .A(y[806]), .B(x[806]), .Z(n22057) );
  XOR U26753 ( .A(y[805]), .B(x[805]), .Z(n22058) );
  XOR U26754 ( .A(y[804]), .B(x[804]), .Z(n22056) );
  XNOR U26755 ( .A(n22049), .B(n22048), .Z(n22051) );
  XNOR U26756 ( .A(n22045), .B(n22044), .Z(n22048) );
  XOR U26757 ( .A(n22047), .B(n22046), .Z(n22044) );
  XOR U26758 ( .A(y[803]), .B(x[803]), .Z(n22046) );
  XOR U26759 ( .A(y[802]), .B(x[802]), .Z(n22047) );
  XOR U26760 ( .A(y[801]), .B(x[801]), .Z(n22045) );
  XOR U26761 ( .A(n22039), .B(n22038), .Z(n22049) );
  XOR U26762 ( .A(n22041), .B(n22040), .Z(n22038) );
  XOR U26763 ( .A(y[800]), .B(x[800]), .Z(n22040) );
  XOR U26764 ( .A(y[799]), .B(x[799]), .Z(n22041) );
  XOR U26765 ( .A(y[798]), .B(x[798]), .Z(n22039) );
  NAND U26766 ( .A(n22102), .B(n22103), .Z(N28329) );
  NAND U26767 ( .A(n22104), .B(n22105), .Z(n22103) );
  NANDN U26768 ( .A(n22106), .B(n22107), .Z(n22105) );
  NANDN U26769 ( .A(n22107), .B(n22106), .Z(n22102) );
  XOR U26770 ( .A(n22106), .B(n22108), .Z(N28328) );
  XNOR U26771 ( .A(n22104), .B(n22107), .Z(n22108) );
  NAND U26772 ( .A(n22109), .B(n22110), .Z(n22107) );
  NAND U26773 ( .A(n22111), .B(n22112), .Z(n22110) );
  NANDN U26774 ( .A(n22113), .B(n22114), .Z(n22112) );
  NANDN U26775 ( .A(n22114), .B(n22113), .Z(n22109) );
  AND U26776 ( .A(n22115), .B(n22116), .Z(n22104) );
  NAND U26777 ( .A(n22117), .B(n22118), .Z(n22116) );
  OR U26778 ( .A(n22119), .B(n22120), .Z(n22118) );
  NAND U26779 ( .A(n22120), .B(n22119), .Z(n22115) );
  IV U26780 ( .A(n22121), .Z(n22120) );
  AND U26781 ( .A(n22122), .B(n22123), .Z(n22106) );
  NAND U26782 ( .A(n22124), .B(n22125), .Z(n22123) );
  NANDN U26783 ( .A(n22126), .B(n22127), .Z(n22125) );
  NANDN U26784 ( .A(n22127), .B(n22126), .Z(n22122) );
  XOR U26785 ( .A(n22119), .B(n22128), .Z(N28327) );
  XOR U26786 ( .A(n22117), .B(n22121), .Z(n22128) );
  XNOR U26787 ( .A(n22114), .B(n22129), .Z(n22121) );
  XNOR U26788 ( .A(n22111), .B(n22113), .Z(n22129) );
  AND U26789 ( .A(n22130), .B(n22131), .Z(n22113) );
  NANDN U26790 ( .A(n22132), .B(n22133), .Z(n22131) );
  NANDN U26791 ( .A(n22134), .B(n22135), .Z(n22133) );
  IV U26792 ( .A(n22136), .Z(n22135) );
  NAND U26793 ( .A(n22136), .B(n22134), .Z(n22130) );
  AND U26794 ( .A(n22137), .B(n22138), .Z(n22111) );
  NAND U26795 ( .A(n22139), .B(n22140), .Z(n22138) );
  OR U26796 ( .A(n22141), .B(n22142), .Z(n22140) );
  NAND U26797 ( .A(n22142), .B(n22141), .Z(n22137) );
  IV U26798 ( .A(n22143), .Z(n22142) );
  NAND U26799 ( .A(n22144), .B(n22145), .Z(n22114) );
  NANDN U26800 ( .A(n22146), .B(n22147), .Z(n22145) );
  NAND U26801 ( .A(n22148), .B(n22149), .Z(n22147) );
  OR U26802 ( .A(n22149), .B(n22148), .Z(n22144) );
  IV U26803 ( .A(n22150), .Z(n22148) );
  AND U26804 ( .A(n22151), .B(n22152), .Z(n22117) );
  NAND U26805 ( .A(n22153), .B(n22154), .Z(n22152) );
  NANDN U26806 ( .A(n22155), .B(n22156), .Z(n22154) );
  NANDN U26807 ( .A(n22156), .B(n22155), .Z(n22151) );
  XOR U26808 ( .A(n22127), .B(n22157), .Z(n22119) );
  XNOR U26809 ( .A(n22124), .B(n22126), .Z(n22157) );
  AND U26810 ( .A(n22158), .B(n22159), .Z(n22126) );
  NANDN U26811 ( .A(n22160), .B(n22161), .Z(n22159) );
  NANDN U26812 ( .A(n22162), .B(n22163), .Z(n22161) );
  IV U26813 ( .A(n22164), .Z(n22163) );
  NAND U26814 ( .A(n22164), .B(n22162), .Z(n22158) );
  AND U26815 ( .A(n22165), .B(n22166), .Z(n22124) );
  NAND U26816 ( .A(n22167), .B(n22168), .Z(n22166) );
  OR U26817 ( .A(n22169), .B(n22170), .Z(n22168) );
  NAND U26818 ( .A(n22170), .B(n22169), .Z(n22165) );
  IV U26819 ( .A(n22171), .Z(n22170) );
  NAND U26820 ( .A(n22172), .B(n22173), .Z(n22127) );
  NANDN U26821 ( .A(n22174), .B(n22175), .Z(n22173) );
  NAND U26822 ( .A(n22176), .B(n22177), .Z(n22175) );
  OR U26823 ( .A(n22177), .B(n22176), .Z(n22172) );
  IV U26824 ( .A(n22178), .Z(n22176) );
  XOR U26825 ( .A(n22153), .B(n22179), .Z(N28326) );
  XNOR U26826 ( .A(n22156), .B(n22155), .Z(n22179) );
  XNOR U26827 ( .A(n22167), .B(n22180), .Z(n22155) );
  XOR U26828 ( .A(n22171), .B(n22169), .Z(n22180) );
  XOR U26829 ( .A(n22177), .B(n22181), .Z(n22169) );
  XOR U26830 ( .A(n22174), .B(n22178), .Z(n22181) );
  NAND U26831 ( .A(n22182), .B(n22183), .Z(n22178) );
  NAND U26832 ( .A(n22184), .B(n22185), .Z(n22183) );
  NAND U26833 ( .A(n22186), .B(n22187), .Z(n22182) );
  AND U26834 ( .A(n22188), .B(n22189), .Z(n22174) );
  NAND U26835 ( .A(n22190), .B(n22191), .Z(n22189) );
  NAND U26836 ( .A(n22192), .B(n22193), .Z(n22188) );
  NANDN U26837 ( .A(n22194), .B(n22195), .Z(n22177) );
  NANDN U26838 ( .A(n22196), .B(n22197), .Z(n22171) );
  XNOR U26839 ( .A(n22162), .B(n22198), .Z(n22167) );
  XOR U26840 ( .A(n22160), .B(n22164), .Z(n22198) );
  NAND U26841 ( .A(n22199), .B(n22200), .Z(n22164) );
  NAND U26842 ( .A(n22201), .B(n22202), .Z(n22200) );
  NAND U26843 ( .A(n22203), .B(n22204), .Z(n22199) );
  AND U26844 ( .A(n22205), .B(n22206), .Z(n22160) );
  NAND U26845 ( .A(n22207), .B(n22208), .Z(n22206) );
  NAND U26846 ( .A(n22209), .B(n22210), .Z(n22205) );
  AND U26847 ( .A(n22211), .B(n22212), .Z(n22162) );
  NAND U26848 ( .A(n22213), .B(n22214), .Z(n22156) );
  XNOR U26849 ( .A(n22139), .B(n22215), .Z(n22153) );
  XOR U26850 ( .A(n22143), .B(n22141), .Z(n22215) );
  XOR U26851 ( .A(n22149), .B(n22216), .Z(n22141) );
  XOR U26852 ( .A(n22146), .B(n22150), .Z(n22216) );
  NAND U26853 ( .A(n22217), .B(n22218), .Z(n22150) );
  NAND U26854 ( .A(n22219), .B(n22220), .Z(n22218) );
  NAND U26855 ( .A(n22221), .B(n22222), .Z(n22217) );
  AND U26856 ( .A(n22223), .B(n22224), .Z(n22146) );
  NAND U26857 ( .A(n22225), .B(n22226), .Z(n22224) );
  NAND U26858 ( .A(n22227), .B(n22228), .Z(n22223) );
  NANDN U26859 ( .A(n22229), .B(n22230), .Z(n22149) );
  NANDN U26860 ( .A(n22231), .B(n22232), .Z(n22143) );
  XNOR U26861 ( .A(n22134), .B(n22233), .Z(n22139) );
  XOR U26862 ( .A(n22132), .B(n22136), .Z(n22233) );
  NAND U26863 ( .A(n22234), .B(n22235), .Z(n22136) );
  NAND U26864 ( .A(n22236), .B(n22237), .Z(n22235) );
  NAND U26865 ( .A(n22238), .B(n22239), .Z(n22234) );
  AND U26866 ( .A(n22240), .B(n22241), .Z(n22132) );
  NAND U26867 ( .A(n22242), .B(n22243), .Z(n22241) );
  NAND U26868 ( .A(n22244), .B(n22245), .Z(n22240) );
  AND U26869 ( .A(n22246), .B(n22247), .Z(n22134) );
  XOR U26870 ( .A(n22214), .B(n22213), .Z(N28325) );
  XNOR U26871 ( .A(n22232), .B(n22231), .Z(n22213) );
  XNOR U26872 ( .A(n22246), .B(n22247), .Z(n22231) );
  XOR U26873 ( .A(n22243), .B(n22242), .Z(n22247) );
  XOR U26874 ( .A(y[795]), .B(x[795]), .Z(n22242) );
  XOR U26875 ( .A(n22245), .B(n22244), .Z(n22243) );
  XOR U26876 ( .A(y[797]), .B(x[797]), .Z(n22244) );
  XOR U26877 ( .A(y[796]), .B(x[796]), .Z(n22245) );
  XOR U26878 ( .A(n22237), .B(n22236), .Z(n22246) );
  XOR U26879 ( .A(n22239), .B(n22238), .Z(n22236) );
  XOR U26880 ( .A(y[794]), .B(x[794]), .Z(n22238) );
  XOR U26881 ( .A(y[793]), .B(x[793]), .Z(n22239) );
  XOR U26882 ( .A(y[792]), .B(x[792]), .Z(n22237) );
  XNOR U26883 ( .A(n22230), .B(n22229), .Z(n22232) );
  XNOR U26884 ( .A(n22226), .B(n22225), .Z(n22229) );
  XOR U26885 ( .A(n22228), .B(n22227), .Z(n22225) );
  XOR U26886 ( .A(y[791]), .B(x[791]), .Z(n22227) );
  XOR U26887 ( .A(y[790]), .B(x[790]), .Z(n22228) );
  XOR U26888 ( .A(y[789]), .B(x[789]), .Z(n22226) );
  XOR U26889 ( .A(n22220), .B(n22219), .Z(n22230) );
  XOR U26890 ( .A(n22222), .B(n22221), .Z(n22219) );
  XOR U26891 ( .A(y[788]), .B(x[788]), .Z(n22221) );
  XOR U26892 ( .A(y[787]), .B(x[787]), .Z(n22222) );
  XOR U26893 ( .A(y[786]), .B(x[786]), .Z(n22220) );
  XNOR U26894 ( .A(n22197), .B(n22196), .Z(n22214) );
  XNOR U26895 ( .A(n22211), .B(n22212), .Z(n22196) );
  XOR U26896 ( .A(n22208), .B(n22207), .Z(n22212) );
  XOR U26897 ( .A(y[783]), .B(x[783]), .Z(n22207) );
  XOR U26898 ( .A(n22210), .B(n22209), .Z(n22208) );
  XOR U26899 ( .A(y[785]), .B(x[785]), .Z(n22209) );
  XOR U26900 ( .A(y[784]), .B(x[784]), .Z(n22210) );
  XOR U26901 ( .A(n22202), .B(n22201), .Z(n22211) );
  XOR U26902 ( .A(n22204), .B(n22203), .Z(n22201) );
  XOR U26903 ( .A(y[782]), .B(x[782]), .Z(n22203) );
  XOR U26904 ( .A(y[781]), .B(x[781]), .Z(n22204) );
  XOR U26905 ( .A(y[780]), .B(x[780]), .Z(n22202) );
  XNOR U26906 ( .A(n22195), .B(n22194), .Z(n22197) );
  XNOR U26907 ( .A(n22191), .B(n22190), .Z(n22194) );
  XOR U26908 ( .A(n22193), .B(n22192), .Z(n22190) );
  XOR U26909 ( .A(y[779]), .B(x[779]), .Z(n22192) );
  XOR U26910 ( .A(y[778]), .B(x[778]), .Z(n22193) );
  XOR U26911 ( .A(y[777]), .B(x[777]), .Z(n22191) );
  XOR U26912 ( .A(n22185), .B(n22184), .Z(n22195) );
  XOR U26913 ( .A(n22187), .B(n22186), .Z(n22184) );
  XOR U26914 ( .A(y[776]), .B(x[776]), .Z(n22186) );
  XOR U26915 ( .A(y[775]), .B(x[775]), .Z(n22187) );
  XOR U26916 ( .A(y[774]), .B(x[774]), .Z(n22185) );
  NAND U26917 ( .A(n22248), .B(n22249), .Z(N28317) );
  NAND U26918 ( .A(n22250), .B(n22251), .Z(n22249) );
  NANDN U26919 ( .A(n22252), .B(n22253), .Z(n22251) );
  NANDN U26920 ( .A(n22253), .B(n22252), .Z(n22248) );
  XOR U26921 ( .A(n22252), .B(n22254), .Z(N28316) );
  XNOR U26922 ( .A(n22250), .B(n22253), .Z(n22254) );
  NAND U26923 ( .A(n22255), .B(n22256), .Z(n22253) );
  NAND U26924 ( .A(n22257), .B(n22258), .Z(n22256) );
  NANDN U26925 ( .A(n22259), .B(n22260), .Z(n22258) );
  NANDN U26926 ( .A(n22260), .B(n22259), .Z(n22255) );
  AND U26927 ( .A(n22261), .B(n22262), .Z(n22250) );
  NAND U26928 ( .A(n22263), .B(n22264), .Z(n22262) );
  OR U26929 ( .A(n22265), .B(n22266), .Z(n22264) );
  NAND U26930 ( .A(n22266), .B(n22265), .Z(n22261) );
  IV U26931 ( .A(n22267), .Z(n22266) );
  AND U26932 ( .A(n22268), .B(n22269), .Z(n22252) );
  NAND U26933 ( .A(n22270), .B(n22271), .Z(n22269) );
  NANDN U26934 ( .A(n22272), .B(n22273), .Z(n22271) );
  NANDN U26935 ( .A(n22273), .B(n22272), .Z(n22268) );
  XOR U26936 ( .A(n22265), .B(n22274), .Z(N28315) );
  XOR U26937 ( .A(n22263), .B(n22267), .Z(n22274) );
  XNOR U26938 ( .A(n22260), .B(n22275), .Z(n22267) );
  XNOR U26939 ( .A(n22257), .B(n22259), .Z(n22275) );
  AND U26940 ( .A(n22276), .B(n22277), .Z(n22259) );
  NANDN U26941 ( .A(n22278), .B(n22279), .Z(n22277) );
  NANDN U26942 ( .A(n22280), .B(n22281), .Z(n22279) );
  IV U26943 ( .A(n22282), .Z(n22281) );
  NAND U26944 ( .A(n22282), .B(n22280), .Z(n22276) );
  AND U26945 ( .A(n22283), .B(n22284), .Z(n22257) );
  NAND U26946 ( .A(n22285), .B(n22286), .Z(n22284) );
  OR U26947 ( .A(n22287), .B(n22288), .Z(n22286) );
  NAND U26948 ( .A(n22288), .B(n22287), .Z(n22283) );
  IV U26949 ( .A(n22289), .Z(n22288) );
  NAND U26950 ( .A(n22290), .B(n22291), .Z(n22260) );
  NANDN U26951 ( .A(n22292), .B(n22293), .Z(n22291) );
  NAND U26952 ( .A(n22294), .B(n22295), .Z(n22293) );
  OR U26953 ( .A(n22295), .B(n22294), .Z(n22290) );
  IV U26954 ( .A(n22296), .Z(n22294) );
  AND U26955 ( .A(n22297), .B(n22298), .Z(n22263) );
  NAND U26956 ( .A(n22299), .B(n22300), .Z(n22298) );
  NANDN U26957 ( .A(n22301), .B(n22302), .Z(n22300) );
  NANDN U26958 ( .A(n22302), .B(n22301), .Z(n22297) );
  XOR U26959 ( .A(n22273), .B(n22303), .Z(n22265) );
  XNOR U26960 ( .A(n22270), .B(n22272), .Z(n22303) );
  AND U26961 ( .A(n22304), .B(n22305), .Z(n22272) );
  NANDN U26962 ( .A(n22306), .B(n22307), .Z(n22305) );
  NANDN U26963 ( .A(n22308), .B(n22309), .Z(n22307) );
  IV U26964 ( .A(n22310), .Z(n22309) );
  NAND U26965 ( .A(n22310), .B(n22308), .Z(n22304) );
  AND U26966 ( .A(n22311), .B(n22312), .Z(n22270) );
  NAND U26967 ( .A(n22313), .B(n22314), .Z(n22312) );
  OR U26968 ( .A(n22315), .B(n22316), .Z(n22314) );
  NAND U26969 ( .A(n22316), .B(n22315), .Z(n22311) );
  IV U26970 ( .A(n22317), .Z(n22316) );
  NAND U26971 ( .A(n22318), .B(n22319), .Z(n22273) );
  NANDN U26972 ( .A(n22320), .B(n22321), .Z(n22319) );
  NAND U26973 ( .A(n22322), .B(n22323), .Z(n22321) );
  OR U26974 ( .A(n22323), .B(n22322), .Z(n22318) );
  IV U26975 ( .A(n22324), .Z(n22322) );
  XOR U26976 ( .A(n22299), .B(n22325), .Z(N28314) );
  XNOR U26977 ( .A(n22302), .B(n22301), .Z(n22325) );
  XNOR U26978 ( .A(n22313), .B(n22326), .Z(n22301) );
  XOR U26979 ( .A(n22317), .B(n22315), .Z(n22326) );
  XOR U26980 ( .A(n22323), .B(n22327), .Z(n22315) );
  XOR U26981 ( .A(n22320), .B(n22324), .Z(n22327) );
  NAND U26982 ( .A(n22328), .B(n22329), .Z(n22324) );
  NAND U26983 ( .A(n22330), .B(n22331), .Z(n22329) );
  NAND U26984 ( .A(n22332), .B(n22333), .Z(n22328) );
  AND U26985 ( .A(n22334), .B(n22335), .Z(n22320) );
  NAND U26986 ( .A(n22336), .B(n22337), .Z(n22335) );
  NAND U26987 ( .A(n22338), .B(n22339), .Z(n22334) );
  NANDN U26988 ( .A(n22340), .B(n22341), .Z(n22323) );
  NANDN U26989 ( .A(n22342), .B(n22343), .Z(n22317) );
  XNOR U26990 ( .A(n22308), .B(n22344), .Z(n22313) );
  XOR U26991 ( .A(n22306), .B(n22310), .Z(n22344) );
  NAND U26992 ( .A(n22345), .B(n22346), .Z(n22310) );
  NAND U26993 ( .A(n22347), .B(n22348), .Z(n22346) );
  NAND U26994 ( .A(n22349), .B(n22350), .Z(n22345) );
  AND U26995 ( .A(n22351), .B(n22352), .Z(n22306) );
  NAND U26996 ( .A(n22353), .B(n22354), .Z(n22352) );
  NAND U26997 ( .A(n22355), .B(n22356), .Z(n22351) );
  AND U26998 ( .A(n22357), .B(n22358), .Z(n22308) );
  NAND U26999 ( .A(n22359), .B(n22360), .Z(n22302) );
  XNOR U27000 ( .A(n22285), .B(n22361), .Z(n22299) );
  XOR U27001 ( .A(n22289), .B(n22287), .Z(n22361) );
  XOR U27002 ( .A(n22295), .B(n22362), .Z(n22287) );
  XOR U27003 ( .A(n22292), .B(n22296), .Z(n22362) );
  NAND U27004 ( .A(n22363), .B(n22364), .Z(n22296) );
  NAND U27005 ( .A(n22365), .B(n22366), .Z(n22364) );
  NAND U27006 ( .A(n22367), .B(n22368), .Z(n22363) );
  AND U27007 ( .A(n22369), .B(n22370), .Z(n22292) );
  NAND U27008 ( .A(n22371), .B(n22372), .Z(n22370) );
  NAND U27009 ( .A(n22373), .B(n22374), .Z(n22369) );
  NANDN U27010 ( .A(n22375), .B(n22376), .Z(n22295) );
  NANDN U27011 ( .A(n22377), .B(n22378), .Z(n22289) );
  XNOR U27012 ( .A(n22280), .B(n22379), .Z(n22285) );
  XOR U27013 ( .A(n22278), .B(n22282), .Z(n22379) );
  NAND U27014 ( .A(n22380), .B(n22381), .Z(n22282) );
  NAND U27015 ( .A(n22382), .B(n22383), .Z(n22381) );
  NAND U27016 ( .A(n22384), .B(n22385), .Z(n22380) );
  AND U27017 ( .A(n22386), .B(n22387), .Z(n22278) );
  NAND U27018 ( .A(n22388), .B(n22389), .Z(n22387) );
  NAND U27019 ( .A(n22390), .B(n22391), .Z(n22386) );
  AND U27020 ( .A(n22392), .B(n22393), .Z(n22280) );
  XOR U27021 ( .A(n22360), .B(n22359), .Z(N28313) );
  XNOR U27022 ( .A(n22378), .B(n22377), .Z(n22359) );
  XNOR U27023 ( .A(n22392), .B(n22393), .Z(n22377) );
  XOR U27024 ( .A(n22389), .B(n22388), .Z(n22393) );
  XOR U27025 ( .A(y[771]), .B(x[771]), .Z(n22388) );
  XOR U27026 ( .A(n22391), .B(n22390), .Z(n22389) );
  XOR U27027 ( .A(y[773]), .B(x[773]), .Z(n22390) );
  XOR U27028 ( .A(y[772]), .B(x[772]), .Z(n22391) );
  XOR U27029 ( .A(n22383), .B(n22382), .Z(n22392) );
  XOR U27030 ( .A(n22385), .B(n22384), .Z(n22382) );
  XOR U27031 ( .A(y[770]), .B(x[770]), .Z(n22384) );
  XOR U27032 ( .A(y[769]), .B(x[769]), .Z(n22385) );
  XOR U27033 ( .A(y[768]), .B(x[768]), .Z(n22383) );
  XNOR U27034 ( .A(n22376), .B(n22375), .Z(n22378) );
  XNOR U27035 ( .A(n22372), .B(n22371), .Z(n22375) );
  XOR U27036 ( .A(n22374), .B(n22373), .Z(n22371) );
  XOR U27037 ( .A(y[767]), .B(x[767]), .Z(n22373) );
  XOR U27038 ( .A(y[766]), .B(x[766]), .Z(n22374) );
  XOR U27039 ( .A(y[765]), .B(x[765]), .Z(n22372) );
  XOR U27040 ( .A(n22366), .B(n22365), .Z(n22376) );
  XOR U27041 ( .A(n22368), .B(n22367), .Z(n22365) );
  XOR U27042 ( .A(y[764]), .B(x[764]), .Z(n22367) );
  XOR U27043 ( .A(y[763]), .B(x[763]), .Z(n22368) );
  XOR U27044 ( .A(y[762]), .B(x[762]), .Z(n22366) );
  XNOR U27045 ( .A(n22343), .B(n22342), .Z(n22360) );
  XNOR U27046 ( .A(n22357), .B(n22358), .Z(n22342) );
  XOR U27047 ( .A(n22354), .B(n22353), .Z(n22358) );
  XOR U27048 ( .A(y[759]), .B(x[759]), .Z(n22353) );
  XOR U27049 ( .A(n22356), .B(n22355), .Z(n22354) );
  XOR U27050 ( .A(y[761]), .B(x[761]), .Z(n22355) );
  XOR U27051 ( .A(y[760]), .B(x[760]), .Z(n22356) );
  XOR U27052 ( .A(n22348), .B(n22347), .Z(n22357) );
  XOR U27053 ( .A(n22350), .B(n22349), .Z(n22347) );
  XOR U27054 ( .A(y[758]), .B(x[758]), .Z(n22349) );
  XOR U27055 ( .A(y[757]), .B(x[757]), .Z(n22350) );
  XOR U27056 ( .A(y[756]), .B(x[756]), .Z(n22348) );
  XNOR U27057 ( .A(n22341), .B(n22340), .Z(n22343) );
  XNOR U27058 ( .A(n22337), .B(n22336), .Z(n22340) );
  XOR U27059 ( .A(n22339), .B(n22338), .Z(n22336) );
  XOR U27060 ( .A(y[755]), .B(x[755]), .Z(n22338) );
  XOR U27061 ( .A(y[754]), .B(x[754]), .Z(n22339) );
  XOR U27062 ( .A(y[753]), .B(x[753]), .Z(n22337) );
  XOR U27063 ( .A(n22331), .B(n22330), .Z(n22341) );
  XOR U27064 ( .A(n22333), .B(n22332), .Z(n22330) );
  XOR U27065 ( .A(y[752]), .B(x[752]), .Z(n22332) );
  XOR U27066 ( .A(y[751]), .B(x[751]), .Z(n22333) );
  XOR U27067 ( .A(y[750]), .B(x[750]), .Z(n22331) );
  NAND U27068 ( .A(n22394), .B(n22395), .Z(N28305) );
  NAND U27069 ( .A(n22396), .B(n22397), .Z(n22395) );
  NANDN U27070 ( .A(n22398), .B(n22399), .Z(n22397) );
  NANDN U27071 ( .A(n22399), .B(n22398), .Z(n22394) );
  XOR U27072 ( .A(n22398), .B(n22400), .Z(N28304) );
  XNOR U27073 ( .A(n22396), .B(n22399), .Z(n22400) );
  NAND U27074 ( .A(n22401), .B(n22402), .Z(n22399) );
  NAND U27075 ( .A(n22403), .B(n22404), .Z(n22402) );
  NANDN U27076 ( .A(n22405), .B(n22406), .Z(n22404) );
  NANDN U27077 ( .A(n22406), .B(n22405), .Z(n22401) );
  AND U27078 ( .A(n22407), .B(n22408), .Z(n22396) );
  NAND U27079 ( .A(n22409), .B(n22410), .Z(n22408) );
  OR U27080 ( .A(n22411), .B(n22412), .Z(n22410) );
  NAND U27081 ( .A(n22412), .B(n22411), .Z(n22407) );
  IV U27082 ( .A(n22413), .Z(n22412) );
  AND U27083 ( .A(n22414), .B(n22415), .Z(n22398) );
  NAND U27084 ( .A(n22416), .B(n22417), .Z(n22415) );
  NANDN U27085 ( .A(n22418), .B(n22419), .Z(n22417) );
  NANDN U27086 ( .A(n22419), .B(n22418), .Z(n22414) );
  XOR U27087 ( .A(n22411), .B(n22420), .Z(N28303) );
  XOR U27088 ( .A(n22409), .B(n22413), .Z(n22420) );
  XNOR U27089 ( .A(n22406), .B(n22421), .Z(n22413) );
  XNOR U27090 ( .A(n22403), .B(n22405), .Z(n22421) );
  AND U27091 ( .A(n22422), .B(n22423), .Z(n22405) );
  NANDN U27092 ( .A(n22424), .B(n22425), .Z(n22423) );
  NANDN U27093 ( .A(n22426), .B(n22427), .Z(n22425) );
  IV U27094 ( .A(n22428), .Z(n22427) );
  NAND U27095 ( .A(n22428), .B(n22426), .Z(n22422) );
  AND U27096 ( .A(n22429), .B(n22430), .Z(n22403) );
  NAND U27097 ( .A(n22431), .B(n22432), .Z(n22430) );
  OR U27098 ( .A(n22433), .B(n22434), .Z(n22432) );
  NAND U27099 ( .A(n22434), .B(n22433), .Z(n22429) );
  IV U27100 ( .A(n22435), .Z(n22434) );
  NAND U27101 ( .A(n22436), .B(n22437), .Z(n22406) );
  NANDN U27102 ( .A(n22438), .B(n22439), .Z(n22437) );
  NAND U27103 ( .A(n22440), .B(n22441), .Z(n22439) );
  OR U27104 ( .A(n22441), .B(n22440), .Z(n22436) );
  IV U27105 ( .A(n22442), .Z(n22440) );
  AND U27106 ( .A(n22443), .B(n22444), .Z(n22409) );
  NAND U27107 ( .A(n22445), .B(n22446), .Z(n22444) );
  NANDN U27108 ( .A(n22447), .B(n22448), .Z(n22446) );
  NANDN U27109 ( .A(n22448), .B(n22447), .Z(n22443) );
  XOR U27110 ( .A(n22419), .B(n22449), .Z(n22411) );
  XNOR U27111 ( .A(n22416), .B(n22418), .Z(n22449) );
  AND U27112 ( .A(n22450), .B(n22451), .Z(n22418) );
  NANDN U27113 ( .A(n22452), .B(n22453), .Z(n22451) );
  NANDN U27114 ( .A(n22454), .B(n22455), .Z(n22453) );
  IV U27115 ( .A(n22456), .Z(n22455) );
  NAND U27116 ( .A(n22456), .B(n22454), .Z(n22450) );
  AND U27117 ( .A(n22457), .B(n22458), .Z(n22416) );
  NAND U27118 ( .A(n22459), .B(n22460), .Z(n22458) );
  OR U27119 ( .A(n22461), .B(n22462), .Z(n22460) );
  NAND U27120 ( .A(n22462), .B(n22461), .Z(n22457) );
  IV U27121 ( .A(n22463), .Z(n22462) );
  NAND U27122 ( .A(n22464), .B(n22465), .Z(n22419) );
  NANDN U27123 ( .A(n22466), .B(n22467), .Z(n22465) );
  NAND U27124 ( .A(n22468), .B(n22469), .Z(n22467) );
  OR U27125 ( .A(n22469), .B(n22468), .Z(n22464) );
  IV U27126 ( .A(n22470), .Z(n22468) );
  XOR U27127 ( .A(n22445), .B(n22471), .Z(N28302) );
  XNOR U27128 ( .A(n22448), .B(n22447), .Z(n22471) );
  XNOR U27129 ( .A(n22459), .B(n22472), .Z(n22447) );
  XOR U27130 ( .A(n22463), .B(n22461), .Z(n22472) );
  XOR U27131 ( .A(n22469), .B(n22473), .Z(n22461) );
  XOR U27132 ( .A(n22466), .B(n22470), .Z(n22473) );
  NAND U27133 ( .A(n22474), .B(n22475), .Z(n22470) );
  NAND U27134 ( .A(n22476), .B(n22477), .Z(n22475) );
  NAND U27135 ( .A(n22478), .B(n22479), .Z(n22474) );
  AND U27136 ( .A(n22480), .B(n22481), .Z(n22466) );
  NAND U27137 ( .A(n22482), .B(n22483), .Z(n22481) );
  NAND U27138 ( .A(n22484), .B(n22485), .Z(n22480) );
  NANDN U27139 ( .A(n22486), .B(n22487), .Z(n22469) );
  NANDN U27140 ( .A(n22488), .B(n22489), .Z(n22463) );
  XNOR U27141 ( .A(n22454), .B(n22490), .Z(n22459) );
  XOR U27142 ( .A(n22452), .B(n22456), .Z(n22490) );
  NAND U27143 ( .A(n22491), .B(n22492), .Z(n22456) );
  NAND U27144 ( .A(n22493), .B(n22494), .Z(n22492) );
  NAND U27145 ( .A(n22495), .B(n22496), .Z(n22491) );
  AND U27146 ( .A(n22497), .B(n22498), .Z(n22452) );
  NAND U27147 ( .A(n22499), .B(n22500), .Z(n22498) );
  NAND U27148 ( .A(n22501), .B(n22502), .Z(n22497) );
  AND U27149 ( .A(n22503), .B(n22504), .Z(n22454) );
  NAND U27150 ( .A(n22505), .B(n22506), .Z(n22448) );
  XNOR U27151 ( .A(n22431), .B(n22507), .Z(n22445) );
  XOR U27152 ( .A(n22435), .B(n22433), .Z(n22507) );
  XOR U27153 ( .A(n22441), .B(n22508), .Z(n22433) );
  XOR U27154 ( .A(n22438), .B(n22442), .Z(n22508) );
  NAND U27155 ( .A(n22509), .B(n22510), .Z(n22442) );
  NAND U27156 ( .A(n22511), .B(n22512), .Z(n22510) );
  NAND U27157 ( .A(n22513), .B(n22514), .Z(n22509) );
  AND U27158 ( .A(n22515), .B(n22516), .Z(n22438) );
  NAND U27159 ( .A(n22517), .B(n22518), .Z(n22516) );
  NAND U27160 ( .A(n22519), .B(n22520), .Z(n22515) );
  NANDN U27161 ( .A(n22521), .B(n22522), .Z(n22441) );
  NANDN U27162 ( .A(n22523), .B(n22524), .Z(n22435) );
  XNOR U27163 ( .A(n22426), .B(n22525), .Z(n22431) );
  XOR U27164 ( .A(n22424), .B(n22428), .Z(n22525) );
  NAND U27165 ( .A(n22526), .B(n22527), .Z(n22428) );
  NAND U27166 ( .A(n22528), .B(n22529), .Z(n22527) );
  NAND U27167 ( .A(n22530), .B(n22531), .Z(n22526) );
  AND U27168 ( .A(n22532), .B(n22533), .Z(n22424) );
  NAND U27169 ( .A(n22534), .B(n22535), .Z(n22533) );
  NAND U27170 ( .A(n22536), .B(n22537), .Z(n22532) );
  AND U27171 ( .A(n22538), .B(n22539), .Z(n22426) );
  XOR U27172 ( .A(n22506), .B(n22505), .Z(N28301) );
  XNOR U27173 ( .A(n22524), .B(n22523), .Z(n22505) );
  XNOR U27174 ( .A(n22538), .B(n22539), .Z(n22523) );
  XOR U27175 ( .A(n22535), .B(n22534), .Z(n22539) );
  XOR U27176 ( .A(y[747]), .B(x[747]), .Z(n22534) );
  XOR U27177 ( .A(n22537), .B(n22536), .Z(n22535) );
  XOR U27178 ( .A(y[749]), .B(x[749]), .Z(n22536) );
  XOR U27179 ( .A(y[748]), .B(x[748]), .Z(n22537) );
  XOR U27180 ( .A(n22529), .B(n22528), .Z(n22538) );
  XOR U27181 ( .A(n22531), .B(n22530), .Z(n22528) );
  XOR U27182 ( .A(y[746]), .B(x[746]), .Z(n22530) );
  XOR U27183 ( .A(y[745]), .B(x[745]), .Z(n22531) );
  XOR U27184 ( .A(y[744]), .B(x[744]), .Z(n22529) );
  XNOR U27185 ( .A(n22522), .B(n22521), .Z(n22524) );
  XNOR U27186 ( .A(n22518), .B(n22517), .Z(n22521) );
  XOR U27187 ( .A(n22520), .B(n22519), .Z(n22517) );
  XOR U27188 ( .A(y[743]), .B(x[743]), .Z(n22519) );
  XOR U27189 ( .A(y[742]), .B(x[742]), .Z(n22520) );
  XOR U27190 ( .A(y[741]), .B(x[741]), .Z(n22518) );
  XOR U27191 ( .A(n22512), .B(n22511), .Z(n22522) );
  XOR U27192 ( .A(n22514), .B(n22513), .Z(n22511) );
  XOR U27193 ( .A(y[740]), .B(x[740]), .Z(n22513) );
  XOR U27194 ( .A(y[739]), .B(x[739]), .Z(n22514) );
  XOR U27195 ( .A(y[738]), .B(x[738]), .Z(n22512) );
  XNOR U27196 ( .A(n22489), .B(n22488), .Z(n22506) );
  XNOR U27197 ( .A(n22503), .B(n22504), .Z(n22488) );
  XOR U27198 ( .A(n22500), .B(n22499), .Z(n22504) );
  XOR U27199 ( .A(y[735]), .B(x[735]), .Z(n22499) );
  XOR U27200 ( .A(n22502), .B(n22501), .Z(n22500) );
  XOR U27201 ( .A(y[737]), .B(x[737]), .Z(n22501) );
  XOR U27202 ( .A(y[736]), .B(x[736]), .Z(n22502) );
  XOR U27203 ( .A(n22494), .B(n22493), .Z(n22503) );
  XOR U27204 ( .A(n22496), .B(n22495), .Z(n22493) );
  XOR U27205 ( .A(y[734]), .B(x[734]), .Z(n22495) );
  XOR U27206 ( .A(y[733]), .B(x[733]), .Z(n22496) );
  XOR U27207 ( .A(y[732]), .B(x[732]), .Z(n22494) );
  XNOR U27208 ( .A(n22487), .B(n22486), .Z(n22489) );
  XNOR U27209 ( .A(n22483), .B(n22482), .Z(n22486) );
  XOR U27210 ( .A(n22485), .B(n22484), .Z(n22482) );
  XOR U27211 ( .A(y[731]), .B(x[731]), .Z(n22484) );
  XOR U27212 ( .A(y[730]), .B(x[730]), .Z(n22485) );
  XOR U27213 ( .A(y[729]), .B(x[729]), .Z(n22483) );
  XOR U27214 ( .A(n22477), .B(n22476), .Z(n22487) );
  XOR U27215 ( .A(n22479), .B(n22478), .Z(n22476) );
  XOR U27216 ( .A(y[728]), .B(x[728]), .Z(n22478) );
  XOR U27217 ( .A(y[727]), .B(x[727]), .Z(n22479) );
  XOR U27218 ( .A(y[726]), .B(x[726]), .Z(n22477) );
  NAND U27219 ( .A(n22540), .B(n22541), .Z(N28293) );
  NAND U27220 ( .A(n22542), .B(n22543), .Z(n22541) );
  NANDN U27221 ( .A(n22544), .B(n22545), .Z(n22543) );
  NANDN U27222 ( .A(n22545), .B(n22544), .Z(n22540) );
  XOR U27223 ( .A(n22544), .B(n22546), .Z(N28292) );
  XNOR U27224 ( .A(n22542), .B(n22545), .Z(n22546) );
  NAND U27225 ( .A(n22547), .B(n22548), .Z(n22545) );
  NAND U27226 ( .A(n22549), .B(n22550), .Z(n22548) );
  NANDN U27227 ( .A(n22551), .B(n22552), .Z(n22550) );
  NANDN U27228 ( .A(n22552), .B(n22551), .Z(n22547) );
  AND U27229 ( .A(n22553), .B(n22554), .Z(n22542) );
  NAND U27230 ( .A(n22555), .B(n22556), .Z(n22554) );
  OR U27231 ( .A(n22557), .B(n22558), .Z(n22556) );
  NAND U27232 ( .A(n22558), .B(n22557), .Z(n22553) );
  IV U27233 ( .A(n22559), .Z(n22558) );
  AND U27234 ( .A(n22560), .B(n22561), .Z(n22544) );
  NAND U27235 ( .A(n22562), .B(n22563), .Z(n22561) );
  NANDN U27236 ( .A(n22564), .B(n22565), .Z(n22563) );
  NANDN U27237 ( .A(n22565), .B(n22564), .Z(n22560) );
  XOR U27238 ( .A(n22557), .B(n22566), .Z(N28291) );
  XOR U27239 ( .A(n22555), .B(n22559), .Z(n22566) );
  XNOR U27240 ( .A(n22552), .B(n22567), .Z(n22559) );
  XNOR U27241 ( .A(n22549), .B(n22551), .Z(n22567) );
  AND U27242 ( .A(n22568), .B(n22569), .Z(n22551) );
  NANDN U27243 ( .A(n22570), .B(n22571), .Z(n22569) );
  NANDN U27244 ( .A(n22572), .B(n22573), .Z(n22571) );
  IV U27245 ( .A(n22574), .Z(n22573) );
  NAND U27246 ( .A(n22574), .B(n22572), .Z(n22568) );
  AND U27247 ( .A(n22575), .B(n22576), .Z(n22549) );
  NAND U27248 ( .A(n22577), .B(n22578), .Z(n22576) );
  OR U27249 ( .A(n22579), .B(n22580), .Z(n22578) );
  NAND U27250 ( .A(n22580), .B(n22579), .Z(n22575) );
  IV U27251 ( .A(n22581), .Z(n22580) );
  NAND U27252 ( .A(n22582), .B(n22583), .Z(n22552) );
  NANDN U27253 ( .A(n22584), .B(n22585), .Z(n22583) );
  NAND U27254 ( .A(n22586), .B(n22587), .Z(n22585) );
  OR U27255 ( .A(n22587), .B(n22586), .Z(n22582) );
  IV U27256 ( .A(n22588), .Z(n22586) );
  AND U27257 ( .A(n22589), .B(n22590), .Z(n22555) );
  NAND U27258 ( .A(n22591), .B(n22592), .Z(n22590) );
  NANDN U27259 ( .A(n22593), .B(n22594), .Z(n22592) );
  NANDN U27260 ( .A(n22594), .B(n22593), .Z(n22589) );
  XOR U27261 ( .A(n22565), .B(n22595), .Z(n22557) );
  XNOR U27262 ( .A(n22562), .B(n22564), .Z(n22595) );
  AND U27263 ( .A(n22596), .B(n22597), .Z(n22564) );
  NANDN U27264 ( .A(n22598), .B(n22599), .Z(n22597) );
  NANDN U27265 ( .A(n22600), .B(n22601), .Z(n22599) );
  IV U27266 ( .A(n22602), .Z(n22601) );
  NAND U27267 ( .A(n22602), .B(n22600), .Z(n22596) );
  AND U27268 ( .A(n22603), .B(n22604), .Z(n22562) );
  NAND U27269 ( .A(n22605), .B(n22606), .Z(n22604) );
  OR U27270 ( .A(n22607), .B(n22608), .Z(n22606) );
  NAND U27271 ( .A(n22608), .B(n22607), .Z(n22603) );
  IV U27272 ( .A(n22609), .Z(n22608) );
  NAND U27273 ( .A(n22610), .B(n22611), .Z(n22565) );
  NANDN U27274 ( .A(n22612), .B(n22613), .Z(n22611) );
  NAND U27275 ( .A(n22614), .B(n22615), .Z(n22613) );
  OR U27276 ( .A(n22615), .B(n22614), .Z(n22610) );
  IV U27277 ( .A(n22616), .Z(n22614) );
  XOR U27278 ( .A(n22591), .B(n22617), .Z(N28290) );
  XNOR U27279 ( .A(n22594), .B(n22593), .Z(n22617) );
  XNOR U27280 ( .A(n22605), .B(n22618), .Z(n22593) );
  XOR U27281 ( .A(n22609), .B(n22607), .Z(n22618) );
  XOR U27282 ( .A(n22615), .B(n22619), .Z(n22607) );
  XOR U27283 ( .A(n22612), .B(n22616), .Z(n22619) );
  NAND U27284 ( .A(n22620), .B(n22621), .Z(n22616) );
  NAND U27285 ( .A(n22622), .B(n22623), .Z(n22621) );
  NAND U27286 ( .A(n22624), .B(n22625), .Z(n22620) );
  AND U27287 ( .A(n22626), .B(n22627), .Z(n22612) );
  NAND U27288 ( .A(n22628), .B(n22629), .Z(n22627) );
  NAND U27289 ( .A(n22630), .B(n22631), .Z(n22626) );
  NANDN U27290 ( .A(n22632), .B(n22633), .Z(n22615) );
  NANDN U27291 ( .A(n22634), .B(n22635), .Z(n22609) );
  XNOR U27292 ( .A(n22600), .B(n22636), .Z(n22605) );
  XOR U27293 ( .A(n22598), .B(n22602), .Z(n22636) );
  NAND U27294 ( .A(n22637), .B(n22638), .Z(n22602) );
  NAND U27295 ( .A(n22639), .B(n22640), .Z(n22638) );
  NAND U27296 ( .A(n22641), .B(n22642), .Z(n22637) );
  AND U27297 ( .A(n22643), .B(n22644), .Z(n22598) );
  NAND U27298 ( .A(n22645), .B(n22646), .Z(n22644) );
  NAND U27299 ( .A(n22647), .B(n22648), .Z(n22643) );
  AND U27300 ( .A(n22649), .B(n22650), .Z(n22600) );
  NAND U27301 ( .A(n22651), .B(n22652), .Z(n22594) );
  XNOR U27302 ( .A(n22577), .B(n22653), .Z(n22591) );
  XOR U27303 ( .A(n22581), .B(n22579), .Z(n22653) );
  XOR U27304 ( .A(n22587), .B(n22654), .Z(n22579) );
  XOR U27305 ( .A(n22584), .B(n22588), .Z(n22654) );
  NAND U27306 ( .A(n22655), .B(n22656), .Z(n22588) );
  NAND U27307 ( .A(n22657), .B(n22658), .Z(n22656) );
  NAND U27308 ( .A(n22659), .B(n22660), .Z(n22655) );
  AND U27309 ( .A(n22661), .B(n22662), .Z(n22584) );
  NAND U27310 ( .A(n22663), .B(n22664), .Z(n22662) );
  NAND U27311 ( .A(n22665), .B(n22666), .Z(n22661) );
  NANDN U27312 ( .A(n22667), .B(n22668), .Z(n22587) );
  NANDN U27313 ( .A(n22669), .B(n22670), .Z(n22581) );
  XNOR U27314 ( .A(n22572), .B(n22671), .Z(n22577) );
  XOR U27315 ( .A(n22570), .B(n22574), .Z(n22671) );
  NAND U27316 ( .A(n22672), .B(n22673), .Z(n22574) );
  NAND U27317 ( .A(n22674), .B(n22675), .Z(n22673) );
  NAND U27318 ( .A(n22676), .B(n22677), .Z(n22672) );
  AND U27319 ( .A(n22678), .B(n22679), .Z(n22570) );
  NAND U27320 ( .A(n22680), .B(n22681), .Z(n22679) );
  NAND U27321 ( .A(n22682), .B(n22683), .Z(n22678) );
  AND U27322 ( .A(n22684), .B(n22685), .Z(n22572) );
  XOR U27323 ( .A(n22652), .B(n22651), .Z(N28289) );
  XNOR U27324 ( .A(n22670), .B(n22669), .Z(n22651) );
  XNOR U27325 ( .A(n22684), .B(n22685), .Z(n22669) );
  XOR U27326 ( .A(n22681), .B(n22680), .Z(n22685) );
  XOR U27327 ( .A(y[723]), .B(x[723]), .Z(n22680) );
  XOR U27328 ( .A(n22683), .B(n22682), .Z(n22681) );
  XOR U27329 ( .A(y[725]), .B(x[725]), .Z(n22682) );
  XOR U27330 ( .A(y[724]), .B(x[724]), .Z(n22683) );
  XOR U27331 ( .A(n22675), .B(n22674), .Z(n22684) );
  XOR U27332 ( .A(n22677), .B(n22676), .Z(n22674) );
  XOR U27333 ( .A(y[722]), .B(x[722]), .Z(n22676) );
  XOR U27334 ( .A(y[721]), .B(x[721]), .Z(n22677) );
  XOR U27335 ( .A(y[720]), .B(x[720]), .Z(n22675) );
  XNOR U27336 ( .A(n22668), .B(n22667), .Z(n22670) );
  XNOR U27337 ( .A(n22664), .B(n22663), .Z(n22667) );
  XOR U27338 ( .A(n22666), .B(n22665), .Z(n22663) );
  XOR U27339 ( .A(y[719]), .B(x[719]), .Z(n22665) );
  XOR U27340 ( .A(y[718]), .B(x[718]), .Z(n22666) );
  XOR U27341 ( .A(y[717]), .B(x[717]), .Z(n22664) );
  XOR U27342 ( .A(n22658), .B(n22657), .Z(n22668) );
  XOR U27343 ( .A(n22660), .B(n22659), .Z(n22657) );
  XOR U27344 ( .A(y[716]), .B(x[716]), .Z(n22659) );
  XOR U27345 ( .A(y[715]), .B(x[715]), .Z(n22660) );
  XOR U27346 ( .A(y[714]), .B(x[714]), .Z(n22658) );
  XNOR U27347 ( .A(n22635), .B(n22634), .Z(n22652) );
  XNOR U27348 ( .A(n22649), .B(n22650), .Z(n22634) );
  XOR U27349 ( .A(n22646), .B(n22645), .Z(n22650) );
  XOR U27350 ( .A(y[711]), .B(x[711]), .Z(n22645) );
  XOR U27351 ( .A(n22648), .B(n22647), .Z(n22646) );
  XOR U27352 ( .A(y[713]), .B(x[713]), .Z(n22647) );
  XOR U27353 ( .A(y[712]), .B(x[712]), .Z(n22648) );
  XOR U27354 ( .A(n22640), .B(n22639), .Z(n22649) );
  XOR U27355 ( .A(n22642), .B(n22641), .Z(n22639) );
  XOR U27356 ( .A(y[710]), .B(x[710]), .Z(n22641) );
  XOR U27357 ( .A(y[709]), .B(x[709]), .Z(n22642) );
  XOR U27358 ( .A(y[708]), .B(x[708]), .Z(n22640) );
  XNOR U27359 ( .A(n22633), .B(n22632), .Z(n22635) );
  XNOR U27360 ( .A(n22629), .B(n22628), .Z(n22632) );
  XOR U27361 ( .A(n22631), .B(n22630), .Z(n22628) );
  XOR U27362 ( .A(y[707]), .B(x[707]), .Z(n22630) );
  XOR U27363 ( .A(y[706]), .B(x[706]), .Z(n22631) );
  XOR U27364 ( .A(y[705]), .B(x[705]), .Z(n22629) );
  XOR U27365 ( .A(n22623), .B(n22622), .Z(n22633) );
  XOR U27366 ( .A(n22625), .B(n22624), .Z(n22622) );
  XOR U27367 ( .A(y[704]), .B(x[704]), .Z(n22624) );
  XOR U27368 ( .A(y[703]), .B(x[703]), .Z(n22625) );
  XOR U27369 ( .A(y[702]), .B(x[702]), .Z(n22623) );
  NAND U27370 ( .A(n22686), .B(n22687), .Z(N28281) );
  NAND U27371 ( .A(n22688), .B(n22689), .Z(n22687) );
  NANDN U27372 ( .A(n22690), .B(n22691), .Z(n22689) );
  NANDN U27373 ( .A(n22691), .B(n22690), .Z(n22686) );
  XOR U27374 ( .A(n22690), .B(n22692), .Z(N28280) );
  XNOR U27375 ( .A(n22688), .B(n22691), .Z(n22692) );
  NAND U27376 ( .A(n22693), .B(n22694), .Z(n22691) );
  NAND U27377 ( .A(n22695), .B(n22696), .Z(n22694) );
  NANDN U27378 ( .A(n22697), .B(n22698), .Z(n22696) );
  NANDN U27379 ( .A(n22698), .B(n22697), .Z(n22693) );
  AND U27380 ( .A(n22699), .B(n22700), .Z(n22688) );
  NAND U27381 ( .A(n22701), .B(n22702), .Z(n22700) );
  OR U27382 ( .A(n22703), .B(n22704), .Z(n22702) );
  NAND U27383 ( .A(n22704), .B(n22703), .Z(n22699) );
  IV U27384 ( .A(n22705), .Z(n22704) );
  AND U27385 ( .A(n22706), .B(n22707), .Z(n22690) );
  NAND U27386 ( .A(n22708), .B(n22709), .Z(n22707) );
  NANDN U27387 ( .A(n22710), .B(n22711), .Z(n22709) );
  NANDN U27388 ( .A(n22711), .B(n22710), .Z(n22706) );
  XOR U27389 ( .A(n22703), .B(n22712), .Z(N28279) );
  XOR U27390 ( .A(n22701), .B(n22705), .Z(n22712) );
  XNOR U27391 ( .A(n22698), .B(n22713), .Z(n22705) );
  XNOR U27392 ( .A(n22695), .B(n22697), .Z(n22713) );
  AND U27393 ( .A(n22714), .B(n22715), .Z(n22697) );
  NANDN U27394 ( .A(n22716), .B(n22717), .Z(n22715) );
  NANDN U27395 ( .A(n22718), .B(n22719), .Z(n22717) );
  IV U27396 ( .A(n22720), .Z(n22719) );
  NAND U27397 ( .A(n22720), .B(n22718), .Z(n22714) );
  AND U27398 ( .A(n22721), .B(n22722), .Z(n22695) );
  NAND U27399 ( .A(n22723), .B(n22724), .Z(n22722) );
  OR U27400 ( .A(n22725), .B(n22726), .Z(n22724) );
  NAND U27401 ( .A(n22726), .B(n22725), .Z(n22721) );
  IV U27402 ( .A(n22727), .Z(n22726) );
  NAND U27403 ( .A(n22728), .B(n22729), .Z(n22698) );
  NANDN U27404 ( .A(n22730), .B(n22731), .Z(n22729) );
  NAND U27405 ( .A(n22732), .B(n22733), .Z(n22731) );
  OR U27406 ( .A(n22733), .B(n22732), .Z(n22728) );
  IV U27407 ( .A(n22734), .Z(n22732) );
  AND U27408 ( .A(n22735), .B(n22736), .Z(n22701) );
  NAND U27409 ( .A(n22737), .B(n22738), .Z(n22736) );
  NANDN U27410 ( .A(n22739), .B(n22740), .Z(n22738) );
  NANDN U27411 ( .A(n22740), .B(n22739), .Z(n22735) );
  XOR U27412 ( .A(n22711), .B(n22741), .Z(n22703) );
  XNOR U27413 ( .A(n22708), .B(n22710), .Z(n22741) );
  AND U27414 ( .A(n22742), .B(n22743), .Z(n22710) );
  NANDN U27415 ( .A(n22744), .B(n22745), .Z(n22743) );
  NANDN U27416 ( .A(n22746), .B(n22747), .Z(n22745) );
  IV U27417 ( .A(n22748), .Z(n22747) );
  NAND U27418 ( .A(n22748), .B(n22746), .Z(n22742) );
  AND U27419 ( .A(n22749), .B(n22750), .Z(n22708) );
  NAND U27420 ( .A(n22751), .B(n22752), .Z(n22750) );
  OR U27421 ( .A(n22753), .B(n22754), .Z(n22752) );
  NAND U27422 ( .A(n22754), .B(n22753), .Z(n22749) );
  IV U27423 ( .A(n22755), .Z(n22754) );
  NAND U27424 ( .A(n22756), .B(n22757), .Z(n22711) );
  NANDN U27425 ( .A(n22758), .B(n22759), .Z(n22757) );
  NAND U27426 ( .A(n22760), .B(n22761), .Z(n22759) );
  OR U27427 ( .A(n22761), .B(n22760), .Z(n22756) );
  IV U27428 ( .A(n22762), .Z(n22760) );
  XOR U27429 ( .A(n22737), .B(n22763), .Z(N28278) );
  XNOR U27430 ( .A(n22740), .B(n22739), .Z(n22763) );
  XNOR U27431 ( .A(n22751), .B(n22764), .Z(n22739) );
  XOR U27432 ( .A(n22755), .B(n22753), .Z(n22764) );
  XOR U27433 ( .A(n22761), .B(n22765), .Z(n22753) );
  XOR U27434 ( .A(n22758), .B(n22762), .Z(n22765) );
  NAND U27435 ( .A(n22766), .B(n22767), .Z(n22762) );
  NAND U27436 ( .A(n22768), .B(n22769), .Z(n22767) );
  NAND U27437 ( .A(n22770), .B(n22771), .Z(n22766) );
  AND U27438 ( .A(n22772), .B(n22773), .Z(n22758) );
  NAND U27439 ( .A(n22774), .B(n22775), .Z(n22773) );
  NAND U27440 ( .A(n22776), .B(n22777), .Z(n22772) );
  NANDN U27441 ( .A(n22778), .B(n22779), .Z(n22761) );
  NANDN U27442 ( .A(n22780), .B(n22781), .Z(n22755) );
  XNOR U27443 ( .A(n22746), .B(n22782), .Z(n22751) );
  XOR U27444 ( .A(n22744), .B(n22748), .Z(n22782) );
  NAND U27445 ( .A(n22783), .B(n22784), .Z(n22748) );
  NAND U27446 ( .A(n22785), .B(n22786), .Z(n22784) );
  NAND U27447 ( .A(n22787), .B(n22788), .Z(n22783) );
  AND U27448 ( .A(n22789), .B(n22790), .Z(n22744) );
  NAND U27449 ( .A(n22791), .B(n22792), .Z(n22790) );
  NAND U27450 ( .A(n22793), .B(n22794), .Z(n22789) );
  AND U27451 ( .A(n22795), .B(n22796), .Z(n22746) );
  NAND U27452 ( .A(n22797), .B(n22798), .Z(n22740) );
  XNOR U27453 ( .A(n22723), .B(n22799), .Z(n22737) );
  XOR U27454 ( .A(n22727), .B(n22725), .Z(n22799) );
  XOR U27455 ( .A(n22733), .B(n22800), .Z(n22725) );
  XOR U27456 ( .A(n22730), .B(n22734), .Z(n22800) );
  NAND U27457 ( .A(n22801), .B(n22802), .Z(n22734) );
  NAND U27458 ( .A(n22803), .B(n22804), .Z(n22802) );
  NAND U27459 ( .A(n22805), .B(n22806), .Z(n22801) );
  AND U27460 ( .A(n22807), .B(n22808), .Z(n22730) );
  NAND U27461 ( .A(n22809), .B(n22810), .Z(n22808) );
  NAND U27462 ( .A(n22811), .B(n22812), .Z(n22807) );
  NANDN U27463 ( .A(n22813), .B(n22814), .Z(n22733) );
  NANDN U27464 ( .A(n22815), .B(n22816), .Z(n22727) );
  XNOR U27465 ( .A(n22718), .B(n22817), .Z(n22723) );
  XOR U27466 ( .A(n22716), .B(n22720), .Z(n22817) );
  NAND U27467 ( .A(n22818), .B(n22819), .Z(n22720) );
  NAND U27468 ( .A(n22820), .B(n22821), .Z(n22819) );
  NAND U27469 ( .A(n22822), .B(n22823), .Z(n22818) );
  AND U27470 ( .A(n22824), .B(n22825), .Z(n22716) );
  NAND U27471 ( .A(n22826), .B(n22827), .Z(n22825) );
  NAND U27472 ( .A(n22828), .B(n22829), .Z(n22824) );
  AND U27473 ( .A(n22830), .B(n22831), .Z(n22718) );
  XOR U27474 ( .A(n22798), .B(n22797), .Z(N28277) );
  XNOR U27475 ( .A(n22816), .B(n22815), .Z(n22797) );
  XNOR U27476 ( .A(n22830), .B(n22831), .Z(n22815) );
  XOR U27477 ( .A(n22827), .B(n22826), .Z(n22831) );
  XOR U27478 ( .A(y[699]), .B(x[699]), .Z(n22826) );
  XOR U27479 ( .A(n22829), .B(n22828), .Z(n22827) );
  XOR U27480 ( .A(y[701]), .B(x[701]), .Z(n22828) );
  XOR U27481 ( .A(y[700]), .B(x[700]), .Z(n22829) );
  XOR U27482 ( .A(n22821), .B(n22820), .Z(n22830) );
  XOR U27483 ( .A(n22823), .B(n22822), .Z(n22820) );
  XOR U27484 ( .A(y[698]), .B(x[698]), .Z(n22822) );
  XOR U27485 ( .A(y[697]), .B(x[697]), .Z(n22823) );
  XOR U27486 ( .A(y[696]), .B(x[696]), .Z(n22821) );
  XNOR U27487 ( .A(n22814), .B(n22813), .Z(n22816) );
  XNOR U27488 ( .A(n22810), .B(n22809), .Z(n22813) );
  XOR U27489 ( .A(n22812), .B(n22811), .Z(n22809) );
  XOR U27490 ( .A(y[695]), .B(x[695]), .Z(n22811) );
  XOR U27491 ( .A(y[694]), .B(x[694]), .Z(n22812) );
  XOR U27492 ( .A(y[693]), .B(x[693]), .Z(n22810) );
  XOR U27493 ( .A(n22804), .B(n22803), .Z(n22814) );
  XOR U27494 ( .A(n22806), .B(n22805), .Z(n22803) );
  XOR U27495 ( .A(y[692]), .B(x[692]), .Z(n22805) );
  XOR U27496 ( .A(y[691]), .B(x[691]), .Z(n22806) );
  XOR U27497 ( .A(y[690]), .B(x[690]), .Z(n22804) );
  XNOR U27498 ( .A(n22781), .B(n22780), .Z(n22798) );
  XNOR U27499 ( .A(n22795), .B(n22796), .Z(n22780) );
  XOR U27500 ( .A(n22792), .B(n22791), .Z(n22796) );
  XOR U27501 ( .A(y[687]), .B(x[687]), .Z(n22791) );
  XOR U27502 ( .A(n22794), .B(n22793), .Z(n22792) );
  XOR U27503 ( .A(y[689]), .B(x[689]), .Z(n22793) );
  XOR U27504 ( .A(y[688]), .B(x[688]), .Z(n22794) );
  XOR U27505 ( .A(n22786), .B(n22785), .Z(n22795) );
  XOR U27506 ( .A(n22788), .B(n22787), .Z(n22785) );
  XOR U27507 ( .A(y[686]), .B(x[686]), .Z(n22787) );
  XOR U27508 ( .A(y[685]), .B(x[685]), .Z(n22788) );
  XOR U27509 ( .A(y[684]), .B(x[684]), .Z(n22786) );
  XNOR U27510 ( .A(n22779), .B(n22778), .Z(n22781) );
  XNOR U27511 ( .A(n22775), .B(n22774), .Z(n22778) );
  XOR U27512 ( .A(n22777), .B(n22776), .Z(n22774) );
  XOR U27513 ( .A(y[683]), .B(x[683]), .Z(n22776) );
  XOR U27514 ( .A(y[682]), .B(x[682]), .Z(n22777) );
  XOR U27515 ( .A(y[681]), .B(x[681]), .Z(n22775) );
  XOR U27516 ( .A(n22769), .B(n22768), .Z(n22779) );
  XOR U27517 ( .A(n22771), .B(n22770), .Z(n22768) );
  XOR U27518 ( .A(y[680]), .B(x[680]), .Z(n22770) );
  XOR U27519 ( .A(y[679]), .B(x[679]), .Z(n22771) );
  XOR U27520 ( .A(y[678]), .B(x[678]), .Z(n22769) );
  NAND U27521 ( .A(n22832), .B(n22833), .Z(N28269) );
  NAND U27522 ( .A(n22834), .B(n22835), .Z(n22833) );
  NANDN U27523 ( .A(n22836), .B(n22837), .Z(n22835) );
  NANDN U27524 ( .A(n22837), .B(n22836), .Z(n22832) );
  XOR U27525 ( .A(n22836), .B(n22838), .Z(N28268) );
  XNOR U27526 ( .A(n22834), .B(n22837), .Z(n22838) );
  NAND U27527 ( .A(n22839), .B(n22840), .Z(n22837) );
  NAND U27528 ( .A(n22841), .B(n22842), .Z(n22840) );
  NANDN U27529 ( .A(n22843), .B(n22844), .Z(n22842) );
  NANDN U27530 ( .A(n22844), .B(n22843), .Z(n22839) );
  AND U27531 ( .A(n22845), .B(n22846), .Z(n22834) );
  NAND U27532 ( .A(n22847), .B(n22848), .Z(n22846) );
  OR U27533 ( .A(n22849), .B(n22850), .Z(n22848) );
  NAND U27534 ( .A(n22850), .B(n22849), .Z(n22845) );
  IV U27535 ( .A(n22851), .Z(n22850) );
  AND U27536 ( .A(n22852), .B(n22853), .Z(n22836) );
  NAND U27537 ( .A(n22854), .B(n22855), .Z(n22853) );
  NANDN U27538 ( .A(n22856), .B(n22857), .Z(n22855) );
  NANDN U27539 ( .A(n22857), .B(n22856), .Z(n22852) );
  XOR U27540 ( .A(n22849), .B(n22858), .Z(N28267) );
  XOR U27541 ( .A(n22847), .B(n22851), .Z(n22858) );
  XNOR U27542 ( .A(n22844), .B(n22859), .Z(n22851) );
  XNOR U27543 ( .A(n22841), .B(n22843), .Z(n22859) );
  AND U27544 ( .A(n22860), .B(n22861), .Z(n22843) );
  NANDN U27545 ( .A(n22862), .B(n22863), .Z(n22861) );
  NANDN U27546 ( .A(n22864), .B(n22865), .Z(n22863) );
  IV U27547 ( .A(n22866), .Z(n22865) );
  NAND U27548 ( .A(n22866), .B(n22864), .Z(n22860) );
  AND U27549 ( .A(n22867), .B(n22868), .Z(n22841) );
  NAND U27550 ( .A(n22869), .B(n22870), .Z(n22868) );
  OR U27551 ( .A(n22871), .B(n22872), .Z(n22870) );
  NAND U27552 ( .A(n22872), .B(n22871), .Z(n22867) );
  IV U27553 ( .A(n22873), .Z(n22872) );
  NAND U27554 ( .A(n22874), .B(n22875), .Z(n22844) );
  NANDN U27555 ( .A(n22876), .B(n22877), .Z(n22875) );
  NAND U27556 ( .A(n22878), .B(n22879), .Z(n22877) );
  OR U27557 ( .A(n22879), .B(n22878), .Z(n22874) );
  IV U27558 ( .A(n22880), .Z(n22878) );
  AND U27559 ( .A(n22881), .B(n22882), .Z(n22847) );
  NAND U27560 ( .A(n22883), .B(n22884), .Z(n22882) );
  NANDN U27561 ( .A(n22885), .B(n22886), .Z(n22884) );
  NANDN U27562 ( .A(n22886), .B(n22885), .Z(n22881) );
  XOR U27563 ( .A(n22857), .B(n22887), .Z(n22849) );
  XNOR U27564 ( .A(n22854), .B(n22856), .Z(n22887) );
  AND U27565 ( .A(n22888), .B(n22889), .Z(n22856) );
  NANDN U27566 ( .A(n22890), .B(n22891), .Z(n22889) );
  NANDN U27567 ( .A(n22892), .B(n22893), .Z(n22891) );
  IV U27568 ( .A(n22894), .Z(n22893) );
  NAND U27569 ( .A(n22894), .B(n22892), .Z(n22888) );
  AND U27570 ( .A(n22895), .B(n22896), .Z(n22854) );
  NAND U27571 ( .A(n22897), .B(n22898), .Z(n22896) );
  OR U27572 ( .A(n22899), .B(n22900), .Z(n22898) );
  NAND U27573 ( .A(n22900), .B(n22899), .Z(n22895) );
  IV U27574 ( .A(n22901), .Z(n22900) );
  NAND U27575 ( .A(n22902), .B(n22903), .Z(n22857) );
  NANDN U27576 ( .A(n22904), .B(n22905), .Z(n22903) );
  NAND U27577 ( .A(n22906), .B(n22907), .Z(n22905) );
  OR U27578 ( .A(n22907), .B(n22906), .Z(n22902) );
  IV U27579 ( .A(n22908), .Z(n22906) );
  XOR U27580 ( .A(n22883), .B(n22909), .Z(N28266) );
  XNOR U27581 ( .A(n22886), .B(n22885), .Z(n22909) );
  XNOR U27582 ( .A(n22897), .B(n22910), .Z(n22885) );
  XOR U27583 ( .A(n22901), .B(n22899), .Z(n22910) );
  XOR U27584 ( .A(n22907), .B(n22911), .Z(n22899) );
  XOR U27585 ( .A(n22904), .B(n22908), .Z(n22911) );
  NAND U27586 ( .A(n22912), .B(n22913), .Z(n22908) );
  NAND U27587 ( .A(n22914), .B(n22915), .Z(n22913) );
  NAND U27588 ( .A(n22916), .B(n22917), .Z(n22912) );
  AND U27589 ( .A(n22918), .B(n22919), .Z(n22904) );
  NAND U27590 ( .A(n22920), .B(n22921), .Z(n22919) );
  NAND U27591 ( .A(n22922), .B(n22923), .Z(n22918) );
  NANDN U27592 ( .A(n22924), .B(n22925), .Z(n22907) );
  NANDN U27593 ( .A(n22926), .B(n22927), .Z(n22901) );
  XNOR U27594 ( .A(n22892), .B(n22928), .Z(n22897) );
  XOR U27595 ( .A(n22890), .B(n22894), .Z(n22928) );
  NAND U27596 ( .A(n22929), .B(n22930), .Z(n22894) );
  NAND U27597 ( .A(n22931), .B(n22932), .Z(n22930) );
  NAND U27598 ( .A(n22933), .B(n22934), .Z(n22929) );
  AND U27599 ( .A(n22935), .B(n22936), .Z(n22890) );
  NAND U27600 ( .A(n22937), .B(n22938), .Z(n22936) );
  NAND U27601 ( .A(n22939), .B(n22940), .Z(n22935) );
  AND U27602 ( .A(n22941), .B(n22942), .Z(n22892) );
  NAND U27603 ( .A(n22943), .B(n22944), .Z(n22886) );
  XNOR U27604 ( .A(n22869), .B(n22945), .Z(n22883) );
  XOR U27605 ( .A(n22873), .B(n22871), .Z(n22945) );
  XOR U27606 ( .A(n22879), .B(n22946), .Z(n22871) );
  XOR U27607 ( .A(n22876), .B(n22880), .Z(n22946) );
  NAND U27608 ( .A(n22947), .B(n22948), .Z(n22880) );
  NAND U27609 ( .A(n22949), .B(n22950), .Z(n22948) );
  NAND U27610 ( .A(n22951), .B(n22952), .Z(n22947) );
  AND U27611 ( .A(n22953), .B(n22954), .Z(n22876) );
  NAND U27612 ( .A(n22955), .B(n22956), .Z(n22954) );
  NAND U27613 ( .A(n22957), .B(n22958), .Z(n22953) );
  NANDN U27614 ( .A(n22959), .B(n22960), .Z(n22879) );
  NANDN U27615 ( .A(n22961), .B(n22962), .Z(n22873) );
  XNOR U27616 ( .A(n22864), .B(n22963), .Z(n22869) );
  XOR U27617 ( .A(n22862), .B(n22866), .Z(n22963) );
  NAND U27618 ( .A(n22964), .B(n22965), .Z(n22866) );
  NAND U27619 ( .A(n22966), .B(n22967), .Z(n22965) );
  NAND U27620 ( .A(n22968), .B(n22969), .Z(n22964) );
  AND U27621 ( .A(n22970), .B(n22971), .Z(n22862) );
  NAND U27622 ( .A(n22972), .B(n22973), .Z(n22971) );
  NAND U27623 ( .A(n22974), .B(n22975), .Z(n22970) );
  AND U27624 ( .A(n22976), .B(n22977), .Z(n22864) );
  XOR U27625 ( .A(n22944), .B(n22943), .Z(N28265) );
  XNOR U27626 ( .A(n22962), .B(n22961), .Z(n22943) );
  XNOR U27627 ( .A(n22976), .B(n22977), .Z(n22961) );
  XOR U27628 ( .A(n22973), .B(n22972), .Z(n22977) );
  XOR U27629 ( .A(y[675]), .B(x[675]), .Z(n22972) );
  XOR U27630 ( .A(n22975), .B(n22974), .Z(n22973) );
  XOR U27631 ( .A(y[677]), .B(x[677]), .Z(n22974) );
  XOR U27632 ( .A(y[676]), .B(x[676]), .Z(n22975) );
  XOR U27633 ( .A(n22967), .B(n22966), .Z(n22976) );
  XOR U27634 ( .A(n22969), .B(n22968), .Z(n22966) );
  XOR U27635 ( .A(y[674]), .B(x[674]), .Z(n22968) );
  XOR U27636 ( .A(y[673]), .B(x[673]), .Z(n22969) );
  XOR U27637 ( .A(y[672]), .B(x[672]), .Z(n22967) );
  XNOR U27638 ( .A(n22960), .B(n22959), .Z(n22962) );
  XNOR U27639 ( .A(n22956), .B(n22955), .Z(n22959) );
  XOR U27640 ( .A(n22958), .B(n22957), .Z(n22955) );
  XOR U27641 ( .A(y[671]), .B(x[671]), .Z(n22957) );
  XOR U27642 ( .A(y[670]), .B(x[670]), .Z(n22958) );
  XOR U27643 ( .A(y[669]), .B(x[669]), .Z(n22956) );
  XOR U27644 ( .A(n22950), .B(n22949), .Z(n22960) );
  XOR U27645 ( .A(n22952), .B(n22951), .Z(n22949) );
  XOR U27646 ( .A(y[668]), .B(x[668]), .Z(n22951) );
  XOR U27647 ( .A(y[667]), .B(x[667]), .Z(n22952) );
  XOR U27648 ( .A(y[666]), .B(x[666]), .Z(n22950) );
  XNOR U27649 ( .A(n22927), .B(n22926), .Z(n22944) );
  XNOR U27650 ( .A(n22941), .B(n22942), .Z(n22926) );
  XOR U27651 ( .A(n22938), .B(n22937), .Z(n22942) );
  XOR U27652 ( .A(y[663]), .B(x[663]), .Z(n22937) );
  XOR U27653 ( .A(n22940), .B(n22939), .Z(n22938) );
  XOR U27654 ( .A(y[665]), .B(x[665]), .Z(n22939) );
  XOR U27655 ( .A(y[664]), .B(x[664]), .Z(n22940) );
  XOR U27656 ( .A(n22932), .B(n22931), .Z(n22941) );
  XOR U27657 ( .A(n22934), .B(n22933), .Z(n22931) );
  XOR U27658 ( .A(y[662]), .B(x[662]), .Z(n22933) );
  XOR U27659 ( .A(y[661]), .B(x[661]), .Z(n22934) );
  XOR U27660 ( .A(y[660]), .B(x[660]), .Z(n22932) );
  XNOR U27661 ( .A(n22925), .B(n22924), .Z(n22927) );
  XNOR U27662 ( .A(n22921), .B(n22920), .Z(n22924) );
  XOR U27663 ( .A(n22923), .B(n22922), .Z(n22920) );
  XOR U27664 ( .A(y[659]), .B(x[659]), .Z(n22922) );
  XOR U27665 ( .A(y[658]), .B(x[658]), .Z(n22923) );
  XOR U27666 ( .A(y[657]), .B(x[657]), .Z(n22921) );
  XOR U27667 ( .A(n22915), .B(n22914), .Z(n22925) );
  XOR U27668 ( .A(n22917), .B(n22916), .Z(n22914) );
  XOR U27669 ( .A(y[656]), .B(x[656]), .Z(n22916) );
  XOR U27670 ( .A(y[655]), .B(x[655]), .Z(n22917) );
  XOR U27671 ( .A(y[654]), .B(x[654]), .Z(n22915) );
  NAND U27672 ( .A(n22978), .B(n22979), .Z(N28257) );
  NAND U27673 ( .A(n22980), .B(n22981), .Z(n22979) );
  NANDN U27674 ( .A(n22982), .B(n22983), .Z(n22981) );
  NANDN U27675 ( .A(n22983), .B(n22982), .Z(n22978) );
  XOR U27676 ( .A(n22982), .B(n22984), .Z(N28256) );
  XNOR U27677 ( .A(n22980), .B(n22983), .Z(n22984) );
  NAND U27678 ( .A(n22985), .B(n22986), .Z(n22983) );
  NAND U27679 ( .A(n22987), .B(n22988), .Z(n22986) );
  NANDN U27680 ( .A(n22989), .B(n22990), .Z(n22988) );
  NANDN U27681 ( .A(n22990), .B(n22989), .Z(n22985) );
  AND U27682 ( .A(n22991), .B(n22992), .Z(n22980) );
  NAND U27683 ( .A(n22993), .B(n22994), .Z(n22992) );
  OR U27684 ( .A(n22995), .B(n22996), .Z(n22994) );
  NAND U27685 ( .A(n22996), .B(n22995), .Z(n22991) );
  IV U27686 ( .A(n22997), .Z(n22996) );
  AND U27687 ( .A(n22998), .B(n22999), .Z(n22982) );
  NAND U27688 ( .A(n23000), .B(n23001), .Z(n22999) );
  NANDN U27689 ( .A(n23002), .B(n23003), .Z(n23001) );
  NANDN U27690 ( .A(n23003), .B(n23002), .Z(n22998) );
  XOR U27691 ( .A(n22995), .B(n23004), .Z(N28255) );
  XOR U27692 ( .A(n22993), .B(n22997), .Z(n23004) );
  XNOR U27693 ( .A(n22990), .B(n23005), .Z(n22997) );
  XNOR U27694 ( .A(n22987), .B(n22989), .Z(n23005) );
  AND U27695 ( .A(n23006), .B(n23007), .Z(n22989) );
  NANDN U27696 ( .A(n23008), .B(n23009), .Z(n23007) );
  NANDN U27697 ( .A(n23010), .B(n23011), .Z(n23009) );
  IV U27698 ( .A(n23012), .Z(n23011) );
  NAND U27699 ( .A(n23012), .B(n23010), .Z(n23006) );
  AND U27700 ( .A(n23013), .B(n23014), .Z(n22987) );
  NAND U27701 ( .A(n23015), .B(n23016), .Z(n23014) );
  OR U27702 ( .A(n23017), .B(n23018), .Z(n23016) );
  NAND U27703 ( .A(n23018), .B(n23017), .Z(n23013) );
  IV U27704 ( .A(n23019), .Z(n23018) );
  NAND U27705 ( .A(n23020), .B(n23021), .Z(n22990) );
  NANDN U27706 ( .A(n23022), .B(n23023), .Z(n23021) );
  NAND U27707 ( .A(n23024), .B(n23025), .Z(n23023) );
  OR U27708 ( .A(n23025), .B(n23024), .Z(n23020) );
  IV U27709 ( .A(n23026), .Z(n23024) );
  AND U27710 ( .A(n23027), .B(n23028), .Z(n22993) );
  NAND U27711 ( .A(n23029), .B(n23030), .Z(n23028) );
  NANDN U27712 ( .A(n23031), .B(n23032), .Z(n23030) );
  NANDN U27713 ( .A(n23032), .B(n23031), .Z(n23027) );
  XOR U27714 ( .A(n23003), .B(n23033), .Z(n22995) );
  XNOR U27715 ( .A(n23000), .B(n23002), .Z(n23033) );
  AND U27716 ( .A(n23034), .B(n23035), .Z(n23002) );
  NANDN U27717 ( .A(n23036), .B(n23037), .Z(n23035) );
  NANDN U27718 ( .A(n23038), .B(n23039), .Z(n23037) );
  IV U27719 ( .A(n23040), .Z(n23039) );
  NAND U27720 ( .A(n23040), .B(n23038), .Z(n23034) );
  AND U27721 ( .A(n23041), .B(n23042), .Z(n23000) );
  NAND U27722 ( .A(n23043), .B(n23044), .Z(n23042) );
  OR U27723 ( .A(n23045), .B(n23046), .Z(n23044) );
  NAND U27724 ( .A(n23046), .B(n23045), .Z(n23041) );
  IV U27725 ( .A(n23047), .Z(n23046) );
  NAND U27726 ( .A(n23048), .B(n23049), .Z(n23003) );
  NANDN U27727 ( .A(n23050), .B(n23051), .Z(n23049) );
  NAND U27728 ( .A(n23052), .B(n23053), .Z(n23051) );
  OR U27729 ( .A(n23053), .B(n23052), .Z(n23048) );
  IV U27730 ( .A(n23054), .Z(n23052) );
  XOR U27731 ( .A(n23029), .B(n23055), .Z(N28254) );
  XNOR U27732 ( .A(n23032), .B(n23031), .Z(n23055) );
  XNOR U27733 ( .A(n23043), .B(n23056), .Z(n23031) );
  XOR U27734 ( .A(n23047), .B(n23045), .Z(n23056) );
  XOR U27735 ( .A(n23053), .B(n23057), .Z(n23045) );
  XOR U27736 ( .A(n23050), .B(n23054), .Z(n23057) );
  NAND U27737 ( .A(n23058), .B(n23059), .Z(n23054) );
  NAND U27738 ( .A(n23060), .B(n23061), .Z(n23059) );
  NAND U27739 ( .A(n23062), .B(n23063), .Z(n23058) );
  AND U27740 ( .A(n23064), .B(n23065), .Z(n23050) );
  NAND U27741 ( .A(n23066), .B(n23067), .Z(n23065) );
  NAND U27742 ( .A(n23068), .B(n23069), .Z(n23064) );
  NANDN U27743 ( .A(n23070), .B(n23071), .Z(n23053) );
  NANDN U27744 ( .A(n23072), .B(n23073), .Z(n23047) );
  XNOR U27745 ( .A(n23038), .B(n23074), .Z(n23043) );
  XOR U27746 ( .A(n23036), .B(n23040), .Z(n23074) );
  NAND U27747 ( .A(n23075), .B(n23076), .Z(n23040) );
  NAND U27748 ( .A(n23077), .B(n23078), .Z(n23076) );
  NAND U27749 ( .A(n23079), .B(n23080), .Z(n23075) );
  AND U27750 ( .A(n23081), .B(n23082), .Z(n23036) );
  NAND U27751 ( .A(n23083), .B(n23084), .Z(n23082) );
  NAND U27752 ( .A(n23085), .B(n23086), .Z(n23081) );
  AND U27753 ( .A(n23087), .B(n23088), .Z(n23038) );
  NAND U27754 ( .A(n23089), .B(n23090), .Z(n23032) );
  XNOR U27755 ( .A(n23015), .B(n23091), .Z(n23029) );
  XOR U27756 ( .A(n23019), .B(n23017), .Z(n23091) );
  XOR U27757 ( .A(n23025), .B(n23092), .Z(n23017) );
  XOR U27758 ( .A(n23022), .B(n23026), .Z(n23092) );
  NAND U27759 ( .A(n23093), .B(n23094), .Z(n23026) );
  NAND U27760 ( .A(n23095), .B(n23096), .Z(n23094) );
  NAND U27761 ( .A(n23097), .B(n23098), .Z(n23093) );
  AND U27762 ( .A(n23099), .B(n23100), .Z(n23022) );
  NAND U27763 ( .A(n23101), .B(n23102), .Z(n23100) );
  NAND U27764 ( .A(n23103), .B(n23104), .Z(n23099) );
  NANDN U27765 ( .A(n23105), .B(n23106), .Z(n23025) );
  NANDN U27766 ( .A(n23107), .B(n23108), .Z(n23019) );
  XNOR U27767 ( .A(n23010), .B(n23109), .Z(n23015) );
  XOR U27768 ( .A(n23008), .B(n23012), .Z(n23109) );
  NAND U27769 ( .A(n23110), .B(n23111), .Z(n23012) );
  NAND U27770 ( .A(n23112), .B(n23113), .Z(n23111) );
  NAND U27771 ( .A(n23114), .B(n23115), .Z(n23110) );
  AND U27772 ( .A(n23116), .B(n23117), .Z(n23008) );
  NAND U27773 ( .A(n23118), .B(n23119), .Z(n23117) );
  NAND U27774 ( .A(n23120), .B(n23121), .Z(n23116) );
  AND U27775 ( .A(n23122), .B(n23123), .Z(n23010) );
  XOR U27776 ( .A(n23090), .B(n23089), .Z(N28253) );
  XNOR U27777 ( .A(n23108), .B(n23107), .Z(n23089) );
  XNOR U27778 ( .A(n23122), .B(n23123), .Z(n23107) );
  XOR U27779 ( .A(n23119), .B(n23118), .Z(n23123) );
  XOR U27780 ( .A(y[651]), .B(x[651]), .Z(n23118) );
  XOR U27781 ( .A(n23121), .B(n23120), .Z(n23119) );
  XOR U27782 ( .A(y[653]), .B(x[653]), .Z(n23120) );
  XOR U27783 ( .A(y[652]), .B(x[652]), .Z(n23121) );
  XOR U27784 ( .A(n23113), .B(n23112), .Z(n23122) );
  XOR U27785 ( .A(n23115), .B(n23114), .Z(n23112) );
  XOR U27786 ( .A(y[650]), .B(x[650]), .Z(n23114) );
  XOR U27787 ( .A(y[649]), .B(x[649]), .Z(n23115) );
  XOR U27788 ( .A(y[648]), .B(x[648]), .Z(n23113) );
  XNOR U27789 ( .A(n23106), .B(n23105), .Z(n23108) );
  XNOR U27790 ( .A(n23102), .B(n23101), .Z(n23105) );
  XOR U27791 ( .A(n23104), .B(n23103), .Z(n23101) );
  XOR U27792 ( .A(y[647]), .B(x[647]), .Z(n23103) );
  XOR U27793 ( .A(y[646]), .B(x[646]), .Z(n23104) );
  XOR U27794 ( .A(y[645]), .B(x[645]), .Z(n23102) );
  XOR U27795 ( .A(n23096), .B(n23095), .Z(n23106) );
  XOR U27796 ( .A(n23098), .B(n23097), .Z(n23095) );
  XOR U27797 ( .A(y[644]), .B(x[644]), .Z(n23097) );
  XOR U27798 ( .A(y[643]), .B(x[643]), .Z(n23098) );
  XOR U27799 ( .A(y[642]), .B(x[642]), .Z(n23096) );
  XNOR U27800 ( .A(n23073), .B(n23072), .Z(n23090) );
  XNOR U27801 ( .A(n23087), .B(n23088), .Z(n23072) );
  XOR U27802 ( .A(n23084), .B(n23083), .Z(n23088) );
  XOR U27803 ( .A(y[639]), .B(x[639]), .Z(n23083) );
  XOR U27804 ( .A(n23086), .B(n23085), .Z(n23084) );
  XOR U27805 ( .A(y[641]), .B(x[641]), .Z(n23085) );
  XOR U27806 ( .A(y[640]), .B(x[640]), .Z(n23086) );
  XOR U27807 ( .A(n23078), .B(n23077), .Z(n23087) );
  XOR U27808 ( .A(n23080), .B(n23079), .Z(n23077) );
  XOR U27809 ( .A(y[638]), .B(x[638]), .Z(n23079) );
  XOR U27810 ( .A(y[637]), .B(x[637]), .Z(n23080) );
  XOR U27811 ( .A(y[636]), .B(x[636]), .Z(n23078) );
  XNOR U27812 ( .A(n23071), .B(n23070), .Z(n23073) );
  XNOR U27813 ( .A(n23067), .B(n23066), .Z(n23070) );
  XOR U27814 ( .A(n23069), .B(n23068), .Z(n23066) );
  XOR U27815 ( .A(y[635]), .B(x[635]), .Z(n23068) );
  XOR U27816 ( .A(y[634]), .B(x[634]), .Z(n23069) );
  XOR U27817 ( .A(y[633]), .B(x[633]), .Z(n23067) );
  XOR U27818 ( .A(n23061), .B(n23060), .Z(n23071) );
  XOR U27819 ( .A(n23063), .B(n23062), .Z(n23060) );
  XOR U27820 ( .A(y[632]), .B(x[632]), .Z(n23062) );
  XOR U27821 ( .A(y[631]), .B(x[631]), .Z(n23063) );
  XOR U27822 ( .A(y[630]), .B(x[630]), .Z(n23061) );
  NAND U27823 ( .A(n23124), .B(n23125), .Z(N28245) );
  NAND U27824 ( .A(n23126), .B(n23127), .Z(n23125) );
  NANDN U27825 ( .A(n23128), .B(n23129), .Z(n23127) );
  NANDN U27826 ( .A(n23129), .B(n23128), .Z(n23124) );
  XOR U27827 ( .A(n23128), .B(n23130), .Z(N28244) );
  XNOR U27828 ( .A(n23126), .B(n23129), .Z(n23130) );
  NAND U27829 ( .A(n23131), .B(n23132), .Z(n23129) );
  NAND U27830 ( .A(n23133), .B(n23134), .Z(n23132) );
  NANDN U27831 ( .A(n23135), .B(n23136), .Z(n23134) );
  NANDN U27832 ( .A(n23136), .B(n23135), .Z(n23131) );
  AND U27833 ( .A(n23137), .B(n23138), .Z(n23126) );
  NAND U27834 ( .A(n23139), .B(n23140), .Z(n23138) );
  OR U27835 ( .A(n23141), .B(n23142), .Z(n23140) );
  NAND U27836 ( .A(n23142), .B(n23141), .Z(n23137) );
  IV U27837 ( .A(n23143), .Z(n23142) );
  AND U27838 ( .A(n23144), .B(n23145), .Z(n23128) );
  NAND U27839 ( .A(n23146), .B(n23147), .Z(n23145) );
  NANDN U27840 ( .A(n23148), .B(n23149), .Z(n23147) );
  NANDN U27841 ( .A(n23149), .B(n23148), .Z(n23144) );
  XOR U27842 ( .A(n23141), .B(n23150), .Z(N28243) );
  XOR U27843 ( .A(n23139), .B(n23143), .Z(n23150) );
  XNOR U27844 ( .A(n23136), .B(n23151), .Z(n23143) );
  XNOR U27845 ( .A(n23133), .B(n23135), .Z(n23151) );
  AND U27846 ( .A(n23152), .B(n23153), .Z(n23135) );
  NANDN U27847 ( .A(n23154), .B(n23155), .Z(n23153) );
  NANDN U27848 ( .A(n23156), .B(n23157), .Z(n23155) );
  IV U27849 ( .A(n23158), .Z(n23157) );
  NAND U27850 ( .A(n23158), .B(n23156), .Z(n23152) );
  AND U27851 ( .A(n23159), .B(n23160), .Z(n23133) );
  NAND U27852 ( .A(n23161), .B(n23162), .Z(n23160) );
  OR U27853 ( .A(n23163), .B(n23164), .Z(n23162) );
  NAND U27854 ( .A(n23164), .B(n23163), .Z(n23159) );
  IV U27855 ( .A(n23165), .Z(n23164) );
  NAND U27856 ( .A(n23166), .B(n23167), .Z(n23136) );
  NANDN U27857 ( .A(n23168), .B(n23169), .Z(n23167) );
  NAND U27858 ( .A(n23170), .B(n23171), .Z(n23169) );
  OR U27859 ( .A(n23171), .B(n23170), .Z(n23166) );
  IV U27860 ( .A(n23172), .Z(n23170) );
  AND U27861 ( .A(n23173), .B(n23174), .Z(n23139) );
  NAND U27862 ( .A(n23175), .B(n23176), .Z(n23174) );
  NANDN U27863 ( .A(n23177), .B(n23178), .Z(n23176) );
  NANDN U27864 ( .A(n23178), .B(n23177), .Z(n23173) );
  XOR U27865 ( .A(n23149), .B(n23179), .Z(n23141) );
  XNOR U27866 ( .A(n23146), .B(n23148), .Z(n23179) );
  AND U27867 ( .A(n23180), .B(n23181), .Z(n23148) );
  NANDN U27868 ( .A(n23182), .B(n23183), .Z(n23181) );
  NANDN U27869 ( .A(n23184), .B(n23185), .Z(n23183) );
  IV U27870 ( .A(n23186), .Z(n23185) );
  NAND U27871 ( .A(n23186), .B(n23184), .Z(n23180) );
  AND U27872 ( .A(n23187), .B(n23188), .Z(n23146) );
  NAND U27873 ( .A(n23189), .B(n23190), .Z(n23188) );
  OR U27874 ( .A(n23191), .B(n23192), .Z(n23190) );
  NAND U27875 ( .A(n23192), .B(n23191), .Z(n23187) );
  IV U27876 ( .A(n23193), .Z(n23192) );
  NAND U27877 ( .A(n23194), .B(n23195), .Z(n23149) );
  NANDN U27878 ( .A(n23196), .B(n23197), .Z(n23195) );
  NAND U27879 ( .A(n23198), .B(n23199), .Z(n23197) );
  OR U27880 ( .A(n23199), .B(n23198), .Z(n23194) );
  IV U27881 ( .A(n23200), .Z(n23198) );
  XOR U27882 ( .A(n23175), .B(n23201), .Z(N28242) );
  XNOR U27883 ( .A(n23178), .B(n23177), .Z(n23201) );
  XNOR U27884 ( .A(n23189), .B(n23202), .Z(n23177) );
  XOR U27885 ( .A(n23193), .B(n23191), .Z(n23202) );
  XOR U27886 ( .A(n23199), .B(n23203), .Z(n23191) );
  XOR U27887 ( .A(n23196), .B(n23200), .Z(n23203) );
  NAND U27888 ( .A(n23204), .B(n23205), .Z(n23200) );
  NAND U27889 ( .A(n23206), .B(n23207), .Z(n23205) );
  NAND U27890 ( .A(n23208), .B(n23209), .Z(n23204) );
  AND U27891 ( .A(n23210), .B(n23211), .Z(n23196) );
  NAND U27892 ( .A(n23212), .B(n23213), .Z(n23211) );
  NAND U27893 ( .A(n23214), .B(n23215), .Z(n23210) );
  NANDN U27894 ( .A(n23216), .B(n23217), .Z(n23199) );
  NANDN U27895 ( .A(n23218), .B(n23219), .Z(n23193) );
  XNOR U27896 ( .A(n23184), .B(n23220), .Z(n23189) );
  XOR U27897 ( .A(n23182), .B(n23186), .Z(n23220) );
  NAND U27898 ( .A(n23221), .B(n23222), .Z(n23186) );
  NAND U27899 ( .A(n23223), .B(n23224), .Z(n23222) );
  NAND U27900 ( .A(n23225), .B(n23226), .Z(n23221) );
  AND U27901 ( .A(n23227), .B(n23228), .Z(n23182) );
  NAND U27902 ( .A(n23229), .B(n23230), .Z(n23228) );
  NAND U27903 ( .A(n23231), .B(n23232), .Z(n23227) );
  AND U27904 ( .A(n23233), .B(n23234), .Z(n23184) );
  NAND U27905 ( .A(n23235), .B(n23236), .Z(n23178) );
  XNOR U27906 ( .A(n23161), .B(n23237), .Z(n23175) );
  XOR U27907 ( .A(n23165), .B(n23163), .Z(n23237) );
  XOR U27908 ( .A(n23171), .B(n23238), .Z(n23163) );
  XOR U27909 ( .A(n23168), .B(n23172), .Z(n23238) );
  NAND U27910 ( .A(n23239), .B(n23240), .Z(n23172) );
  NAND U27911 ( .A(n23241), .B(n23242), .Z(n23240) );
  NAND U27912 ( .A(n23243), .B(n23244), .Z(n23239) );
  AND U27913 ( .A(n23245), .B(n23246), .Z(n23168) );
  NAND U27914 ( .A(n23247), .B(n23248), .Z(n23246) );
  NAND U27915 ( .A(n23249), .B(n23250), .Z(n23245) );
  NANDN U27916 ( .A(n23251), .B(n23252), .Z(n23171) );
  NANDN U27917 ( .A(n23253), .B(n23254), .Z(n23165) );
  XNOR U27918 ( .A(n23156), .B(n23255), .Z(n23161) );
  XOR U27919 ( .A(n23154), .B(n23158), .Z(n23255) );
  NAND U27920 ( .A(n23256), .B(n23257), .Z(n23158) );
  NAND U27921 ( .A(n23258), .B(n23259), .Z(n23257) );
  NAND U27922 ( .A(n23260), .B(n23261), .Z(n23256) );
  AND U27923 ( .A(n23262), .B(n23263), .Z(n23154) );
  NAND U27924 ( .A(n23264), .B(n23265), .Z(n23263) );
  NAND U27925 ( .A(n23266), .B(n23267), .Z(n23262) );
  AND U27926 ( .A(n23268), .B(n23269), .Z(n23156) );
  XOR U27927 ( .A(n23236), .B(n23235), .Z(N28241) );
  XNOR U27928 ( .A(n23254), .B(n23253), .Z(n23235) );
  XNOR U27929 ( .A(n23268), .B(n23269), .Z(n23253) );
  XOR U27930 ( .A(n23265), .B(n23264), .Z(n23269) );
  XOR U27931 ( .A(y[627]), .B(x[627]), .Z(n23264) );
  XOR U27932 ( .A(n23267), .B(n23266), .Z(n23265) );
  XOR U27933 ( .A(y[629]), .B(x[629]), .Z(n23266) );
  XOR U27934 ( .A(y[628]), .B(x[628]), .Z(n23267) );
  XOR U27935 ( .A(n23259), .B(n23258), .Z(n23268) );
  XOR U27936 ( .A(n23261), .B(n23260), .Z(n23258) );
  XOR U27937 ( .A(y[626]), .B(x[626]), .Z(n23260) );
  XOR U27938 ( .A(y[625]), .B(x[625]), .Z(n23261) );
  XOR U27939 ( .A(y[624]), .B(x[624]), .Z(n23259) );
  XNOR U27940 ( .A(n23252), .B(n23251), .Z(n23254) );
  XNOR U27941 ( .A(n23248), .B(n23247), .Z(n23251) );
  XOR U27942 ( .A(n23250), .B(n23249), .Z(n23247) );
  XOR U27943 ( .A(y[623]), .B(x[623]), .Z(n23249) );
  XOR U27944 ( .A(y[622]), .B(x[622]), .Z(n23250) );
  XOR U27945 ( .A(y[621]), .B(x[621]), .Z(n23248) );
  XOR U27946 ( .A(n23242), .B(n23241), .Z(n23252) );
  XOR U27947 ( .A(n23244), .B(n23243), .Z(n23241) );
  XOR U27948 ( .A(y[620]), .B(x[620]), .Z(n23243) );
  XOR U27949 ( .A(y[619]), .B(x[619]), .Z(n23244) );
  XOR U27950 ( .A(y[618]), .B(x[618]), .Z(n23242) );
  XNOR U27951 ( .A(n23219), .B(n23218), .Z(n23236) );
  XNOR U27952 ( .A(n23233), .B(n23234), .Z(n23218) );
  XOR U27953 ( .A(n23230), .B(n23229), .Z(n23234) );
  XOR U27954 ( .A(y[615]), .B(x[615]), .Z(n23229) );
  XOR U27955 ( .A(n23232), .B(n23231), .Z(n23230) );
  XOR U27956 ( .A(y[617]), .B(x[617]), .Z(n23231) );
  XOR U27957 ( .A(y[616]), .B(x[616]), .Z(n23232) );
  XOR U27958 ( .A(n23224), .B(n23223), .Z(n23233) );
  XOR U27959 ( .A(n23226), .B(n23225), .Z(n23223) );
  XOR U27960 ( .A(y[614]), .B(x[614]), .Z(n23225) );
  XOR U27961 ( .A(y[613]), .B(x[613]), .Z(n23226) );
  XOR U27962 ( .A(y[612]), .B(x[612]), .Z(n23224) );
  XNOR U27963 ( .A(n23217), .B(n23216), .Z(n23219) );
  XNOR U27964 ( .A(n23213), .B(n23212), .Z(n23216) );
  XOR U27965 ( .A(n23215), .B(n23214), .Z(n23212) );
  XOR U27966 ( .A(y[611]), .B(x[611]), .Z(n23214) );
  XOR U27967 ( .A(y[610]), .B(x[610]), .Z(n23215) );
  XOR U27968 ( .A(y[609]), .B(x[609]), .Z(n23213) );
  XOR U27969 ( .A(n23207), .B(n23206), .Z(n23217) );
  XOR U27970 ( .A(n23209), .B(n23208), .Z(n23206) );
  XOR U27971 ( .A(y[608]), .B(x[608]), .Z(n23208) );
  XOR U27972 ( .A(y[607]), .B(x[607]), .Z(n23209) );
  XOR U27973 ( .A(y[606]), .B(x[606]), .Z(n23207) );
  NAND U27974 ( .A(n23270), .B(n23271), .Z(N28233) );
  NAND U27975 ( .A(n23272), .B(n23273), .Z(n23271) );
  NANDN U27976 ( .A(n23274), .B(n23275), .Z(n23273) );
  NANDN U27977 ( .A(n23275), .B(n23274), .Z(n23270) );
  XOR U27978 ( .A(n23274), .B(n23276), .Z(N28232) );
  XNOR U27979 ( .A(n23272), .B(n23275), .Z(n23276) );
  NAND U27980 ( .A(n23277), .B(n23278), .Z(n23275) );
  NAND U27981 ( .A(n23279), .B(n23280), .Z(n23278) );
  NANDN U27982 ( .A(n23281), .B(n23282), .Z(n23280) );
  NANDN U27983 ( .A(n23282), .B(n23281), .Z(n23277) );
  AND U27984 ( .A(n23283), .B(n23284), .Z(n23272) );
  NAND U27985 ( .A(n23285), .B(n23286), .Z(n23284) );
  OR U27986 ( .A(n23287), .B(n23288), .Z(n23286) );
  NAND U27987 ( .A(n23288), .B(n23287), .Z(n23283) );
  IV U27988 ( .A(n23289), .Z(n23288) );
  AND U27989 ( .A(n23290), .B(n23291), .Z(n23274) );
  NAND U27990 ( .A(n23292), .B(n23293), .Z(n23291) );
  NANDN U27991 ( .A(n23294), .B(n23295), .Z(n23293) );
  NANDN U27992 ( .A(n23295), .B(n23294), .Z(n23290) );
  XOR U27993 ( .A(n23287), .B(n23296), .Z(N28231) );
  XOR U27994 ( .A(n23285), .B(n23289), .Z(n23296) );
  XNOR U27995 ( .A(n23282), .B(n23297), .Z(n23289) );
  XNOR U27996 ( .A(n23279), .B(n23281), .Z(n23297) );
  AND U27997 ( .A(n23298), .B(n23299), .Z(n23281) );
  NANDN U27998 ( .A(n23300), .B(n23301), .Z(n23299) );
  NANDN U27999 ( .A(n23302), .B(n23303), .Z(n23301) );
  IV U28000 ( .A(n23304), .Z(n23303) );
  NAND U28001 ( .A(n23304), .B(n23302), .Z(n23298) );
  AND U28002 ( .A(n23305), .B(n23306), .Z(n23279) );
  NAND U28003 ( .A(n23307), .B(n23308), .Z(n23306) );
  OR U28004 ( .A(n23309), .B(n23310), .Z(n23308) );
  NAND U28005 ( .A(n23310), .B(n23309), .Z(n23305) );
  IV U28006 ( .A(n23311), .Z(n23310) );
  NAND U28007 ( .A(n23312), .B(n23313), .Z(n23282) );
  NANDN U28008 ( .A(n23314), .B(n23315), .Z(n23313) );
  NAND U28009 ( .A(n23316), .B(n23317), .Z(n23315) );
  OR U28010 ( .A(n23317), .B(n23316), .Z(n23312) );
  IV U28011 ( .A(n23318), .Z(n23316) );
  AND U28012 ( .A(n23319), .B(n23320), .Z(n23285) );
  NAND U28013 ( .A(n23321), .B(n23322), .Z(n23320) );
  NANDN U28014 ( .A(n23323), .B(n23324), .Z(n23322) );
  NANDN U28015 ( .A(n23324), .B(n23323), .Z(n23319) );
  XOR U28016 ( .A(n23295), .B(n23325), .Z(n23287) );
  XNOR U28017 ( .A(n23292), .B(n23294), .Z(n23325) );
  AND U28018 ( .A(n23326), .B(n23327), .Z(n23294) );
  NANDN U28019 ( .A(n23328), .B(n23329), .Z(n23327) );
  NANDN U28020 ( .A(n23330), .B(n23331), .Z(n23329) );
  IV U28021 ( .A(n23332), .Z(n23331) );
  NAND U28022 ( .A(n23332), .B(n23330), .Z(n23326) );
  AND U28023 ( .A(n23333), .B(n23334), .Z(n23292) );
  NAND U28024 ( .A(n23335), .B(n23336), .Z(n23334) );
  OR U28025 ( .A(n23337), .B(n23338), .Z(n23336) );
  NAND U28026 ( .A(n23338), .B(n23337), .Z(n23333) );
  IV U28027 ( .A(n23339), .Z(n23338) );
  NAND U28028 ( .A(n23340), .B(n23341), .Z(n23295) );
  NANDN U28029 ( .A(n23342), .B(n23343), .Z(n23341) );
  NAND U28030 ( .A(n23344), .B(n23345), .Z(n23343) );
  OR U28031 ( .A(n23345), .B(n23344), .Z(n23340) );
  IV U28032 ( .A(n23346), .Z(n23344) );
  XOR U28033 ( .A(n23321), .B(n23347), .Z(N28230) );
  XNOR U28034 ( .A(n23324), .B(n23323), .Z(n23347) );
  XNOR U28035 ( .A(n23335), .B(n23348), .Z(n23323) );
  XOR U28036 ( .A(n23339), .B(n23337), .Z(n23348) );
  XOR U28037 ( .A(n23345), .B(n23349), .Z(n23337) );
  XOR U28038 ( .A(n23342), .B(n23346), .Z(n23349) );
  NAND U28039 ( .A(n23350), .B(n23351), .Z(n23346) );
  NAND U28040 ( .A(n23352), .B(n23353), .Z(n23351) );
  NAND U28041 ( .A(n23354), .B(n23355), .Z(n23350) );
  AND U28042 ( .A(n23356), .B(n23357), .Z(n23342) );
  NAND U28043 ( .A(n23358), .B(n23359), .Z(n23357) );
  NAND U28044 ( .A(n23360), .B(n23361), .Z(n23356) );
  NANDN U28045 ( .A(n23362), .B(n23363), .Z(n23345) );
  NANDN U28046 ( .A(n23364), .B(n23365), .Z(n23339) );
  XNOR U28047 ( .A(n23330), .B(n23366), .Z(n23335) );
  XOR U28048 ( .A(n23328), .B(n23332), .Z(n23366) );
  NAND U28049 ( .A(n23367), .B(n23368), .Z(n23332) );
  NAND U28050 ( .A(n23369), .B(n23370), .Z(n23368) );
  NAND U28051 ( .A(n23371), .B(n23372), .Z(n23367) );
  AND U28052 ( .A(n23373), .B(n23374), .Z(n23328) );
  NAND U28053 ( .A(n23375), .B(n23376), .Z(n23374) );
  NAND U28054 ( .A(n23377), .B(n23378), .Z(n23373) );
  AND U28055 ( .A(n23379), .B(n23380), .Z(n23330) );
  NAND U28056 ( .A(n23381), .B(n23382), .Z(n23324) );
  XNOR U28057 ( .A(n23307), .B(n23383), .Z(n23321) );
  XOR U28058 ( .A(n23311), .B(n23309), .Z(n23383) );
  XOR U28059 ( .A(n23317), .B(n23384), .Z(n23309) );
  XOR U28060 ( .A(n23314), .B(n23318), .Z(n23384) );
  NAND U28061 ( .A(n23385), .B(n23386), .Z(n23318) );
  NAND U28062 ( .A(n23387), .B(n23388), .Z(n23386) );
  NAND U28063 ( .A(n23389), .B(n23390), .Z(n23385) );
  AND U28064 ( .A(n23391), .B(n23392), .Z(n23314) );
  NAND U28065 ( .A(n23393), .B(n23394), .Z(n23392) );
  NAND U28066 ( .A(n23395), .B(n23396), .Z(n23391) );
  NANDN U28067 ( .A(n23397), .B(n23398), .Z(n23317) );
  NANDN U28068 ( .A(n23399), .B(n23400), .Z(n23311) );
  XNOR U28069 ( .A(n23302), .B(n23401), .Z(n23307) );
  XOR U28070 ( .A(n23300), .B(n23304), .Z(n23401) );
  NAND U28071 ( .A(n23402), .B(n23403), .Z(n23304) );
  NAND U28072 ( .A(n23404), .B(n23405), .Z(n23403) );
  NAND U28073 ( .A(n23406), .B(n23407), .Z(n23402) );
  AND U28074 ( .A(n23408), .B(n23409), .Z(n23300) );
  NAND U28075 ( .A(n23410), .B(n23411), .Z(n23409) );
  NAND U28076 ( .A(n23412), .B(n23413), .Z(n23408) );
  AND U28077 ( .A(n23414), .B(n23415), .Z(n23302) );
  XOR U28078 ( .A(n23382), .B(n23381), .Z(N28229) );
  XNOR U28079 ( .A(n23400), .B(n23399), .Z(n23381) );
  XNOR U28080 ( .A(n23414), .B(n23415), .Z(n23399) );
  XOR U28081 ( .A(n23411), .B(n23410), .Z(n23415) );
  XOR U28082 ( .A(y[603]), .B(x[603]), .Z(n23410) );
  XOR U28083 ( .A(n23413), .B(n23412), .Z(n23411) );
  XOR U28084 ( .A(y[605]), .B(x[605]), .Z(n23412) );
  XOR U28085 ( .A(y[604]), .B(x[604]), .Z(n23413) );
  XOR U28086 ( .A(n23405), .B(n23404), .Z(n23414) );
  XOR U28087 ( .A(n23407), .B(n23406), .Z(n23404) );
  XOR U28088 ( .A(y[602]), .B(x[602]), .Z(n23406) );
  XOR U28089 ( .A(y[601]), .B(x[601]), .Z(n23407) );
  XOR U28090 ( .A(y[600]), .B(x[600]), .Z(n23405) );
  XNOR U28091 ( .A(n23398), .B(n23397), .Z(n23400) );
  XNOR U28092 ( .A(n23394), .B(n23393), .Z(n23397) );
  XOR U28093 ( .A(n23396), .B(n23395), .Z(n23393) );
  XOR U28094 ( .A(y[599]), .B(x[599]), .Z(n23395) );
  XOR U28095 ( .A(y[598]), .B(x[598]), .Z(n23396) );
  XOR U28096 ( .A(y[597]), .B(x[597]), .Z(n23394) );
  XOR U28097 ( .A(n23388), .B(n23387), .Z(n23398) );
  XOR U28098 ( .A(n23390), .B(n23389), .Z(n23387) );
  XOR U28099 ( .A(y[596]), .B(x[596]), .Z(n23389) );
  XOR U28100 ( .A(y[595]), .B(x[595]), .Z(n23390) );
  XOR U28101 ( .A(y[594]), .B(x[594]), .Z(n23388) );
  XNOR U28102 ( .A(n23365), .B(n23364), .Z(n23382) );
  XNOR U28103 ( .A(n23379), .B(n23380), .Z(n23364) );
  XOR U28104 ( .A(n23376), .B(n23375), .Z(n23380) );
  XOR U28105 ( .A(y[591]), .B(x[591]), .Z(n23375) );
  XOR U28106 ( .A(n23378), .B(n23377), .Z(n23376) );
  XOR U28107 ( .A(y[593]), .B(x[593]), .Z(n23377) );
  XOR U28108 ( .A(y[592]), .B(x[592]), .Z(n23378) );
  XOR U28109 ( .A(n23370), .B(n23369), .Z(n23379) );
  XOR U28110 ( .A(n23372), .B(n23371), .Z(n23369) );
  XOR U28111 ( .A(y[590]), .B(x[590]), .Z(n23371) );
  XOR U28112 ( .A(y[589]), .B(x[589]), .Z(n23372) );
  XOR U28113 ( .A(y[588]), .B(x[588]), .Z(n23370) );
  XNOR U28114 ( .A(n23363), .B(n23362), .Z(n23365) );
  XNOR U28115 ( .A(n23359), .B(n23358), .Z(n23362) );
  XOR U28116 ( .A(n23361), .B(n23360), .Z(n23358) );
  XOR U28117 ( .A(y[587]), .B(x[587]), .Z(n23360) );
  XOR U28118 ( .A(y[586]), .B(x[586]), .Z(n23361) );
  XOR U28119 ( .A(y[585]), .B(x[585]), .Z(n23359) );
  XOR U28120 ( .A(n23353), .B(n23352), .Z(n23363) );
  XOR U28121 ( .A(n23355), .B(n23354), .Z(n23352) );
  XOR U28122 ( .A(y[584]), .B(x[584]), .Z(n23354) );
  XOR U28123 ( .A(y[583]), .B(x[583]), .Z(n23355) );
  XOR U28124 ( .A(y[582]), .B(x[582]), .Z(n23353) );
  NAND U28125 ( .A(n23416), .B(n23417), .Z(N28221) );
  NAND U28126 ( .A(n23418), .B(n23419), .Z(n23417) );
  NANDN U28127 ( .A(n23420), .B(n23421), .Z(n23419) );
  NANDN U28128 ( .A(n23421), .B(n23420), .Z(n23416) );
  XOR U28129 ( .A(n23420), .B(n23422), .Z(N28220) );
  XNOR U28130 ( .A(n23418), .B(n23421), .Z(n23422) );
  NAND U28131 ( .A(n23423), .B(n23424), .Z(n23421) );
  NAND U28132 ( .A(n23425), .B(n23426), .Z(n23424) );
  NANDN U28133 ( .A(n23427), .B(n23428), .Z(n23426) );
  NANDN U28134 ( .A(n23428), .B(n23427), .Z(n23423) );
  AND U28135 ( .A(n23429), .B(n23430), .Z(n23418) );
  NAND U28136 ( .A(n23431), .B(n23432), .Z(n23430) );
  OR U28137 ( .A(n23433), .B(n23434), .Z(n23432) );
  NAND U28138 ( .A(n23434), .B(n23433), .Z(n23429) );
  IV U28139 ( .A(n23435), .Z(n23434) );
  AND U28140 ( .A(n23436), .B(n23437), .Z(n23420) );
  NAND U28141 ( .A(n23438), .B(n23439), .Z(n23437) );
  NANDN U28142 ( .A(n23440), .B(n23441), .Z(n23439) );
  NANDN U28143 ( .A(n23441), .B(n23440), .Z(n23436) );
  XOR U28144 ( .A(n23433), .B(n23442), .Z(N28219) );
  XOR U28145 ( .A(n23431), .B(n23435), .Z(n23442) );
  XNOR U28146 ( .A(n23428), .B(n23443), .Z(n23435) );
  XNOR U28147 ( .A(n23425), .B(n23427), .Z(n23443) );
  AND U28148 ( .A(n23444), .B(n23445), .Z(n23427) );
  NANDN U28149 ( .A(n23446), .B(n23447), .Z(n23445) );
  NANDN U28150 ( .A(n23448), .B(n23449), .Z(n23447) );
  IV U28151 ( .A(n23450), .Z(n23449) );
  NAND U28152 ( .A(n23450), .B(n23448), .Z(n23444) );
  AND U28153 ( .A(n23451), .B(n23452), .Z(n23425) );
  NAND U28154 ( .A(n23453), .B(n23454), .Z(n23452) );
  OR U28155 ( .A(n23455), .B(n23456), .Z(n23454) );
  NAND U28156 ( .A(n23456), .B(n23455), .Z(n23451) );
  IV U28157 ( .A(n23457), .Z(n23456) );
  NAND U28158 ( .A(n23458), .B(n23459), .Z(n23428) );
  NANDN U28159 ( .A(n23460), .B(n23461), .Z(n23459) );
  NAND U28160 ( .A(n23462), .B(n23463), .Z(n23461) );
  OR U28161 ( .A(n23463), .B(n23462), .Z(n23458) );
  IV U28162 ( .A(n23464), .Z(n23462) );
  AND U28163 ( .A(n23465), .B(n23466), .Z(n23431) );
  NAND U28164 ( .A(n23467), .B(n23468), .Z(n23466) );
  NANDN U28165 ( .A(n23469), .B(n23470), .Z(n23468) );
  NANDN U28166 ( .A(n23470), .B(n23469), .Z(n23465) );
  XOR U28167 ( .A(n23441), .B(n23471), .Z(n23433) );
  XNOR U28168 ( .A(n23438), .B(n23440), .Z(n23471) );
  AND U28169 ( .A(n23472), .B(n23473), .Z(n23440) );
  NANDN U28170 ( .A(n23474), .B(n23475), .Z(n23473) );
  NANDN U28171 ( .A(n23476), .B(n23477), .Z(n23475) );
  IV U28172 ( .A(n23478), .Z(n23477) );
  NAND U28173 ( .A(n23478), .B(n23476), .Z(n23472) );
  AND U28174 ( .A(n23479), .B(n23480), .Z(n23438) );
  NAND U28175 ( .A(n23481), .B(n23482), .Z(n23480) );
  OR U28176 ( .A(n23483), .B(n23484), .Z(n23482) );
  NAND U28177 ( .A(n23484), .B(n23483), .Z(n23479) );
  IV U28178 ( .A(n23485), .Z(n23484) );
  NAND U28179 ( .A(n23486), .B(n23487), .Z(n23441) );
  NANDN U28180 ( .A(n23488), .B(n23489), .Z(n23487) );
  NAND U28181 ( .A(n23490), .B(n23491), .Z(n23489) );
  OR U28182 ( .A(n23491), .B(n23490), .Z(n23486) );
  IV U28183 ( .A(n23492), .Z(n23490) );
  XOR U28184 ( .A(n23467), .B(n23493), .Z(N28218) );
  XNOR U28185 ( .A(n23470), .B(n23469), .Z(n23493) );
  XNOR U28186 ( .A(n23481), .B(n23494), .Z(n23469) );
  XOR U28187 ( .A(n23485), .B(n23483), .Z(n23494) );
  XOR U28188 ( .A(n23491), .B(n23495), .Z(n23483) );
  XOR U28189 ( .A(n23488), .B(n23492), .Z(n23495) );
  NAND U28190 ( .A(n23496), .B(n23497), .Z(n23492) );
  NAND U28191 ( .A(n23498), .B(n23499), .Z(n23497) );
  NAND U28192 ( .A(n23500), .B(n23501), .Z(n23496) );
  AND U28193 ( .A(n23502), .B(n23503), .Z(n23488) );
  NAND U28194 ( .A(n23504), .B(n23505), .Z(n23503) );
  NAND U28195 ( .A(n23506), .B(n23507), .Z(n23502) );
  NANDN U28196 ( .A(n23508), .B(n23509), .Z(n23491) );
  NANDN U28197 ( .A(n23510), .B(n23511), .Z(n23485) );
  XNOR U28198 ( .A(n23476), .B(n23512), .Z(n23481) );
  XOR U28199 ( .A(n23474), .B(n23478), .Z(n23512) );
  NAND U28200 ( .A(n23513), .B(n23514), .Z(n23478) );
  NAND U28201 ( .A(n23515), .B(n23516), .Z(n23514) );
  NAND U28202 ( .A(n23517), .B(n23518), .Z(n23513) );
  AND U28203 ( .A(n23519), .B(n23520), .Z(n23474) );
  NAND U28204 ( .A(n23521), .B(n23522), .Z(n23520) );
  NAND U28205 ( .A(n23523), .B(n23524), .Z(n23519) );
  AND U28206 ( .A(n23525), .B(n23526), .Z(n23476) );
  NAND U28207 ( .A(n23527), .B(n23528), .Z(n23470) );
  XNOR U28208 ( .A(n23453), .B(n23529), .Z(n23467) );
  XOR U28209 ( .A(n23457), .B(n23455), .Z(n23529) );
  XOR U28210 ( .A(n23463), .B(n23530), .Z(n23455) );
  XOR U28211 ( .A(n23460), .B(n23464), .Z(n23530) );
  NAND U28212 ( .A(n23531), .B(n23532), .Z(n23464) );
  NAND U28213 ( .A(n23533), .B(n23534), .Z(n23532) );
  NAND U28214 ( .A(n23535), .B(n23536), .Z(n23531) );
  AND U28215 ( .A(n23537), .B(n23538), .Z(n23460) );
  NAND U28216 ( .A(n23539), .B(n23540), .Z(n23538) );
  NAND U28217 ( .A(n23541), .B(n23542), .Z(n23537) );
  NANDN U28218 ( .A(n23543), .B(n23544), .Z(n23463) );
  NANDN U28219 ( .A(n23545), .B(n23546), .Z(n23457) );
  XNOR U28220 ( .A(n23448), .B(n23547), .Z(n23453) );
  XOR U28221 ( .A(n23446), .B(n23450), .Z(n23547) );
  NAND U28222 ( .A(n23548), .B(n23549), .Z(n23450) );
  NAND U28223 ( .A(n23550), .B(n23551), .Z(n23549) );
  NAND U28224 ( .A(n23552), .B(n23553), .Z(n23548) );
  AND U28225 ( .A(n23554), .B(n23555), .Z(n23446) );
  NAND U28226 ( .A(n23556), .B(n23557), .Z(n23555) );
  NAND U28227 ( .A(n23558), .B(n23559), .Z(n23554) );
  AND U28228 ( .A(n23560), .B(n23561), .Z(n23448) );
  XOR U28229 ( .A(n23528), .B(n23527), .Z(N28217) );
  XNOR U28230 ( .A(n23546), .B(n23545), .Z(n23527) );
  XNOR U28231 ( .A(n23560), .B(n23561), .Z(n23545) );
  XOR U28232 ( .A(n23557), .B(n23556), .Z(n23561) );
  XOR U28233 ( .A(y[579]), .B(x[579]), .Z(n23556) );
  XOR U28234 ( .A(n23559), .B(n23558), .Z(n23557) );
  XOR U28235 ( .A(y[581]), .B(x[581]), .Z(n23558) );
  XOR U28236 ( .A(y[580]), .B(x[580]), .Z(n23559) );
  XOR U28237 ( .A(n23551), .B(n23550), .Z(n23560) );
  XOR U28238 ( .A(n23553), .B(n23552), .Z(n23550) );
  XOR U28239 ( .A(y[578]), .B(x[578]), .Z(n23552) );
  XOR U28240 ( .A(y[577]), .B(x[577]), .Z(n23553) );
  XOR U28241 ( .A(y[576]), .B(x[576]), .Z(n23551) );
  XNOR U28242 ( .A(n23544), .B(n23543), .Z(n23546) );
  XNOR U28243 ( .A(n23540), .B(n23539), .Z(n23543) );
  XOR U28244 ( .A(n23542), .B(n23541), .Z(n23539) );
  XOR U28245 ( .A(y[575]), .B(x[575]), .Z(n23541) );
  XOR U28246 ( .A(y[574]), .B(x[574]), .Z(n23542) );
  XOR U28247 ( .A(y[573]), .B(x[573]), .Z(n23540) );
  XOR U28248 ( .A(n23534), .B(n23533), .Z(n23544) );
  XOR U28249 ( .A(n23536), .B(n23535), .Z(n23533) );
  XOR U28250 ( .A(y[572]), .B(x[572]), .Z(n23535) );
  XOR U28251 ( .A(y[571]), .B(x[571]), .Z(n23536) );
  XOR U28252 ( .A(y[570]), .B(x[570]), .Z(n23534) );
  XNOR U28253 ( .A(n23511), .B(n23510), .Z(n23528) );
  XNOR U28254 ( .A(n23525), .B(n23526), .Z(n23510) );
  XOR U28255 ( .A(n23522), .B(n23521), .Z(n23526) );
  XOR U28256 ( .A(y[567]), .B(x[567]), .Z(n23521) );
  XOR U28257 ( .A(n23524), .B(n23523), .Z(n23522) );
  XOR U28258 ( .A(y[569]), .B(x[569]), .Z(n23523) );
  XOR U28259 ( .A(y[568]), .B(x[568]), .Z(n23524) );
  XOR U28260 ( .A(n23516), .B(n23515), .Z(n23525) );
  XOR U28261 ( .A(n23518), .B(n23517), .Z(n23515) );
  XOR U28262 ( .A(y[566]), .B(x[566]), .Z(n23517) );
  XOR U28263 ( .A(y[565]), .B(x[565]), .Z(n23518) );
  XOR U28264 ( .A(y[564]), .B(x[564]), .Z(n23516) );
  XNOR U28265 ( .A(n23509), .B(n23508), .Z(n23511) );
  XNOR U28266 ( .A(n23505), .B(n23504), .Z(n23508) );
  XOR U28267 ( .A(n23507), .B(n23506), .Z(n23504) );
  XOR U28268 ( .A(y[563]), .B(x[563]), .Z(n23506) );
  XOR U28269 ( .A(y[562]), .B(x[562]), .Z(n23507) );
  XOR U28270 ( .A(y[561]), .B(x[561]), .Z(n23505) );
  XOR U28271 ( .A(n23499), .B(n23498), .Z(n23509) );
  XOR U28272 ( .A(n23501), .B(n23500), .Z(n23498) );
  XOR U28273 ( .A(y[560]), .B(x[560]), .Z(n23500) );
  XOR U28274 ( .A(y[559]), .B(x[559]), .Z(n23501) );
  XOR U28275 ( .A(y[558]), .B(x[558]), .Z(n23499) );
  NAND U28276 ( .A(n23562), .B(n23563), .Z(N28209) );
  NAND U28277 ( .A(n23564), .B(n23565), .Z(n23563) );
  NANDN U28278 ( .A(n23566), .B(n23567), .Z(n23565) );
  NANDN U28279 ( .A(n23567), .B(n23566), .Z(n23562) );
  XOR U28280 ( .A(n23566), .B(n23568), .Z(N28208) );
  XNOR U28281 ( .A(n23564), .B(n23567), .Z(n23568) );
  NAND U28282 ( .A(n23569), .B(n23570), .Z(n23567) );
  NAND U28283 ( .A(n23571), .B(n23572), .Z(n23570) );
  NANDN U28284 ( .A(n23573), .B(n23574), .Z(n23572) );
  NANDN U28285 ( .A(n23574), .B(n23573), .Z(n23569) );
  AND U28286 ( .A(n23575), .B(n23576), .Z(n23564) );
  NAND U28287 ( .A(n23577), .B(n23578), .Z(n23576) );
  OR U28288 ( .A(n23579), .B(n23580), .Z(n23578) );
  NAND U28289 ( .A(n23580), .B(n23579), .Z(n23575) );
  IV U28290 ( .A(n23581), .Z(n23580) );
  AND U28291 ( .A(n23582), .B(n23583), .Z(n23566) );
  NAND U28292 ( .A(n23584), .B(n23585), .Z(n23583) );
  NANDN U28293 ( .A(n23586), .B(n23587), .Z(n23585) );
  NANDN U28294 ( .A(n23587), .B(n23586), .Z(n23582) );
  XOR U28295 ( .A(n23579), .B(n23588), .Z(N28207) );
  XOR U28296 ( .A(n23577), .B(n23581), .Z(n23588) );
  XNOR U28297 ( .A(n23574), .B(n23589), .Z(n23581) );
  XNOR U28298 ( .A(n23571), .B(n23573), .Z(n23589) );
  AND U28299 ( .A(n23590), .B(n23591), .Z(n23573) );
  NANDN U28300 ( .A(n23592), .B(n23593), .Z(n23591) );
  NANDN U28301 ( .A(n23594), .B(n23595), .Z(n23593) );
  IV U28302 ( .A(n23596), .Z(n23595) );
  NAND U28303 ( .A(n23596), .B(n23594), .Z(n23590) );
  AND U28304 ( .A(n23597), .B(n23598), .Z(n23571) );
  NAND U28305 ( .A(n23599), .B(n23600), .Z(n23598) );
  OR U28306 ( .A(n23601), .B(n23602), .Z(n23600) );
  NAND U28307 ( .A(n23602), .B(n23601), .Z(n23597) );
  IV U28308 ( .A(n23603), .Z(n23602) );
  NAND U28309 ( .A(n23604), .B(n23605), .Z(n23574) );
  NANDN U28310 ( .A(n23606), .B(n23607), .Z(n23605) );
  NAND U28311 ( .A(n23608), .B(n23609), .Z(n23607) );
  OR U28312 ( .A(n23609), .B(n23608), .Z(n23604) );
  IV U28313 ( .A(n23610), .Z(n23608) );
  AND U28314 ( .A(n23611), .B(n23612), .Z(n23577) );
  NAND U28315 ( .A(n23613), .B(n23614), .Z(n23612) );
  NANDN U28316 ( .A(n23615), .B(n23616), .Z(n23614) );
  NANDN U28317 ( .A(n23616), .B(n23615), .Z(n23611) );
  XOR U28318 ( .A(n23587), .B(n23617), .Z(n23579) );
  XNOR U28319 ( .A(n23584), .B(n23586), .Z(n23617) );
  AND U28320 ( .A(n23618), .B(n23619), .Z(n23586) );
  NANDN U28321 ( .A(n23620), .B(n23621), .Z(n23619) );
  NANDN U28322 ( .A(n23622), .B(n23623), .Z(n23621) );
  IV U28323 ( .A(n23624), .Z(n23623) );
  NAND U28324 ( .A(n23624), .B(n23622), .Z(n23618) );
  AND U28325 ( .A(n23625), .B(n23626), .Z(n23584) );
  NAND U28326 ( .A(n23627), .B(n23628), .Z(n23626) );
  OR U28327 ( .A(n23629), .B(n23630), .Z(n23628) );
  NAND U28328 ( .A(n23630), .B(n23629), .Z(n23625) );
  IV U28329 ( .A(n23631), .Z(n23630) );
  NAND U28330 ( .A(n23632), .B(n23633), .Z(n23587) );
  NANDN U28331 ( .A(n23634), .B(n23635), .Z(n23633) );
  NAND U28332 ( .A(n23636), .B(n23637), .Z(n23635) );
  OR U28333 ( .A(n23637), .B(n23636), .Z(n23632) );
  IV U28334 ( .A(n23638), .Z(n23636) );
  XOR U28335 ( .A(n23613), .B(n23639), .Z(N28206) );
  XNOR U28336 ( .A(n23616), .B(n23615), .Z(n23639) );
  XNOR U28337 ( .A(n23627), .B(n23640), .Z(n23615) );
  XOR U28338 ( .A(n23631), .B(n23629), .Z(n23640) );
  XOR U28339 ( .A(n23637), .B(n23641), .Z(n23629) );
  XOR U28340 ( .A(n23634), .B(n23638), .Z(n23641) );
  NAND U28341 ( .A(n23642), .B(n23643), .Z(n23638) );
  NAND U28342 ( .A(n23644), .B(n23645), .Z(n23643) );
  NAND U28343 ( .A(n23646), .B(n23647), .Z(n23642) );
  AND U28344 ( .A(n23648), .B(n23649), .Z(n23634) );
  NAND U28345 ( .A(n23650), .B(n23651), .Z(n23649) );
  NAND U28346 ( .A(n23652), .B(n23653), .Z(n23648) );
  NANDN U28347 ( .A(n23654), .B(n23655), .Z(n23637) );
  NANDN U28348 ( .A(n23656), .B(n23657), .Z(n23631) );
  XNOR U28349 ( .A(n23622), .B(n23658), .Z(n23627) );
  XOR U28350 ( .A(n23620), .B(n23624), .Z(n23658) );
  NAND U28351 ( .A(n23659), .B(n23660), .Z(n23624) );
  NAND U28352 ( .A(n23661), .B(n23662), .Z(n23660) );
  NAND U28353 ( .A(n23663), .B(n23664), .Z(n23659) );
  AND U28354 ( .A(n23665), .B(n23666), .Z(n23620) );
  NAND U28355 ( .A(n23667), .B(n23668), .Z(n23666) );
  NAND U28356 ( .A(n23669), .B(n23670), .Z(n23665) );
  AND U28357 ( .A(n23671), .B(n23672), .Z(n23622) );
  NAND U28358 ( .A(n23673), .B(n23674), .Z(n23616) );
  XNOR U28359 ( .A(n23599), .B(n23675), .Z(n23613) );
  XOR U28360 ( .A(n23603), .B(n23601), .Z(n23675) );
  XOR U28361 ( .A(n23609), .B(n23676), .Z(n23601) );
  XOR U28362 ( .A(n23606), .B(n23610), .Z(n23676) );
  NAND U28363 ( .A(n23677), .B(n23678), .Z(n23610) );
  NAND U28364 ( .A(n23679), .B(n23680), .Z(n23678) );
  NAND U28365 ( .A(n23681), .B(n23682), .Z(n23677) );
  AND U28366 ( .A(n23683), .B(n23684), .Z(n23606) );
  NAND U28367 ( .A(n23685), .B(n23686), .Z(n23684) );
  NAND U28368 ( .A(n23687), .B(n23688), .Z(n23683) );
  NANDN U28369 ( .A(n23689), .B(n23690), .Z(n23609) );
  NANDN U28370 ( .A(n23691), .B(n23692), .Z(n23603) );
  XNOR U28371 ( .A(n23594), .B(n23693), .Z(n23599) );
  XOR U28372 ( .A(n23592), .B(n23596), .Z(n23693) );
  NAND U28373 ( .A(n23694), .B(n23695), .Z(n23596) );
  NAND U28374 ( .A(n23696), .B(n23697), .Z(n23695) );
  NAND U28375 ( .A(n23698), .B(n23699), .Z(n23694) );
  AND U28376 ( .A(n23700), .B(n23701), .Z(n23592) );
  NAND U28377 ( .A(n23702), .B(n23703), .Z(n23701) );
  NAND U28378 ( .A(n23704), .B(n23705), .Z(n23700) );
  AND U28379 ( .A(n23706), .B(n23707), .Z(n23594) );
  XOR U28380 ( .A(n23674), .B(n23673), .Z(N28205) );
  XNOR U28381 ( .A(n23692), .B(n23691), .Z(n23673) );
  XNOR U28382 ( .A(n23706), .B(n23707), .Z(n23691) );
  XOR U28383 ( .A(n23703), .B(n23702), .Z(n23707) );
  XOR U28384 ( .A(y[555]), .B(x[555]), .Z(n23702) );
  XOR U28385 ( .A(n23705), .B(n23704), .Z(n23703) );
  XOR U28386 ( .A(y[557]), .B(x[557]), .Z(n23704) );
  XOR U28387 ( .A(y[556]), .B(x[556]), .Z(n23705) );
  XOR U28388 ( .A(n23697), .B(n23696), .Z(n23706) );
  XOR U28389 ( .A(n23699), .B(n23698), .Z(n23696) );
  XOR U28390 ( .A(y[554]), .B(x[554]), .Z(n23698) );
  XOR U28391 ( .A(y[553]), .B(x[553]), .Z(n23699) );
  XOR U28392 ( .A(y[552]), .B(x[552]), .Z(n23697) );
  XNOR U28393 ( .A(n23690), .B(n23689), .Z(n23692) );
  XNOR U28394 ( .A(n23686), .B(n23685), .Z(n23689) );
  XOR U28395 ( .A(n23688), .B(n23687), .Z(n23685) );
  XOR U28396 ( .A(y[551]), .B(x[551]), .Z(n23687) );
  XOR U28397 ( .A(y[550]), .B(x[550]), .Z(n23688) );
  XOR U28398 ( .A(y[549]), .B(x[549]), .Z(n23686) );
  XOR U28399 ( .A(n23680), .B(n23679), .Z(n23690) );
  XOR U28400 ( .A(n23682), .B(n23681), .Z(n23679) );
  XOR U28401 ( .A(y[548]), .B(x[548]), .Z(n23681) );
  XOR U28402 ( .A(y[547]), .B(x[547]), .Z(n23682) );
  XOR U28403 ( .A(y[546]), .B(x[546]), .Z(n23680) );
  XNOR U28404 ( .A(n23657), .B(n23656), .Z(n23674) );
  XNOR U28405 ( .A(n23671), .B(n23672), .Z(n23656) );
  XOR U28406 ( .A(n23668), .B(n23667), .Z(n23672) );
  XOR U28407 ( .A(y[543]), .B(x[543]), .Z(n23667) );
  XOR U28408 ( .A(n23670), .B(n23669), .Z(n23668) );
  XOR U28409 ( .A(y[545]), .B(x[545]), .Z(n23669) );
  XOR U28410 ( .A(y[544]), .B(x[544]), .Z(n23670) );
  XOR U28411 ( .A(n23662), .B(n23661), .Z(n23671) );
  XOR U28412 ( .A(n23664), .B(n23663), .Z(n23661) );
  XOR U28413 ( .A(y[542]), .B(x[542]), .Z(n23663) );
  XOR U28414 ( .A(y[541]), .B(x[541]), .Z(n23664) );
  XOR U28415 ( .A(y[540]), .B(x[540]), .Z(n23662) );
  XNOR U28416 ( .A(n23655), .B(n23654), .Z(n23657) );
  XNOR U28417 ( .A(n23651), .B(n23650), .Z(n23654) );
  XOR U28418 ( .A(n23653), .B(n23652), .Z(n23650) );
  XOR U28419 ( .A(y[539]), .B(x[539]), .Z(n23652) );
  XOR U28420 ( .A(y[538]), .B(x[538]), .Z(n23653) );
  XOR U28421 ( .A(y[537]), .B(x[537]), .Z(n23651) );
  XOR U28422 ( .A(n23645), .B(n23644), .Z(n23655) );
  XOR U28423 ( .A(n23647), .B(n23646), .Z(n23644) );
  XOR U28424 ( .A(y[536]), .B(x[536]), .Z(n23646) );
  XOR U28425 ( .A(y[535]), .B(x[535]), .Z(n23647) );
  XOR U28426 ( .A(y[534]), .B(x[534]), .Z(n23645) );
  NAND U28427 ( .A(n23708), .B(n23709), .Z(N28197) );
  NAND U28428 ( .A(n23710), .B(n23711), .Z(n23709) );
  NANDN U28429 ( .A(n23712), .B(n23713), .Z(n23711) );
  NANDN U28430 ( .A(n23713), .B(n23712), .Z(n23708) );
  XOR U28431 ( .A(n23712), .B(n23714), .Z(N28196) );
  XNOR U28432 ( .A(n23710), .B(n23713), .Z(n23714) );
  NAND U28433 ( .A(n23715), .B(n23716), .Z(n23713) );
  NAND U28434 ( .A(n23717), .B(n23718), .Z(n23716) );
  NANDN U28435 ( .A(n23719), .B(n23720), .Z(n23718) );
  NANDN U28436 ( .A(n23720), .B(n23719), .Z(n23715) );
  AND U28437 ( .A(n23721), .B(n23722), .Z(n23710) );
  NAND U28438 ( .A(n23723), .B(n23724), .Z(n23722) );
  OR U28439 ( .A(n23725), .B(n23726), .Z(n23724) );
  NAND U28440 ( .A(n23726), .B(n23725), .Z(n23721) );
  IV U28441 ( .A(n23727), .Z(n23726) );
  AND U28442 ( .A(n23728), .B(n23729), .Z(n23712) );
  NAND U28443 ( .A(n23730), .B(n23731), .Z(n23729) );
  NANDN U28444 ( .A(n23732), .B(n23733), .Z(n23731) );
  NANDN U28445 ( .A(n23733), .B(n23732), .Z(n23728) );
  XOR U28446 ( .A(n23725), .B(n23734), .Z(N28195) );
  XOR U28447 ( .A(n23723), .B(n23727), .Z(n23734) );
  XNOR U28448 ( .A(n23720), .B(n23735), .Z(n23727) );
  XNOR U28449 ( .A(n23717), .B(n23719), .Z(n23735) );
  AND U28450 ( .A(n23736), .B(n23737), .Z(n23719) );
  NANDN U28451 ( .A(n23738), .B(n23739), .Z(n23737) );
  NANDN U28452 ( .A(n23740), .B(n23741), .Z(n23739) );
  IV U28453 ( .A(n23742), .Z(n23741) );
  NAND U28454 ( .A(n23742), .B(n23740), .Z(n23736) );
  AND U28455 ( .A(n23743), .B(n23744), .Z(n23717) );
  NAND U28456 ( .A(n23745), .B(n23746), .Z(n23744) );
  OR U28457 ( .A(n23747), .B(n23748), .Z(n23746) );
  NAND U28458 ( .A(n23748), .B(n23747), .Z(n23743) );
  IV U28459 ( .A(n23749), .Z(n23748) );
  NAND U28460 ( .A(n23750), .B(n23751), .Z(n23720) );
  NANDN U28461 ( .A(n23752), .B(n23753), .Z(n23751) );
  NAND U28462 ( .A(n23754), .B(n23755), .Z(n23753) );
  OR U28463 ( .A(n23755), .B(n23754), .Z(n23750) );
  IV U28464 ( .A(n23756), .Z(n23754) );
  AND U28465 ( .A(n23757), .B(n23758), .Z(n23723) );
  NAND U28466 ( .A(n23759), .B(n23760), .Z(n23758) );
  NANDN U28467 ( .A(n23761), .B(n23762), .Z(n23760) );
  NANDN U28468 ( .A(n23762), .B(n23761), .Z(n23757) );
  XOR U28469 ( .A(n23733), .B(n23763), .Z(n23725) );
  XNOR U28470 ( .A(n23730), .B(n23732), .Z(n23763) );
  AND U28471 ( .A(n23764), .B(n23765), .Z(n23732) );
  NANDN U28472 ( .A(n23766), .B(n23767), .Z(n23765) );
  NANDN U28473 ( .A(n23768), .B(n23769), .Z(n23767) );
  IV U28474 ( .A(n23770), .Z(n23769) );
  NAND U28475 ( .A(n23770), .B(n23768), .Z(n23764) );
  AND U28476 ( .A(n23771), .B(n23772), .Z(n23730) );
  NAND U28477 ( .A(n23773), .B(n23774), .Z(n23772) );
  OR U28478 ( .A(n23775), .B(n23776), .Z(n23774) );
  NAND U28479 ( .A(n23776), .B(n23775), .Z(n23771) );
  IV U28480 ( .A(n23777), .Z(n23776) );
  NAND U28481 ( .A(n23778), .B(n23779), .Z(n23733) );
  NANDN U28482 ( .A(n23780), .B(n23781), .Z(n23779) );
  NAND U28483 ( .A(n23782), .B(n23783), .Z(n23781) );
  OR U28484 ( .A(n23783), .B(n23782), .Z(n23778) );
  IV U28485 ( .A(n23784), .Z(n23782) );
  XOR U28486 ( .A(n23759), .B(n23785), .Z(N28194) );
  XNOR U28487 ( .A(n23762), .B(n23761), .Z(n23785) );
  XNOR U28488 ( .A(n23773), .B(n23786), .Z(n23761) );
  XOR U28489 ( .A(n23777), .B(n23775), .Z(n23786) );
  XOR U28490 ( .A(n23783), .B(n23787), .Z(n23775) );
  XOR U28491 ( .A(n23780), .B(n23784), .Z(n23787) );
  NAND U28492 ( .A(n23788), .B(n23789), .Z(n23784) );
  NAND U28493 ( .A(n23790), .B(n23791), .Z(n23789) );
  NAND U28494 ( .A(n23792), .B(n23793), .Z(n23788) );
  AND U28495 ( .A(n23794), .B(n23795), .Z(n23780) );
  NAND U28496 ( .A(n23796), .B(n23797), .Z(n23795) );
  NAND U28497 ( .A(n23798), .B(n23799), .Z(n23794) );
  NANDN U28498 ( .A(n23800), .B(n23801), .Z(n23783) );
  NANDN U28499 ( .A(n23802), .B(n23803), .Z(n23777) );
  XNOR U28500 ( .A(n23768), .B(n23804), .Z(n23773) );
  XOR U28501 ( .A(n23766), .B(n23770), .Z(n23804) );
  NAND U28502 ( .A(n23805), .B(n23806), .Z(n23770) );
  NAND U28503 ( .A(n23807), .B(n23808), .Z(n23806) );
  NAND U28504 ( .A(n23809), .B(n23810), .Z(n23805) );
  AND U28505 ( .A(n23811), .B(n23812), .Z(n23766) );
  NAND U28506 ( .A(n23813), .B(n23814), .Z(n23812) );
  NAND U28507 ( .A(n23815), .B(n23816), .Z(n23811) );
  AND U28508 ( .A(n23817), .B(n23818), .Z(n23768) );
  NAND U28509 ( .A(n23819), .B(n23820), .Z(n23762) );
  XNOR U28510 ( .A(n23745), .B(n23821), .Z(n23759) );
  XOR U28511 ( .A(n23749), .B(n23747), .Z(n23821) );
  XOR U28512 ( .A(n23755), .B(n23822), .Z(n23747) );
  XOR U28513 ( .A(n23752), .B(n23756), .Z(n23822) );
  NAND U28514 ( .A(n23823), .B(n23824), .Z(n23756) );
  NAND U28515 ( .A(n23825), .B(n23826), .Z(n23824) );
  NAND U28516 ( .A(n23827), .B(n23828), .Z(n23823) );
  AND U28517 ( .A(n23829), .B(n23830), .Z(n23752) );
  NAND U28518 ( .A(n23831), .B(n23832), .Z(n23830) );
  NAND U28519 ( .A(n23833), .B(n23834), .Z(n23829) );
  NANDN U28520 ( .A(n23835), .B(n23836), .Z(n23755) );
  NANDN U28521 ( .A(n23837), .B(n23838), .Z(n23749) );
  XNOR U28522 ( .A(n23740), .B(n23839), .Z(n23745) );
  XOR U28523 ( .A(n23738), .B(n23742), .Z(n23839) );
  NAND U28524 ( .A(n23840), .B(n23841), .Z(n23742) );
  NAND U28525 ( .A(n23842), .B(n23843), .Z(n23841) );
  NAND U28526 ( .A(n23844), .B(n23845), .Z(n23840) );
  AND U28527 ( .A(n23846), .B(n23847), .Z(n23738) );
  NAND U28528 ( .A(n23848), .B(n23849), .Z(n23847) );
  NAND U28529 ( .A(n23850), .B(n23851), .Z(n23846) );
  AND U28530 ( .A(n23852), .B(n23853), .Z(n23740) );
  XOR U28531 ( .A(n23820), .B(n23819), .Z(N28193) );
  XNOR U28532 ( .A(n23838), .B(n23837), .Z(n23819) );
  XNOR U28533 ( .A(n23852), .B(n23853), .Z(n23837) );
  XOR U28534 ( .A(n23849), .B(n23848), .Z(n23853) );
  XOR U28535 ( .A(y[531]), .B(x[531]), .Z(n23848) );
  XOR U28536 ( .A(n23851), .B(n23850), .Z(n23849) );
  XOR U28537 ( .A(y[533]), .B(x[533]), .Z(n23850) );
  XOR U28538 ( .A(y[532]), .B(x[532]), .Z(n23851) );
  XOR U28539 ( .A(n23843), .B(n23842), .Z(n23852) );
  XOR U28540 ( .A(n23845), .B(n23844), .Z(n23842) );
  XOR U28541 ( .A(y[530]), .B(x[530]), .Z(n23844) );
  XOR U28542 ( .A(y[529]), .B(x[529]), .Z(n23845) );
  XOR U28543 ( .A(y[528]), .B(x[528]), .Z(n23843) );
  XNOR U28544 ( .A(n23836), .B(n23835), .Z(n23838) );
  XNOR U28545 ( .A(n23832), .B(n23831), .Z(n23835) );
  XOR U28546 ( .A(n23834), .B(n23833), .Z(n23831) );
  XOR U28547 ( .A(y[527]), .B(x[527]), .Z(n23833) );
  XOR U28548 ( .A(y[526]), .B(x[526]), .Z(n23834) );
  XOR U28549 ( .A(y[525]), .B(x[525]), .Z(n23832) );
  XOR U28550 ( .A(n23826), .B(n23825), .Z(n23836) );
  XOR U28551 ( .A(n23828), .B(n23827), .Z(n23825) );
  XOR U28552 ( .A(y[524]), .B(x[524]), .Z(n23827) );
  XOR U28553 ( .A(y[523]), .B(x[523]), .Z(n23828) );
  XOR U28554 ( .A(y[522]), .B(x[522]), .Z(n23826) );
  XNOR U28555 ( .A(n23803), .B(n23802), .Z(n23820) );
  XNOR U28556 ( .A(n23817), .B(n23818), .Z(n23802) );
  XOR U28557 ( .A(n23814), .B(n23813), .Z(n23818) );
  XOR U28558 ( .A(y[519]), .B(x[519]), .Z(n23813) );
  XOR U28559 ( .A(n23816), .B(n23815), .Z(n23814) );
  XOR U28560 ( .A(y[521]), .B(x[521]), .Z(n23815) );
  XOR U28561 ( .A(y[520]), .B(x[520]), .Z(n23816) );
  XOR U28562 ( .A(n23808), .B(n23807), .Z(n23817) );
  XOR U28563 ( .A(n23810), .B(n23809), .Z(n23807) );
  XOR U28564 ( .A(y[518]), .B(x[518]), .Z(n23809) );
  XOR U28565 ( .A(y[517]), .B(x[517]), .Z(n23810) );
  XOR U28566 ( .A(y[516]), .B(x[516]), .Z(n23808) );
  XNOR U28567 ( .A(n23801), .B(n23800), .Z(n23803) );
  XNOR U28568 ( .A(n23797), .B(n23796), .Z(n23800) );
  XOR U28569 ( .A(n23799), .B(n23798), .Z(n23796) );
  XOR U28570 ( .A(y[515]), .B(x[515]), .Z(n23798) );
  XOR U28571 ( .A(y[514]), .B(x[514]), .Z(n23799) );
  XOR U28572 ( .A(y[513]), .B(x[513]), .Z(n23797) );
  XOR U28573 ( .A(n23791), .B(n23790), .Z(n23801) );
  XOR U28574 ( .A(n23793), .B(n23792), .Z(n23790) );
  XOR U28575 ( .A(y[512]), .B(x[512]), .Z(n23792) );
  XOR U28576 ( .A(y[511]), .B(x[511]), .Z(n23793) );
  XOR U28577 ( .A(y[510]), .B(x[510]), .Z(n23791) );
  NAND U28578 ( .A(n23854), .B(n23855), .Z(N28185) );
  NAND U28579 ( .A(n23856), .B(n23857), .Z(n23855) );
  NANDN U28580 ( .A(n23858), .B(n23859), .Z(n23857) );
  NANDN U28581 ( .A(n23859), .B(n23858), .Z(n23854) );
  XOR U28582 ( .A(n23858), .B(n23860), .Z(N28184) );
  XNOR U28583 ( .A(n23856), .B(n23859), .Z(n23860) );
  NAND U28584 ( .A(n23861), .B(n23862), .Z(n23859) );
  NAND U28585 ( .A(n23863), .B(n23864), .Z(n23862) );
  NANDN U28586 ( .A(n23865), .B(n23866), .Z(n23864) );
  NANDN U28587 ( .A(n23866), .B(n23865), .Z(n23861) );
  AND U28588 ( .A(n23867), .B(n23868), .Z(n23856) );
  NAND U28589 ( .A(n23869), .B(n23870), .Z(n23868) );
  OR U28590 ( .A(n23871), .B(n23872), .Z(n23870) );
  NAND U28591 ( .A(n23872), .B(n23871), .Z(n23867) );
  IV U28592 ( .A(n23873), .Z(n23872) );
  AND U28593 ( .A(n23874), .B(n23875), .Z(n23858) );
  NAND U28594 ( .A(n23876), .B(n23877), .Z(n23875) );
  NANDN U28595 ( .A(n23878), .B(n23879), .Z(n23877) );
  NANDN U28596 ( .A(n23879), .B(n23878), .Z(n23874) );
  XOR U28597 ( .A(n23871), .B(n23880), .Z(N28183) );
  XOR U28598 ( .A(n23869), .B(n23873), .Z(n23880) );
  XNOR U28599 ( .A(n23866), .B(n23881), .Z(n23873) );
  XNOR U28600 ( .A(n23863), .B(n23865), .Z(n23881) );
  AND U28601 ( .A(n23882), .B(n23883), .Z(n23865) );
  NANDN U28602 ( .A(n23884), .B(n23885), .Z(n23883) );
  NANDN U28603 ( .A(n23886), .B(n23887), .Z(n23885) );
  IV U28604 ( .A(n23888), .Z(n23887) );
  NAND U28605 ( .A(n23888), .B(n23886), .Z(n23882) );
  AND U28606 ( .A(n23889), .B(n23890), .Z(n23863) );
  NAND U28607 ( .A(n23891), .B(n23892), .Z(n23890) );
  OR U28608 ( .A(n23893), .B(n23894), .Z(n23892) );
  NAND U28609 ( .A(n23894), .B(n23893), .Z(n23889) );
  IV U28610 ( .A(n23895), .Z(n23894) );
  NAND U28611 ( .A(n23896), .B(n23897), .Z(n23866) );
  NANDN U28612 ( .A(n23898), .B(n23899), .Z(n23897) );
  NAND U28613 ( .A(n23900), .B(n23901), .Z(n23899) );
  OR U28614 ( .A(n23901), .B(n23900), .Z(n23896) );
  IV U28615 ( .A(n23902), .Z(n23900) );
  AND U28616 ( .A(n23903), .B(n23904), .Z(n23869) );
  NAND U28617 ( .A(n23905), .B(n23906), .Z(n23904) );
  NANDN U28618 ( .A(n23907), .B(n23908), .Z(n23906) );
  NANDN U28619 ( .A(n23908), .B(n23907), .Z(n23903) );
  XOR U28620 ( .A(n23879), .B(n23909), .Z(n23871) );
  XNOR U28621 ( .A(n23876), .B(n23878), .Z(n23909) );
  AND U28622 ( .A(n23910), .B(n23911), .Z(n23878) );
  NANDN U28623 ( .A(n23912), .B(n23913), .Z(n23911) );
  NANDN U28624 ( .A(n23914), .B(n23915), .Z(n23913) );
  IV U28625 ( .A(n23916), .Z(n23915) );
  NAND U28626 ( .A(n23916), .B(n23914), .Z(n23910) );
  AND U28627 ( .A(n23917), .B(n23918), .Z(n23876) );
  NAND U28628 ( .A(n23919), .B(n23920), .Z(n23918) );
  OR U28629 ( .A(n23921), .B(n23922), .Z(n23920) );
  NAND U28630 ( .A(n23922), .B(n23921), .Z(n23917) );
  IV U28631 ( .A(n23923), .Z(n23922) );
  NAND U28632 ( .A(n23924), .B(n23925), .Z(n23879) );
  NANDN U28633 ( .A(n23926), .B(n23927), .Z(n23925) );
  NAND U28634 ( .A(n23928), .B(n23929), .Z(n23927) );
  OR U28635 ( .A(n23929), .B(n23928), .Z(n23924) );
  IV U28636 ( .A(n23930), .Z(n23928) );
  XOR U28637 ( .A(n23905), .B(n23931), .Z(N28182) );
  XNOR U28638 ( .A(n23908), .B(n23907), .Z(n23931) );
  XNOR U28639 ( .A(n23919), .B(n23932), .Z(n23907) );
  XOR U28640 ( .A(n23923), .B(n23921), .Z(n23932) );
  XOR U28641 ( .A(n23929), .B(n23933), .Z(n23921) );
  XOR U28642 ( .A(n23926), .B(n23930), .Z(n23933) );
  NAND U28643 ( .A(n23934), .B(n23935), .Z(n23930) );
  NAND U28644 ( .A(n23936), .B(n23937), .Z(n23935) );
  NAND U28645 ( .A(n23938), .B(n23939), .Z(n23934) );
  AND U28646 ( .A(n23940), .B(n23941), .Z(n23926) );
  NAND U28647 ( .A(n23942), .B(n23943), .Z(n23941) );
  NAND U28648 ( .A(n23944), .B(n23945), .Z(n23940) );
  NANDN U28649 ( .A(n23946), .B(n23947), .Z(n23929) );
  NANDN U28650 ( .A(n23948), .B(n23949), .Z(n23923) );
  XNOR U28651 ( .A(n23914), .B(n23950), .Z(n23919) );
  XOR U28652 ( .A(n23912), .B(n23916), .Z(n23950) );
  NAND U28653 ( .A(n23951), .B(n23952), .Z(n23916) );
  NAND U28654 ( .A(n23953), .B(n23954), .Z(n23952) );
  NAND U28655 ( .A(n23955), .B(n23956), .Z(n23951) );
  AND U28656 ( .A(n23957), .B(n23958), .Z(n23912) );
  NAND U28657 ( .A(n23959), .B(n23960), .Z(n23958) );
  NAND U28658 ( .A(n23961), .B(n23962), .Z(n23957) );
  AND U28659 ( .A(n23963), .B(n23964), .Z(n23914) );
  NAND U28660 ( .A(n23965), .B(n23966), .Z(n23908) );
  XNOR U28661 ( .A(n23891), .B(n23967), .Z(n23905) );
  XOR U28662 ( .A(n23895), .B(n23893), .Z(n23967) );
  XOR U28663 ( .A(n23901), .B(n23968), .Z(n23893) );
  XOR U28664 ( .A(n23898), .B(n23902), .Z(n23968) );
  NAND U28665 ( .A(n23969), .B(n23970), .Z(n23902) );
  NAND U28666 ( .A(n23971), .B(n23972), .Z(n23970) );
  NAND U28667 ( .A(n23973), .B(n23974), .Z(n23969) );
  AND U28668 ( .A(n23975), .B(n23976), .Z(n23898) );
  NAND U28669 ( .A(n23977), .B(n23978), .Z(n23976) );
  NAND U28670 ( .A(n23979), .B(n23980), .Z(n23975) );
  NANDN U28671 ( .A(n23981), .B(n23982), .Z(n23901) );
  NANDN U28672 ( .A(n23983), .B(n23984), .Z(n23895) );
  XNOR U28673 ( .A(n23886), .B(n23985), .Z(n23891) );
  XOR U28674 ( .A(n23884), .B(n23888), .Z(n23985) );
  NAND U28675 ( .A(n23986), .B(n23987), .Z(n23888) );
  NAND U28676 ( .A(n23988), .B(n23989), .Z(n23987) );
  NAND U28677 ( .A(n23990), .B(n23991), .Z(n23986) );
  AND U28678 ( .A(n23992), .B(n23993), .Z(n23884) );
  NAND U28679 ( .A(n23994), .B(n23995), .Z(n23993) );
  NAND U28680 ( .A(n23996), .B(n23997), .Z(n23992) );
  AND U28681 ( .A(n23998), .B(n23999), .Z(n23886) );
  XOR U28682 ( .A(n23966), .B(n23965), .Z(N28181) );
  XNOR U28683 ( .A(n23984), .B(n23983), .Z(n23965) );
  XNOR U28684 ( .A(n23998), .B(n23999), .Z(n23983) );
  XOR U28685 ( .A(n23995), .B(n23994), .Z(n23999) );
  XOR U28686 ( .A(y[507]), .B(x[507]), .Z(n23994) );
  XOR U28687 ( .A(n23997), .B(n23996), .Z(n23995) );
  XOR U28688 ( .A(y[509]), .B(x[509]), .Z(n23996) );
  XOR U28689 ( .A(y[508]), .B(x[508]), .Z(n23997) );
  XOR U28690 ( .A(n23989), .B(n23988), .Z(n23998) );
  XOR U28691 ( .A(n23991), .B(n23990), .Z(n23988) );
  XOR U28692 ( .A(y[506]), .B(x[506]), .Z(n23990) );
  XOR U28693 ( .A(y[505]), .B(x[505]), .Z(n23991) );
  XOR U28694 ( .A(y[504]), .B(x[504]), .Z(n23989) );
  XNOR U28695 ( .A(n23982), .B(n23981), .Z(n23984) );
  XNOR U28696 ( .A(n23978), .B(n23977), .Z(n23981) );
  XOR U28697 ( .A(n23980), .B(n23979), .Z(n23977) );
  XOR U28698 ( .A(y[503]), .B(x[503]), .Z(n23979) );
  XOR U28699 ( .A(y[502]), .B(x[502]), .Z(n23980) );
  XOR U28700 ( .A(y[501]), .B(x[501]), .Z(n23978) );
  XOR U28701 ( .A(n23972), .B(n23971), .Z(n23982) );
  XOR U28702 ( .A(n23974), .B(n23973), .Z(n23971) );
  XOR U28703 ( .A(y[500]), .B(x[500]), .Z(n23973) );
  XOR U28704 ( .A(y[499]), .B(x[499]), .Z(n23974) );
  XOR U28705 ( .A(y[498]), .B(x[498]), .Z(n23972) );
  XNOR U28706 ( .A(n23949), .B(n23948), .Z(n23966) );
  XNOR U28707 ( .A(n23963), .B(n23964), .Z(n23948) );
  XOR U28708 ( .A(n23960), .B(n23959), .Z(n23964) );
  XOR U28709 ( .A(y[495]), .B(x[495]), .Z(n23959) );
  XOR U28710 ( .A(n23962), .B(n23961), .Z(n23960) );
  XOR U28711 ( .A(y[497]), .B(x[497]), .Z(n23961) );
  XOR U28712 ( .A(y[496]), .B(x[496]), .Z(n23962) );
  XOR U28713 ( .A(n23954), .B(n23953), .Z(n23963) );
  XOR U28714 ( .A(n23956), .B(n23955), .Z(n23953) );
  XOR U28715 ( .A(y[494]), .B(x[494]), .Z(n23955) );
  XOR U28716 ( .A(y[493]), .B(x[493]), .Z(n23956) );
  XOR U28717 ( .A(y[492]), .B(x[492]), .Z(n23954) );
  XNOR U28718 ( .A(n23947), .B(n23946), .Z(n23949) );
  XNOR U28719 ( .A(n23943), .B(n23942), .Z(n23946) );
  XOR U28720 ( .A(n23945), .B(n23944), .Z(n23942) );
  XOR U28721 ( .A(y[491]), .B(x[491]), .Z(n23944) );
  XOR U28722 ( .A(y[490]), .B(x[490]), .Z(n23945) );
  XOR U28723 ( .A(y[489]), .B(x[489]), .Z(n23943) );
  XOR U28724 ( .A(n23937), .B(n23936), .Z(n23947) );
  XOR U28725 ( .A(n23939), .B(n23938), .Z(n23936) );
  XOR U28726 ( .A(y[488]), .B(x[488]), .Z(n23938) );
  XOR U28727 ( .A(y[487]), .B(x[487]), .Z(n23939) );
  XOR U28728 ( .A(y[486]), .B(x[486]), .Z(n23937) );
  NAND U28729 ( .A(n24000), .B(n24001), .Z(N28173) );
  NAND U28730 ( .A(n24002), .B(n24003), .Z(n24001) );
  NANDN U28731 ( .A(n24004), .B(n24005), .Z(n24003) );
  NANDN U28732 ( .A(n24005), .B(n24004), .Z(n24000) );
  XOR U28733 ( .A(n24004), .B(n24006), .Z(N28172) );
  XNOR U28734 ( .A(n24002), .B(n24005), .Z(n24006) );
  NAND U28735 ( .A(n24007), .B(n24008), .Z(n24005) );
  NAND U28736 ( .A(n24009), .B(n24010), .Z(n24008) );
  NANDN U28737 ( .A(n24011), .B(n24012), .Z(n24010) );
  NANDN U28738 ( .A(n24012), .B(n24011), .Z(n24007) );
  AND U28739 ( .A(n24013), .B(n24014), .Z(n24002) );
  NAND U28740 ( .A(n24015), .B(n24016), .Z(n24014) );
  OR U28741 ( .A(n24017), .B(n24018), .Z(n24016) );
  NAND U28742 ( .A(n24018), .B(n24017), .Z(n24013) );
  IV U28743 ( .A(n24019), .Z(n24018) );
  AND U28744 ( .A(n24020), .B(n24021), .Z(n24004) );
  NAND U28745 ( .A(n24022), .B(n24023), .Z(n24021) );
  NANDN U28746 ( .A(n24024), .B(n24025), .Z(n24023) );
  NANDN U28747 ( .A(n24025), .B(n24024), .Z(n24020) );
  XOR U28748 ( .A(n24017), .B(n24026), .Z(N28171) );
  XOR U28749 ( .A(n24015), .B(n24019), .Z(n24026) );
  XNOR U28750 ( .A(n24012), .B(n24027), .Z(n24019) );
  XNOR U28751 ( .A(n24009), .B(n24011), .Z(n24027) );
  AND U28752 ( .A(n24028), .B(n24029), .Z(n24011) );
  NANDN U28753 ( .A(n24030), .B(n24031), .Z(n24029) );
  NANDN U28754 ( .A(n24032), .B(n24033), .Z(n24031) );
  IV U28755 ( .A(n24034), .Z(n24033) );
  NAND U28756 ( .A(n24034), .B(n24032), .Z(n24028) );
  AND U28757 ( .A(n24035), .B(n24036), .Z(n24009) );
  NAND U28758 ( .A(n24037), .B(n24038), .Z(n24036) );
  OR U28759 ( .A(n24039), .B(n24040), .Z(n24038) );
  NAND U28760 ( .A(n24040), .B(n24039), .Z(n24035) );
  IV U28761 ( .A(n24041), .Z(n24040) );
  NAND U28762 ( .A(n24042), .B(n24043), .Z(n24012) );
  NANDN U28763 ( .A(n24044), .B(n24045), .Z(n24043) );
  NAND U28764 ( .A(n24046), .B(n24047), .Z(n24045) );
  OR U28765 ( .A(n24047), .B(n24046), .Z(n24042) );
  IV U28766 ( .A(n24048), .Z(n24046) );
  AND U28767 ( .A(n24049), .B(n24050), .Z(n24015) );
  NAND U28768 ( .A(n24051), .B(n24052), .Z(n24050) );
  NANDN U28769 ( .A(n24053), .B(n24054), .Z(n24052) );
  NANDN U28770 ( .A(n24054), .B(n24053), .Z(n24049) );
  XOR U28771 ( .A(n24025), .B(n24055), .Z(n24017) );
  XNOR U28772 ( .A(n24022), .B(n24024), .Z(n24055) );
  AND U28773 ( .A(n24056), .B(n24057), .Z(n24024) );
  NANDN U28774 ( .A(n24058), .B(n24059), .Z(n24057) );
  NANDN U28775 ( .A(n24060), .B(n24061), .Z(n24059) );
  IV U28776 ( .A(n24062), .Z(n24061) );
  NAND U28777 ( .A(n24062), .B(n24060), .Z(n24056) );
  AND U28778 ( .A(n24063), .B(n24064), .Z(n24022) );
  NAND U28779 ( .A(n24065), .B(n24066), .Z(n24064) );
  OR U28780 ( .A(n24067), .B(n24068), .Z(n24066) );
  NAND U28781 ( .A(n24068), .B(n24067), .Z(n24063) );
  IV U28782 ( .A(n24069), .Z(n24068) );
  NAND U28783 ( .A(n24070), .B(n24071), .Z(n24025) );
  NANDN U28784 ( .A(n24072), .B(n24073), .Z(n24071) );
  NAND U28785 ( .A(n24074), .B(n24075), .Z(n24073) );
  OR U28786 ( .A(n24075), .B(n24074), .Z(n24070) );
  IV U28787 ( .A(n24076), .Z(n24074) );
  XOR U28788 ( .A(n24051), .B(n24077), .Z(N28170) );
  XNOR U28789 ( .A(n24054), .B(n24053), .Z(n24077) );
  XNOR U28790 ( .A(n24065), .B(n24078), .Z(n24053) );
  XOR U28791 ( .A(n24069), .B(n24067), .Z(n24078) );
  XOR U28792 ( .A(n24075), .B(n24079), .Z(n24067) );
  XOR U28793 ( .A(n24072), .B(n24076), .Z(n24079) );
  NAND U28794 ( .A(n24080), .B(n24081), .Z(n24076) );
  NAND U28795 ( .A(n24082), .B(n24083), .Z(n24081) );
  NAND U28796 ( .A(n24084), .B(n24085), .Z(n24080) );
  AND U28797 ( .A(n24086), .B(n24087), .Z(n24072) );
  NAND U28798 ( .A(n24088), .B(n24089), .Z(n24087) );
  NAND U28799 ( .A(n24090), .B(n24091), .Z(n24086) );
  NANDN U28800 ( .A(n24092), .B(n24093), .Z(n24075) );
  NANDN U28801 ( .A(n24094), .B(n24095), .Z(n24069) );
  XNOR U28802 ( .A(n24060), .B(n24096), .Z(n24065) );
  XOR U28803 ( .A(n24058), .B(n24062), .Z(n24096) );
  NAND U28804 ( .A(n24097), .B(n24098), .Z(n24062) );
  NAND U28805 ( .A(n24099), .B(n24100), .Z(n24098) );
  NAND U28806 ( .A(n24101), .B(n24102), .Z(n24097) );
  AND U28807 ( .A(n24103), .B(n24104), .Z(n24058) );
  NAND U28808 ( .A(n24105), .B(n24106), .Z(n24104) );
  NAND U28809 ( .A(n24107), .B(n24108), .Z(n24103) );
  AND U28810 ( .A(n24109), .B(n24110), .Z(n24060) );
  NAND U28811 ( .A(n24111), .B(n24112), .Z(n24054) );
  XNOR U28812 ( .A(n24037), .B(n24113), .Z(n24051) );
  XOR U28813 ( .A(n24041), .B(n24039), .Z(n24113) );
  XOR U28814 ( .A(n24047), .B(n24114), .Z(n24039) );
  XOR U28815 ( .A(n24044), .B(n24048), .Z(n24114) );
  NAND U28816 ( .A(n24115), .B(n24116), .Z(n24048) );
  NAND U28817 ( .A(n24117), .B(n24118), .Z(n24116) );
  NAND U28818 ( .A(n24119), .B(n24120), .Z(n24115) );
  AND U28819 ( .A(n24121), .B(n24122), .Z(n24044) );
  NAND U28820 ( .A(n24123), .B(n24124), .Z(n24122) );
  NAND U28821 ( .A(n24125), .B(n24126), .Z(n24121) );
  NANDN U28822 ( .A(n24127), .B(n24128), .Z(n24047) );
  NANDN U28823 ( .A(n24129), .B(n24130), .Z(n24041) );
  XNOR U28824 ( .A(n24032), .B(n24131), .Z(n24037) );
  XOR U28825 ( .A(n24030), .B(n24034), .Z(n24131) );
  NAND U28826 ( .A(n24132), .B(n24133), .Z(n24034) );
  NAND U28827 ( .A(n24134), .B(n24135), .Z(n24133) );
  NAND U28828 ( .A(n24136), .B(n24137), .Z(n24132) );
  AND U28829 ( .A(n24138), .B(n24139), .Z(n24030) );
  NAND U28830 ( .A(n24140), .B(n24141), .Z(n24139) );
  NAND U28831 ( .A(n24142), .B(n24143), .Z(n24138) );
  AND U28832 ( .A(n24144), .B(n24145), .Z(n24032) );
  XOR U28833 ( .A(n24112), .B(n24111), .Z(N28169) );
  XNOR U28834 ( .A(n24130), .B(n24129), .Z(n24111) );
  XNOR U28835 ( .A(n24144), .B(n24145), .Z(n24129) );
  XOR U28836 ( .A(n24141), .B(n24140), .Z(n24145) );
  XOR U28837 ( .A(y[483]), .B(x[483]), .Z(n24140) );
  XOR U28838 ( .A(n24143), .B(n24142), .Z(n24141) );
  XOR U28839 ( .A(y[485]), .B(x[485]), .Z(n24142) );
  XOR U28840 ( .A(y[484]), .B(x[484]), .Z(n24143) );
  XOR U28841 ( .A(n24135), .B(n24134), .Z(n24144) );
  XOR U28842 ( .A(n24137), .B(n24136), .Z(n24134) );
  XOR U28843 ( .A(y[482]), .B(x[482]), .Z(n24136) );
  XOR U28844 ( .A(y[481]), .B(x[481]), .Z(n24137) );
  XOR U28845 ( .A(y[480]), .B(x[480]), .Z(n24135) );
  XNOR U28846 ( .A(n24128), .B(n24127), .Z(n24130) );
  XNOR U28847 ( .A(n24124), .B(n24123), .Z(n24127) );
  XOR U28848 ( .A(n24126), .B(n24125), .Z(n24123) );
  XOR U28849 ( .A(y[479]), .B(x[479]), .Z(n24125) );
  XOR U28850 ( .A(y[478]), .B(x[478]), .Z(n24126) );
  XOR U28851 ( .A(y[477]), .B(x[477]), .Z(n24124) );
  XOR U28852 ( .A(n24118), .B(n24117), .Z(n24128) );
  XOR U28853 ( .A(n24120), .B(n24119), .Z(n24117) );
  XOR U28854 ( .A(y[476]), .B(x[476]), .Z(n24119) );
  XOR U28855 ( .A(y[475]), .B(x[475]), .Z(n24120) );
  XOR U28856 ( .A(y[474]), .B(x[474]), .Z(n24118) );
  XNOR U28857 ( .A(n24095), .B(n24094), .Z(n24112) );
  XNOR U28858 ( .A(n24109), .B(n24110), .Z(n24094) );
  XOR U28859 ( .A(n24106), .B(n24105), .Z(n24110) );
  XOR U28860 ( .A(y[471]), .B(x[471]), .Z(n24105) );
  XOR U28861 ( .A(n24108), .B(n24107), .Z(n24106) );
  XOR U28862 ( .A(y[473]), .B(x[473]), .Z(n24107) );
  XOR U28863 ( .A(y[472]), .B(x[472]), .Z(n24108) );
  XOR U28864 ( .A(n24100), .B(n24099), .Z(n24109) );
  XOR U28865 ( .A(n24102), .B(n24101), .Z(n24099) );
  XOR U28866 ( .A(y[470]), .B(x[470]), .Z(n24101) );
  XOR U28867 ( .A(y[469]), .B(x[469]), .Z(n24102) );
  XOR U28868 ( .A(y[468]), .B(x[468]), .Z(n24100) );
  XNOR U28869 ( .A(n24093), .B(n24092), .Z(n24095) );
  XNOR U28870 ( .A(n24089), .B(n24088), .Z(n24092) );
  XOR U28871 ( .A(n24091), .B(n24090), .Z(n24088) );
  XOR U28872 ( .A(y[467]), .B(x[467]), .Z(n24090) );
  XOR U28873 ( .A(y[466]), .B(x[466]), .Z(n24091) );
  XOR U28874 ( .A(y[465]), .B(x[465]), .Z(n24089) );
  XOR U28875 ( .A(n24083), .B(n24082), .Z(n24093) );
  XOR U28876 ( .A(n24085), .B(n24084), .Z(n24082) );
  XOR U28877 ( .A(y[464]), .B(x[464]), .Z(n24084) );
  XOR U28878 ( .A(y[463]), .B(x[463]), .Z(n24085) );
  XOR U28879 ( .A(y[462]), .B(x[462]), .Z(n24083) );
  NAND U28880 ( .A(n24146), .B(n24147), .Z(N28161) );
  NAND U28881 ( .A(n24148), .B(n24149), .Z(n24147) );
  NANDN U28882 ( .A(n24150), .B(n24151), .Z(n24149) );
  NANDN U28883 ( .A(n24151), .B(n24150), .Z(n24146) );
  XOR U28884 ( .A(n24150), .B(n24152), .Z(N28160) );
  XNOR U28885 ( .A(n24148), .B(n24151), .Z(n24152) );
  NAND U28886 ( .A(n24153), .B(n24154), .Z(n24151) );
  NAND U28887 ( .A(n24155), .B(n24156), .Z(n24154) );
  NANDN U28888 ( .A(n24157), .B(n24158), .Z(n24156) );
  NANDN U28889 ( .A(n24158), .B(n24157), .Z(n24153) );
  AND U28890 ( .A(n24159), .B(n24160), .Z(n24148) );
  NAND U28891 ( .A(n24161), .B(n24162), .Z(n24160) );
  OR U28892 ( .A(n24163), .B(n24164), .Z(n24162) );
  NAND U28893 ( .A(n24164), .B(n24163), .Z(n24159) );
  IV U28894 ( .A(n24165), .Z(n24164) );
  AND U28895 ( .A(n24166), .B(n24167), .Z(n24150) );
  NAND U28896 ( .A(n24168), .B(n24169), .Z(n24167) );
  NANDN U28897 ( .A(n24170), .B(n24171), .Z(n24169) );
  NANDN U28898 ( .A(n24171), .B(n24170), .Z(n24166) );
  XOR U28899 ( .A(n24163), .B(n24172), .Z(N28159) );
  XOR U28900 ( .A(n24161), .B(n24165), .Z(n24172) );
  XNOR U28901 ( .A(n24158), .B(n24173), .Z(n24165) );
  XNOR U28902 ( .A(n24155), .B(n24157), .Z(n24173) );
  AND U28903 ( .A(n24174), .B(n24175), .Z(n24157) );
  NANDN U28904 ( .A(n24176), .B(n24177), .Z(n24175) );
  NANDN U28905 ( .A(n24178), .B(n24179), .Z(n24177) );
  IV U28906 ( .A(n24180), .Z(n24179) );
  NAND U28907 ( .A(n24180), .B(n24178), .Z(n24174) );
  AND U28908 ( .A(n24181), .B(n24182), .Z(n24155) );
  NAND U28909 ( .A(n24183), .B(n24184), .Z(n24182) );
  OR U28910 ( .A(n24185), .B(n24186), .Z(n24184) );
  NAND U28911 ( .A(n24186), .B(n24185), .Z(n24181) );
  IV U28912 ( .A(n24187), .Z(n24186) );
  NAND U28913 ( .A(n24188), .B(n24189), .Z(n24158) );
  NANDN U28914 ( .A(n24190), .B(n24191), .Z(n24189) );
  NAND U28915 ( .A(n24192), .B(n24193), .Z(n24191) );
  OR U28916 ( .A(n24193), .B(n24192), .Z(n24188) );
  IV U28917 ( .A(n24194), .Z(n24192) );
  AND U28918 ( .A(n24195), .B(n24196), .Z(n24161) );
  NAND U28919 ( .A(n24197), .B(n24198), .Z(n24196) );
  NANDN U28920 ( .A(n24199), .B(n24200), .Z(n24198) );
  NANDN U28921 ( .A(n24200), .B(n24199), .Z(n24195) );
  XOR U28922 ( .A(n24171), .B(n24201), .Z(n24163) );
  XNOR U28923 ( .A(n24168), .B(n24170), .Z(n24201) );
  AND U28924 ( .A(n24202), .B(n24203), .Z(n24170) );
  NANDN U28925 ( .A(n24204), .B(n24205), .Z(n24203) );
  NANDN U28926 ( .A(n24206), .B(n24207), .Z(n24205) );
  IV U28927 ( .A(n24208), .Z(n24207) );
  NAND U28928 ( .A(n24208), .B(n24206), .Z(n24202) );
  AND U28929 ( .A(n24209), .B(n24210), .Z(n24168) );
  NAND U28930 ( .A(n24211), .B(n24212), .Z(n24210) );
  OR U28931 ( .A(n24213), .B(n24214), .Z(n24212) );
  NAND U28932 ( .A(n24214), .B(n24213), .Z(n24209) );
  IV U28933 ( .A(n24215), .Z(n24214) );
  NAND U28934 ( .A(n24216), .B(n24217), .Z(n24171) );
  NANDN U28935 ( .A(n24218), .B(n24219), .Z(n24217) );
  NAND U28936 ( .A(n24220), .B(n24221), .Z(n24219) );
  OR U28937 ( .A(n24221), .B(n24220), .Z(n24216) );
  IV U28938 ( .A(n24222), .Z(n24220) );
  XOR U28939 ( .A(n24197), .B(n24223), .Z(N28158) );
  XNOR U28940 ( .A(n24200), .B(n24199), .Z(n24223) );
  XNOR U28941 ( .A(n24211), .B(n24224), .Z(n24199) );
  XOR U28942 ( .A(n24215), .B(n24213), .Z(n24224) );
  XOR U28943 ( .A(n24221), .B(n24225), .Z(n24213) );
  XOR U28944 ( .A(n24218), .B(n24222), .Z(n24225) );
  NAND U28945 ( .A(n24226), .B(n24227), .Z(n24222) );
  NAND U28946 ( .A(n24228), .B(n24229), .Z(n24227) );
  NAND U28947 ( .A(n24230), .B(n24231), .Z(n24226) );
  AND U28948 ( .A(n24232), .B(n24233), .Z(n24218) );
  NAND U28949 ( .A(n24234), .B(n24235), .Z(n24233) );
  NAND U28950 ( .A(n24236), .B(n24237), .Z(n24232) );
  NANDN U28951 ( .A(n24238), .B(n24239), .Z(n24221) );
  NANDN U28952 ( .A(n24240), .B(n24241), .Z(n24215) );
  XNOR U28953 ( .A(n24206), .B(n24242), .Z(n24211) );
  XOR U28954 ( .A(n24204), .B(n24208), .Z(n24242) );
  NAND U28955 ( .A(n24243), .B(n24244), .Z(n24208) );
  NAND U28956 ( .A(n24245), .B(n24246), .Z(n24244) );
  NAND U28957 ( .A(n24247), .B(n24248), .Z(n24243) );
  AND U28958 ( .A(n24249), .B(n24250), .Z(n24204) );
  NAND U28959 ( .A(n24251), .B(n24252), .Z(n24250) );
  NAND U28960 ( .A(n24253), .B(n24254), .Z(n24249) );
  AND U28961 ( .A(n24255), .B(n24256), .Z(n24206) );
  NAND U28962 ( .A(n24257), .B(n24258), .Z(n24200) );
  XNOR U28963 ( .A(n24183), .B(n24259), .Z(n24197) );
  XOR U28964 ( .A(n24187), .B(n24185), .Z(n24259) );
  XOR U28965 ( .A(n24193), .B(n24260), .Z(n24185) );
  XOR U28966 ( .A(n24190), .B(n24194), .Z(n24260) );
  NAND U28967 ( .A(n24261), .B(n24262), .Z(n24194) );
  NAND U28968 ( .A(n24263), .B(n24264), .Z(n24262) );
  NAND U28969 ( .A(n24265), .B(n24266), .Z(n24261) );
  AND U28970 ( .A(n24267), .B(n24268), .Z(n24190) );
  NAND U28971 ( .A(n24269), .B(n24270), .Z(n24268) );
  NAND U28972 ( .A(n24271), .B(n24272), .Z(n24267) );
  NANDN U28973 ( .A(n24273), .B(n24274), .Z(n24193) );
  NANDN U28974 ( .A(n24275), .B(n24276), .Z(n24187) );
  XNOR U28975 ( .A(n24178), .B(n24277), .Z(n24183) );
  XOR U28976 ( .A(n24176), .B(n24180), .Z(n24277) );
  NAND U28977 ( .A(n24278), .B(n24279), .Z(n24180) );
  NAND U28978 ( .A(n24280), .B(n24281), .Z(n24279) );
  NAND U28979 ( .A(n24282), .B(n24283), .Z(n24278) );
  AND U28980 ( .A(n24284), .B(n24285), .Z(n24176) );
  NAND U28981 ( .A(n24286), .B(n24287), .Z(n24285) );
  NAND U28982 ( .A(n24288), .B(n24289), .Z(n24284) );
  AND U28983 ( .A(n24290), .B(n24291), .Z(n24178) );
  XOR U28984 ( .A(n24258), .B(n24257), .Z(N28157) );
  XNOR U28985 ( .A(n24276), .B(n24275), .Z(n24257) );
  XNOR U28986 ( .A(n24290), .B(n24291), .Z(n24275) );
  XOR U28987 ( .A(n24287), .B(n24286), .Z(n24291) );
  XOR U28988 ( .A(y[459]), .B(x[459]), .Z(n24286) );
  XOR U28989 ( .A(n24289), .B(n24288), .Z(n24287) );
  XOR U28990 ( .A(y[461]), .B(x[461]), .Z(n24288) );
  XOR U28991 ( .A(y[460]), .B(x[460]), .Z(n24289) );
  XOR U28992 ( .A(n24281), .B(n24280), .Z(n24290) );
  XOR U28993 ( .A(n24283), .B(n24282), .Z(n24280) );
  XOR U28994 ( .A(y[458]), .B(x[458]), .Z(n24282) );
  XOR U28995 ( .A(y[457]), .B(x[457]), .Z(n24283) );
  XOR U28996 ( .A(y[456]), .B(x[456]), .Z(n24281) );
  XNOR U28997 ( .A(n24274), .B(n24273), .Z(n24276) );
  XNOR U28998 ( .A(n24270), .B(n24269), .Z(n24273) );
  XOR U28999 ( .A(n24272), .B(n24271), .Z(n24269) );
  XOR U29000 ( .A(y[455]), .B(x[455]), .Z(n24271) );
  XOR U29001 ( .A(y[454]), .B(x[454]), .Z(n24272) );
  XOR U29002 ( .A(y[453]), .B(x[453]), .Z(n24270) );
  XOR U29003 ( .A(n24264), .B(n24263), .Z(n24274) );
  XOR U29004 ( .A(n24266), .B(n24265), .Z(n24263) );
  XOR U29005 ( .A(y[452]), .B(x[452]), .Z(n24265) );
  XOR U29006 ( .A(y[451]), .B(x[451]), .Z(n24266) );
  XOR U29007 ( .A(y[450]), .B(x[450]), .Z(n24264) );
  XNOR U29008 ( .A(n24241), .B(n24240), .Z(n24258) );
  XNOR U29009 ( .A(n24255), .B(n24256), .Z(n24240) );
  XOR U29010 ( .A(n24252), .B(n24251), .Z(n24256) );
  XOR U29011 ( .A(y[447]), .B(x[447]), .Z(n24251) );
  XOR U29012 ( .A(n24254), .B(n24253), .Z(n24252) );
  XOR U29013 ( .A(y[449]), .B(x[449]), .Z(n24253) );
  XOR U29014 ( .A(y[448]), .B(x[448]), .Z(n24254) );
  XOR U29015 ( .A(n24246), .B(n24245), .Z(n24255) );
  XOR U29016 ( .A(n24248), .B(n24247), .Z(n24245) );
  XOR U29017 ( .A(y[446]), .B(x[446]), .Z(n24247) );
  XOR U29018 ( .A(y[445]), .B(x[445]), .Z(n24248) );
  XOR U29019 ( .A(y[444]), .B(x[444]), .Z(n24246) );
  XNOR U29020 ( .A(n24239), .B(n24238), .Z(n24241) );
  XNOR U29021 ( .A(n24235), .B(n24234), .Z(n24238) );
  XOR U29022 ( .A(n24237), .B(n24236), .Z(n24234) );
  XOR U29023 ( .A(y[443]), .B(x[443]), .Z(n24236) );
  XOR U29024 ( .A(y[442]), .B(x[442]), .Z(n24237) );
  XOR U29025 ( .A(y[441]), .B(x[441]), .Z(n24235) );
  XOR U29026 ( .A(n24229), .B(n24228), .Z(n24239) );
  XOR U29027 ( .A(n24231), .B(n24230), .Z(n24228) );
  XOR U29028 ( .A(y[440]), .B(x[440]), .Z(n24230) );
  XOR U29029 ( .A(y[439]), .B(x[439]), .Z(n24231) );
  XOR U29030 ( .A(y[438]), .B(x[438]), .Z(n24229) );
  NAND U29031 ( .A(n24292), .B(n24293), .Z(N28149) );
  NAND U29032 ( .A(n24294), .B(n24295), .Z(n24293) );
  NANDN U29033 ( .A(n24296), .B(n24297), .Z(n24295) );
  NANDN U29034 ( .A(n24297), .B(n24296), .Z(n24292) );
  XOR U29035 ( .A(n24296), .B(n24298), .Z(N28148) );
  XNOR U29036 ( .A(n24294), .B(n24297), .Z(n24298) );
  NAND U29037 ( .A(n24299), .B(n24300), .Z(n24297) );
  NAND U29038 ( .A(n24301), .B(n24302), .Z(n24300) );
  NANDN U29039 ( .A(n24303), .B(n24304), .Z(n24302) );
  NANDN U29040 ( .A(n24304), .B(n24303), .Z(n24299) );
  AND U29041 ( .A(n24305), .B(n24306), .Z(n24294) );
  NAND U29042 ( .A(n24307), .B(n24308), .Z(n24306) );
  OR U29043 ( .A(n24309), .B(n24310), .Z(n24308) );
  NAND U29044 ( .A(n24310), .B(n24309), .Z(n24305) );
  IV U29045 ( .A(n24311), .Z(n24310) );
  AND U29046 ( .A(n24312), .B(n24313), .Z(n24296) );
  NAND U29047 ( .A(n24314), .B(n24315), .Z(n24313) );
  NANDN U29048 ( .A(n24316), .B(n24317), .Z(n24315) );
  NANDN U29049 ( .A(n24317), .B(n24316), .Z(n24312) );
  XOR U29050 ( .A(n24309), .B(n24318), .Z(N28147) );
  XOR U29051 ( .A(n24307), .B(n24311), .Z(n24318) );
  XNOR U29052 ( .A(n24304), .B(n24319), .Z(n24311) );
  XNOR U29053 ( .A(n24301), .B(n24303), .Z(n24319) );
  AND U29054 ( .A(n24320), .B(n24321), .Z(n24303) );
  NANDN U29055 ( .A(n24322), .B(n24323), .Z(n24321) );
  NANDN U29056 ( .A(n24324), .B(n24325), .Z(n24323) );
  IV U29057 ( .A(n24326), .Z(n24325) );
  NAND U29058 ( .A(n24326), .B(n24324), .Z(n24320) );
  AND U29059 ( .A(n24327), .B(n24328), .Z(n24301) );
  NAND U29060 ( .A(n24329), .B(n24330), .Z(n24328) );
  OR U29061 ( .A(n24331), .B(n24332), .Z(n24330) );
  NAND U29062 ( .A(n24332), .B(n24331), .Z(n24327) );
  IV U29063 ( .A(n24333), .Z(n24332) );
  NAND U29064 ( .A(n24334), .B(n24335), .Z(n24304) );
  NANDN U29065 ( .A(n24336), .B(n24337), .Z(n24335) );
  NAND U29066 ( .A(n24338), .B(n24339), .Z(n24337) );
  OR U29067 ( .A(n24339), .B(n24338), .Z(n24334) );
  IV U29068 ( .A(n24340), .Z(n24338) );
  AND U29069 ( .A(n24341), .B(n24342), .Z(n24307) );
  NAND U29070 ( .A(n24343), .B(n24344), .Z(n24342) );
  NANDN U29071 ( .A(n24345), .B(n24346), .Z(n24344) );
  NANDN U29072 ( .A(n24346), .B(n24345), .Z(n24341) );
  XOR U29073 ( .A(n24317), .B(n24347), .Z(n24309) );
  XNOR U29074 ( .A(n24314), .B(n24316), .Z(n24347) );
  AND U29075 ( .A(n24348), .B(n24349), .Z(n24316) );
  NANDN U29076 ( .A(n24350), .B(n24351), .Z(n24349) );
  NANDN U29077 ( .A(n24352), .B(n24353), .Z(n24351) );
  IV U29078 ( .A(n24354), .Z(n24353) );
  NAND U29079 ( .A(n24354), .B(n24352), .Z(n24348) );
  AND U29080 ( .A(n24355), .B(n24356), .Z(n24314) );
  NAND U29081 ( .A(n24357), .B(n24358), .Z(n24356) );
  OR U29082 ( .A(n24359), .B(n24360), .Z(n24358) );
  NAND U29083 ( .A(n24360), .B(n24359), .Z(n24355) );
  IV U29084 ( .A(n24361), .Z(n24360) );
  NAND U29085 ( .A(n24362), .B(n24363), .Z(n24317) );
  NANDN U29086 ( .A(n24364), .B(n24365), .Z(n24363) );
  NAND U29087 ( .A(n24366), .B(n24367), .Z(n24365) );
  OR U29088 ( .A(n24367), .B(n24366), .Z(n24362) );
  IV U29089 ( .A(n24368), .Z(n24366) );
  XOR U29090 ( .A(n24343), .B(n24369), .Z(N28146) );
  XNOR U29091 ( .A(n24346), .B(n24345), .Z(n24369) );
  XNOR U29092 ( .A(n24357), .B(n24370), .Z(n24345) );
  XOR U29093 ( .A(n24361), .B(n24359), .Z(n24370) );
  XOR U29094 ( .A(n24367), .B(n24371), .Z(n24359) );
  XOR U29095 ( .A(n24364), .B(n24368), .Z(n24371) );
  NAND U29096 ( .A(n24372), .B(n24373), .Z(n24368) );
  NAND U29097 ( .A(n24374), .B(n24375), .Z(n24373) );
  NAND U29098 ( .A(n24376), .B(n24377), .Z(n24372) );
  AND U29099 ( .A(n24378), .B(n24379), .Z(n24364) );
  NAND U29100 ( .A(n24380), .B(n24381), .Z(n24379) );
  NAND U29101 ( .A(n24382), .B(n24383), .Z(n24378) );
  NANDN U29102 ( .A(n24384), .B(n24385), .Z(n24367) );
  NANDN U29103 ( .A(n24386), .B(n24387), .Z(n24361) );
  XNOR U29104 ( .A(n24352), .B(n24388), .Z(n24357) );
  XOR U29105 ( .A(n24350), .B(n24354), .Z(n24388) );
  NAND U29106 ( .A(n24389), .B(n24390), .Z(n24354) );
  NAND U29107 ( .A(n24391), .B(n24392), .Z(n24390) );
  NAND U29108 ( .A(n24393), .B(n24394), .Z(n24389) );
  AND U29109 ( .A(n24395), .B(n24396), .Z(n24350) );
  NAND U29110 ( .A(n24397), .B(n24398), .Z(n24396) );
  NAND U29111 ( .A(n24399), .B(n24400), .Z(n24395) );
  AND U29112 ( .A(n24401), .B(n24402), .Z(n24352) );
  NAND U29113 ( .A(n24403), .B(n24404), .Z(n24346) );
  XNOR U29114 ( .A(n24329), .B(n24405), .Z(n24343) );
  XOR U29115 ( .A(n24333), .B(n24331), .Z(n24405) );
  XOR U29116 ( .A(n24339), .B(n24406), .Z(n24331) );
  XOR U29117 ( .A(n24336), .B(n24340), .Z(n24406) );
  NAND U29118 ( .A(n24407), .B(n24408), .Z(n24340) );
  NAND U29119 ( .A(n24409), .B(n24410), .Z(n24408) );
  NAND U29120 ( .A(n24411), .B(n24412), .Z(n24407) );
  AND U29121 ( .A(n24413), .B(n24414), .Z(n24336) );
  NAND U29122 ( .A(n24415), .B(n24416), .Z(n24414) );
  NAND U29123 ( .A(n24417), .B(n24418), .Z(n24413) );
  NANDN U29124 ( .A(n24419), .B(n24420), .Z(n24339) );
  NANDN U29125 ( .A(n24421), .B(n24422), .Z(n24333) );
  XNOR U29126 ( .A(n24324), .B(n24423), .Z(n24329) );
  XOR U29127 ( .A(n24322), .B(n24326), .Z(n24423) );
  NAND U29128 ( .A(n24424), .B(n24425), .Z(n24326) );
  NAND U29129 ( .A(n24426), .B(n24427), .Z(n24425) );
  NAND U29130 ( .A(n24428), .B(n24429), .Z(n24424) );
  AND U29131 ( .A(n24430), .B(n24431), .Z(n24322) );
  NAND U29132 ( .A(n24432), .B(n24433), .Z(n24431) );
  NAND U29133 ( .A(n24434), .B(n24435), .Z(n24430) );
  AND U29134 ( .A(n24436), .B(n24437), .Z(n24324) );
  XOR U29135 ( .A(n24404), .B(n24403), .Z(N28145) );
  XNOR U29136 ( .A(n24422), .B(n24421), .Z(n24403) );
  XNOR U29137 ( .A(n24436), .B(n24437), .Z(n24421) );
  XOR U29138 ( .A(n24433), .B(n24432), .Z(n24437) );
  XOR U29139 ( .A(y[435]), .B(x[435]), .Z(n24432) );
  XOR U29140 ( .A(n24435), .B(n24434), .Z(n24433) );
  XOR U29141 ( .A(y[437]), .B(x[437]), .Z(n24434) );
  XOR U29142 ( .A(y[436]), .B(x[436]), .Z(n24435) );
  XOR U29143 ( .A(n24427), .B(n24426), .Z(n24436) );
  XOR U29144 ( .A(n24429), .B(n24428), .Z(n24426) );
  XOR U29145 ( .A(y[434]), .B(x[434]), .Z(n24428) );
  XOR U29146 ( .A(y[433]), .B(x[433]), .Z(n24429) );
  XOR U29147 ( .A(y[432]), .B(x[432]), .Z(n24427) );
  XNOR U29148 ( .A(n24420), .B(n24419), .Z(n24422) );
  XNOR U29149 ( .A(n24416), .B(n24415), .Z(n24419) );
  XOR U29150 ( .A(n24418), .B(n24417), .Z(n24415) );
  XOR U29151 ( .A(y[431]), .B(x[431]), .Z(n24417) );
  XOR U29152 ( .A(y[430]), .B(x[430]), .Z(n24418) );
  XOR U29153 ( .A(y[429]), .B(x[429]), .Z(n24416) );
  XOR U29154 ( .A(n24410), .B(n24409), .Z(n24420) );
  XOR U29155 ( .A(n24412), .B(n24411), .Z(n24409) );
  XOR U29156 ( .A(y[428]), .B(x[428]), .Z(n24411) );
  XOR U29157 ( .A(y[427]), .B(x[427]), .Z(n24412) );
  XOR U29158 ( .A(y[426]), .B(x[426]), .Z(n24410) );
  XNOR U29159 ( .A(n24387), .B(n24386), .Z(n24404) );
  XNOR U29160 ( .A(n24401), .B(n24402), .Z(n24386) );
  XOR U29161 ( .A(n24398), .B(n24397), .Z(n24402) );
  XOR U29162 ( .A(y[423]), .B(x[423]), .Z(n24397) );
  XOR U29163 ( .A(n24400), .B(n24399), .Z(n24398) );
  XOR U29164 ( .A(y[425]), .B(x[425]), .Z(n24399) );
  XOR U29165 ( .A(y[424]), .B(x[424]), .Z(n24400) );
  XOR U29166 ( .A(n24392), .B(n24391), .Z(n24401) );
  XOR U29167 ( .A(n24394), .B(n24393), .Z(n24391) );
  XOR U29168 ( .A(y[422]), .B(x[422]), .Z(n24393) );
  XOR U29169 ( .A(y[421]), .B(x[421]), .Z(n24394) );
  XOR U29170 ( .A(y[420]), .B(x[420]), .Z(n24392) );
  XNOR U29171 ( .A(n24385), .B(n24384), .Z(n24387) );
  XNOR U29172 ( .A(n24381), .B(n24380), .Z(n24384) );
  XOR U29173 ( .A(n24383), .B(n24382), .Z(n24380) );
  XOR U29174 ( .A(y[419]), .B(x[419]), .Z(n24382) );
  XOR U29175 ( .A(y[418]), .B(x[418]), .Z(n24383) );
  XOR U29176 ( .A(y[417]), .B(x[417]), .Z(n24381) );
  XOR U29177 ( .A(n24375), .B(n24374), .Z(n24385) );
  XOR U29178 ( .A(n24377), .B(n24376), .Z(n24374) );
  XOR U29179 ( .A(y[416]), .B(x[416]), .Z(n24376) );
  XOR U29180 ( .A(y[415]), .B(x[415]), .Z(n24377) );
  XOR U29181 ( .A(y[414]), .B(x[414]), .Z(n24375) );
  NAND U29182 ( .A(n24438), .B(n24439), .Z(N28137) );
  NAND U29183 ( .A(n24440), .B(n24441), .Z(n24439) );
  NANDN U29184 ( .A(n24442), .B(n24443), .Z(n24441) );
  NANDN U29185 ( .A(n24443), .B(n24442), .Z(n24438) );
  XOR U29186 ( .A(n24442), .B(n24444), .Z(N28136) );
  XNOR U29187 ( .A(n24440), .B(n24443), .Z(n24444) );
  NAND U29188 ( .A(n24445), .B(n24446), .Z(n24443) );
  NAND U29189 ( .A(n24447), .B(n24448), .Z(n24446) );
  NANDN U29190 ( .A(n24449), .B(n24450), .Z(n24448) );
  NANDN U29191 ( .A(n24450), .B(n24449), .Z(n24445) );
  AND U29192 ( .A(n24451), .B(n24452), .Z(n24440) );
  NAND U29193 ( .A(n24453), .B(n24454), .Z(n24452) );
  OR U29194 ( .A(n24455), .B(n24456), .Z(n24454) );
  NAND U29195 ( .A(n24456), .B(n24455), .Z(n24451) );
  IV U29196 ( .A(n24457), .Z(n24456) );
  AND U29197 ( .A(n24458), .B(n24459), .Z(n24442) );
  NAND U29198 ( .A(n24460), .B(n24461), .Z(n24459) );
  NANDN U29199 ( .A(n24462), .B(n24463), .Z(n24461) );
  NANDN U29200 ( .A(n24463), .B(n24462), .Z(n24458) );
  XOR U29201 ( .A(n24455), .B(n24464), .Z(N28135) );
  XOR U29202 ( .A(n24453), .B(n24457), .Z(n24464) );
  XNOR U29203 ( .A(n24450), .B(n24465), .Z(n24457) );
  XNOR U29204 ( .A(n24447), .B(n24449), .Z(n24465) );
  AND U29205 ( .A(n24466), .B(n24467), .Z(n24449) );
  NANDN U29206 ( .A(n24468), .B(n24469), .Z(n24467) );
  NANDN U29207 ( .A(n24470), .B(n24471), .Z(n24469) );
  IV U29208 ( .A(n24472), .Z(n24471) );
  NAND U29209 ( .A(n24472), .B(n24470), .Z(n24466) );
  AND U29210 ( .A(n24473), .B(n24474), .Z(n24447) );
  NAND U29211 ( .A(n24475), .B(n24476), .Z(n24474) );
  OR U29212 ( .A(n24477), .B(n24478), .Z(n24476) );
  NAND U29213 ( .A(n24478), .B(n24477), .Z(n24473) );
  IV U29214 ( .A(n24479), .Z(n24478) );
  NAND U29215 ( .A(n24480), .B(n24481), .Z(n24450) );
  NANDN U29216 ( .A(n24482), .B(n24483), .Z(n24481) );
  NAND U29217 ( .A(n24484), .B(n24485), .Z(n24483) );
  OR U29218 ( .A(n24485), .B(n24484), .Z(n24480) );
  IV U29219 ( .A(n24486), .Z(n24484) );
  AND U29220 ( .A(n24487), .B(n24488), .Z(n24453) );
  NAND U29221 ( .A(n24489), .B(n24490), .Z(n24488) );
  NANDN U29222 ( .A(n24491), .B(n24492), .Z(n24490) );
  NANDN U29223 ( .A(n24492), .B(n24491), .Z(n24487) );
  XOR U29224 ( .A(n24463), .B(n24493), .Z(n24455) );
  XNOR U29225 ( .A(n24460), .B(n24462), .Z(n24493) );
  AND U29226 ( .A(n24494), .B(n24495), .Z(n24462) );
  NANDN U29227 ( .A(n24496), .B(n24497), .Z(n24495) );
  NANDN U29228 ( .A(n24498), .B(n24499), .Z(n24497) );
  IV U29229 ( .A(n24500), .Z(n24499) );
  NAND U29230 ( .A(n24500), .B(n24498), .Z(n24494) );
  AND U29231 ( .A(n24501), .B(n24502), .Z(n24460) );
  NAND U29232 ( .A(n24503), .B(n24504), .Z(n24502) );
  OR U29233 ( .A(n24505), .B(n24506), .Z(n24504) );
  NAND U29234 ( .A(n24506), .B(n24505), .Z(n24501) );
  IV U29235 ( .A(n24507), .Z(n24506) );
  NAND U29236 ( .A(n24508), .B(n24509), .Z(n24463) );
  NANDN U29237 ( .A(n24510), .B(n24511), .Z(n24509) );
  NAND U29238 ( .A(n24512), .B(n24513), .Z(n24511) );
  OR U29239 ( .A(n24513), .B(n24512), .Z(n24508) );
  IV U29240 ( .A(n24514), .Z(n24512) );
  XOR U29241 ( .A(n24489), .B(n24515), .Z(N28134) );
  XNOR U29242 ( .A(n24492), .B(n24491), .Z(n24515) );
  XNOR U29243 ( .A(n24503), .B(n24516), .Z(n24491) );
  XOR U29244 ( .A(n24507), .B(n24505), .Z(n24516) );
  XOR U29245 ( .A(n24513), .B(n24517), .Z(n24505) );
  XOR U29246 ( .A(n24510), .B(n24514), .Z(n24517) );
  NAND U29247 ( .A(n24518), .B(n24519), .Z(n24514) );
  NAND U29248 ( .A(n24520), .B(n24521), .Z(n24519) );
  NAND U29249 ( .A(n24522), .B(n24523), .Z(n24518) );
  AND U29250 ( .A(n24524), .B(n24525), .Z(n24510) );
  NAND U29251 ( .A(n24526), .B(n24527), .Z(n24525) );
  NAND U29252 ( .A(n24528), .B(n24529), .Z(n24524) );
  NANDN U29253 ( .A(n24530), .B(n24531), .Z(n24513) );
  NANDN U29254 ( .A(n24532), .B(n24533), .Z(n24507) );
  XNOR U29255 ( .A(n24498), .B(n24534), .Z(n24503) );
  XOR U29256 ( .A(n24496), .B(n24500), .Z(n24534) );
  NAND U29257 ( .A(n24535), .B(n24536), .Z(n24500) );
  NAND U29258 ( .A(n24537), .B(n24538), .Z(n24536) );
  NAND U29259 ( .A(n24539), .B(n24540), .Z(n24535) );
  AND U29260 ( .A(n24541), .B(n24542), .Z(n24496) );
  NAND U29261 ( .A(n24543), .B(n24544), .Z(n24542) );
  NAND U29262 ( .A(n24545), .B(n24546), .Z(n24541) );
  AND U29263 ( .A(n24547), .B(n24548), .Z(n24498) );
  NAND U29264 ( .A(n24549), .B(n24550), .Z(n24492) );
  XNOR U29265 ( .A(n24475), .B(n24551), .Z(n24489) );
  XOR U29266 ( .A(n24479), .B(n24477), .Z(n24551) );
  XOR U29267 ( .A(n24485), .B(n24552), .Z(n24477) );
  XOR U29268 ( .A(n24482), .B(n24486), .Z(n24552) );
  NAND U29269 ( .A(n24553), .B(n24554), .Z(n24486) );
  NAND U29270 ( .A(n24555), .B(n24556), .Z(n24554) );
  NAND U29271 ( .A(n24557), .B(n24558), .Z(n24553) );
  AND U29272 ( .A(n24559), .B(n24560), .Z(n24482) );
  NAND U29273 ( .A(n24561), .B(n24562), .Z(n24560) );
  NAND U29274 ( .A(n24563), .B(n24564), .Z(n24559) );
  NANDN U29275 ( .A(n24565), .B(n24566), .Z(n24485) );
  NANDN U29276 ( .A(n24567), .B(n24568), .Z(n24479) );
  XNOR U29277 ( .A(n24470), .B(n24569), .Z(n24475) );
  XOR U29278 ( .A(n24468), .B(n24472), .Z(n24569) );
  NAND U29279 ( .A(n24570), .B(n24571), .Z(n24472) );
  NAND U29280 ( .A(n24572), .B(n24573), .Z(n24571) );
  NAND U29281 ( .A(n24574), .B(n24575), .Z(n24570) );
  AND U29282 ( .A(n24576), .B(n24577), .Z(n24468) );
  NAND U29283 ( .A(n24578), .B(n24579), .Z(n24577) );
  NAND U29284 ( .A(n24580), .B(n24581), .Z(n24576) );
  AND U29285 ( .A(n24582), .B(n24583), .Z(n24470) );
  XOR U29286 ( .A(n24550), .B(n24549), .Z(N28133) );
  XNOR U29287 ( .A(n24568), .B(n24567), .Z(n24549) );
  XNOR U29288 ( .A(n24582), .B(n24583), .Z(n24567) );
  XOR U29289 ( .A(n24579), .B(n24578), .Z(n24583) );
  XOR U29290 ( .A(y[411]), .B(x[411]), .Z(n24578) );
  XOR U29291 ( .A(n24581), .B(n24580), .Z(n24579) );
  XOR U29292 ( .A(y[413]), .B(x[413]), .Z(n24580) );
  XOR U29293 ( .A(y[412]), .B(x[412]), .Z(n24581) );
  XOR U29294 ( .A(n24573), .B(n24572), .Z(n24582) );
  XOR U29295 ( .A(n24575), .B(n24574), .Z(n24572) );
  XOR U29296 ( .A(y[410]), .B(x[410]), .Z(n24574) );
  XOR U29297 ( .A(y[409]), .B(x[409]), .Z(n24575) );
  XOR U29298 ( .A(y[408]), .B(x[408]), .Z(n24573) );
  XNOR U29299 ( .A(n24566), .B(n24565), .Z(n24568) );
  XNOR U29300 ( .A(n24562), .B(n24561), .Z(n24565) );
  XOR U29301 ( .A(n24564), .B(n24563), .Z(n24561) );
  XOR U29302 ( .A(y[407]), .B(x[407]), .Z(n24563) );
  XOR U29303 ( .A(y[406]), .B(x[406]), .Z(n24564) );
  XOR U29304 ( .A(y[405]), .B(x[405]), .Z(n24562) );
  XOR U29305 ( .A(n24556), .B(n24555), .Z(n24566) );
  XOR U29306 ( .A(n24558), .B(n24557), .Z(n24555) );
  XOR U29307 ( .A(y[404]), .B(x[404]), .Z(n24557) );
  XOR U29308 ( .A(y[403]), .B(x[403]), .Z(n24558) );
  XOR U29309 ( .A(y[402]), .B(x[402]), .Z(n24556) );
  XNOR U29310 ( .A(n24533), .B(n24532), .Z(n24550) );
  XNOR U29311 ( .A(n24547), .B(n24548), .Z(n24532) );
  XOR U29312 ( .A(n24544), .B(n24543), .Z(n24548) );
  XOR U29313 ( .A(y[399]), .B(x[399]), .Z(n24543) );
  XOR U29314 ( .A(n24546), .B(n24545), .Z(n24544) );
  XOR U29315 ( .A(y[401]), .B(x[401]), .Z(n24545) );
  XOR U29316 ( .A(y[400]), .B(x[400]), .Z(n24546) );
  XOR U29317 ( .A(n24538), .B(n24537), .Z(n24547) );
  XOR U29318 ( .A(n24540), .B(n24539), .Z(n24537) );
  XOR U29319 ( .A(y[398]), .B(x[398]), .Z(n24539) );
  XOR U29320 ( .A(y[397]), .B(x[397]), .Z(n24540) );
  XOR U29321 ( .A(y[396]), .B(x[396]), .Z(n24538) );
  XNOR U29322 ( .A(n24531), .B(n24530), .Z(n24533) );
  XNOR U29323 ( .A(n24527), .B(n24526), .Z(n24530) );
  XOR U29324 ( .A(n24529), .B(n24528), .Z(n24526) );
  XOR U29325 ( .A(y[395]), .B(x[395]), .Z(n24528) );
  XOR U29326 ( .A(y[394]), .B(x[394]), .Z(n24529) );
  XOR U29327 ( .A(y[393]), .B(x[393]), .Z(n24527) );
  XOR U29328 ( .A(n24521), .B(n24520), .Z(n24531) );
  XOR U29329 ( .A(n24523), .B(n24522), .Z(n24520) );
  XOR U29330 ( .A(y[392]), .B(x[392]), .Z(n24522) );
  XOR U29331 ( .A(y[391]), .B(x[391]), .Z(n24523) );
  XOR U29332 ( .A(y[390]), .B(x[390]), .Z(n24521) );
  NAND U29333 ( .A(n24584), .B(n24585), .Z(N28125) );
  NAND U29334 ( .A(n24586), .B(n24587), .Z(n24585) );
  NANDN U29335 ( .A(n24588), .B(n24589), .Z(n24587) );
  NANDN U29336 ( .A(n24589), .B(n24588), .Z(n24584) );
  XOR U29337 ( .A(n24588), .B(n24590), .Z(N28124) );
  XNOR U29338 ( .A(n24586), .B(n24589), .Z(n24590) );
  NAND U29339 ( .A(n24591), .B(n24592), .Z(n24589) );
  NAND U29340 ( .A(n24593), .B(n24594), .Z(n24592) );
  NANDN U29341 ( .A(n24595), .B(n24596), .Z(n24594) );
  NANDN U29342 ( .A(n24596), .B(n24595), .Z(n24591) );
  AND U29343 ( .A(n24597), .B(n24598), .Z(n24586) );
  NAND U29344 ( .A(n24599), .B(n24600), .Z(n24598) );
  OR U29345 ( .A(n24601), .B(n24602), .Z(n24600) );
  NAND U29346 ( .A(n24602), .B(n24601), .Z(n24597) );
  IV U29347 ( .A(n24603), .Z(n24602) );
  AND U29348 ( .A(n24604), .B(n24605), .Z(n24588) );
  NAND U29349 ( .A(n24606), .B(n24607), .Z(n24605) );
  NANDN U29350 ( .A(n24608), .B(n24609), .Z(n24607) );
  NANDN U29351 ( .A(n24609), .B(n24608), .Z(n24604) );
  XOR U29352 ( .A(n24601), .B(n24610), .Z(N28123) );
  XOR U29353 ( .A(n24599), .B(n24603), .Z(n24610) );
  XNOR U29354 ( .A(n24596), .B(n24611), .Z(n24603) );
  XNOR U29355 ( .A(n24593), .B(n24595), .Z(n24611) );
  AND U29356 ( .A(n24612), .B(n24613), .Z(n24595) );
  NANDN U29357 ( .A(n24614), .B(n24615), .Z(n24613) );
  NANDN U29358 ( .A(n24616), .B(n24617), .Z(n24615) );
  IV U29359 ( .A(n24618), .Z(n24617) );
  NAND U29360 ( .A(n24618), .B(n24616), .Z(n24612) );
  AND U29361 ( .A(n24619), .B(n24620), .Z(n24593) );
  NAND U29362 ( .A(n24621), .B(n24622), .Z(n24620) );
  OR U29363 ( .A(n24623), .B(n24624), .Z(n24622) );
  NAND U29364 ( .A(n24624), .B(n24623), .Z(n24619) );
  IV U29365 ( .A(n24625), .Z(n24624) );
  NAND U29366 ( .A(n24626), .B(n24627), .Z(n24596) );
  NANDN U29367 ( .A(n24628), .B(n24629), .Z(n24627) );
  NAND U29368 ( .A(n24630), .B(n24631), .Z(n24629) );
  OR U29369 ( .A(n24631), .B(n24630), .Z(n24626) );
  IV U29370 ( .A(n24632), .Z(n24630) );
  AND U29371 ( .A(n24633), .B(n24634), .Z(n24599) );
  NAND U29372 ( .A(n24635), .B(n24636), .Z(n24634) );
  NANDN U29373 ( .A(n24637), .B(n24638), .Z(n24636) );
  NANDN U29374 ( .A(n24638), .B(n24637), .Z(n24633) );
  XOR U29375 ( .A(n24609), .B(n24639), .Z(n24601) );
  XNOR U29376 ( .A(n24606), .B(n24608), .Z(n24639) );
  AND U29377 ( .A(n24640), .B(n24641), .Z(n24608) );
  NANDN U29378 ( .A(n24642), .B(n24643), .Z(n24641) );
  NANDN U29379 ( .A(n24644), .B(n24645), .Z(n24643) );
  IV U29380 ( .A(n24646), .Z(n24645) );
  NAND U29381 ( .A(n24646), .B(n24644), .Z(n24640) );
  AND U29382 ( .A(n24647), .B(n24648), .Z(n24606) );
  NAND U29383 ( .A(n24649), .B(n24650), .Z(n24648) );
  OR U29384 ( .A(n24651), .B(n24652), .Z(n24650) );
  NAND U29385 ( .A(n24652), .B(n24651), .Z(n24647) );
  IV U29386 ( .A(n24653), .Z(n24652) );
  NAND U29387 ( .A(n24654), .B(n24655), .Z(n24609) );
  NANDN U29388 ( .A(n24656), .B(n24657), .Z(n24655) );
  NAND U29389 ( .A(n24658), .B(n24659), .Z(n24657) );
  OR U29390 ( .A(n24659), .B(n24658), .Z(n24654) );
  IV U29391 ( .A(n24660), .Z(n24658) );
  XOR U29392 ( .A(n24635), .B(n24661), .Z(N28122) );
  XNOR U29393 ( .A(n24638), .B(n24637), .Z(n24661) );
  XNOR U29394 ( .A(n24649), .B(n24662), .Z(n24637) );
  XOR U29395 ( .A(n24653), .B(n24651), .Z(n24662) );
  XOR U29396 ( .A(n24659), .B(n24663), .Z(n24651) );
  XOR U29397 ( .A(n24656), .B(n24660), .Z(n24663) );
  NAND U29398 ( .A(n24664), .B(n24665), .Z(n24660) );
  NAND U29399 ( .A(n24666), .B(n24667), .Z(n24665) );
  NAND U29400 ( .A(n24668), .B(n24669), .Z(n24664) );
  AND U29401 ( .A(n24670), .B(n24671), .Z(n24656) );
  NAND U29402 ( .A(n24672), .B(n24673), .Z(n24671) );
  NAND U29403 ( .A(n24674), .B(n24675), .Z(n24670) );
  NANDN U29404 ( .A(n24676), .B(n24677), .Z(n24659) );
  NANDN U29405 ( .A(n24678), .B(n24679), .Z(n24653) );
  XNOR U29406 ( .A(n24644), .B(n24680), .Z(n24649) );
  XOR U29407 ( .A(n24642), .B(n24646), .Z(n24680) );
  NAND U29408 ( .A(n24681), .B(n24682), .Z(n24646) );
  NAND U29409 ( .A(n24683), .B(n24684), .Z(n24682) );
  NAND U29410 ( .A(n24685), .B(n24686), .Z(n24681) );
  AND U29411 ( .A(n24687), .B(n24688), .Z(n24642) );
  NAND U29412 ( .A(n24689), .B(n24690), .Z(n24688) );
  NAND U29413 ( .A(n24691), .B(n24692), .Z(n24687) );
  AND U29414 ( .A(n24693), .B(n24694), .Z(n24644) );
  NAND U29415 ( .A(n24695), .B(n24696), .Z(n24638) );
  XNOR U29416 ( .A(n24621), .B(n24697), .Z(n24635) );
  XOR U29417 ( .A(n24625), .B(n24623), .Z(n24697) );
  XOR U29418 ( .A(n24631), .B(n24698), .Z(n24623) );
  XOR U29419 ( .A(n24628), .B(n24632), .Z(n24698) );
  NAND U29420 ( .A(n24699), .B(n24700), .Z(n24632) );
  NAND U29421 ( .A(n24701), .B(n24702), .Z(n24700) );
  NAND U29422 ( .A(n24703), .B(n24704), .Z(n24699) );
  AND U29423 ( .A(n24705), .B(n24706), .Z(n24628) );
  NAND U29424 ( .A(n24707), .B(n24708), .Z(n24706) );
  NAND U29425 ( .A(n24709), .B(n24710), .Z(n24705) );
  NANDN U29426 ( .A(n24711), .B(n24712), .Z(n24631) );
  NANDN U29427 ( .A(n24713), .B(n24714), .Z(n24625) );
  XNOR U29428 ( .A(n24616), .B(n24715), .Z(n24621) );
  XOR U29429 ( .A(n24614), .B(n24618), .Z(n24715) );
  NAND U29430 ( .A(n24716), .B(n24717), .Z(n24618) );
  NAND U29431 ( .A(n24718), .B(n24719), .Z(n24717) );
  NAND U29432 ( .A(n24720), .B(n24721), .Z(n24716) );
  AND U29433 ( .A(n24722), .B(n24723), .Z(n24614) );
  NAND U29434 ( .A(n24724), .B(n24725), .Z(n24723) );
  NAND U29435 ( .A(n24726), .B(n24727), .Z(n24722) );
  AND U29436 ( .A(n24728), .B(n24729), .Z(n24616) );
  XOR U29437 ( .A(n24696), .B(n24695), .Z(N28121) );
  XNOR U29438 ( .A(n24714), .B(n24713), .Z(n24695) );
  XNOR U29439 ( .A(n24728), .B(n24729), .Z(n24713) );
  XOR U29440 ( .A(n24725), .B(n24724), .Z(n24729) );
  XOR U29441 ( .A(y[387]), .B(x[387]), .Z(n24724) );
  XOR U29442 ( .A(n24727), .B(n24726), .Z(n24725) );
  XOR U29443 ( .A(y[389]), .B(x[389]), .Z(n24726) );
  XOR U29444 ( .A(y[388]), .B(x[388]), .Z(n24727) );
  XOR U29445 ( .A(n24719), .B(n24718), .Z(n24728) );
  XOR U29446 ( .A(n24721), .B(n24720), .Z(n24718) );
  XOR U29447 ( .A(y[386]), .B(x[386]), .Z(n24720) );
  XOR U29448 ( .A(y[385]), .B(x[385]), .Z(n24721) );
  XOR U29449 ( .A(y[384]), .B(x[384]), .Z(n24719) );
  XNOR U29450 ( .A(n24712), .B(n24711), .Z(n24714) );
  XNOR U29451 ( .A(n24708), .B(n24707), .Z(n24711) );
  XOR U29452 ( .A(n24710), .B(n24709), .Z(n24707) );
  XOR U29453 ( .A(y[383]), .B(x[383]), .Z(n24709) );
  XOR U29454 ( .A(y[382]), .B(x[382]), .Z(n24710) );
  XOR U29455 ( .A(y[381]), .B(x[381]), .Z(n24708) );
  XOR U29456 ( .A(n24702), .B(n24701), .Z(n24712) );
  XOR U29457 ( .A(n24704), .B(n24703), .Z(n24701) );
  XOR U29458 ( .A(y[380]), .B(x[380]), .Z(n24703) );
  XOR U29459 ( .A(y[379]), .B(x[379]), .Z(n24704) );
  XOR U29460 ( .A(y[378]), .B(x[378]), .Z(n24702) );
  XNOR U29461 ( .A(n24679), .B(n24678), .Z(n24696) );
  XNOR U29462 ( .A(n24693), .B(n24694), .Z(n24678) );
  XOR U29463 ( .A(n24690), .B(n24689), .Z(n24694) );
  XOR U29464 ( .A(y[375]), .B(x[375]), .Z(n24689) );
  XOR U29465 ( .A(n24692), .B(n24691), .Z(n24690) );
  XOR U29466 ( .A(y[377]), .B(x[377]), .Z(n24691) );
  XOR U29467 ( .A(y[376]), .B(x[376]), .Z(n24692) );
  XOR U29468 ( .A(n24684), .B(n24683), .Z(n24693) );
  XOR U29469 ( .A(n24686), .B(n24685), .Z(n24683) );
  XOR U29470 ( .A(y[374]), .B(x[374]), .Z(n24685) );
  XOR U29471 ( .A(y[373]), .B(x[373]), .Z(n24686) );
  XOR U29472 ( .A(y[372]), .B(x[372]), .Z(n24684) );
  XNOR U29473 ( .A(n24677), .B(n24676), .Z(n24679) );
  XNOR U29474 ( .A(n24673), .B(n24672), .Z(n24676) );
  XOR U29475 ( .A(n24675), .B(n24674), .Z(n24672) );
  XOR U29476 ( .A(y[371]), .B(x[371]), .Z(n24674) );
  XOR U29477 ( .A(y[370]), .B(x[370]), .Z(n24675) );
  XOR U29478 ( .A(y[369]), .B(x[369]), .Z(n24673) );
  XOR U29479 ( .A(n24667), .B(n24666), .Z(n24677) );
  XOR U29480 ( .A(n24669), .B(n24668), .Z(n24666) );
  XOR U29481 ( .A(y[368]), .B(x[368]), .Z(n24668) );
  XOR U29482 ( .A(y[367]), .B(x[367]), .Z(n24669) );
  XOR U29483 ( .A(y[366]), .B(x[366]), .Z(n24667) );
  NAND U29484 ( .A(n24730), .B(n24731), .Z(N28113) );
  NAND U29485 ( .A(n24732), .B(n24733), .Z(n24731) );
  NANDN U29486 ( .A(n24734), .B(n24735), .Z(n24733) );
  NANDN U29487 ( .A(n24735), .B(n24734), .Z(n24730) );
  XOR U29488 ( .A(n24734), .B(n24736), .Z(N28112) );
  XNOR U29489 ( .A(n24732), .B(n24735), .Z(n24736) );
  NAND U29490 ( .A(n24737), .B(n24738), .Z(n24735) );
  NAND U29491 ( .A(n24739), .B(n24740), .Z(n24738) );
  NANDN U29492 ( .A(n24741), .B(n24742), .Z(n24740) );
  NANDN U29493 ( .A(n24742), .B(n24741), .Z(n24737) );
  AND U29494 ( .A(n24743), .B(n24744), .Z(n24732) );
  NAND U29495 ( .A(n24745), .B(n24746), .Z(n24744) );
  OR U29496 ( .A(n24747), .B(n24748), .Z(n24746) );
  NAND U29497 ( .A(n24748), .B(n24747), .Z(n24743) );
  IV U29498 ( .A(n24749), .Z(n24748) );
  AND U29499 ( .A(n24750), .B(n24751), .Z(n24734) );
  NAND U29500 ( .A(n24752), .B(n24753), .Z(n24751) );
  NANDN U29501 ( .A(n24754), .B(n24755), .Z(n24753) );
  NANDN U29502 ( .A(n24755), .B(n24754), .Z(n24750) );
  XOR U29503 ( .A(n24747), .B(n24756), .Z(N28111) );
  XOR U29504 ( .A(n24745), .B(n24749), .Z(n24756) );
  XNOR U29505 ( .A(n24742), .B(n24757), .Z(n24749) );
  XNOR U29506 ( .A(n24739), .B(n24741), .Z(n24757) );
  AND U29507 ( .A(n24758), .B(n24759), .Z(n24741) );
  NANDN U29508 ( .A(n24760), .B(n24761), .Z(n24759) );
  NANDN U29509 ( .A(n24762), .B(n24763), .Z(n24761) );
  IV U29510 ( .A(n24764), .Z(n24763) );
  NAND U29511 ( .A(n24764), .B(n24762), .Z(n24758) );
  AND U29512 ( .A(n24765), .B(n24766), .Z(n24739) );
  NAND U29513 ( .A(n24767), .B(n24768), .Z(n24766) );
  OR U29514 ( .A(n24769), .B(n24770), .Z(n24768) );
  NAND U29515 ( .A(n24770), .B(n24769), .Z(n24765) );
  IV U29516 ( .A(n24771), .Z(n24770) );
  NAND U29517 ( .A(n24772), .B(n24773), .Z(n24742) );
  NANDN U29518 ( .A(n24774), .B(n24775), .Z(n24773) );
  NAND U29519 ( .A(n24776), .B(n24777), .Z(n24775) );
  OR U29520 ( .A(n24777), .B(n24776), .Z(n24772) );
  IV U29521 ( .A(n24778), .Z(n24776) );
  AND U29522 ( .A(n24779), .B(n24780), .Z(n24745) );
  NAND U29523 ( .A(n24781), .B(n24782), .Z(n24780) );
  NANDN U29524 ( .A(n24783), .B(n24784), .Z(n24782) );
  NANDN U29525 ( .A(n24784), .B(n24783), .Z(n24779) );
  XOR U29526 ( .A(n24755), .B(n24785), .Z(n24747) );
  XNOR U29527 ( .A(n24752), .B(n24754), .Z(n24785) );
  AND U29528 ( .A(n24786), .B(n24787), .Z(n24754) );
  NANDN U29529 ( .A(n24788), .B(n24789), .Z(n24787) );
  NANDN U29530 ( .A(n24790), .B(n24791), .Z(n24789) );
  IV U29531 ( .A(n24792), .Z(n24791) );
  NAND U29532 ( .A(n24792), .B(n24790), .Z(n24786) );
  AND U29533 ( .A(n24793), .B(n24794), .Z(n24752) );
  NAND U29534 ( .A(n24795), .B(n24796), .Z(n24794) );
  OR U29535 ( .A(n24797), .B(n24798), .Z(n24796) );
  NAND U29536 ( .A(n24798), .B(n24797), .Z(n24793) );
  IV U29537 ( .A(n24799), .Z(n24798) );
  NAND U29538 ( .A(n24800), .B(n24801), .Z(n24755) );
  NANDN U29539 ( .A(n24802), .B(n24803), .Z(n24801) );
  NAND U29540 ( .A(n24804), .B(n24805), .Z(n24803) );
  OR U29541 ( .A(n24805), .B(n24804), .Z(n24800) );
  IV U29542 ( .A(n24806), .Z(n24804) );
  XOR U29543 ( .A(n24781), .B(n24807), .Z(N28110) );
  XNOR U29544 ( .A(n24784), .B(n24783), .Z(n24807) );
  XNOR U29545 ( .A(n24795), .B(n24808), .Z(n24783) );
  XOR U29546 ( .A(n24799), .B(n24797), .Z(n24808) );
  XOR U29547 ( .A(n24805), .B(n24809), .Z(n24797) );
  XOR U29548 ( .A(n24802), .B(n24806), .Z(n24809) );
  NAND U29549 ( .A(n24810), .B(n24811), .Z(n24806) );
  NAND U29550 ( .A(n24812), .B(n24813), .Z(n24811) );
  NAND U29551 ( .A(n24814), .B(n24815), .Z(n24810) );
  AND U29552 ( .A(n24816), .B(n24817), .Z(n24802) );
  NAND U29553 ( .A(n24818), .B(n24819), .Z(n24817) );
  NAND U29554 ( .A(n24820), .B(n24821), .Z(n24816) );
  NANDN U29555 ( .A(n24822), .B(n24823), .Z(n24805) );
  NANDN U29556 ( .A(n24824), .B(n24825), .Z(n24799) );
  XNOR U29557 ( .A(n24790), .B(n24826), .Z(n24795) );
  XOR U29558 ( .A(n24788), .B(n24792), .Z(n24826) );
  NAND U29559 ( .A(n24827), .B(n24828), .Z(n24792) );
  NAND U29560 ( .A(n24829), .B(n24830), .Z(n24828) );
  NAND U29561 ( .A(n24831), .B(n24832), .Z(n24827) );
  AND U29562 ( .A(n24833), .B(n24834), .Z(n24788) );
  NAND U29563 ( .A(n24835), .B(n24836), .Z(n24834) );
  NAND U29564 ( .A(n24837), .B(n24838), .Z(n24833) );
  AND U29565 ( .A(n24839), .B(n24840), .Z(n24790) );
  NAND U29566 ( .A(n24841), .B(n24842), .Z(n24784) );
  XNOR U29567 ( .A(n24767), .B(n24843), .Z(n24781) );
  XOR U29568 ( .A(n24771), .B(n24769), .Z(n24843) );
  XOR U29569 ( .A(n24777), .B(n24844), .Z(n24769) );
  XOR U29570 ( .A(n24774), .B(n24778), .Z(n24844) );
  NAND U29571 ( .A(n24845), .B(n24846), .Z(n24778) );
  NAND U29572 ( .A(n24847), .B(n24848), .Z(n24846) );
  NAND U29573 ( .A(n24849), .B(n24850), .Z(n24845) );
  AND U29574 ( .A(n24851), .B(n24852), .Z(n24774) );
  NAND U29575 ( .A(n24853), .B(n24854), .Z(n24852) );
  NAND U29576 ( .A(n24855), .B(n24856), .Z(n24851) );
  NANDN U29577 ( .A(n24857), .B(n24858), .Z(n24777) );
  NANDN U29578 ( .A(n24859), .B(n24860), .Z(n24771) );
  XNOR U29579 ( .A(n24762), .B(n24861), .Z(n24767) );
  XOR U29580 ( .A(n24760), .B(n24764), .Z(n24861) );
  NAND U29581 ( .A(n24862), .B(n24863), .Z(n24764) );
  NAND U29582 ( .A(n24864), .B(n24865), .Z(n24863) );
  NAND U29583 ( .A(n24866), .B(n24867), .Z(n24862) );
  AND U29584 ( .A(n24868), .B(n24869), .Z(n24760) );
  NAND U29585 ( .A(n24870), .B(n24871), .Z(n24869) );
  NAND U29586 ( .A(n24872), .B(n24873), .Z(n24868) );
  AND U29587 ( .A(n24874), .B(n24875), .Z(n24762) );
  XOR U29588 ( .A(n24842), .B(n24841), .Z(N28109) );
  XNOR U29589 ( .A(n24860), .B(n24859), .Z(n24841) );
  XNOR U29590 ( .A(n24874), .B(n24875), .Z(n24859) );
  XOR U29591 ( .A(n24871), .B(n24870), .Z(n24875) );
  XOR U29592 ( .A(y[363]), .B(x[363]), .Z(n24870) );
  XOR U29593 ( .A(n24873), .B(n24872), .Z(n24871) );
  XOR U29594 ( .A(y[365]), .B(x[365]), .Z(n24872) );
  XOR U29595 ( .A(y[364]), .B(x[364]), .Z(n24873) );
  XOR U29596 ( .A(n24865), .B(n24864), .Z(n24874) );
  XOR U29597 ( .A(n24867), .B(n24866), .Z(n24864) );
  XOR U29598 ( .A(y[362]), .B(x[362]), .Z(n24866) );
  XOR U29599 ( .A(y[361]), .B(x[361]), .Z(n24867) );
  XOR U29600 ( .A(y[360]), .B(x[360]), .Z(n24865) );
  XNOR U29601 ( .A(n24858), .B(n24857), .Z(n24860) );
  XNOR U29602 ( .A(n24854), .B(n24853), .Z(n24857) );
  XOR U29603 ( .A(n24856), .B(n24855), .Z(n24853) );
  XOR U29604 ( .A(y[359]), .B(x[359]), .Z(n24855) );
  XOR U29605 ( .A(y[358]), .B(x[358]), .Z(n24856) );
  XOR U29606 ( .A(y[357]), .B(x[357]), .Z(n24854) );
  XOR U29607 ( .A(n24848), .B(n24847), .Z(n24858) );
  XOR U29608 ( .A(n24850), .B(n24849), .Z(n24847) );
  XOR U29609 ( .A(y[356]), .B(x[356]), .Z(n24849) );
  XOR U29610 ( .A(y[355]), .B(x[355]), .Z(n24850) );
  XOR U29611 ( .A(y[354]), .B(x[354]), .Z(n24848) );
  XNOR U29612 ( .A(n24825), .B(n24824), .Z(n24842) );
  XNOR U29613 ( .A(n24839), .B(n24840), .Z(n24824) );
  XOR U29614 ( .A(n24836), .B(n24835), .Z(n24840) );
  XOR U29615 ( .A(y[351]), .B(x[351]), .Z(n24835) );
  XOR U29616 ( .A(n24838), .B(n24837), .Z(n24836) );
  XOR U29617 ( .A(y[353]), .B(x[353]), .Z(n24837) );
  XOR U29618 ( .A(y[352]), .B(x[352]), .Z(n24838) );
  XOR U29619 ( .A(n24830), .B(n24829), .Z(n24839) );
  XOR U29620 ( .A(n24832), .B(n24831), .Z(n24829) );
  XOR U29621 ( .A(y[350]), .B(x[350]), .Z(n24831) );
  XOR U29622 ( .A(y[349]), .B(x[349]), .Z(n24832) );
  XOR U29623 ( .A(y[348]), .B(x[348]), .Z(n24830) );
  XNOR U29624 ( .A(n24823), .B(n24822), .Z(n24825) );
  XNOR U29625 ( .A(n24819), .B(n24818), .Z(n24822) );
  XOR U29626 ( .A(n24821), .B(n24820), .Z(n24818) );
  XOR U29627 ( .A(y[347]), .B(x[347]), .Z(n24820) );
  XOR U29628 ( .A(y[346]), .B(x[346]), .Z(n24821) );
  XOR U29629 ( .A(y[345]), .B(x[345]), .Z(n24819) );
  XOR U29630 ( .A(n24813), .B(n24812), .Z(n24823) );
  XOR U29631 ( .A(n24815), .B(n24814), .Z(n24812) );
  XOR U29632 ( .A(y[344]), .B(x[344]), .Z(n24814) );
  XOR U29633 ( .A(y[343]), .B(x[343]), .Z(n24815) );
  XOR U29634 ( .A(y[342]), .B(x[342]), .Z(n24813) );
  NAND U29635 ( .A(n24876), .B(n24877), .Z(N28101) );
  NAND U29636 ( .A(n24878), .B(n24879), .Z(n24877) );
  NANDN U29637 ( .A(n24880), .B(n24881), .Z(n24879) );
  NANDN U29638 ( .A(n24881), .B(n24880), .Z(n24876) );
  XOR U29639 ( .A(n24880), .B(n24882), .Z(N28100) );
  XNOR U29640 ( .A(n24878), .B(n24881), .Z(n24882) );
  NAND U29641 ( .A(n24883), .B(n24884), .Z(n24881) );
  NAND U29642 ( .A(n24885), .B(n24886), .Z(n24884) );
  NANDN U29643 ( .A(n24887), .B(n24888), .Z(n24886) );
  NANDN U29644 ( .A(n24888), .B(n24887), .Z(n24883) );
  AND U29645 ( .A(n24889), .B(n24890), .Z(n24878) );
  NAND U29646 ( .A(n24891), .B(n24892), .Z(n24890) );
  OR U29647 ( .A(n24893), .B(n24894), .Z(n24892) );
  NAND U29648 ( .A(n24894), .B(n24893), .Z(n24889) );
  IV U29649 ( .A(n24895), .Z(n24894) );
  AND U29650 ( .A(n24896), .B(n24897), .Z(n24880) );
  NAND U29651 ( .A(n24898), .B(n24899), .Z(n24897) );
  NANDN U29652 ( .A(n24900), .B(n24901), .Z(n24899) );
  NANDN U29653 ( .A(n24901), .B(n24900), .Z(n24896) );
  XOR U29654 ( .A(n24893), .B(n24902), .Z(N28099) );
  XOR U29655 ( .A(n24891), .B(n24895), .Z(n24902) );
  XNOR U29656 ( .A(n24888), .B(n24903), .Z(n24895) );
  XNOR U29657 ( .A(n24885), .B(n24887), .Z(n24903) );
  AND U29658 ( .A(n24904), .B(n24905), .Z(n24887) );
  NANDN U29659 ( .A(n24906), .B(n24907), .Z(n24905) );
  NANDN U29660 ( .A(n24908), .B(n24909), .Z(n24907) );
  IV U29661 ( .A(n24910), .Z(n24909) );
  NAND U29662 ( .A(n24910), .B(n24908), .Z(n24904) );
  AND U29663 ( .A(n24911), .B(n24912), .Z(n24885) );
  NAND U29664 ( .A(n24913), .B(n24914), .Z(n24912) );
  OR U29665 ( .A(n24915), .B(n24916), .Z(n24914) );
  NAND U29666 ( .A(n24916), .B(n24915), .Z(n24911) );
  IV U29667 ( .A(n24917), .Z(n24916) );
  NAND U29668 ( .A(n24918), .B(n24919), .Z(n24888) );
  NANDN U29669 ( .A(n24920), .B(n24921), .Z(n24919) );
  NAND U29670 ( .A(n24922), .B(n24923), .Z(n24921) );
  OR U29671 ( .A(n24923), .B(n24922), .Z(n24918) );
  IV U29672 ( .A(n24924), .Z(n24922) );
  AND U29673 ( .A(n24925), .B(n24926), .Z(n24891) );
  NAND U29674 ( .A(n24927), .B(n24928), .Z(n24926) );
  NANDN U29675 ( .A(n24929), .B(n24930), .Z(n24928) );
  NANDN U29676 ( .A(n24930), .B(n24929), .Z(n24925) );
  XOR U29677 ( .A(n24901), .B(n24931), .Z(n24893) );
  XNOR U29678 ( .A(n24898), .B(n24900), .Z(n24931) );
  AND U29679 ( .A(n24932), .B(n24933), .Z(n24900) );
  NANDN U29680 ( .A(n24934), .B(n24935), .Z(n24933) );
  NANDN U29681 ( .A(n24936), .B(n24937), .Z(n24935) );
  IV U29682 ( .A(n24938), .Z(n24937) );
  NAND U29683 ( .A(n24938), .B(n24936), .Z(n24932) );
  AND U29684 ( .A(n24939), .B(n24940), .Z(n24898) );
  NAND U29685 ( .A(n24941), .B(n24942), .Z(n24940) );
  OR U29686 ( .A(n24943), .B(n24944), .Z(n24942) );
  NAND U29687 ( .A(n24944), .B(n24943), .Z(n24939) );
  IV U29688 ( .A(n24945), .Z(n24944) );
  NAND U29689 ( .A(n24946), .B(n24947), .Z(n24901) );
  NANDN U29690 ( .A(n24948), .B(n24949), .Z(n24947) );
  NAND U29691 ( .A(n24950), .B(n24951), .Z(n24949) );
  OR U29692 ( .A(n24951), .B(n24950), .Z(n24946) );
  IV U29693 ( .A(n24952), .Z(n24950) );
  XOR U29694 ( .A(n24927), .B(n24953), .Z(N28098) );
  XNOR U29695 ( .A(n24930), .B(n24929), .Z(n24953) );
  XNOR U29696 ( .A(n24941), .B(n24954), .Z(n24929) );
  XOR U29697 ( .A(n24945), .B(n24943), .Z(n24954) );
  XOR U29698 ( .A(n24951), .B(n24955), .Z(n24943) );
  XOR U29699 ( .A(n24948), .B(n24952), .Z(n24955) );
  NAND U29700 ( .A(n24956), .B(n24957), .Z(n24952) );
  NAND U29701 ( .A(n24958), .B(n24959), .Z(n24957) );
  NAND U29702 ( .A(n24960), .B(n24961), .Z(n24956) );
  AND U29703 ( .A(n24962), .B(n24963), .Z(n24948) );
  NAND U29704 ( .A(n24964), .B(n24965), .Z(n24963) );
  NAND U29705 ( .A(n24966), .B(n24967), .Z(n24962) );
  NANDN U29706 ( .A(n24968), .B(n24969), .Z(n24951) );
  NANDN U29707 ( .A(n24970), .B(n24971), .Z(n24945) );
  XNOR U29708 ( .A(n24936), .B(n24972), .Z(n24941) );
  XOR U29709 ( .A(n24934), .B(n24938), .Z(n24972) );
  NAND U29710 ( .A(n24973), .B(n24974), .Z(n24938) );
  NAND U29711 ( .A(n24975), .B(n24976), .Z(n24974) );
  NAND U29712 ( .A(n24977), .B(n24978), .Z(n24973) );
  AND U29713 ( .A(n24979), .B(n24980), .Z(n24934) );
  NAND U29714 ( .A(n24981), .B(n24982), .Z(n24980) );
  NAND U29715 ( .A(n24983), .B(n24984), .Z(n24979) );
  AND U29716 ( .A(n24985), .B(n24986), .Z(n24936) );
  NAND U29717 ( .A(n24987), .B(n24988), .Z(n24930) );
  XNOR U29718 ( .A(n24913), .B(n24989), .Z(n24927) );
  XOR U29719 ( .A(n24917), .B(n24915), .Z(n24989) );
  XOR U29720 ( .A(n24923), .B(n24990), .Z(n24915) );
  XOR U29721 ( .A(n24920), .B(n24924), .Z(n24990) );
  NAND U29722 ( .A(n24991), .B(n24992), .Z(n24924) );
  NAND U29723 ( .A(n24993), .B(n24994), .Z(n24992) );
  NAND U29724 ( .A(n24995), .B(n24996), .Z(n24991) );
  AND U29725 ( .A(n24997), .B(n24998), .Z(n24920) );
  NAND U29726 ( .A(n24999), .B(n25000), .Z(n24998) );
  NAND U29727 ( .A(n25001), .B(n25002), .Z(n24997) );
  NANDN U29728 ( .A(n25003), .B(n25004), .Z(n24923) );
  NANDN U29729 ( .A(n25005), .B(n25006), .Z(n24917) );
  XNOR U29730 ( .A(n24908), .B(n25007), .Z(n24913) );
  XOR U29731 ( .A(n24906), .B(n24910), .Z(n25007) );
  NAND U29732 ( .A(n25008), .B(n25009), .Z(n24910) );
  NAND U29733 ( .A(n25010), .B(n25011), .Z(n25009) );
  NAND U29734 ( .A(n25012), .B(n25013), .Z(n25008) );
  AND U29735 ( .A(n25014), .B(n25015), .Z(n24906) );
  NAND U29736 ( .A(n25016), .B(n25017), .Z(n25015) );
  NAND U29737 ( .A(n25018), .B(n25019), .Z(n25014) );
  AND U29738 ( .A(n25020), .B(n25021), .Z(n24908) );
  XOR U29739 ( .A(n24988), .B(n24987), .Z(N28097) );
  XNOR U29740 ( .A(n25006), .B(n25005), .Z(n24987) );
  XNOR U29741 ( .A(n25020), .B(n25021), .Z(n25005) );
  XOR U29742 ( .A(n25017), .B(n25016), .Z(n25021) );
  XOR U29743 ( .A(y[339]), .B(x[339]), .Z(n25016) );
  XOR U29744 ( .A(n25019), .B(n25018), .Z(n25017) );
  XOR U29745 ( .A(y[341]), .B(x[341]), .Z(n25018) );
  XOR U29746 ( .A(y[340]), .B(x[340]), .Z(n25019) );
  XOR U29747 ( .A(n25011), .B(n25010), .Z(n25020) );
  XOR U29748 ( .A(n25013), .B(n25012), .Z(n25010) );
  XOR U29749 ( .A(y[338]), .B(x[338]), .Z(n25012) );
  XOR U29750 ( .A(y[337]), .B(x[337]), .Z(n25013) );
  XOR U29751 ( .A(y[336]), .B(x[336]), .Z(n25011) );
  XNOR U29752 ( .A(n25004), .B(n25003), .Z(n25006) );
  XNOR U29753 ( .A(n25000), .B(n24999), .Z(n25003) );
  XOR U29754 ( .A(n25002), .B(n25001), .Z(n24999) );
  XOR U29755 ( .A(y[335]), .B(x[335]), .Z(n25001) );
  XOR U29756 ( .A(y[334]), .B(x[334]), .Z(n25002) );
  XOR U29757 ( .A(y[333]), .B(x[333]), .Z(n25000) );
  XOR U29758 ( .A(n24994), .B(n24993), .Z(n25004) );
  XOR U29759 ( .A(n24996), .B(n24995), .Z(n24993) );
  XOR U29760 ( .A(y[332]), .B(x[332]), .Z(n24995) );
  XOR U29761 ( .A(y[331]), .B(x[331]), .Z(n24996) );
  XOR U29762 ( .A(y[330]), .B(x[330]), .Z(n24994) );
  XNOR U29763 ( .A(n24971), .B(n24970), .Z(n24988) );
  XNOR U29764 ( .A(n24985), .B(n24986), .Z(n24970) );
  XOR U29765 ( .A(n24982), .B(n24981), .Z(n24986) );
  XOR U29766 ( .A(y[327]), .B(x[327]), .Z(n24981) );
  XOR U29767 ( .A(n24984), .B(n24983), .Z(n24982) );
  XOR U29768 ( .A(y[329]), .B(x[329]), .Z(n24983) );
  XOR U29769 ( .A(y[328]), .B(x[328]), .Z(n24984) );
  XOR U29770 ( .A(n24976), .B(n24975), .Z(n24985) );
  XOR U29771 ( .A(n24978), .B(n24977), .Z(n24975) );
  XOR U29772 ( .A(y[326]), .B(x[326]), .Z(n24977) );
  XOR U29773 ( .A(y[325]), .B(x[325]), .Z(n24978) );
  XOR U29774 ( .A(y[324]), .B(x[324]), .Z(n24976) );
  XNOR U29775 ( .A(n24969), .B(n24968), .Z(n24971) );
  XNOR U29776 ( .A(n24965), .B(n24964), .Z(n24968) );
  XOR U29777 ( .A(n24967), .B(n24966), .Z(n24964) );
  XOR U29778 ( .A(y[323]), .B(x[323]), .Z(n24966) );
  XOR U29779 ( .A(y[322]), .B(x[322]), .Z(n24967) );
  XOR U29780 ( .A(y[321]), .B(x[321]), .Z(n24965) );
  XOR U29781 ( .A(n24959), .B(n24958), .Z(n24969) );
  XOR U29782 ( .A(n24961), .B(n24960), .Z(n24958) );
  XOR U29783 ( .A(y[320]), .B(x[320]), .Z(n24960) );
  XOR U29784 ( .A(y[319]), .B(x[319]), .Z(n24961) );
  XOR U29785 ( .A(y[318]), .B(x[318]), .Z(n24959) );
  NAND U29786 ( .A(n25022), .B(n25023), .Z(N28089) );
  NAND U29787 ( .A(n25024), .B(n25025), .Z(n25023) );
  NANDN U29788 ( .A(n25026), .B(n25027), .Z(n25025) );
  NANDN U29789 ( .A(n25027), .B(n25026), .Z(n25022) );
  XOR U29790 ( .A(n25026), .B(n25028), .Z(N28088) );
  XNOR U29791 ( .A(n25024), .B(n25027), .Z(n25028) );
  NAND U29792 ( .A(n25029), .B(n25030), .Z(n25027) );
  NAND U29793 ( .A(n25031), .B(n25032), .Z(n25030) );
  NANDN U29794 ( .A(n25033), .B(n25034), .Z(n25032) );
  NANDN U29795 ( .A(n25034), .B(n25033), .Z(n25029) );
  AND U29796 ( .A(n25035), .B(n25036), .Z(n25024) );
  NAND U29797 ( .A(n25037), .B(n25038), .Z(n25036) );
  OR U29798 ( .A(n25039), .B(n25040), .Z(n25038) );
  NAND U29799 ( .A(n25040), .B(n25039), .Z(n25035) );
  IV U29800 ( .A(n25041), .Z(n25040) );
  AND U29801 ( .A(n25042), .B(n25043), .Z(n25026) );
  NAND U29802 ( .A(n25044), .B(n25045), .Z(n25043) );
  NANDN U29803 ( .A(n25046), .B(n25047), .Z(n25045) );
  NANDN U29804 ( .A(n25047), .B(n25046), .Z(n25042) );
  XOR U29805 ( .A(n25039), .B(n25048), .Z(N28087) );
  XOR U29806 ( .A(n25037), .B(n25041), .Z(n25048) );
  XNOR U29807 ( .A(n25034), .B(n25049), .Z(n25041) );
  XNOR U29808 ( .A(n25031), .B(n25033), .Z(n25049) );
  AND U29809 ( .A(n25050), .B(n25051), .Z(n25033) );
  NANDN U29810 ( .A(n25052), .B(n25053), .Z(n25051) );
  NANDN U29811 ( .A(n25054), .B(n25055), .Z(n25053) );
  IV U29812 ( .A(n25056), .Z(n25055) );
  NAND U29813 ( .A(n25056), .B(n25054), .Z(n25050) );
  AND U29814 ( .A(n25057), .B(n25058), .Z(n25031) );
  NAND U29815 ( .A(n25059), .B(n25060), .Z(n25058) );
  OR U29816 ( .A(n25061), .B(n25062), .Z(n25060) );
  NAND U29817 ( .A(n25062), .B(n25061), .Z(n25057) );
  IV U29818 ( .A(n25063), .Z(n25062) );
  NAND U29819 ( .A(n25064), .B(n25065), .Z(n25034) );
  NANDN U29820 ( .A(n25066), .B(n25067), .Z(n25065) );
  NAND U29821 ( .A(n25068), .B(n25069), .Z(n25067) );
  OR U29822 ( .A(n25069), .B(n25068), .Z(n25064) );
  IV U29823 ( .A(n25070), .Z(n25068) );
  AND U29824 ( .A(n25071), .B(n25072), .Z(n25037) );
  NAND U29825 ( .A(n25073), .B(n25074), .Z(n25072) );
  NANDN U29826 ( .A(n25075), .B(n25076), .Z(n25074) );
  NANDN U29827 ( .A(n25076), .B(n25075), .Z(n25071) );
  XOR U29828 ( .A(n25047), .B(n25077), .Z(n25039) );
  XNOR U29829 ( .A(n25044), .B(n25046), .Z(n25077) );
  AND U29830 ( .A(n25078), .B(n25079), .Z(n25046) );
  NANDN U29831 ( .A(n25080), .B(n25081), .Z(n25079) );
  NANDN U29832 ( .A(n25082), .B(n25083), .Z(n25081) );
  IV U29833 ( .A(n25084), .Z(n25083) );
  NAND U29834 ( .A(n25084), .B(n25082), .Z(n25078) );
  AND U29835 ( .A(n25085), .B(n25086), .Z(n25044) );
  NAND U29836 ( .A(n25087), .B(n25088), .Z(n25086) );
  OR U29837 ( .A(n25089), .B(n25090), .Z(n25088) );
  NAND U29838 ( .A(n25090), .B(n25089), .Z(n25085) );
  IV U29839 ( .A(n25091), .Z(n25090) );
  NAND U29840 ( .A(n25092), .B(n25093), .Z(n25047) );
  NANDN U29841 ( .A(n25094), .B(n25095), .Z(n25093) );
  NAND U29842 ( .A(n25096), .B(n25097), .Z(n25095) );
  OR U29843 ( .A(n25097), .B(n25096), .Z(n25092) );
  IV U29844 ( .A(n25098), .Z(n25096) );
  XOR U29845 ( .A(n25073), .B(n25099), .Z(N28086) );
  XNOR U29846 ( .A(n25076), .B(n25075), .Z(n25099) );
  XNOR U29847 ( .A(n25087), .B(n25100), .Z(n25075) );
  XOR U29848 ( .A(n25091), .B(n25089), .Z(n25100) );
  XOR U29849 ( .A(n25097), .B(n25101), .Z(n25089) );
  XOR U29850 ( .A(n25094), .B(n25098), .Z(n25101) );
  NAND U29851 ( .A(n25102), .B(n25103), .Z(n25098) );
  NAND U29852 ( .A(n25104), .B(n25105), .Z(n25103) );
  NAND U29853 ( .A(n25106), .B(n25107), .Z(n25102) );
  AND U29854 ( .A(n25108), .B(n25109), .Z(n25094) );
  NAND U29855 ( .A(n25110), .B(n25111), .Z(n25109) );
  NAND U29856 ( .A(n25112), .B(n25113), .Z(n25108) );
  NANDN U29857 ( .A(n25114), .B(n25115), .Z(n25097) );
  NANDN U29858 ( .A(n25116), .B(n25117), .Z(n25091) );
  XNOR U29859 ( .A(n25082), .B(n25118), .Z(n25087) );
  XOR U29860 ( .A(n25080), .B(n25084), .Z(n25118) );
  NAND U29861 ( .A(n25119), .B(n25120), .Z(n25084) );
  NAND U29862 ( .A(n25121), .B(n25122), .Z(n25120) );
  NAND U29863 ( .A(n25123), .B(n25124), .Z(n25119) );
  AND U29864 ( .A(n25125), .B(n25126), .Z(n25080) );
  NAND U29865 ( .A(n25127), .B(n25128), .Z(n25126) );
  NAND U29866 ( .A(n25129), .B(n25130), .Z(n25125) );
  AND U29867 ( .A(n25131), .B(n25132), .Z(n25082) );
  NAND U29868 ( .A(n25133), .B(n25134), .Z(n25076) );
  XNOR U29869 ( .A(n25059), .B(n25135), .Z(n25073) );
  XOR U29870 ( .A(n25063), .B(n25061), .Z(n25135) );
  XOR U29871 ( .A(n25069), .B(n25136), .Z(n25061) );
  XOR U29872 ( .A(n25066), .B(n25070), .Z(n25136) );
  NAND U29873 ( .A(n25137), .B(n25138), .Z(n25070) );
  NAND U29874 ( .A(n25139), .B(n25140), .Z(n25138) );
  NAND U29875 ( .A(n25141), .B(n25142), .Z(n25137) );
  AND U29876 ( .A(n25143), .B(n25144), .Z(n25066) );
  NAND U29877 ( .A(n25145), .B(n25146), .Z(n25144) );
  NAND U29878 ( .A(n25147), .B(n25148), .Z(n25143) );
  NANDN U29879 ( .A(n25149), .B(n25150), .Z(n25069) );
  NANDN U29880 ( .A(n25151), .B(n25152), .Z(n25063) );
  XNOR U29881 ( .A(n25054), .B(n25153), .Z(n25059) );
  XOR U29882 ( .A(n25052), .B(n25056), .Z(n25153) );
  NAND U29883 ( .A(n25154), .B(n25155), .Z(n25056) );
  NAND U29884 ( .A(n25156), .B(n25157), .Z(n25155) );
  NAND U29885 ( .A(n25158), .B(n25159), .Z(n25154) );
  AND U29886 ( .A(n25160), .B(n25161), .Z(n25052) );
  NAND U29887 ( .A(n25162), .B(n25163), .Z(n25161) );
  NAND U29888 ( .A(n25164), .B(n25165), .Z(n25160) );
  AND U29889 ( .A(n25166), .B(n25167), .Z(n25054) );
  XOR U29890 ( .A(n25134), .B(n25133), .Z(N28085) );
  XNOR U29891 ( .A(n25152), .B(n25151), .Z(n25133) );
  XNOR U29892 ( .A(n25166), .B(n25167), .Z(n25151) );
  XOR U29893 ( .A(n25163), .B(n25162), .Z(n25167) );
  XOR U29894 ( .A(y[315]), .B(x[315]), .Z(n25162) );
  XOR U29895 ( .A(n25165), .B(n25164), .Z(n25163) );
  XOR U29896 ( .A(y[317]), .B(x[317]), .Z(n25164) );
  XOR U29897 ( .A(y[316]), .B(x[316]), .Z(n25165) );
  XOR U29898 ( .A(n25157), .B(n25156), .Z(n25166) );
  XOR U29899 ( .A(n25159), .B(n25158), .Z(n25156) );
  XOR U29900 ( .A(y[314]), .B(x[314]), .Z(n25158) );
  XOR U29901 ( .A(y[313]), .B(x[313]), .Z(n25159) );
  XOR U29902 ( .A(y[312]), .B(x[312]), .Z(n25157) );
  XNOR U29903 ( .A(n25150), .B(n25149), .Z(n25152) );
  XNOR U29904 ( .A(n25146), .B(n25145), .Z(n25149) );
  XOR U29905 ( .A(n25148), .B(n25147), .Z(n25145) );
  XOR U29906 ( .A(y[311]), .B(x[311]), .Z(n25147) );
  XOR U29907 ( .A(y[310]), .B(x[310]), .Z(n25148) );
  XOR U29908 ( .A(y[309]), .B(x[309]), .Z(n25146) );
  XOR U29909 ( .A(n25140), .B(n25139), .Z(n25150) );
  XOR U29910 ( .A(n25142), .B(n25141), .Z(n25139) );
  XOR U29911 ( .A(y[308]), .B(x[308]), .Z(n25141) );
  XOR U29912 ( .A(y[307]), .B(x[307]), .Z(n25142) );
  XOR U29913 ( .A(y[306]), .B(x[306]), .Z(n25140) );
  XNOR U29914 ( .A(n25117), .B(n25116), .Z(n25134) );
  XNOR U29915 ( .A(n25131), .B(n25132), .Z(n25116) );
  XOR U29916 ( .A(n25128), .B(n25127), .Z(n25132) );
  XOR U29917 ( .A(y[303]), .B(x[303]), .Z(n25127) );
  XOR U29918 ( .A(n25130), .B(n25129), .Z(n25128) );
  XOR U29919 ( .A(y[305]), .B(x[305]), .Z(n25129) );
  XOR U29920 ( .A(y[304]), .B(x[304]), .Z(n25130) );
  XOR U29921 ( .A(n25122), .B(n25121), .Z(n25131) );
  XOR U29922 ( .A(n25124), .B(n25123), .Z(n25121) );
  XOR U29923 ( .A(y[302]), .B(x[302]), .Z(n25123) );
  XOR U29924 ( .A(y[301]), .B(x[301]), .Z(n25124) );
  XOR U29925 ( .A(y[300]), .B(x[300]), .Z(n25122) );
  XNOR U29926 ( .A(n25115), .B(n25114), .Z(n25117) );
  XNOR U29927 ( .A(n25111), .B(n25110), .Z(n25114) );
  XOR U29928 ( .A(n25113), .B(n25112), .Z(n25110) );
  XOR U29929 ( .A(y[299]), .B(x[299]), .Z(n25112) );
  XOR U29930 ( .A(y[298]), .B(x[298]), .Z(n25113) );
  XOR U29931 ( .A(y[297]), .B(x[297]), .Z(n25111) );
  XOR U29932 ( .A(n25105), .B(n25104), .Z(n25115) );
  XOR U29933 ( .A(n25107), .B(n25106), .Z(n25104) );
  XOR U29934 ( .A(y[296]), .B(x[296]), .Z(n25106) );
  XOR U29935 ( .A(y[295]), .B(x[295]), .Z(n25107) );
  XOR U29936 ( .A(y[294]), .B(x[294]), .Z(n25105) );
  NAND U29937 ( .A(n25168), .B(n25169), .Z(N28077) );
  NAND U29938 ( .A(n25170), .B(n25171), .Z(n25169) );
  NANDN U29939 ( .A(n25172), .B(n25173), .Z(n25171) );
  NANDN U29940 ( .A(n25173), .B(n25172), .Z(n25168) );
  XOR U29941 ( .A(n25172), .B(n25174), .Z(N28076) );
  XNOR U29942 ( .A(n25170), .B(n25173), .Z(n25174) );
  NAND U29943 ( .A(n25175), .B(n25176), .Z(n25173) );
  NAND U29944 ( .A(n25177), .B(n25178), .Z(n25176) );
  NANDN U29945 ( .A(n25179), .B(n25180), .Z(n25178) );
  NANDN U29946 ( .A(n25180), .B(n25179), .Z(n25175) );
  AND U29947 ( .A(n25181), .B(n25182), .Z(n25170) );
  NAND U29948 ( .A(n25183), .B(n25184), .Z(n25182) );
  OR U29949 ( .A(n25185), .B(n25186), .Z(n25184) );
  NAND U29950 ( .A(n25186), .B(n25185), .Z(n25181) );
  IV U29951 ( .A(n25187), .Z(n25186) );
  AND U29952 ( .A(n25188), .B(n25189), .Z(n25172) );
  NAND U29953 ( .A(n25190), .B(n25191), .Z(n25189) );
  NANDN U29954 ( .A(n25192), .B(n25193), .Z(n25191) );
  NANDN U29955 ( .A(n25193), .B(n25192), .Z(n25188) );
  XOR U29956 ( .A(n25185), .B(n25194), .Z(N28075) );
  XOR U29957 ( .A(n25183), .B(n25187), .Z(n25194) );
  XNOR U29958 ( .A(n25180), .B(n25195), .Z(n25187) );
  XNOR U29959 ( .A(n25177), .B(n25179), .Z(n25195) );
  AND U29960 ( .A(n25196), .B(n25197), .Z(n25179) );
  NANDN U29961 ( .A(n25198), .B(n25199), .Z(n25197) );
  NANDN U29962 ( .A(n25200), .B(n25201), .Z(n25199) );
  IV U29963 ( .A(n25202), .Z(n25201) );
  NAND U29964 ( .A(n25202), .B(n25200), .Z(n25196) );
  AND U29965 ( .A(n25203), .B(n25204), .Z(n25177) );
  NAND U29966 ( .A(n25205), .B(n25206), .Z(n25204) );
  OR U29967 ( .A(n25207), .B(n25208), .Z(n25206) );
  NAND U29968 ( .A(n25208), .B(n25207), .Z(n25203) );
  IV U29969 ( .A(n25209), .Z(n25208) );
  NAND U29970 ( .A(n25210), .B(n25211), .Z(n25180) );
  NANDN U29971 ( .A(n25212), .B(n25213), .Z(n25211) );
  NAND U29972 ( .A(n25214), .B(n25215), .Z(n25213) );
  OR U29973 ( .A(n25215), .B(n25214), .Z(n25210) );
  IV U29974 ( .A(n25216), .Z(n25214) );
  AND U29975 ( .A(n25217), .B(n25218), .Z(n25183) );
  NAND U29976 ( .A(n25219), .B(n25220), .Z(n25218) );
  NANDN U29977 ( .A(n25221), .B(n25222), .Z(n25220) );
  NANDN U29978 ( .A(n25222), .B(n25221), .Z(n25217) );
  XOR U29979 ( .A(n25193), .B(n25223), .Z(n25185) );
  XNOR U29980 ( .A(n25190), .B(n25192), .Z(n25223) );
  AND U29981 ( .A(n25224), .B(n25225), .Z(n25192) );
  NANDN U29982 ( .A(n25226), .B(n25227), .Z(n25225) );
  NANDN U29983 ( .A(n25228), .B(n25229), .Z(n25227) );
  IV U29984 ( .A(n25230), .Z(n25229) );
  NAND U29985 ( .A(n25230), .B(n25228), .Z(n25224) );
  AND U29986 ( .A(n25231), .B(n25232), .Z(n25190) );
  NAND U29987 ( .A(n25233), .B(n25234), .Z(n25232) );
  OR U29988 ( .A(n25235), .B(n25236), .Z(n25234) );
  NAND U29989 ( .A(n25236), .B(n25235), .Z(n25231) );
  IV U29990 ( .A(n25237), .Z(n25236) );
  NAND U29991 ( .A(n25238), .B(n25239), .Z(n25193) );
  NANDN U29992 ( .A(n25240), .B(n25241), .Z(n25239) );
  NAND U29993 ( .A(n25242), .B(n25243), .Z(n25241) );
  OR U29994 ( .A(n25243), .B(n25242), .Z(n25238) );
  IV U29995 ( .A(n25244), .Z(n25242) );
  XOR U29996 ( .A(n25219), .B(n25245), .Z(N28074) );
  XNOR U29997 ( .A(n25222), .B(n25221), .Z(n25245) );
  XNOR U29998 ( .A(n25233), .B(n25246), .Z(n25221) );
  XOR U29999 ( .A(n25237), .B(n25235), .Z(n25246) );
  XOR U30000 ( .A(n25243), .B(n25247), .Z(n25235) );
  XOR U30001 ( .A(n25240), .B(n25244), .Z(n25247) );
  NAND U30002 ( .A(n25248), .B(n25249), .Z(n25244) );
  NAND U30003 ( .A(n25250), .B(n25251), .Z(n25249) );
  NAND U30004 ( .A(n25252), .B(n25253), .Z(n25248) );
  AND U30005 ( .A(n25254), .B(n25255), .Z(n25240) );
  NAND U30006 ( .A(n25256), .B(n25257), .Z(n25255) );
  NAND U30007 ( .A(n25258), .B(n25259), .Z(n25254) );
  NANDN U30008 ( .A(n25260), .B(n25261), .Z(n25243) );
  NANDN U30009 ( .A(n25262), .B(n25263), .Z(n25237) );
  XNOR U30010 ( .A(n25228), .B(n25264), .Z(n25233) );
  XOR U30011 ( .A(n25226), .B(n25230), .Z(n25264) );
  NAND U30012 ( .A(n25265), .B(n25266), .Z(n25230) );
  NAND U30013 ( .A(n25267), .B(n25268), .Z(n25266) );
  NAND U30014 ( .A(n25269), .B(n25270), .Z(n25265) );
  AND U30015 ( .A(n25271), .B(n25272), .Z(n25226) );
  NAND U30016 ( .A(n25273), .B(n25274), .Z(n25272) );
  NAND U30017 ( .A(n25275), .B(n25276), .Z(n25271) );
  AND U30018 ( .A(n25277), .B(n25278), .Z(n25228) );
  NAND U30019 ( .A(n25279), .B(n25280), .Z(n25222) );
  XNOR U30020 ( .A(n25205), .B(n25281), .Z(n25219) );
  XOR U30021 ( .A(n25209), .B(n25207), .Z(n25281) );
  XOR U30022 ( .A(n25215), .B(n25282), .Z(n25207) );
  XOR U30023 ( .A(n25212), .B(n25216), .Z(n25282) );
  NAND U30024 ( .A(n25283), .B(n25284), .Z(n25216) );
  NAND U30025 ( .A(n25285), .B(n25286), .Z(n25284) );
  NAND U30026 ( .A(n25287), .B(n25288), .Z(n25283) );
  AND U30027 ( .A(n25289), .B(n25290), .Z(n25212) );
  NAND U30028 ( .A(n25291), .B(n25292), .Z(n25290) );
  NAND U30029 ( .A(n25293), .B(n25294), .Z(n25289) );
  NANDN U30030 ( .A(n25295), .B(n25296), .Z(n25215) );
  NANDN U30031 ( .A(n25297), .B(n25298), .Z(n25209) );
  XNOR U30032 ( .A(n25200), .B(n25299), .Z(n25205) );
  XOR U30033 ( .A(n25198), .B(n25202), .Z(n25299) );
  NAND U30034 ( .A(n25300), .B(n25301), .Z(n25202) );
  NAND U30035 ( .A(n25302), .B(n25303), .Z(n25301) );
  NAND U30036 ( .A(n25304), .B(n25305), .Z(n25300) );
  AND U30037 ( .A(n25306), .B(n25307), .Z(n25198) );
  NAND U30038 ( .A(n25308), .B(n25309), .Z(n25307) );
  NAND U30039 ( .A(n25310), .B(n25311), .Z(n25306) );
  AND U30040 ( .A(n25312), .B(n25313), .Z(n25200) );
  XOR U30041 ( .A(n25280), .B(n25279), .Z(N28073) );
  XNOR U30042 ( .A(n25298), .B(n25297), .Z(n25279) );
  XNOR U30043 ( .A(n25312), .B(n25313), .Z(n25297) );
  XOR U30044 ( .A(n25309), .B(n25308), .Z(n25313) );
  XOR U30045 ( .A(y[291]), .B(x[291]), .Z(n25308) );
  XOR U30046 ( .A(n25311), .B(n25310), .Z(n25309) );
  XOR U30047 ( .A(y[293]), .B(x[293]), .Z(n25310) );
  XOR U30048 ( .A(y[292]), .B(x[292]), .Z(n25311) );
  XOR U30049 ( .A(n25303), .B(n25302), .Z(n25312) );
  XOR U30050 ( .A(n25305), .B(n25304), .Z(n25302) );
  XOR U30051 ( .A(y[290]), .B(x[290]), .Z(n25304) );
  XOR U30052 ( .A(y[289]), .B(x[289]), .Z(n25305) );
  XOR U30053 ( .A(y[288]), .B(x[288]), .Z(n25303) );
  XNOR U30054 ( .A(n25296), .B(n25295), .Z(n25298) );
  XNOR U30055 ( .A(n25292), .B(n25291), .Z(n25295) );
  XOR U30056 ( .A(n25294), .B(n25293), .Z(n25291) );
  XOR U30057 ( .A(y[287]), .B(x[287]), .Z(n25293) );
  XOR U30058 ( .A(y[286]), .B(x[286]), .Z(n25294) );
  XOR U30059 ( .A(y[285]), .B(x[285]), .Z(n25292) );
  XOR U30060 ( .A(n25286), .B(n25285), .Z(n25296) );
  XOR U30061 ( .A(n25288), .B(n25287), .Z(n25285) );
  XOR U30062 ( .A(y[284]), .B(x[284]), .Z(n25287) );
  XOR U30063 ( .A(y[283]), .B(x[283]), .Z(n25288) );
  XOR U30064 ( .A(y[282]), .B(x[282]), .Z(n25286) );
  XNOR U30065 ( .A(n25263), .B(n25262), .Z(n25280) );
  XNOR U30066 ( .A(n25277), .B(n25278), .Z(n25262) );
  XOR U30067 ( .A(n25274), .B(n25273), .Z(n25278) );
  XOR U30068 ( .A(y[279]), .B(x[279]), .Z(n25273) );
  XOR U30069 ( .A(n25276), .B(n25275), .Z(n25274) );
  XOR U30070 ( .A(y[281]), .B(x[281]), .Z(n25275) );
  XOR U30071 ( .A(y[280]), .B(x[280]), .Z(n25276) );
  XOR U30072 ( .A(n25268), .B(n25267), .Z(n25277) );
  XOR U30073 ( .A(n25270), .B(n25269), .Z(n25267) );
  XOR U30074 ( .A(y[278]), .B(x[278]), .Z(n25269) );
  XOR U30075 ( .A(y[277]), .B(x[277]), .Z(n25270) );
  XOR U30076 ( .A(y[276]), .B(x[276]), .Z(n25268) );
  XNOR U30077 ( .A(n25261), .B(n25260), .Z(n25263) );
  XNOR U30078 ( .A(n25257), .B(n25256), .Z(n25260) );
  XOR U30079 ( .A(n25259), .B(n25258), .Z(n25256) );
  XOR U30080 ( .A(y[275]), .B(x[275]), .Z(n25258) );
  XOR U30081 ( .A(y[274]), .B(x[274]), .Z(n25259) );
  XOR U30082 ( .A(y[273]), .B(x[273]), .Z(n25257) );
  XOR U30083 ( .A(n25251), .B(n25250), .Z(n25261) );
  XOR U30084 ( .A(n25253), .B(n25252), .Z(n25250) );
  XOR U30085 ( .A(y[272]), .B(x[272]), .Z(n25252) );
  XOR U30086 ( .A(y[271]), .B(x[271]), .Z(n25253) );
  XOR U30087 ( .A(y[270]), .B(x[270]), .Z(n25251) );
  NAND U30088 ( .A(n25314), .B(n25315), .Z(N28065) );
  NAND U30089 ( .A(n25316), .B(n25317), .Z(n25315) );
  NANDN U30090 ( .A(n25318), .B(n25319), .Z(n25317) );
  NANDN U30091 ( .A(n25319), .B(n25318), .Z(n25314) );
  XOR U30092 ( .A(n25318), .B(n25320), .Z(N28064) );
  XNOR U30093 ( .A(n25316), .B(n25319), .Z(n25320) );
  NAND U30094 ( .A(n25321), .B(n25322), .Z(n25319) );
  NAND U30095 ( .A(n25323), .B(n25324), .Z(n25322) );
  NANDN U30096 ( .A(n25325), .B(n25326), .Z(n25324) );
  NANDN U30097 ( .A(n25326), .B(n25325), .Z(n25321) );
  AND U30098 ( .A(n25327), .B(n25328), .Z(n25316) );
  NAND U30099 ( .A(n25329), .B(n25330), .Z(n25328) );
  OR U30100 ( .A(n25331), .B(n25332), .Z(n25330) );
  NAND U30101 ( .A(n25332), .B(n25331), .Z(n25327) );
  IV U30102 ( .A(n25333), .Z(n25332) );
  AND U30103 ( .A(n25334), .B(n25335), .Z(n25318) );
  NAND U30104 ( .A(n25336), .B(n25337), .Z(n25335) );
  NANDN U30105 ( .A(n25338), .B(n25339), .Z(n25337) );
  NANDN U30106 ( .A(n25339), .B(n25338), .Z(n25334) );
  XOR U30107 ( .A(n25331), .B(n25340), .Z(N28063) );
  XOR U30108 ( .A(n25329), .B(n25333), .Z(n25340) );
  XNOR U30109 ( .A(n25326), .B(n25341), .Z(n25333) );
  XNOR U30110 ( .A(n25323), .B(n25325), .Z(n25341) );
  AND U30111 ( .A(n25342), .B(n25343), .Z(n25325) );
  NANDN U30112 ( .A(n25344), .B(n25345), .Z(n25343) );
  NANDN U30113 ( .A(n25346), .B(n25347), .Z(n25345) );
  IV U30114 ( .A(n25348), .Z(n25347) );
  NAND U30115 ( .A(n25348), .B(n25346), .Z(n25342) );
  AND U30116 ( .A(n25349), .B(n25350), .Z(n25323) );
  NAND U30117 ( .A(n25351), .B(n25352), .Z(n25350) );
  OR U30118 ( .A(n25353), .B(n25354), .Z(n25352) );
  NAND U30119 ( .A(n25354), .B(n25353), .Z(n25349) );
  IV U30120 ( .A(n25355), .Z(n25354) );
  NAND U30121 ( .A(n25356), .B(n25357), .Z(n25326) );
  NANDN U30122 ( .A(n25358), .B(n25359), .Z(n25357) );
  NAND U30123 ( .A(n25360), .B(n25361), .Z(n25359) );
  OR U30124 ( .A(n25361), .B(n25360), .Z(n25356) );
  IV U30125 ( .A(n25362), .Z(n25360) );
  AND U30126 ( .A(n25363), .B(n25364), .Z(n25329) );
  NAND U30127 ( .A(n25365), .B(n25366), .Z(n25364) );
  NANDN U30128 ( .A(n25367), .B(n25368), .Z(n25366) );
  NANDN U30129 ( .A(n25368), .B(n25367), .Z(n25363) );
  XOR U30130 ( .A(n25339), .B(n25369), .Z(n25331) );
  XNOR U30131 ( .A(n25336), .B(n25338), .Z(n25369) );
  AND U30132 ( .A(n25370), .B(n25371), .Z(n25338) );
  NANDN U30133 ( .A(n25372), .B(n25373), .Z(n25371) );
  NANDN U30134 ( .A(n25374), .B(n25375), .Z(n25373) );
  IV U30135 ( .A(n25376), .Z(n25375) );
  NAND U30136 ( .A(n25376), .B(n25374), .Z(n25370) );
  AND U30137 ( .A(n25377), .B(n25378), .Z(n25336) );
  NAND U30138 ( .A(n25379), .B(n25380), .Z(n25378) );
  OR U30139 ( .A(n25381), .B(n25382), .Z(n25380) );
  NAND U30140 ( .A(n25382), .B(n25381), .Z(n25377) );
  IV U30141 ( .A(n25383), .Z(n25382) );
  NAND U30142 ( .A(n25384), .B(n25385), .Z(n25339) );
  NANDN U30143 ( .A(n25386), .B(n25387), .Z(n25385) );
  NAND U30144 ( .A(n25388), .B(n25389), .Z(n25387) );
  OR U30145 ( .A(n25389), .B(n25388), .Z(n25384) );
  IV U30146 ( .A(n25390), .Z(n25388) );
  XOR U30147 ( .A(n25365), .B(n25391), .Z(N28062) );
  XNOR U30148 ( .A(n25368), .B(n25367), .Z(n25391) );
  XNOR U30149 ( .A(n25379), .B(n25392), .Z(n25367) );
  XOR U30150 ( .A(n25383), .B(n25381), .Z(n25392) );
  XOR U30151 ( .A(n25389), .B(n25393), .Z(n25381) );
  XOR U30152 ( .A(n25386), .B(n25390), .Z(n25393) );
  NAND U30153 ( .A(n25394), .B(n25395), .Z(n25390) );
  NAND U30154 ( .A(n25396), .B(n25397), .Z(n25395) );
  NAND U30155 ( .A(n25398), .B(n25399), .Z(n25394) );
  AND U30156 ( .A(n25400), .B(n25401), .Z(n25386) );
  NAND U30157 ( .A(n25402), .B(n25403), .Z(n25401) );
  NAND U30158 ( .A(n25404), .B(n25405), .Z(n25400) );
  NANDN U30159 ( .A(n25406), .B(n25407), .Z(n25389) );
  NANDN U30160 ( .A(n25408), .B(n25409), .Z(n25383) );
  XNOR U30161 ( .A(n25374), .B(n25410), .Z(n25379) );
  XOR U30162 ( .A(n25372), .B(n25376), .Z(n25410) );
  NAND U30163 ( .A(n25411), .B(n25412), .Z(n25376) );
  NAND U30164 ( .A(n25413), .B(n25414), .Z(n25412) );
  NAND U30165 ( .A(n25415), .B(n25416), .Z(n25411) );
  AND U30166 ( .A(n25417), .B(n25418), .Z(n25372) );
  NAND U30167 ( .A(n25419), .B(n25420), .Z(n25418) );
  NAND U30168 ( .A(n25421), .B(n25422), .Z(n25417) );
  AND U30169 ( .A(n25423), .B(n25424), .Z(n25374) );
  NAND U30170 ( .A(n25425), .B(n25426), .Z(n25368) );
  XNOR U30171 ( .A(n25351), .B(n25427), .Z(n25365) );
  XOR U30172 ( .A(n25355), .B(n25353), .Z(n25427) );
  XOR U30173 ( .A(n25361), .B(n25428), .Z(n25353) );
  XOR U30174 ( .A(n25358), .B(n25362), .Z(n25428) );
  NAND U30175 ( .A(n25429), .B(n25430), .Z(n25362) );
  NAND U30176 ( .A(n25431), .B(n25432), .Z(n25430) );
  NAND U30177 ( .A(n25433), .B(n25434), .Z(n25429) );
  AND U30178 ( .A(n25435), .B(n25436), .Z(n25358) );
  NAND U30179 ( .A(n25437), .B(n25438), .Z(n25436) );
  NAND U30180 ( .A(n25439), .B(n25440), .Z(n25435) );
  NANDN U30181 ( .A(n25441), .B(n25442), .Z(n25361) );
  NANDN U30182 ( .A(n25443), .B(n25444), .Z(n25355) );
  XNOR U30183 ( .A(n25346), .B(n25445), .Z(n25351) );
  XOR U30184 ( .A(n25344), .B(n25348), .Z(n25445) );
  NAND U30185 ( .A(n25446), .B(n25447), .Z(n25348) );
  NAND U30186 ( .A(n25448), .B(n25449), .Z(n25447) );
  NAND U30187 ( .A(n25450), .B(n25451), .Z(n25446) );
  AND U30188 ( .A(n25452), .B(n25453), .Z(n25344) );
  NAND U30189 ( .A(n25454), .B(n25455), .Z(n25453) );
  NAND U30190 ( .A(n25456), .B(n25457), .Z(n25452) );
  AND U30191 ( .A(n25458), .B(n25459), .Z(n25346) );
  XOR U30192 ( .A(n25426), .B(n25425), .Z(N28061) );
  XNOR U30193 ( .A(n25444), .B(n25443), .Z(n25425) );
  XNOR U30194 ( .A(n25458), .B(n25459), .Z(n25443) );
  XOR U30195 ( .A(n25455), .B(n25454), .Z(n25459) );
  XOR U30196 ( .A(y[267]), .B(x[267]), .Z(n25454) );
  XOR U30197 ( .A(n25457), .B(n25456), .Z(n25455) );
  XOR U30198 ( .A(y[269]), .B(x[269]), .Z(n25456) );
  XOR U30199 ( .A(y[268]), .B(x[268]), .Z(n25457) );
  XOR U30200 ( .A(n25449), .B(n25448), .Z(n25458) );
  XOR U30201 ( .A(n25451), .B(n25450), .Z(n25448) );
  XOR U30202 ( .A(y[266]), .B(x[266]), .Z(n25450) );
  XOR U30203 ( .A(y[265]), .B(x[265]), .Z(n25451) );
  XOR U30204 ( .A(y[264]), .B(x[264]), .Z(n25449) );
  XNOR U30205 ( .A(n25442), .B(n25441), .Z(n25444) );
  XNOR U30206 ( .A(n25438), .B(n25437), .Z(n25441) );
  XOR U30207 ( .A(n25440), .B(n25439), .Z(n25437) );
  XOR U30208 ( .A(y[263]), .B(x[263]), .Z(n25439) );
  XOR U30209 ( .A(y[262]), .B(x[262]), .Z(n25440) );
  XOR U30210 ( .A(y[261]), .B(x[261]), .Z(n25438) );
  XOR U30211 ( .A(n25432), .B(n25431), .Z(n25442) );
  XOR U30212 ( .A(n25434), .B(n25433), .Z(n25431) );
  XOR U30213 ( .A(y[260]), .B(x[260]), .Z(n25433) );
  XOR U30214 ( .A(y[259]), .B(x[259]), .Z(n25434) );
  XOR U30215 ( .A(y[258]), .B(x[258]), .Z(n25432) );
  XNOR U30216 ( .A(n25409), .B(n25408), .Z(n25426) );
  XNOR U30217 ( .A(n25423), .B(n25424), .Z(n25408) );
  XOR U30218 ( .A(n25420), .B(n25419), .Z(n25424) );
  XOR U30219 ( .A(y[255]), .B(x[255]), .Z(n25419) );
  XOR U30220 ( .A(n25422), .B(n25421), .Z(n25420) );
  XOR U30221 ( .A(y[257]), .B(x[257]), .Z(n25421) );
  XOR U30222 ( .A(y[256]), .B(x[256]), .Z(n25422) );
  XOR U30223 ( .A(n25414), .B(n25413), .Z(n25423) );
  XOR U30224 ( .A(n25416), .B(n25415), .Z(n25413) );
  XOR U30225 ( .A(y[254]), .B(x[254]), .Z(n25415) );
  XOR U30226 ( .A(y[253]), .B(x[253]), .Z(n25416) );
  XOR U30227 ( .A(y[252]), .B(x[252]), .Z(n25414) );
  XNOR U30228 ( .A(n25407), .B(n25406), .Z(n25409) );
  XNOR U30229 ( .A(n25403), .B(n25402), .Z(n25406) );
  XOR U30230 ( .A(n25405), .B(n25404), .Z(n25402) );
  XOR U30231 ( .A(y[251]), .B(x[251]), .Z(n25404) );
  XOR U30232 ( .A(y[250]), .B(x[250]), .Z(n25405) );
  XOR U30233 ( .A(y[249]), .B(x[249]), .Z(n25403) );
  XOR U30234 ( .A(n25397), .B(n25396), .Z(n25407) );
  XOR U30235 ( .A(n25399), .B(n25398), .Z(n25396) );
  XOR U30236 ( .A(y[248]), .B(x[248]), .Z(n25398) );
  XOR U30237 ( .A(y[247]), .B(x[247]), .Z(n25399) );
  XOR U30238 ( .A(y[246]), .B(x[246]), .Z(n25397) );
  NAND U30239 ( .A(n25460), .B(n25461), .Z(N28053) );
  NAND U30240 ( .A(n25462), .B(n25463), .Z(n25461) );
  NANDN U30241 ( .A(n25464), .B(n25465), .Z(n25463) );
  NANDN U30242 ( .A(n25465), .B(n25464), .Z(n25460) );
  XOR U30243 ( .A(n25464), .B(n25466), .Z(N28052) );
  XNOR U30244 ( .A(n25462), .B(n25465), .Z(n25466) );
  NAND U30245 ( .A(n25467), .B(n25468), .Z(n25465) );
  NAND U30246 ( .A(n25469), .B(n25470), .Z(n25468) );
  NANDN U30247 ( .A(n25471), .B(n25472), .Z(n25470) );
  NANDN U30248 ( .A(n25472), .B(n25471), .Z(n25467) );
  AND U30249 ( .A(n25473), .B(n25474), .Z(n25462) );
  NAND U30250 ( .A(n25475), .B(n25476), .Z(n25474) );
  OR U30251 ( .A(n25477), .B(n25478), .Z(n25476) );
  NAND U30252 ( .A(n25478), .B(n25477), .Z(n25473) );
  IV U30253 ( .A(n25479), .Z(n25478) );
  AND U30254 ( .A(n25480), .B(n25481), .Z(n25464) );
  NAND U30255 ( .A(n25482), .B(n25483), .Z(n25481) );
  NANDN U30256 ( .A(n25484), .B(n25485), .Z(n25483) );
  NANDN U30257 ( .A(n25485), .B(n25484), .Z(n25480) );
  XOR U30258 ( .A(n25477), .B(n25486), .Z(N28051) );
  XOR U30259 ( .A(n25475), .B(n25479), .Z(n25486) );
  XNOR U30260 ( .A(n25472), .B(n25487), .Z(n25479) );
  XNOR U30261 ( .A(n25469), .B(n25471), .Z(n25487) );
  AND U30262 ( .A(n25488), .B(n25489), .Z(n25471) );
  NANDN U30263 ( .A(n25490), .B(n25491), .Z(n25489) );
  NANDN U30264 ( .A(n25492), .B(n25493), .Z(n25491) );
  IV U30265 ( .A(n25494), .Z(n25493) );
  NAND U30266 ( .A(n25494), .B(n25492), .Z(n25488) );
  AND U30267 ( .A(n25495), .B(n25496), .Z(n25469) );
  NAND U30268 ( .A(n25497), .B(n25498), .Z(n25496) );
  OR U30269 ( .A(n25499), .B(n25500), .Z(n25498) );
  NAND U30270 ( .A(n25500), .B(n25499), .Z(n25495) );
  IV U30271 ( .A(n25501), .Z(n25500) );
  NAND U30272 ( .A(n25502), .B(n25503), .Z(n25472) );
  NANDN U30273 ( .A(n25504), .B(n25505), .Z(n25503) );
  NAND U30274 ( .A(n25506), .B(n25507), .Z(n25505) );
  OR U30275 ( .A(n25507), .B(n25506), .Z(n25502) );
  IV U30276 ( .A(n25508), .Z(n25506) );
  AND U30277 ( .A(n25509), .B(n25510), .Z(n25475) );
  NAND U30278 ( .A(n25511), .B(n25512), .Z(n25510) );
  NANDN U30279 ( .A(n25513), .B(n25514), .Z(n25512) );
  NANDN U30280 ( .A(n25514), .B(n25513), .Z(n25509) );
  XOR U30281 ( .A(n25485), .B(n25515), .Z(n25477) );
  XNOR U30282 ( .A(n25482), .B(n25484), .Z(n25515) );
  AND U30283 ( .A(n25516), .B(n25517), .Z(n25484) );
  NANDN U30284 ( .A(n25518), .B(n25519), .Z(n25517) );
  NANDN U30285 ( .A(n25520), .B(n25521), .Z(n25519) );
  IV U30286 ( .A(n25522), .Z(n25521) );
  NAND U30287 ( .A(n25522), .B(n25520), .Z(n25516) );
  AND U30288 ( .A(n25523), .B(n25524), .Z(n25482) );
  NAND U30289 ( .A(n25525), .B(n25526), .Z(n25524) );
  OR U30290 ( .A(n25527), .B(n25528), .Z(n25526) );
  NAND U30291 ( .A(n25528), .B(n25527), .Z(n25523) );
  IV U30292 ( .A(n25529), .Z(n25528) );
  NAND U30293 ( .A(n25530), .B(n25531), .Z(n25485) );
  NANDN U30294 ( .A(n25532), .B(n25533), .Z(n25531) );
  NAND U30295 ( .A(n25534), .B(n25535), .Z(n25533) );
  OR U30296 ( .A(n25535), .B(n25534), .Z(n25530) );
  IV U30297 ( .A(n25536), .Z(n25534) );
  XOR U30298 ( .A(n25511), .B(n25537), .Z(N28050) );
  XNOR U30299 ( .A(n25514), .B(n25513), .Z(n25537) );
  XNOR U30300 ( .A(n25525), .B(n25538), .Z(n25513) );
  XOR U30301 ( .A(n25529), .B(n25527), .Z(n25538) );
  XOR U30302 ( .A(n25535), .B(n25539), .Z(n25527) );
  XOR U30303 ( .A(n25532), .B(n25536), .Z(n25539) );
  NAND U30304 ( .A(n25540), .B(n25541), .Z(n25536) );
  NAND U30305 ( .A(n25542), .B(n25543), .Z(n25541) );
  NAND U30306 ( .A(n25544), .B(n25545), .Z(n25540) );
  AND U30307 ( .A(n25546), .B(n25547), .Z(n25532) );
  NAND U30308 ( .A(n25548), .B(n25549), .Z(n25547) );
  NAND U30309 ( .A(n25550), .B(n25551), .Z(n25546) );
  NANDN U30310 ( .A(n25552), .B(n25553), .Z(n25535) );
  NANDN U30311 ( .A(n25554), .B(n25555), .Z(n25529) );
  XNOR U30312 ( .A(n25520), .B(n25556), .Z(n25525) );
  XOR U30313 ( .A(n25518), .B(n25522), .Z(n25556) );
  NAND U30314 ( .A(n25557), .B(n25558), .Z(n25522) );
  NAND U30315 ( .A(n25559), .B(n25560), .Z(n25558) );
  NAND U30316 ( .A(n25561), .B(n25562), .Z(n25557) );
  AND U30317 ( .A(n25563), .B(n25564), .Z(n25518) );
  NAND U30318 ( .A(n25565), .B(n25566), .Z(n25564) );
  NAND U30319 ( .A(n25567), .B(n25568), .Z(n25563) );
  AND U30320 ( .A(n25569), .B(n25570), .Z(n25520) );
  NAND U30321 ( .A(n25571), .B(n25572), .Z(n25514) );
  XNOR U30322 ( .A(n25497), .B(n25573), .Z(n25511) );
  XOR U30323 ( .A(n25501), .B(n25499), .Z(n25573) );
  XOR U30324 ( .A(n25507), .B(n25574), .Z(n25499) );
  XOR U30325 ( .A(n25504), .B(n25508), .Z(n25574) );
  NAND U30326 ( .A(n25575), .B(n25576), .Z(n25508) );
  NAND U30327 ( .A(n25577), .B(n25578), .Z(n25576) );
  NAND U30328 ( .A(n25579), .B(n25580), .Z(n25575) );
  AND U30329 ( .A(n25581), .B(n25582), .Z(n25504) );
  NAND U30330 ( .A(n25583), .B(n25584), .Z(n25582) );
  NAND U30331 ( .A(n25585), .B(n25586), .Z(n25581) );
  NANDN U30332 ( .A(n25587), .B(n25588), .Z(n25507) );
  NANDN U30333 ( .A(n25589), .B(n25590), .Z(n25501) );
  XNOR U30334 ( .A(n25492), .B(n25591), .Z(n25497) );
  XOR U30335 ( .A(n25490), .B(n25494), .Z(n25591) );
  NAND U30336 ( .A(n25592), .B(n25593), .Z(n25494) );
  NAND U30337 ( .A(n25594), .B(n25595), .Z(n25593) );
  NAND U30338 ( .A(n25596), .B(n25597), .Z(n25592) );
  AND U30339 ( .A(n25598), .B(n25599), .Z(n25490) );
  NAND U30340 ( .A(n25600), .B(n25601), .Z(n25599) );
  NAND U30341 ( .A(n25602), .B(n25603), .Z(n25598) );
  AND U30342 ( .A(n25604), .B(n25605), .Z(n25492) );
  XOR U30343 ( .A(n25572), .B(n25571), .Z(N28049) );
  XNOR U30344 ( .A(n25590), .B(n25589), .Z(n25571) );
  XNOR U30345 ( .A(n25604), .B(n25605), .Z(n25589) );
  XOR U30346 ( .A(n25601), .B(n25600), .Z(n25605) );
  XOR U30347 ( .A(y[243]), .B(x[243]), .Z(n25600) );
  XOR U30348 ( .A(n25603), .B(n25602), .Z(n25601) );
  XOR U30349 ( .A(y[245]), .B(x[245]), .Z(n25602) );
  XOR U30350 ( .A(y[244]), .B(x[244]), .Z(n25603) );
  XOR U30351 ( .A(n25595), .B(n25594), .Z(n25604) );
  XOR U30352 ( .A(n25597), .B(n25596), .Z(n25594) );
  XOR U30353 ( .A(y[242]), .B(x[242]), .Z(n25596) );
  XOR U30354 ( .A(y[241]), .B(x[241]), .Z(n25597) );
  XOR U30355 ( .A(y[240]), .B(x[240]), .Z(n25595) );
  XNOR U30356 ( .A(n25588), .B(n25587), .Z(n25590) );
  XNOR U30357 ( .A(n25584), .B(n25583), .Z(n25587) );
  XOR U30358 ( .A(n25586), .B(n25585), .Z(n25583) );
  XOR U30359 ( .A(y[239]), .B(x[239]), .Z(n25585) );
  XOR U30360 ( .A(y[238]), .B(x[238]), .Z(n25586) );
  XOR U30361 ( .A(y[237]), .B(x[237]), .Z(n25584) );
  XOR U30362 ( .A(n25578), .B(n25577), .Z(n25588) );
  XOR U30363 ( .A(n25580), .B(n25579), .Z(n25577) );
  XOR U30364 ( .A(y[236]), .B(x[236]), .Z(n25579) );
  XOR U30365 ( .A(y[235]), .B(x[235]), .Z(n25580) );
  XOR U30366 ( .A(y[234]), .B(x[234]), .Z(n25578) );
  XNOR U30367 ( .A(n25555), .B(n25554), .Z(n25572) );
  XNOR U30368 ( .A(n25569), .B(n25570), .Z(n25554) );
  XOR U30369 ( .A(n25566), .B(n25565), .Z(n25570) );
  XOR U30370 ( .A(y[231]), .B(x[231]), .Z(n25565) );
  XOR U30371 ( .A(n25568), .B(n25567), .Z(n25566) );
  XOR U30372 ( .A(y[233]), .B(x[233]), .Z(n25567) );
  XOR U30373 ( .A(y[232]), .B(x[232]), .Z(n25568) );
  XOR U30374 ( .A(n25560), .B(n25559), .Z(n25569) );
  XOR U30375 ( .A(n25562), .B(n25561), .Z(n25559) );
  XOR U30376 ( .A(y[230]), .B(x[230]), .Z(n25561) );
  XOR U30377 ( .A(y[229]), .B(x[229]), .Z(n25562) );
  XOR U30378 ( .A(y[228]), .B(x[228]), .Z(n25560) );
  XNOR U30379 ( .A(n25553), .B(n25552), .Z(n25555) );
  XNOR U30380 ( .A(n25549), .B(n25548), .Z(n25552) );
  XOR U30381 ( .A(n25551), .B(n25550), .Z(n25548) );
  XOR U30382 ( .A(y[227]), .B(x[227]), .Z(n25550) );
  XOR U30383 ( .A(y[226]), .B(x[226]), .Z(n25551) );
  XOR U30384 ( .A(y[225]), .B(x[225]), .Z(n25549) );
  XOR U30385 ( .A(n25543), .B(n25542), .Z(n25553) );
  XOR U30386 ( .A(n25545), .B(n25544), .Z(n25542) );
  XOR U30387 ( .A(y[224]), .B(x[224]), .Z(n25544) );
  XOR U30388 ( .A(y[223]), .B(x[223]), .Z(n25545) );
  XOR U30389 ( .A(y[222]), .B(x[222]), .Z(n25543) );
  NAND U30390 ( .A(n25606), .B(n25607), .Z(N28041) );
  NAND U30391 ( .A(n25608), .B(n25609), .Z(n25607) );
  NANDN U30392 ( .A(n25610), .B(n25611), .Z(n25609) );
  NANDN U30393 ( .A(n25611), .B(n25610), .Z(n25606) );
  XOR U30394 ( .A(n25610), .B(n25612), .Z(N28040) );
  XNOR U30395 ( .A(n25608), .B(n25611), .Z(n25612) );
  NAND U30396 ( .A(n25613), .B(n25614), .Z(n25611) );
  NAND U30397 ( .A(n25615), .B(n25616), .Z(n25614) );
  NANDN U30398 ( .A(n25617), .B(n25618), .Z(n25616) );
  NANDN U30399 ( .A(n25618), .B(n25617), .Z(n25613) );
  AND U30400 ( .A(n25619), .B(n25620), .Z(n25608) );
  NAND U30401 ( .A(n25621), .B(n25622), .Z(n25620) );
  OR U30402 ( .A(n25623), .B(n25624), .Z(n25622) );
  NAND U30403 ( .A(n25624), .B(n25623), .Z(n25619) );
  IV U30404 ( .A(n25625), .Z(n25624) );
  AND U30405 ( .A(n25626), .B(n25627), .Z(n25610) );
  NAND U30406 ( .A(n25628), .B(n25629), .Z(n25627) );
  NANDN U30407 ( .A(n25630), .B(n25631), .Z(n25629) );
  NANDN U30408 ( .A(n25631), .B(n25630), .Z(n25626) );
  XOR U30409 ( .A(n25623), .B(n25632), .Z(N28039) );
  XOR U30410 ( .A(n25621), .B(n25625), .Z(n25632) );
  XNOR U30411 ( .A(n25618), .B(n25633), .Z(n25625) );
  XNOR U30412 ( .A(n25615), .B(n25617), .Z(n25633) );
  AND U30413 ( .A(n25634), .B(n25635), .Z(n25617) );
  NANDN U30414 ( .A(n25636), .B(n25637), .Z(n25635) );
  NANDN U30415 ( .A(n25638), .B(n25639), .Z(n25637) );
  IV U30416 ( .A(n25640), .Z(n25639) );
  NAND U30417 ( .A(n25640), .B(n25638), .Z(n25634) );
  AND U30418 ( .A(n25641), .B(n25642), .Z(n25615) );
  NAND U30419 ( .A(n25643), .B(n25644), .Z(n25642) );
  OR U30420 ( .A(n25645), .B(n25646), .Z(n25644) );
  NAND U30421 ( .A(n25646), .B(n25645), .Z(n25641) );
  IV U30422 ( .A(n25647), .Z(n25646) );
  NAND U30423 ( .A(n25648), .B(n25649), .Z(n25618) );
  NANDN U30424 ( .A(n25650), .B(n25651), .Z(n25649) );
  NAND U30425 ( .A(n25652), .B(n25653), .Z(n25651) );
  OR U30426 ( .A(n25653), .B(n25652), .Z(n25648) );
  IV U30427 ( .A(n25654), .Z(n25652) );
  AND U30428 ( .A(n25655), .B(n25656), .Z(n25621) );
  NAND U30429 ( .A(n25657), .B(n25658), .Z(n25656) );
  NANDN U30430 ( .A(n25659), .B(n25660), .Z(n25658) );
  NANDN U30431 ( .A(n25660), .B(n25659), .Z(n25655) );
  XOR U30432 ( .A(n25631), .B(n25661), .Z(n25623) );
  XNOR U30433 ( .A(n25628), .B(n25630), .Z(n25661) );
  AND U30434 ( .A(n25662), .B(n25663), .Z(n25630) );
  NANDN U30435 ( .A(n25664), .B(n25665), .Z(n25663) );
  NANDN U30436 ( .A(n25666), .B(n25667), .Z(n25665) );
  IV U30437 ( .A(n25668), .Z(n25667) );
  NAND U30438 ( .A(n25668), .B(n25666), .Z(n25662) );
  AND U30439 ( .A(n25669), .B(n25670), .Z(n25628) );
  NAND U30440 ( .A(n25671), .B(n25672), .Z(n25670) );
  OR U30441 ( .A(n25673), .B(n25674), .Z(n25672) );
  NAND U30442 ( .A(n25674), .B(n25673), .Z(n25669) );
  IV U30443 ( .A(n25675), .Z(n25674) );
  NAND U30444 ( .A(n25676), .B(n25677), .Z(n25631) );
  NANDN U30445 ( .A(n25678), .B(n25679), .Z(n25677) );
  NAND U30446 ( .A(n25680), .B(n25681), .Z(n25679) );
  OR U30447 ( .A(n25681), .B(n25680), .Z(n25676) );
  IV U30448 ( .A(n25682), .Z(n25680) );
  XOR U30449 ( .A(n25657), .B(n25683), .Z(N28038) );
  XNOR U30450 ( .A(n25660), .B(n25659), .Z(n25683) );
  XNOR U30451 ( .A(n25671), .B(n25684), .Z(n25659) );
  XOR U30452 ( .A(n25675), .B(n25673), .Z(n25684) );
  XOR U30453 ( .A(n25681), .B(n25685), .Z(n25673) );
  XOR U30454 ( .A(n25678), .B(n25682), .Z(n25685) );
  NAND U30455 ( .A(n25686), .B(n25687), .Z(n25682) );
  NAND U30456 ( .A(n25688), .B(n25689), .Z(n25687) );
  NAND U30457 ( .A(n25690), .B(n25691), .Z(n25686) );
  AND U30458 ( .A(n25692), .B(n25693), .Z(n25678) );
  NAND U30459 ( .A(n25694), .B(n25695), .Z(n25693) );
  NAND U30460 ( .A(n25696), .B(n25697), .Z(n25692) );
  NANDN U30461 ( .A(n25698), .B(n25699), .Z(n25681) );
  NANDN U30462 ( .A(n25700), .B(n25701), .Z(n25675) );
  XNOR U30463 ( .A(n25666), .B(n25702), .Z(n25671) );
  XOR U30464 ( .A(n25664), .B(n25668), .Z(n25702) );
  NAND U30465 ( .A(n25703), .B(n25704), .Z(n25668) );
  NAND U30466 ( .A(n25705), .B(n25706), .Z(n25704) );
  NAND U30467 ( .A(n25707), .B(n25708), .Z(n25703) );
  AND U30468 ( .A(n25709), .B(n25710), .Z(n25664) );
  NAND U30469 ( .A(n25711), .B(n25712), .Z(n25710) );
  NAND U30470 ( .A(n25713), .B(n25714), .Z(n25709) );
  AND U30471 ( .A(n25715), .B(n25716), .Z(n25666) );
  NAND U30472 ( .A(n25717), .B(n25718), .Z(n25660) );
  XNOR U30473 ( .A(n25643), .B(n25719), .Z(n25657) );
  XOR U30474 ( .A(n25647), .B(n25645), .Z(n25719) );
  XOR U30475 ( .A(n25653), .B(n25720), .Z(n25645) );
  XOR U30476 ( .A(n25650), .B(n25654), .Z(n25720) );
  NAND U30477 ( .A(n25721), .B(n25722), .Z(n25654) );
  NAND U30478 ( .A(n25723), .B(n25724), .Z(n25722) );
  NAND U30479 ( .A(n25725), .B(n25726), .Z(n25721) );
  AND U30480 ( .A(n25727), .B(n25728), .Z(n25650) );
  NAND U30481 ( .A(n25729), .B(n25730), .Z(n25728) );
  NAND U30482 ( .A(n25731), .B(n25732), .Z(n25727) );
  NANDN U30483 ( .A(n25733), .B(n25734), .Z(n25653) );
  NANDN U30484 ( .A(n25735), .B(n25736), .Z(n25647) );
  XNOR U30485 ( .A(n25638), .B(n25737), .Z(n25643) );
  XOR U30486 ( .A(n25636), .B(n25640), .Z(n25737) );
  NAND U30487 ( .A(n25738), .B(n25739), .Z(n25640) );
  NAND U30488 ( .A(n25740), .B(n25741), .Z(n25739) );
  NAND U30489 ( .A(n25742), .B(n25743), .Z(n25738) );
  AND U30490 ( .A(n25744), .B(n25745), .Z(n25636) );
  NAND U30491 ( .A(n25746), .B(n25747), .Z(n25745) );
  NAND U30492 ( .A(n25748), .B(n25749), .Z(n25744) );
  AND U30493 ( .A(n25750), .B(n25751), .Z(n25638) );
  XOR U30494 ( .A(n25718), .B(n25717), .Z(N28037) );
  XNOR U30495 ( .A(n25736), .B(n25735), .Z(n25717) );
  XNOR U30496 ( .A(n25750), .B(n25751), .Z(n25735) );
  XOR U30497 ( .A(n25747), .B(n25746), .Z(n25751) );
  XOR U30498 ( .A(y[219]), .B(x[219]), .Z(n25746) );
  XOR U30499 ( .A(n25749), .B(n25748), .Z(n25747) );
  XOR U30500 ( .A(y[221]), .B(x[221]), .Z(n25748) );
  XOR U30501 ( .A(y[220]), .B(x[220]), .Z(n25749) );
  XOR U30502 ( .A(n25741), .B(n25740), .Z(n25750) );
  XOR U30503 ( .A(n25743), .B(n25742), .Z(n25740) );
  XOR U30504 ( .A(y[218]), .B(x[218]), .Z(n25742) );
  XOR U30505 ( .A(y[217]), .B(x[217]), .Z(n25743) );
  XOR U30506 ( .A(y[216]), .B(x[216]), .Z(n25741) );
  XNOR U30507 ( .A(n25734), .B(n25733), .Z(n25736) );
  XNOR U30508 ( .A(n25730), .B(n25729), .Z(n25733) );
  XOR U30509 ( .A(n25732), .B(n25731), .Z(n25729) );
  XOR U30510 ( .A(y[215]), .B(x[215]), .Z(n25731) );
  XOR U30511 ( .A(y[214]), .B(x[214]), .Z(n25732) );
  XOR U30512 ( .A(y[213]), .B(x[213]), .Z(n25730) );
  XOR U30513 ( .A(n25724), .B(n25723), .Z(n25734) );
  XOR U30514 ( .A(n25726), .B(n25725), .Z(n25723) );
  XOR U30515 ( .A(y[212]), .B(x[212]), .Z(n25725) );
  XOR U30516 ( .A(y[211]), .B(x[211]), .Z(n25726) );
  XOR U30517 ( .A(y[210]), .B(x[210]), .Z(n25724) );
  XNOR U30518 ( .A(n25701), .B(n25700), .Z(n25718) );
  XNOR U30519 ( .A(n25715), .B(n25716), .Z(n25700) );
  XOR U30520 ( .A(n25712), .B(n25711), .Z(n25716) );
  XOR U30521 ( .A(y[207]), .B(x[207]), .Z(n25711) );
  XOR U30522 ( .A(n25714), .B(n25713), .Z(n25712) );
  XOR U30523 ( .A(y[209]), .B(x[209]), .Z(n25713) );
  XOR U30524 ( .A(y[208]), .B(x[208]), .Z(n25714) );
  XOR U30525 ( .A(n25706), .B(n25705), .Z(n25715) );
  XOR U30526 ( .A(n25708), .B(n25707), .Z(n25705) );
  XOR U30527 ( .A(y[206]), .B(x[206]), .Z(n25707) );
  XOR U30528 ( .A(y[205]), .B(x[205]), .Z(n25708) );
  XOR U30529 ( .A(y[204]), .B(x[204]), .Z(n25706) );
  XNOR U30530 ( .A(n25699), .B(n25698), .Z(n25701) );
  XNOR U30531 ( .A(n25695), .B(n25694), .Z(n25698) );
  XOR U30532 ( .A(n25697), .B(n25696), .Z(n25694) );
  XOR U30533 ( .A(y[203]), .B(x[203]), .Z(n25696) );
  XOR U30534 ( .A(y[202]), .B(x[202]), .Z(n25697) );
  XOR U30535 ( .A(y[201]), .B(x[201]), .Z(n25695) );
  XOR U30536 ( .A(n25689), .B(n25688), .Z(n25699) );
  XOR U30537 ( .A(n25691), .B(n25690), .Z(n25688) );
  XOR U30538 ( .A(y[200]), .B(x[200]), .Z(n25690) );
  XOR U30539 ( .A(y[199]), .B(x[199]), .Z(n25691) );
  XOR U30540 ( .A(y[198]), .B(x[198]), .Z(n25689) );
  NAND U30541 ( .A(n25752), .B(n25753), .Z(N28029) );
  NAND U30542 ( .A(n25754), .B(n25755), .Z(n25753) );
  NANDN U30543 ( .A(n25756), .B(n25757), .Z(n25755) );
  NANDN U30544 ( .A(n25757), .B(n25756), .Z(n25752) );
  XOR U30545 ( .A(n25756), .B(n25758), .Z(N28028) );
  XNOR U30546 ( .A(n25754), .B(n25757), .Z(n25758) );
  NAND U30547 ( .A(n25759), .B(n25760), .Z(n25757) );
  NAND U30548 ( .A(n25761), .B(n25762), .Z(n25760) );
  NANDN U30549 ( .A(n25763), .B(n25764), .Z(n25762) );
  NANDN U30550 ( .A(n25764), .B(n25763), .Z(n25759) );
  AND U30551 ( .A(n25765), .B(n25766), .Z(n25754) );
  NAND U30552 ( .A(n25767), .B(n25768), .Z(n25766) );
  OR U30553 ( .A(n25769), .B(n25770), .Z(n25768) );
  NAND U30554 ( .A(n25770), .B(n25769), .Z(n25765) );
  IV U30555 ( .A(n25771), .Z(n25770) );
  AND U30556 ( .A(n25772), .B(n25773), .Z(n25756) );
  NAND U30557 ( .A(n25774), .B(n25775), .Z(n25773) );
  NANDN U30558 ( .A(n25776), .B(n25777), .Z(n25775) );
  NANDN U30559 ( .A(n25777), .B(n25776), .Z(n25772) );
  XOR U30560 ( .A(n25769), .B(n25778), .Z(N28027) );
  XOR U30561 ( .A(n25767), .B(n25771), .Z(n25778) );
  XNOR U30562 ( .A(n25764), .B(n25779), .Z(n25771) );
  XNOR U30563 ( .A(n25761), .B(n25763), .Z(n25779) );
  AND U30564 ( .A(n25780), .B(n25781), .Z(n25763) );
  NANDN U30565 ( .A(n25782), .B(n25783), .Z(n25781) );
  NANDN U30566 ( .A(n25784), .B(n25785), .Z(n25783) );
  IV U30567 ( .A(n25786), .Z(n25785) );
  NAND U30568 ( .A(n25786), .B(n25784), .Z(n25780) );
  AND U30569 ( .A(n25787), .B(n25788), .Z(n25761) );
  NAND U30570 ( .A(n25789), .B(n25790), .Z(n25788) );
  OR U30571 ( .A(n25791), .B(n25792), .Z(n25790) );
  NAND U30572 ( .A(n25792), .B(n25791), .Z(n25787) );
  IV U30573 ( .A(n25793), .Z(n25792) );
  NAND U30574 ( .A(n25794), .B(n25795), .Z(n25764) );
  NANDN U30575 ( .A(n25796), .B(n25797), .Z(n25795) );
  NAND U30576 ( .A(n25798), .B(n25799), .Z(n25797) );
  OR U30577 ( .A(n25799), .B(n25798), .Z(n25794) );
  IV U30578 ( .A(n25800), .Z(n25798) );
  AND U30579 ( .A(n25801), .B(n25802), .Z(n25767) );
  NAND U30580 ( .A(n25803), .B(n25804), .Z(n25802) );
  NANDN U30581 ( .A(n25805), .B(n25806), .Z(n25804) );
  NANDN U30582 ( .A(n25806), .B(n25805), .Z(n25801) );
  XOR U30583 ( .A(n25777), .B(n25807), .Z(n25769) );
  XNOR U30584 ( .A(n25774), .B(n25776), .Z(n25807) );
  AND U30585 ( .A(n25808), .B(n25809), .Z(n25776) );
  NANDN U30586 ( .A(n25810), .B(n25811), .Z(n25809) );
  NANDN U30587 ( .A(n25812), .B(n25813), .Z(n25811) );
  IV U30588 ( .A(n25814), .Z(n25813) );
  NAND U30589 ( .A(n25814), .B(n25812), .Z(n25808) );
  AND U30590 ( .A(n25815), .B(n25816), .Z(n25774) );
  NAND U30591 ( .A(n25817), .B(n25818), .Z(n25816) );
  OR U30592 ( .A(n25819), .B(n25820), .Z(n25818) );
  NAND U30593 ( .A(n25820), .B(n25819), .Z(n25815) );
  IV U30594 ( .A(n25821), .Z(n25820) );
  NAND U30595 ( .A(n25822), .B(n25823), .Z(n25777) );
  NANDN U30596 ( .A(n25824), .B(n25825), .Z(n25823) );
  NAND U30597 ( .A(n25826), .B(n25827), .Z(n25825) );
  OR U30598 ( .A(n25827), .B(n25826), .Z(n25822) );
  IV U30599 ( .A(n25828), .Z(n25826) );
  XOR U30600 ( .A(n25803), .B(n25829), .Z(N28026) );
  XNOR U30601 ( .A(n25806), .B(n25805), .Z(n25829) );
  XNOR U30602 ( .A(n25817), .B(n25830), .Z(n25805) );
  XOR U30603 ( .A(n25821), .B(n25819), .Z(n25830) );
  XOR U30604 ( .A(n25827), .B(n25831), .Z(n25819) );
  XOR U30605 ( .A(n25824), .B(n25828), .Z(n25831) );
  NAND U30606 ( .A(n25832), .B(n25833), .Z(n25828) );
  NAND U30607 ( .A(n25834), .B(n25835), .Z(n25833) );
  NAND U30608 ( .A(n25836), .B(n25837), .Z(n25832) );
  AND U30609 ( .A(n25838), .B(n25839), .Z(n25824) );
  NAND U30610 ( .A(n25840), .B(n25841), .Z(n25839) );
  NAND U30611 ( .A(n25842), .B(n25843), .Z(n25838) );
  NANDN U30612 ( .A(n25844), .B(n25845), .Z(n25827) );
  NANDN U30613 ( .A(n25846), .B(n25847), .Z(n25821) );
  XNOR U30614 ( .A(n25812), .B(n25848), .Z(n25817) );
  XOR U30615 ( .A(n25810), .B(n25814), .Z(n25848) );
  NAND U30616 ( .A(n25849), .B(n25850), .Z(n25814) );
  NAND U30617 ( .A(n25851), .B(n25852), .Z(n25850) );
  NAND U30618 ( .A(n25853), .B(n25854), .Z(n25849) );
  AND U30619 ( .A(n25855), .B(n25856), .Z(n25810) );
  NAND U30620 ( .A(n25857), .B(n25858), .Z(n25856) );
  NAND U30621 ( .A(n25859), .B(n25860), .Z(n25855) );
  AND U30622 ( .A(n25861), .B(n25862), .Z(n25812) );
  NAND U30623 ( .A(n25863), .B(n25864), .Z(n25806) );
  XNOR U30624 ( .A(n25789), .B(n25865), .Z(n25803) );
  XOR U30625 ( .A(n25793), .B(n25791), .Z(n25865) );
  XOR U30626 ( .A(n25799), .B(n25866), .Z(n25791) );
  XOR U30627 ( .A(n25796), .B(n25800), .Z(n25866) );
  NAND U30628 ( .A(n25867), .B(n25868), .Z(n25800) );
  NAND U30629 ( .A(n25869), .B(n25870), .Z(n25868) );
  NAND U30630 ( .A(n25871), .B(n25872), .Z(n25867) );
  AND U30631 ( .A(n25873), .B(n25874), .Z(n25796) );
  NAND U30632 ( .A(n25875), .B(n25876), .Z(n25874) );
  NAND U30633 ( .A(n25877), .B(n25878), .Z(n25873) );
  NANDN U30634 ( .A(n25879), .B(n25880), .Z(n25799) );
  NANDN U30635 ( .A(n25881), .B(n25882), .Z(n25793) );
  XNOR U30636 ( .A(n25784), .B(n25883), .Z(n25789) );
  XOR U30637 ( .A(n25782), .B(n25786), .Z(n25883) );
  NAND U30638 ( .A(n25884), .B(n25885), .Z(n25786) );
  NAND U30639 ( .A(n25886), .B(n25887), .Z(n25885) );
  NAND U30640 ( .A(n25888), .B(n25889), .Z(n25884) );
  AND U30641 ( .A(n25890), .B(n25891), .Z(n25782) );
  NAND U30642 ( .A(n25892), .B(n25893), .Z(n25891) );
  NAND U30643 ( .A(n25894), .B(n25895), .Z(n25890) );
  AND U30644 ( .A(n25896), .B(n25897), .Z(n25784) );
  XOR U30645 ( .A(n25864), .B(n25863), .Z(N28025) );
  XNOR U30646 ( .A(n25882), .B(n25881), .Z(n25863) );
  XNOR U30647 ( .A(n25896), .B(n25897), .Z(n25881) );
  XOR U30648 ( .A(n25893), .B(n25892), .Z(n25897) );
  XOR U30649 ( .A(y[195]), .B(x[195]), .Z(n25892) );
  XOR U30650 ( .A(n25895), .B(n25894), .Z(n25893) );
  XOR U30651 ( .A(y[197]), .B(x[197]), .Z(n25894) );
  XOR U30652 ( .A(y[196]), .B(x[196]), .Z(n25895) );
  XOR U30653 ( .A(n25887), .B(n25886), .Z(n25896) );
  XOR U30654 ( .A(n25889), .B(n25888), .Z(n25886) );
  XOR U30655 ( .A(y[194]), .B(x[194]), .Z(n25888) );
  XOR U30656 ( .A(y[193]), .B(x[193]), .Z(n25889) );
  XOR U30657 ( .A(y[192]), .B(x[192]), .Z(n25887) );
  XNOR U30658 ( .A(n25880), .B(n25879), .Z(n25882) );
  XNOR U30659 ( .A(n25876), .B(n25875), .Z(n25879) );
  XOR U30660 ( .A(n25878), .B(n25877), .Z(n25875) );
  XOR U30661 ( .A(y[191]), .B(x[191]), .Z(n25877) );
  XOR U30662 ( .A(y[190]), .B(x[190]), .Z(n25878) );
  XOR U30663 ( .A(y[189]), .B(x[189]), .Z(n25876) );
  XOR U30664 ( .A(n25870), .B(n25869), .Z(n25880) );
  XOR U30665 ( .A(n25872), .B(n25871), .Z(n25869) );
  XOR U30666 ( .A(y[188]), .B(x[188]), .Z(n25871) );
  XOR U30667 ( .A(y[187]), .B(x[187]), .Z(n25872) );
  XOR U30668 ( .A(y[186]), .B(x[186]), .Z(n25870) );
  XNOR U30669 ( .A(n25847), .B(n25846), .Z(n25864) );
  XNOR U30670 ( .A(n25861), .B(n25862), .Z(n25846) );
  XOR U30671 ( .A(n25858), .B(n25857), .Z(n25862) );
  XOR U30672 ( .A(y[183]), .B(x[183]), .Z(n25857) );
  XOR U30673 ( .A(n25860), .B(n25859), .Z(n25858) );
  XOR U30674 ( .A(y[185]), .B(x[185]), .Z(n25859) );
  XOR U30675 ( .A(y[184]), .B(x[184]), .Z(n25860) );
  XOR U30676 ( .A(n25852), .B(n25851), .Z(n25861) );
  XOR U30677 ( .A(n25854), .B(n25853), .Z(n25851) );
  XOR U30678 ( .A(y[182]), .B(x[182]), .Z(n25853) );
  XOR U30679 ( .A(y[181]), .B(x[181]), .Z(n25854) );
  XOR U30680 ( .A(y[180]), .B(x[180]), .Z(n25852) );
  XNOR U30681 ( .A(n25845), .B(n25844), .Z(n25847) );
  XNOR U30682 ( .A(n25841), .B(n25840), .Z(n25844) );
  XOR U30683 ( .A(n25843), .B(n25842), .Z(n25840) );
  XOR U30684 ( .A(y[179]), .B(x[179]), .Z(n25842) );
  XOR U30685 ( .A(y[178]), .B(x[178]), .Z(n25843) );
  XOR U30686 ( .A(y[177]), .B(x[177]), .Z(n25841) );
  XOR U30687 ( .A(n25835), .B(n25834), .Z(n25845) );
  XOR U30688 ( .A(n25837), .B(n25836), .Z(n25834) );
  XOR U30689 ( .A(y[176]), .B(x[176]), .Z(n25836) );
  XOR U30690 ( .A(y[175]), .B(x[175]), .Z(n25837) );
  XOR U30691 ( .A(y[174]), .B(x[174]), .Z(n25835) );
  NAND U30692 ( .A(n25898), .B(n25899), .Z(N28017) );
  NAND U30693 ( .A(n25900), .B(n25901), .Z(n25899) );
  NANDN U30694 ( .A(n25902), .B(n25903), .Z(n25901) );
  NANDN U30695 ( .A(n25903), .B(n25902), .Z(n25898) );
  XOR U30696 ( .A(n25902), .B(n25904), .Z(N28016) );
  XNOR U30697 ( .A(n25900), .B(n25903), .Z(n25904) );
  NAND U30698 ( .A(n25905), .B(n25906), .Z(n25903) );
  NAND U30699 ( .A(n25907), .B(n25908), .Z(n25906) );
  NANDN U30700 ( .A(n25909), .B(n25910), .Z(n25908) );
  NANDN U30701 ( .A(n25910), .B(n25909), .Z(n25905) );
  AND U30702 ( .A(n25911), .B(n25912), .Z(n25900) );
  NAND U30703 ( .A(n25913), .B(n25914), .Z(n25912) );
  OR U30704 ( .A(n25915), .B(n25916), .Z(n25914) );
  NAND U30705 ( .A(n25916), .B(n25915), .Z(n25911) );
  IV U30706 ( .A(n25917), .Z(n25916) );
  AND U30707 ( .A(n25918), .B(n25919), .Z(n25902) );
  NAND U30708 ( .A(n25920), .B(n25921), .Z(n25919) );
  NANDN U30709 ( .A(n25922), .B(n25923), .Z(n25921) );
  NANDN U30710 ( .A(n25923), .B(n25922), .Z(n25918) );
  XOR U30711 ( .A(n25915), .B(n25924), .Z(N28015) );
  XOR U30712 ( .A(n25913), .B(n25917), .Z(n25924) );
  XNOR U30713 ( .A(n25910), .B(n25925), .Z(n25917) );
  XNOR U30714 ( .A(n25907), .B(n25909), .Z(n25925) );
  AND U30715 ( .A(n25926), .B(n25927), .Z(n25909) );
  NANDN U30716 ( .A(n25928), .B(n25929), .Z(n25927) );
  NANDN U30717 ( .A(n25930), .B(n25931), .Z(n25929) );
  IV U30718 ( .A(n25932), .Z(n25931) );
  NAND U30719 ( .A(n25932), .B(n25930), .Z(n25926) );
  AND U30720 ( .A(n25933), .B(n25934), .Z(n25907) );
  NAND U30721 ( .A(n25935), .B(n25936), .Z(n25934) );
  OR U30722 ( .A(n25937), .B(n25938), .Z(n25936) );
  NAND U30723 ( .A(n25938), .B(n25937), .Z(n25933) );
  IV U30724 ( .A(n25939), .Z(n25938) );
  NAND U30725 ( .A(n25940), .B(n25941), .Z(n25910) );
  NANDN U30726 ( .A(n25942), .B(n25943), .Z(n25941) );
  NAND U30727 ( .A(n25944), .B(n25945), .Z(n25943) );
  OR U30728 ( .A(n25945), .B(n25944), .Z(n25940) );
  IV U30729 ( .A(n25946), .Z(n25944) );
  AND U30730 ( .A(n25947), .B(n25948), .Z(n25913) );
  NAND U30731 ( .A(n25949), .B(n25950), .Z(n25948) );
  NANDN U30732 ( .A(n25951), .B(n25952), .Z(n25950) );
  NANDN U30733 ( .A(n25952), .B(n25951), .Z(n25947) );
  XOR U30734 ( .A(n25923), .B(n25953), .Z(n25915) );
  XNOR U30735 ( .A(n25920), .B(n25922), .Z(n25953) );
  AND U30736 ( .A(n25954), .B(n25955), .Z(n25922) );
  NANDN U30737 ( .A(n25956), .B(n25957), .Z(n25955) );
  NANDN U30738 ( .A(n25958), .B(n25959), .Z(n25957) );
  IV U30739 ( .A(n25960), .Z(n25959) );
  NAND U30740 ( .A(n25960), .B(n25958), .Z(n25954) );
  AND U30741 ( .A(n25961), .B(n25962), .Z(n25920) );
  NAND U30742 ( .A(n25963), .B(n25964), .Z(n25962) );
  OR U30743 ( .A(n25965), .B(n25966), .Z(n25964) );
  NAND U30744 ( .A(n25966), .B(n25965), .Z(n25961) );
  IV U30745 ( .A(n25967), .Z(n25966) );
  NAND U30746 ( .A(n25968), .B(n25969), .Z(n25923) );
  NANDN U30747 ( .A(n25970), .B(n25971), .Z(n25969) );
  NAND U30748 ( .A(n25972), .B(n25973), .Z(n25971) );
  OR U30749 ( .A(n25973), .B(n25972), .Z(n25968) );
  IV U30750 ( .A(n25974), .Z(n25972) );
  XOR U30751 ( .A(n25949), .B(n25975), .Z(N28014) );
  XNOR U30752 ( .A(n25952), .B(n25951), .Z(n25975) );
  XNOR U30753 ( .A(n25963), .B(n25976), .Z(n25951) );
  XOR U30754 ( .A(n25967), .B(n25965), .Z(n25976) );
  XOR U30755 ( .A(n25973), .B(n25977), .Z(n25965) );
  XOR U30756 ( .A(n25970), .B(n25974), .Z(n25977) );
  NAND U30757 ( .A(n25978), .B(n25979), .Z(n25974) );
  NAND U30758 ( .A(n25980), .B(n25981), .Z(n25979) );
  NAND U30759 ( .A(n25982), .B(n25983), .Z(n25978) );
  AND U30760 ( .A(n25984), .B(n25985), .Z(n25970) );
  NAND U30761 ( .A(n25986), .B(n25987), .Z(n25985) );
  NAND U30762 ( .A(n25988), .B(n25989), .Z(n25984) );
  NANDN U30763 ( .A(n25990), .B(n25991), .Z(n25973) );
  NANDN U30764 ( .A(n25992), .B(n25993), .Z(n25967) );
  XNOR U30765 ( .A(n25958), .B(n25994), .Z(n25963) );
  XOR U30766 ( .A(n25956), .B(n25960), .Z(n25994) );
  NAND U30767 ( .A(n25995), .B(n25996), .Z(n25960) );
  NAND U30768 ( .A(n25997), .B(n25998), .Z(n25996) );
  NAND U30769 ( .A(n25999), .B(n26000), .Z(n25995) );
  AND U30770 ( .A(n26001), .B(n26002), .Z(n25956) );
  NAND U30771 ( .A(n26003), .B(n26004), .Z(n26002) );
  NAND U30772 ( .A(n26005), .B(n26006), .Z(n26001) );
  AND U30773 ( .A(n26007), .B(n26008), .Z(n25958) );
  NAND U30774 ( .A(n26009), .B(n26010), .Z(n25952) );
  XNOR U30775 ( .A(n25935), .B(n26011), .Z(n25949) );
  XOR U30776 ( .A(n25939), .B(n25937), .Z(n26011) );
  XOR U30777 ( .A(n25945), .B(n26012), .Z(n25937) );
  XOR U30778 ( .A(n25942), .B(n25946), .Z(n26012) );
  NAND U30779 ( .A(n26013), .B(n26014), .Z(n25946) );
  NAND U30780 ( .A(n26015), .B(n26016), .Z(n26014) );
  NAND U30781 ( .A(n26017), .B(n26018), .Z(n26013) );
  AND U30782 ( .A(n26019), .B(n26020), .Z(n25942) );
  NAND U30783 ( .A(n26021), .B(n26022), .Z(n26020) );
  NAND U30784 ( .A(n26023), .B(n26024), .Z(n26019) );
  NANDN U30785 ( .A(n26025), .B(n26026), .Z(n25945) );
  NANDN U30786 ( .A(n26027), .B(n26028), .Z(n25939) );
  XNOR U30787 ( .A(n25930), .B(n26029), .Z(n25935) );
  XOR U30788 ( .A(n25928), .B(n25932), .Z(n26029) );
  NAND U30789 ( .A(n26030), .B(n26031), .Z(n25932) );
  NAND U30790 ( .A(n26032), .B(n26033), .Z(n26031) );
  NAND U30791 ( .A(n26034), .B(n26035), .Z(n26030) );
  AND U30792 ( .A(n26036), .B(n26037), .Z(n25928) );
  NAND U30793 ( .A(n26038), .B(n26039), .Z(n26037) );
  NAND U30794 ( .A(n26040), .B(n26041), .Z(n26036) );
  AND U30795 ( .A(n26042), .B(n26043), .Z(n25930) );
  XOR U30796 ( .A(n26010), .B(n26009), .Z(N28013) );
  XNOR U30797 ( .A(n26028), .B(n26027), .Z(n26009) );
  XNOR U30798 ( .A(n26042), .B(n26043), .Z(n26027) );
  XOR U30799 ( .A(n26039), .B(n26038), .Z(n26043) );
  XOR U30800 ( .A(y[171]), .B(x[171]), .Z(n26038) );
  XOR U30801 ( .A(n26041), .B(n26040), .Z(n26039) );
  XOR U30802 ( .A(y[173]), .B(x[173]), .Z(n26040) );
  XOR U30803 ( .A(y[172]), .B(x[172]), .Z(n26041) );
  XOR U30804 ( .A(n26033), .B(n26032), .Z(n26042) );
  XOR U30805 ( .A(n26035), .B(n26034), .Z(n26032) );
  XOR U30806 ( .A(y[170]), .B(x[170]), .Z(n26034) );
  XOR U30807 ( .A(y[169]), .B(x[169]), .Z(n26035) );
  XOR U30808 ( .A(y[168]), .B(x[168]), .Z(n26033) );
  XNOR U30809 ( .A(n26026), .B(n26025), .Z(n26028) );
  XNOR U30810 ( .A(n26022), .B(n26021), .Z(n26025) );
  XOR U30811 ( .A(n26024), .B(n26023), .Z(n26021) );
  XOR U30812 ( .A(y[167]), .B(x[167]), .Z(n26023) );
  XOR U30813 ( .A(y[166]), .B(x[166]), .Z(n26024) );
  XOR U30814 ( .A(y[165]), .B(x[165]), .Z(n26022) );
  XOR U30815 ( .A(n26016), .B(n26015), .Z(n26026) );
  XOR U30816 ( .A(n26018), .B(n26017), .Z(n26015) );
  XOR U30817 ( .A(y[164]), .B(x[164]), .Z(n26017) );
  XOR U30818 ( .A(y[163]), .B(x[163]), .Z(n26018) );
  XOR U30819 ( .A(y[162]), .B(x[162]), .Z(n26016) );
  XNOR U30820 ( .A(n25993), .B(n25992), .Z(n26010) );
  XNOR U30821 ( .A(n26007), .B(n26008), .Z(n25992) );
  XOR U30822 ( .A(n26004), .B(n26003), .Z(n26008) );
  XOR U30823 ( .A(y[159]), .B(x[159]), .Z(n26003) );
  XOR U30824 ( .A(n26006), .B(n26005), .Z(n26004) );
  XOR U30825 ( .A(y[161]), .B(x[161]), .Z(n26005) );
  XOR U30826 ( .A(y[160]), .B(x[160]), .Z(n26006) );
  XOR U30827 ( .A(n25998), .B(n25997), .Z(n26007) );
  XOR U30828 ( .A(n26000), .B(n25999), .Z(n25997) );
  XOR U30829 ( .A(y[158]), .B(x[158]), .Z(n25999) );
  XOR U30830 ( .A(y[157]), .B(x[157]), .Z(n26000) );
  XOR U30831 ( .A(y[156]), .B(x[156]), .Z(n25998) );
  XNOR U30832 ( .A(n25991), .B(n25990), .Z(n25993) );
  XNOR U30833 ( .A(n25987), .B(n25986), .Z(n25990) );
  XOR U30834 ( .A(n25989), .B(n25988), .Z(n25986) );
  XOR U30835 ( .A(y[155]), .B(x[155]), .Z(n25988) );
  XOR U30836 ( .A(y[154]), .B(x[154]), .Z(n25989) );
  XOR U30837 ( .A(y[153]), .B(x[153]), .Z(n25987) );
  XOR U30838 ( .A(n25981), .B(n25980), .Z(n25991) );
  XOR U30839 ( .A(n25983), .B(n25982), .Z(n25980) );
  XOR U30840 ( .A(y[152]), .B(x[152]), .Z(n25982) );
  XOR U30841 ( .A(y[151]), .B(x[151]), .Z(n25983) );
  XOR U30842 ( .A(y[150]), .B(x[150]), .Z(n25981) );
  NAND U30843 ( .A(n26044), .B(n26045), .Z(N28005) );
  NAND U30844 ( .A(n26046), .B(n26047), .Z(n26045) );
  NANDN U30845 ( .A(n26048), .B(n26049), .Z(n26047) );
  NANDN U30846 ( .A(n26049), .B(n26048), .Z(n26044) );
  XOR U30847 ( .A(n26048), .B(n26050), .Z(N28004) );
  XNOR U30848 ( .A(n26046), .B(n26049), .Z(n26050) );
  NAND U30849 ( .A(n26051), .B(n26052), .Z(n26049) );
  NAND U30850 ( .A(n26053), .B(n26054), .Z(n26052) );
  NANDN U30851 ( .A(n26055), .B(n26056), .Z(n26054) );
  NANDN U30852 ( .A(n26056), .B(n26055), .Z(n26051) );
  AND U30853 ( .A(n26057), .B(n26058), .Z(n26046) );
  NAND U30854 ( .A(n26059), .B(n26060), .Z(n26058) );
  OR U30855 ( .A(n26061), .B(n26062), .Z(n26060) );
  NAND U30856 ( .A(n26062), .B(n26061), .Z(n26057) );
  IV U30857 ( .A(n26063), .Z(n26062) );
  AND U30858 ( .A(n26064), .B(n26065), .Z(n26048) );
  NAND U30859 ( .A(n26066), .B(n26067), .Z(n26065) );
  NANDN U30860 ( .A(n26068), .B(n26069), .Z(n26067) );
  NANDN U30861 ( .A(n26069), .B(n26068), .Z(n26064) );
  XOR U30862 ( .A(n26061), .B(n26070), .Z(N28003) );
  XOR U30863 ( .A(n26059), .B(n26063), .Z(n26070) );
  XNOR U30864 ( .A(n26056), .B(n26071), .Z(n26063) );
  XNOR U30865 ( .A(n26053), .B(n26055), .Z(n26071) );
  AND U30866 ( .A(n26072), .B(n26073), .Z(n26055) );
  NANDN U30867 ( .A(n26074), .B(n26075), .Z(n26073) );
  NANDN U30868 ( .A(n26076), .B(n26077), .Z(n26075) );
  IV U30869 ( .A(n26078), .Z(n26077) );
  NAND U30870 ( .A(n26078), .B(n26076), .Z(n26072) );
  AND U30871 ( .A(n26079), .B(n26080), .Z(n26053) );
  NAND U30872 ( .A(n26081), .B(n26082), .Z(n26080) );
  OR U30873 ( .A(n26083), .B(n26084), .Z(n26082) );
  NAND U30874 ( .A(n26084), .B(n26083), .Z(n26079) );
  IV U30875 ( .A(n26085), .Z(n26084) );
  NAND U30876 ( .A(n26086), .B(n26087), .Z(n26056) );
  NANDN U30877 ( .A(n26088), .B(n26089), .Z(n26087) );
  NAND U30878 ( .A(n26090), .B(n26091), .Z(n26089) );
  OR U30879 ( .A(n26091), .B(n26090), .Z(n26086) );
  IV U30880 ( .A(n26092), .Z(n26090) );
  AND U30881 ( .A(n26093), .B(n26094), .Z(n26059) );
  NAND U30882 ( .A(n26095), .B(n26096), .Z(n26094) );
  NANDN U30883 ( .A(n26097), .B(n26098), .Z(n26096) );
  NANDN U30884 ( .A(n26098), .B(n26097), .Z(n26093) );
  XOR U30885 ( .A(n26069), .B(n26099), .Z(n26061) );
  XNOR U30886 ( .A(n26066), .B(n26068), .Z(n26099) );
  AND U30887 ( .A(n26100), .B(n26101), .Z(n26068) );
  NANDN U30888 ( .A(n26102), .B(n26103), .Z(n26101) );
  NANDN U30889 ( .A(n26104), .B(n26105), .Z(n26103) );
  IV U30890 ( .A(n26106), .Z(n26105) );
  NAND U30891 ( .A(n26106), .B(n26104), .Z(n26100) );
  AND U30892 ( .A(n26107), .B(n26108), .Z(n26066) );
  NAND U30893 ( .A(n26109), .B(n26110), .Z(n26108) );
  OR U30894 ( .A(n26111), .B(n26112), .Z(n26110) );
  NAND U30895 ( .A(n26112), .B(n26111), .Z(n26107) );
  IV U30896 ( .A(n26113), .Z(n26112) );
  NAND U30897 ( .A(n26114), .B(n26115), .Z(n26069) );
  NANDN U30898 ( .A(n26116), .B(n26117), .Z(n26115) );
  NAND U30899 ( .A(n26118), .B(n26119), .Z(n26117) );
  OR U30900 ( .A(n26119), .B(n26118), .Z(n26114) );
  IV U30901 ( .A(n26120), .Z(n26118) );
  XOR U30902 ( .A(n26095), .B(n26121), .Z(N28002) );
  XNOR U30903 ( .A(n26098), .B(n26097), .Z(n26121) );
  XNOR U30904 ( .A(n26109), .B(n26122), .Z(n26097) );
  XOR U30905 ( .A(n26113), .B(n26111), .Z(n26122) );
  XOR U30906 ( .A(n26119), .B(n26123), .Z(n26111) );
  XOR U30907 ( .A(n26116), .B(n26120), .Z(n26123) );
  NAND U30908 ( .A(n26124), .B(n26125), .Z(n26120) );
  NAND U30909 ( .A(n26126), .B(n26127), .Z(n26125) );
  NAND U30910 ( .A(n26128), .B(n26129), .Z(n26124) );
  AND U30911 ( .A(n26130), .B(n26131), .Z(n26116) );
  NAND U30912 ( .A(n26132), .B(n26133), .Z(n26131) );
  NAND U30913 ( .A(n26134), .B(n26135), .Z(n26130) );
  NANDN U30914 ( .A(n26136), .B(n26137), .Z(n26119) );
  NANDN U30915 ( .A(n26138), .B(n26139), .Z(n26113) );
  XNOR U30916 ( .A(n26104), .B(n26140), .Z(n26109) );
  XOR U30917 ( .A(n26102), .B(n26106), .Z(n26140) );
  NAND U30918 ( .A(n26141), .B(n26142), .Z(n26106) );
  NAND U30919 ( .A(n26143), .B(n26144), .Z(n26142) );
  NAND U30920 ( .A(n26145), .B(n26146), .Z(n26141) );
  AND U30921 ( .A(n26147), .B(n26148), .Z(n26102) );
  NAND U30922 ( .A(n26149), .B(n26150), .Z(n26148) );
  NAND U30923 ( .A(n26151), .B(n26152), .Z(n26147) );
  AND U30924 ( .A(n26153), .B(n26154), .Z(n26104) );
  NAND U30925 ( .A(n26155), .B(n26156), .Z(n26098) );
  XNOR U30926 ( .A(n26081), .B(n26157), .Z(n26095) );
  XOR U30927 ( .A(n26085), .B(n26083), .Z(n26157) );
  XOR U30928 ( .A(n26091), .B(n26158), .Z(n26083) );
  XOR U30929 ( .A(n26088), .B(n26092), .Z(n26158) );
  NAND U30930 ( .A(n26159), .B(n26160), .Z(n26092) );
  NAND U30931 ( .A(n26161), .B(n26162), .Z(n26160) );
  NAND U30932 ( .A(n26163), .B(n26164), .Z(n26159) );
  AND U30933 ( .A(n26165), .B(n26166), .Z(n26088) );
  NAND U30934 ( .A(n26167), .B(n26168), .Z(n26166) );
  NAND U30935 ( .A(n26169), .B(n26170), .Z(n26165) );
  NANDN U30936 ( .A(n26171), .B(n26172), .Z(n26091) );
  NANDN U30937 ( .A(n26173), .B(n26174), .Z(n26085) );
  XNOR U30938 ( .A(n26076), .B(n26175), .Z(n26081) );
  XOR U30939 ( .A(n26074), .B(n26078), .Z(n26175) );
  NAND U30940 ( .A(n26176), .B(n26177), .Z(n26078) );
  NAND U30941 ( .A(n26178), .B(n26179), .Z(n26177) );
  NAND U30942 ( .A(n26180), .B(n26181), .Z(n26176) );
  AND U30943 ( .A(n26182), .B(n26183), .Z(n26074) );
  NAND U30944 ( .A(n26184), .B(n26185), .Z(n26183) );
  NAND U30945 ( .A(n26186), .B(n26187), .Z(n26182) );
  AND U30946 ( .A(n26188), .B(n26189), .Z(n26076) );
  XOR U30947 ( .A(n26156), .B(n26155), .Z(N28001) );
  XNOR U30948 ( .A(n26174), .B(n26173), .Z(n26155) );
  XNOR U30949 ( .A(n26188), .B(n26189), .Z(n26173) );
  XOR U30950 ( .A(n26185), .B(n26184), .Z(n26189) );
  XOR U30951 ( .A(y[147]), .B(x[147]), .Z(n26184) );
  XOR U30952 ( .A(n26187), .B(n26186), .Z(n26185) );
  XOR U30953 ( .A(y[149]), .B(x[149]), .Z(n26186) );
  XOR U30954 ( .A(y[148]), .B(x[148]), .Z(n26187) );
  XOR U30955 ( .A(n26179), .B(n26178), .Z(n26188) );
  XOR U30956 ( .A(n26181), .B(n26180), .Z(n26178) );
  XOR U30957 ( .A(y[146]), .B(x[146]), .Z(n26180) );
  XOR U30958 ( .A(y[145]), .B(x[145]), .Z(n26181) );
  XOR U30959 ( .A(y[144]), .B(x[144]), .Z(n26179) );
  XNOR U30960 ( .A(n26172), .B(n26171), .Z(n26174) );
  XNOR U30961 ( .A(n26168), .B(n26167), .Z(n26171) );
  XOR U30962 ( .A(n26170), .B(n26169), .Z(n26167) );
  XOR U30963 ( .A(y[143]), .B(x[143]), .Z(n26169) );
  XOR U30964 ( .A(y[142]), .B(x[142]), .Z(n26170) );
  XOR U30965 ( .A(y[141]), .B(x[141]), .Z(n26168) );
  XOR U30966 ( .A(n26162), .B(n26161), .Z(n26172) );
  XOR U30967 ( .A(n26164), .B(n26163), .Z(n26161) );
  XOR U30968 ( .A(y[140]), .B(x[140]), .Z(n26163) );
  XOR U30969 ( .A(y[139]), .B(x[139]), .Z(n26164) );
  XOR U30970 ( .A(y[138]), .B(x[138]), .Z(n26162) );
  XNOR U30971 ( .A(n26139), .B(n26138), .Z(n26156) );
  XNOR U30972 ( .A(n26153), .B(n26154), .Z(n26138) );
  XOR U30973 ( .A(n26150), .B(n26149), .Z(n26154) );
  XOR U30974 ( .A(y[135]), .B(x[135]), .Z(n26149) );
  XOR U30975 ( .A(n26152), .B(n26151), .Z(n26150) );
  XOR U30976 ( .A(y[137]), .B(x[137]), .Z(n26151) );
  XOR U30977 ( .A(y[136]), .B(x[136]), .Z(n26152) );
  XOR U30978 ( .A(n26144), .B(n26143), .Z(n26153) );
  XOR U30979 ( .A(n26146), .B(n26145), .Z(n26143) );
  XOR U30980 ( .A(y[134]), .B(x[134]), .Z(n26145) );
  XOR U30981 ( .A(y[133]), .B(x[133]), .Z(n26146) );
  XOR U30982 ( .A(y[132]), .B(x[132]), .Z(n26144) );
  XNOR U30983 ( .A(n26137), .B(n26136), .Z(n26139) );
  XNOR U30984 ( .A(n26133), .B(n26132), .Z(n26136) );
  XOR U30985 ( .A(n26135), .B(n26134), .Z(n26132) );
  XOR U30986 ( .A(y[131]), .B(x[131]), .Z(n26134) );
  XOR U30987 ( .A(y[130]), .B(x[130]), .Z(n26135) );
  XOR U30988 ( .A(y[129]), .B(x[129]), .Z(n26133) );
  XOR U30989 ( .A(n26127), .B(n26126), .Z(n26137) );
  XOR U30990 ( .A(n26129), .B(n26128), .Z(n26126) );
  XOR U30991 ( .A(y[128]), .B(x[128]), .Z(n26128) );
  XOR U30992 ( .A(y[127]), .B(x[127]), .Z(n26129) );
  XOR U30993 ( .A(y[126]), .B(x[126]), .Z(n26127) );
  NAND U30994 ( .A(n26190), .B(n26191), .Z(N27993) );
  NAND U30995 ( .A(n26192), .B(n26193), .Z(n26191) );
  NANDN U30996 ( .A(n26194), .B(n26195), .Z(n26193) );
  NANDN U30997 ( .A(n26195), .B(n26194), .Z(n26190) );
  XOR U30998 ( .A(n26194), .B(n26196), .Z(N27992) );
  XNOR U30999 ( .A(n26192), .B(n26195), .Z(n26196) );
  NAND U31000 ( .A(n26197), .B(n26198), .Z(n26195) );
  NAND U31001 ( .A(n26199), .B(n26200), .Z(n26198) );
  NANDN U31002 ( .A(n26201), .B(n26202), .Z(n26200) );
  NANDN U31003 ( .A(n26202), .B(n26201), .Z(n26197) );
  AND U31004 ( .A(n26203), .B(n26204), .Z(n26192) );
  NAND U31005 ( .A(n26205), .B(n26206), .Z(n26204) );
  OR U31006 ( .A(n26207), .B(n26208), .Z(n26206) );
  NAND U31007 ( .A(n26208), .B(n26207), .Z(n26203) );
  IV U31008 ( .A(n26209), .Z(n26208) );
  AND U31009 ( .A(n26210), .B(n26211), .Z(n26194) );
  NAND U31010 ( .A(n26212), .B(n26213), .Z(n26211) );
  NANDN U31011 ( .A(n26214), .B(n26215), .Z(n26213) );
  NANDN U31012 ( .A(n26215), .B(n26214), .Z(n26210) );
  XOR U31013 ( .A(n26207), .B(n26216), .Z(N27991) );
  XOR U31014 ( .A(n26205), .B(n26209), .Z(n26216) );
  XNOR U31015 ( .A(n26202), .B(n26217), .Z(n26209) );
  XNOR U31016 ( .A(n26199), .B(n26201), .Z(n26217) );
  AND U31017 ( .A(n26218), .B(n26219), .Z(n26201) );
  NANDN U31018 ( .A(n26220), .B(n26221), .Z(n26219) );
  NANDN U31019 ( .A(n26222), .B(n26223), .Z(n26221) );
  IV U31020 ( .A(n26224), .Z(n26223) );
  NAND U31021 ( .A(n26224), .B(n26222), .Z(n26218) );
  AND U31022 ( .A(n26225), .B(n26226), .Z(n26199) );
  NAND U31023 ( .A(n26227), .B(n26228), .Z(n26226) );
  OR U31024 ( .A(n26229), .B(n26230), .Z(n26228) );
  NAND U31025 ( .A(n26230), .B(n26229), .Z(n26225) );
  IV U31026 ( .A(n26231), .Z(n26230) );
  NAND U31027 ( .A(n26232), .B(n26233), .Z(n26202) );
  NANDN U31028 ( .A(n26234), .B(n26235), .Z(n26233) );
  NAND U31029 ( .A(n26236), .B(n26237), .Z(n26235) );
  OR U31030 ( .A(n26237), .B(n26236), .Z(n26232) );
  IV U31031 ( .A(n26238), .Z(n26236) );
  AND U31032 ( .A(n26239), .B(n26240), .Z(n26205) );
  NAND U31033 ( .A(n26241), .B(n26242), .Z(n26240) );
  NANDN U31034 ( .A(n26243), .B(n26244), .Z(n26242) );
  NANDN U31035 ( .A(n26244), .B(n26243), .Z(n26239) );
  XOR U31036 ( .A(n26215), .B(n26245), .Z(n26207) );
  XNOR U31037 ( .A(n26212), .B(n26214), .Z(n26245) );
  AND U31038 ( .A(n26246), .B(n26247), .Z(n26214) );
  NANDN U31039 ( .A(n26248), .B(n26249), .Z(n26247) );
  NANDN U31040 ( .A(n26250), .B(n26251), .Z(n26249) );
  IV U31041 ( .A(n26252), .Z(n26251) );
  NAND U31042 ( .A(n26252), .B(n26250), .Z(n26246) );
  AND U31043 ( .A(n26253), .B(n26254), .Z(n26212) );
  NAND U31044 ( .A(n26255), .B(n26256), .Z(n26254) );
  OR U31045 ( .A(n26257), .B(n26258), .Z(n26256) );
  NAND U31046 ( .A(n26258), .B(n26257), .Z(n26253) );
  IV U31047 ( .A(n26259), .Z(n26258) );
  NAND U31048 ( .A(n26260), .B(n26261), .Z(n26215) );
  NANDN U31049 ( .A(n26262), .B(n26263), .Z(n26261) );
  NAND U31050 ( .A(n26264), .B(n26265), .Z(n26263) );
  OR U31051 ( .A(n26265), .B(n26264), .Z(n26260) );
  IV U31052 ( .A(n26266), .Z(n26264) );
  XOR U31053 ( .A(n26241), .B(n26267), .Z(N27990) );
  XNOR U31054 ( .A(n26244), .B(n26243), .Z(n26267) );
  XNOR U31055 ( .A(n26255), .B(n26268), .Z(n26243) );
  XOR U31056 ( .A(n26259), .B(n26257), .Z(n26268) );
  XOR U31057 ( .A(n26265), .B(n26269), .Z(n26257) );
  XOR U31058 ( .A(n26262), .B(n26266), .Z(n26269) );
  NAND U31059 ( .A(n26270), .B(n26271), .Z(n26266) );
  NAND U31060 ( .A(n26272), .B(n26273), .Z(n26271) );
  NAND U31061 ( .A(n26274), .B(n26275), .Z(n26270) );
  AND U31062 ( .A(n26276), .B(n26277), .Z(n26262) );
  NAND U31063 ( .A(n26278), .B(n26279), .Z(n26277) );
  NAND U31064 ( .A(n26280), .B(n26281), .Z(n26276) );
  NANDN U31065 ( .A(n26282), .B(n26283), .Z(n26265) );
  NANDN U31066 ( .A(n26284), .B(n26285), .Z(n26259) );
  XNOR U31067 ( .A(n26250), .B(n26286), .Z(n26255) );
  XOR U31068 ( .A(n26248), .B(n26252), .Z(n26286) );
  NAND U31069 ( .A(n26287), .B(n26288), .Z(n26252) );
  NAND U31070 ( .A(n26289), .B(n26290), .Z(n26288) );
  NAND U31071 ( .A(n26291), .B(n26292), .Z(n26287) );
  AND U31072 ( .A(n26293), .B(n26294), .Z(n26248) );
  NAND U31073 ( .A(n26295), .B(n26296), .Z(n26294) );
  NAND U31074 ( .A(n26297), .B(n26298), .Z(n26293) );
  AND U31075 ( .A(n26299), .B(n26300), .Z(n26250) );
  NAND U31076 ( .A(n26301), .B(n26302), .Z(n26244) );
  XNOR U31077 ( .A(n26227), .B(n26303), .Z(n26241) );
  XOR U31078 ( .A(n26231), .B(n26229), .Z(n26303) );
  XOR U31079 ( .A(n26237), .B(n26304), .Z(n26229) );
  XOR U31080 ( .A(n26234), .B(n26238), .Z(n26304) );
  NAND U31081 ( .A(n26305), .B(n26306), .Z(n26238) );
  NAND U31082 ( .A(n26307), .B(n26308), .Z(n26306) );
  NAND U31083 ( .A(n26309), .B(n26310), .Z(n26305) );
  AND U31084 ( .A(n26311), .B(n26312), .Z(n26234) );
  NAND U31085 ( .A(n26313), .B(n26314), .Z(n26312) );
  NAND U31086 ( .A(n26315), .B(n26316), .Z(n26311) );
  NANDN U31087 ( .A(n26317), .B(n26318), .Z(n26237) );
  NANDN U31088 ( .A(n26319), .B(n26320), .Z(n26231) );
  XNOR U31089 ( .A(n26222), .B(n26321), .Z(n26227) );
  XOR U31090 ( .A(n26220), .B(n26224), .Z(n26321) );
  NAND U31091 ( .A(n26322), .B(n26323), .Z(n26224) );
  NAND U31092 ( .A(n26324), .B(n26325), .Z(n26323) );
  NAND U31093 ( .A(n26326), .B(n26327), .Z(n26322) );
  AND U31094 ( .A(n26328), .B(n26329), .Z(n26220) );
  NAND U31095 ( .A(n26330), .B(n26331), .Z(n26329) );
  NAND U31096 ( .A(n26332), .B(n26333), .Z(n26328) );
  AND U31097 ( .A(n26334), .B(n26335), .Z(n26222) );
  XOR U31098 ( .A(n26302), .B(n26301), .Z(N27989) );
  XNOR U31099 ( .A(n26320), .B(n26319), .Z(n26301) );
  XNOR U31100 ( .A(n26334), .B(n26335), .Z(n26319) );
  XOR U31101 ( .A(n26331), .B(n26330), .Z(n26335) );
  XOR U31102 ( .A(y[123]), .B(x[123]), .Z(n26330) );
  XOR U31103 ( .A(n26333), .B(n26332), .Z(n26331) );
  XOR U31104 ( .A(y[125]), .B(x[125]), .Z(n26332) );
  XOR U31105 ( .A(y[124]), .B(x[124]), .Z(n26333) );
  XOR U31106 ( .A(n26325), .B(n26324), .Z(n26334) );
  XOR U31107 ( .A(n26327), .B(n26326), .Z(n26324) );
  XOR U31108 ( .A(y[122]), .B(x[122]), .Z(n26326) );
  XOR U31109 ( .A(y[121]), .B(x[121]), .Z(n26327) );
  XOR U31110 ( .A(y[120]), .B(x[120]), .Z(n26325) );
  XNOR U31111 ( .A(n26318), .B(n26317), .Z(n26320) );
  XNOR U31112 ( .A(n26314), .B(n26313), .Z(n26317) );
  XOR U31113 ( .A(n26316), .B(n26315), .Z(n26313) );
  XOR U31114 ( .A(y[119]), .B(x[119]), .Z(n26315) );
  XOR U31115 ( .A(y[118]), .B(x[118]), .Z(n26316) );
  XOR U31116 ( .A(y[117]), .B(x[117]), .Z(n26314) );
  XOR U31117 ( .A(n26308), .B(n26307), .Z(n26318) );
  XOR U31118 ( .A(n26310), .B(n26309), .Z(n26307) );
  XOR U31119 ( .A(y[116]), .B(x[116]), .Z(n26309) );
  XOR U31120 ( .A(y[115]), .B(x[115]), .Z(n26310) );
  XOR U31121 ( .A(y[114]), .B(x[114]), .Z(n26308) );
  XNOR U31122 ( .A(n26285), .B(n26284), .Z(n26302) );
  XNOR U31123 ( .A(n26299), .B(n26300), .Z(n26284) );
  XOR U31124 ( .A(n26296), .B(n26295), .Z(n26300) );
  XOR U31125 ( .A(y[111]), .B(x[111]), .Z(n26295) );
  XOR U31126 ( .A(n26298), .B(n26297), .Z(n26296) );
  XOR U31127 ( .A(y[113]), .B(x[113]), .Z(n26297) );
  XOR U31128 ( .A(y[112]), .B(x[112]), .Z(n26298) );
  XOR U31129 ( .A(n26290), .B(n26289), .Z(n26299) );
  XOR U31130 ( .A(n26292), .B(n26291), .Z(n26289) );
  XOR U31131 ( .A(y[110]), .B(x[110]), .Z(n26291) );
  XOR U31132 ( .A(y[109]), .B(x[109]), .Z(n26292) );
  XOR U31133 ( .A(y[108]), .B(x[108]), .Z(n26290) );
  XNOR U31134 ( .A(n26283), .B(n26282), .Z(n26285) );
  XNOR U31135 ( .A(n26279), .B(n26278), .Z(n26282) );
  XOR U31136 ( .A(n26281), .B(n26280), .Z(n26278) );
  XOR U31137 ( .A(y[107]), .B(x[107]), .Z(n26280) );
  XOR U31138 ( .A(y[106]), .B(x[106]), .Z(n26281) );
  XOR U31139 ( .A(y[105]), .B(x[105]), .Z(n26279) );
  XOR U31140 ( .A(n26273), .B(n26272), .Z(n26283) );
  XOR U31141 ( .A(n26275), .B(n26274), .Z(n26272) );
  XOR U31142 ( .A(y[104]), .B(x[104]), .Z(n26274) );
  XOR U31143 ( .A(y[103]), .B(x[103]), .Z(n26275) );
  XOR U31144 ( .A(y[102]), .B(x[102]), .Z(n26273) );
  NAND U31145 ( .A(n26336), .B(n26337), .Z(N27981) );
  NAND U31146 ( .A(n26338), .B(n26339), .Z(n26337) );
  NANDN U31147 ( .A(n26340), .B(n26341), .Z(n26339) );
  NANDN U31148 ( .A(n26341), .B(n26340), .Z(n26336) );
  XOR U31149 ( .A(n26340), .B(n26342), .Z(N27980) );
  XNOR U31150 ( .A(n26338), .B(n26341), .Z(n26342) );
  NAND U31151 ( .A(n26343), .B(n26344), .Z(n26341) );
  NAND U31152 ( .A(n26345), .B(n26346), .Z(n26344) );
  NANDN U31153 ( .A(n26347), .B(n26348), .Z(n26346) );
  NANDN U31154 ( .A(n26348), .B(n26347), .Z(n26343) );
  AND U31155 ( .A(n26349), .B(n26350), .Z(n26338) );
  NAND U31156 ( .A(n26351), .B(n26352), .Z(n26350) );
  OR U31157 ( .A(n26353), .B(n26354), .Z(n26352) );
  NAND U31158 ( .A(n26354), .B(n26353), .Z(n26349) );
  IV U31159 ( .A(n26355), .Z(n26354) );
  AND U31160 ( .A(n26356), .B(n26357), .Z(n26340) );
  NAND U31161 ( .A(n26358), .B(n26359), .Z(n26357) );
  NANDN U31162 ( .A(n26360), .B(n26361), .Z(n26359) );
  NANDN U31163 ( .A(n26361), .B(n26360), .Z(n26356) );
  XOR U31164 ( .A(n26353), .B(n26362), .Z(N27979) );
  XOR U31165 ( .A(n26351), .B(n26355), .Z(n26362) );
  XNOR U31166 ( .A(n26348), .B(n26363), .Z(n26355) );
  XNOR U31167 ( .A(n26345), .B(n26347), .Z(n26363) );
  AND U31168 ( .A(n26364), .B(n26365), .Z(n26347) );
  NANDN U31169 ( .A(n26366), .B(n26367), .Z(n26365) );
  NANDN U31170 ( .A(n26368), .B(n26369), .Z(n26367) );
  IV U31171 ( .A(n26370), .Z(n26369) );
  NAND U31172 ( .A(n26370), .B(n26368), .Z(n26364) );
  AND U31173 ( .A(n26371), .B(n26372), .Z(n26345) );
  NAND U31174 ( .A(n26373), .B(n26374), .Z(n26372) );
  OR U31175 ( .A(n26375), .B(n26376), .Z(n26374) );
  NAND U31176 ( .A(n26376), .B(n26375), .Z(n26371) );
  IV U31177 ( .A(n26377), .Z(n26376) );
  NAND U31178 ( .A(n26378), .B(n26379), .Z(n26348) );
  NANDN U31179 ( .A(n26380), .B(n26381), .Z(n26379) );
  NAND U31180 ( .A(n26382), .B(n26383), .Z(n26381) );
  OR U31181 ( .A(n26383), .B(n26382), .Z(n26378) );
  IV U31182 ( .A(n26384), .Z(n26382) );
  AND U31183 ( .A(n26385), .B(n26386), .Z(n26351) );
  NAND U31184 ( .A(n26387), .B(n26388), .Z(n26386) );
  NANDN U31185 ( .A(n26389), .B(n26390), .Z(n26388) );
  NANDN U31186 ( .A(n26390), .B(n26389), .Z(n26385) );
  XOR U31187 ( .A(n26361), .B(n26391), .Z(n26353) );
  XNOR U31188 ( .A(n26358), .B(n26360), .Z(n26391) );
  AND U31189 ( .A(n26392), .B(n26393), .Z(n26360) );
  NANDN U31190 ( .A(n26394), .B(n26395), .Z(n26393) );
  NANDN U31191 ( .A(n26396), .B(n26397), .Z(n26395) );
  IV U31192 ( .A(n26398), .Z(n26397) );
  NAND U31193 ( .A(n26398), .B(n26396), .Z(n26392) );
  AND U31194 ( .A(n26399), .B(n26400), .Z(n26358) );
  NAND U31195 ( .A(n26401), .B(n26402), .Z(n26400) );
  OR U31196 ( .A(n26403), .B(n26404), .Z(n26402) );
  NAND U31197 ( .A(n26404), .B(n26403), .Z(n26399) );
  IV U31198 ( .A(n26405), .Z(n26404) );
  NAND U31199 ( .A(n26406), .B(n26407), .Z(n26361) );
  NANDN U31200 ( .A(n26408), .B(n26409), .Z(n26407) );
  NAND U31201 ( .A(n26410), .B(n26411), .Z(n26409) );
  OR U31202 ( .A(n26411), .B(n26410), .Z(n26406) );
  IV U31203 ( .A(n26412), .Z(n26410) );
  XOR U31204 ( .A(n26387), .B(n26413), .Z(N27978) );
  XNOR U31205 ( .A(n26390), .B(n26389), .Z(n26413) );
  XNOR U31206 ( .A(n26401), .B(n26414), .Z(n26389) );
  XOR U31207 ( .A(n26405), .B(n26403), .Z(n26414) );
  XOR U31208 ( .A(n26411), .B(n26415), .Z(n26403) );
  XOR U31209 ( .A(n26408), .B(n26412), .Z(n26415) );
  NAND U31210 ( .A(n26416), .B(n26417), .Z(n26412) );
  NAND U31211 ( .A(n26418), .B(n26419), .Z(n26417) );
  NAND U31212 ( .A(n26420), .B(n26421), .Z(n26416) );
  AND U31213 ( .A(n26422), .B(n26423), .Z(n26408) );
  NAND U31214 ( .A(n26424), .B(n26425), .Z(n26423) );
  NAND U31215 ( .A(n26426), .B(n26427), .Z(n26422) );
  NANDN U31216 ( .A(n26428), .B(n26429), .Z(n26411) );
  NANDN U31217 ( .A(n26430), .B(n26431), .Z(n26405) );
  XNOR U31218 ( .A(n26396), .B(n26432), .Z(n26401) );
  XOR U31219 ( .A(n26394), .B(n26398), .Z(n26432) );
  NAND U31220 ( .A(n26433), .B(n26434), .Z(n26398) );
  NAND U31221 ( .A(n26435), .B(n26436), .Z(n26434) );
  NAND U31222 ( .A(n26437), .B(n26438), .Z(n26433) );
  AND U31223 ( .A(n26439), .B(n26440), .Z(n26394) );
  NAND U31224 ( .A(n26441), .B(n26442), .Z(n26440) );
  NAND U31225 ( .A(n26443), .B(n26444), .Z(n26439) );
  AND U31226 ( .A(n26445), .B(n26446), .Z(n26396) );
  NAND U31227 ( .A(n26447), .B(n26448), .Z(n26390) );
  XNOR U31228 ( .A(n26373), .B(n26449), .Z(n26387) );
  XOR U31229 ( .A(n26377), .B(n26375), .Z(n26449) );
  XOR U31230 ( .A(n26383), .B(n26450), .Z(n26375) );
  XOR U31231 ( .A(n26380), .B(n26384), .Z(n26450) );
  NAND U31232 ( .A(n26451), .B(n26452), .Z(n26384) );
  NAND U31233 ( .A(n26453), .B(n26454), .Z(n26452) );
  NAND U31234 ( .A(n26455), .B(n26456), .Z(n26451) );
  AND U31235 ( .A(n26457), .B(n26458), .Z(n26380) );
  NAND U31236 ( .A(n26459), .B(n26460), .Z(n26458) );
  NAND U31237 ( .A(n26461), .B(n26462), .Z(n26457) );
  NANDN U31238 ( .A(n26463), .B(n26464), .Z(n26383) );
  NANDN U31239 ( .A(n26465), .B(n26466), .Z(n26377) );
  XNOR U31240 ( .A(n26368), .B(n26467), .Z(n26373) );
  XOR U31241 ( .A(n26366), .B(n26370), .Z(n26467) );
  NAND U31242 ( .A(n26468), .B(n26469), .Z(n26370) );
  NAND U31243 ( .A(n26470), .B(n26471), .Z(n26469) );
  NAND U31244 ( .A(n26472), .B(n26473), .Z(n26468) );
  AND U31245 ( .A(n26474), .B(n26475), .Z(n26366) );
  NAND U31246 ( .A(n26476), .B(n26477), .Z(n26475) );
  NAND U31247 ( .A(n26478), .B(n26479), .Z(n26474) );
  AND U31248 ( .A(n26480), .B(n26481), .Z(n26368) );
  XOR U31249 ( .A(n26448), .B(n26447), .Z(N27977) );
  XNOR U31250 ( .A(n26466), .B(n26465), .Z(n26447) );
  XNOR U31251 ( .A(n26480), .B(n26481), .Z(n26465) );
  XOR U31252 ( .A(n26477), .B(n26476), .Z(n26481) );
  XOR U31253 ( .A(y[99]), .B(x[99]), .Z(n26476) );
  XOR U31254 ( .A(n26479), .B(n26478), .Z(n26477) );
  XOR U31255 ( .A(y[101]), .B(x[101]), .Z(n26478) );
  XOR U31256 ( .A(y[100]), .B(x[100]), .Z(n26479) );
  XOR U31257 ( .A(n26471), .B(n26470), .Z(n26480) );
  XOR U31258 ( .A(n26473), .B(n26472), .Z(n26470) );
  XOR U31259 ( .A(y[98]), .B(x[98]), .Z(n26472) );
  XOR U31260 ( .A(y[97]), .B(x[97]), .Z(n26473) );
  XOR U31261 ( .A(y[96]), .B(x[96]), .Z(n26471) );
  XNOR U31262 ( .A(n26464), .B(n26463), .Z(n26466) );
  XNOR U31263 ( .A(n26460), .B(n26459), .Z(n26463) );
  XOR U31264 ( .A(n26462), .B(n26461), .Z(n26459) );
  XOR U31265 ( .A(y[95]), .B(x[95]), .Z(n26461) );
  XOR U31266 ( .A(y[94]), .B(x[94]), .Z(n26462) );
  XOR U31267 ( .A(y[93]), .B(x[93]), .Z(n26460) );
  XOR U31268 ( .A(n26454), .B(n26453), .Z(n26464) );
  XOR U31269 ( .A(n26456), .B(n26455), .Z(n26453) );
  XOR U31270 ( .A(y[92]), .B(x[92]), .Z(n26455) );
  XOR U31271 ( .A(y[91]), .B(x[91]), .Z(n26456) );
  XOR U31272 ( .A(y[90]), .B(x[90]), .Z(n26454) );
  XNOR U31273 ( .A(n26431), .B(n26430), .Z(n26448) );
  XNOR U31274 ( .A(n26445), .B(n26446), .Z(n26430) );
  XOR U31275 ( .A(n26442), .B(n26441), .Z(n26446) );
  XOR U31276 ( .A(y[87]), .B(x[87]), .Z(n26441) );
  XOR U31277 ( .A(n26444), .B(n26443), .Z(n26442) );
  XOR U31278 ( .A(y[89]), .B(x[89]), .Z(n26443) );
  XOR U31279 ( .A(y[88]), .B(x[88]), .Z(n26444) );
  XOR U31280 ( .A(n26436), .B(n26435), .Z(n26445) );
  XOR U31281 ( .A(n26438), .B(n26437), .Z(n26435) );
  XOR U31282 ( .A(y[86]), .B(x[86]), .Z(n26437) );
  XOR U31283 ( .A(y[85]), .B(x[85]), .Z(n26438) );
  XOR U31284 ( .A(y[84]), .B(x[84]), .Z(n26436) );
  XNOR U31285 ( .A(n26429), .B(n26428), .Z(n26431) );
  XNOR U31286 ( .A(n26425), .B(n26424), .Z(n26428) );
  XOR U31287 ( .A(n26427), .B(n26426), .Z(n26424) );
  XOR U31288 ( .A(y[83]), .B(x[83]), .Z(n26426) );
  XOR U31289 ( .A(y[82]), .B(x[82]), .Z(n26427) );
  XOR U31290 ( .A(y[81]), .B(x[81]), .Z(n26425) );
  XOR U31291 ( .A(n26419), .B(n26418), .Z(n26429) );
  XOR U31292 ( .A(n26421), .B(n26420), .Z(n26418) );
  XOR U31293 ( .A(y[80]), .B(x[80]), .Z(n26420) );
  XOR U31294 ( .A(y[79]), .B(x[79]), .Z(n26421) );
  XOR U31295 ( .A(y[78]), .B(x[78]), .Z(n26419) );
  NAND U31296 ( .A(n26482), .B(n26483), .Z(N27969) );
  NAND U31297 ( .A(n26484), .B(n26485), .Z(n26483) );
  NANDN U31298 ( .A(n26486), .B(n26487), .Z(n26485) );
  NANDN U31299 ( .A(n26487), .B(n26486), .Z(n26482) );
  XOR U31300 ( .A(n26486), .B(n26488), .Z(N27968) );
  XNOR U31301 ( .A(n26484), .B(n26487), .Z(n26488) );
  NAND U31302 ( .A(n26489), .B(n26490), .Z(n26487) );
  NAND U31303 ( .A(n26491), .B(n26492), .Z(n26490) );
  NANDN U31304 ( .A(n26493), .B(n26494), .Z(n26492) );
  NANDN U31305 ( .A(n26494), .B(n26493), .Z(n26489) );
  AND U31306 ( .A(n26495), .B(n26496), .Z(n26484) );
  NAND U31307 ( .A(n26497), .B(n26498), .Z(n26496) );
  OR U31308 ( .A(n26499), .B(n26500), .Z(n26498) );
  NAND U31309 ( .A(n26500), .B(n26499), .Z(n26495) );
  IV U31310 ( .A(n26501), .Z(n26500) );
  AND U31311 ( .A(n26502), .B(n26503), .Z(n26486) );
  NAND U31312 ( .A(n26504), .B(n26505), .Z(n26503) );
  NANDN U31313 ( .A(n26506), .B(n26507), .Z(n26505) );
  NANDN U31314 ( .A(n26507), .B(n26506), .Z(n26502) );
  XOR U31315 ( .A(n26499), .B(n26508), .Z(N27967) );
  XOR U31316 ( .A(n26497), .B(n26501), .Z(n26508) );
  XNOR U31317 ( .A(n26494), .B(n26509), .Z(n26501) );
  XNOR U31318 ( .A(n26491), .B(n26493), .Z(n26509) );
  AND U31319 ( .A(n26510), .B(n26511), .Z(n26493) );
  NANDN U31320 ( .A(n26512), .B(n26513), .Z(n26511) );
  NANDN U31321 ( .A(n26514), .B(n26515), .Z(n26513) );
  IV U31322 ( .A(n26516), .Z(n26515) );
  NAND U31323 ( .A(n26516), .B(n26514), .Z(n26510) );
  AND U31324 ( .A(n26517), .B(n26518), .Z(n26491) );
  NAND U31325 ( .A(n26519), .B(n26520), .Z(n26518) );
  OR U31326 ( .A(n26521), .B(n26522), .Z(n26520) );
  NAND U31327 ( .A(n26522), .B(n26521), .Z(n26517) );
  IV U31328 ( .A(n26523), .Z(n26522) );
  NAND U31329 ( .A(n26524), .B(n26525), .Z(n26494) );
  NANDN U31330 ( .A(n26526), .B(n26527), .Z(n26525) );
  NAND U31331 ( .A(n26528), .B(n26529), .Z(n26527) );
  OR U31332 ( .A(n26529), .B(n26528), .Z(n26524) );
  IV U31333 ( .A(n26530), .Z(n26528) );
  AND U31334 ( .A(n26531), .B(n26532), .Z(n26497) );
  NAND U31335 ( .A(n26533), .B(n26534), .Z(n26532) );
  NANDN U31336 ( .A(n26535), .B(n26536), .Z(n26534) );
  NANDN U31337 ( .A(n26536), .B(n26535), .Z(n26531) );
  XOR U31338 ( .A(n26507), .B(n26537), .Z(n26499) );
  XNOR U31339 ( .A(n26504), .B(n26506), .Z(n26537) );
  AND U31340 ( .A(n26538), .B(n26539), .Z(n26506) );
  NANDN U31341 ( .A(n26540), .B(n26541), .Z(n26539) );
  NANDN U31342 ( .A(n26542), .B(n26543), .Z(n26541) );
  IV U31343 ( .A(n26544), .Z(n26543) );
  NAND U31344 ( .A(n26544), .B(n26542), .Z(n26538) );
  AND U31345 ( .A(n26545), .B(n26546), .Z(n26504) );
  NAND U31346 ( .A(n26547), .B(n26548), .Z(n26546) );
  OR U31347 ( .A(n26549), .B(n26550), .Z(n26548) );
  NAND U31348 ( .A(n26550), .B(n26549), .Z(n26545) );
  IV U31349 ( .A(n26551), .Z(n26550) );
  NAND U31350 ( .A(n26552), .B(n26553), .Z(n26507) );
  NANDN U31351 ( .A(n26554), .B(n26555), .Z(n26553) );
  NAND U31352 ( .A(n26556), .B(n26557), .Z(n26555) );
  OR U31353 ( .A(n26557), .B(n26556), .Z(n26552) );
  IV U31354 ( .A(n26558), .Z(n26556) );
  XOR U31355 ( .A(n26533), .B(n26559), .Z(N27966) );
  XNOR U31356 ( .A(n26536), .B(n26535), .Z(n26559) );
  XNOR U31357 ( .A(n26547), .B(n26560), .Z(n26535) );
  XOR U31358 ( .A(n26551), .B(n26549), .Z(n26560) );
  XOR U31359 ( .A(n26557), .B(n26561), .Z(n26549) );
  XOR U31360 ( .A(n26554), .B(n26558), .Z(n26561) );
  NAND U31361 ( .A(n26562), .B(n26563), .Z(n26558) );
  NAND U31362 ( .A(n26564), .B(n26565), .Z(n26563) );
  NAND U31363 ( .A(n26566), .B(n26567), .Z(n26562) );
  AND U31364 ( .A(n26568), .B(n26569), .Z(n26554) );
  NAND U31365 ( .A(n26570), .B(n26571), .Z(n26569) );
  NAND U31366 ( .A(n26572), .B(n26573), .Z(n26568) );
  NANDN U31367 ( .A(n26574), .B(n26575), .Z(n26557) );
  NANDN U31368 ( .A(n26576), .B(n26577), .Z(n26551) );
  XNOR U31369 ( .A(n26542), .B(n26578), .Z(n26547) );
  XOR U31370 ( .A(n26540), .B(n26544), .Z(n26578) );
  NAND U31371 ( .A(n26579), .B(n26580), .Z(n26544) );
  NAND U31372 ( .A(n26581), .B(n26582), .Z(n26580) );
  NAND U31373 ( .A(n26583), .B(n26584), .Z(n26579) );
  AND U31374 ( .A(n26585), .B(n26586), .Z(n26540) );
  NAND U31375 ( .A(n26587), .B(n26588), .Z(n26586) );
  NAND U31376 ( .A(n26589), .B(n26590), .Z(n26585) );
  AND U31377 ( .A(n26591), .B(n26592), .Z(n26542) );
  NAND U31378 ( .A(n26593), .B(n26594), .Z(n26536) );
  XNOR U31379 ( .A(n26519), .B(n26595), .Z(n26533) );
  XOR U31380 ( .A(n26523), .B(n26521), .Z(n26595) );
  XOR U31381 ( .A(n26529), .B(n26596), .Z(n26521) );
  XOR U31382 ( .A(n26526), .B(n26530), .Z(n26596) );
  NAND U31383 ( .A(n26597), .B(n26598), .Z(n26530) );
  NAND U31384 ( .A(n26599), .B(n26600), .Z(n26598) );
  NAND U31385 ( .A(n26601), .B(n26602), .Z(n26597) );
  AND U31386 ( .A(n26603), .B(n26604), .Z(n26526) );
  NAND U31387 ( .A(n26605), .B(n26606), .Z(n26604) );
  NAND U31388 ( .A(n26607), .B(n26608), .Z(n26603) );
  NANDN U31389 ( .A(n26609), .B(n26610), .Z(n26529) );
  NANDN U31390 ( .A(n26611), .B(n26612), .Z(n26523) );
  XNOR U31391 ( .A(n26514), .B(n26613), .Z(n26519) );
  XOR U31392 ( .A(n26512), .B(n26516), .Z(n26613) );
  NAND U31393 ( .A(n26614), .B(n26615), .Z(n26516) );
  NAND U31394 ( .A(n26616), .B(n26617), .Z(n26615) );
  NAND U31395 ( .A(n26618), .B(n26619), .Z(n26614) );
  AND U31396 ( .A(n26620), .B(n26621), .Z(n26512) );
  NAND U31397 ( .A(n26622), .B(n26623), .Z(n26621) );
  NAND U31398 ( .A(n26624), .B(n26625), .Z(n26620) );
  AND U31399 ( .A(n26626), .B(n26627), .Z(n26514) );
  XOR U31400 ( .A(n26594), .B(n26593), .Z(N27965) );
  XNOR U31401 ( .A(n26612), .B(n26611), .Z(n26593) );
  XNOR U31402 ( .A(n26626), .B(n26627), .Z(n26611) );
  XOR U31403 ( .A(n26623), .B(n26622), .Z(n26627) );
  XOR U31404 ( .A(y[75]), .B(x[75]), .Z(n26622) );
  XOR U31405 ( .A(n26625), .B(n26624), .Z(n26623) );
  XOR U31406 ( .A(y[77]), .B(x[77]), .Z(n26624) );
  XOR U31407 ( .A(y[76]), .B(x[76]), .Z(n26625) );
  XOR U31408 ( .A(n26617), .B(n26616), .Z(n26626) );
  XOR U31409 ( .A(n26619), .B(n26618), .Z(n26616) );
  XOR U31410 ( .A(y[74]), .B(x[74]), .Z(n26618) );
  XOR U31411 ( .A(y[73]), .B(x[73]), .Z(n26619) );
  XOR U31412 ( .A(y[72]), .B(x[72]), .Z(n26617) );
  XNOR U31413 ( .A(n26610), .B(n26609), .Z(n26612) );
  XNOR U31414 ( .A(n26606), .B(n26605), .Z(n26609) );
  XOR U31415 ( .A(n26608), .B(n26607), .Z(n26605) );
  XOR U31416 ( .A(y[71]), .B(x[71]), .Z(n26607) );
  XOR U31417 ( .A(y[70]), .B(x[70]), .Z(n26608) );
  XOR U31418 ( .A(y[69]), .B(x[69]), .Z(n26606) );
  XOR U31419 ( .A(n26600), .B(n26599), .Z(n26610) );
  XOR U31420 ( .A(n26602), .B(n26601), .Z(n26599) );
  XOR U31421 ( .A(y[68]), .B(x[68]), .Z(n26601) );
  XOR U31422 ( .A(y[67]), .B(x[67]), .Z(n26602) );
  XOR U31423 ( .A(y[66]), .B(x[66]), .Z(n26600) );
  XNOR U31424 ( .A(n26577), .B(n26576), .Z(n26594) );
  XNOR U31425 ( .A(n26591), .B(n26592), .Z(n26576) );
  XOR U31426 ( .A(n26588), .B(n26587), .Z(n26592) );
  XOR U31427 ( .A(y[63]), .B(x[63]), .Z(n26587) );
  XOR U31428 ( .A(n26590), .B(n26589), .Z(n26588) );
  XOR U31429 ( .A(y[65]), .B(x[65]), .Z(n26589) );
  XOR U31430 ( .A(y[64]), .B(x[64]), .Z(n26590) );
  XOR U31431 ( .A(n26582), .B(n26581), .Z(n26591) );
  XOR U31432 ( .A(n26584), .B(n26583), .Z(n26581) );
  XOR U31433 ( .A(y[62]), .B(x[62]), .Z(n26583) );
  XOR U31434 ( .A(y[61]), .B(x[61]), .Z(n26584) );
  XOR U31435 ( .A(y[60]), .B(x[60]), .Z(n26582) );
  XNOR U31436 ( .A(n26575), .B(n26574), .Z(n26577) );
  XNOR U31437 ( .A(n26571), .B(n26570), .Z(n26574) );
  XOR U31438 ( .A(n26573), .B(n26572), .Z(n26570) );
  XOR U31439 ( .A(y[59]), .B(x[59]), .Z(n26572) );
  XOR U31440 ( .A(y[58]), .B(x[58]), .Z(n26573) );
  XOR U31441 ( .A(y[57]), .B(x[57]), .Z(n26571) );
  XOR U31442 ( .A(n26565), .B(n26564), .Z(n26575) );
  XOR U31443 ( .A(n26567), .B(n26566), .Z(n26564) );
  XOR U31444 ( .A(y[56]), .B(x[56]), .Z(n26566) );
  XOR U31445 ( .A(y[55]), .B(x[55]), .Z(n26567) );
  XOR U31446 ( .A(y[54]), .B(x[54]), .Z(n26565) );
  NAND U31447 ( .A(n26628), .B(n26629), .Z(N27957) );
  NAND U31448 ( .A(n26630), .B(n26631), .Z(n26629) );
  NANDN U31449 ( .A(n26632), .B(n26633), .Z(n26631) );
  NANDN U31450 ( .A(n26633), .B(n26632), .Z(n26628) );
  XOR U31451 ( .A(n26632), .B(n26634), .Z(N27956) );
  XNOR U31452 ( .A(n26630), .B(n26633), .Z(n26634) );
  NAND U31453 ( .A(n26635), .B(n26636), .Z(n26633) );
  NAND U31454 ( .A(n26637), .B(n26638), .Z(n26636) );
  NANDN U31455 ( .A(n26639), .B(n26640), .Z(n26638) );
  NANDN U31456 ( .A(n26640), .B(n26639), .Z(n26635) );
  AND U31457 ( .A(n26641), .B(n26642), .Z(n26630) );
  NAND U31458 ( .A(n26643), .B(n26644), .Z(n26642) );
  OR U31459 ( .A(n26645), .B(n26646), .Z(n26644) );
  NAND U31460 ( .A(n26646), .B(n26645), .Z(n26641) );
  IV U31461 ( .A(n26647), .Z(n26646) );
  AND U31462 ( .A(n26648), .B(n26649), .Z(n26632) );
  NAND U31463 ( .A(n26650), .B(n26651), .Z(n26649) );
  NANDN U31464 ( .A(n26652), .B(n26653), .Z(n26651) );
  NANDN U31465 ( .A(n26653), .B(n26652), .Z(n26648) );
  XOR U31466 ( .A(n26645), .B(n26654), .Z(N27955) );
  XOR U31467 ( .A(n26643), .B(n26647), .Z(n26654) );
  XNOR U31468 ( .A(n26640), .B(n26655), .Z(n26647) );
  XNOR U31469 ( .A(n26637), .B(n26639), .Z(n26655) );
  AND U31470 ( .A(n26656), .B(n26657), .Z(n26639) );
  NANDN U31471 ( .A(n26658), .B(n26659), .Z(n26657) );
  NANDN U31472 ( .A(n26660), .B(n26661), .Z(n26659) );
  IV U31473 ( .A(n26662), .Z(n26661) );
  NAND U31474 ( .A(n26662), .B(n26660), .Z(n26656) );
  AND U31475 ( .A(n26663), .B(n26664), .Z(n26637) );
  NAND U31476 ( .A(n26665), .B(n26666), .Z(n26664) );
  OR U31477 ( .A(n26667), .B(n26668), .Z(n26666) );
  NAND U31478 ( .A(n26668), .B(n26667), .Z(n26663) );
  IV U31479 ( .A(n26669), .Z(n26668) );
  NAND U31480 ( .A(n26670), .B(n26671), .Z(n26640) );
  NANDN U31481 ( .A(n26672), .B(n26673), .Z(n26671) );
  NAND U31482 ( .A(n26674), .B(n26675), .Z(n26673) );
  OR U31483 ( .A(n26675), .B(n26674), .Z(n26670) );
  IV U31484 ( .A(n26676), .Z(n26674) );
  AND U31485 ( .A(n26677), .B(n26678), .Z(n26643) );
  NAND U31486 ( .A(n26679), .B(n26680), .Z(n26678) );
  NANDN U31487 ( .A(n26681), .B(n26682), .Z(n26680) );
  NANDN U31488 ( .A(n26682), .B(n26681), .Z(n26677) );
  XOR U31489 ( .A(n26653), .B(n26683), .Z(n26645) );
  XNOR U31490 ( .A(n26650), .B(n26652), .Z(n26683) );
  AND U31491 ( .A(n26684), .B(n26685), .Z(n26652) );
  NANDN U31492 ( .A(n26686), .B(n26687), .Z(n26685) );
  NANDN U31493 ( .A(n26688), .B(n26689), .Z(n26687) );
  IV U31494 ( .A(n26690), .Z(n26689) );
  NAND U31495 ( .A(n26690), .B(n26688), .Z(n26684) );
  AND U31496 ( .A(n26691), .B(n26692), .Z(n26650) );
  NAND U31497 ( .A(n26693), .B(n26694), .Z(n26692) );
  OR U31498 ( .A(n26695), .B(n26696), .Z(n26694) );
  NAND U31499 ( .A(n26696), .B(n26695), .Z(n26691) );
  IV U31500 ( .A(n26697), .Z(n26696) );
  NAND U31501 ( .A(n26698), .B(n26699), .Z(n26653) );
  NANDN U31502 ( .A(n26700), .B(n26701), .Z(n26699) );
  NAND U31503 ( .A(n26702), .B(n26703), .Z(n26701) );
  OR U31504 ( .A(n26703), .B(n26702), .Z(n26698) );
  IV U31505 ( .A(n26704), .Z(n26702) );
  XOR U31506 ( .A(n26679), .B(n26705), .Z(N27954) );
  XNOR U31507 ( .A(n26682), .B(n26681), .Z(n26705) );
  XNOR U31508 ( .A(n26693), .B(n26706), .Z(n26681) );
  XOR U31509 ( .A(n26697), .B(n26695), .Z(n26706) );
  XOR U31510 ( .A(n26703), .B(n26707), .Z(n26695) );
  XOR U31511 ( .A(n26700), .B(n26704), .Z(n26707) );
  NAND U31512 ( .A(n26708), .B(n26709), .Z(n26704) );
  NAND U31513 ( .A(n26710), .B(n26711), .Z(n26709) );
  NAND U31514 ( .A(n26712), .B(n26713), .Z(n26708) );
  AND U31515 ( .A(n26714), .B(n26715), .Z(n26700) );
  NAND U31516 ( .A(n26716), .B(n26717), .Z(n26715) );
  NAND U31517 ( .A(n26718), .B(n26719), .Z(n26714) );
  NANDN U31518 ( .A(n26720), .B(n26721), .Z(n26703) );
  NANDN U31519 ( .A(n26722), .B(n26723), .Z(n26697) );
  XNOR U31520 ( .A(n26688), .B(n26724), .Z(n26693) );
  XOR U31521 ( .A(n26686), .B(n26690), .Z(n26724) );
  NAND U31522 ( .A(n26725), .B(n26726), .Z(n26690) );
  NAND U31523 ( .A(n26727), .B(n26728), .Z(n26726) );
  NAND U31524 ( .A(n26729), .B(n26730), .Z(n26725) );
  AND U31525 ( .A(n26731), .B(n26732), .Z(n26686) );
  NAND U31526 ( .A(n26733), .B(n26734), .Z(n26732) );
  NAND U31527 ( .A(n26735), .B(n26736), .Z(n26731) );
  AND U31528 ( .A(n26737), .B(n26738), .Z(n26688) );
  NAND U31529 ( .A(n26739), .B(n26740), .Z(n26682) );
  XNOR U31530 ( .A(n26665), .B(n26741), .Z(n26679) );
  XOR U31531 ( .A(n26669), .B(n26667), .Z(n26741) );
  XOR U31532 ( .A(n26675), .B(n26742), .Z(n26667) );
  XOR U31533 ( .A(n26672), .B(n26676), .Z(n26742) );
  NAND U31534 ( .A(n26743), .B(n26744), .Z(n26676) );
  NAND U31535 ( .A(n26745), .B(n26746), .Z(n26744) );
  NAND U31536 ( .A(n26747), .B(n26748), .Z(n26743) );
  AND U31537 ( .A(n26749), .B(n26750), .Z(n26672) );
  NAND U31538 ( .A(n26751), .B(n26752), .Z(n26750) );
  NAND U31539 ( .A(n26753), .B(n26754), .Z(n26749) );
  NANDN U31540 ( .A(n26755), .B(n26756), .Z(n26675) );
  NANDN U31541 ( .A(n26757), .B(n26758), .Z(n26669) );
  XNOR U31542 ( .A(n26660), .B(n26759), .Z(n26665) );
  XOR U31543 ( .A(n26658), .B(n26662), .Z(n26759) );
  NAND U31544 ( .A(n26760), .B(n26761), .Z(n26662) );
  NAND U31545 ( .A(n26762), .B(n26763), .Z(n26761) );
  NAND U31546 ( .A(n26764), .B(n26765), .Z(n26760) );
  AND U31547 ( .A(n26766), .B(n26767), .Z(n26658) );
  NAND U31548 ( .A(n26768), .B(n26769), .Z(n26767) );
  NAND U31549 ( .A(n26770), .B(n26771), .Z(n26766) );
  AND U31550 ( .A(n26772), .B(n26773), .Z(n26660) );
  XOR U31551 ( .A(n26740), .B(n26739), .Z(N27953) );
  XNOR U31552 ( .A(n26758), .B(n26757), .Z(n26739) );
  XNOR U31553 ( .A(n26772), .B(n26773), .Z(n26757) );
  XOR U31554 ( .A(n26769), .B(n26768), .Z(n26773) );
  XOR U31555 ( .A(y[51]), .B(x[51]), .Z(n26768) );
  XOR U31556 ( .A(n26771), .B(n26770), .Z(n26769) );
  XOR U31557 ( .A(y[53]), .B(x[53]), .Z(n26770) );
  XOR U31558 ( .A(y[52]), .B(x[52]), .Z(n26771) );
  XOR U31559 ( .A(n26763), .B(n26762), .Z(n26772) );
  XOR U31560 ( .A(n26765), .B(n26764), .Z(n26762) );
  XOR U31561 ( .A(y[50]), .B(x[50]), .Z(n26764) );
  XOR U31562 ( .A(y[49]), .B(x[49]), .Z(n26765) );
  XOR U31563 ( .A(y[48]), .B(x[48]), .Z(n26763) );
  XNOR U31564 ( .A(n26756), .B(n26755), .Z(n26758) );
  XNOR U31565 ( .A(n26752), .B(n26751), .Z(n26755) );
  XOR U31566 ( .A(n26754), .B(n26753), .Z(n26751) );
  XOR U31567 ( .A(y[47]), .B(x[47]), .Z(n26753) );
  XOR U31568 ( .A(y[46]), .B(x[46]), .Z(n26754) );
  XOR U31569 ( .A(y[45]), .B(x[45]), .Z(n26752) );
  XOR U31570 ( .A(n26746), .B(n26745), .Z(n26756) );
  XOR U31571 ( .A(n26748), .B(n26747), .Z(n26745) );
  XOR U31572 ( .A(y[44]), .B(x[44]), .Z(n26747) );
  XOR U31573 ( .A(y[43]), .B(x[43]), .Z(n26748) );
  XOR U31574 ( .A(y[42]), .B(x[42]), .Z(n26746) );
  XNOR U31575 ( .A(n26723), .B(n26722), .Z(n26740) );
  XNOR U31576 ( .A(n26737), .B(n26738), .Z(n26722) );
  XOR U31577 ( .A(n26734), .B(n26733), .Z(n26738) );
  XOR U31578 ( .A(y[39]), .B(x[39]), .Z(n26733) );
  XOR U31579 ( .A(n26736), .B(n26735), .Z(n26734) );
  XOR U31580 ( .A(y[41]), .B(x[41]), .Z(n26735) );
  XOR U31581 ( .A(y[40]), .B(x[40]), .Z(n26736) );
  XOR U31582 ( .A(n26728), .B(n26727), .Z(n26737) );
  XOR U31583 ( .A(n26730), .B(n26729), .Z(n26727) );
  XOR U31584 ( .A(y[38]), .B(x[38]), .Z(n26729) );
  XOR U31585 ( .A(y[37]), .B(x[37]), .Z(n26730) );
  XOR U31586 ( .A(y[36]), .B(x[36]), .Z(n26728) );
  XNOR U31587 ( .A(n26721), .B(n26720), .Z(n26723) );
  XNOR U31588 ( .A(n26717), .B(n26716), .Z(n26720) );
  XOR U31589 ( .A(n26719), .B(n26718), .Z(n26716) );
  XOR U31590 ( .A(y[35]), .B(x[35]), .Z(n26718) );
  XOR U31591 ( .A(y[34]), .B(x[34]), .Z(n26719) );
  XOR U31592 ( .A(y[33]), .B(x[33]), .Z(n26717) );
  XOR U31593 ( .A(n26711), .B(n26710), .Z(n26721) );
  XOR U31594 ( .A(n26713), .B(n26712), .Z(n26710) );
  XOR U31595 ( .A(y[32]), .B(x[32]), .Z(n26712) );
  XOR U31596 ( .A(y[31]), .B(x[31]), .Z(n26713) );
  XOR U31597 ( .A(y[30]), .B(x[30]), .Z(n26711) );
  NAND U31598 ( .A(n26774), .B(n26775), .Z(N27945) );
  NAND U31599 ( .A(n26776), .B(n26777), .Z(n26775) );
  NANDN U31600 ( .A(n26778), .B(n26779), .Z(n26777) );
  NANDN U31601 ( .A(n26779), .B(n26778), .Z(n26774) );
  XOR U31602 ( .A(n26778), .B(n26780), .Z(N27944) );
  XNOR U31603 ( .A(n26776), .B(n26779), .Z(n26780) );
  NAND U31604 ( .A(n26781), .B(n26782), .Z(n26779) );
  NAND U31605 ( .A(n26783), .B(n26784), .Z(n26782) );
  NANDN U31606 ( .A(n26785), .B(n26786), .Z(n26784) );
  NANDN U31607 ( .A(n26786), .B(n26785), .Z(n26781) );
  AND U31608 ( .A(n26787), .B(n26788), .Z(n26776) );
  NAND U31609 ( .A(n26789), .B(n26790), .Z(n26788) );
  OR U31610 ( .A(n26791), .B(n26792), .Z(n26790) );
  NAND U31611 ( .A(n26792), .B(n26791), .Z(n26787) );
  IV U31612 ( .A(n26793), .Z(n26792) );
  AND U31613 ( .A(n26794), .B(n26795), .Z(n26778) );
  NAND U31614 ( .A(n26796), .B(n26797), .Z(n26795) );
  NANDN U31615 ( .A(n26798), .B(n26799), .Z(n26797) );
  NANDN U31616 ( .A(n26799), .B(n26798), .Z(n26794) );
  XOR U31617 ( .A(n26791), .B(n26800), .Z(N27943) );
  XOR U31618 ( .A(n26789), .B(n26793), .Z(n26800) );
  XNOR U31619 ( .A(n26786), .B(n26801), .Z(n26793) );
  XNOR U31620 ( .A(n26783), .B(n26785), .Z(n26801) );
  AND U31621 ( .A(n26802), .B(n26803), .Z(n26785) );
  NANDN U31622 ( .A(n26804), .B(n26805), .Z(n26803) );
  NANDN U31623 ( .A(n26806), .B(n26807), .Z(n26805) );
  IV U31624 ( .A(n26808), .Z(n26807) );
  NAND U31625 ( .A(n26808), .B(n26806), .Z(n26802) );
  AND U31626 ( .A(n26809), .B(n26810), .Z(n26783) );
  NAND U31627 ( .A(n26811), .B(n26812), .Z(n26810) );
  OR U31628 ( .A(n26813), .B(n26814), .Z(n26812) );
  NAND U31629 ( .A(n26814), .B(n26813), .Z(n26809) );
  IV U31630 ( .A(n26815), .Z(n26814) );
  NAND U31631 ( .A(n26816), .B(n26817), .Z(n26786) );
  NANDN U31632 ( .A(n26818), .B(n26819), .Z(n26817) );
  NAND U31633 ( .A(n26820), .B(n26821), .Z(n26819) );
  OR U31634 ( .A(n26821), .B(n26820), .Z(n26816) );
  IV U31635 ( .A(n26822), .Z(n26820) );
  AND U31636 ( .A(n26823), .B(n26824), .Z(n26789) );
  NAND U31637 ( .A(n26825), .B(n26826), .Z(n26824) );
  NANDN U31638 ( .A(n26827), .B(n26828), .Z(n26826) );
  NANDN U31639 ( .A(n26828), .B(n26827), .Z(n26823) );
  XOR U31640 ( .A(n26799), .B(n26829), .Z(n26791) );
  XNOR U31641 ( .A(n26796), .B(n26798), .Z(n26829) );
  AND U31642 ( .A(n26830), .B(n26831), .Z(n26798) );
  NANDN U31643 ( .A(n26832), .B(n26833), .Z(n26831) );
  NANDN U31644 ( .A(n26834), .B(n26835), .Z(n26833) );
  IV U31645 ( .A(n26836), .Z(n26835) );
  NAND U31646 ( .A(n26836), .B(n26834), .Z(n26830) );
  AND U31647 ( .A(n26837), .B(n26838), .Z(n26796) );
  NAND U31648 ( .A(n26839), .B(n26840), .Z(n26838) );
  OR U31649 ( .A(n26841), .B(n26842), .Z(n26840) );
  NAND U31650 ( .A(n26842), .B(n26841), .Z(n26837) );
  IV U31651 ( .A(n26843), .Z(n26842) );
  NAND U31652 ( .A(n26844), .B(n26845), .Z(n26799) );
  NANDN U31653 ( .A(n26846), .B(n26847), .Z(n26845) );
  AND U31654 ( .A(n26848), .B(n26849), .Z(n26847) );
  NAND U31655 ( .A(n26850), .B(n26851), .Z(n26849) );
  OR U31656 ( .A(n26851), .B(n26850), .Z(n26844) );
  IV U31657 ( .A(n26852), .Z(n26850) );
  XOR U31658 ( .A(n26825), .B(n26853), .Z(N27942) );
  XNOR U31659 ( .A(n26828), .B(n26827), .Z(n26853) );
  XNOR U31660 ( .A(n26839), .B(n26854), .Z(n26827) );
  XOR U31661 ( .A(n26843), .B(n26841), .Z(n26854) );
  XNOR U31662 ( .A(n26855), .B(n26856), .Z(n26841) );
  XOR U31663 ( .A(n26851), .B(n26852), .Z(n26856) );
  NAND U31664 ( .A(n26857), .B(n26858), .Z(n26852) );
  NAND U31665 ( .A(n26859), .B(n26860), .Z(n26858) );
  NANDN U31666 ( .A(n26861), .B(n26862), .Z(n26857) );
  AND U31667 ( .A(n26863), .B(n26864), .Z(n26851) );
  NANDN U31668 ( .A(n26865), .B(n26866), .Z(n26864) );
  NAND U31669 ( .A(n26867), .B(n26868), .Z(n26863) );
  ANDN U31670 ( .B(n26848), .A(n26846), .Z(n26855) );
  NANDN U31671 ( .A(n26869), .B(n26870), .Z(n26843) );
  XNOR U31672 ( .A(n26834), .B(n26871), .Z(n26839) );
  XOR U31673 ( .A(n26832), .B(n26836), .Z(n26871) );
  NAND U31674 ( .A(n26872), .B(n26873), .Z(n26836) );
  NAND U31675 ( .A(n26874), .B(n26875), .Z(n26873) );
  NAND U31676 ( .A(n26876), .B(n26877), .Z(n26872) );
  AND U31677 ( .A(n26878), .B(n26879), .Z(n26832) );
  NAND U31678 ( .A(n26880), .B(n26881), .Z(n26879) );
  NAND U31679 ( .A(n26882), .B(n26883), .Z(n26878) );
  AND U31680 ( .A(n26884), .B(n26885), .Z(n26834) );
  NAND U31681 ( .A(n26886), .B(n26887), .Z(n26828) );
  XNOR U31682 ( .A(n26811), .B(n26888), .Z(n26825) );
  XOR U31683 ( .A(n26815), .B(n26813), .Z(n26888) );
  XOR U31684 ( .A(n26821), .B(n26889), .Z(n26813) );
  XOR U31685 ( .A(n26818), .B(n26822), .Z(n26889) );
  NAND U31686 ( .A(n26890), .B(n26891), .Z(n26822) );
  NAND U31687 ( .A(n26892), .B(n26893), .Z(n26891) );
  NAND U31688 ( .A(n26894), .B(n26895), .Z(n26890) );
  AND U31689 ( .A(n26896), .B(n26897), .Z(n26818) );
  NAND U31690 ( .A(n26898), .B(n26899), .Z(n26897) );
  NAND U31691 ( .A(n26900), .B(n26901), .Z(n26896) );
  NANDN U31692 ( .A(n26902), .B(n26903), .Z(n26821) );
  NANDN U31693 ( .A(n26904), .B(n26905), .Z(n26815) );
  XNOR U31694 ( .A(n26806), .B(n26906), .Z(n26811) );
  XOR U31695 ( .A(n26804), .B(n26808), .Z(n26906) );
  NAND U31696 ( .A(n26907), .B(n26908), .Z(n26808) );
  NAND U31697 ( .A(n26909), .B(n26910), .Z(n26908) );
  NAND U31698 ( .A(n26911), .B(n26912), .Z(n26907) );
  AND U31699 ( .A(n26913), .B(n26914), .Z(n26804) );
  NAND U31700 ( .A(n26915), .B(n26916), .Z(n26914) );
  NAND U31701 ( .A(n26917), .B(n26918), .Z(n26913) );
  AND U31702 ( .A(n26919), .B(n26920), .Z(n26806) );
  XOR U31703 ( .A(n26887), .B(n26886), .Z(N27941) );
  XNOR U31704 ( .A(n26905), .B(n26904), .Z(n26886) );
  XNOR U31705 ( .A(n26919), .B(n26920), .Z(n26904) );
  XOR U31706 ( .A(n26916), .B(n26915), .Z(n26920) );
  XOR U31707 ( .A(y[27]), .B(x[27]), .Z(n26915) );
  XOR U31708 ( .A(n26918), .B(n26917), .Z(n26916) );
  XOR U31709 ( .A(y[29]), .B(x[29]), .Z(n26917) );
  XOR U31710 ( .A(y[28]), .B(x[28]), .Z(n26918) );
  XOR U31711 ( .A(n26910), .B(n26909), .Z(n26919) );
  XOR U31712 ( .A(n26912), .B(n26911), .Z(n26909) );
  XOR U31713 ( .A(y[26]), .B(x[26]), .Z(n26911) );
  XOR U31714 ( .A(y[25]), .B(x[25]), .Z(n26912) );
  XOR U31715 ( .A(y[24]), .B(x[24]), .Z(n26910) );
  XNOR U31716 ( .A(n26903), .B(n26902), .Z(n26905) );
  XNOR U31717 ( .A(n26899), .B(n26898), .Z(n26902) );
  XOR U31718 ( .A(n26901), .B(n26900), .Z(n26898) );
  XOR U31719 ( .A(y[23]), .B(x[23]), .Z(n26900) );
  XOR U31720 ( .A(y[22]), .B(x[22]), .Z(n26901) );
  XOR U31721 ( .A(y[21]), .B(x[21]), .Z(n26899) );
  XOR U31722 ( .A(n26893), .B(n26892), .Z(n26903) );
  XOR U31723 ( .A(n26895), .B(n26894), .Z(n26892) );
  XOR U31724 ( .A(y[20]), .B(x[20]), .Z(n26894) );
  XOR U31725 ( .A(y[19]), .B(x[19]), .Z(n26895) );
  XOR U31726 ( .A(y[18]), .B(x[18]), .Z(n26893) );
  XNOR U31727 ( .A(n26870), .B(n26869), .Z(n26887) );
  XNOR U31728 ( .A(n26884), .B(n26885), .Z(n26869) );
  XOR U31729 ( .A(n26881), .B(n26880), .Z(n26885) );
  XOR U31730 ( .A(y[15]), .B(x[15]), .Z(n26880) );
  XOR U31731 ( .A(n26883), .B(n26882), .Z(n26881) );
  XOR U31732 ( .A(y[17]), .B(x[17]), .Z(n26882) );
  XOR U31733 ( .A(y[16]), .B(x[16]), .Z(n26883) );
  XOR U31734 ( .A(n26875), .B(n26874), .Z(n26884) );
  XOR U31735 ( .A(n26877), .B(n26876), .Z(n26874) );
  XOR U31736 ( .A(y[14]), .B(x[14]), .Z(n26876) );
  XOR U31737 ( .A(y[13]), .B(x[13]), .Z(n26877) );
  XOR U31738 ( .A(y[12]), .B(x[12]), .Z(n26875) );
  XNOR U31739 ( .A(n26848), .B(n26846), .Z(n26870) );
  XNOR U31740 ( .A(n26860), .B(n26859), .Z(n26846) );
  XNOR U31741 ( .A(n26862), .B(n26861), .Z(n26859) );
  XNOR U31742 ( .A(y[8]), .B(x[8]), .Z(n26861) );
  XOR U31743 ( .A(y[7]), .B(x[7]), .Z(n26862) );
  XOR U31744 ( .A(y[6]), .B(x[6]), .Z(n26860) );
  XNOR U31745 ( .A(n26866), .B(n26865), .Z(n26848) );
  XNOR U31746 ( .A(n26868), .B(n26867), .Z(n26865) );
  XOR U31747 ( .A(y[11]), .B(x[11]), .Z(n26867) );
  XOR U31748 ( .A(y[10]), .B(x[10]), .Z(n26868) );
  XOR U31749 ( .A(y[9]), .B(x[9]), .Z(n26866) );
  AND U31750 ( .A(n26921), .B(n26922), .Z(N27933) );
  XOR U31751 ( .A(n26922), .B(n26921), .Z(N27932) );
  AND U31752 ( .A(n26923), .B(n26924), .Z(n26921) );
  AND U31753 ( .A(n26925), .B(n26926), .Z(n26922) );
  NAND U31754 ( .A(n26927), .B(n26928), .Z(n26926) );
  NANDN U31755 ( .A(n26929), .B(n26930), .Z(n26928) );
  NANDN U31756 ( .A(n26930), .B(n26929), .Z(n26925) );
  XOR U31757 ( .A(n26930), .B(n26931), .Z(N27931) );
  XOR U31758 ( .A(n26927), .B(n26929), .Z(n26931) );
  AND U31759 ( .A(n26932), .B(n26933), .Z(n26929) );
  NANDN U31760 ( .A(n26934), .B(n26935), .Z(n26933) );
  NAND U31761 ( .A(n26936), .B(n26937), .Z(n26935) );
  OR U31762 ( .A(n26937), .B(n26936), .Z(n26932) );
  IV U31763 ( .A(n26938), .Z(n26936) );
  AND U31764 ( .A(n26939), .B(n26940), .Z(n26927) );
  NAND U31765 ( .A(n26941), .B(n26942), .Z(n26940) );
  NANDN U31766 ( .A(n26943), .B(n26944), .Z(n26942) );
  NANDN U31767 ( .A(n26944), .B(n26943), .Z(n26939) );
  XNOR U31768 ( .A(n26945), .B(n26923), .Z(n26930) );
  NAND U31769 ( .A(n26946), .B(n26947), .Z(n26923) );
  NANDN U31770 ( .A(n26948), .B(n26949), .Z(n26947) );
  NANDN U31771 ( .A(n26950), .B(n26951), .Z(n26946) );
  IV U31772 ( .A(n26924), .Z(n26945) );
  NAND U31773 ( .A(n26952), .B(n26953), .Z(n26924) );
  NANDN U31774 ( .A(n26954), .B(n26955), .Z(n26953) );
  NANDN U31775 ( .A(n26956), .B(n26957), .Z(n26955) );
  NANDN U31776 ( .A(n26957), .B(n26956), .Z(n26952) );
  XOR U31777 ( .A(n26941), .B(n26958), .Z(N27930) );
  XNOR U31778 ( .A(n26944), .B(n26943), .Z(n26958) );
  XOR U31779 ( .A(n26937), .B(n26959), .Z(n26943) );
  XOR U31780 ( .A(n26934), .B(n26938), .Z(n26959) );
  NAND U31781 ( .A(n26960), .B(n26961), .Z(n26938) );
  NAND U31782 ( .A(n26962), .B(n26963), .Z(n26961) );
  NAND U31783 ( .A(n26964), .B(n26965), .Z(n26960) );
  AND U31784 ( .A(n26966), .B(n26967), .Z(n26934) );
  NAND U31785 ( .A(n26968), .B(n26969), .Z(n26967) );
  NAND U31786 ( .A(n26970), .B(n26971), .Z(n26966) );
  NANDN U31787 ( .A(n26972), .B(n26973), .Z(n26937) );
  NAND U31788 ( .A(n26974), .B(n26975), .Z(n26944) );
  XNOR U31789 ( .A(n26954), .B(n26976), .Z(n26941) );
  XNOR U31790 ( .A(n26957), .B(n26956), .Z(n26976) );
  ANDN U31791 ( .B(n26977), .A(n26978), .Z(n26956) );
  AND U31792 ( .A(n26979), .B(n26980), .Z(n26957) );
  NAND U31793 ( .A(n26981), .B(n26982), .Z(n26980) );
  NAND U31794 ( .A(n26983), .B(n26984), .Z(n26979) );
  XOR U31795 ( .A(n26948), .B(n26949), .Z(n26954) );
  XNOR U31796 ( .A(n26950), .B(n26951), .Z(n26949) );
  NAND U31797 ( .A(n26985), .B(n26986), .Z(n26951) );
  NANDN U31798 ( .A(n26987), .B(n26988), .Z(n26986) );
  NANDN U31799 ( .A(n26989), .B(n26990), .Z(n26985) );
  AND U31800 ( .A(n26991), .B(n26992), .Z(n26950) );
  NAND U31801 ( .A(n26993), .B(n26994), .Z(n26992) );
  IV U31802 ( .A(n26995), .Z(n26993) );
  NANDN U31803 ( .A(n26996), .B(n26997), .Z(n26991) );
  AND U31804 ( .A(n26998), .B(n26999), .Z(n26948) );
  NAND U31805 ( .A(n27000), .B(n27001), .Z(n26999) );
  NAND U31806 ( .A(n27002), .B(n27003), .Z(n26998) );
  XOR U31807 ( .A(n26975), .B(n26974), .Z(N27929) );
  XNOR U31808 ( .A(n26977), .B(n26978), .Z(n26974) );
  XNOR U31809 ( .A(n27003), .B(n27002), .Z(n26978) );
  XOR U31810 ( .A(y[3999]), .B(x[3999]), .Z(n27002) );
  XOR U31811 ( .A(n27001), .B(n27000), .Z(n27003) );
  XNOR U31812 ( .A(n26994), .B(n26995), .Z(n27000) );
  XNOR U31813 ( .A(y[3]), .B(x[3]), .Z(n26995) );
  XNOR U31814 ( .A(n26997), .B(n26996), .Z(n26994) );
  XNOR U31815 ( .A(y[5]), .B(x[5]), .Z(n26996) );
  XOR U31816 ( .A(y[4]), .B(x[4]), .Z(n26997) );
  XNOR U31817 ( .A(n26988), .B(n26987), .Z(n27001) );
  XNOR U31818 ( .A(y[0]), .B(x[0]), .Z(n26987) );
  XNOR U31819 ( .A(n26990), .B(n26989), .Z(n26988) );
  XNOR U31820 ( .A(y[2]), .B(x[2]), .Z(n26989) );
  XOR U31821 ( .A(y[1]), .B(x[1]), .Z(n26990) );
  XOR U31822 ( .A(n26982), .B(n26981), .Z(n26977) );
  XOR U31823 ( .A(n26984), .B(n26983), .Z(n26981) );
  XOR U31824 ( .A(y[3998]), .B(x[3998]), .Z(n26983) );
  XOR U31825 ( .A(y[3997]), .B(x[3997]), .Z(n26984) );
  XOR U31826 ( .A(y[3996]), .B(x[3996]), .Z(n26982) );
  XNOR U31827 ( .A(n26973), .B(n26972), .Z(n26975) );
  XNOR U31828 ( .A(n26969), .B(n26968), .Z(n26972) );
  XOR U31829 ( .A(y[3993]), .B(x[3993]), .Z(n26968) );
  XOR U31830 ( .A(n26971), .B(n26970), .Z(n26969) );
  XOR U31831 ( .A(y[3995]), .B(x[3995]), .Z(n26970) );
  XOR U31832 ( .A(y[3994]), .B(x[3994]), .Z(n26971) );
  XOR U31833 ( .A(n26963), .B(n26962), .Z(n26973) );
  XOR U31834 ( .A(n26965), .B(n26964), .Z(n26962) );
  XOR U31835 ( .A(y[3992]), .B(x[3992]), .Z(n26964) );
  XOR U31836 ( .A(y[3991]), .B(x[3991]), .Z(n26965) );
  XOR U31837 ( .A(y[3990]), .B(x[3990]), .Z(n26963) );
endmodule

