
module stackMachine_N16 ( clk, rst, x, opcode, o );
  input [15:0] x;
  input [2:0] opcode;
  output [15:0] o;
  input clk, rst;
  wire   \stack[7][15] , \stack[7][14] , \stack[7][13] , \stack[7][12] ,
         \stack[7][11] , \stack[7][10] , \stack[7][9] , \stack[7][8] ,
         \stack[7][7] , \stack[7][6] , \stack[7][5] , \stack[7][4] ,
         \stack[7][3] , \stack[7][2] , \stack[7][1] , \stack[7][0] ,
         \stack[6][15] , \stack[6][14] , \stack[6][13] , \stack[6][12] ,
         \stack[6][11] , \stack[6][10] , \stack[6][9] , \stack[6][8] ,
         \stack[6][7] , \stack[6][6] , \stack[6][5] , \stack[6][4] ,
         \stack[6][3] , \stack[6][2] , \stack[6][1] , \stack[6][0] ,
         \stack[5][15] , \stack[5][14] , \stack[5][13] , \stack[5][12] ,
         \stack[5][11] , \stack[5][10] , \stack[5][9] , \stack[5][8] ,
         \stack[5][7] , \stack[5][6] , \stack[5][5] , \stack[5][4] ,
         \stack[5][3] , \stack[5][2] , \stack[5][1] , \stack[5][0] ,
         \stack[4][15] , \stack[4][14] , \stack[4][13] , \stack[4][12] ,
         \stack[4][11] , \stack[4][10] , \stack[4][9] , \stack[4][8] ,
         \stack[4][7] , \stack[4][6] , \stack[4][5] , \stack[4][4] ,
         \stack[4][3] , \stack[4][2] , \stack[4][1] , \stack[4][0] ,
         \stack[3][15] , \stack[3][14] , \stack[3][13] , \stack[3][12] ,
         \stack[3][11] , \stack[3][10] , \stack[3][9] , \stack[3][8] ,
         \stack[3][7] , \stack[3][6] , \stack[3][5] , \stack[3][4] ,
         \stack[3][3] , \stack[3][2] , \stack[3][1] , \stack[3][0] ,
         \stack[2][15] , \stack[2][14] , \stack[2][13] , \stack[2][12] ,
         \stack[2][11] , \stack[2][10] , \stack[2][9] , \stack[2][8] ,
         \stack[2][7] , \stack[2][6] , \stack[2][5] , \stack[2][4] ,
         \stack[2][3] , \stack[2][2] , \stack[2][1] , \stack[2][0] ,
         \stack[1][15] , \stack[1][14] , \stack[1][13] , \stack[1][12] ,
         \stack[1][11] , \stack[1][10] , \stack[1][9] , \stack[1][8] ,
         \stack[1][7] , \stack[1][6] , \stack[1][5] , \stack[1][4] ,
         \stack[1][3] , \stack[1][2] , \stack[1][1] , \stack[1][0] ,
         \C3/DATA5_0 , \C3/DATA5_2 , \C3/DATA5_3 , \C3/DATA5_4 , \C3/DATA5_5 ,
         \C3/DATA5_6 , \C3/DATA5_7 , \C3/DATA5_8 , \C3/DATA5_9 , \C3/DATA5_10 ,
         \C3/DATA5_11 , \C3/DATA5_12 , \C3/DATA5_13 , \C3/DATA5_14 ,
         \C3/DATA5_15 , n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, \C1/Z_0 ,
         \U1/RSOP_16/C3/Z_15 , \U1/RSOP_16/C3/Z_14 , \U1/RSOP_16/C3/Z_13 ,
         \U1/RSOP_16/C3/Z_12 , \U1/RSOP_16/C3/Z_11 , \U1/RSOP_16/C3/Z_10 ,
         \U1/RSOP_16/C3/Z_9 , \U1/RSOP_16/C3/Z_8 , \U1/RSOP_16/C3/Z_7 ,
         \U1/RSOP_16/C3/Z_6 , \U1/RSOP_16/C3/Z_5 , \U1/RSOP_16/C3/Z_4 ,
         \U1/RSOP_16/C3/Z_3 , \U1/RSOP_16/C3/Z_2 , \U1/RSOP_16/C3/Z_1 ,
         \U1/RSOP_16/C3/Z_0 , \U1/RSOP_16/C2/Z_15 , \U1/RSOP_16/C2/Z_14 ,
         \U1/RSOP_16/C2/Z_13 , \U1/RSOP_16/C2/Z_12 , \U1/RSOP_16/C2/Z_11 ,
         \U1/RSOP_16/C2/Z_10 , \U1/RSOP_16/C2/Z_9 , \U1/RSOP_16/C2/Z_8 ,
         \U1/RSOP_16/C2/Z_7 , \U1/RSOP_16/C2/Z_6 , \U1/RSOP_16/C2/Z_5 ,
         \U1/RSOP_16/C2/Z_4 , \U1/RSOP_16/C2/Z_3 , \U1/RSOP_16/C2/Z_2 ,
         \U1/RSOP_16/C2/Z_1 , \U1/RSOP_16/C2/Z_0 , \DP_OP_25_64_3291/n169 ,
         \DP_OP_25_64_3291/n168 , \DP_OP_25_64_3291/n167 ,
         \DP_OP_25_64_3291/n166 , \DP_OP_25_64_3291/n165 ,
         \DP_OP_25_64_3291/n164 , \DP_OP_25_64_3291/n163 ,
         \DP_OP_25_64_3291/n162 , \DP_OP_25_64_3291/n161 ,
         \DP_OP_25_64_3291/n160 , \DP_OP_25_64_3291/n159 ,
         \DP_OP_25_64_3291/n158 , \DP_OP_25_64_3291/n157 ,
         \DP_OP_25_64_3291/n156 , \DP_OP_25_64_3291/n155 ,
         \DP_OP_25_64_3291/n154 , \DP_OP_25_64_3291/n149 ,
         \DP_OP_25_64_3291/n148 , \DP_OP_25_64_3291/n147 ,
         \DP_OP_25_64_3291/n146 , \DP_OP_25_64_3291/n145 ,
         \DP_OP_25_64_3291/n144 , \DP_OP_25_64_3291/n143 ,
         \DP_OP_25_64_3291/n142 , \DP_OP_25_64_3291/n141 ,
         \DP_OP_25_64_3291/n140 , \DP_OP_25_64_3291/n139 ,
         \DP_OP_25_64_3291/n138 , \DP_OP_25_64_3291/n137 ,
         \DP_OP_25_64_3291/n136 , \DP_OP_25_64_3291/n135 ,
         \DP_OP_25_64_3291/n134 , \DP_OP_25_64_3291/n133 ,
         \DP_OP_25_64_3291/n132 , \DP_OP_25_64_3291/n131 ,
         \DP_OP_25_64_3291/n130 , \DP_OP_25_64_3291/n129 ,
         \DP_OP_25_64_3291/n128 , \DP_OP_25_64_3291/n127 ,
         \DP_OP_25_64_3291/n126 , \DP_OP_25_64_3291/n125 ,
         \DP_OP_25_64_3291/n124 , \DP_OP_25_64_3291/n123 ,
         \DP_OP_25_64_3291/n122 , \DP_OP_25_64_3291/n121 ,
         \DP_OP_25_64_3291/n120 , \DP_OP_25_64_3291/n119 ,
         \DP_OP_25_64_3291/n117 , \DP_OP_25_64_3291/n116 ,
         \DP_OP_25_64_3291/n110 , \DP_OP_25_64_3291/n109 ,
         \DP_OP_25_64_3291/n103 , \DP_OP_25_64_3291/n102 ,
         \DP_OP_25_64_3291/n96 , \DP_OP_25_64_3291/n95 ,
         \DP_OP_25_64_3291/n89 , \DP_OP_25_64_3291/n88 ,
         \DP_OP_25_64_3291/n82 , \DP_OP_25_64_3291/n81 ,
         \DP_OP_25_64_3291/n70 , \DP_OP_25_64_3291/n69 ,
         \DP_OP_25_64_3291/n57 , \DP_OP_25_64_3291/n56 ,
         \DP_OP_25_64_3291/n50 , \DP_OP_25_64_3291/n49 ,
         \DP_OP_25_64_3291/n43 , \DP_OP_25_64_3291/n42 ,
         \DP_OP_25_64_3291/n36 , \DP_OP_25_64_3291/n35 ,
         \DP_OP_25_64_3291/n29 , \DP_OP_25_64_3291/n28 ,
         \DP_OP_25_64_3291/n22 , \DP_OP_25_64_3291/n21 ,
         \DP_OP_25_64_3291/n15 , \DP_OP_25_64_3291/n14 , \DP_OP_25_64_3291/n8 ,
         \DP_OP_25_64_3291/n5 , n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101;

  DFF \stack_reg[0][0]  ( .D(n649), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \stack_reg[1][0]  ( .D(n648), .CLK(clk), .RST(rst), .Q(\stack[1][0] ) );
  DFF \stack_reg[0][1]  ( .D(n647), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \stack_reg[1][1]  ( .D(n646), .CLK(clk), .RST(rst), .Q(\stack[1][1] ) );
  DFF \stack_reg[2][1]  ( .D(n645), .CLK(clk), .RST(rst), .Q(\stack[2][1] ) );
  DFF \stack_reg[3][1]  ( .D(n644), .CLK(clk), .RST(rst), .Q(\stack[3][1] ) );
  DFF \stack_reg[4][1]  ( .D(n643), .CLK(clk), .RST(rst), .Q(\stack[4][1] ) );
  DFF \stack_reg[5][1]  ( .D(n642), .CLK(clk), .RST(rst), .Q(\stack[5][1] ) );
  DFF \stack_reg[6][1]  ( .D(n641), .CLK(clk), .RST(rst), .Q(\stack[6][1] ) );
  DFF \stack_reg[7][1]  ( .D(n640), .CLK(clk), .RST(rst), .Q(\stack[7][1] ) );
  DFF \stack_reg[0][2]  ( .D(n639), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \stack_reg[1][2]  ( .D(n638), .CLK(clk), .RST(rst), .Q(\stack[1][2] ) );
  DFF \stack_reg[2][2]  ( .D(n637), .CLK(clk), .RST(rst), .Q(\stack[2][2] ) );
  DFF \stack_reg[3][2]  ( .D(n636), .CLK(clk), .RST(rst), .Q(\stack[3][2] ) );
  DFF \stack_reg[4][2]  ( .D(n635), .CLK(clk), .RST(rst), .Q(\stack[4][2] ) );
  DFF \stack_reg[5][2]  ( .D(n634), .CLK(clk), .RST(rst), .Q(\stack[5][2] ) );
  DFF \stack_reg[6][2]  ( .D(n633), .CLK(clk), .RST(rst), .Q(\stack[6][2] ) );
  DFF \stack_reg[7][2]  ( .D(n632), .CLK(clk), .RST(rst), .Q(\stack[7][2] ) );
  DFF \stack_reg[0][3]  ( .D(n631), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \stack_reg[1][3]  ( .D(n630), .CLK(clk), .RST(rst), .Q(\stack[1][3] ) );
  DFF \stack_reg[2][3]  ( .D(n629), .CLK(clk), .RST(rst), .Q(\stack[2][3] ) );
  DFF \stack_reg[3][3]  ( .D(n628), .CLK(clk), .RST(rst), .Q(\stack[3][3] ) );
  DFF \stack_reg[4][3]  ( .D(n627), .CLK(clk), .RST(rst), .Q(\stack[4][3] ) );
  DFF \stack_reg[5][3]  ( .D(n626), .CLK(clk), .RST(rst), .Q(\stack[5][3] ) );
  DFF \stack_reg[6][3]  ( .D(n625), .CLK(clk), .RST(rst), .Q(\stack[6][3] ) );
  DFF \stack_reg[7][3]  ( .D(n624), .CLK(clk), .RST(rst), .Q(\stack[7][3] ) );
  DFF \stack_reg[0][4]  ( .D(n623), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \stack_reg[1][4]  ( .D(n622), .CLK(clk), .RST(rst), .Q(\stack[1][4] ) );
  DFF \stack_reg[2][4]  ( .D(n621), .CLK(clk), .RST(rst), .Q(\stack[2][4] ) );
  DFF \stack_reg[3][4]  ( .D(n620), .CLK(clk), .RST(rst), .Q(\stack[3][4] ) );
  DFF \stack_reg[4][4]  ( .D(n619), .CLK(clk), .RST(rst), .Q(\stack[4][4] ) );
  DFF \stack_reg[5][4]  ( .D(n618), .CLK(clk), .RST(rst), .Q(\stack[5][4] ) );
  DFF \stack_reg[6][4]  ( .D(n617), .CLK(clk), .RST(rst), .Q(\stack[6][4] ) );
  DFF \stack_reg[7][4]  ( .D(n616), .CLK(clk), .RST(rst), .Q(\stack[7][4] ) );
  DFF \stack_reg[0][5]  ( .D(n615), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \stack_reg[1][5]  ( .D(n614), .CLK(clk), .RST(rst), .Q(\stack[1][5] ) );
  DFF \stack_reg[2][5]  ( .D(n613), .CLK(clk), .RST(rst), .Q(\stack[2][5] ) );
  DFF \stack_reg[3][5]  ( .D(n612), .CLK(clk), .RST(rst), .Q(\stack[3][5] ) );
  DFF \stack_reg[4][5]  ( .D(n611), .CLK(clk), .RST(rst), .Q(\stack[4][5] ) );
  DFF \stack_reg[5][5]  ( .D(n610), .CLK(clk), .RST(rst), .Q(\stack[5][5] ) );
  DFF \stack_reg[6][5]  ( .D(n609), .CLK(clk), .RST(rst), .Q(\stack[6][5] ) );
  DFF \stack_reg[7][5]  ( .D(n608), .CLK(clk), .RST(rst), .Q(\stack[7][5] ) );
  DFF \stack_reg[0][6]  ( .D(n607), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \stack_reg[1][6]  ( .D(n606), .CLK(clk), .RST(rst), .Q(\stack[1][6] ) );
  DFF \stack_reg[2][6]  ( .D(n605), .CLK(clk), .RST(rst), .Q(\stack[2][6] ) );
  DFF \stack_reg[3][6]  ( .D(n604), .CLK(clk), .RST(rst), .Q(\stack[3][6] ) );
  DFF \stack_reg[4][6]  ( .D(n603), .CLK(clk), .RST(rst), .Q(\stack[4][6] ) );
  DFF \stack_reg[5][6]  ( .D(n602), .CLK(clk), .RST(rst), .Q(\stack[5][6] ) );
  DFF \stack_reg[6][6]  ( .D(n601), .CLK(clk), .RST(rst), .Q(\stack[6][6] ) );
  DFF \stack_reg[7][6]  ( .D(n600), .CLK(clk), .RST(rst), .Q(\stack[7][6] ) );
  DFF \stack_reg[0][7]  ( .D(n599), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \stack_reg[1][7]  ( .D(n598), .CLK(clk), .RST(rst), .Q(\stack[1][7] ) );
  DFF \stack_reg[2][7]  ( .D(n597), .CLK(clk), .RST(rst), .Q(\stack[2][7] ) );
  DFF \stack_reg[3][7]  ( .D(n596), .CLK(clk), .RST(rst), .Q(\stack[3][7] ) );
  DFF \stack_reg[4][7]  ( .D(n595), .CLK(clk), .RST(rst), .Q(\stack[4][7] ) );
  DFF \stack_reg[5][7]  ( .D(n594), .CLK(clk), .RST(rst), .Q(\stack[5][7] ) );
  DFF \stack_reg[6][7]  ( .D(n593), .CLK(clk), .RST(rst), .Q(\stack[6][7] ) );
  DFF \stack_reg[7][7]  ( .D(n592), .CLK(clk), .RST(rst), .Q(\stack[7][7] ) );
  DFF \stack_reg[0][8]  ( .D(n591), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \stack_reg[1][8]  ( .D(n590), .CLK(clk), .RST(rst), .Q(\stack[1][8] ) );
  DFF \stack_reg[2][8]  ( .D(n589), .CLK(clk), .RST(rst), .Q(\stack[2][8] ) );
  DFF \stack_reg[3][8]  ( .D(n588), .CLK(clk), .RST(rst), .Q(\stack[3][8] ) );
  DFF \stack_reg[4][8]  ( .D(n587), .CLK(clk), .RST(rst), .Q(\stack[4][8] ) );
  DFF \stack_reg[5][8]  ( .D(n586), .CLK(clk), .RST(rst), .Q(\stack[5][8] ) );
  DFF \stack_reg[6][8]  ( .D(n585), .CLK(clk), .RST(rst), .Q(\stack[6][8] ) );
  DFF \stack_reg[7][8]  ( .D(n584), .CLK(clk), .RST(rst), .Q(\stack[7][8] ) );
  DFF \stack_reg[0][9]  ( .D(n583), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \stack_reg[1][9]  ( .D(n582), .CLK(clk), .RST(rst), .Q(\stack[1][9] ) );
  DFF \stack_reg[2][9]  ( .D(n581), .CLK(clk), .RST(rst), .Q(\stack[2][9] ) );
  DFF \stack_reg[3][9]  ( .D(n580), .CLK(clk), .RST(rst), .Q(\stack[3][9] ) );
  DFF \stack_reg[4][9]  ( .D(n579), .CLK(clk), .RST(rst), .Q(\stack[4][9] ) );
  DFF \stack_reg[5][9]  ( .D(n578), .CLK(clk), .RST(rst), .Q(\stack[5][9] ) );
  DFF \stack_reg[6][9]  ( .D(n577), .CLK(clk), .RST(rst), .Q(\stack[6][9] ) );
  DFF \stack_reg[7][9]  ( .D(n576), .CLK(clk), .RST(rst), .Q(\stack[7][9] ) );
  DFF \stack_reg[0][10]  ( .D(n575), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \stack_reg[1][10]  ( .D(n574), .CLK(clk), .RST(rst), .Q(\stack[1][10] )
         );
  DFF \stack_reg[2][10]  ( .D(n573), .CLK(clk), .RST(rst), .Q(\stack[2][10] )
         );
  DFF \stack_reg[3][10]  ( .D(n572), .CLK(clk), .RST(rst), .Q(\stack[3][10] )
         );
  DFF \stack_reg[4][10]  ( .D(n571), .CLK(clk), .RST(rst), .Q(\stack[4][10] )
         );
  DFF \stack_reg[5][10]  ( .D(n570), .CLK(clk), .RST(rst), .Q(\stack[5][10] )
         );
  DFF \stack_reg[6][10]  ( .D(n569), .CLK(clk), .RST(rst), .Q(\stack[6][10] )
         );
  DFF \stack_reg[7][10]  ( .D(n568), .CLK(clk), .RST(rst), .Q(\stack[7][10] )
         );
  DFF \stack_reg[0][11]  ( .D(n567), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \stack_reg[1][11]  ( .D(n566), .CLK(clk), .RST(rst), .Q(\stack[1][11] )
         );
  DFF \stack_reg[2][11]  ( .D(n565), .CLK(clk), .RST(rst), .Q(\stack[2][11] )
         );
  DFF \stack_reg[3][11]  ( .D(n564), .CLK(clk), .RST(rst), .Q(\stack[3][11] )
         );
  DFF \stack_reg[4][11]  ( .D(n563), .CLK(clk), .RST(rst), .Q(\stack[4][11] )
         );
  DFF \stack_reg[5][11]  ( .D(n562), .CLK(clk), .RST(rst), .Q(\stack[5][11] )
         );
  DFF \stack_reg[6][11]  ( .D(n561), .CLK(clk), .RST(rst), .Q(\stack[6][11] )
         );
  DFF \stack_reg[7][11]  ( .D(n560), .CLK(clk), .RST(rst), .Q(\stack[7][11] )
         );
  DFF \stack_reg[0][12]  ( .D(n559), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \stack_reg[1][12]  ( .D(n558), .CLK(clk), .RST(rst), .Q(\stack[1][12] )
         );
  DFF \stack_reg[2][12]  ( .D(n557), .CLK(clk), .RST(rst), .Q(\stack[2][12] )
         );
  DFF \stack_reg[3][12]  ( .D(n556), .CLK(clk), .RST(rst), .Q(\stack[3][12] )
         );
  DFF \stack_reg[4][12]  ( .D(n555), .CLK(clk), .RST(rst), .Q(\stack[4][12] )
         );
  DFF \stack_reg[5][12]  ( .D(n554), .CLK(clk), .RST(rst), .Q(\stack[5][12] )
         );
  DFF \stack_reg[6][12]  ( .D(n553), .CLK(clk), .RST(rst), .Q(\stack[6][12] )
         );
  DFF \stack_reg[7][12]  ( .D(n552), .CLK(clk), .RST(rst), .Q(\stack[7][12] )
         );
  DFF \stack_reg[0][13]  ( .D(n551), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \stack_reg[1][13]  ( .D(n550), .CLK(clk), .RST(rst), .Q(\stack[1][13] )
         );
  DFF \stack_reg[2][13]  ( .D(n549), .CLK(clk), .RST(rst), .Q(\stack[2][13] )
         );
  DFF \stack_reg[3][13]  ( .D(n548), .CLK(clk), .RST(rst), .Q(\stack[3][13] )
         );
  DFF \stack_reg[4][13]  ( .D(n547), .CLK(clk), .RST(rst), .Q(\stack[4][13] )
         );
  DFF \stack_reg[5][13]  ( .D(n546), .CLK(clk), .RST(rst), .Q(\stack[5][13] )
         );
  DFF \stack_reg[6][13]  ( .D(n545), .CLK(clk), .RST(rst), .Q(\stack[6][13] )
         );
  DFF \stack_reg[7][13]  ( .D(n544), .CLK(clk), .RST(rst), .Q(\stack[7][13] )
         );
  DFF \stack_reg[0][14]  ( .D(n543), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \stack_reg[1][14]  ( .D(n542), .CLK(clk), .RST(rst), .Q(\stack[1][14] )
         );
  DFF \stack_reg[2][14]  ( .D(n541), .CLK(clk), .RST(rst), .Q(\stack[2][14] )
         );
  DFF \stack_reg[3][14]  ( .D(n540), .CLK(clk), .RST(rst), .Q(\stack[3][14] )
         );
  DFF \stack_reg[4][14]  ( .D(n539), .CLK(clk), .RST(rst), .Q(\stack[4][14] )
         );
  DFF \stack_reg[5][14]  ( .D(n538), .CLK(clk), .RST(rst), .Q(\stack[5][14] )
         );
  DFF \stack_reg[6][14]  ( .D(n537), .CLK(clk), .RST(rst), .Q(\stack[6][14] )
         );
  DFF \stack_reg[7][14]  ( .D(n536), .CLK(clk), .RST(rst), .Q(\stack[7][14] )
         );
  DFF \stack_reg[0][15]  ( .D(n535), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \stack_reg[1][15]  ( .D(n534), .CLK(clk), .RST(rst), .Q(\stack[1][15] )
         );
  DFF \stack_reg[2][15]  ( .D(n533), .CLK(clk), .RST(rst), .Q(\stack[2][15] )
         );
  DFF \stack_reg[3][15]  ( .D(n532), .CLK(clk), .RST(rst), .Q(\stack[3][15] )
         );
  DFF \stack_reg[4][15]  ( .D(n531), .CLK(clk), .RST(rst), .Q(\stack[4][15] )
         );
  DFF \stack_reg[5][15]  ( .D(n530), .CLK(clk), .RST(rst), .Q(\stack[5][15] )
         );
  DFF \stack_reg[6][15]  ( .D(n529), .CLK(clk), .RST(rst), .Q(\stack[6][15] )
         );
  DFF \stack_reg[7][15]  ( .D(n528), .CLK(clk), .RST(rst), .Q(\stack[7][15] )
         );
  DFF \stack_reg[2][0]  ( .D(n527), .CLK(clk), .RST(rst), .Q(\stack[2][0] ) );
  DFF \stack_reg[3][0]  ( .D(n526), .CLK(clk), .RST(rst), .Q(\stack[3][0] ) );
  DFF \stack_reg[4][0]  ( .D(n525), .CLK(clk), .RST(rst), .Q(\stack[4][0] ) );
  DFF \stack_reg[5][0]  ( .D(n524), .CLK(clk), .RST(rst), .Q(\stack[5][0] ) );
  DFF \stack_reg[6][0]  ( .D(n523), .CLK(clk), .RST(rst), .Q(\stack[6][0] ) );
  DFF \stack_reg[7][0]  ( .D(n522), .CLK(clk), .RST(rst), .Q(\stack[7][0] ) );
  XOR \DP_OP_25_64_3291/U80  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_0 ), .Z(
        \DP_OP_25_64_3291/n169 ) );
  XOR \DP_OP_25_64_3291/U79  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_1 ), .Z(
        \DP_OP_25_64_3291/n168 ) );
  XOR \DP_OP_25_64_3291/U78  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_2 ), .Z(
        \DP_OP_25_64_3291/n167 ) );
  XOR \DP_OP_25_64_3291/U77  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_3 ), .Z(
        \DP_OP_25_64_3291/n166 ) );
  XOR \DP_OP_25_64_3291/U76  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_4 ), .Z(
        \DP_OP_25_64_3291/n165 ) );
  XOR \DP_OP_25_64_3291/U75  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_5 ), .Z(
        \DP_OP_25_64_3291/n164 ) );
  XOR \DP_OP_25_64_3291/U74  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_6 ), .Z(
        \DP_OP_25_64_3291/n163 ) );
  XOR \DP_OP_25_64_3291/U73  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_7 ), .Z(
        \DP_OP_25_64_3291/n162 ) );
  XOR \DP_OP_25_64_3291/U72  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_8 ), .Z(
        \DP_OP_25_64_3291/n161 ) );
  XOR \DP_OP_25_64_3291/U71  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_9 ), .Z(
        \DP_OP_25_64_3291/n160 ) );
  XOR \DP_OP_25_64_3291/U70  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_10 ), .Z(
        \DP_OP_25_64_3291/n159 ) );
  XOR \DP_OP_25_64_3291/U69  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_11 ), .Z(
        \DP_OP_25_64_3291/n158 ) );
  XOR \DP_OP_25_64_3291/U68  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_12 ), .Z(
        \DP_OP_25_64_3291/n157 ) );
  XOR \DP_OP_25_64_3291/U67  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_13 ), .Z(
        \DP_OP_25_64_3291/n156 ) );
  XOR \DP_OP_25_64_3291/U66  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_14 ), .Z(
        \DP_OP_25_64_3291/n155 ) );
  XOR \DP_OP_25_64_3291/U65  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_15 ), .Z(
        \DP_OP_25_64_3291/n154 ) );
  XOR \DP_OP_25_64_3291/U62  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_3291/n134 ) );
  XOR \DP_OP_25_64_3291/U61  ( .A(\DP_OP_25_64_3291/n134 ), .B(
        \DP_OP_25_64_3291/n169 ), .Z(\C3/DATA5_0 ) );
  XOR \DP_OP_25_64_3291/U60  ( .A(\DP_OP_25_64_3291/n168 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_3291/n133 ) );
  XOR \DP_OP_25_64_3291/U58  ( .A(\DP_OP_25_64_3291/n167 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_3291/n132 ) );
  XOR \DP_OP_25_64_3291/U57  ( .A(\DP_OP_25_64_3291/n148 ), .B(
        \DP_OP_25_64_3291/n132 ), .Z(\C3/DATA5_2 ) );
  XOR \DP_OP_25_64_3291/U56  ( .A(\DP_OP_25_64_3291/n166 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_3291/n131 ) );
  XOR \DP_OP_25_64_3291/U55  ( .A(\DP_OP_25_64_3291/n147 ), .B(
        \DP_OP_25_64_3291/n131 ), .Z(\C3/DATA5_3 ) );
  XOR \DP_OP_25_64_3291/U54  ( .A(\DP_OP_25_64_3291/n165 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_3291/n130 ) );
  XOR \DP_OP_25_64_3291/U53  ( .A(\DP_OP_25_64_3291/n146 ), .B(
        \DP_OP_25_64_3291/n130 ), .Z(\C3/DATA5_4 ) );
  XOR \DP_OP_25_64_3291/U52  ( .A(\DP_OP_25_64_3291/n164 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_3291/n129 ) );
  XOR \DP_OP_25_64_3291/U51  ( .A(\DP_OP_25_64_3291/n145 ), .B(
        \DP_OP_25_64_3291/n129 ), .Z(\C3/DATA5_5 ) );
  XOR \DP_OP_25_64_3291/U50  ( .A(\DP_OP_25_64_3291/n163 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_3291/n128 ) );
  XOR \DP_OP_25_64_3291/U49  ( .A(\DP_OP_25_64_3291/n144 ), .B(
        \DP_OP_25_64_3291/n128 ), .Z(\C3/DATA5_6 ) );
  XOR \DP_OP_25_64_3291/U48  ( .A(\DP_OP_25_64_3291/n162 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_3291/n127 ) );
  XOR \DP_OP_25_64_3291/U47  ( .A(\DP_OP_25_64_3291/n143 ), .B(
        \DP_OP_25_64_3291/n127 ), .Z(\C3/DATA5_7 ) );
  XOR \DP_OP_25_64_3291/U46  ( .A(\DP_OP_25_64_3291/n161 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_3291/n126 ) );
  XOR \DP_OP_25_64_3291/U45  ( .A(\DP_OP_25_64_3291/n142 ), .B(
        \DP_OP_25_64_3291/n126 ), .Z(\C3/DATA5_8 ) );
  XOR \DP_OP_25_64_3291/U44  ( .A(\DP_OP_25_64_3291/n160 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_3291/n125 ) );
  XOR \DP_OP_25_64_3291/U43  ( .A(\DP_OP_25_64_3291/n141 ), .B(
        \DP_OP_25_64_3291/n125 ), .Z(\C3/DATA5_9 ) );
  XOR \DP_OP_25_64_3291/U42  ( .A(\DP_OP_25_64_3291/n159 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_3291/n124 ) );
  XOR \DP_OP_25_64_3291/U41  ( .A(\DP_OP_25_64_3291/n140 ), .B(
        \DP_OP_25_64_3291/n124 ), .Z(\C3/DATA5_10 ) );
  XOR \DP_OP_25_64_3291/U40  ( .A(\DP_OP_25_64_3291/n158 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_3291/n123 ) );
  XOR \DP_OP_25_64_3291/U30  ( .A(\DP_OP_25_64_3291/n139 ), .B(
        \DP_OP_25_64_3291/n123 ), .Z(\C3/DATA5_11 ) );
  XOR \DP_OP_25_64_3291/U20  ( .A(\DP_OP_25_64_3291/n157 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_3291/n122 ) );
  XOR \DP_OP_25_64_3291/U10  ( .A(\DP_OP_25_64_3291/n138 ), .B(
        \DP_OP_25_64_3291/n122 ), .Z(\C3/DATA5_12 ) );
  XOR \DP_OP_25_64_3291/U9  ( .A(\DP_OP_25_64_3291/n156 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_3291/n121 ) );
  XOR \DP_OP_25_64_3291/U8  ( .A(\DP_OP_25_64_3291/n137 ), .B(
        \DP_OP_25_64_3291/n121 ), .Z(\C3/DATA5_13 ) );
  XOR \DP_OP_25_64_3291/U7  ( .A(\DP_OP_25_64_3291/n155 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_3291/n120 ) );
  XOR \DP_OP_25_64_3291/U6  ( .A(\DP_OP_25_64_3291/n136 ), .B(
        \DP_OP_25_64_3291/n120 ), .Z(\C3/DATA5_14 ) );
  XOR \DP_OP_25_64_3291/U5  ( .A(\DP_OP_25_64_3291/n154 ), .B(
        \U1/RSOP_16/C2/Z_15 ), .Z(\DP_OP_25_64_3291/n119 ) );
  XOR \DP_OP_25_64_3291/U4  ( .A(\DP_OP_25_64_3291/n135 ), .B(
        \DP_OP_25_64_3291/n119 ), .Z(\C3/DATA5_15 ) );
  NAND \DP_OP_25_64_3291/U114  ( .A(\DP_OP_25_64_3291/n155 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_3291/n5 ) );
  NAND \DP_OP_25_64_3291/U214  ( .A(\DP_OP_25_64_3291/n136 ), .B(
        \DP_OP_25_64_3291/n120 ), .Z(\DP_OP_25_64_3291/n8 ) );
  NAND \DP_OP_25_64_3291/U314  ( .A(\DP_OP_25_64_3291/n5 ), .B(
        \DP_OP_25_64_3291/n8 ), .Z(\DP_OP_25_64_3291/n135 ) );
  NAND \DP_OP_25_64_3291/U113  ( .A(\DP_OP_25_64_3291/n156 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_3291/n14 ) );
  NAND \DP_OP_25_64_3291/U213  ( .A(\DP_OP_25_64_3291/n137 ), .B(
        \DP_OP_25_64_3291/n121 ), .Z(\DP_OP_25_64_3291/n15 ) );
  NAND \DP_OP_25_64_3291/U313  ( .A(\DP_OP_25_64_3291/n14 ), .B(
        \DP_OP_25_64_3291/n15 ), .Z(\DP_OP_25_64_3291/n136 ) );
  NAND \DP_OP_25_64_3291/U112  ( .A(\DP_OP_25_64_3291/n157 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_3291/n21 ) );
  NAND \DP_OP_25_64_3291/U212  ( .A(\DP_OP_25_64_3291/n138 ), .B(
        \DP_OP_25_64_3291/n122 ), .Z(\DP_OP_25_64_3291/n22 ) );
  NAND \DP_OP_25_64_3291/U312  ( .A(\DP_OP_25_64_3291/n21 ), .B(
        \DP_OP_25_64_3291/n22 ), .Z(\DP_OP_25_64_3291/n137 ) );
  NAND \DP_OP_25_64_3291/U111  ( .A(\DP_OP_25_64_3291/n158 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_3291/n28 ) );
  NAND \DP_OP_25_64_3291/U211  ( .A(\DP_OP_25_64_3291/n139 ), .B(
        \DP_OP_25_64_3291/n123 ), .Z(\DP_OP_25_64_3291/n29 ) );
  NAND \DP_OP_25_64_3291/U311  ( .A(\DP_OP_25_64_3291/n28 ), .B(
        \DP_OP_25_64_3291/n29 ), .Z(\DP_OP_25_64_3291/n138 ) );
  NAND \DP_OP_25_64_3291/U110  ( .A(\DP_OP_25_64_3291/n159 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_3291/n35 ) );
  NAND \DP_OP_25_64_3291/U210  ( .A(\DP_OP_25_64_3291/n140 ), .B(
        \DP_OP_25_64_3291/n124 ), .Z(\DP_OP_25_64_3291/n36 ) );
  NAND \DP_OP_25_64_3291/U310  ( .A(\DP_OP_25_64_3291/n35 ), .B(
        \DP_OP_25_64_3291/n36 ), .Z(\DP_OP_25_64_3291/n139 ) );
  NAND \DP_OP_25_64_3291/U19  ( .A(\DP_OP_25_64_3291/n160 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_3291/n42 ) );
  NAND \DP_OP_25_64_3291/U29  ( .A(\DP_OP_25_64_3291/n141 ), .B(
        \DP_OP_25_64_3291/n125 ), .Z(\DP_OP_25_64_3291/n43 ) );
  NAND \DP_OP_25_64_3291/U39  ( .A(\DP_OP_25_64_3291/n42 ), .B(
        \DP_OP_25_64_3291/n43 ), .Z(\DP_OP_25_64_3291/n140 ) );
  NAND \DP_OP_25_64_3291/U18  ( .A(\DP_OP_25_64_3291/n161 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_3291/n49 ) );
  NAND \DP_OP_25_64_3291/U28  ( .A(\DP_OP_25_64_3291/n142 ), .B(
        \DP_OP_25_64_3291/n126 ), .Z(\DP_OP_25_64_3291/n50 ) );
  NAND \DP_OP_25_64_3291/U38  ( .A(\DP_OP_25_64_3291/n49 ), .B(
        \DP_OP_25_64_3291/n50 ), .Z(\DP_OP_25_64_3291/n141 ) );
  NAND \DP_OP_25_64_3291/U17  ( .A(\DP_OP_25_64_3291/n162 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_3291/n56 ) );
  NAND \DP_OP_25_64_3291/U27  ( .A(\DP_OP_25_64_3291/n143 ), .B(
        \DP_OP_25_64_3291/n127 ), .Z(\DP_OP_25_64_3291/n57 ) );
  NAND \DP_OP_25_64_3291/U37  ( .A(\DP_OP_25_64_3291/n56 ), .B(
        \DP_OP_25_64_3291/n57 ), .Z(\DP_OP_25_64_3291/n142 ) );
  NAND \DP_OP_25_64_3291/U16  ( .A(\DP_OP_25_64_3291/n163 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_3291/n69 ) );
  NAND \DP_OP_25_64_3291/U26  ( .A(\DP_OP_25_64_3291/n144 ), .B(
        \DP_OP_25_64_3291/n128 ), .Z(\DP_OP_25_64_3291/n70 ) );
  NAND \DP_OP_25_64_3291/U36  ( .A(\DP_OP_25_64_3291/n69 ), .B(
        \DP_OP_25_64_3291/n70 ), .Z(\DP_OP_25_64_3291/n143 ) );
  NAND \DP_OP_25_64_3291/U15  ( .A(\DP_OP_25_64_3291/n164 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_3291/n81 ) );
  NAND \DP_OP_25_64_3291/U25  ( .A(\DP_OP_25_64_3291/n145 ), .B(
        \DP_OP_25_64_3291/n129 ), .Z(\DP_OP_25_64_3291/n82 ) );
  NAND \DP_OP_25_64_3291/U35  ( .A(\DP_OP_25_64_3291/n81 ), .B(
        \DP_OP_25_64_3291/n82 ), .Z(\DP_OP_25_64_3291/n144 ) );
  NAND \DP_OP_25_64_3291/U14  ( .A(\DP_OP_25_64_3291/n165 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_3291/n88 ) );
  NAND \DP_OP_25_64_3291/U24  ( .A(\DP_OP_25_64_3291/n146 ), .B(
        \DP_OP_25_64_3291/n130 ), .Z(\DP_OP_25_64_3291/n89 ) );
  NAND \DP_OP_25_64_3291/U34  ( .A(\DP_OP_25_64_3291/n88 ), .B(
        \DP_OP_25_64_3291/n89 ), .Z(\DP_OP_25_64_3291/n145 ) );
  NAND \DP_OP_25_64_3291/U13  ( .A(\DP_OP_25_64_3291/n166 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_3291/n95 ) );
  NAND \DP_OP_25_64_3291/U23  ( .A(\DP_OP_25_64_3291/n147 ), .B(
        \DP_OP_25_64_3291/n131 ), .Z(\DP_OP_25_64_3291/n96 ) );
  NAND \DP_OP_25_64_3291/U33  ( .A(\DP_OP_25_64_3291/n95 ), .B(
        \DP_OP_25_64_3291/n96 ), .Z(\DP_OP_25_64_3291/n146 ) );
  NAND \DP_OP_25_64_3291/U12  ( .A(\DP_OP_25_64_3291/n167 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_3291/n102 ) );
  NAND \DP_OP_25_64_3291/U22  ( .A(\DP_OP_25_64_3291/n148 ), .B(
        \DP_OP_25_64_3291/n132 ), .Z(\DP_OP_25_64_3291/n103 ) );
  NAND \DP_OP_25_64_3291/U32  ( .A(\DP_OP_25_64_3291/n102 ), .B(
        \DP_OP_25_64_3291/n103 ), .Z(\DP_OP_25_64_3291/n147 ) );
  NAND \DP_OP_25_64_3291/U11  ( .A(\DP_OP_25_64_3291/n168 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_3291/n109 ) );
  NAND \DP_OP_25_64_3291/U21  ( .A(\DP_OP_25_64_3291/n149 ), .B(
        \DP_OP_25_64_3291/n133 ), .Z(\DP_OP_25_64_3291/n110 ) );
  NAND \DP_OP_25_64_3291/U31  ( .A(\DP_OP_25_64_3291/n109 ), .B(
        \DP_OP_25_64_3291/n110 ), .Z(\DP_OP_25_64_3291/n148 ) );
  NAND \DP_OP_25_64_3291/U1  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_3291/n116 ) );
  NAND \DP_OP_25_64_3291/U2  ( .A(\DP_OP_25_64_3291/n134 ), .B(
        \DP_OP_25_64_3291/n169 ), .Z(\DP_OP_25_64_3291/n117 ) );
  NAND \DP_OP_25_64_3291/U3  ( .A(\DP_OP_25_64_3291/n116 ), .B(
        \DP_OP_25_64_3291/n117 ), .Z(\DP_OP_25_64_3291/n149 ) );
  AND U760 ( .A(o[2]), .B(\stack[1][7] ), .Z(n988) );
  NAND U761 ( .A(n1509), .B(n1511), .Z(n759) );
  XOR U762 ( .A(n1511), .B(n1509), .Z(n760) );
  NANDN U763 ( .A(n1508), .B(n760), .Z(n761) );
  NAND U764 ( .A(n759), .B(n761), .Z(n1235) );
  AND U765 ( .A(o[2]), .B(\stack[1][9] ), .Z(n1055) );
  XOR U766 ( .A(n1107), .B(n1108), .Z(n762) );
  NANDN U767 ( .A(n1109), .B(n762), .Z(n763) );
  NAND U768 ( .A(n1107), .B(n1108), .Z(n764) );
  AND U769 ( .A(n763), .B(n764), .Z(n965) );
  NAND U770 ( .A(n1467), .B(n1469), .Z(n765) );
  XOR U771 ( .A(n1469), .B(n1467), .Z(n766) );
  NAND U772 ( .A(n766), .B(n1466), .Z(n767) );
  NAND U773 ( .A(n765), .B(n767), .Z(n1205) );
  AND U774 ( .A(o[2]), .B(\stack[1][10] ), .Z(n1157) );
  XOR U775 ( .A(n1217), .B(n1218), .Z(n768) );
  NANDN U776 ( .A(n1219), .B(n768), .Z(n769) );
  NAND U777 ( .A(n1217), .B(n1218), .Z(n770) );
  AND U778 ( .A(n769), .B(n770), .Z(n1106) );
  XOR U779 ( .A(n1118), .B(n1119), .Z(n771) );
  XNOR U780 ( .A(n1120), .B(n771), .Z(n1184) );
  XOR U781 ( .A(n1328), .B(n1329), .Z(n1438) );
  NAND U782 ( .A(n1523), .B(n1525), .Z(n772) );
  XOR U783 ( .A(n1525), .B(n1523), .Z(n773) );
  NANDN U784 ( .A(n1522), .B(n773), .Z(n774) );
  NAND U785 ( .A(n772), .B(n774), .Z(n1319) );
  AND U786 ( .A(o[2]), .B(\stack[1][11] ), .Z(n1302) );
  XOR U787 ( .A(n1118), .B(n1119), .Z(n775) );
  NANDN U788 ( .A(n1120), .B(n775), .Z(n776) );
  NAND U789 ( .A(n1118), .B(n1119), .Z(n777) );
  AND U790 ( .A(n776), .B(n777), .Z(n1177) );
  XNOR U791 ( .A(n1343), .B(n1342), .Z(n1389) );
  XOR U792 ( .A(n1217), .B(n1218), .Z(n778) );
  XNOR U793 ( .A(n1219), .B(n778), .Z(n1486) );
  XNOR U794 ( .A(n1514), .B(n1515), .Z(n1516) );
  XNOR U795 ( .A(n1500), .B(n1501), .Z(n1502) );
  XNOR U796 ( .A(n1472), .B(n1473), .Z(n1474) );
  XNOR U797 ( .A(n1458), .B(n1459), .Z(n1460) );
  XNOR U798 ( .A(n1528), .B(n1529), .Z(n1532) );
  XOR U799 ( .A(n1338), .B(n1339), .Z(n1342) );
  XOR U800 ( .A(n1394), .B(n1395), .Z(n1411) );
  XOR U801 ( .A(n1107), .B(n1108), .Z(n779) );
  XNOR U802 ( .A(n1109), .B(n779), .Z(n1186) );
  XOR U803 ( .A(n1322), .B(n1323), .Z(n1426) );
  XNOR U804 ( .A(n1188), .B(n1189), .Z(n1480) );
  XNOR U805 ( .A(n1532), .B(n1531), .Z(n1578) );
  XOR U806 ( .A(n1516), .B(n1517), .Z(n1655) );
  XOR U807 ( .A(n1502), .B(n1503), .Z(n1732) );
  XOR U808 ( .A(n1488), .B(n1489), .Z(n1809) );
  XOR U809 ( .A(n1474), .B(n1475), .Z(n1887) );
  XOR U810 ( .A(n1460), .B(n1461), .Z(n1965) );
  ANDN U811 ( .B(n852), .A(opcode[0]), .Z(n780) );
  NAND U812 ( .A(n780), .B(opcode[2]), .Z(n795) );
  XOR U813 ( .A(\DP_OP_25_64_3291/n149 ), .B(\DP_OP_25_64_3291/n133 ), .Z(n781) );
  NAND U814 ( .A(n781), .B(n849), .Z(n782) );
  NAND U815 ( .A(\stack[1][1] ), .B(n2093), .Z(n783) );
  NANDN U816 ( .A(n2081), .B(n2082), .Z(n784) );
  AND U817 ( .A(n783), .B(n784), .Z(n785) );
  NAND U818 ( .A(x[1]), .B(n796), .Z(n786) );
  ANDN U819 ( .B(n2081), .A(n2080), .Z(n787) );
  NAND U820 ( .A(n787), .B(n2092), .Z(n788) );
  AND U821 ( .A(n786), .B(n788), .Z(n789) );
  NAND U822 ( .A(n785), .B(n2083), .Z(n790) );
  NAND U823 ( .A(n790), .B(o[1]), .Z(n791) );
  AND U824 ( .A(n789), .B(n791), .Z(n792) );
  AND U825 ( .A(n782), .B(n792), .Z(n793) );
  NANDN U826 ( .A(n2096), .B(\stack[1][1] ), .Z(n794) );
  NAND U827 ( .A(n793), .B(n794), .Z(n647) );
  IV U828 ( .A(n795), .Z(n796) );
  IV U829 ( .A(opcode[1]), .Z(n852) );
  IV U830 ( .A(opcode[2]), .Z(n851) );
  NOR U831 ( .A(opcode[0]), .B(opcode[2]), .Z(n797) );
  NAND U832 ( .A(opcode[1]), .B(n797), .Z(n833) );
  ANDN U833 ( .B(opcode[0]), .A(opcode[1]), .Z(n834) );
  NANDN U834 ( .A(opcode[2]), .B(n834), .Z(n798) );
  NAND U835 ( .A(n833), .B(n798), .Z(n829) );
  AND U836 ( .A(o[15]), .B(n829), .Z(\U1/RSOP_16/C2/Z_15 ) );
  AND U837 ( .A(o[14]), .B(n829), .Z(\U1/RSOP_16/C2/Z_14 ) );
  AND U838 ( .A(o[13]), .B(n829), .Z(\U1/RSOP_16/C2/Z_13 ) );
  AND U839 ( .A(o[12]), .B(n829), .Z(\U1/RSOP_16/C2/Z_12 ) );
  AND U840 ( .A(o[11]), .B(n829), .Z(\U1/RSOP_16/C2/Z_11 ) );
  AND U841 ( .A(o[10]), .B(n829), .Z(\U1/RSOP_16/C2/Z_10 ) );
  AND U842 ( .A(o[9]), .B(n829), .Z(\U1/RSOP_16/C2/Z_9 ) );
  AND U843 ( .A(o[8]), .B(n829), .Z(\U1/RSOP_16/C2/Z_8 ) );
  AND U844 ( .A(o[7]), .B(n829), .Z(\U1/RSOP_16/C2/Z_7 ) );
  AND U845 ( .A(o[6]), .B(n829), .Z(\U1/RSOP_16/C2/Z_6 ) );
  AND U846 ( .A(o[5]), .B(n829), .Z(\U1/RSOP_16/C2/Z_5 ) );
  AND U847 ( .A(o[4]), .B(n829), .Z(\U1/RSOP_16/C2/Z_4 ) );
  AND U848 ( .A(o[3]), .B(n829), .Z(\U1/RSOP_16/C2/Z_3 ) );
  AND U849 ( .A(o[2]), .B(n829), .Z(\U1/RSOP_16/C2/Z_2 ) );
  AND U850 ( .A(o[1]), .B(n829), .Z(\U1/RSOP_16/C2/Z_1 ) );
  AND U851 ( .A(o[0]), .B(n829), .Z(\U1/RSOP_16/C2/Z_0 ) );
  AND U852 ( .A(n834), .B(opcode[2]), .Z(n832) );
  NAND U853 ( .A(n832), .B(o[15]), .Z(n800) );
  NAND U854 ( .A(\stack[1][15] ), .B(n829), .Z(n799) );
  NAND U855 ( .A(n800), .B(n799), .Z(\U1/RSOP_16/C3/Z_15 ) );
  NAND U856 ( .A(n832), .B(o[14]), .Z(n802) );
  NAND U857 ( .A(\stack[1][14] ), .B(n829), .Z(n801) );
  NAND U858 ( .A(n802), .B(n801), .Z(\U1/RSOP_16/C3/Z_14 ) );
  NAND U859 ( .A(n832), .B(o[13]), .Z(n804) );
  NAND U860 ( .A(\stack[1][13] ), .B(n829), .Z(n803) );
  NAND U861 ( .A(n804), .B(n803), .Z(\U1/RSOP_16/C3/Z_13 ) );
  NAND U862 ( .A(n832), .B(o[12]), .Z(n806) );
  NAND U863 ( .A(\stack[1][12] ), .B(n829), .Z(n805) );
  NAND U864 ( .A(n806), .B(n805), .Z(\U1/RSOP_16/C3/Z_12 ) );
  NAND U865 ( .A(n832), .B(o[11]), .Z(n808) );
  NAND U866 ( .A(\stack[1][11] ), .B(n829), .Z(n807) );
  NAND U867 ( .A(n808), .B(n807), .Z(\U1/RSOP_16/C3/Z_11 ) );
  NAND U868 ( .A(n832), .B(o[10]), .Z(n810) );
  NAND U869 ( .A(\stack[1][10] ), .B(n829), .Z(n809) );
  NAND U870 ( .A(n810), .B(n809), .Z(\U1/RSOP_16/C3/Z_10 ) );
  NAND U871 ( .A(n832), .B(o[9]), .Z(n812) );
  NAND U872 ( .A(\stack[1][9] ), .B(n829), .Z(n811) );
  NAND U873 ( .A(n812), .B(n811), .Z(\U1/RSOP_16/C3/Z_9 ) );
  NAND U874 ( .A(n832), .B(o[8]), .Z(n814) );
  NAND U875 ( .A(\stack[1][8] ), .B(n829), .Z(n813) );
  NAND U876 ( .A(n814), .B(n813), .Z(\U1/RSOP_16/C3/Z_8 ) );
  NAND U877 ( .A(n832), .B(o[7]), .Z(n816) );
  NAND U878 ( .A(\stack[1][7] ), .B(n829), .Z(n815) );
  NAND U879 ( .A(n816), .B(n815), .Z(\U1/RSOP_16/C3/Z_7 ) );
  NAND U880 ( .A(n832), .B(o[6]), .Z(n818) );
  NAND U881 ( .A(\stack[1][6] ), .B(n829), .Z(n817) );
  NAND U882 ( .A(n818), .B(n817), .Z(\U1/RSOP_16/C3/Z_6 ) );
  NAND U883 ( .A(n832), .B(o[5]), .Z(n820) );
  NAND U884 ( .A(\stack[1][5] ), .B(n829), .Z(n819) );
  NAND U885 ( .A(n820), .B(n819), .Z(\U1/RSOP_16/C3/Z_5 ) );
  NAND U886 ( .A(n832), .B(o[4]), .Z(n822) );
  NAND U887 ( .A(\stack[1][4] ), .B(n829), .Z(n821) );
  NAND U888 ( .A(n822), .B(n821), .Z(\U1/RSOP_16/C3/Z_4 ) );
  NAND U889 ( .A(n832), .B(o[3]), .Z(n824) );
  NAND U890 ( .A(\stack[1][3] ), .B(n829), .Z(n823) );
  NAND U891 ( .A(n824), .B(n823), .Z(\U1/RSOP_16/C3/Z_3 ) );
  NAND U892 ( .A(n832), .B(o[2]), .Z(n826) );
  NAND U893 ( .A(\stack[1][2] ), .B(n829), .Z(n825) );
  NAND U894 ( .A(n826), .B(n825), .Z(\U1/RSOP_16/C3/Z_2 ) );
  NAND U895 ( .A(n832), .B(o[1]), .Z(n828) );
  NAND U896 ( .A(\stack[1][1] ), .B(n829), .Z(n827) );
  NAND U897 ( .A(n828), .B(n827), .Z(\U1/RSOP_16/C3/Z_1 ) );
  NAND U898 ( .A(n832), .B(o[0]), .Z(n831) );
  NAND U899 ( .A(\stack[1][0] ), .B(n829), .Z(n830) );
  NAND U900 ( .A(n831), .B(n830), .Z(\U1/RSOP_16/C3/Z_0 ) );
  NANDN U901 ( .A(n832), .B(n833), .Z(\C1/Z_0 ) );
  NANDN U902 ( .A(n834), .B(n833), .Z(n849) );
  NAND U903 ( .A(\C3/DATA5_15 ), .B(n849), .Z(n835) );
  AND U904 ( .A(n1537), .B(n835), .Z(n1538) );
  NAND U905 ( .A(\C3/DATA5_14 ), .B(n849), .Z(n836) );
  AND U906 ( .A(n1576), .B(n836), .Z(n1588) );
  NAND U907 ( .A(\C3/DATA5_12 ), .B(n849), .Z(n837) );
  AND U908 ( .A(n1654), .B(n837), .Z(n1665) );
  NAND U909 ( .A(\C3/DATA5_10 ), .B(n849), .Z(n838) );
  AND U910 ( .A(n1731), .B(n838), .Z(n1742) );
  NAND U911 ( .A(\C3/DATA5_8 ), .B(n849), .Z(n839) );
  AND U912 ( .A(n1808), .B(n839), .Z(n1819) );
  NAND U913 ( .A(\C3/DATA5_7 ), .B(n849), .Z(n840) );
  AND U914 ( .A(n1846), .B(n840), .Z(n1851) );
  NAND U915 ( .A(\C3/DATA5_6 ), .B(n849), .Z(n841) );
  AND U916 ( .A(n1886), .B(n841), .Z(n1897) );
  NAND U917 ( .A(\C3/DATA5_5 ), .B(n849), .Z(n842) );
  AND U918 ( .A(n1924), .B(n842), .Z(n1929) );
  NAND U919 ( .A(\C3/DATA5_4 ), .B(n849), .Z(n843) );
  AND U920 ( .A(n1964), .B(n843), .Z(n1975) );
  NAND U921 ( .A(\C3/DATA5_3 ), .B(n849), .Z(n844) );
  AND U922 ( .A(n2008), .B(n844), .Z(n2009) );
  NAND U923 ( .A(\C3/DATA5_2 ), .B(n849), .Z(n845) );
  AND U924 ( .A(n2041), .B(n845), .Z(n2046) );
  NAND U925 ( .A(\C3/DATA5_0 ), .B(n849), .Z(n846) );
  AND U926 ( .A(n2091), .B(n846), .Z(n2101) );
  NAND U927 ( .A(\C3/DATA5_13 ), .B(n849), .Z(n847) );
  NAND U928 ( .A(n1626), .B(n847), .Z(n551) );
  NAND U929 ( .A(\C3/DATA5_11 ), .B(n849), .Z(n848) );
  NAND U930 ( .A(n1703), .B(n848), .Z(n567) );
  NAND U931 ( .A(\C3/DATA5_9 ), .B(n849), .Z(n850) );
  NAND U932 ( .A(n1780), .B(n850), .Z(n583) );
  NAND U933 ( .A(n796), .B(\stack[6][0] ), .Z(n854) );
  NAND U934 ( .A(n795), .B(\stack[7][0] ), .Z(n853) );
  NAND U935 ( .A(n854), .B(n853), .Z(n522) );
  NAND U936 ( .A(n796), .B(\stack[5][0] ), .Z(n857) );
  NAND U937 ( .A(opcode[0]), .B(n851), .Z(n855) );
  AND U938 ( .A(n855), .B(n852), .Z(n2084) );
  NANDN U939 ( .A(n2084), .B(\stack[7][0] ), .Z(n856) );
  AND U940 ( .A(n857), .B(n856), .Z(n859) );
  XNOR U941 ( .A(opcode[2]), .B(opcode[0]), .Z(n1541) );
  NAND U942 ( .A(n852), .B(n1541), .Z(n2087) );
  NANDN U943 ( .A(n2087), .B(\stack[6][0] ), .Z(n858) );
  NAND U944 ( .A(n859), .B(n858), .Z(n523) );
  NAND U945 ( .A(n796), .B(\stack[4][0] ), .Z(n861) );
  NANDN U946 ( .A(n2084), .B(\stack[6][0] ), .Z(n860) );
  AND U947 ( .A(n861), .B(n860), .Z(n863) );
  NANDN U948 ( .A(n2087), .B(\stack[5][0] ), .Z(n862) );
  NAND U949 ( .A(n863), .B(n862), .Z(n524) );
  NAND U950 ( .A(n796), .B(\stack[3][0] ), .Z(n865) );
  NANDN U951 ( .A(n2084), .B(\stack[5][0] ), .Z(n864) );
  AND U952 ( .A(n865), .B(n864), .Z(n867) );
  NANDN U953 ( .A(n2087), .B(\stack[4][0] ), .Z(n866) );
  NAND U954 ( .A(n867), .B(n866), .Z(n525) );
  NAND U955 ( .A(n796), .B(\stack[2][0] ), .Z(n869) );
  NANDN U956 ( .A(n2084), .B(\stack[4][0] ), .Z(n868) );
  AND U957 ( .A(n869), .B(n868), .Z(n871) );
  NANDN U958 ( .A(n2087), .B(\stack[3][0] ), .Z(n870) );
  NAND U959 ( .A(n871), .B(n870), .Z(n526) );
  NAND U960 ( .A(\stack[1][0] ), .B(n796), .Z(n873) );
  NANDN U961 ( .A(n2084), .B(\stack[3][0] ), .Z(n872) );
  AND U962 ( .A(n873), .B(n872), .Z(n875) );
  NANDN U963 ( .A(n2087), .B(\stack[2][0] ), .Z(n874) );
  NAND U964 ( .A(n875), .B(n874), .Z(n527) );
  NAND U965 ( .A(n796), .B(\stack[6][15] ), .Z(n877) );
  NAND U966 ( .A(n795), .B(\stack[7][15] ), .Z(n876) );
  NAND U967 ( .A(n877), .B(n876), .Z(n528) );
  NAND U968 ( .A(n796), .B(\stack[5][15] ), .Z(n879) );
  NANDN U969 ( .A(n2084), .B(\stack[7][15] ), .Z(n878) );
  AND U970 ( .A(n879), .B(n878), .Z(n881) );
  NANDN U971 ( .A(n2087), .B(\stack[6][15] ), .Z(n880) );
  NAND U972 ( .A(n881), .B(n880), .Z(n529) );
  NAND U973 ( .A(n796), .B(\stack[4][15] ), .Z(n883) );
  NANDN U974 ( .A(n2084), .B(\stack[6][15] ), .Z(n882) );
  AND U975 ( .A(n883), .B(n882), .Z(n885) );
  NANDN U976 ( .A(n2087), .B(\stack[5][15] ), .Z(n884) );
  NAND U977 ( .A(n885), .B(n884), .Z(n530) );
  NAND U978 ( .A(n796), .B(\stack[3][15] ), .Z(n887) );
  NANDN U979 ( .A(n2084), .B(\stack[5][15] ), .Z(n886) );
  AND U980 ( .A(n887), .B(n886), .Z(n889) );
  NANDN U981 ( .A(n2087), .B(\stack[4][15] ), .Z(n888) );
  NAND U982 ( .A(n889), .B(n888), .Z(n531) );
  NAND U983 ( .A(n796), .B(\stack[2][15] ), .Z(n891) );
  NANDN U984 ( .A(n2084), .B(\stack[4][15] ), .Z(n890) );
  AND U985 ( .A(n891), .B(n890), .Z(n893) );
  NANDN U986 ( .A(n2087), .B(\stack[3][15] ), .Z(n892) );
  NAND U987 ( .A(n893), .B(n892), .Z(n532) );
  NAND U988 ( .A(n796), .B(\stack[1][15] ), .Z(n895) );
  NANDN U989 ( .A(n2084), .B(\stack[3][15] ), .Z(n894) );
  AND U990 ( .A(n895), .B(n894), .Z(n897) );
  NANDN U991 ( .A(n2087), .B(\stack[2][15] ), .Z(n896) );
  NAND U992 ( .A(n897), .B(n896), .Z(n533) );
  NAND U993 ( .A(n796), .B(o[15]), .Z(n899) );
  NANDN U994 ( .A(n2084), .B(\stack[2][15] ), .Z(n898) );
  AND U995 ( .A(n899), .B(n898), .Z(n901) );
  NANDN U996 ( .A(n2087), .B(\stack[1][15] ), .Z(n900) );
  NAND U997 ( .A(n901), .B(n900), .Z(n534) );
  IV U998 ( .A(\stack[1][3] ), .Z(n1256) );
  ANDN U999 ( .B(o[7]), .A(n1256), .Z(n964) );
  ANDN U1000 ( .B(o[5]), .A(n1256), .Z(n923) );
  IV U1001 ( .A(o[0]), .Z(n1445) );
  ANDN U1002 ( .B(\stack[1][6] ), .A(n1445), .Z(n904) );
  NAND U1003 ( .A(\stack[1][5] ), .B(o[1]), .Z(n905) );
  ANDN U1004 ( .B(n904), .A(n905), .Z(n933) );
  IV U1005 ( .A(\stack[1][5] ), .Z(n1270) );
  ANDN U1006 ( .B(o[2]), .A(n1270), .Z(n934) );
  XNOR U1007 ( .A(n933), .B(n934), .Z(n936) );
  NAND U1008 ( .A(\stack[1][6] ), .B(o[1]), .Z(n931) );
  ANDN U1009 ( .B(\stack[1][7] ), .A(n1445), .Z(n932) );
  XNOR U1010 ( .A(n931), .B(n932), .Z(n935) );
  XNOR U1011 ( .A(n936), .B(n935), .Z(n928) );
  IV U1012 ( .A(\stack[1][4] ), .Z(n1316) );
  ANDN U1013 ( .B(o[2]), .A(n1316), .Z(n902) );
  ANDN U1014 ( .B(\stack[1][5] ), .A(n1445), .Z(n910) );
  NAND U1015 ( .A(\stack[1][4] ), .B(o[1]), .Z(n911) );
  ANDN U1016 ( .B(n910), .A(n911), .Z(n903) );
  OR U1017 ( .A(n902), .B(n903), .Z(n907) );
  XNOR U1018 ( .A(n903), .B(n902), .Z(n915) );
  XNOR U1019 ( .A(n905), .B(n904), .Z(n914) );
  OR U1020 ( .A(n915), .B(n914), .Z(n906) );
  AND U1021 ( .A(n907), .B(n906), .Z(n926) );
  NAND U1022 ( .A(\stack[1][4] ), .B(o[3]), .Z(n925) );
  XOR U1023 ( .A(n926), .B(n925), .Z(n927) );
  XNOR U1024 ( .A(n928), .B(n927), .Z(n919) );
  IV U1025 ( .A(n919), .Z(n1097) );
  ANDN U1026 ( .B(o[2]), .A(n1256), .Z(n908) );
  ANDN U1027 ( .B(\stack[1][4] ), .A(n1445), .Z(n1078) );
  NAND U1028 ( .A(\stack[1][3] ), .B(o[1]), .Z(n1079) );
  ANDN U1029 ( .B(n1078), .A(n1079), .Z(n909) );
  OR U1030 ( .A(n908), .B(n909), .Z(n913) );
  XNOR U1031 ( .A(n909), .B(n908), .Z(n1083) );
  XNOR U1032 ( .A(n911), .B(n910), .Z(n1082) );
  OR U1033 ( .A(n1083), .B(n1082), .Z(n912) );
  AND U1034 ( .A(n913), .B(n912), .Z(n916) );
  ANDN U1035 ( .B(o[3]), .A(n1256), .Z(n2002) );
  OR U1036 ( .A(n916), .B(n2002), .Z(n918) );
  XNOR U1037 ( .A(n915), .B(n914), .Z(n1089) );
  XNOR U1038 ( .A(n2002), .B(n916), .Z(n1088) );
  OR U1039 ( .A(n1089), .B(n1088), .Z(n917) );
  NAND U1040 ( .A(n918), .B(n917), .Z(n1100) );
  NAND U1041 ( .A(n1097), .B(n1100), .Z(n922) );
  ANDN U1042 ( .B(n919), .A(n1100), .Z(n920) );
  NAND U1043 ( .A(\stack[1][3] ), .B(o[4]), .Z(n1098) );
  NANDN U1044 ( .A(n920), .B(n1098), .Z(n921) );
  NAND U1045 ( .A(n922), .B(n921), .Z(n924) );
  NANDN U1046 ( .A(n923), .B(n924), .Z(n941) );
  XOR U1047 ( .A(n924), .B(n923), .Z(n1104) );
  NANDN U1048 ( .A(n926), .B(n925), .Z(n930) );
  OR U1049 ( .A(n928), .B(n927), .Z(n929) );
  AND U1050 ( .A(n930), .B(n929), .Z(n944) );
  NAND U1051 ( .A(\stack[1][4] ), .B(o[4]), .Z(n945) );
  ANDN U1052 ( .B(n932), .A(n931), .Z(n957) );
  IV U1053 ( .A(\stack[1][6] ), .Z(n1315) );
  ANDN U1054 ( .B(o[2]), .A(n1315), .Z(n958) );
  XNOR U1055 ( .A(n957), .B(n958), .Z(n960) );
  NAND U1056 ( .A(\stack[1][7] ), .B(o[1]), .Z(n955) );
  ANDN U1057 ( .B(\stack[1][8] ), .A(n1445), .Z(n956) );
  XNOR U1058 ( .A(n955), .B(n956), .Z(n959) );
  XNOR U1059 ( .A(n960), .B(n959), .Z(n952) );
  OR U1060 ( .A(n934), .B(n933), .Z(n938) );
  OR U1061 ( .A(n936), .B(n935), .Z(n937) );
  AND U1062 ( .A(n938), .B(n937), .Z(n950) );
  NAND U1063 ( .A(\stack[1][5] ), .B(o[3]), .Z(n949) );
  XOR U1064 ( .A(n950), .B(n949), .Z(n951) );
  XNOR U1065 ( .A(n952), .B(n951), .Z(n943) );
  IV U1066 ( .A(n943), .Z(n942) );
  XOR U1067 ( .A(n945), .B(n942), .Z(n939) );
  XOR U1068 ( .A(n944), .B(n939), .Z(n1103) );
  OR U1069 ( .A(n1104), .B(n1103), .Z(n940) );
  AND U1070 ( .A(n941), .B(n940), .Z(n1108) );
  NANDN U1071 ( .A(n944), .B(n942), .Z(n948) );
  AND U1072 ( .A(n944), .B(n943), .Z(n946) );
  NANDN U1073 ( .A(n946), .B(n945), .Z(n947) );
  NAND U1074 ( .A(n948), .B(n947), .Z(n966) );
  ANDN U1075 ( .B(o[5]), .A(n1316), .Z(n967) );
  XOR U1076 ( .A(n966), .B(n967), .Z(n969) );
  NANDN U1077 ( .A(n950), .B(n949), .Z(n954) );
  OR U1078 ( .A(n952), .B(n951), .Z(n953) );
  AND U1079 ( .A(n954), .B(n953), .Z(n974) );
  NAND U1080 ( .A(\stack[1][5] ), .B(o[4]), .Z(n975) );
  ANDN U1081 ( .B(n956), .A(n955), .Z(n987) );
  XNOR U1082 ( .A(n987), .B(n988), .Z(n990) );
  NAND U1083 ( .A(\stack[1][8] ), .B(o[1]), .Z(n985) );
  ANDN U1084 ( .B(\stack[1][9] ), .A(n1445), .Z(n986) );
  XNOR U1085 ( .A(n985), .B(n986), .Z(n989) );
  XNOR U1086 ( .A(n990), .B(n989), .Z(n982) );
  OR U1087 ( .A(n958), .B(n957), .Z(n962) );
  OR U1088 ( .A(n960), .B(n959), .Z(n961) );
  AND U1089 ( .A(n962), .B(n961), .Z(n980) );
  NAND U1090 ( .A(\stack[1][6] ), .B(o[3]), .Z(n979) );
  XOR U1091 ( .A(n980), .B(n979), .Z(n981) );
  XNOR U1092 ( .A(n982), .B(n981), .Z(n973) );
  IV U1093 ( .A(n973), .Z(n972) );
  XOR U1094 ( .A(n975), .B(n972), .Z(n963) );
  XOR U1095 ( .A(n974), .B(n963), .Z(n968) );
  XNOR U1096 ( .A(n969), .B(n968), .Z(n1107) );
  NAND U1097 ( .A(\stack[1][3] ), .B(o[6]), .Z(n1109) );
  NANDN U1098 ( .A(n964), .B(n965), .Z(n996) );
  XOR U1099 ( .A(n965), .B(n964), .Z(n1076) );
  NANDN U1100 ( .A(n967), .B(n966), .Z(n971) );
  OR U1101 ( .A(n969), .B(n968), .Z(n970) );
  AND U1102 ( .A(n971), .B(n970), .Z(n999) );
  NAND U1103 ( .A(\stack[1][4] ), .B(o[6]), .Z(n1000) );
  NANDN U1104 ( .A(n974), .B(n972), .Z(n978) );
  AND U1105 ( .A(n974), .B(n973), .Z(n976) );
  NANDN U1106 ( .A(n976), .B(n975), .Z(n977) );
  NAND U1107 ( .A(n978), .B(n977), .Z(n1026) );
  NAND U1108 ( .A(\stack[1][5] ), .B(o[5]), .Z(n1930) );
  XNOR U1109 ( .A(n1026), .B(n1930), .Z(n1028) );
  NANDN U1110 ( .A(n980), .B(n979), .Z(n984) );
  OR U1111 ( .A(n982), .B(n981), .Z(n983) );
  AND U1112 ( .A(n984), .B(n983), .Z(n1006) );
  NAND U1113 ( .A(\stack[1][6] ), .B(o[4]), .Z(n1007) );
  ANDN U1114 ( .B(n986), .A(n985), .Z(n1019) );
  IV U1115 ( .A(\stack[1][8] ), .Z(n1284) );
  ANDN U1116 ( .B(o[2]), .A(n1284), .Z(n1020) );
  XNOR U1117 ( .A(n1019), .B(n1020), .Z(n1022) );
  NAND U1118 ( .A(\stack[1][9] ), .B(o[1]), .Z(n1017) );
  ANDN U1119 ( .B(\stack[1][10] ), .A(n1445), .Z(n1018) );
  XNOR U1120 ( .A(n1017), .B(n1018), .Z(n1021) );
  XNOR U1121 ( .A(n1022), .B(n1021), .Z(n1014) );
  OR U1122 ( .A(n988), .B(n987), .Z(n992) );
  OR U1123 ( .A(n990), .B(n989), .Z(n991) );
  AND U1124 ( .A(n992), .B(n991), .Z(n1012) );
  NAND U1125 ( .A(\stack[1][7] ), .B(o[3]), .Z(n1011) );
  XOR U1126 ( .A(n1012), .B(n1011), .Z(n1013) );
  XNOR U1127 ( .A(n1014), .B(n1013), .Z(n1005) );
  IV U1128 ( .A(n1005), .Z(n1004) );
  XOR U1129 ( .A(n1007), .B(n1004), .Z(n993) );
  XOR U1130 ( .A(n1006), .B(n993), .Z(n1027) );
  XNOR U1131 ( .A(n1028), .B(n1027), .Z(n998) );
  IV U1132 ( .A(n998), .Z(n997) );
  XOR U1133 ( .A(n1000), .B(n997), .Z(n994) );
  XOR U1134 ( .A(n999), .B(n994), .Z(n1075) );
  OR U1135 ( .A(n1076), .B(n1075), .Z(n995) );
  AND U1136 ( .A(n996), .B(n995), .Z(n1119) );
  NANDN U1137 ( .A(n999), .B(n997), .Z(n1003) );
  AND U1138 ( .A(n999), .B(n998), .Z(n1001) );
  NANDN U1139 ( .A(n1001), .B(n1000), .Z(n1002) );
  NAND U1140 ( .A(n1003), .B(n1002), .Z(n1068) );
  ANDN U1141 ( .B(o[7]), .A(n1316), .Z(n1069) );
  XOR U1142 ( .A(n1068), .B(n1069), .Z(n1071) );
  NAND U1143 ( .A(\stack[1][5] ), .B(o[6]), .Z(n1035) );
  NANDN U1144 ( .A(n1006), .B(n1004), .Z(n1010) );
  AND U1145 ( .A(n1006), .B(n1005), .Z(n1008) );
  NANDN U1146 ( .A(n1008), .B(n1007), .Z(n1009) );
  NAND U1147 ( .A(n1010), .B(n1009), .Z(n1061) );
  IV U1148 ( .A(o[5]), .Z(n1292) );
  ANDN U1149 ( .B(\stack[1][6] ), .A(n1292), .Z(n1062) );
  XOR U1150 ( .A(n1061), .B(n1062), .Z(n1064) );
  NANDN U1151 ( .A(n1012), .B(n1011), .Z(n1016) );
  OR U1152 ( .A(n1014), .B(n1013), .Z(n1015) );
  AND U1153 ( .A(n1016), .B(n1015), .Z(n1041) );
  NAND U1154 ( .A(\stack[1][7] ), .B(o[4]), .Z(n1042) );
  ANDN U1155 ( .B(n1018), .A(n1017), .Z(n1054) );
  XNOR U1156 ( .A(n1054), .B(n1055), .Z(n1057) );
  NAND U1157 ( .A(\stack[1][10] ), .B(o[1]), .Z(n1052) );
  ANDN U1158 ( .B(\stack[1][11] ), .A(n1445), .Z(n1053) );
  XNOR U1159 ( .A(n1052), .B(n1053), .Z(n1056) );
  XNOR U1160 ( .A(n1057), .B(n1056), .Z(n1049) );
  OR U1161 ( .A(n1020), .B(n1019), .Z(n1024) );
  OR U1162 ( .A(n1022), .B(n1021), .Z(n1023) );
  AND U1163 ( .A(n1024), .B(n1023), .Z(n1047) );
  NAND U1164 ( .A(\stack[1][8] ), .B(o[3]), .Z(n1046) );
  XOR U1165 ( .A(n1047), .B(n1046), .Z(n1048) );
  XNOR U1166 ( .A(n1049), .B(n1048), .Z(n1040) );
  IV U1167 ( .A(n1040), .Z(n1039) );
  XOR U1168 ( .A(n1042), .B(n1039), .Z(n1025) );
  XOR U1169 ( .A(n1041), .B(n1025), .Z(n1063) );
  XNOR U1170 ( .A(n1064), .B(n1063), .Z(n1033) );
  IV U1171 ( .A(n1033), .Z(n1032) );
  NAND U1172 ( .A(n1930), .B(n1026), .Z(n1030) );
  OR U1173 ( .A(n1028), .B(n1027), .Z(n1029) );
  AND U1174 ( .A(n1030), .B(n1029), .Z(n1034) );
  XOR U1175 ( .A(n1032), .B(n1034), .Z(n1031) );
  XOR U1176 ( .A(n1035), .B(n1031), .Z(n1070) );
  XNOR U1177 ( .A(n1071), .B(n1070), .Z(n1118) );
  NAND U1178 ( .A(\stack[1][3] ), .B(o[8]), .Z(n1120) );
  ANDN U1179 ( .B(o[9]), .A(n1256), .Z(n1178) );
  XOR U1180 ( .A(n1177), .B(n1178), .Z(n1180) );
  NAND U1181 ( .A(\stack[1][4] ), .B(o[8]), .Z(n1130) );
  NANDN U1182 ( .A(n1034), .B(n1032), .Z(n1038) );
  AND U1183 ( .A(n1034), .B(n1033), .Z(n1036) );
  NANDN U1184 ( .A(n1036), .B(n1035), .Z(n1037) );
  NAND U1185 ( .A(n1038), .B(n1037), .Z(n1170) );
  ANDN U1186 ( .B(o[7]), .A(n1270), .Z(n1171) );
  XOR U1187 ( .A(n1170), .B(n1171), .Z(n1173) );
  NAND U1188 ( .A(\stack[1][6] ), .B(o[6]), .Z(n1137) );
  NANDN U1189 ( .A(n1041), .B(n1039), .Z(n1045) );
  AND U1190 ( .A(n1041), .B(n1040), .Z(n1043) );
  NANDN U1191 ( .A(n1043), .B(n1042), .Z(n1044) );
  NAND U1192 ( .A(n1045), .B(n1044), .Z(n1163) );
  ANDN U1193 ( .B(\stack[1][7] ), .A(n1292), .Z(n1164) );
  XOR U1194 ( .A(n1163), .B(n1164), .Z(n1166) );
  NANDN U1195 ( .A(n1047), .B(n1046), .Z(n1051) );
  OR U1196 ( .A(n1049), .B(n1048), .Z(n1050) );
  AND U1197 ( .A(n1051), .B(n1050), .Z(n1143) );
  NAND U1198 ( .A(\stack[1][8] ), .B(o[4]), .Z(n1144) );
  ANDN U1199 ( .B(n1053), .A(n1052), .Z(n1156) );
  XNOR U1200 ( .A(n1156), .B(n1157), .Z(n1159) );
  NAND U1201 ( .A(\stack[1][11] ), .B(o[1]), .Z(n1154) );
  ANDN U1202 ( .B(\stack[1][12] ), .A(n1445), .Z(n1155) );
  XNOR U1203 ( .A(n1154), .B(n1155), .Z(n1158) );
  XNOR U1204 ( .A(n1159), .B(n1158), .Z(n1151) );
  OR U1205 ( .A(n1055), .B(n1054), .Z(n1059) );
  OR U1206 ( .A(n1057), .B(n1056), .Z(n1058) );
  AND U1207 ( .A(n1059), .B(n1058), .Z(n1149) );
  NAND U1208 ( .A(\stack[1][9] ), .B(o[3]), .Z(n1148) );
  XOR U1209 ( .A(n1149), .B(n1148), .Z(n1150) );
  XNOR U1210 ( .A(n1151), .B(n1150), .Z(n1142) );
  IV U1211 ( .A(n1142), .Z(n1141) );
  XOR U1212 ( .A(n1144), .B(n1141), .Z(n1060) );
  XOR U1213 ( .A(n1143), .B(n1060), .Z(n1165) );
  XNOR U1214 ( .A(n1166), .B(n1165), .Z(n1135) );
  IV U1215 ( .A(n1135), .Z(n1134) );
  NANDN U1216 ( .A(n1062), .B(n1061), .Z(n1066) );
  OR U1217 ( .A(n1064), .B(n1063), .Z(n1065) );
  AND U1218 ( .A(n1066), .B(n1065), .Z(n1136) );
  XOR U1219 ( .A(n1134), .B(n1136), .Z(n1067) );
  XOR U1220 ( .A(n1137), .B(n1067), .Z(n1172) );
  XNOR U1221 ( .A(n1173), .B(n1172), .Z(n1128) );
  IV U1222 ( .A(n1128), .Z(n1127) );
  NANDN U1223 ( .A(n1069), .B(n1068), .Z(n1073) );
  OR U1224 ( .A(n1071), .B(n1070), .Z(n1072) );
  AND U1225 ( .A(n1073), .B(n1072), .Z(n1129) );
  XOR U1226 ( .A(n1127), .B(n1129), .Z(n1074) );
  XOR U1227 ( .A(n1130), .B(n1074), .Z(n1179) );
  XNOR U1228 ( .A(n1180), .B(n1179), .Z(n1123) );
  IV U1229 ( .A(n1123), .Z(n1236) );
  IV U1230 ( .A(\stack[1][2] ), .Z(n1317) );
  ANDN U1231 ( .B(o[9]), .A(n1317), .Z(n1116) );
  XNOR U1232 ( .A(n1076), .B(n1075), .Z(n1112) );
  IV U1233 ( .A(n1112), .Z(n1228) );
  ANDN U1234 ( .B(o[7]), .A(n1317), .Z(n1105) );
  ANDN U1235 ( .B(o[5]), .A(n1317), .Z(n1095) );
  ANDN U1236 ( .B(o[3]), .A(n1317), .Z(n1084) );
  NAND U1237 ( .A(\stack[1][2] ), .B(o[1]), .Z(n1195) );
  NAND U1238 ( .A(o[0]), .B(\stack[1][3] ), .Z(n1194) );
  NOR U1239 ( .A(n1195), .B(n1194), .Z(n1077) );
  NAND U1240 ( .A(\stack[1][2] ), .B(o[2]), .Z(n2047) );
  NANDN U1241 ( .A(n1077), .B(n2047), .Z(n1081) );
  XOR U1242 ( .A(n1077), .B(n2047), .Z(n1199) );
  XNOR U1243 ( .A(n1079), .B(n1078), .Z(n1198) );
  OR U1244 ( .A(n1199), .B(n1198), .Z(n1080) );
  AND U1245 ( .A(n1081), .B(n1080), .Z(n1085) );
  OR U1246 ( .A(n1084), .B(n1085), .Z(n1087) );
  XNOR U1247 ( .A(n1083), .B(n1082), .Z(n1191) );
  XNOR U1248 ( .A(n1085), .B(n1084), .Z(n1190) );
  OR U1249 ( .A(n1191), .B(n1190), .Z(n1086) );
  NAND U1250 ( .A(n1087), .B(n1086), .Z(n1090) );
  XNOR U1251 ( .A(n1089), .B(n1088), .Z(n1091) );
  IV U1252 ( .A(n1091), .Z(n1209) );
  NAND U1253 ( .A(n1090), .B(n1209), .Z(n1094) );
  IV U1254 ( .A(n1090), .Z(n1207) );
  AND U1255 ( .A(n1091), .B(n1207), .Z(n1092) );
  NAND U1256 ( .A(\stack[1][2] ), .B(o[4]), .Z(n1206) );
  NANDN U1257 ( .A(n1092), .B(n1206), .Z(n1093) );
  NAND U1258 ( .A(n1094), .B(n1093), .Z(n1096) );
  NANDN U1259 ( .A(n1095), .B(n1096), .Z(n1102) );
  XOR U1260 ( .A(n1096), .B(n1095), .Z(n1189) );
  XOR U1261 ( .A(n1098), .B(n1097), .Z(n1099) );
  XOR U1262 ( .A(n1100), .B(n1099), .Z(n1188) );
  NANDN U1263 ( .A(n1189), .B(n1188), .Z(n1101) );
  AND U1264 ( .A(n1102), .B(n1101), .Z(n1218) );
  XNOR U1265 ( .A(n1104), .B(n1103), .Z(n1217) );
  NAND U1266 ( .A(\stack[1][2] ), .B(o[6]), .Z(n1219) );
  NANDN U1267 ( .A(n1105), .B(n1106), .Z(n1111) );
  XOR U1268 ( .A(n1106), .B(n1105), .Z(n1187) );
  OR U1269 ( .A(n1187), .B(n1186), .Z(n1110) );
  NAND U1270 ( .A(n1111), .B(n1110), .Z(n1231) );
  NAND U1271 ( .A(n1228), .B(n1231), .Z(n1115) );
  ANDN U1272 ( .B(n1112), .A(n1231), .Z(n1113) );
  NAND U1273 ( .A(\stack[1][2] ), .B(o[8]), .Z(n1229) );
  NANDN U1274 ( .A(n1113), .B(n1229), .Z(n1114) );
  NAND U1275 ( .A(n1115), .B(n1114), .Z(n1117) );
  NANDN U1276 ( .A(n1116), .B(n1117), .Z(n1122) );
  XOR U1277 ( .A(n1117), .B(n1116), .Z(n1185) );
  OR U1278 ( .A(n1185), .B(n1184), .Z(n1121) );
  NAND U1279 ( .A(n1122), .B(n1121), .Z(n1239) );
  NAND U1280 ( .A(n1236), .B(n1239), .Z(n1126) );
  ANDN U1281 ( .B(n1123), .A(n1239), .Z(n1124) );
  NAND U1282 ( .A(\stack[1][2] ), .B(o[10]), .Z(n1237) );
  NANDN U1283 ( .A(n1124), .B(n1237), .Z(n1125) );
  NAND U1284 ( .A(n1126), .B(n1125), .Z(n1243) );
  ANDN U1285 ( .B(o[11]), .A(n1317), .Z(n1244) );
  XOR U1286 ( .A(n1243), .B(n1244), .Z(n1246) );
  NAND U1287 ( .A(\stack[1][3] ), .B(o[10]), .Z(n1252) );
  NANDN U1288 ( .A(n1129), .B(n1127), .Z(n1133) );
  AND U1289 ( .A(n1129), .B(n1128), .Z(n1131) );
  NANDN U1290 ( .A(n1131), .B(n1130), .Z(n1132) );
  NAND U1291 ( .A(n1133), .B(n1132), .Z(n1257) );
  ANDN U1292 ( .B(o[9]), .A(n1316), .Z(n1258) );
  XOR U1293 ( .A(n1257), .B(n1258), .Z(n1260) );
  NAND U1294 ( .A(\stack[1][5] ), .B(o[8]), .Z(n1266) );
  NANDN U1295 ( .A(n1136), .B(n1134), .Z(n1140) );
  AND U1296 ( .A(n1136), .B(n1135), .Z(n1138) );
  NANDN U1297 ( .A(n1138), .B(n1137), .Z(n1139) );
  NAND U1298 ( .A(n1140), .B(n1139), .Z(n1271) );
  ANDN U1299 ( .B(o[7]), .A(n1315), .Z(n1272) );
  XOR U1300 ( .A(n1271), .B(n1272), .Z(n1274) );
  NAND U1301 ( .A(\stack[1][7] ), .B(o[6]), .Z(n1280) );
  NANDN U1302 ( .A(n1143), .B(n1141), .Z(n1147) );
  AND U1303 ( .A(n1143), .B(n1142), .Z(n1145) );
  NANDN U1304 ( .A(n1145), .B(n1144), .Z(n1146) );
  NAND U1305 ( .A(n1147), .B(n1146), .Z(n1308) );
  ANDN U1306 ( .B(\stack[1][8] ), .A(n1292), .Z(n1309) );
  XOR U1307 ( .A(n1308), .B(n1309), .Z(n1311) );
  NANDN U1308 ( .A(n1149), .B(n1148), .Z(n1153) );
  OR U1309 ( .A(n1151), .B(n1150), .Z(n1152) );
  AND U1310 ( .A(n1153), .B(n1152), .Z(n1287) );
  NAND U1311 ( .A(\stack[1][9] ), .B(o[4]), .Z(n1288) );
  ANDN U1312 ( .B(n1155), .A(n1154), .Z(n1301) );
  XNOR U1313 ( .A(n1301), .B(n1302), .Z(n1304) );
  NAND U1314 ( .A(\stack[1][12] ), .B(o[1]), .Z(n1299) );
  ANDN U1315 ( .B(\stack[1][13] ), .A(n1445), .Z(n1300) );
  XNOR U1316 ( .A(n1299), .B(n1300), .Z(n1303) );
  XNOR U1317 ( .A(n1304), .B(n1303), .Z(n1296) );
  OR U1318 ( .A(n1157), .B(n1156), .Z(n1161) );
  OR U1319 ( .A(n1159), .B(n1158), .Z(n1160) );
  AND U1320 ( .A(n1161), .B(n1160), .Z(n1294) );
  NAND U1321 ( .A(\stack[1][10] ), .B(o[3]), .Z(n1293) );
  XOR U1322 ( .A(n1294), .B(n1293), .Z(n1295) );
  XNOR U1323 ( .A(n1296), .B(n1295), .Z(n1286) );
  IV U1324 ( .A(n1286), .Z(n1285) );
  XOR U1325 ( .A(n1288), .B(n1285), .Z(n1162) );
  XOR U1326 ( .A(n1287), .B(n1162), .Z(n1310) );
  XNOR U1327 ( .A(n1311), .B(n1310), .Z(n1278) );
  IV U1328 ( .A(n1278), .Z(n1277) );
  NANDN U1329 ( .A(n1164), .B(n1163), .Z(n1168) );
  OR U1330 ( .A(n1166), .B(n1165), .Z(n1167) );
  AND U1331 ( .A(n1168), .B(n1167), .Z(n1279) );
  XOR U1332 ( .A(n1277), .B(n1279), .Z(n1169) );
  XOR U1333 ( .A(n1280), .B(n1169), .Z(n1273) );
  XNOR U1334 ( .A(n1274), .B(n1273), .Z(n1264) );
  IV U1335 ( .A(n1264), .Z(n1263) );
  NANDN U1336 ( .A(n1171), .B(n1170), .Z(n1175) );
  OR U1337 ( .A(n1173), .B(n1172), .Z(n1174) );
  AND U1338 ( .A(n1175), .B(n1174), .Z(n1265) );
  XOR U1339 ( .A(n1263), .B(n1265), .Z(n1176) );
  XOR U1340 ( .A(n1266), .B(n1176), .Z(n1259) );
  XNOR U1341 ( .A(n1260), .B(n1259), .Z(n1251) );
  IV U1342 ( .A(n1251), .Z(n1249) );
  NANDN U1343 ( .A(n1178), .B(n1177), .Z(n1182) );
  OR U1344 ( .A(n1180), .B(n1179), .Z(n1181) );
  NAND U1345 ( .A(n1182), .B(n1181), .Z(n1250) );
  XOR U1346 ( .A(n1249), .B(n1250), .Z(n1183) );
  XNOR U1347 ( .A(n1252), .B(n1183), .Z(n1245) );
  XNOR U1348 ( .A(n1246), .B(n1245), .Z(n1522) );
  IV U1349 ( .A(\stack[1][1] ), .Z(n1242) );
  ANDN U1350 ( .B(o[11]), .A(n1242), .Z(n1234) );
  XNOR U1351 ( .A(n1185), .B(n1184), .Z(n1508) );
  ANDN U1352 ( .B(o[9]), .A(n1242), .Z(n1226) );
  XNOR U1353 ( .A(n1187), .B(n1186), .Z(n1495) );
  ANDN U1354 ( .B(o[7]), .A(n1242), .Z(n1215) );
  ANDN U1355 ( .B(o[5]), .A(n1242), .Z(n1204) );
  XOR U1356 ( .A(n1191), .B(n1190), .Z(n1466) );
  ANDN U1357 ( .B(o[3]), .A(n1242), .Z(n1200) );
  ANDN U1358 ( .B(o[2]), .A(n1242), .Z(n1192) );
  NAND U1359 ( .A(\stack[1][1] ), .B(o[1]), .Z(n1449) );
  NAND U1360 ( .A(o[0]), .B(\stack[1][2] ), .Z(n1448) );
  OR U1361 ( .A(n1449), .B(n1448), .Z(n1193) );
  NANDN U1362 ( .A(n1192), .B(n1193), .Z(n1197) );
  XOR U1363 ( .A(n1193), .B(n1192), .Z(n1455) );
  XOR U1364 ( .A(n1195), .B(n1194), .Z(n1454) );
  OR U1365 ( .A(n1455), .B(n1454), .Z(n1196) );
  AND U1366 ( .A(n1197), .B(n1196), .Z(n1201) );
  OR U1367 ( .A(n1200), .B(n1201), .Z(n1203) );
  XNOR U1368 ( .A(n1199), .B(n1198), .Z(n1459) );
  XOR U1369 ( .A(n1201), .B(n1200), .Z(n1458) );
  NANDN U1370 ( .A(n1459), .B(n1458), .Z(n1202) );
  NAND U1371 ( .A(n1203), .B(n1202), .Z(n1469) );
  NAND U1372 ( .A(\stack[1][1] ), .B(o[4]), .Z(n1467) );
  NANDN U1373 ( .A(n1204), .B(n1205), .Z(n1211) );
  XOR U1374 ( .A(n1205), .B(n1204), .Z(n1473) );
  XNOR U1375 ( .A(n1207), .B(n1206), .Z(n1208) );
  XOR U1376 ( .A(n1209), .B(n1208), .Z(n1472) );
  NANDN U1377 ( .A(n1473), .B(n1472), .Z(n1210) );
  NAND U1378 ( .A(n1211), .B(n1210), .Z(n1483) );
  NAND U1379 ( .A(n1480), .B(n1483), .Z(n1214) );
  NOR U1380 ( .A(n1483), .B(n1480), .Z(n1212) );
  NAND U1381 ( .A(\stack[1][1] ), .B(o[6]), .Z(n1481) );
  NANDN U1382 ( .A(n1212), .B(n1481), .Z(n1213) );
  NAND U1383 ( .A(n1214), .B(n1213), .Z(n1216) );
  NANDN U1384 ( .A(n1215), .B(n1216), .Z(n1221) );
  XOR U1385 ( .A(n1216), .B(n1215), .Z(n1487) );
  OR U1386 ( .A(n1487), .B(n1486), .Z(n1220) );
  NAND U1387 ( .A(n1221), .B(n1220), .Z(n1222) );
  NANDN U1388 ( .A(n1495), .B(n1222), .Z(n1225) );
  IV U1389 ( .A(n1222), .Z(n1494) );
  AND U1390 ( .A(n1495), .B(n1494), .Z(n1223) );
  NAND U1391 ( .A(\stack[1][1] ), .B(o[8]), .Z(n1497) );
  NANDN U1392 ( .A(n1223), .B(n1497), .Z(n1224) );
  NAND U1393 ( .A(n1225), .B(n1224), .Z(n1227) );
  NANDN U1394 ( .A(n1226), .B(n1227), .Z(n1233) );
  XOR U1395 ( .A(n1227), .B(n1226), .Z(n1501) );
  XOR U1396 ( .A(n1229), .B(n1228), .Z(n1230) );
  XOR U1397 ( .A(n1231), .B(n1230), .Z(n1500) );
  NANDN U1398 ( .A(n1501), .B(n1500), .Z(n1232) );
  NAND U1399 ( .A(n1233), .B(n1232), .Z(n1511) );
  NAND U1400 ( .A(\stack[1][1] ), .B(o[10]), .Z(n1509) );
  NANDN U1401 ( .A(n1234), .B(n1235), .Z(n1241) );
  XOR U1402 ( .A(n1235), .B(n1234), .Z(n1515) );
  XOR U1403 ( .A(n1237), .B(n1236), .Z(n1238) );
  XOR U1404 ( .A(n1239), .B(n1238), .Z(n1514) );
  NANDN U1405 ( .A(n1515), .B(n1514), .Z(n1240) );
  NAND U1406 ( .A(n1241), .B(n1240), .Z(n1525) );
  NAND U1407 ( .A(\stack[1][1] ), .B(o[12]), .Z(n1523) );
  ANDN U1408 ( .B(o[13]), .A(n1242), .Z(n1318) );
  XOR U1409 ( .A(n1319), .B(n1318), .Z(n1529) );
  NANDN U1410 ( .A(n1244), .B(n1243), .Z(n1248) );
  OR U1411 ( .A(n1246), .B(n1245), .Z(n1247) );
  NAND U1412 ( .A(n1248), .B(n1247), .Z(n1440) );
  AND U1413 ( .A(n1250), .B(n1249), .Z(n1255) );
  ANDN U1414 ( .B(n1251), .A(n1250), .Z(n1253) );
  NANDN U1415 ( .A(n1253), .B(n1252), .Z(n1254) );
  NANDN U1416 ( .A(n1255), .B(n1254), .Z(n1330) );
  ANDN U1417 ( .B(o[11]), .A(n1256), .Z(n1331) );
  XOR U1418 ( .A(n1330), .B(n1331), .Z(n1329) );
  NANDN U1419 ( .A(n1258), .B(n1257), .Z(n1262) );
  OR U1420 ( .A(n1260), .B(n1259), .Z(n1261) );
  NAND U1421 ( .A(n1262), .B(n1261), .Z(n1428) );
  NANDN U1422 ( .A(n1265), .B(n1263), .Z(n1269) );
  AND U1423 ( .A(n1265), .B(n1264), .Z(n1267) );
  NANDN U1424 ( .A(n1267), .B(n1266), .Z(n1268) );
  NAND U1425 ( .A(n1269), .B(n1268), .Z(n1324) );
  ANDN U1426 ( .B(o[9]), .A(n1270), .Z(n1325) );
  XOR U1427 ( .A(n1324), .B(n1325), .Z(n1323) );
  NANDN U1428 ( .A(n1272), .B(n1271), .Z(n1276) );
  OR U1429 ( .A(n1274), .B(n1273), .Z(n1275) );
  NAND U1430 ( .A(n1276), .B(n1275), .Z(n1405) );
  NANDN U1431 ( .A(n1279), .B(n1277), .Z(n1283) );
  AND U1432 ( .A(n1279), .B(n1278), .Z(n1281) );
  NANDN U1433 ( .A(n1281), .B(n1280), .Z(n1282) );
  NAND U1434 ( .A(n1283), .B(n1282), .Z(n1420) );
  NAND U1435 ( .A(\stack[1][7] ), .B(o[7]), .Z(n1852) );
  XNOR U1436 ( .A(n1420), .B(n1852), .Z(n1419) );
  ANDN U1437 ( .B(o[6]), .A(n1284), .Z(n1410) );
  NANDN U1438 ( .A(n1287), .B(n1285), .Z(n1291) );
  AND U1439 ( .A(n1287), .B(n1286), .Z(n1289) );
  NANDN U1440 ( .A(n1289), .B(n1288), .Z(n1290) );
  NAND U1441 ( .A(n1291), .B(n1290), .Z(n1392) );
  ANDN U1442 ( .B(\stack[1][9] ), .A(n1292), .Z(n1393) );
  XOR U1443 ( .A(n1392), .B(n1393), .Z(n1395) );
  NANDN U1444 ( .A(n1294), .B(n1293), .Z(n1298) );
  OR U1445 ( .A(n1296), .B(n1295), .Z(n1297) );
  AND U1446 ( .A(n1298), .B(n1297), .Z(n1378) );
  NAND U1447 ( .A(\stack[1][10] ), .B(o[4]), .Z(n1381) );
  AND U1448 ( .A(o[2]), .B(\stack[1][12] ), .Z(n1338) );
  ANDN U1449 ( .B(n1300), .A(n1299), .Z(n1339) );
  NAND U1450 ( .A(\stack[1][13] ), .B(o[1]), .Z(n1336) );
  AND U1451 ( .A(\stack[1][14] ), .B(o[0]), .Z(n1337) );
  XNOR U1452 ( .A(n1336), .B(n1337), .Z(n1343) );
  OR U1453 ( .A(n1302), .B(n1301), .Z(n1306) );
  OR U1454 ( .A(n1304), .B(n1303), .Z(n1305) );
  AND U1455 ( .A(n1306), .B(n1305), .Z(n1386) );
  NAND U1456 ( .A(\stack[1][11] ), .B(o[3]), .Z(n1387) );
  XOR U1457 ( .A(n1386), .B(n1387), .Z(n1388) );
  XOR U1458 ( .A(n1389), .B(n1388), .Z(n1379) );
  XNOR U1459 ( .A(n1381), .B(n1379), .Z(n1307) );
  XNOR U1460 ( .A(n1378), .B(n1307), .Z(n1394) );
  NANDN U1461 ( .A(n1309), .B(n1308), .Z(n1313) );
  OR U1462 ( .A(n1311), .B(n1310), .Z(n1312) );
  NAND U1463 ( .A(n1313), .B(n1312), .Z(n1413) );
  XOR U1464 ( .A(n1411), .B(n1413), .Z(n1314) );
  XNOR U1465 ( .A(n1410), .B(n1314), .Z(n1418) );
  XNOR U1466 ( .A(n1419), .B(n1418), .Z(n1403) );
  ANDN U1467 ( .B(o[8]), .A(n1315), .Z(n1402) );
  XOR U1468 ( .A(n1403), .B(n1402), .Z(n1404) );
  XOR U1469 ( .A(n1405), .B(n1404), .Z(n1322) );
  ANDN U1470 ( .B(o[10]), .A(n1316), .Z(n1425) );
  XOR U1471 ( .A(n1426), .B(n1425), .Z(n1427) );
  XOR U1472 ( .A(n1428), .B(n1427), .Z(n1328) );
  ANDN U1473 ( .B(o[12]), .A(n1317), .Z(n1437) );
  XOR U1474 ( .A(n1438), .B(n1437), .Z(n1439) );
  XOR U1475 ( .A(n1440), .B(n1439), .Z(n1528) );
  NANDN U1476 ( .A(n1529), .B(n1528), .Z(n1321) );
  ANDN U1477 ( .B(n1319), .A(n1318), .Z(n1320) );
  ANDN U1478 ( .B(n1321), .A(n1320), .Z(n1436) );
  NANDN U1479 ( .A(n1323), .B(n1322), .Z(n1327) );
  NANDN U1480 ( .A(n1325), .B(n1324), .Z(n1326) );
  AND U1481 ( .A(n1327), .B(n1326), .Z(n1335) );
  NANDN U1482 ( .A(n1329), .B(n1328), .Z(n1333) );
  NANDN U1483 ( .A(n1331), .B(n1330), .Z(n1332) );
  NAND U1484 ( .A(n1333), .B(n1332), .Z(n1334) );
  XNOR U1485 ( .A(n1335), .B(n1334), .Z(n1434) );
  ANDN U1486 ( .B(n1337), .A(n1336), .Z(n1341) );
  AND U1487 ( .A(n1339), .B(n1338), .Z(n1340) );
  XNOR U1488 ( .A(n1341), .B(n1340), .Z(n1345) );
  NAND U1489 ( .A(n1343), .B(n1342), .Z(n1344) );
  NAND U1490 ( .A(n1345), .B(n1344), .Z(n1377) );
  AND U1491 ( .A(o[7]), .B(\stack[1][8] ), .Z(n1347) );
  NAND U1492 ( .A(\stack[1][5] ), .B(o[10]), .Z(n1346) );
  XNOR U1493 ( .A(n1347), .B(n1346), .Z(n1351) );
  AND U1494 ( .A(o[11]), .B(\stack[1][4] ), .Z(n1349) );
  NAND U1495 ( .A(\stack[1][3] ), .B(o[12]), .Z(n1348) );
  XNOR U1496 ( .A(n1349), .B(n1348), .Z(n1350) );
  XOR U1497 ( .A(n1351), .B(n1350), .Z(n1359) );
  AND U1498 ( .A(o[9]), .B(\stack[1][6] ), .Z(n1353) );
  NAND U1499 ( .A(\stack[1][11] ), .B(o[4]), .Z(n1352) );
  XNOR U1500 ( .A(n1353), .B(n1352), .Z(n1357) );
  AND U1501 ( .A(o[6]), .B(\stack[1][9] ), .Z(n1355) );
  NAND U1502 ( .A(o[5]), .B(\stack[1][10] ), .Z(n1354) );
  XNOR U1503 ( .A(n1355), .B(n1354), .Z(n1356) );
  XNOR U1504 ( .A(n1357), .B(n1356), .Z(n1358) );
  XNOR U1505 ( .A(n1359), .B(n1358), .Z(n1375) );
  AND U1506 ( .A(o[8]), .B(\stack[1][7] ), .Z(n1361) );
  NAND U1507 ( .A(o[3]), .B(\stack[1][12] ), .Z(n1360) );
  XNOR U1508 ( .A(n1361), .B(n1360), .Z(n1365) );
  AND U1509 ( .A(o[2]), .B(\stack[1][13] ), .Z(n1363) );
  NAND U1510 ( .A(o[0]), .B(\stack[1][15] ), .Z(n1362) );
  XNOR U1511 ( .A(n1363), .B(n1362), .Z(n1364) );
  XOR U1512 ( .A(n1365), .B(n1364), .Z(n1373) );
  AND U1513 ( .A(\stack[1][14] ), .B(o[1]), .Z(n1367) );
  NAND U1514 ( .A(\stack[1][0] ), .B(o[15]), .Z(n1366) );
  XNOR U1515 ( .A(n1367), .B(n1366), .Z(n1371) );
  AND U1516 ( .A(o[13]), .B(\stack[1][2] ), .Z(n1369) );
  NAND U1517 ( .A(\stack[1][1] ), .B(o[14]), .Z(n1368) );
  XNOR U1518 ( .A(n1369), .B(n1368), .Z(n1370) );
  XNOR U1519 ( .A(n1371), .B(n1370), .Z(n1372) );
  XNOR U1520 ( .A(n1373), .B(n1372), .Z(n1374) );
  XNOR U1521 ( .A(n1375), .B(n1374), .Z(n1376) );
  XNOR U1522 ( .A(n1377), .B(n1376), .Z(n1385) );
  NAND U1523 ( .A(n1379), .B(n1378), .Z(n1383) );
  XOR U1524 ( .A(n1379), .B(n1378), .Z(n1380) );
  NANDN U1525 ( .A(n1381), .B(n1380), .Z(n1382) );
  NAND U1526 ( .A(n1383), .B(n1382), .Z(n1384) );
  XNOR U1527 ( .A(n1385), .B(n1384), .Z(n1401) );
  ANDN U1528 ( .B(n1387), .A(n1386), .Z(n1391) );
  ANDN U1529 ( .B(n1389), .A(n1388), .Z(n1390) );
  NOR U1530 ( .A(n1391), .B(n1390), .Z(n1399) );
  NANDN U1531 ( .A(n1393), .B(n1392), .Z(n1397) );
  NANDN U1532 ( .A(n1395), .B(n1394), .Z(n1396) );
  AND U1533 ( .A(n1397), .B(n1396), .Z(n1398) );
  XNOR U1534 ( .A(n1399), .B(n1398), .Z(n1400) );
  XNOR U1535 ( .A(n1401), .B(n1400), .Z(n1409) );
  NAND U1536 ( .A(n1403), .B(n1402), .Z(n1407) );
  NANDN U1537 ( .A(n1405), .B(n1404), .Z(n1406) );
  AND U1538 ( .A(n1407), .B(n1406), .Z(n1408) );
  XNOR U1539 ( .A(n1409), .B(n1408), .Z(n1417) );
  NAND U1540 ( .A(n1411), .B(n1410), .Z(n1415) );
  XOR U1541 ( .A(n1411), .B(n1410), .Z(n1412) );
  NANDN U1542 ( .A(n1413), .B(n1412), .Z(n1414) );
  AND U1543 ( .A(n1415), .B(n1414), .Z(n1416) );
  XNOR U1544 ( .A(n1417), .B(n1416), .Z(n1424) );
  OR U1545 ( .A(n1419), .B(n1418), .Z(n1422) );
  NAND U1546 ( .A(n1852), .B(n1420), .Z(n1421) );
  NAND U1547 ( .A(n1422), .B(n1421), .Z(n1423) );
  XNOR U1548 ( .A(n1424), .B(n1423), .Z(n1432) );
  NAND U1549 ( .A(n1426), .B(n1425), .Z(n1430) );
  NANDN U1550 ( .A(n1428), .B(n1427), .Z(n1429) );
  AND U1551 ( .A(n1430), .B(n1429), .Z(n1431) );
  XNOR U1552 ( .A(n1432), .B(n1431), .Z(n1433) );
  XNOR U1553 ( .A(n1434), .B(n1433), .Z(n1435) );
  XNOR U1554 ( .A(n1436), .B(n1435), .Z(n1444) );
  NAND U1555 ( .A(n1438), .B(n1437), .Z(n1442) );
  NANDN U1556 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U1557 ( .A(n1442), .B(n1441), .Z(n1443) );
  XNOR U1558 ( .A(n1444), .B(n1443), .Z(n1535) );
  NAND U1559 ( .A(\stack[1][0] ), .B(o[14]), .Z(n1530) );
  IV U1560 ( .A(\stack[1][0] ), .Z(n1577) );
  ANDN U1561 ( .B(o[13]), .A(n1577), .Z(n1520) );
  ANDN U1562 ( .B(o[11]), .A(n1577), .Z(n1506) );
  ANDN U1563 ( .B(o[9]), .A(n1577), .Z(n1492) );
  ANDN U1564 ( .B(o[7]), .A(n1577), .Z(n1478) );
  ANDN U1565 ( .B(o[5]), .A(n1577), .Z(n1464) );
  ANDN U1566 ( .B(o[3]), .A(n1577), .Z(n1452) );
  ANDN U1567 ( .B(o[2]), .A(n1577), .Z(n1446) );
  ANDN U1568 ( .B(o[1]), .A(n1577), .Z(n2080) );
  ANDN U1569 ( .B(\stack[1][1] ), .A(n1445), .Z(n2081) );
  AND U1570 ( .A(n2080), .B(n2081), .Z(n1447) );
  OR U1571 ( .A(n1446), .B(n1447), .Z(n1451) );
  XNOR U1572 ( .A(n1447), .B(n1446), .Z(n2042) );
  XOR U1573 ( .A(n1449), .B(n1448), .Z(n2043) );
  OR U1574 ( .A(n2042), .B(n2043), .Z(n1450) );
  AND U1575 ( .A(n1451), .B(n1450), .Z(n1453) );
  OR U1576 ( .A(n1452), .B(n1453), .Z(n1457) );
  XNOR U1577 ( .A(n1453), .B(n1452), .Z(n2005) );
  XOR U1578 ( .A(n1455), .B(n1454), .Z(n2006) );
  NANDN U1579 ( .A(n2005), .B(n2006), .Z(n1456) );
  AND U1580 ( .A(n1457), .B(n1456), .Z(n1461) );
  NANDN U1581 ( .A(n1461), .B(n1460), .Z(n1463) );
  NAND U1582 ( .A(\stack[1][0] ), .B(o[4]), .Z(n1462) );
  NANDN U1583 ( .A(n1965), .B(n1462), .Z(n1963) );
  NAND U1584 ( .A(n1463), .B(n1963), .Z(n1465) );
  NANDN U1585 ( .A(n1464), .B(n1465), .Z(n1471) );
  XOR U1586 ( .A(n1465), .B(n1464), .Z(n1925) );
  XOR U1587 ( .A(n1467), .B(n1466), .Z(n1468) );
  XOR U1588 ( .A(n1469), .B(n1468), .Z(n1926) );
  NANDN U1589 ( .A(n1925), .B(n1926), .Z(n1470) );
  AND U1590 ( .A(n1471), .B(n1470), .Z(n1475) );
  NANDN U1591 ( .A(n1475), .B(n1474), .Z(n1477) );
  NAND U1592 ( .A(\stack[1][0] ), .B(o[6]), .Z(n1476) );
  NANDN U1593 ( .A(n1887), .B(n1476), .Z(n1885) );
  NAND U1594 ( .A(n1477), .B(n1885), .Z(n1479) );
  NANDN U1595 ( .A(n1478), .B(n1479), .Z(n1485) );
  XOR U1596 ( .A(n1479), .B(n1478), .Z(n1847) );
  XOR U1597 ( .A(n1481), .B(n1480), .Z(n1482) );
  XOR U1598 ( .A(n1483), .B(n1482), .Z(n1848) );
  NANDN U1599 ( .A(n1847), .B(n1848), .Z(n1484) );
  AND U1600 ( .A(n1485), .B(n1484), .Z(n1489) );
  XOR U1601 ( .A(n1487), .B(n1486), .Z(n1488) );
  NANDN U1602 ( .A(n1489), .B(n1488), .Z(n1491) );
  NAND U1603 ( .A(\stack[1][0] ), .B(o[8]), .Z(n1490) );
  NANDN U1604 ( .A(n1809), .B(n1490), .Z(n1807) );
  NAND U1605 ( .A(n1491), .B(n1807), .Z(n1493) );
  NANDN U1606 ( .A(n1492), .B(n1493), .Z(n1499) );
  XOR U1607 ( .A(n1493), .B(n1492), .Z(n1774) );
  XOR U1608 ( .A(n1495), .B(n1494), .Z(n1496) );
  XNOR U1609 ( .A(n1497), .B(n1496), .Z(n1773) );
  OR U1610 ( .A(n1774), .B(n1773), .Z(n1498) );
  AND U1611 ( .A(n1499), .B(n1498), .Z(n1503) );
  NANDN U1612 ( .A(n1503), .B(n1502), .Z(n1505) );
  NAND U1613 ( .A(\stack[1][0] ), .B(o[10]), .Z(n1504) );
  NANDN U1614 ( .A(n1732), .B(n1504), .Z(n1730) );
  NAND U1615 ( .A(n1505), .B(n1730), .Z(n1507) );
  NANDN U1616 ( .A(n1506), .B(n1507), .Z(n1513) );
  XOR U1617 ( .A(n1507), .B(n1506), .Z(n1697) );
  XNOR U1618 ( .A(n1509), .B(n1508), .Z(n1510) );
  XOR U1619 ( .A(n1511), .B(n1510), .Z(n1696) );
  NANDN U1620 ( .A(n1697), .B(n1696), .Z(n1512) );
  AND U1621 ( .A(n1513), .B(n1512), .Z(n1517) );
  NANDN U1622 ( .A(n1517), .B(n1516), .Z(n1519) );
  NAND U1623 ( .A(\stack[1][0] ), .B(o[12]), .Z(n1518) );
  NANDN U1624 ( .A(n1655), .B(n1518), .Z(n1653) );
  NAND U1625 ( .A(n1519), .B(n1653), .Z(n1521) );
  NANDN U1626 ( .A(n1520), .B(n1521), .Z(n1527) );
  XOR U1627 ( .A(n1521), .B(n1520), .Z(n1620) );
  XNOR U1628 ( .A(n1523), .B(n1522), .Z(n1524) );
  XOR U1629 ( .A(n1525), .B(n1524), .Z(n1619) );
  NANDN U1630 ( .A(n1620), .B(n1619), .Z(n1526) );
  AND U1631 ( .A(n1527), .B(n1526), .Z(n1531) );
  NAND U1632 ( .A(n1530), .B(n1578), .Z(n1575) );
  ANDN U1633 ( .B(n1532), .A(n1531), .Z(n1533) );
  ANDN U1634 ( .B(n1575), .A(n1533), .Z(n1534) );
  XNOR U1635 ( .A(n1535), .B(n1534), .Z(n1536) );
  NAND U1636 ( .A(opcode[1]), .B(opcode[0]), .Z(n1544) );
  ANDN U1637 ( .B(n851), .A(n1544), .Z(n2092) );
  NAND U1638 ( .A(n1536), .B(n2092), .Z(n1539) );
  NAND U1639 ( .A(n796), .B(x[15]), .Z(n1537) );
  AND U1640 ( .A(n1539), .B(n1538), .Z(n1543) );
  XNOR U1641 ( .A(opcode[2]), .B(opcode[1]), .Z(n1540) );
  AND U1642 ( .A(n1541), .B(n1540), .Z(n2090) );
  NAND U1643 ( .A(n2090), .B(o[15]), .Z(n1542) );
  AND U1644 ( .A(n1543), .B(n1542), .Z(n1548) );
  AND U1645 ( .A(opcode[2]), .B(opcode[1]), .Z(n2093) );
  NAND U1646 ( .A(o[15]), .B(n2093), .Z(n1545) );
  NANDN U1647 ( .A(n1544), .B(opcode[2]), .Z(n2096) );
  NAND U1648 ( .A(n1545), .B(n2096), .Z(n1546) );
  NAND U1649 ( .A(n1546), .B(\stack[1][15] ), .Z(n1547) );
  NAND U1650 ( .A(n1548), .B(n1547), .Z(n535) );
  NAND U1651 ( .A(n796), .B(\stack[6][14] ), .Z(n1550) );
  NAND U1652 ( .A(n795), .B(\stack[7][14] ), .Z(n1549) );
  NAND U1653 ( .A(n1550), .B(n1549), .Z(n536) );
  NAND U1654 ( .A(n796), .B(\stack[5][14] ), .Z(n1552) );
  NANDN U1655 ( .A(n2084), .B(\stack[7][14] ), .Z(n1551) );
  AND U1656 ( .A(n1552), .B(n1551), .Z(n1554) );
  NANDN U1657 ( .A(n2087), .B(\stack[6][14] ), .Z(n1553) );
  NAND U1658 ( .A(n1554), .B(n1553), .Z(n537) );
  NAND U1659 ( .A(n796), .B(\stack[4][14] ), .Z(n1556) );
  NANDN U1660 ( .A(n2084), .B(\stack[6][14] ), .Z(n1555) );
  AND U1661 ( .A(n1556), .B(n1555), .Z(n1558) );
  NANDN U1662 ( .A(n2087), .B(\stack[5][14] ), .Z(n1557) );
  NAND U1663 ( .A(n1558), .B(n1557), .Z(n538) );
  NAND U1664 ( .A(n796), .B(\stack[3][14] ), .Z(n1560) );
  NANDN U1665 ( .A(n2084), .B(\stack[5][14] ), .Z(n1559) );
  AND U1666 ( .A(n1560), .B(n1559), .Z(n1562) );
  NANDN U1667 ( .A(n2087), .B(\stack[4][14] ), .Z(n1561) );
  NAND U1668 ( .A(n1562), .B(n1561), .Z(n539) );
  NAND U1669 ( .A(n796), .B(\stack[2][14] ), .Z(n1564) );
  NANDN U1670 ( .A(n2084), .B(\stack[4][14] ), .Z(n1563) );
  AND U1671 ( .A(n1564), .B(n1563), .Z(n1566) );
  NANDN U1672 ( .A(n2087), .B(\stack[3][14] ), .Z(n1565) );
  NAND U1673 ( .A(n1566), .B(n1565), .Z(n540) );
  NAND U1674 ( .A(n796), .B(\stack[1][14] ), .Z(n1568) );
  NANDN U1675 ( .A(n2084), .B(\stack[3][14] ), .Z(n1567) );
  AND U1676 ( .A(n1568), .B(n1567), .Z(n1570) );
  NANDN U1677 ( .A(n2087), .B(\stack[2][14] ), .Z(n1569) );
  NAND U1678 ( .A(n1570), .B(n1569), .Z(n541) );
  NAND U1679 ( .A(n796), .B(o[14]), .Z(n1572) );
  NANDN U1680 ( .A(n2084), .B(\stack[2][14] ), .Z(n1571) );
  AND U1681 ( .A(n1572), .B(n1571), .Z(n1574) );
  NANDN U1682 ( .A(n2087), .B(\stack[1][14] ), .Z(n1573) );
  NAND U1683 ( .A(n1574), .B(n1573), .Z(n542) );
  NANDN U1684 ( .A(n1575), .B(n2092), .Z(n1576) );
  IV U1685 ( .A(n2090), .Z(n2083) );
  NAND U1686 ( .A(\stack[1][14] ), .B(n2093), .Z(n1580) );
  ANDN U1687 ( .B(n2092), .A(n1577), .Z(n2082) );
  NANDN U1688 ( .A(n1578), .B(n2082), .Z(n1579) );
  AND U1689 ( .A(n1580), .B(n1579), .Z(n1581) );
  NAND U1690 ( .A(n2083), .B(n1581), .Z(n1582) );
  NAND U1691 ( .A(n1582), .B(o[14]), .Z(n1586) );
  NAND U1692 ( .A(n796), .B(x[14]), .Z(n1584) );
  NANDN U1693 ( .A(n2096), .B(\stack[1][14] ), .Z(n1583) );
  NAND U1694 ( .A(n1584), .B(n1583), .Z(n1585) );
  ANDN U1695 ( .B(n1586), .A(n1585), .Z(n1587) );
  NAND U1696 ( .A(n1588), .B(n1587), .Z(n543) );
  NAND U1697 ( .A(n796), .B(\stack[6][13] ), .Z(n1590) );
  NAND U1698 ( .A(n795), .B(\stack[7][13] ), .Z(n1589) );
  NAND U1699 ( .A(n1590), .B(n1589), .Z(n544) );
  NAND U1700 ( .A(n796), .B(\stack[5][13] ), .Z(n1592) );
  NANDN U1701 ( .A(n2084), .B(\stack[7][13] ), .Z(n1591) );
  AND U1702 ( .A(n1592), .B(n1591), .Z(n1594) );
  NANDN U1703 ( .A(n2087), .B(\stack[6][13] ), .Z(n1593) );
  NAND U1704 ( .A(n1594), .B(n1593), .Z(n545) );
  NAND U1705 ( .A(n796), .B(\stack[4][13] ), .Z(n1596) );
  NANDN U1706 ( .A(n2084), .B(\stack[6][13] ), .Z(n1595) );
  AND U1707 ( .A(n1596), .B(n1595), .Z(n1598) );
  NANDN U1708 ( .A(n2087), .B(\stack[5][13] ), .Z(n1597) );
  NAND U1709 ( .A(n1598), .B(n1597), .Z(n546) );
  NAND U1710 ( .A(n796), .B(\stack[3][13] ), .Z(n1600) );
  NANDN U1711 ( .A(n2084), .B(\stack[5][13] ), .Z(n1599) );
  AND U1712 ( .A(n1600), .B(n1599), .Z(n1602) );
  NANDN U1713 ( .A(n2087), .B(\stack[4][13] ), .Z(n1601) );
  NAND U1714 ( .A(n1602), .B(n1601), .Z(n547) );
  NAND U1715 ( .A(n796), .B(\stack[2][13] ), .Z(n1604) );
  NANDN U1716 ( .A(n2084), .B(\stack[4][13] ), .Z(n1603) );
  AND U1717 ( .A(n1604), .B(n1603), .Z(n1606) );
  NANDN U1718 ( .A(n2087), .B(\stack[3][13] ), .Z(n1605) );
  NAND U1719 ( .A(n1606), .B(n1605), .Z(n548) );
  NAND U1720 ( .A(n796), .B(\stack[1][13] ), .Z(n1608) );
  NANDN U1721 ( .A(n2084), .B(\stack[3][13] ), .Z(n1607) );
  AND U1722 ( .A(n1608), .B(n1607), .Z(n1610) );
  NANDN U1723 ( .A(n2087), .B(\stack[2][13] ), .Z(n1609) );
  NAND U1724 ( .A(n1610), .B(n1609), .Z(n549) );
  NAND U1725 ( .A(n796), .B(o[13]), .Z(n1612) );
  NANDN U1726 ( .A(n2084), .B(\stack[2][13] ), .Z(n1611) );
  AND U1727 ( .A(n1612), .B(n1611), .Z(n1614) );
  NANDN U1728 ( .A(n2087), .B(\stack[1][13] ), .Z(n1613) );
  NAND U1729 ( .A(n1614), .B(n1613), .Z(n550) );
  NAND U1730 ( .A(\stack[1][13] ), .B(n2093), .Z(n1615) );
  NAND U1731 ( .A(n2083), .B(n1615), .Z(n1616) );
  AND U1732 ( .A(n1616), .B(o[13]), .Z(n1625) );
  NAND U1733 ( .A(n796), .B(x[13]), .Z(n1618) );
  NANDN U1734 ( .A(n2096), .B(\stack[1][13] ), .Z(n1617) );
  NAND U1735 ( .A(n1618), .B(n1617), .Z(n1623) );
  XOR U1736 ( .A(n1620), .B(n1619), .Z(n1621) );
  NAND U1737 ( .A(n1621), .B(n2092), .Z(n1622) );
  NANDN U1738 ( .A(n1623), .B(n1622), .Z(n1624) );
  NOR U1739 ( .A(n1625), .B(n1624), .Z(n1626) );
  NAND U1740 ( .A(n796), .B(\stack[6][12] ), .Z(n1628) );
  NAND U1741 ( .A(n795), .B(\stack[7][12] ), .Z(n1627) );
  NAND U1742 ( .A(n1628), .B(n1627), .Z(n552) );
  NAND U1743 ( .A(n796), .B(\stack[5][12] ), .Z(n1630) );
  NANDN U1744 ( .A(n2084), .B(\stack[7][12] ), .Z(n1629) );
  AND U1745 ( .A(n1630), .B(n1629), .Z(n1632) );
  NANDN U1746 ( .A(n2087), .B(\stack[6][12] ), .Z(n1631) );
  NAND U1747 ( .A(n1632), .B(n1631), .Z(n553) );
  NAND U1748 ( .A(n796), .B(\stack[4][12] ), .Z(n1634) );
  NANDN U1749 ( .A(n2084), .B(\stack[6][12] ), .Z(n1633) );
  AND U1750 ( .A(n1634), .B(n1633), .Z(n1636) );
  NANDN U1751 ( .A(n2087), .B(\stack[5][12] ), .Z(n1635) );
  NAND U1752 ( .A(n1636), .B(n1635), .Z(n554) );
  NAND U1753 ( .A(n796), .B(\stack[3][12] ), .Z(n1638) );
  NANDN U1754 ( .A(n2084), .B(\stack[5][12] ), .Z(n1637) );
  AND U1755 ( .A(n1638), .B(n1637), .Z(n1640) );
  NANDN U1756 ( .A(n2087), .B(\stack[4][12] ), .Z(n1639) );
  NAND U1757 ( .A(n1640), .B(n1639), .Z(n555) );
  NAND U1758 ( .A(n796), .B(\stack[2][12] ), .Z(n1642) );
  NANDN U1759 ( .A(n2084), .B(\stack[4][12] ), .Z(n1641) );
  AND U1760 ( .A(n1642), .B(n1641), .Z(n1644) );
  NANDN U1761 ( .A(n2087), .B(\stack[3][12] ), .Z(n1643) );
  NAND U1762 ( .A(n1644), .B(n1643), .Z(n556) );
  NAND U1763 ( .A(n796), .B(\stack[1][12] ), .Z(n1646) );
  NANDN U1764 ( .A(n2084), .B(\stack[3][12] ), .Z(n1645) );
  AND U1765 ( .A(n1646), .B(n1645), .Z(n1648) );
  NANDN U1766 ( .A(n2087), .B(\stack[2][12] ), .Z(n1647) );
  NAND U1767 ( .A(n1648), .B(n1647), .Z(n557) );
  NAND U1768 ( .A(n796), .B(o[12]), .Z(n1650) );
  NANDN U1769 ( .A(n2084), .B(\stack[2][12] ), .Z(n1649) );
  AND U1770 ( .A(n1650), .B(n1649), .Z(n1652) );
  NANDN U1771 ( .A(n2087), .B(\stack[1][12] ), .Z(n1651) );
  NAND U1772 ( .A(n1652), .B(n1651), .Z(n558) );
  NANDN U1773 ( .A(n1653), .B(n2092), .Z(n1654) );
  NAND U1774 ( .A(\stack[1][12] ), .B(n2093), .Z(n1657) );
  NAND U1775 ( .A(n1655), .B(n2082), .Z(n1656) );
  AND U1776 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U1777 ( .A(n2083), .B(n1658), .Z(n1659) );
  NAND U1778 ( .A(n1659), .B(o[12]), .Z(n1663) );
  NAND U1779 ( .A(n796), .B(x[12]), .Z(n1661) );
  NANDN U1780 ( .A(n2096), .B(\stack[1][12] ), .Z(n1660) );
  NAND U1781 ( .A(n1661), .B(n1660), .Z(n1662) );
  ANDN U1782 ( .B(n1663), .A(n1662), .Z(n1664) );
  NAND U1783 ( .A(n1665), .B(n1664), .Z(n559) );
  NAND U1784 ( .A(n796), .B(\stack[6][11] ), .Z(n1667) );
  NAND U1785 ( .A(n795), .B(\stack[7][11] ), .Z(n1666) );
  NAND U1786 ( .A(n1667), .B(n1666), .Z(n560) );
  NAND U1787 ( .A(n796), .B(\stack[5][11] ), .Z(n1669) );
  NANDN U1788 ( .A(n2084), .B(\stack[7][11] ), .Z(n1668) );
  AND U1789 ( .A(n1669), .B(n1668), .Z(n1671) );
  NANDN U1790 ( .A(n2087), .B(\stack[6][11] ), .Z(n1670) );
  NAND U1791 ( .A(n1671), .B(n1670), .Z(n561) );
  NAND U1792 ( .A(n796), .B(\stack[4][11] ), .Z(n1673) );
  NANDN U1793 ( .A(n2084), .B(\stack[6][11] ), .Z(n1672) );
  AND U1794 ( .A(n1673), .B(n1672), .Z(n1675) );
  NANDN U1795 ( .A(n2087), .B(\stack[5][11] ), .Z(n1674) );
  NAND U1796 ( .A(n1675), .B(n1674), .Z(n562) );
  NAND U1797 ( .A(n796), .B(\stack[3][11] ), .Z(n1677) );
  NANDN U1798 ( .A(n2084), .B(\stack[5][11] ), .Z(n1676) );
  AND U1799 ( .A(n1677), .B(n1676), .Z(n1679) );
  NANDN U1800 ( .A(n2087), .B(\stack[4][11] ), .Z(n1678) );
  NAND U1801 ( .A(n1679), .B(n1678), .Z(n563) );
  NAND U1802 ( .A(n796), .B(\stack[2][11] ), .Z(n1681) );
  NANDN U1803 ( .A(n2084), .B(\stack[4][11] ), .Z(n1680) );
  AND U1804 ( .A(n1681), .B(n1680), .Z(n1683) );
  NANDN U1805 ( .A(n2087), .B(\stack[3][11] ), .Z(n1682) );
  NAND U1806 ( .A(n1683), .B(n1682), .Z(n564) );
  NAND U1807 ( .A(\stack[1][11] ), .B(n796), .Z(n1685) );
  NANDN U1808 ( .A(n2084), .B(\stack[3][11] ), .Z(n1684) );
  AND U1809 ( .A(n1685), .B(n1684), .Z(n1687) );
  NANDN U1810 ( .A(n2087), .B(\stack[2][11] ), .Z(n1686) );
  NAND U1811 ( .A(n1687), .B(n1686), .Z(n565) );
  NAND U1812 ( .A(n796), .B(o[11]), .Z(n1689) );
  NANDN U1813 ( .A(n2084), .B(\stack[2][11] ), .Z(n1688) );
  AND U1814 ( .A(n1689), .B(n1688), .Z(n1691) );
  NANDN U1815 ( .A(n2087), .B(\stack[1][11] ), .Z(n1690) );
  NAND U1816 ( .A(n1691), .B(n1690), .Z(n566) );
  NAND U1817 ( .A(\stack[1][11] ), .B(n2093), .Z(n1692) );
  NAND U1818 ( .A(n2083), .B(n1692), .Z(n1693) );
  AND U1819 ( .A(n1693), .B(o[11]), .Z(n1702) );
  NAND U1820 ( .A(n796), .B(x[11]), .Z(n1695) );
  NANDN U1821 ( .A(n2096), .B(\stack[1][11] ), .Z(n1694) );
  NAND U1822 ( .A(n1695), .B(n1694), .Z(n1700) );
  XOR U1823 ( .A(n1697), .B(n1696), .Z(n1698) );
  NAND U1824 ( .A(n1698), .B(n2092), .Z(n1699) );
  NANDN U1825 ( .A(n1700), .B(n1699), .Z(n1701) );
  NOR U1826 ( .A(n1702), .B(n1701), .Z(n1703) );
  NAND U1827 ( .A(n796), .B(\stack[6][10] ), .Z(n1705) );
  NAND U1828 ( .A(n795), .B(\stack[7][10] ), .Z(n1704) );
  NAND U1829 ( .A(n1705), .B(n1704), .Z(n568) );
  NAND U1830 ( .A(n796), .B(\stack[5][10] ), .Z(n1707) );
  NANDN U1831 ( .A(n2084), .B(\stack[7][10] ), .Z(n1706) );
  AND U1832 ( .A(n1707), .B(n1706), .Z(n1709) );
  NANDN U1833 ( .A(n2087), .B(\stack[6][10] ), .Z(n1708) );
  NAND U1834 ( .A(n1709), .B(n1708), .Z(n569) );
  NAND U1835 ( .A(n796), .B(\stack[4][10] ), .Z(n1711) );
  NANDN U1836 ( .A(n2084), .B(\stack[6][10] ), .Z(n1710) );
  AND U1837 ( .A(n1711), .B(n1710), .Z(n1713) );
  NANDN U1838 ( .A(n2087), .B(\stack[5][10] ), .Z(n1712) );
  NAND U1839 ( .A(n1713), .B(n1712), .Z(n570) );
  NAND U1840 ( .A(n796), .B(\stack[3][10] ), .Z(n1715) );
  NANDN U1841 ( .A(n2084), .B(\stack[5][10] ), .Z(n1714) );
  AND U1842 ( .A(n1715), .B(n1714), .Z(n1717) );
  NANDN U1843 ( .A(n2087), .B(\stack[4][10] ), .Z(n1716) );
  NAND U1844 ( .A(n1717), .B(n1716), .Z(n571) );
  NAND U1845 ( .A(n796), .B(\stack[2][10] ), .Z(n1719) );
  NANDN U1846 ( .A(n2084), .B(\stack[4][10] ), .Z(n1718) );
  AND U1847 ( .A(n1719), .B(n1718), .Z(n1721) );
  NANDN U1848 ( .A(n2087), .B(\stack[3][10] ), .Z(n1720) );
  NAND U1849 ( .A(n1721), .B(n1720), .Z(n572) );
  NAND U1850 ( .A(\stack[1][10] ), .B(n796), .Z(n1723) );
  NANDN U1851 ( .A(n2084), .B(\stack[3][10] ), .Z(n1722) );
  AND U1852 ( .A(n1723), .B(n1722), .Z(n1725) );
  NANDN U1853 ( .A(n2087), .B(\stack[2][10] ), .Z(n1724) );
  NAND U1854 ( .A(n1725), .B(n1724), .Z(n573) );
  NAND U1855 ( .A(n796), .B(o[10]), .Z(n1727) );
  NANDN U1856 ( .A(n2084), .B(\stack[2][10] ), .Z(n1726) );
  AND U1857 ( .A(n1727), .B(n1726), .Z(n1729) );
  NANDN U1858 ( .A(n2087), .B(\stack[1][10] ), .Z(n1728) );
  NAND U1859 ( .A(n1729), .B(n1728), .Z(n574) );
  NANDN U1860 ( .A(n1730), .B(n2092), .Z(n1731) );
  NAND U1861 ( .A(\stack[1][10] ), .B(n2093), .Z(n1734) );
  NAND U1862 ( .A(n2082), .B(n1732), .Z(n1733) );
  AND U1863 ( .A(n1734), .B(n1733), .Z(n1735) );
  NAND U1864 ( .A(n2083), .B(n1735), .Z(n1736) );
  NAND U1865 ( .A(n1736), .B(o[10]), .Z(n1740) );
  NAND U1866 ( .A(n796), .B(x[10]), .Z(n1738) );
  NANDN U1867 ( .A(n2096), .B(\stack[1][10] ), .Z(n1737) );
  NAND U1868 ( .A(n1738), .B(n1737), .Z(n1739) );
  ANDN U1869 ( .B(n1740), .A(n1739), .Z(n1741) );
  NAND U1870 ( .A(n1742), .B(n1741), .Z(n575) );
  NAND U1871 ( .A(n796), .B(\stack[6][9] ), .Z(n1744) );
  NAND U1872 ( .A(n795), .B(\stack[7][9] ), .Z(n1743) );
  NAND U1873 ( .A(n1744), .B(n1743), .Z(n576) );
  NAND U1874 ( .A(n796), .B(\stack[5][9] ), .Z(n1746) );
  NANDN U1875 ( .A(n2084), .B(\stack[7][9] ), .Z(n1745) );
  AND U1876 ( .A(n1746), .B(n1745), .Z(n1748) );
  NANDN U1877 ( .A(n2087), .B(\stack[6][9] ), .Z(n1747) );
  NAND U1878 ( .A(n1748), .B(n1747), .Z(n577) );
  NAND U1879 ( .A(n796), .B(\stack[4][9] ), .Z(n1750) );
  NANDN U1880 ( .A(n2084), .B(\stack[6][9] ), .Z(n1749) );
  AND U1881 ( .A(n1750), .B(n1749), .Z(n1752) );
  NANDN U1882 ( .A(n2087), .B(\stack[5][9] ), .Z(n1751) );
  NAND U1883 ( .A(n1752), .B(n1751), .Z(n578) );
  NAND U1884 ( .A(n796), .B(\stack[3][9] ), .Z(n1754) );
  NANDN U1885 ( .A(n2084), .B(\stack[5][9] ), .Z(n1753) );
  AND U1886 ( .A(n1754), .B(n1753), .Z(n1756) );
  NANDN U1887 ( .A(n2087), .B(\stack[4][9] ), .Z(n1755) );
  NAND U1888 ( .A(n1756), .B(n1755), .Z(n579) );
  NAND U1889 ( .A(n796), .B(\stack[2][9] ), .Z(n1758) );
  NANDN U1890 ( .A(n2084), .B(\stack[4][9] ), .Z(n1757) );
  AND U1891 ( .A(n1758), .B(n1757), .Z(n1760) );
  NANDN U1892 ( .A(n2087), .B(\stack[3][9] ), .Z(n1759) );
  NAND U1893 ( .A(n1760), .B(n1759), .Z(n580) );
  NAND U1894 ( .A(\stack[1][9] ), .B(n796), .Z(n1762) );
  NANDN U1895 ( .A(n2084), .B(\stack[3][9] ), .Z(n1761) );
  AND U1896 ( .A(n1762), .B(n1761), .Z(n1764) );
  NANDN U1897 ( .A(n2087), .B(\stack[2][9] ), .Z(n1763) );
  NAND U1898 ( .A(n1764), .B(n1763), .Z(n581) );
  NAND U1899 ( .A(n796), .B(o[9]), .Z(n1766) );
  NANDN U1900 ( .A(n2084), .B(\stack[2][9] ), .Z(n1765) );
  AND U1901 ( .A(n1766), .B(n1765), .Z(n1768) );
  NANDN U1902 ( .A(n2087), .B(\stack[1][9] ), .Z(n1767) );
  NAND U1903 ( .A(n1768), .B(n1767), .Z(n582) );
  NAND U1904 ( .A(\stack[1][9] ), .B(n2093), .Z(n1769) );
  NAND U1905 ( .A(n2083), .B(n1769), .Z(n1770) );
  AND U1906 ( .A(n1770), .B(o[9]), .Z(n1779) );
  NAND U1907 ( .A(n796), .B(x[9]), .Z(n1772) );
  NANDN U1908 ( .A(n2096), .B(\stack[1][9] ), .Z(n1771) );
  NAND U1909 ( .A(n1772), .B(n1771), .Z(n1777) );
  XNOR U1910 ( .A(n1774), .B(n1773), .Z(n1775) );
  NAND U1911 ( .A(n1775), .B(n2092), .Z(n1776) );
  NANDN U1912 ( .A(n1777), .B(n1776), .Z(n1778) );
  NOR U1913 ( .A(n1779), .B(n1778), .Z(n1780) );
  NAND U1914 ( .A(n796), .B(\stack[6][8] ), .Z(n1782) );
  NAND U1915 ( .A(n795), .B(\stack[7][8] ), .Z(n1781) );
  NAND U1916 ( .A(n1782), .B(n1781), .Z(n584) );
  NAND U1917 ( .A(n796), .B(\stack[5][8] ), .Z(n1784) );
  NANDN U1918 ( .A(n2084), .B(\stack[7][8] ), .Z(n1783) );
  AND U1919 ( .A(n1784), .B(n1783), .Z(n1786) );
  NANDN U1920 ( .A(n2087), .B(\stack[6][8] ), .Z(n1785) );
  NAND U1921 ( .A(n1786), .B(n1785), .Z(n585) );
  NAND U1922 ( .A(n796), .B(\stack[4][8] ), .Z(n1788) );
  NANDN U1923 ( .A(n2084), .B(\stack[6][8] ), .Z(n1787) );
  AND U1924 ( .A(n1788), .B(n1787), .Z(n1790) );
  NANDN U1925 ( .A(n2087), .B(\stack[5][8] ), .Z(n1789) );
  NAND U1926 ( .A(n1790), .B(n1789), .Z(n586) );
  NAND U1927 ( .A(n796), .B(\stack[3][8] ), .Z(n1792) );
  NANDN U1928 ( .A(n2084), .B(\stack[5][8] ), .Z(n1791) );
  AND U1929 ( .A(n1792), .B(n1791), .Z(n1794) );
  NANDN U1930 ( .A(n2087), .B(\stack[4][8] ), .Z(n1793) );
  NAND U1931 ( .A(n1794), .B(n1793), .Z(n587) );
  NAND U1932 ( .A(n796), .B(\stack[2][8] ), .Z(n1796) );
  NANDN U1933 ( .A(n2084), .B(\stack[4][8] ), .Z(n1795) );
  AND U1934 ( .A(n1796), .B(n1795), .Z(n1798) );
  NANDN U1935 ( .A(n2087), .B(\stack[3][8] ), .Z(n1797) );
  NAND U1936 ( .A(n1798), .B(n1797), .Z(n588) );
  NAND U1937 ( .A(\stack[1][8] ), .B(n796), .Z(n1800) );
  NANDN U1938 ( .A(n2084), .B(\stack[3][8] ), .Z(n1799) );
  AND U1939 ( .A(n1800), .B(n1799), .Z(n1802) );
  NANDN U1940 ( .A(n2087), .B(\stack[2][8] ), .Z(n1801) );
  NAND U1941 ( .A(n1802), .B(n1801), .Z(n589) );
  NAND U1942 ( .A(n796), .B(o[8]), .Z(n1804) );
  NANDN U1943 ( .A(n2084), .B(\stack[2][8] ), .Z(n1803) );
  AND U1944 ( .A(n1804), .B(n1803), .Z(n1806) );
  NANDN U1945 ( .A(n2087), .B(\stack[1][8] ), .Z(n1805) );
  NAND U1946 ( .A(n1806), .B(n1805), .Z(n590) );
  NANDN U1947 ( .A(n1807), .B(n2092), .Z(n1808) );
  NAND U1948 ( .A(\stack[1][8] ), .B(n2093), .Z(n1811) );
  NAND U1949 ( .A(n2082), .B(n1809), .Z(n1810) );
  AND U1950 ( .A(n1811), .B(n1810), .Z(n1812) );
  NAND U1951 ( .A(n2083), .B(n1812), .Z(n1813) );
  NAND U1952 ( .A(n1813), .B(o[8]), .Z(n1817) );
  NAND U1953 ( .A(n796), .B(x[8]), .Z(n1815) );
  NANDN U1954 ( .A(n2096), .B(\stack[1][8] ), .Z(n1814) );
  NAND U1955 ( .A(n1815), .B(n1814), .Z(n1816) );
  ANDN U1956 ( .B(n1817), .A(n1816), .Z(n1818) );
  NAND U1957 ( .A(n1819), .B(n1818), .Z(n591) );
  NAND U1958 ( .A(n796), .B(\stack[6][7] ), .Z(n1821) );
  NAND U1959 ( .A(n795), .B(\stack[7][7] ), .Z(n1820) );
  NAND U1960 ( .A(n1821), .B(n1820), .Z(n592) );
  NAND U1961 ( .A(n796), .B(\stack[5][7] ), .Z(n1823) );
  NANDN U1962 ( .A(n2084), .B(\stack[7][7] ), .Z(n1822) );
  AND U1963 ( .A(n1823), .B(n1822), .Z(n1825) );
  NANDN U1964 ( .A(n2087), .B(\stack[6][7] ), .Z(n1824) );
  NAND U1965 ( .A(n1825), .B(n1824), .Z(n593) );
  NAND U1966 ( .A(n796), .B(\stack[4][7] ), .Z(n1827) );
  NANDN U1967 ( .A(n2084), .B(\stack[6][7] ), .Z(n1826) );
  AND U1968 ( .A(n1827), .B(n1826), .Z(n1829) );
  NANDN U1969 ( .A(n2087), .B(\stack[5][7] ), .Z(n1828) );
  NAND U1970 ( .A(n1829), .B(n1828), .Z(n594) );
  NAND U1971 ( .A(n796), .B(\stack[3][7] ), .Z(n1831) );
  NANDN U1972 ( .A(n2084), .B(\stack[5][7] ), .Z(n1830) );
  AND U1973 ( .A(n1831), .B(n1830), .Z(n1833) );
  NANDN U1974 ( .A(n2087), .B(\stack[4][7] ), .Z(n1832) );
  NAND U1975 ( .A(n1833), .B(n1832), .Z(n595) );
  NAND U1976 ( .A(n796), .B(\stack[2][7] ), .Z(n1835) );
  NANDN U1977 ( .A(n2084), .B(\stack[4][7] ), .Z(n1834) );
  AND U1978 ( .A(n1835), .B(n1834), .Z(n1837) );
  NANDN U1979 ( .A(n2087), .B(\stack[3][7] ), .Z(n1836) );
  NAND U1980 ( .A(n1837), .B(n1836), .Z(n596) );
  NAND U1981 ( .A(\stack[1][7] ), .B(n796), .Z(n1839) );
  NANDN U1982 ( .A(n2084), .B(\stack[3][7] ), .Z(n1838) );
  AND U1983 ( .A(n1839), .B(n1838), .Z(n1841) );
  NANDN U1984 ( .A(n2087), .B(\stack[2][7] ), .Z(n1840) );
  NAND U1985 ( .A(n1841), .B(n1840), .Z(n597) );
  NAND U1986 ( .A(n796), .B(o[7]), .Z(n1843) );
  NANDN U1987 ( .A(n2084), .B(\stack[2][7] ), .Z(n1842) );
  AND U1988 ( .A(n1843), .B(n1842), .Z(n1845) );
  NANDN U1989 ( .A(n2087), .B(\stack[1][7] ), .Z(n1844) );
  NAND U1990 ( .A(n1845), .B(n1844), .Z(n598) );
  NANDN U1991 ( .A(n2096), .B(\stack[1][7] ), .Z(n1846) );
  XOR U1992 ( .A(n1848), .B(n1847), .Z(n1849) );
  NAND U1993 ( .A(n1849), .B(n2092), .Z(n1850) );
  AND U1994 ( .A(n1851), .B(n1850), .Z(n1856) );
  NANDN U1995 ( .A(n1852), .B(n2093), .Z(n1854) );
  NAND U1996 ( .A(n796), .B(x[7]), .Z(n1853) );
  NAND U1997 ( .A(n1854), .B(n1853), .Z(n1855) );
  ANDN U1998 ( .B(n1856), .A(n1855), .Z(n1858) );
  NAND U1999 ( .A(n2090), .B(o[7]), .Z(n1857) );
  NAND U2000 ( .A(n1858), .B(n1857), .Z(n599) );
  NAND U2001 ( .A(n796), .B(\stack[6][6] ), .Z(n1860) );
  NAND U2002 ( .A(n795), .B(\stack[7][6] ), .Z(n1859) );
  NAND U2003 ( .A(n1860), .B(n1859), .Z(n600) );
  NAND U2004 ( .A(n796), .B(\stack[5][6] ), .Z(n1862) );
  NANDN U2005 ( .A(n2084), .B(\stack[7][6] ), .Z(n1861) );
  AND U2006 ( .A(n1862), .B(n1861), .Z(n1864) );
  NANDN U2007 ( .A(n2087), .B(\stack[6][6] ), .Z(n1863) );
  NAND U2008 ( .A(n1864), .B(n1863), .Z(n601) );
  NAND U2009 ( .A(n796), .B(\stack[4][6] ), .Z(n1866) );
  NANDN U2010 ( .A(n2084), .B(\stack[6][6] ), .Z(n1865) );
  AND U2011 ( .A(n1866), .B(n1865), .Z(n1868) );
  NANDN U2012 ( .A(n2087), .B(\stack[5][6] ), .Z(n1867) );
  NAND U2013 ( .A(n1868), .B(n1867), .Z(n602) );
  NAND U2014 ( .A(n796), .B(\stack[3][6] ), .Z(n1870) );
  NANDN U2015 ( .A(n2084), .B(\stack[5][6] ), .Z(n1869) );
  AND U2016 ( .A(n1870), .B(n1869), .Z(n1872) );
  NANDN U2017 ( .A(n2087), .B(\stack[4][6] ), .Z(n1871) );
  NAND U2018 ( .A(n1872), .B(n1871), .Z(n603) );
  NAND U2019 ( .A(n796), .B(\stack[2][6] ), .Z(n1874) );
  NANDN U2020 ( .A(n2084), .B(\stack[4][6] ), .Z(n1873) );
  AND U2021 ( .A(n1874), .B(n1873), .Z(n1876) );
  NANDN U2022 ( .A(n2087), .B(\stack[3][6] ), .Z(n1875) );
  NAND U2023 ( .A(n1876), .B(n1875), .Z(n604) );
  NAND U2024 ( .A(\stack[1][6] ), .B(n796), .Z(n1878) );
  NANDN U2025 ( .A(n2084), .B(\stack[3][6] ), .Z(n1877) );
  AND U2026 ( .A(n1878), .B(n1877), .Z(n1880) );
  NANDN U2027 ( .A(n2087), .B(\stack[2][6] ), .Z(n1879) );
  NAND U2028 ( .A(n1880), .B(n1879), .Z(n605) );
  NAND U2029 ( .A(n796), .B(o[6]), .Z(n1882) );
  NANDN U2030 ( .A(n2084), .B(\stack[2][6] ), .Z(n1881) );
  AND U2031 ( .A(n1882), .B(n1881), .Z(n1884) );
  NANDN U2032 ( .A(n2087), .B(\stack[1][6] ), .Z(n1883) );
  NAND U2033 ( .A(n1884), .B(n1883), .Z(n606) );
  NANDN U2034 ( .A(n1885), .B(n2092), .Z(n1886) );
  NAND U2035 ( .A(\stack[1][6] ), .B(n2093), .Z(n1889) );
  NAND U2036 ( .A(n2082), .B(n1887), .Z(n1888) );
  AND U2037 ( .A(n1889), .B(n1888), .Z(n1890) );
  NAND U2038 ( .A(n2083), .B(n1890), .Z(n1891) );
  NAND U2039 ( .A(o[6]), .B(n1891), .Z(n1895) );
  NAND U2040 ( .A(n796), .B(x[6]), .Z(n1893) );
  NANDN U2041 ( .A(n2096), .B(\stack[1][6] ), .Z(n1892) );
  NAND U2042 ( .A(n1893), .B(n1892), .Z(n1894) );
  ANDN U2043 ( .B(n1895), .A(n1894), .Z(n1896) );
  NAND U2044 ( .A(n1897), .B(n1896), .Z(n607) );
  NAND U2045 ( .A(n796), .B(\stack[6][5] ), .Z(n1899) );
  NAND U2046 ( .A(n795), .B(\stack[7][5] ), .Z(n1898) );
  NAND U2047 ( .A(n1899), .B(n1898), .Z(n608) );
  NAND U2048 ( .A(n796), .B(\stack[5][5] ), .Z(n1901) );
  NANDN U2049 ( .A(n2084), .B(\stack[7][5] ), .Z(n1900) );
  AND U2050 ( .A(n1901), .B(n1900), .Z(n1903) );
  NANDN U2051 ( .A(n2087), .B(\stack[6][5] ), .Z(n1902) );
  NAND U2052 ( .A(n1903), .B(n1902), .Z(n609) );
  NAND U2053 ( .A(n796), .B(\stack[4][5] ), .Z(n1905) );
  NANDN U2054 ( .A(n2084), .B(\stack[6][5] ), .Z(n1904) );
  AND U2055 ( .A(n1905), .B(n1904), .Z(n1907) );
  NANDN U2056 ( .A(n2087), .B(\stack[5][5] ), .Z(n1906) );
  NAND U2057 ( .A(n1907), .B(n1906), .Z(n610) );
  NAND U2058 ( .A(n796), .B(\stack[3][5] ), .Z(n1909) );
  NANDN U2059 ( .A(n2084), .B(\stack[5][5] ), .Z(n1908) );
  AND U2060 ( .A(n1909), .B(n1908), .Z(n1911) );
  NANDN U2061 ( .A(n2087), .B(\stack[4][5] ), .Z(n1910) );
  NAND U2062 ( .A(n1911), .B(n1910), .Z(n611) );
  NAND U2063 ( .A(n796), .B(\stack[2][5] ), .Z(n1913) );
  NANDN U2064 ( .A(n2084), .B(\stack[4][5] ), .Z(n1912) );
  AND U2065 ( .A(n1913), .B(n1912), .Z(n1915) );
  NANDN U2066 ( .A(n2087), .B(\stack[3][5] ), .Z(n1914) );
  NAND U2067 ( .A(n1915), .B(n1914), .Z(n612) );
  NAND U2068 ( .A(\stack[1][5] ), .B(n796), .Z(n1917) );
  NANDN U2069 ( .A(n2084), .B(\stack[3][5] ), .Z(n1916) );
  AND U2070 ( .A(n1917), .B(n1916), .Z(n1919) );
  NANDN U2071 ( .A(n2087), .B(\stack[2][5] ), .Z(n1918) );
  NAND U2072 ( .A(n1919), .B(n1918), .Z(n613) );
  NAND U2073 ( .A(o[5]), .B(n796), .Z(n1921) );
  NANDN U2074 ( .A(n2084), .B(\stack[2][5] ), .Z(n1920) );
  AND U2075 ( .A(n1921), .B(n1920), .Z(n1923) );
  NANDN U2076 ( .A(n2087), .B(\stack[1][5] ), .Z(n1922) );
  NAND U2077 ( .A(n1923), .B(n1922), .Z(n614) );
  NANDN U2078 ( .A(n2096), .B(\stack[1][5] ), .Z(n1924) );
  XOR U2079 ( .A(n1926), .B(n1925), .Z(n1927) );
  NAND U2080 ( .A(n1927), .B(n2092), .Z(n1928) );
  AND U2081 ( .A(n1929), .B(n1928), .Z(n1934) );
  NANDN U2082 ( .A(n1930), .B(n2093), .Z(n1932) );
  NAND U2083 ( .A(n796), .B(x[5]), .Z(n1931) );
  NAND U2084 ( .A(n1932), .B(n1931), .Z(n1933) );
  ANDN U2085 ( .B(n1934), .A(n1933), .Z(n1936) );
  NAND U2086 ( .A(o[5]), .B(n2090), .Z(n1935) );
  NAND U2087 ( .A(n1936), .B(n1935), .Z(n615) );
  NAND U2088 ( .A(n796), .B(\stack[6][4] ), .Z(n1938) );
  NAND U2089 ( .A(n795), .B(\stack[7][4] ), .Z(n1937) );
  NAND U2090 ( .A(n1938), .B(n1937), .Z(n616) );
  NAND U2091 ( .A(n796), .B(\stack[5][4] ), .Z(n1940) );
  NANDN U2092 ( .A(n2084), .B(\stack[7][4] ), .Z(n1939) );
  AND U2093 ( .A(n1940), .B(n1939), .Z(n1942) );
  NANDN U2094 ( .A(n2087), .B(\stack[6][4] ), .Z(n1941) );
  NAND U2095 ( .A(n1942), .B(n1941), .Z(n617) );
  NAND U2096 ( .A(n796), .B(\stack[4][4] ), .Z(n1944) );
  NANDN U2097 ( .A(n2084), .B(\stack[6][4] ), .Z(n1943) );
  AND U2098 ( .A(n1944), .B(n1943), .Z(n1946) );
  NANDN U2099 ( .A(n2087), .B(\stack[5][4] ), .Z(n1945) );
  NAND U2100 ( .A(n1946), .B(n1945), .Z(n618) );
  NAND U2101 ( .A(n796), .B(\stack[3][4] ), .Z(n1948) );
  NANDN U2102 ( .A(n2084), .B(\stack[5][4] ), .Z(n1947) );
  AND U2103 ( .A(n1948), .B(n1947), .Z(n1950) );
  NANDN U2104 ( .A(n2087), .B(\stack[4][4] ), .Z(n1949) );
  NAND U2105 ( .A(n1950), .B(n1949), .Z(n619) );
  NAND U2106 ( .A(n796), .B(\stack[2][4] ), .Z(n1952) );
  NANDN U2107 ( .A(n2084), .B(\stack[4][4] ), .Z(n1951) );
  AND U2108 ( .A(n1952), .B(n1951), .Z(n1954) );
  NANDN U2109 ( .A(n2087), .B(\stack[3][4] ), .Z(n1953) );
  NAND U2110 ( .A(n1954), .B(n1953), .Z(n620) );
  NAND U2111 ( .A(\stack[1][4] ), .B(n796), .Z(n1956) );
  NANDN U2112 ( .A(n2084), .B(\stack[3][4] ), .Z(n1955) );
  AND U2113 ( .A(n1956), .B(n1955), .Z(n1958) );
  NANDN U2114 ( .A(n2087), .B(\stack[2][4] ), .Z(n1957) );
  NAND U2115 ( .A(n1958), .B(n1957), .Z(n621) );
  NAND U2116 ( .A(n796), .B(o[4]), .Z(n1960) );
  NANDN U2117 ( .A(n2084), .B(\stack[2][4] ), .Z(n1959) );
  AND U2118 ( .A(n1960), .B(n1959), .Z(n1962) );
  NANDN U2119 ( .A(n2087), .B(\stack[1][4] ), .Z(n1961) );
  NAND U2120 ( .A(n1962), .B(n1961), .Z(n622) );
  NANDN U2121 ( .A(n1963), .B(n2092), .Z(n1964) );
  NAND U2122 ( .A(\stack[1][4] ), .B(n2093), .Z(n1967) );
  NAND U2123 ( .A(n2082), .B(n1965), .Z(n1966) );
  AND U2124 ( .A(n1967), .B(n1966), .Z(n1968) );
  NAND U2125 ( .A(n2083), .B(n1968), .Z(n1969) );
  NAND U2126 ( .A(n1969), .B(o[4]), .Z(n1973) );
  NAND U2127 ( .A(n796), .B(x[4]), .Z(n1971) );
  NANDN U2128 ( .A(n2096), .B(\stack[1][4] ), .Z(n1970) );
  NAND U2129 ( .A(n1971), .B(n1970), .Z(n1972) );
  ANDN U2130 ( .B(n1973), .A(n1972), .Z(n1974) );
  NAND U2131 ( .A(n1975), .B(n1974), .Z(n623) );
  NAND U2132 ( .A(n796), .B(\stack[6][3] ), .Z(n1977) );
  NAND U2133 ( .A(n795), .B(\stack[7][3] ), .Z(n1976) );
  NAND U2134 ( .A(n1977), .B(n1976), .Z(n624) );
  NAND U2135 ( .A(n796), .B(\stack[5][3] ), .Z(n1979) );
  NANDN U2136 ( .A(n2084), .B(\stack[7][3] ), .Z(n1978) );
  AND U2137 ( .A(n1979), .B(n1978), .Z(n1981) );
  NANDN U2138 ( .A(n2087), .B(\stack[6][3] ), .Z(n1980) );
  NAND U2139 ( .A(n1981), .B(n1980), .Z(n625) );
  NAND U2140 ( .A(n796), .B(\stack[4][3] ), .Z(n1983) );
  NANDN U2141 ( .A(n2084), .B(\stack[6][3] ), .Z(n1982) );
  AND U2142 ( .A(n1983), .B(n1982), .Z(n1985) );
  NANDN U2143 ( .A(n2087), .B(\stack[5][3] ), .Z(n1984) );
  NAND U2144 ( .A(n1985), .B(n1984), .Z(n626) );
  NAND U2145 ( .A(n796), .B(\stack[3][3] ), .Z(n1987) );
  NANDN U2146 ( .A(n2084), .B(\stack[5][3] ), .Z(n1986) );
  AND U2147 ( .A(n1987), .B(n1986), .Z(n1989) );
  NANDN U2148 ( .A(n2087), .B(\stack[4][3] ), .Z(n1988) );
  NAND U2149 ( .A(n1989), .B(n1988), .Z(n627) );
  NAND U2150 ( .A(n796), .B(\stack[2][3] ), .Z(n1991) );
  NANDN U2151 ( .A(n2084), .B(\stack[4][3] ), .Z(n1990) );
  AND U2152 ( .A(n1991), .B(n1990), .Z(n1993) );
  NANDN U2153 ( .A(n2087), .B(\stack[3][3] ), .Z(n1992) );
  NAND U2154 ( .A(n1993), .B(n1992), .Z(n628) );
  NAND U2155 ( .A(\stack[1][3] ), .B(n796), .Z(n1995) );
  NANDN U2156 ( .A(n2084), .B(\stack[3][3] ), .Z(n1994) );
  AND U2157 ( .A(n1995), .B(n1994), .Z(n1997) );
  NANDN U2158 ( .A(n2087), .B(\stack[2][3] ), .Z(n1996) );
  NAND U2159 ( .A(n1997), .B(n1996), .Z(n629) );
  NAND U2160 ( .A(n796), .B(o[3]), .Z(n1999) );
  NANDN U2161 ( .A(n2084), .B(\stack[2][3] ), .Z(n1998) );
  AND U2162 ( .A(n1999), .B(n1998), .Z(n2001) );
  NANDN U2163 ( .A(n2087), .B(\stack[1][3] ), .Z(n2000) );
  NAND U2164 ( .A(n2001), .B(n2000), .Z(n630) );
  NAND U2165 ( .A(n796), .B(x[3]), .Z(n2004) );
  NAND U2166 ( .A(n2002), .B(n2093), .Z(n2003) );
  NAND U2167 ( .A(n2004), .B(n2003), .Z(n2012) );
  XOR U2168 ( .A(n2006), .B(n2005), .Z(n2007) );
  NAND U2169 ( .A(n2007), .B(n2092), .Z(n2010) );
  NANDN U2170 ( .A(n2096), .B(\stack[1][3] ), .Z(n2008) );
  NAND U2171 ( .A(n2010), .B(n2009), .Z(n2011) );
  NOR U2172 ( .A(n2012), .B(n2011), .Z(n2014) );
  NAND U2173 ( .A(n2090), .B(o[3]), .Z(n2013) );
  NAND U2174 ( .A(n2014), .B(n2013), .Z(n631) );
  NAND U2175 ( .A(n796), .B(\stack[6][2] ), .Z(n2016) );
  NAND U2176 ( .A(n795), .B(\stack[7][2] ), .Z(n2015) );
  NAND U2177 ( .A(n2016), .B(n2015), .Z(n632) );
  NAND U2178 ( .A(n796), .B(\stack[5][2] ), .Z(n2018) );
  NANDN U2179 ( .A(n2084), .B(\stack[7][2] ), .Z(n2017) );
  AND U2180 ( .A(n2018), .B(n2017), .Z(n2020) );
  NANDN U2181 ( .A(n2087), .B(\stack[6][2] ), .Z(n2019) );
  NAND U2182 ( .A(n2020), .B(n2019), .Z(n633) );
  NAND U2183 ( .A(n796), .B(\stack[4][2] ), .Z(n2022) );
  NANDN U2184 ( .A(n2084), .B(\stack[6][2] ), .Z(n2021) );
  AND U2185 ( .A(n2022), .B(n2021), .Z(n2024) );
  NANDN U2186 ( .A(n2087), .B(\stack[5][2] ), .Z(n2023) );
  NAND U2187 ( .A(n2024), .B(n2023), .Z(n634) );
  NAND U2188 ( .A(n796), .B(\stack[3][2] ), .Z(n2026) );
  NANDN U2189 ( .A(n2084), .B(\stack[5][2] ), .Z(n2025) );
  AND U2190 ( .A(n2026), .B(n2025), .Z(n2028) );
  NANDN U2191 ( .A(n2087), .B(\stack[4][2] ), .Z(n2027) );
  NAND U2192 ( .A(n2028), .B(n2027), .Z(n635) );
  NAND U2193 ( .A(n796), .B(\stack[2][2] ), .Z(n2030) );
  NANDN U2194 ( .A(n2084), .B(\stack[4][2] ), .Z(n2029) );
  AND U2195 ( .A(n2030), .B(n2029), .Z(n2032) );
  NANDN U2196 ( .A(n2087), .B(\stack[3][2] ), .Z(n2031) );
  NAND U2197 ( .A(n2032), .B(n2031), .Z(n636) );
  NAND U2198 ( .A(\stack[1][2] ), .B(n796), .Z(n2034) );
  NANDN U2199 ( .A(n2084), .B(\stack[3][2] ), .Z(n2033) );
  AND U2200 ( .A(n2034), .B(n2033), .Z(n2036) );
  NANDN U2201 ( .A(n2087), .B(\stack[2][2] ), .Z(n2035) );
  NAND U2202 ( .A(n2036), .B(n2035), .Z(n637) );
  NAND U2203 ( .A(n796), .B(o[2]), .Z(n2038) );
  NANDN U2204 ( .A(n2084), .B(\stack[2][2] ), .Z(n2037) );
  AND U2205 ( .A(n2038), .B(n2037), .Z(n2040) );
  NANDN U2206 ( .A(n2087), .B(\stack[1][2] ), .Z(n2039) );
  NAND U2207 ( .A(n2040), .B(n2039), .Z(n638) );
  NANDN U2208 ( .A(n2096), .B(\stack[1][2] ), .Z(n2041) );
  XNOR U2209 ( .A(n2043), .B(n2042), .Z(n2044) );
  NAND U2210 ( .A(n2044), .B(n2092), .Z(n2045) );
  AND U2211 ( .A(n2046), .B(n2045), .Z(n2051) );
  NANDN U2212 ( .A(n2047), .B(n2093), .Z(n2049) );
  NAND U2213 ( .A(n796), .B(x[2]), .Z(n2048) );
  NAND U2214 ( .A(n2049), .B(n2048), .Z(n2050) );
  ANDN U2215 ( .B(n2051), .A(n2050), .Z(n2053) );
  NAND U2216 ( .A(n2090), .B(o[2]), .Z(n2052) );
  NAND U2217 ( .A(n2053), .B(n2052), .Z(n639) );
  NAND U2218 ( .A(n796), .B(\stack[6][1] ), .Z(n2055) );
  NAND U2219 ( .A(n795), .B(\stack[7][1] ), .Z(n2054) );
  NAND U2220 ( .A(n2055), .B(n2054), .Z(n640) );
  NAND U2221 ( .A(n796), .B(\stack[5][1] ), .Z(n2057) );
  NANDN U2222 ( .A(n2084), .B(\stack[7][1] ), .Z(n2056) );
  AND U2223 ( .A(n2057), .B(n2056), .Z(n2059) );
  NANDN U2224 ( .A(n2087), .B(\stack[6][1] ), .Z(n2058) );
  NAND U2225 ( .A(n2059), .B(n2058), .Z(n641) );
  NAND U2226 ( .A(n796), .B(\stack[4][1] ), .Z(n2061) );
  NANDN U2227 ( .A(n2084), .B(\stack[6][1] ), .Z(n2060) );
  AND U2228 ( .A(n2061), .B(n2060), .Z(n2063) );
  NANDN U2229 ( .A(n2087), .B(\stack[5][1] ), .Z(n2062) );
  NAND U2230 ( .A(n2063), .B(n2062), .Z(n642) );
  NAND U2231 ( .A(n796), .B(\stack[3][1] ), .Z(n2065) );
  NANDN U2232 ( .A(n2084), .B(\stack[5][1] ), .Z(n2064) );
  AND U2233 ( .A(n2065), .B(n2064), .Z(n2067) );
  NANDN U2234 ( .A(n2087), .B(\stack[4][1] ), .Z(n2066) );
  NAND U2235 ( .A(n2067), .B(n2066), .Z(n643) );
  NAND U2236 ( .A(n796), .B(\stack[2][1] ), .Z(n2069) );
  NANDN U2237 ( .A(n2084), .B(\stack[4][1] ), .Z(n2068) );
  AND U2238 ( .A(n2069), .B(n2068), .Z(n2071) );
  NANDN U2239 ( .A(n2087), .B(\stack[3][1] ), .Z(n2070) );
  NAND U2240 ( .A(n2071), .B(n2070), .Z(n644) );
  NAND U2241 ( .A(\stack[1][1] ), .B(n796), .Z(n2073) );
  NANDN U2242 ( .A(n2084), .B(\stack[3][1] ), .Z(n2072) );
  AND U2243 ( .A(n2073), .B(n2072), .Z(n2075) );
  NANDN U2244 ( .A(n2087), .B(\stack[2][1] ), .Z(n2074) );
  NAND U2245 ( .A(n2075), .B(n2074), .Z(n645) );
  NAND U2246 ( .A(n796), .B(o[1]), .Z(n2077) );
  NANDN U2247 ( .A(n2084), .B(\stack[2][1] ), .Z(n2076) );
  AND U2248 ( .A(n2077), .B(n2076), .Z(n2079) );
  NANDN U2249 ( .A(n2087), .B(\stack[1][1] ), .Z(n2078) );
  NAND U2250 ( .A(n2079), .B(n2078), .Z(n646) );
  NAND U2251 ( .A(o[0]), .B(n796), .Z(n2086) );
  NANDN U2252 ( .A(n2084), .B(\stack[2][0] ), .Z(n2085) );
  AND U2253 ( .A(n2086), .B(n2085), .Z(n2089) );
  NANDN U2254 ( .A(n2087), .B(\stack[1][0] ), .Z(n2088) );
  NAND U2255 ( .A(n2089), .B(n2088), .Z(n648) );
  NAND U2256 ( .A(o[0]), .B(n2090), .Z(n2091) );
  NAND U2257 ( .A(n796), .B(x[0]), .Z(n2099) );
  OR U2258 ( .A(n2093), .B(n2092), .Z(n2094) );
  NAND U2259 ( .A(o[0]), .B(n2094), .Z(n2095) );
  AND U2260 ( .A(n2096), .B(n2095), .Z(n2097) );
  NANDN U2261 ( .A(n2097), .B(\stack[1][0] ), .Z(n2098) );
  AND U2262 ( .A(n2099), .B(n2098), .Z(n2100) );
  NAND U2263 ( .A(n2101), .B(n2100), .Z(n649) );
endmodule

