
module hamming_N160_CC4 ( clk, rst, x, y, o );
  input [39:0] x;
  input [39:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244;
  wire   [7:0] oglobal;

  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NANDN U43 ( .A(n135), .B(n134), .Z(n1) );
  NANDN U44 ( .A(n137), .B(n136), .Z(n2) );
  AND U45 ( .A(n1), .B(n2), .Z(n178) );
  NANDN U46 ( .A(n75), .B(n74), .Z(n3) );
  NANDN U47 ( .A(n73), .B(n72), .Z(n4) );
  NAND U48 ( .A(n3), .B(n4), .Z(n176) );
  NANDN U49 ( .A(n148), .B(n147), .Z(n5) );
  NANDN U50 ( .A(n150), .B(n149), .Z(n6) );
  AND U51 ( .A(n5), .B(n6), .Z(n168) );
  NAND U52 ( .A(n174), .B(n172), .Z(n7) );
  XOR U53 ( .A(n172), .B(n174), .Z(n8) );
  NANDN U54 ( .A(n173), .B(n8), .Z(n9) );
  NAND U55 ( .A(n7), .B(n9), .Z(n209) );
  NANDN U56 ( .A(n133), .B(n132), .Z(n10) );
  NANDN U57 ( .A(n131), .B(n130), .Z(n11) );
  NAND U58 ( .A(n10), .B(n11), .Z(n177) );
  XOR U59 ( .A(oglobal[1]), .B(n175), .Z(n12) );
  NAND U60 ( .A(n12), .B(n176), .Z(n13) );
  NAND U61 ( .A(oglobal[1]), .B(n175), .Z(n14) );
  AND U62 ( .A(n13), .B(n14), .Z(n215) );
  NAND U63 ( .A(n170), .B(n169), .Z(n15) );
  XOR U64 ( .A(n169), .B(n170), .Z(n16) );
  NAND U65 ( .A(n16), .B(n168), .Z(n17) );
  NAND U66 ( .A(n15), .B(n17), .Z(n219) );
  NAND U67 ( .A(n61), .B(n60), .Z(n18) );
  NANDN U68 ( .A(n59), .B(n58), .Z(n19) );
  AND U69 ( .A(n18), .B(n19), .Z(n173) );
  XOR U70 ( .A(oglobal[2]), .B(n216), .Z(n20) );
  NANDN U71 ( .A(n215), .B(n20), .Z(n21) );
  NAND U72 ( .A(oglobal[2]), .B(n216), .Z(n22) );
  AND U73 ( .A(n21), .B(n22), .Z(n221) );
  XOR U74 ( .A(n70), .B(n69), .Z(n23) );
  NANDN U75 ( .A(n68), .B(n23), .Z(n24) );
  NAND U76 ( .A(n70), .B(n69), .Z(n25) );
  AND U77 ( .A(n24), .B(n25), .Z(n172) );
  NAND U78 ( .A(n186), .B(n184), .Z(n26) );
  XOR U79 ( .A(n184), .B(n186), .Z(n27) );
  NANDN U80 ( .A(n185), .B(n27), .Z(n28) );
  NAND U81 ( .A(n26), .B(n28), .Z(n202) );
  NAND U82 ( .A(n218), .B(n217), .Z(n29) );
  XOR U83 ( .A(n217), .B(n218), .Z(n30) );
  NANDN U84 ( .A(n219), .B(n30), .Z(n31) );
  NAND U85 ( .A(n29), .B(n31), .Z(n222) );
  NANDN U86 ( .A(n129), .B(n128), .Z(n32) );
  NANDN U87 ( .A(n127), .B(n126), .Z(n33) );
  NAND U88 ( .A(n32), .B(n33), .Z(n180) );
  NANDN U89 ( .A(n79), .B(n78), .Z(n34) );
  NANDN U90 ( .A(n77), .B(n76), .Z(n35) );
  NAND U91 ( .A(n34), .B(n35), .Z(n175) );
  NANDN U92 ( .A(n113), .B(n112), .Z(n36) );
  NANDN U93 ( .A(n111), .B(n110), .Z(n37) );
  NAND U94 ( .A(n36), .B(n37), .Z(n163) );
  NANDN U95 ( .A(n139), .B(n138), .Z(n38) );
  NANDN U96 ( .A(n141), .B(n140), .Z(n39) );
  AND U97 ( .A(n38), .B(n39), .Z(n170) );
  NANDN U98 ( .A(n96), .B(n95), .Z(n40) );
  NANDN U99 ( .A(n94), .B(n93), .Z(n41) );
  NAND U100 ( .A(n40), .B(n41), .Z(n156) );
  XOR U101 ( .A(n155), .B(n154), .Z(n42) );
  NANDN U102 ( .A(n153), .B(n42), .Z(n43) );
  NAND U103 ( .A(n155), .B(n154), .Z(n44) );
  AND U104 ( .A(n43), .B(n44), .Z(n203) );
  NAND U105 ( .A(n202), .B(n200), .Z(n45) );
  XOR U106 ( .A(n200), .B(n202), .Z(n46) );
  NANDN U107 ( .A(n201), .B(n46), .Z(n47) );
  NAND U108 ( .A(n45), .B(n47), .Z(n225) );
  NAND U109 ( .A(n224), .B(n223), .Z(n48) );
  XOR U110 ( .A(n223), .B(n224), .Z(n49) );
  NAND U111 ( .A(n49), .B(n222), .Z(n50) );
  NAND U112 ( .A(n48), .B(n50), .Z(n232) );
  XNOR U113 ( .A(x[35]), .B(y[35]), .Z(n94) );
  XOR U114 ( .A(x[33]), .B(y[33]), .Z(n93) );
  XNOR U115 ( .A(n94), .B(n93), .Z(n95) );
  XNOR U116 ( .A(x[27]), .B(y[27]), .Z(n75) );
  XNOR U117 ( .A(x[39]), .B(y[39]), .Z(n73) );
  XOR U118 ( .A(x[25]), .B(y[25]), .Z(n72) );
  XNOR U119 ( .A(n73), .B(n72), .Z(n74) );
  XOR U120 ( .A(n75), .B(n74), .Z(n96) );
  XNOR U121 ( .A(n95), .B(n96), .Z(n62) );
  XNOR U122 ( .A(x[5]), .B(y[5]), .Z(n123) );
  XNOR U123 ( .A(x[3]), .B(y[3]), .Z(n121) );
  XNOR U124 ( .A(x[1]), .B(y[1]), .Z(n120) );
  XOR U125 ( .A(n121), .B(n120), .Z(n122) );
  XOR U126 ( .A(n123), .B(n122), .Z(n63) );
  XNOR U127 ( .A(n62), .B(n63), .Z(n64) );
  XNOR U128 ( .A(x[17]), .B(y[17]), .Z(n90) );
  XNOR U129 ( .A(x[15]), .B(y[15]), .Z(n88) );
  XNOR U130 ( .A(x[13]), .B(y[13]), .Z(n87) );
  XOR U131 ( .A(n88), .B(n87), .Z(n89) );
  XOR U132 ( .A(n90), .B(n89), .Z(n65) );
  XNOR U133 ( .A(n64), .B(n65), .Z(n52) );
  XNOR U134 ( .A(x[18]), .B(y[18]), .Z(n150) );
  XNOR U135 ( .A(x[22]), .B(y[22]), .Z(n148) );
  XOR U136 ( .A(x[20]), .B(y[20]), .Z(n147) );
  XNOR U137 ( .A(n148), .B(n147), .Z(n149) );
  XOR U138 ( .A(n150), .B(n149), .Z(n84) );
  XNOR U139 ( .A(x[24]), .B(y[24]), .Z(n141) );
  XNOR U140 ( .A(x[28]), .B(y[28]), .Z(n139) );
  XOR U141 ( .A(x[26]), .B(y[26]), .Z(n138) );
  XNOR U142 ( .A(n139), .B(n138), .Z(n140) );
  XOR U143 ( .A(n141), .B(n140), .Z(n81) );
  XNOR U144 ( .A(x[30]), .B(y[30]), .Z(n144) );
  XOR U145 ( .A(x[32]), .B(y[32]), .Z(n142) );
  XNOR U146 ( .A(oglobal[0]), .B(n142), .Z(n143) );
  XOR U147 ( .A(n144), .B(n143), .Z(n82) );
  XNOR U148 ( .A(n81), .B(n82), .Z(n83) );
  XNOR U149 ( .A(n84), .B(n83), .Z(n53) );
  XOR U150 ( .A(n52), .B(n53), .Z(n54) );
  XNOR U151 ( .A(x[6]), .B(y[6]), .Z(n137) );
  XNOR U152 ( .A(x[10]), .B(y[10]), .Z(n135) );
  XOR U153 ( .A(x[8]), .B(y[8]), .Z(n134) );
  XNOR U154 ( .A(n135), .B(n134), .Z(n136) );
  XOR U155 ( .A(n137), .B(n136), .Z(n70) );
  XNOR U156 ( .A(x[0]), .B(y[0]), .Z(n113) );
  XNOR U157 ( .A(x[4]), .B(y[4]), .Z(n111) );
  XOR U158 ( .A(x[2]), .B(y[2]), .Z(n110) );
  XNOR U159 ( .A(n111), .B(n110), .Z(n112) );
  XNOR U160 ( .A(n113), .B(n112), .Z(n68) );
  XNOR U161 ( .A(x[12]), .B(y[12]), .Z(n133) );
  XNOR U162 ( .A(x[16]), .B(y[16]), .Z(n131) );
  XOR U163 ( .A(x[14]), .B(y[14]), .Z(n130) );
  XNOR U164 ( .A(n131), .B(n130), .Z(n132) );
  XOR U165 ( .A(n133), .B(n132), .Z(n69) );
  XOR U166 ( .A(n68), .B(n69), .Z(n51) );
  XNOR U167 ( .A(n70), .B(n51), .Z(n107) );
  XNOR U168 ( .A(x[31]), .B(y[31]), .Z(n100) );
  XNOR U169 ( .A(x[37]), .B(y[37]), .Z(n98) );
  XNOR U170 ( .A(x[29]), .B(y[29]), .Z(n97) );
  XOR U171 ( .A(n98), .B(n97), .Z(n99) );
  XNOR U172 ( .A(n100), .B(n99), .Z(n60) );
  XNOR U173 ( .A(x[11]), .B(y[11]), .Z(n117) );
  XNOR U174 ( .A(x[9]), .B(y[9]), .Z(n115) );
  XNOR U175 ( .A(x[7]), .B(y[7]), .Z(n114) );
  XOR U176 ( .A(n115), .B(n114), .Z(n116) );
  XNOR U177 ( .A(n117), .B(n116), .Z(n58) );
  XNOR U178 ( .A(x[23]), .B(y[23]), .Z(n79) );
  XNOR U179 ( .A(x[21]), .B(y[21]), .Z(n77) );
  XOR U180 ( .A(x[19]), .B(y[19]), .Z(n76) );
  XNOR U181 ( .A(n77), .B(n76), .Z(n78) );
  XOR U182 ( .A(n79), .B(n78), .Z(n59) );
  XNOR U183 ( .A(n58), .B(n59), .Z(n61) );
  XOR U184 ( .A(n60), .B(n61), .Z(n104) );
  XNOR U185 ( .A(x[34]), .B(y[34]), .Z(n129) );
  XNOR U186 ( .A(x[38]), .B(y[38]), .Z(n127) );
  XOR U187 ( .A(x[36]), .B(y[36]), .Z(n126) );
  XNOR U188 ( .A(n127), .B(n126), .Z(n128) );
  XNOR U189 ( .A(n129), .B(n128), .Z(n105) );
  XOR U190 ( .A(n104), .B(n105), .Z(n106) );
  XOR U191 ( .A(n107), .B(n106), .Z(n55) );
  XNOR U192 ( .A(n54), .B(n55), .Z(o[0]) );
  NAND U193 ( .A(n53), .B(n52), .Z(n57) );
  NANDN U194 ( .A(n55), .B(n54), .Z(n56) );
  AND U195 ( .A(n57), .B(n56), .Z(n154) );
  NANDN U196 ( .A(n63), .B(n62), .Z(n67) );
  NANDN U197 ( .A(n65), .B(n64), .Z(n66) );
  NAND U198 ( .A(n67), .B(n66), .Z(n174) );
  XNOR U199 ( .A(n174), .B(n172), .Z(n71) );
  XNOR U200 ( .A(n173), .B(n71), .Z(n155) );
  XOR U201 ( .A(n175), .B(oglobal[1]), .Z(n80) );
  XOR U202 ( .A(n176), .B(n80), .Z(n186) );
  NANDN U203 ( .A(n82), .B(n81), .Z(n86) );
  NAND U204 ( .A(n84), .B(n83), .Z(n85) );
  NAND U205 ( .A(n86), .B(n85), .Z(n185) );
  OR U206 ( .A(n88), .B(n87), .Z(n92) );
  NANDN U207 ( .A(n90), .B(n89), .Z(n91) );
  NAND U208 ( .A(n92), .B(n91), .Z(n159) );
  OR U209 ( .A(n98), .B(n97), .Z(n102) );
  NANDN U210 ( .A(n100), .B(n99), .Z(n101) );
  AND U211 ( .A(n102), .B(n101), .Z(n157) );
  XNOR U212 ( .A(n156), .B(n157), .Z(n158) );
  XOR U213 ( .A(n159), .B(n158), .Z(n184) );
  XOR U214 ( .A(n185), .B(n184), .Z(n103) );
  XOR U215 ( .A(n186), .B(n103), .Z(n190) );
  OR U216 ( .A(n105), .B(n104), .Z(n109) );
  NAND U217 ( .A(n107), .B(n106), .Z(n108) );
  NAND U218 ( .A(n109), .B(n108), .Z(n187) );
  OR U219 ( .A(n115), .B(n114), .Z(n119) );
  NANDN U220 ( .A(n117), .B(n116), .Z(n118) );
  AND U221 ( .A(n119), .B(n118), .Z(n162) );
  XNOR U222 ( .A(n163), .B(n162), .Z(n164) );
  OR U223 ( .A(n121), .B(n120), .Z(n125) );
  NANDN U224 ( .A(n123), .B(n122), .Z(n124) );
  NAND U225 ( .A(n125), .B(n124), .Z(n165) );
  XNOR U226 ( .A(n164), .B(n165), .Z(n193) );
  XNOR U227 ( .A(n177), .B(n178), .Z(n179) );
  XNOR U228 ( .A(n180), .B(n179), .Z(n194) );
  XNOR U229 ( .A(n193), .B(n194), .Z(n196) );
  NAND U230 ( .A(n142), .B(oglobal[0]), .Z(n146) );
  OR U231 ( .A(n144), .B(n143), .Z(n145) );
  AND U232 ( .A(n146), .B(n145), .Z(n169) );
  XNOR U233 ( .A(n169), .B(n168), .Z(n151) );
  XOR U234 ( .A(n170), .B(n151), .Z(n195) );
  XNOR U235 ( .A(n196), .B(n195), .Z(n188) );
  XNOR U236 ( .A(n187), .B(n188), .Z(n189) );
  XNOR U237 ( .A(n190), .B(n189), .Z(n153) );
  XNOR U238 ( .A(n155), .B(n153), .Z(n152) );
  XNOR U239 ( .A(n154), .B(n152), .Z(o[1]) );
  NANDN U240 ( .A(n157), .B(n156), .Z(n161) );
  NAND U241 ( .A(n159), .B(n158), .Z(n160) );
  NAND U242 ( .A(n161), .B(n160), .Z(n217) );
  NANDN U243 ( .A(n163), .B(n162), .Z(n167) );
  NANDN U244 ( .A(n165), .B(n164), .Z(n166) );
  AND U245 ( .A(n167), .B(n166), .Z(n218) );
  XOR U246 ( .A(n218), .B(n219), .Z(n171) );
  XNOR U247 ( .A(n217), .B(n171), .Z(n211) );
  NANDN U248 ( .A(n178), .B(n177), .Z(n182) );
  NAND U249 ( .A(n180), .B(n179), .Z(n181) );
  NAND U250 ( .A(n182), .B(n181), .Z(n216) );
  XOR U251 ( .A(n215), .B(n216), .Z(n183) );
  XOR U252 ( .A(oglobal[2]), .B(n183), .Z(n210) );
  XOR U253 ( .A(n209), .B(n210), .Z(n212) );
  XNOR U254 ( .A(n211), .B(n212), .Z(n204) );
  XOR U255 ( .A(n203), .B(n204), .Z(n205) );
  NANDN U256 ( .A(n188), .B(n187), .Z(n192) );
  NAND U257 ( .A(n190), .B(n189), .Z(n191) );
  AND U258 ( .A(n192), .B(n191), .Z(n200) );
  OR U259 ( .A(n194), .B(n193), .Z(n198) );
  NANDN U260 ( .A(n196), .B(n195), .Z(n197) );
  AND U261 ( .A(n198), .B(n197), .Z(n201) );
  XNOR U262 ( .A(n200), .B(n201), .Z(n199) );
  XOR U263 ( .A(n202), .B(n199), .Z(n206) );
  XOR U264 ( .A(n205), .B(n206), .Z(o[2]) );
  NAND U265 ( .A(n204), .B(n203), .Z(n208) );
  NAND U266 ( .A(n206), .B(n205), .Z(n207) );
  AND U267 ( .A(n208), .B(n207), .Z(n226) );
  XNOR U268 ( .A(n225), .B(n226), .Z(n227) );
  NANDN U269 ( .A(n210), .B(n209), .Z(n214) );
  NANDN U270 ( .A(n212), .B(n211), .Z(n213) );
  NAND U271 ( .A(n214), .B(n213), .Z(n224) );
  XNOR U272 ( .A(oglobal[3]), .B(n221), .Z(n223) );
  XOR U273 ( .A(n223), .B(n222), .Z(n220) );
  XOR U274 ( .A(n224), .B(n220), .Z(n228) );
  XOR U275 ( .A(n227), .B(n228), .Z(o[3]) );
  NANDN U276 ( .A(n221), .B(oglobal[3]), .Z(n231) );
  XOR U277 ( .A(oglobal[4]), .B(n231), .Z(n233) );
  XOR U278 ( .A(n233), .B(n232), .Z(n235) );
  NANDN U279 ( .A(n226), .B(n225), .Z(n230) );
  NAND U280 ( .A(n228), .B(n227), .Z(n229) );
  AND U281 ( .A(n230), .B(n229), .Z(n234) );
  XOR U282 ( .A(n235), .B(n234), .Z(o[4]) );
  NANDN U283 ( .A(n231), .B(oglobal[4]), .Z(n238) );
  XOR U284 ( .A(oglobal[5]), .B(n238), .Z(n240) );
  NANDN U285 ( .A(n233), .B(n232), .Z(n237) );
  OR U286 ( .A(n235), .B(n234), .Z(n236) );
  AND U287 ( .A(n237), .B(n236), .Z(n239) );
  XOR U288 ( .A(n240), .B(n239), .Z(o[5]) );
  NANDN U289 ( .A(n238), .B(oglobal[5]), .Z(n242) );
  OR U290 ( .A(n240), .B(n239), .Z(n241) );
  NAND U291 ( .A(n242), .B(n241), .Z(n243) );
  XOR U292 ( .A(n243), .B(oglobal[6]), .Z(o[6]) );
  NAND U293 ( .A(oglobal[6]), .B(n243), .Z(n244) );
  XNOR U294 ( .A(oglobal[7]), .B(n244), .Z(o[7]) );
endmodule

