
module mult_N256_CC8 ( clk, rst, a, b, c );
  input [255:0] a;
  input [31:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
         n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
         n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553,
         n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
         n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
         n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577,
         n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
         n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
         n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
         n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
         n38610;
  wire   [511:0] sreg;

  DFF \sreg_reg[479]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U35 ( .A(n3829), .B(n3828), .Z(n1) );
  NANDN U36 ( .A(n3827), .B(n3826), .Z(n2) );
  AND U37 ( .A(n1), .B(n2), .Z(n3981) );
  NAND U38 ( .A(n3822), .B(n3823), .Z(n3) );
  NANDN U39 ( .A(n3825), .B(n3824), .Z(n4) );
  NAND U40 ( .A(n3), .B(n4), .Z(n3982) );
  NAND U41 ( .A(n17089), .B(n17090), .Z(n5) );
  NANDN U42 ( .A(n17088), .B(n17087), .Z(n6) );
  NAND U43 ( .A(n5), .B(n6), .Z(n17274) );
  NAND U44 ( .A(n17555), .B(n17554), .Z(n7) );
  NANDN U45 ( .A(n17553), .B(n17552), .Z(n8) );
  AND U46 ( .A(n7), .B(n8), .Z(n17655) );
  NAND U47 ( .A(n34650), .B(n34651), .Z(n9) );
  NANDN U48 ( .A(n34649), .B(n34648), .Z(n10) );
  NAND U49 ( .A(n9), .B(n10), .Z(n34823) );
  NAND U50 ( .A(n37646), .B(n37645), .Z(n11) );
  NANDN U51 ( .A(n37644), .B(n37643), .Z(n12) );
  AND U52 ( .A(n11), .B(n12), .Z(n37728) );
  NAND U53 ( .A(n36878), .B(n36877), .Z(n13) );
  NANDN U54 ( .A(n36876), .B(n36875), .Z(n14) );
  AND U55 ( .A(n13), .B(n14), .Z(n36886) );
  NAND U56 ( .A(n37532), .B(n37531), .Z(n15) );
  NANDN U57 ( .A(n37530), .B(n37529), .Z(n16) );
  AND U58 ( .A(n15), .B(n16), .Z(n37548) );
  NAND U59 ( .A(n37715), .B(n37714), .Z(n17) );
  NANDN U60 ( .A(n37713), .B(n37712), .Z(n18) );
  AND U61 ( .A(n17), .B(n18), .Z(n37727) );
  XNOR U62 ( .A(n4254), .B(n4253), .Z(n4255) );
  XNOR U63 ( .A(n4684), .B(n4683), .Z(n4685) );
  XNOR U64 ( .A(n5977), .B(n5976), .Z(n5978) );
  XNOR U65 ( .A(n6269), .B(n6268), .Z(n6270) );
  XNOR U66 ( .A(n8200), .B(n8199), .Z(n8201) );
  XNOR U67 ( .A(n10115), .B(n10114), .Z(n10116) );
  XNOR U68 ( .A(n10679), .B(n10678), .Z(n10680) );
  XNOR U69 ( .A(n12733), .B(n12732), .Z(n12734) );
  XNOR U70 ( .A(n14198), .B(n14197), .Z(n14199) );
  XNOR U71 ( .A(n14794), .B(n14793), .Z(n14795) );
  XNOR U72 ( .A(n16551), .B(n16550), .Z(n16552) );
  XNOR U73 ( .A(n18268), .B(n18267), .Z(n18269) );
  XNOR U74 ( .A(n18556), .B(n18555), .Z(n18557) );
  XNOR U75 ( .A(n19709), .B(n19708), .Z(n19710) );
  XNOR U76 ( .A(n20149), .B(n20148), .Z(n20150) );
  XNOR U77 ( .A(n20722), .B(n20721), .Z(n20723) );
  XNOR U78 ( .A(n21304), .B(n21303), .Z(n21305) );
  XNOR U79 ( .A(n21739), .B(n21738), .Z(n21740) );
  XNOR U80 ( .A(n22919), .B(n22918), .Z(n22920) );
  XNOR U81 ( .A(n23193), .B(n23192), .Z(n23194) );
  XNOR U82 ( .A(n24353), .B(n24352), .Z(n24354) );
  XNOR U83 ( .A(n25081), .B(n25080), .Z(n25082) );
  XNOR U84 ( .A(n26260), .B(n26259), .Z(n26261) );
  XNOR U85 ( .A(n27851), .B(n27850), .Z(n27852) );
  XNOR U86 ( .A(n29166), .B(n29165), .Z(n29167) );
  XNOR U87 ( .A(n29452), .B(n29451), .Z(n29453) );
  XNOR U88 ( .A(n29746), .B(n29745), .Z(n29747) );
  XNOR U89 ( .A(n30022), .B(n30021), .Z(n30023) );
  XNOR U90 ( .A(n30745), .B(n30744), .Z(n30746) );
  XNOR U91 ( .A(n31909), .B(n31908), .Z(n31910) );
  XNOR U92 ( .A(n33652), .B(n33651), .Z(n33653) );
  XNOR U93 ( .A(n35259), .B(n35258), .Z(n35260) );
  NAND U94 ( .A(n2670), .B(n2669), .Z(n19) );
  NANDN U95 ( .A(n2668), .B(n2667), .Z(n20) );
  NAND U96 ( .A(n19), .B(n20), .Z(n2720) );
  NAND U97 ( .A(n3669), .B(n3670), .Z(n21) );
  NANDN U98 ( .A(n3672), .B(n3671), .Z(n22) );
  AND U99 ( .A(n21), .B(n22), .Z(n3890) );
  NANDN U100 ( .A(n3819), .B(n3818), .Z(n23) );
  NANDN U101 ( .A(n3821), .B(n3820), .Z(n24) );
  NAND U102 ( .A(n23), .B(n24), .Z(n3983) );
  NAND U103 ( .A(n4249), .B(n4250), .Z(n25) );
  NANDN U104 ( .A(n4252), .B(n4251), .Z(n26) );
  AND U105 ( .A(n25), .B(n26), .Z(n4415) );
  NAND U106 ( .A(n4414), .B(n4413), .Z(n27) );
  NANDN U107 ( .A(n4412), .B(n4411), .Z(n28) );
  AND U108 ( .A(n27), .B(n28), .Z(n4500) );
  NAND U109 ( .A(n4603), .B(n4602), .Z(n29) );
  NANDN U110 ( .A(n4601), .B(n4600), .Z(n30) );
  AND U111 ( .A(n29), .B(n30), .Z(n4689) );
  NAND U112 ( .A(n4679), .B(n4680), .Z(n31) );
  NANDN U113 ( .A(n4682), .B(n4681), .Z(n32) );
  AND U114 ( .A(n31), .B(n32), .Z(n4836) );
  NAND U115 ( .A(n4826), .B(n4827), .Z(n33) );
  NANDN U116 ( .A(n4829), .B(n4828), .Z(n34) );
  AND U117 ( .A(n33), .B(n34), .Z(n4975) );
  NAND U118 ( .A(n4974), .B(n4973), .Z(n35) );
  NANDN U119 ( .A(n4972), .B(n4971), .Z(n36) );
  AND U120 ( .A(n35), .B(n36), .Z(n5108) );
  NAND U121 ( .A(n5972), .B(n5973), .Z(n37) );
  NANDN U122 ( .A(n5975), .B(n5974), .Z(n38) );
  AND U123 ( .A(n37), .B(n38), .Z(n6141) );
  NAND U124 ( .A(n6264), .B(n6265), .Z(n39) );
  NANDN U125 ( .A(n6267), .B(n6266), .Z(n40) );
  AND U126 ( .A(n39), .B(n40), .Z(n6433) );
  NAND U127 ( .A(n8195), .B(n8196), .Z(n41) );
  NANDN U128 ( .A(n8198), .B(n8197), .Z(n42) );
  AND U129 ( .A(n41), .B(n42), .Z(n8352) );
  XNOR U130 ( .A(n9825), .B(n9826), .Z(n9828) );
  NAND U131 ( .A(n10110), .B(n10111), .Z(n43) );
  NANDN U132 ( .A(n10113), .B(n10112), .Z(n44) );
  AND U133 ( .A(n43), .B(n44), .Z(n10265) );
  NAND U134 ( .A(n10264), .B(n10263), .Z(n45) );
  NANDN U135 ( .A(n10262), .B(n10261), .Z(n46) );
  AND U136 ( .A(n45), .B(n46), .Z(n10398) );
  XOR U137 ( .A(n10737), .B(n10738), .Z(n10739) );
  NAND U138 ( .A(n10674), .B(n10675), .Z(n47) );
  NANDN U139 ( .A(n10677), .B(n10676), .Z(n48) );
  AND U140 ( .A(n47), .B(n48), .Z(n10840) );
  NAND U141 ( .A(n11563), .B(n11562), .Z(n49) );
  NANDN U142 ( .A(n11561), .B(n11560), .Z(n50) );
  AND U143 ( .A(n49), .B(n50), .Z(n11713) );
  NAND U144 ( .A(n12590), .B(n12589), .Z(n51) );
  NANDN U145 ( .A(n12588), .B(n12587), .Z(n52) );
  AND U146 ( .A(n51), .B(n52), .Z(n12738) );
  NAND U147 ( .A(n12728), .B(n12729), .Z(n53) );
  NANDN U148 ( .A(n12731), .B(n12730), .Z(n54) );
  AND U149 ( .A(n53), .B(n54), .Z(n12893) );
  NAND U150 ( .A(n14193), .B(n14194), .Z(n55) );
  NANDN U151 ( .A(n14196), .B(n14195), .Z(n56) );
  AND U152 ( .A(n55), .B(n56), .Z(n14360) );
  XNOR U153 ( .A(n14642), .B(n14643), .Z(n14645) );
  NAND U154 ( .A(n14789), .B(n14790), .Z(n57) );
  NANDN U155 ( .A(n14792), .B(n14791), .Z(n58) );
  AND U156 ( .A(n57), .B(n58), .Z(n14942) );
  NAND U157 ( .A(n14941), .B(n14940), .Z(n59) );
  NANDN U158 ( .A(n14939), .B(n14938), .Z(n60) );
  AND U159 ( .A(n59), .B(n60), .Z(n15027) );
  NAND U160 ( .A(n16093), .B(n16094), .Z(n61) );
  NANDN U161 ( .A(n16096), .B(n16095), .Z(n62) );
  AND U162 ( .A(n61), .B(n62), .Z(n16262) );
  NAND U163 ( .A(n16546), .B(n16547), .Z(n63) );
  NANDN U164 ( .A(n16549), .B(n16548), .Z(n64) );
  AND U165 ( .A(n63), .B(n64), .Z(n16699) );
  NAND U166 ( .A(n16698), .B(n16697), .Z(n65) );
  NANDN U167 ( .A(n16696), .B(n16695), .Z(n66) );
  AND U168 ( .A(n65), .B(n66), .Z(n16832) );
  NAND U169 ( .A(n17085), .B(n17086), .Z(n67) );
  NANDN U170 ( .A(n17084), .B(n17083), .Z(n68) );
  NAND U171 ( .A(n67), .B(n68), .Z(n17275) );
  NAND U172 ( .A(n17756), .B(n17755), .Z(n69) );
  NANDN U173 ( .A(n17754), .B(n17753), .Z(n70) );
  AND U174 ( .A(n69), .B(n70), .Z(n17843) );
  NAND U175 ( .A(n18263), .B(n18264), .Z(n71) );
  NANDN U176 ( .A(n18266), .B(n18265), .Z(n72) );
  AND U177 ( .A(n71), .B(n72), .Z(n18430) );
  NAND U178 ( .A(n18429), .B(n18428), .Z(n73) );
  NANDN U179 ( .A(n18427), .B(n18426), .Z(n74) );
  AND U180 ( .A(n73), .B(n74), .Z(n18561) );
  NAND U181 ( .A(n18551), .B(n18552), .Z(n75) );
  NANDN U182 ( .A(n18554), .B(n18553), .Z(n76) );
  AND U183 ( .A(n75), .B(n76), .Z(n18712) );
  NAND U184 ( .A(n18702), .B(n18703), .Z(n77) );
  NANDN U185 ( .A(n18705), .B(n18704), .Z(n78) );
  AND U186 ( .A(n77), .B(n78), .Z(n18851) );
  NAND U187 ( .A(n18850), .B(n18849), .Z(n79) );
  NANDN U188 ( .A(n18848), .B(n18847), .Z(n80) );
  AND U189 ( .A(n79), .B(n80), .Z(n18936) );
  NAND U190 ( .A(n19566), .B(n19565), .Z(n81) );
  NANDN U191 ( .A(n19564), .B(n19563), .Z(n82) );
  AND U192 ( .A(n81), .B(n82), .Z(n19714) );
  NAND U193 ( .A(n19704), .B(n19705), .Z(n83) );
  NANDN U194 ( .A(n19707), .B(n19706), .Z(n84) );
  AND U195 ( .A(n83), .B(n84), .Z(n19865) );
  NAND U196 ( .A(n20144), .B(n20145), .Z(n85) );
  NANDN U197 ( .A(n20147), .B(n20146), .Z(n86) );
  AND U198 ( .A(n85), .B(n86), .Z(n20302) );
  NAND U199 ( .A(n20717), .B(n20718), .Z(n87) );
  NANDN U200 ( .A(n20720), .B(n20719), .Z(n88) );
  AND U201 ( .A(n87), .B(n88), .Z(n20884) );
  NAND U202 ( .A(n21299), .B(n21300), .Z(n89) );
  NANDN U203 ( .A(n21302), .B(n21301), .Z(n90) );
  AND U204 ( .A(n89), .B(n90), .Z(n21466) );
  NAND U205 ( .A(n21734), .B(n21735), .Z(n91) );
  NANDN U206 ( .A(n21737), .B(n21736), .Z(n92) );
  AND U207 ( .A(n91), .B(n92), .Z(n21899) );
  NAND U208 ( .A(n21898), .B(n21897), .Z(n93) );
  NANDN U209 ( .A(n21896), .B(n21895), .Z(n94) );
  AND U210 ( .A(n93), .B(n94), .Z(n22032) );
  NAND U211 ( .A(n22914), .B(n22915), .Z(n95) );
  NANDN U212 ( .A(n22917), .B(n22916), .Z(n96) );
  AND U213 ( .A(n95), .B(n96), .Z(n23067) );
  NAND U214 ( .A(n23066), .B(n23065), .Z(n97) );
  NANDN U215 ( .A(n23064), .B(n23063), .Z(n98) );
  AND U216 ( .A(n97), .B(n98), .Z(n23198) );
  NAND U217 ( .A(n23188), .B(n23189), .Z(n99) );
  NANDN U218 ( .A(n23191), .B(n23190), .Z(n100) );
  AND U219 ( .A(n99), .B(n100), .Z(n23349) );
  NAND U220 ( .A(n23348), .B(n23347), .Z(n101) );
  NANDN U221 ( .A(n23346), .B(n23345), .Z(n102) );
  AND U222 ( .A(n101), .B(n102), .Z(n23433) );
  NAND U223 ( .A(n23534), .B(n23533), .Z(n103) );
  NANDN U224 ( .A(n23532), .B(n23531), .Z(n104) );
  AND U225 ( .A(n103), .B(n104), .Z(n23622) );
  NAND U226 ( .A(n24210), .B(n24209), .Z(n105) );
  NANDN U227 ( .A(n24208), .B(n24207), .Z(n106) );
  AND U228 ( .A(n105), .B(n106), .Z(n24358) );
  NAND U229 ( .A(n24348), .B(n24349), .Z(n107) );
  NANDN U230 ( .A(n24351), .B(n24350), .Z(n108) );
  AND U231 ( .A(n107), .B(n108), .Z(n24513) );
  NAND U232 ( .A(n25076), .B(n25077), .Z(n109) );
  NANDN U233 ( .A(n25079), .B(n25078), .Z(n110) );
  AND U234 ( .A(n109), .B(n110), .Z(n25244) );
  NAND U235 ( .A(n25683), .B(n25682), .Z(n111) );
  NANDN U236 ( .A(n25681), .B(n25680), .Z(n112) );
  AND U237 ( .A(n111), .B(n112), .Z(n25821) );
  NAND U238 ( .A(n26255), .B(n26256), .Z(n113) );
  NANDN U239 ( .A(n26258), .B(n26257), .Z(n114) );
  AND U240 ( .A(n113), .B(n114), .Z(n26410) );
  NAND U241 ( .A(n26409), .B(n26408), .Z(n115) );
  NANDN U242 ( .A(n26407), .B(n26406), .Z(n116) );
  AND U243 ( .A(n115), .B(n116), .Z(n26495) );
  NAND U244 ( .A(n26596), .B(n26595), .Z(n117) );
  NANDN U245 ( .A(n26594), .B(n26593), .Z(n118) );
  AND U246 ( .A(n117), .B(n118), .Z(n26684) );
  NAND U247 ( .A(n27846), .B(n27847), .Z(n119) );
  NANDN U248 ( .A(n27849), .B(n27848), .Z(n120) );
  AND U249 ( .A(n119), .B(n120), .Z(n28015) );
  NAND U250 ( .A(n28751), .B(n28750), .Z(n121) );
  NANDN U251 ( .A(n28749), .B(n28748), .Z(n122) );
  AND U252 ( .A(n121), .B(n122), .Z(n28839) );
  XNOR U253 ( .A(n29171), .B(n29172), .Z(n29174) );
  NAND U254 ( .A(n29161), .B(n29162), .Z(n123) );
  NANDN U255 ( .A(n29164), .B(n29163), .Z(n124) );
  AND U256 ( .A(n123), .B(n124), .Z(n29326) );
  NAND U257 ( .A(n29325), .B(n29324), .Z(n125) );
  NANDN U258 ( .A(n29323), .B(n29322), .Z(n126) );
  AND U259 ( .A(n125), .B(n126), .Z(n29457) );
  NAND U260 ( .A(n29447), .B(n29448), .Z(n127) );
  NANDN U261 ( .A(n29450), .B(n29449), .Z(n128) );
  AND U262 ( .A(n127), .B(n128), .Z(n29610) );
  NAND U263 ( .A(n29741), .B(n29742), .Z(n129) );
  NANDN U264 ( .A(n29744), .B(n29743), .Z(n130) );
  AND U265 ( .A(n129), .B(n130), .Z(n29896) );
  NAND U266 ( .A(n30017), .B(n30018), .Z(n131) );
  NANDN U267 ( .A(n30020), .B(n30019), .Z(n132) );
  AND U268 ( .A(n131), .B(n132), .Z(n30182) );
  NAND U269 ( .A(n30181), .B(n30180), .Z(n133) );
  NANDN U270 ( .A(n30179), .B(n30178), .Z(n134) );
  AND U271 ( .A(n133), .B(n134), .Z(n30267) );
  NAND U272 ( .A(n30368), .B(n30367), .Z(n135) );
  NANDN U273 ( .A(n30366), .B(n30365), .Z(n136) );
  AND U274 ( .A(n135), .B(n136), .Z(n30456) );
  NAND U275 ( .A(n30740), .B(n30741), .Z(n137) );
  NANDN U276 ( .A(n30743), .B(n30742), .Z(n138) );
  AND U277 ( .A(n137), .B(n138), .Z(n30895) );
  NAND U278 ( .A(n31185), .B(n31184), .Z(n139) );
  NANDN U279 ( .A(n31183), .B(n31182), .Z(n140) );
  AND U280 ( .A(n139), .B(n140), .Z(n31323) );
  NAND U281 ( .A(n31904), .B(n31905), .Z(n141) );
  NANDN U282 ( .A(n31907), .B(n31906), .Z(n142) );
  AND U283 ( .A(n141), .B(n142), .Z(n32059) );
  NAND U284 ( .A(n32049), .B(n32050), .Z(n143) );
  NANDN U285 ( .A(n32052), .B(n32051), .Z(n144) );
  AND U286 ( .A(n143), .B(n144), .Z(n32202) );
  XNOR U287 ( .A(n33082), .B(n33083), .Z(n33085) );
  NAND U288 ( .A(n33511), .B(n33510), .Z(n145) );
  NANDN U289 ( .A(n33509), .B(n33508), .Z(n146) );
  AND U290 ( .A(n145), .B(n146), .Z(n33657) );
  NAND U291 ( .A(n33647), .B(n33648), .Z(n147) );
  NANDN U292 ( .A(n33650), .B(n33649), .Z(n148) );
  AND U293 ( .A(n147), .B(n148), .Z(n33806) );
  NAND U294 ( .A(n33805), .B(n33804), .Z(n149) );
  NANDN U295 ( .A(n33803), .B(n33802), .Z(n150) );
  AND U296 ( .A(n149), .B(n150), .Z(n33937) );
  NAND U297 ( .A(n34646), .B(n34647), .Z(n151) );
  NANDN U298 ( .A(n34645), .B(n34644), .Z(n152) );
  NAND U299 ( .A(n151), .B(n152), .Z(n34824) );
  NAND U300 ( .A(n35254), .B(n35255), .Z(n153) );
  NANDN U301 ( .A(n35257), .B(n35256), .Z(n154) );
  AND U302 ( .A(n153), .B(n154), .Z(n35410) );
  XNOR U303 ( .A(n35651), .B(n35650), .Z(n35652) );
  NAND U304 ( .A(n35400), .B(n35401), .Z(n155) );
  NANDN U305 ( .A(n35403), .B(n35402), .Z(n156) );
  AND U306 ( .A(n155), .B(n156), .Z(n35553) );
  NAND U307 ( .A(n36420), .B(n36419), .Z(n157) );
  NAND U308 ( .A(n36417), .B(n36418), .Z(n158) );
  NAND U309 ( .A(n157), .B(n158), .Z(n36538) );
  NAND U310 ( .A(n1613), .B(n1612), .Z(n159) );
  NANDN U311 ( .A(n1611), .B(n1610), .Z(n160) );
  NAND U312 ( .A(n159), .B(n160), .Z(n1649) );
  NAND U313 ( .A(n1847), .B(n1846), .Z(n161) );
  NANDN U314 ( .A(n1845), .B(n1844), .Z(n162) );
  AND U315 ( .A(n161), .B(n162), .Z(n1870) );
  NAND U316 ( .A(n17912), .B(n17913), .Z(n163) );
  NANDN U317 ( .A(n17911), .B(n17910), .Z(n164) );
  NAND U318 ( .A(n163), .B(n164), .Z(n17929) );
  NAND U319 ( .A(n37480), .B(n37479), .Z(n165) );
  NAND U320 ( .A(n37477), .B(n37478), .Z(n166) );
  NAND U321 ( .A(n165), .B(n166), .Z(n37561) );
  NAND U322 ( .A(n37462), .B(n37461), .Z(n167) );
  NANDN U323 ( .A(n37460), .B(n37459), .Z(n168) );
  AND U324 ( .A(n167), .B(n168), .Z(n37555) );
  NAND U325 ( .A(n37642), .B(n37641), .Z(n169) );
  NANDN U326 ( .A(n37640), .B(n37639), .Z(n170) );
  NAND U327 ( .A(n169), .B(n170), .Z(n37729) );
  NAND U328 ( .A(n37860), .B(n37859), .Z(n171) );
  NANDN U329 ( .A(n37858), .B(n37857), .Z(n172) );
  NAND U330 ( .A(n171), .B(n172), .Z(n37893) );
  NAND U331 ( .A(n38198), .B(n38197), .Z(n173) );
  NANDN U332 ( .A(n38196), .B(n38290), .Z(n174) );
  NAND U333 ( .A(n173), .B(n174), .Z(n38247) );
  XOR U334 ( .A(n1110), .B(n1109), .Z(n175) );
  NANDN U335 ( .A(n1108), .B(n175), .Z(n176) );
  NAND U336 ( .A(n1110), .B(n1109), .Z(n177) );
  AND U337 ( .A(n176), .B(n177), .Z(n1137) );
  NAND U338 ( .A(n5635), .B(n5634), .Z(n178) );
  NAND U339 ( .A(n5632), .B(n5633), .Z(n179) );
  NAND U340 ( .A(n178), .B(n179), .Z(n5782) );
  NAND U341 ( .A(n17787), .B(n17786), .Z(n180) );
  NAND U342 ( .A(n17784), .B(n17785), .Z(n181) );
  NAND U343 ( .A(n180), .B(n181), .Z(n17928) );
  NAND U344 ( .A(n37454), .B(n37453), .Z(n182) );
  NANDN U345 ( .A(n37452), .B(n37451), .Z(n183) );
  NAND U346 ( .A(n182), .B(n183), .Z(n37551) );
  NAND U347 ( .A(n36882), .B(n36881), .Z(n184) );
  NANDN U348 ( .A(n36880), .B(n36879), .Z(n185) );
  AND U349 ( .A(n184), .B(n185), .Z(n37002) );
  NANDN U350 ( .A(n37802), .B(n37800), .Z(n186) );
  NAND U351 ( .A(n37802), .B(n37799), .Z(n187) );
  NANDN U352 ( .A(n37801), .B(n187), .Z(n188) );
  NAND U353 ( .A(n186), .B(n188), .Z(n37806) );
  NAND U354 ( .A(n3291), .B(n3290), .Z(n189) );
  NANDN U355 ( .A(n3289), .B(n3288), .Z(n190) );
  AND U356 ( .A(n189), .B(n190), .Z(n3412) );
  XNOR U357 ( .A(n4114), .B(n4115), .Z(n4117) );
  XNOR U358 ( .A(n4583), .B(n4582), .Z(n4584) );
  XNOR U359 ( .A(n4831), .B(n4830), .Z(n4832) );
  XNOR U360 ( .A(n5384), .B(n5385), .Z(n5387) );
  XNOR U361 ( .A(n5513), .B(n5514), .Z(n5516) );
  XNOR U362 ( .A(n5507), .B(n5508), .Z(n5510) );
  XNOR U363 ( .A(n5660), .B(n5661), .Z(n5663) );
  XNOR U364 ( .A(n5654), .B(n5655), .Z(n5657) );
  XNOR U365 ( .A(n5807), .B(n5808), .Z(n5810) );
  XNOR U366 ( .A(n5801), .B(n5802), .Z(n5804) );
  XNOR U367 ( .A(n6111), .B(n6112), .Z(n6114) );
  XNOR U368 ( .A(n6105), .B(n6106), .Z(n6108) );
  XNOR U369 ( .A(n6566), .B(n6567), .Z(n6569) );
  XNOR U370 ( .A(n7011), .B(n7012), .Z(n7014) );
  XOR U371 ( .A(n7115), .B(n7116), .Z(n7117) );
  XOR U372 ( .A(n7109), .B(n7110), .Z(n7111) );
  XNOR U373 ( .A(n7602), .B(n7603), .Z(n7605) );
  XNOR U374 ( .A(n7731), .B(n7732), .Z(n7734) );
  XNOR U375 ( .A(n7725), .B(n7726), .Z(n7728) );
  XNOR U376 ( .A(n8028), .B(n8029), .Z(n8031) );
  XNOR U377 ( .A(n8022), .B(n8023), .Z(n8025) );
  XNOR U378 ( .A(n8777), .B(n8778), .Z(n8780) );
  XNOR U379 ( .A(n9223), .B(n9224), .Z(n9226) );
  XNOR U380 ( .A(n9350), .B(n9351), .Z(n9353) );
  XNOR U381 ( .A(n9344), .B(n9345), .Z(n9347) );
  XNOR U382 ( .A(n9813), .B(n9814), .Z(n9816) );
  XNOR U383 ( .A(n9943), .B(n9944), .Z(n9946) );
  XNOR U384 ( .A(n9937), .B(n9938), .Z(n9940) );
  XNOR U385 ( .A(n10386), .B(n10387), .Z(n10389) );
  XNOR U386 ( .A(n11124), .B(n11125), .Z(n11127) );
  XNOR U387 ( .A(n11241), .B(n11242), .Z(n11244) );
  XNOR U388 ( .A(n11235), .B(n11236), .Z(n11238) );
  XNOR U389 ( .A(n11389), .B(n11390), .Z(n11392) );
  XNOR U390 ( .A(n11383), .B(n11384), .Z(n11386) );
  XNOR U391 ( .A(n11543), .B(n11542), .Z(n11544) );
  XNOR U392 ( .A(n11701), .B(n11702), .Z(n11704) );
  XNOR U393 ( .A(n11999), .B(n12000), .Z(n12002) );
  XNOR U394 ( .A(n12296), .B(n12297), .Z(n12299) );
  XNOR U395 ( .A(n12415), .B(n12416), .Z(n12418) );
  XNOR U396 ( .A(n12409), .B(n12410), .Z(n12412) );
  XNOR U397 ( .A(n12881), .B(n12882), .Z(n12884) );
  XNOR U398 ( .A(n13159), .B(n13160), .Z(n13162) );
  XNOR U399 ( .A(n13605), .B(n13606), .Z(n13608) );
  XNOR U400 ( .A(n14048), .B(n14049), .Z(n14051) );
  XNOR U401 ( .A(n14630), .B(n14631), .Z(n14633) );
  XNOR U402 ( .A(n15364), .B(n15365), .Z(n15367) );
  XOR U403 ( .A(n15472), .B(n15473), .Z(n15474) );
  XOR U404 ( .A(n15466), .B(n15467), .Z(n15468) );
  XNOR U405 ( .A(n15807), .B(n15808), .Z(n15810) );
  XNOR U406 ( .A(n15938), .B(n15939), .Z(n15941) );
  XNOR U407 ( .A(n15932), .B(n15933), .Z(n15935) );
  XNOR U408 ( .A(n16397), .B(n16398), .Z(n16400) );
  XNOR U409 ( .A(n16973), .B(n16974), .Z(n16976) );
  XOR U410 ( .A(n17379), .B(n17380), .Z(n17381) );
  XNOR U411 ( .A(n17374), .B(n17373), .Z(n17375) );
  XNOR U412 ( .A(n17831), .B(n17832), .Z(n17834) );
  XOR U413 ( .A(n17941), .B(n17942), .Z(n17943) );
  XOR U414 ( .A(n17935), .B(n17936), .Z(n17937) );
  XNOR U415 ( .A(n18110), .B(n18111), .Z(n18113) );
  XNOR U416 ( .A(n18104), .B(n18105), .Z(n18107) );
  XNOR U417 ( .A(n18707), .B(n18706), .Z(n18708) );
  XNOR U418 ( .A(n19273), .B(n19274), .Z(n19276) );
  XNOR U419 ( .A(n19392), .B(n19393), .Z(n19395) );
  XNOR U420 ( .A(n19386), .B(n19387), .Z(n19389) );
  XOR U421 ( .A(n19853), .B(n19854), .Z(n19855) );
  XNOR U422 ( .A(n19859), .B(n19860), .Z(n19862) );
  XNOR U423 ( .A(n19967), .B(n19968), .Z(n19970) );
  XNOR U424 ( .A(n19961), .B(n19962), .Z(n19964) );
  XNOR U425 ( .A(n20582), .B(n20583), .Z(n20585) );
  XNOR U426 ( .A(n21152), .B(n21153), .Z(n21155) );
  XNOR U427 ( .A(n21599), .B(n21600), .Z(n21602) );
  XNOR U428 ( .A(n22163), .B(n22164), .Z(n22166) );
  XOR U429 ( .A(n22291), .B(n22292), .Z(n22293) );
  XOR U430 ( .A(n22285), .B(n22286), .Z(n22287) );
  XNOR U431 ( .A(n22440), .B(n22441), .Z(n22443) );
  XNOR U432 ( .A(n22434), .B(n22435), .Z(n22437) );
  XNOR U433 ( .A(n22765), .B(n22766), .Z(n22768) );
  XNOR U434 ( .A(n23610), .B(n23611), .Z(n23613) );
  XNOR U435 ( .A(n23901), .B(n23902), .Z(n23904) );
  XNOR U436 ( .A(n24045), .B(n24046), .Z(n24048) );
  XNOR U437 ( .A(n24039), .B(n24040), .Z(n24042) );
  XOR U438 ( .A(n24615), .B(n24616), .Z(n24617) );
  XOR U439 ( .A(n24609), .B(n24610), .Z(n24611) );
  XNOR U440 ( .A(n24927), .B(n24928), .Z(n24930) );
  XNOR U441 ( .A(n25377), .B(n25378), .Z(n25380) );
  XNOR U442 ( .A(n25507), .B(n25508), .Z(n25510) );
  XNOR U443 ( .A(n25501), .B(n25502), .Z(n25504) );
  XNOR U444 ( .A(n25809), .B(n25810), .Z(n25812) );
  XOR U445 ( .A(n25931), .B(n25932), .Z(n25933) );
  XOR U446 ( .A(n25925), .B(n25926), .Z(n25927) );
  XNOR U447 ( .A(n26080), .B(n26081), .Z(n26083) );
  XNOR U448 ( .A(n26074), .B(n26075), .Z(n26077) );
  XNOR U449 ( .A(n26576), .B(n26575), .Z(n26577) );
  XNOR U450 ( .A(n26811), .B(n26812), .Z(n26814) );
  XNOR U451 ( .A(n27118), .B(n27119), .Z(n27121) );
  XNOR U452 ( .A(n27564), .B(n27565), .Z(n27567) );
  XNOR U453 ( .A(n27681), .B(n27682), .Z(n27684) );
  XNOR U454 ( .A(n27675), .B(n27676), .Z(n27678) );
  XNOR U455 ( .A(n28003), .B(n28004), .Z(n28006) );
  XNOR U456 ( .A(n28130), .B(n28131), .Z(n28133) );
  XNOR U457 ( .A(n28124), .B(n28125), .Z(n28127) );
  XNOR U458 ( .A(n28583), .B(n28584), .Z(n28586) );
  XNOR U459 ( .A(n28731), .B(n28730), .Z(n28732) );
  XOR U460 ( .A(n28996), .B(n28997), .Z(n28998) );
  XNOR U461 ( .A(n28991), .B(n28990), .Z(n28992) );
  XNOR U462 ( .A(n29598), .B(n29599), .Z(n29601) );
  XNOR U463 ( .A(n29884), .B(n29885), .Z(n29887) );
  XNOR U464 ( .A(n30348), .B(n30347), .Z(n30349) );
  XNOR U465 ( .A(n30593), .B(n30594), .Z(n30596) );
  XNOR U466 ( .A(n30883), .B(n30884), .Z(n30886) );
  XNOR U467 ( .A(n30999), .B(n31000), .Z(n31002) );
  XNOR U468 ( .A(n30993), .B(n30994), .Z(n30996) );
  XNOR U469 ( .A(n31165), .B(n31164), .Z(n31166) );
  XNOR U470 ( .A(n31453), .B(n31454), .Z(n31456) );
  XOR U471 ( .A(n31569), .B(n31570), .Z(n31571) );
  XOR U472 ( .A(n31563), .B(n31564), .Z(n31565) );
  XNOR U473 ( .A(n31729), .B(n31730), .Z(n31732) );
  XNOR U474 ( .A(n31723), .B(n31724), .Z(n31726) );
  XNOR U475 ( .A(n32054), .B(n32053), .Z(n32055) );
  XNOR U476 ( .A(n32190), .B(n32191), .Z(n32193) );
  XNOR U477 ( .A(n32632), .B(n32633), .Z(n32635) );
  XNOR U478 ( .A(n33070), .B(n33071), .Z(n33073) );
  XNOR U479 ( .A(n33365), .B(n33366), .Z(n33368) );
  XNOR U480 ( .A(n34213), .B(n34214), .Z(n34216) );
  XNOR U481 ( .A(n34509), .B(n34510), .Z(n34512) );
  XNOR U482 ( .A(n34813), .B(n34814), .Z(n34805) );
  XNOR U483 ( .A(n34958), .B(n34959), .Z(n34961) );
  XNOR U484 ( .A(n35077), .B(n35078), .Z(n35080) );
  XNOR U485 ( .A(n35071), .B(n35072), .Z(n35074) );
  NAND U486 ( .A(n2795), .B(n2794), .Z(n191) );
  NANDN U487 ( .A(n2793), .B(n2792), .Z(n192) );
  AND U488 ( .A(n191), .B(n192), .Z(n2833) );
  NAND U489 ( .A(n3272), .B(n3271), .Z(n193) );
  NANDN U490 ( .A(n3270), .B(n3269), .Z(n194) );
  NAND U491 ( .A(n193), .B(n194), .Z(n3364) );
  XOR U492 ( .A(n3697), .B(n3698), .Z(n3699) );
  XOR U493 ( .A(n4126), .B(n4127), .Z(n4128) );
  NAND U494 ( .A(n3994), .B(n3993), .Z(n195) );
  NANDN U495 ( .A(n3992), .B(n3991), .Z(n196) );
  NAND U496 ( .A(n195), .B(n196), .Z(n4190) );
  NAND U497 ( .A(n4428), .B(n4427), .Z(n197) );
  NANDN U498 ( .A(n4426), .B(n4425), .Z(n198) );
  NAND U499 ( .A(n197), .B(n198), .Z(n4604) );
  NAND U500 ( .A(n4702), .B(n4701), .Z(n199) );
  NANDN U501 ( .A(n4700), .B(n4699), .Z(n200) );
  NAND U502 ( .A(n199), .B(n200), .Z(n4781) );
  NAND U503 ( .A(n4988), .B(n4987), .Z(n201) );
  NANDN U504 ( .A(n4986), .B(n4985), .Z(n202) );
  NAND U505 ( .A(n201), .B(n202), .Z(n5164) );
  XOR U506 ( .A(n5261), .B(n5262), .Z(n5263) );
  NAND U507 ( .A(n5121), .B(n5120), .Z(n203) );
  NANDN U508 ( .A(n5119), .B(n5118), .Z(n204) );
  NAND U509 ( .A(n203), .B(n204), .Z(n5325) );
  XOR U510 ( .A(n5396), .B(n5397), .Z(n5398) );
  XOR U511 ( .A(n6578), .B(n6579), .Z(n6580) );
  NAND U512 ( .A(n6446), .B(n6445), .Z(n205) );
  NANDN U513 ( .A(n6444), .B(n6443), .Z(n206) );
  NAND U514 ( .A(n205), .B(n206), .Z(n6642) );
  XNOR U515 ( .A(n6862), .B(n6863), .Z(n6865) );
  XOR U516 ( .A(n7023), .B(n7024), .Z(n7025) );
  XNOR U517 ( .A(n7317), .B(n7318), .Z(n7320) );
  XNOR U518 ( .A(n7465), .B(n7466), .Z(n7468) );
  XOR U519 ( .A(n7614), .B(n7615), .Z(n7616) );
  XOR U520 ( .A(n8495), .B(n8496), .Z(n8497) );
  NAND U521 ( .A(n8365), .B(n8364), .Z(n207) );
  NANDN U522 ( .A(n8363), .B(n8362), .Z(n208) );
  NAND U523 ( .A(n207), .B(n208), .Z(n8560) );
  XOR U524 ( .A(n8642), .B(n8643), .Z(n8644) );
  XOR U525 ( .A(n8789), .B(n8790), .Z(n8791) );
  XNOR U526 ( .A(n9074), .B(n9075), .Z(n9077) );
  XOR U527 ( .A(n9235), .B(n9236), .Z(n9237) );
  NAND U528 ( .A(n10278), .B(n10277), .Z(n209) );
  NANDN U529 ( .A(n10276), .B(n10275), .Z(n210) );
  NAND U530 ( .A(n209), .B(n210), .Z(n10454) );
  NAND U531 ( .A(n10411), .B(n10410), .Z(n211) );
  NANDN U532 ( .A(n10409), .B(n10408), .Z(n212) );
  NAND U533 ( .A(n211), .B(n212), .Z(n10605) );
  NAND U534 ( .A(n10693), .B(n10692), .Z(n213) );
  NANDN U535 ( .A(n10691), .B(n10690), .Z(n214) );
  NAND U536 ( .A(n213), .B(n214), .Z(n10783) );
  XNOR U537 ( .A(n10975), .B(n10976), .Z(n10978) );
  XOR U538 ( .A(n11136), .B(n11137), .Z(n11138) );
  NAND U539 ( .A(n11726), .B(n11725), .Z(n215) );
  NANDN U540 ( .A(n11724), .B(n11723), .Z(n216) );
  NAND U541 ( .A(n215), .B(n216), .Z(n11921) );
  XNOR U542 ( .A(n12011), .B(n12012), .Z(n12014) );
  XNOR U543 ( .A(n12308), .B(n12309), .Z(n12311) );
  XNOR U544 ( .A(n13171), .B(n13172), .Z(n13174) );
  XNOR U545 ( .A(n13480), .B(n13481), .Z(n13483) );
  XOR U546 ( .A(n13617), .B(n13618), .Z(n13619) );
  XNOR U547 ( .A(n13911), .B(n13912), .Z(n13914) );
  XOR U548 ( .A(n14060), .B(n14061), .Z(n14062) );
  NAND U549 ( .A(n14373), .B(n14372), .Z(n217) );
  NANDN U550 ( .A(n14371), .B(n14370), .Z(n218) );
  NAND U551 ( .A(n217), .B(n218), .Z(n14452) );
  NAND U552 ( .A(n14955), .B(n14954), .Z(n219) );
  NANDN U553 ( .A(n14953), .B(n14952), .Z(n220) );
  NAND U554 ( .A(n219), .B(n220), .Z(n15132) );
  NAND U555 ( .A(n15040), .B(n15039), .Z(n221) );
  NANDN U556 ( .A(n15038), .B(n15037), .Z(n222) );
  NAND U557 ( .A(n221), .B(n222), .Z(n15176) );
  XNOR U558 ( .A(n15376), .B(n15377), .Z(n15379) );
  XNOR U559 ( .A(n15662), .B(n15663), .Z(n15665) );
  XNOR U560 ( .A(n15819), .B(n15820), .Z(n15822) );
  XNOR U561 ( .A(n16409), .B(n16410), .Z(n16412) );
  NAND U562 ( .A(n16712), .B(n16711), .Z(n223) );
  NANDN U563 ( .A(n16710), .B(n16709), .Z(n224) );
  NAND U564 ( .A(n223), .B(n224), .Z(n16888) );
  XOR U565 ( .A(n16985), .B(n16986), .Z(n16987) );
  NANDN U566 ( .A(n17080), .B(n17079), .Z(n225) );
  NANDN U567 ( .A(n17082), .B(n17081), .Z(n226) );
  NAND U568 ( .A(n225), .B(n226), .Z(n17276) );
  XNOR U569 ( .A(n17556), .B(n17557), .Z(n17559) );
  XNOR U570 ( .A(n18140), .B(n18141), .Z(n18143) );
  NAND U571 ( .A(n18443), .B(n18442), .Z(n227) );
  NANDN U572 ( .A(n18441), .B(n18440), .Z(n228) );
  NAND U573 ( .A(n227), .B(n228), .Z(n18618) );
  NAND U574 ( .A(n18574), .B(n18573), .Z(n229) );
  NANDN U575 ( .A(n18572), .B(n18571), .Z(n230) );
  NAND U576 ( .A(n229), .B(n230), .Z(n18657) );
  NAND U577 ( .A(n18864), .B(n18863), .Z(n231) );
  NANDN U578 ( .A(n18862), .B(n18861), .Z(n232) );
  NAND U579 ( .A(n231), .B(n232), .Z(n19041) );
  NAND U580 ( .A(n18949), .B(n18948), .Z(n233) );
  NANDN U581 ( .A(n18947), .B(n18946), .Z(n234) );
  NAND U582 ( .A(n233), .B(n234), .Z(n19085) );
  XNOR U583 ( .A(n19285), .B(n19286), .Z(n19288) );
  NAND U584 ( .A(n19878), .B(n19877), .Z(n235) );
  NANDN U585 ( .A(n19876), .B(n19875), .Z(n236) );
  NAND U586 ( .A(n235), .B(n236), .Z(n20064) );
  XOR U587 ( .A(n20447), .B(n20448), .Z(n20449) );
  NAND U588 ( .A(n20315), .B(n20314), .Z(n237) );
  NANDN U589 ( .A(n20313), .B(n20312), .Z(n238) );
  NAND U590 ( .A(n237), .B(n238), .Z(n20511) );
  XOR U591 ( .A(n20594), .B(n20595), .Z(n20596) );
  XOR U592 ( .A(n21029), .B(n21030), .Z(n21031) );
  NAND U593 ( .A(n20897), .B(n20896), .Z(n239) );
  NANDN U594 ( .A(n20895), .B(n20894), .Z(n240) );
  NAND U595 ( .A(n239), .B(n240), .Z(n21093) );
  XOR U596 ( .A(n21164), .B(n21165), .Z(n21166) );
  XOR U597 ( .A(n21611), .B(n21612), .Z(n21613) );
  NAND U598 ( .A(n21479), .B(n21478), .Z(n241) );
  NANDN U599 ( .A(n21477), .B(n21476), .Z(n242) );
  NAND U600 ( .A(n241), .B(n242), .Z(n21675) );
  NAND U601 ( .A(n21912), .B(n21911), .Z(n243) );
  NANDN U602 ( .A(n21910), .B(n21909), .Z(n244) );
  NAND U603 ( .A(n243), .B(n244), .Z(n22088) );
  XOR U604 ( .A(n22175), .B(n22176), .Z(n22177) );
  NAND U605 ( .A(n22045), .B(n22044), .Z(n245) );
  NANDN U606 ( .A(n22043), .B(n22042), .Z(n246) );
  NAND U607 ( .A(n245), .B(n246), .Z(n22240) );
  XNOR U608 ( .A(n22470), .B(n22471), .Z(n22473) );
  XNOR U609 ( .A(n22777), .B(n22778), .Z(n22780) );
  NAND U610 ( .A(n23080), .B(n23079), .Z(n247) );
  NANDN U611 ( .A(n23078), .B(n23077), .Z(n248) );
  NAND U612 ( .A(n247), .B(n248), .Z(n23255) );
  NAND U613 ( .A(n23211), .B(n23210), .Z(n249) );
  NANDN U614 ( .A(n23209), .B(n23208), .Z(n250) );
  NAND U615 ( .A(n249), .B(n250), .Z(n23294) );
  XNOR U616 ( .A(n23913), .B(n23914), .Z(n23916) );
  XNOR U617 ( .A(n24794), .B(n24795), .Z(n24797) );
  XNOR U618 ( .A(n24939), .B(n24940), .Z(n24942) );
  XOR U619 ( .A(n25389), .B(n25390), .Z(n25391) );
  NAND U620 ( .A(n25257), .B(n25256), .Z(n251) );
  NANDN U621 ( .A(n25255), .B(n25254), .Z(n252) );
  NAND U622 ( .A(n251), .B(n252), .Z(n25454) );
  XNOR U623 ( .A(n26110), .B(n26111), .Z(n26113) );
  NAND U624 ( .A(n26423), .B(n26422), .Z(n253) );
  NANDN U625 ( .A(n26421), .B(n26420), .Z(n254) );
  NAND U626 ( .A(n253), .B(n254), .Z(n26598) );
  XOR U627 ( .A(n26823), .B(n26824), .Z(n26825) );
  NAND U628 ( .A(n26697), .B(n26696), .Z(n255) );
  NANDN U629 ( .A(n26695), .B(n26694), .Z(n256) );
  NAND U630 ( .A(n255), .B(n256), .Z(n26889) );
  XNOR U631 ( .A(n27130), .B(n27131), .Z(n27133) );
  XNOR U632 ( .A(n27415), .B(n27416), .Z(n27418) );
  XOR U633 ( .A(n27576), .B(n27577), .Z(n27578) );
  NAND U634 ( .A(n28028), .B(n28027), .Z(n257) );
  NANDN U635 ( .A(n28026), .B(n28025), .Z(n258) );
  NAND U636 ( .A(n257), .B(n258), .Z(n28227) );
  XNOR U637 ( .A(n28458), .B(n28459), .Z(n28461) );
  XOR U638 ( .A(n28595), .B(n28596), .Z(n28597) );
  NAND U639 ( .A(n28852), .B(n28851), .Z(n259) );
  NANDN U640 ( .A(n28850), .B(n28849), .Z(n260) );
  NAND U641 ( .A(n259), .B(n260), .Z(n28985) );
  NAND U642 ( .A(n29339), .B(n29338), .Z(n261) );
  NANDN U643 ( .A(n29337), .B(n29336), .Z(n262) );
  NAND U644 ( .A(n261), .B(n262), .Z(n29513) );
  NAND U645 ( .A(n29470), .B(n29469), .Z(n263) );
  NANDN U646 ( .A(n29468), .B(n29467), .Z(n264) );
  NAND U647 ( .A(n263), .B(n264), .Z(n29553) );
  NAND U648 ( .A(n29909), .B(n29908), .Z(n265) );
  NANDN U649 ( .A(n29907), .B(n29906), .Z(n266) );
  NAND U650 ( .A(n265), .B(n266), .Z(n30092) );
  NAND U651 ( .A(n30195), .B(n30194), .Z(n267) );
  NANDN U652 ( .A(n30193), .B(n30192), .Z(n268) );
  NAND U653 ( .A(n267), .B(n268), .Z(n30370) );
  XOR U654 ( .A(n30605), .B(n30606), .Z(n30607) );
  NAND U655 ( .A(n30469), .B(n30468), .Z(n269) );
  NANDN U656 ( .A(n30467), .B(n30466), .Z(n270) );
  NAND U657 ( .A(n269), .B(n270), .Z(n30669) );
  NAND U658 ( .A(n30908), .B(n30907), .Z(n271) );
  NANDN U659 ( .A(n30906), .B(n30905), .Z(n272) );
  NAND U660 ( .A(n271), .B(n272), .Z(n31096) );
  XOR U661 ( .A(n31465), .B(n31466), .Z(n31467) );
  NAND U662 ( .A(n31336), .B(n31335), .Z(n273) );
  NANDN U663 ( .A(n31334), .B(n31333), .Z(n274) );
  NAND U664 ( .A(n273), .B(n274), .Z(n31530) );
  XNOR U665 ( .A(n31759), .B(n31760), .Z(n31762) );
  NAND U666 ( .A(n32072), .B(n32071), .Z(n275) );
  NANDN U667 ( .A(n32070), .B(n32069), .Z(n276) );
  NAND U668 ( .A(n275), .B(n276), .Z(n32144) );
  NAND U669 ( .A(n32215), .B(n32214), .Z(n277) );
  NANDN U670 ( .A(n32213), .B(n32212), .Z(n278) );
  NAND U671 ( .A(n277), .B(n278), .Z(n32403) );
  XNOR U672 ( .A(n32483), .B(n32484), .Z(n32486) );
  XOR U673 ( .A(n32644), .B(n32645), .Z(n32646) );
  NAND U674 ( .A(n32777), .B(n32776), .Z(n279) );
  NANDN U675 ( .A(n32775), .B(n32774), .Z(n280) );
  AND U676 ( .A(n279), .B(n280), .Z(n32925) );
  XNOR U677 ( .A(n33377), .B(n33378), .Z(n33380) );
  NAND U678 ( .A(n33819), .B(n33818), .Z(n281) );
  NANDN U679 ( .A(n33817), .B(n33816), .Z(n282) );
  NAND U680 ( .A(n281), .B(n282), .Z(n33993) );
  XOR U681 ( .A(n34090), .B(n34091), .Z(n34092) );
  NAND U682 ( .A(n33950), .B(n33949), .Z(n283) );
  NANDN U683 ( .A(n33948), .B(n33947), .Z(n284) );
  NAND U684 ( .A(n283), .B(n284), .Z(n34154) );
  XOR U685 ( .A(n34225), .B(n34226), .Z(n34227) );
  XNOR U686 ( .A(n34521), .B(n34522), .Z(n34524) );
  NANDN U687 ( .A(n34641), .B(n34640), .Z(n285) );
  NANDN U688 ( .A(n34643), .B(n34642), .Z(n286) );
  NAND U689 ( .A(n285), .B(n286), .Z(n34825) );
  XNOR U690 ( .A(n35405), .B(n35404), .Z(n35406) );
  XNOR U691 ( .A(n2078), .B(n2079), .Z(n2083) );
  NAND U692 ( .A(n3892), .B(n3893), .Z(n287) );
  NANDN U693 ( .A(n3891), .B(n3890), .Z(n288) );
  NAND U694 ( .A(n287), .B(n288), .Z(n4044) );
  NAND U695 ( .A(n3983), .B(n3984), .Z(n289) );
  NANDN U696 ( .A(n3982), .B(n3981), .Z(n290) );
  NAND U697 ( .A(n289), .B(n290), .Z(n4073) );
  XNOR U698 ( .A(n4479), .B(n4480), .Z(n4474) );
  NAND U699 ( .A(n4417), .B(n4418), .Z(n291) );
  NANDN U700 ( .A(n4416), .B(n4415), .Z(n292) );
  NAND U701 ( .A(n291), .B(n292), .Z(n4623) );
  OR U702 ( .A(n4691), .B(n4692), .Z(n293) );
  NAND U703 ( .A(n4690), .B(n4689), .Z(n294) );
  NAND U704 ( .A(n293), .B(n294), .Z(n4892) );
  NAND U705 ( .A(n4789), .B(n4788), .Z(n295) );
  NAND U706 ( .A(n4786), .B(n4787), .Z(n296) );
  NAND U707 ( .A(n295), .B(n296), .Z(n5032) );
  NAND U708 ( .A(n4977), .B(n4978), .Z(n297) );
  NANDN U709 ( .A(n4976), .B(n4975), .Z(n298) );
  NAND U710 ( .A(n297), .B(n298), .Z(n5183) );
  OR U711 ( .A(n5110), .B(n5111), .Z(n299) );
  NAND U712 ( .A(n5109), .B(n5108), .Z(n300) );
  NAND U713 ( .A(n299), .B(n300), .Z(n5203) );
  XNOR U714 ( .A(n6207), .B(n6208), .Z(n6202) );
  NAND U715 ( .A(n6143), .B(n6144), .Z(n301) );
  NANDN U716 ( .A(n6142), .B(n6141), .Z(n302) );
  NAND U717 ( .A(n301), .B(n302), .Z(n6353) );
  XNOR U718 ( .A(n6497), .B(n6498), .Z(n6492) );
  NAND U719 ( .A(n6435), .B(n6436), .Z(n303) );
  NANDN U720 ( .A(n6434), .B(n6433), .Z(n304) );
  NAND U721 ( .A(n303), .B(n304), .Z(n6525) );
  OR U722 ( .A(n7090), .B(n7091), .Z(n305) );
  NAND U723 ( .A(n7089), .B(n7088), .Z(n306) );
  NAND U724 ( .A(n305), .B(n306), .Z(n7231) );
  XNOR U725 ( .A(n8416), .B(n8417), .Z(n8411) );
  NAND U726 ( .A(n8354), .B(n8355), .Z(n307) );
  NANDN U727 ( .A(n8353), .B(n8352), .Z(n308) );
  NAND U728 ( .A(n307), .B(n308), .Z(n8444) );
  OR U729 ( .A(n9301), .B(n9302), .Z(n309) );
  NAND U730 ( .A(n9300), .B(n9299), .Z(n310) );
  NAND U731 ( .A(n309), .B(n310), .Z(n9321) );
  NAND U732 ( .A(n9889), .B(n9888), .Z(n311) );
  NANDN U733 ( .A(n9887), .B(n9886), .Z(n312) );
  NAND U734 ( .A(n311), .B(n312), .Z(n9914) );
  XNOR U735 ( .A(n10329), .B(n10330), .Z(n10324) );
  NAND U736 ( .A(n10267), .B(n10268), .Z(n313) );
  NANDN U737 ( .A(n10266), .B(n10265), .Z(n314) );
  NAND U738 ( .A(n313), .B(n314), .Z(n10473) );
  OR U739 ( .A(n10400), .B(n10401), .Z(n315) );
  NAND U740 ( .A(n10399), .B(n10398), .Z(n316) );
  NAND U741 ( .A(n315), .B(n316), .Z(n10611) );
  XNOR U742 ( .A(n10906), .B(n10907), .Z(n10901) );
  NAND U743 ( .A(n10842), .B(n10843), .Z(n317) );
  NANDN U744 ( .A(n10841), .B(n10840), .Z(n318) );
  NAND U745 ( .A(n317), .B(n318), .Z(n11054) );
  OR U746 ( .A(n11715), .B(n11716), .Z(n319) );
  NAND U747 ( .A(n11714), .B(n11713), .Z(n320) );
  NAND U748 ( .A(n319), .B(n320), .Z(n11926) );
  OR U749 ( .A(n12740), .B(n12741), .Z(n321) );
  NAND U750 ( .A(n12739), .B(n12738), .Z(n322) );
  NAND U751 ( .A(n321), .B(n322), .Z(n12949) );
  NAND U752 ( .A(n12844), .B(n12843), .Z(n323) );
  NAND U753 ( .A(n12841), .B(n12842), .Z(n324) );
  NAND U754 ( .A(n323), .B(n324), .Z(n13097) );
  OR U755 ( .A(n14126), .B(n14127), .Z(n325) );
  NAND U756 ( .A(n14125), .B(n14124), .Z(n326) );
  NAND U757 ( .A(n325), .B(n326), .Z(n14274) );
  XNOR U758 ( .A(n14424), .B(n14425), .Z(n14419) );
  NAND U759 ( .A(n14362), .B(n14363), .Z(n327) );
  NANDN U760 ( .A(n14361), .B(n14360), .Z(n328) );
  NAND U761 ( .A(n327), .B(n328), .Z(n14572) );
  NAND U762 ( .A(n14705), .B(n14704), .Z(n329) );
  NANDN U763 ( .A(n14703), .B(n14702), .Z(n330) );
  NAND U764 ( .A(n329), .B(n330), .Z(n14742) );
  XNOR U765 ( .A(n15006), .B(n15007), .Z(n15001) );
  NAND U766 ( .A(n14944), .B(n14945), .Z(n331) );
  NANDN U767 ( .A(n14943), .B(n14942), .Z(n332) );
  NAND U768 ( .A(n331), .B(n332), .Z(n15151) );
  OR U769 ( .A(n15029), .B(n15030), .Z(n333) );
  NAND U770 ( .A(n15028), .B(n15027), .Z(n334) );
  NAND U771 ( .A(n333), .B(n334), .Z(n15289) );
  NANDN U772 ( .A(n15174), .B(n15173), .Z(n335) );
  NANDN U773 ( .A(n15172), .B(n15171), .Z(n336) );
  NAND U774 ( .A(n335), .B(n336), .Z(n15322) );
  XNOR U775 ( .A(n16328), .B(n16329), .Z(n16323) );
  NAND U776 ( .A(n16264), .B(n16265), .Z(n337) );
  NANDN U777 ( .A(n16263), .B(n16262), .Z(n338) );
  NAND U778 ( .A(n337), .B(n338), .Z(n16356) );
  XNOR U779 ( .A(n16763), .B(n16764), .Z(n16758) );
  NAND U780 ( .A(n16701), .B(n16702), .Z(n339) );
  NANDN U781 ( .A(n16700), .B(n16699), .Z(n340) );
  NAND U782 ( .A(n339), .B(n340), .Z(n16907) );
  NAND U783 ( .A(n17766), .B(n17765), .Z(n341) );
  NANDN U784 ( .A(n17764), .B(n17763), .Z(n342) );
  NAND U785 ( .A(n341), .B(n342), .Z(n17915) );
  NAND U786 ( .A(n17909), .B(n17908), .Z(n343) );
  NANDN U787 ( .A(n17907), .B(n17906), .Z(n344) );
  NAND U788 ( .A(n343), .B(n344), .Z(n18060) );
  XNOR U789 ( .A(n18494), .B(n18495), .Z(n18489) );
  NAND U790 ( .A(n18432), .B(n18433), .Z(n345) );
  NANDN U791 ( .A(n18431), .B(n18430), .Z(n346) );
  NAND U792 ( .A(n345), .B(n346), .Z(n18636) );
  OR U793 ( .A(n18563), .B(n18564), .Z(n347) );
  NAND U794 ( .A(n18562), .B(n18561), .Z(n348) );
  NAND U795 ( .A(n347), .B(n348), .Z(n18768) );
  NAND U796 ( .A(n18665), .B(n18664), .Z(n349) );
  NAND U797 ( .A(n18662), .B(n18663), .Z(n350) );
  NAND U798 ( .A(n349), .B(n350), .Z(n18908) );
  NAND U799 ( .A(n18853), .B(n18854), .Z(n351) );
  NANDN U800 ( .A(n18852), .B(n18851), .Z(n352) );
  NAND U801 ( .A(n351), .B(n352), .Z(n19060) );
  OR U802 ( .A(n18938), .B(n18939), .Z(n353) );
  NAND U803 ( .A(n18937), .B(n18936), .Z(n354) );
  NAND U804 ( .A(n353), .B(n354), .Z(n19198) );
  NANDN U805 ( .A(n19083), .B(n19082), .Z(n355) );
  NANDN U806 ( .A(n19081), .B(n19080), .Z(n356) );
  NAND U807 ( .A(n355), .B(n356), .Z(n19231) );
  NAND U808 ( .A(n19779), .B(n19778), .Z(n357) );
  NANDN U809 ( .A(n19777), .B(n19776), .Z(n358) );
  NAND U810 ( .A(n357), .B(n358), .Z(n19927) );
  NAND U811 ( .A(n19867), .B(n19868), .Z(n359) );
  NANDN U812 ( .A(n19866), .B(n19865), .Z(n360) );
  NAND U813 ( .A(n359), .B(n360), .Z(n20076) );
  XNOR U814 ( .A(n20366), .B(n20367), .Z(n20361) );
  NAND U815 ( .A(n20304), .B(n20305), .Z(n361) );
  NANDN U816 ( .A(n20303), .B(n20302), .Z(n362) );
  NAND U817 ( .A(n361), .B(n362), .Z(n20394) );
  XNOR U818 ( .A(n20948), .B(n20949), .Z(n20943) );
  NAND U819 ( .A(n20886), .B(n20887), .Z(n363) );
  NANDN U820 ( .A(n20885), .B(n20884), .Z(n364) );
  NAND U821 ( .A(n363), .B(n364), .Z(n20976) );
  XNOR U822 ( .A(n21530), .B(n21531), .Z(n21525) );
  NAND U823 ( .A(n21468), .B(n21469), .Z(n365) );
  NANDN U824 ( .A(n21467), .B(n21466), .Z(n366) );
  NAND U825 ( .A(n365), .B(n366), .Z(n21558) );
  XNOR U826 ( .A(n21963), .B(n21964), .Z(n21958) );
  NAND U827 ( .A(n21901), .B(n21902), .Z(n367) );
  NANDN U828 ( .A(n21900), .B(n21899), .Z(n368) );
  NAND U829 ( .A(n367), .B(n368), .Z(n22107) );
  OR U830 ( .A(n22034), .B(n22035), .Z(n369) );
  NAND U831 ( .A(n22033), .B(n22032), .Z(n370) );
  NAND U832 ( .A(n369), .B(n370), .Z(n22246) );
  XNOR U833 ( .A(n23131), .B(n23132), .Z(n23126) );
  NAND U834 ( .A(n23069), .B(n23070), .Z(n371) );
  NANDN U835 ( .A(n23068), .B(n23067), .Z(n372) );
  NAND U836 ( .A(n371), .B(n372), .Z(n23273) );
  OR U837 ( .A(n23200), .B(n23201), .Z(n373) );
  NAND U838 ( .A(n23199), .B(n23198), .Z(n374) );
  NAND U839 ( .A(n373), .B(n374), .Z(n23406) );
  NAND U840 ( .A(n23302), .B(n23301), .Z(n375) );
  NAND U841 ( .A(n23299), .B(n23300), .Z(n376) );
  NAND U842 ( .A(n375), .B(n376), .Z(n23548) );
  OR U843 ( .A(n23624), .B(n23625), .Z(n377) );
  NAND U844 ( .A(n23623), .B(n23622), .Z(n378) );
  NAND U845 ( .A(n377), .B(n378), .Z(n23718) );
  OR U846 ( .A(n24360), .B(n24361), .Z(n379) );
  NAND U847 ( .A(n24359), .B(n24358), .Z(n380) );
  NAND U848 ( .A(n379), .B(n380), .Z(n24570) );
  NAND U849 ( .A(n24464), .B(n24463), .Z(n381) );
  NAND U850 ( .A(n24461), .B(n24462), .Z(n382) );
  NAND U851 ( .A(n381), .B(n382), .Z(n24718) );
  XNOR U852 ( .A(n25308), .B(n25309), .Z(n25303) );
  NAND U853 ( .A(n25246), .B(n25247), .Z(n383) );
  NANDN U854 ( .A(n25245), .B(n25244), .Z(n384) );
  NAND U855 ( .A(n383), .B(n384), .Z(n25336) );
  NAND U856 ( .A(n25887), .B(n25886), .Z(n385) );
  NANDN U857 ( .A(n25885), .B(n25884), .Z(n386) );
  NAND U858 ( .A(n385), .B(n386), .Z(n25920) );
  XNOR U859 ( .A(n26474), .B(n26475), .Z(n26469) );
  NAND U860 ( .A(n26412), .B(n26413), .Z(n387) );
  NANDN U861 ( .A(n26411), .B(n26410), .Z(n388) );
  NAND U862 ( .A(n387), .B(n388), .Z(n26616) );
  OR U863 ( .A(n26686), .B(n26687), .Z(n389) );
  NAND U864 ( .A(n26685), .B(n26684), .Z(n390) );
  NAND U865 ( .A(n389), .B(n390), .Z(n26894) );
  XNOR U866 ( .A(n28079), .B(n28080), .Z(n28074) );
  NAND U867 ( .A(n28017), .B(n28018), .Z(n391) );
  NANDN U868 ( .A(n28016), .B(n28015), .Z(n392) );
  NAND U869 ( .A(n391), .B(n392), .Z(n28107) );
  OR U870 ( .A(n28841), .B(n28842), .Z(n393) );
  NAND U871 ( .A(n28840), .B(n28839), .Z(n394) );
  NAND U872 ( .A(n393), .B(n394), .Z(n29098) );
  NANDN U873 ( .A(n28983), .B(n28982), .Z(n395) );
  NANDN U874 ( .A(n28981), .B(n28980), .Z(n396) );
  NAND U875 ( .A(n395), .B(n396), .Z(n29247) );
  XNOR U876 ( .A(n29390), .B(n29391), .Z(n29385) );
  NAND U877 ( .A(n29328), .B(n29329), .Z(n397) );
  NANDN U878 ( .A(n29327), .B(n29326), .Z(n398) );
  NAND U879 ( .A(n397), .B(n398), .Z(n29532) );
  OR U880 ( .A(n29459), .B(n29460), .Z(n399) );
  NAND U881 ( .A(n29458), .B(n29457), .Z(n400) );
  NAND U882 ( .A(n399), .B(n400), .Z(n29666) );
  NAND U883 ( .A(n29561), .B(n29560), .Z(n401) );
  NAND U884 ( .A(n29558), .B(n29559), .Z(n402) );
  NAND U885 ( .A(n401), .B(n402), .Z(n29694) );
  XNOR U886 ( .A(n29960), .B(n29961), .Z(n29955) );
  NAND U887 ( .A(n29898), .B(n29899), .Z(n403) );
  NANDN U888 ( .A(n29897), .B(n29896), .Z(n404) );
  NAND U889 ( .A(n403), .B(n404), .Z(n30104) );
  XNOR U890 ( .A(n30246), .B(n30247), .Z(n30241) );
  NAND U891 ( .A(n30184), .B(n30185), .Z(n405) );
  NANDN U892 ( .A(n30183), .B(n30182), .Z(n406) );
  NAND U893 ( .A(n405), .B(n406), .Z(n30388) );
  OR U894 ( .A(n30458), .B(n30459), .Z(n407) );
  NAND U895 ( .A(n30457), .B(n30456), .Z(n408) );
  NAND U896 ( .A(n407), .B(n408), .Z(n30547) );
  XNOR U897 ( .A(n30960), .B(n30961), .Z(n30955) );
  NAND U898 ( .A(n30897), .B(n30898), .Z(n409) );
  NANDN U899 ( .A(n30896), .B(n30895), .Z(n410) );
  NAND U900 ( .A(n409), .B(n410), .Z(n31108) );
  OR U901 ( .A(n31325), .B(n31326), .Z(n411) );
  NAND U902 ( .A(n31324), .B(n31323), .Z(n412) );
  NAND U903 ( .A(n411), .B(n412), .Z(n31536) );
  XNOR U904 ( .A(n32123), .B(n32124), .Z(n32118) );
  NAND U905 ( .A(n32061), .B(n32062), .Z(n413) );
  NANDN U906 ( .A(n32060), .B(n32059), .Z(n414) );
  NAND U907 ( .A(n413), .B(n414), .Z(n32266) );
  NAND U908 ( .A(n32204), .B(n32205), .Z(n415) );
  NANDN U909 ( .A(n32203), .B(n32202), .Z(n416) );
  NAND U910 ( .A(n415), .B(n416), .Z(n32415) );
  NAND U911 ( .A(n33146), .B(n33145), .Z(n417) );
  NANDN U912 ( .A(n33144), .B(n33143), .Z(n418) );
  NAND U913 ( .A(n417), .B(n418), .Z(n33291) );
  NAND U914 ( .A(n33722), .B(n33721), .Z(n419) );
  NANDN U915 ( .A(n33720), .B(n33719), .Z(n420) );
  NAND U916 ( .A(n419), .B(n420), .Z(n33867) );
  NAND U917 ( .A(n33808), .B(n33809), .Z(n421) );
  NANDN U918 ( .A(n33807), .B(n33806), .Z(n422) );
  NAND U919 ( .A(n421), .B(n422), .Z(n34012) );
  OR U920 ( .A(n33939), .B(n33940), .Z(n423) );
  NAND U921 ( .A(n33938), .B(n33937), .Z(n424) );
  NAND U922 ( .A(n423), .B(n424), .Z(n34032) );
  XNOR U923 ( .A(n35474), .B(n35475), .Z(n35469) );
  NAND U924 ( .A(n35423), .B(n35422), .Z(n425) );
  NANDN U925 ( .A(n35421), .B(n35420), .Z(n426) );
  NAND U926 ( .A(n425), .B(n426), .Z(n35495) );
  NAND U927 ( .A(n35412), .B(n35413), .Z(n427) );
  NANDN U928 ( .A(n35411), .B(n35410), .Z(n428) );
  NAND U929 ( .A(n427), .B(n428), .Z(n35616) );
  NAND U930 ( .A(n35566), .B(n35565), .Z(n429) );
  NANDN U931 ( .A(n35564), .B(n35563), .Z(n430) );
  NAND U932 ( .A(n429), .B(n430), .Z(n35638) );
  NAND U933 ( .A(n1667), .B(n1666), .Z(n431) );
  NANDN U934 ( .A(n1665), .B(n1664), .Z(n432) );
  NAND U935 ( .A(n431), .B(n432), .Z(n1713) );
  NAND U936 ( .A(n4757), .B(n4758), .Z(n433) );
  NANDN U937 ( .A(n4756), .B(n4755), .Z(n434) );
  NAND U938 ( .A(n433), .B(n434), .Z(n4774) );
  NANDN U939 ( .A(n16928), .B(n16927), .Z(n435) );
  NANDN U940 ( .A(n16930), .B(n16929), .Z(n436) );
  NAND U941 ( .A(n435), .B(n436), .Z(n17067) );
  NANDN U942 ( .A(n18056), .B(n18055), .Z(n437) );
  NANDN U943 ( .A(n18058), .B(n18057), .Z(n438) );
  NAND U944 ( .A(n437), .B(n438), .Z(n18074) );
  NANDN U945 ( .A(n19923), .B(n19922), .Z(n439) );
  NANDN U946 ( .A(n19925), .B(n19924), .Z(n440) );
  NAND U947 ( .A(n439), .B(n440), .Z(n19943) );
  NAND U948 ( .A(n23695), .B(n23696), .Z(n441) );
  NANDN U949 ( .A(n23694), .B(n23693), .Z(n442) );
  NAND U950 ( .A(n441), .B(n442), .Z(n23712) );
  NANDN U951 ( .A(n25916), .B(n25915), .Z(n443) );
  NANDN U952 ( .A(n25918), .B(n25917), .Z(n444) );
  NAND U953 ( .A(n443), .B(n444), .Z(n26056) );
  NAND U954 ( .A(n26752), .B(n26753), .Z(n445) );
  NANDN U955 ( .A(n26751), .B(n26750), .Z(n446) );
  NAND U956 ( .A(n445), .B(n446), .Z(n26769) );
  NAND U957 ( .A(n30524), .B(n30525), .Z(n447) );
  NANDN U958 ( .A(n30523), .B(n30522), .Z(n448) );
  NAND U959 ( .A(n447), .B(n448), .Z(n30541) );
  NANDN U960 ( .A(n33863), .B(n33862), .Z(n449) );
  NANDN U961 ( .A(n33865), .B(n33864), .Z(n450) );
  NAND U962 ( .A(n449), .B(n450), .Z(n33883) );
  NAND U963 ( .A(n35555), .B(n35556), .Z(n451) );
  NANDN U964 ( .A(n35554), .B(n35553), .Z(n452) );
  NAND U965 ( .A(n451), .B(n452), .Z(n35765) );
  NAND U966 ( .A(n35914), .B(n35913), .Z(n453) );
  NANDN U967 ( .A(n35912), .B(n35911), .Z(n454) );
  NAND U968 ( .A(n453), .B(n454), .Z(n35927) );
  NAND U969 ( .A(n36088), .B(n36089), .Z(n455) );
  NANDN U970 ( .A(n36087), .B(n36086), .Z(n456) );
  NAND U971 ( .A(n455), .B(n456), .Z(n36221) );
  NAND U972 ( .A(n36786), .B(n36785), .Z(n457) );
  NANDN U973 ( .A(n36784), .B(n36783), .Z(n458) );
  NAND U974 ( .A(n457), .B(n458), .Z(n36980) );
  NAND U975 ( .A(n37199), .B(n37198), .Z(n459) );
  NANDN U976 ( .A(n37197), .B(n37269), .Z(n460) );
  NAND U977 ( .A(n459), .B(n460), .Z(n37263) );
  NAND U978 ( .A(n37650), .B(n37649), .Z(n461) );
  NANDN U979 ( .A(n37648), .B(n37647), .Z(n462) );
  NAND U980 ( .A(n461), .B(n462), .Z(n37735) );
  NANDN U981 ( .A(n1308), .B(n1307), .Z(n463) );
  NANDN U982 ( .A(n1306), .B(n1305), .Z(n464) );
  NAND U983 ( .A(n463), .B(n464), .Z(n1333) );
  NAND U984 ( .A(n1575), .B(n1574), .Z(n465) );
  NANDN U985 ( .A(n1573), .B(n1572), .Z(n466) );
  NAND U986 ( .A(n465), .B(n466), .Z(n1641) );
  NAND U987 ( .A(n3197), .B(n3196), .Z(n467) );
  NANDN U988 ( .A(n3195), .B(n3194), .Z(n468) );
  AND U989 ( .A(n467), .B(n468), .Z(n3213) );
  NAND U990 ( .A(n36512), .B(n36511), .Z(n469) );
  NANDN U991 ( .A(n36510), .B(n36509), .Z(n470) );
  NAND U992 ( .A(n469), .B(n470), .Z(n36751) );
  NAND U993 ( .A(n37557), .B(n37556), .Z(n471) );
  NANDN U994 ( .A(n37555), .B(n37554), .Z(n472) );
  NAND U995 ( .A(n471), .B(n472), .Z(n37712) );
  NAND U996 ( .A(n1868), .B(n1869), .Z(n473) );
  NANDN U997 ( .A(n1867), .B(n1866), .Z(n474) );
  NAND U998 ( .A(n473), .B(n474), .Z(n1959) );
  NAND U999 ( .A(n3632), .B(n3631), .Z(n475) );
  NANDN U1000 ( .A(n3630), .B(n3629), .Z(n476) );
  NAND U1001 ( .A(n475), .B(n476), .Z(n3777) );
  NAND U1002 ( .A(n4636), .B(n4635), .Z(n477) );
  NAND U1003 ( .A(n4633), .B(n4634), .Z(n478) );
  NAND U1004 ( .A(n477), .B(n478), .Z(n4773) );
  NAND U1005 ( .A(n5782), .B(n5781), .Z(n479) );
  NAND U1006 ( .A(n5779), .B(n5780), .Z(n480) );
  NAND U1007 ( .A(n479), .B(n480), .Z(n5929) );
  NAND U1008 ( .A(n11511), .B(n11510), .Z(n481) );
  NAND U1009 ( .A(n11508), .B(n11509), .Z(n482) );
  NAND U1010 ( .A(n481), .B(n482), .Z(n11656) );
  NAND U1011 ( .A(n11944), .B(n11943), .Z(n483) );
  NAND U1012 ( .A(n11941), .B(n11942), .Z(n484) );
  NAND U1013 ( .A(n483), .B(n484), .Z(n12092) );
  NAND U1014 ( .A(n12538), .B(n12537), .Z(n485) );
  NAND U1015 ( .A(n12535), .B(n12536), .Z(n486) );
  NAND U1016 ( .A(n485), .B(n486), .Z(n12683) );
  NAND U1017 ( .A(n13116), .B(n13115), .Z(n487) );
  NAND U1018 ( .A(n13113), .B(n13114), .Z(n488) );
  NAND U1019 ( .A(n487), .B(n488), .Z(n13264) );
  NAND U1020 ( .A(n15607), .B(n15606), .Z(n489) );
  NAND U1021 ( .A(n15604), .B(n15605), .Z(n490) );
  NAND U1022 ( .A(n489), .B(n490), .Z(n15752) );
  NAND U1023 ( .A(n16920), .B(n16919), .Z(n491) );
  NAND U1024 ( .A(n16917), .B(n16918), .Z(n492) );
  NAND U1025 ( .A(n491), .B(n492), .Z(n17064) );
  NAND U1026 ( .A(n17928), .B(n17927), .Z(n493) );
  NAND U1027 ( .A(n17925), .B(n17926), .Z(n494) );
  NAND U1028 ( .A(n493), .B(n494), .Z(n18073) );
  NAND U1029 ( .A(n19800), .B(n19799), .Z(n495) );
  NAND U1030 ( .A(n19797), .B(n19798), .Z(n496) );
  NAND U1031 ( .A(n495), .B(n496), .Z(n19940) );
  NAND U1032 ( .A(n23567), .B(n23566), .Z(n497) );
  NAND U1033 ( .A(n23564), .B(n23565), .Z(n498) );
  NAND U1034 ( .A(n497), .B(n498), .Z(n23711) );
  NAND U1035 ( .A(n25908), .B(n25907), .Z(n499) );
  NAND U1036 ( .A(n25905), .B(n25906), .Z(n500) );
  NAND U1037 ( .A(n499), .B(n500), .Z(n26053) );
  NAND U1038 ( .A(n26629), .B(n26628), .Z(n501) );
  NAND U1039 ( .A(n26626), .B(n26627), .Z(n502) );
  NAND U1040 ( .A(n501), .B(n502), .Z(n26768) );
  NAND U1041 ( .A(n30401), .B(n30400), .Z(n503) );
  NAND U1042 ( .A(n30398), .B(n30399), .Z(n504) );
  NAND U1043 ( .A(n503), .B(n504), .Z(n30540) );
  NAND U1044 ( .A(n31121), .B(n31120), .Z(n505) );
  NAND U1045 ( .A(n31118), .B(n31119), .Z(n506) );
  NAND U1046 ( .A(n505), .B(n506), .Z(n31266) );
  NAND U1047 ( .A(n31704), .B(n31703), .Z(n507) );
  NAND U1048 ( .A(n31701), .B(n31702), .Z(n508) );
  NAND U1049 ( .A(n507), .B(n508), .Z(n31849) );
  NAND U1050 ( .A(n33015), .B(n33014), .Z(n509) );
  NAND U1051 ( .A(n33012), .B(n33013), .Z(n510) );
  NAND U1052 ( .A(n509), .B(n510), .Z(n33161) );
  NAND U1053 ( .A(n33743), .B(n33742), .Z(n511) );
  NAND U1054 ( .A(n33740), .B(n33741), .Z(n512) );
  NAND U1055 ( .A(n511), .B(n512), .Z(n33880) );
  NAND U1056 ( .A(n37631), .B(n37630), .Z(n513) );
  NANDN U1057 ( .A(n37629), .B(n37628), .Z(n514) );
  NAND U1058 ( .A(n513), .B(n514), .Z(n37636) );
  NAND U1059 ( .A(n37870), .B(n37869), .Z(n515) );
  NANDN U1060 ( .A(n37868), .B(n37867), .Z(n516) );
  AND U1061 ( .A(n515), .B(n516), .Z(n37957) );
  NAND U1062 ( .A(n38391), .B(n38390), .Z(n517) );
  NANDN U1063 ( .A(n38389), .B(n38388), .Z(n518) );
  NAND U1064 ( .A(n517), .B(n518), .Z(n38395) );
  XNOR U1065 ( .A(n38560), .B(n38559), .Z(n38546) );
  XOR U1066 ( .A(n1106), .B(n1105), .Z(n519) );
  NAND U1067 ( .A(n519), .B(n1104), .Z(n520) );
  NAND U1068 ( .A(n1106), .B(n1105), .Z(n521) );
  AND U1069 ( .A(n520), .B(n521), .Z(n1110) );
  NAND U1070 ( .A(n1506), .B(n1505), .Z(n522) );
  NAND U1071 ( .A(n1503), .B(n1504), .Z(n523) );
  NAND U1072 ( .A(n522), .B(n523), .Z(n1563) );
  NAND U1073 ( .A(n37006), .B(n37005), .Z(n524) );
  XOR U1074 ( .A(n37005), .B(n37006), .Z(n525) );
  NANDN U1075 ( .A(n37007), .B(n525), .Z(n526) );
  NAND U1076 ( .A(n524), .B(n526), .Z(n37131) );
  NANDN U1077 ( .A(n37232), .B(n37231), .Z(n527) );
  NANDN U1078 ( .A(n37234), .B(n37233), .Z(n528) );
  NAND U1079 ( .A(n527), .B(n528), .Z(n37237) );
  XOR U1080 ( .A(n37547), .B(n37545), .Z(n529) );
  NANDN U1081 ( .A(n37546), .B(n529), .Z(n530) );
  NAND U1082 ( .A(n37547), .B(n37545), .Z(n531) );
  AND U1083 ( .A(n530), .B(n531), .Z(n37718) );
  NAND U1084 ( .A(n37805), .B(n37804), .Z(n532) );
  XOR U1085 ( .A(n37804), .B(n37805), .Z(n533) );
  NANDN U1086 ( .A(n37806), .B(n533), .Z(n534) );
  NAND U1087 ( .A(n532), .B(n534), .Z(n37890) );
  NAND U1088 ( .A(n38116), .B(n38114), .Z(n535) );
  XOR U1089 ( .A(n38114), .B(n38116), .Z(n536) );
  NANDN U1090 ( .A(n38115), .B(n536), .Z(n537) );
  NAND U1091 ( .A(n535), .B(n537), .Z(n38183) );
  NAND U1092 ( .A(n38307), .B(n38306), .Z(n538) );
  NANDN U1093 ( .A(n38305), .B(n38304), .Z(n539) );
  NAND U1094 ( .A(n538), .B(n539), .Z(n38347) );
  NAND U1095 ( .A(n38480), .B(n38479), .Z(n540) );
  XOR U1096 ( .A(n38479), .B(n38480), .Z(n541) );
  NAND U1097 ( .A(n541), .B(n38478), .Z(n542) );
  NAND U1098 ( .A(n540), .B(n542), .Z(n38512) );
  NANDN U1099 ( .A(n3393), .B(b[29]), .Z(n543) );
  ANDN U1100 ( .B(n543), .A(n1059), .Z(n544) );
  XNOR U1101 ( .A(b[29]), .B(n3393), .Z(n545) );
  NAND U1102 ( .A(n545), .B(b[30]), .Z(n546) );
  NAND U1103 ( .A(n544), .B(n546), .Z(n3376) );
  XNOR U1104 ( .A(n3969), .B(n3970), .Z(n3972) );
  XOR U1105 ( .A(n4393), .B(n4394), .Z(n4395) );
  XNOR U1106 ( .A(n4954), .B(n4953), .Z(n4955) );
  XNOR U1107 ( .A(n5096), .B(n5097), .Z(n5099) );
  XNOR U1108 ( .A(n5249), .B(n5250), .Z(n5252) );
  XOR U1109 ( .A(n5501), .B(n5502), .Z(n5503) );
  XNOR U1110 ( .A(n5496), .B(n5495), .Z(n5497) );
  XOR U1111 ( .A(n5648), .B(n5649), .Z(n5650) );
  XNOR U1112 ( .A(n5643), .B(n5642), .Z(n5644) );
  XOR U1113 ( .A(n5795), .B(n5796), .Z(n5797) );
  XNOR U1114 ( .A(n5790), .B(n5789), .Z(n5791) );
  XOR U1115 ( .A(n6099), .B(n6100), .Z(n6101) );
  XNOR U1116 ( .A(n6094), .B(n6093), .Z(n6095) );
  XNOR U1117 ( .A(n6421), .B(n6422), .Z(n6424) );
  XNOR U1118 ( .A(n6695), .B(n6696), .Z(n6698) );
  XNOR U1119 ( .A(n6689), .B(n6690), .Z(n6692) );
  XOR U1120 ( .A(n6683), .B(n6684), .Z(n6685) );
  XNOR U1121 ( .A(n6678), .B(n6677), .Z(n6679) );
  XNOR U1122 ( .A(n6850), .B(n6851), .Z(n6853) );
  XNOR U1123 ( .A(n7127), .B(n7128), .Z(n7130) );
  XNOR U1124 ( .A(n7121), .B(n7122), .Z(n7124) );
  XNOR U1125 ( .A(n7287), .B(n7288), .Z(n7290) );
  XNOR U1126 ( .A(n7281), .B(n7282), .Z(n7284) );
  XOR U1127 ( .A(n7275), .B(n7276), .Z(n7277) );
  XOR U1128 ( .A(n7269), .B(n7270), .Z(n7271) );
  XNOR U1129 ( .A(n7453), .B(n7454), .Z(n7456) );
  XOR U1130 ( .A(n7719), .B(n7720), .Z(n7721) );
  XNOR U1131 ( .A(n7714), .B(n7713), .Z(n7715) );
  XNOR U1132 ( .A(n7904), .B(n7905), .Z(n7907) );
  XOR U1133 ( .A(n8016), .B(n8017), .Z(n8018) );
  XOR U1134 ( .A(n8010), .B(n8011), .Z(n8012) );
  XNOR U1135 ( .A(n8340), .B(n8341), .Z(n8343) );
  XNOR U1136 ( .A(n8483), .B(n8484), .Z(n8486) );
  XNOR U1137 ( .A(n8630), .B(n8631), .Z(n8633) );
  XNOR U1138 ( .A(n8907), .B(n8908), .Z(n8910) );
  XNOR U1139 ( .A(n8901), .B(n8902), .Z(n8904) );
  XOR U1140 ( .A(n8895), .B(n8896), .Z(n8897) );
  XOR U1141 ( .A(n8889), .B(n8890), .Z(n8891) );
  XNOR U1142 ( .A(n9062), .B(n9063), .Z(n9065) );
  XOR U1143 ( .A(n9338), .B(n9339), .Z(n9340) );
  XNOR U1144 ( .A(n9333), .B(n9332), .Z(n9334) );
  XNOR U1145 ( .A(n9511), .B(n9512), .Z(n9514) );
  XNOR U1146 ( .A(n9646), .B(n9647), .Z(n9649) );
  XNOR U1147 ( .A(n9640), .B(n9641), .Z(n9643) );
  XOR U1148 ( .A(n9634), .B(n9635), .Z(n9636) );
  XNOR U1149 ( .A(n9629), .B(n9628), .Z(n9630) );
  XOR U1150 ( .A(n9931), .B(n9932), .Z(n9933) );
  XOR U1151 ( .A(n9925), .B(n9926), .Z(n9927) );
  XNOR U1152 ( .A(n10244), .B(n10243), .Z(n10245) );
  XOR U1153 ( .A(n10529), .B(n10530), .Z(n10531) );
  XNOR U1154 ( .A(n10535), .B(n10536), .Z(n10538) );
  XNOR U1155 ( .A(n10810), .B(n10811), .Z(n10813) );
  XNOR U1156 ( .A(n10804), .B(n10805), .Z(n10807) );
  XOR U1157 ( .A(n10798), .B(n10799), .Z(n10800) );
  XOR U1158 ( .A(n10792), .B(n10793), .Z(n10794) );
  XNOR U1159 ( .A(n10963), .B(n10964), .Z(n10966) );
  XOR U1160 ( .A(n11229), .B(n11230), .Z(n11231) );
  XNOR U1161 ( .A(n11224), .B(n11223), .Z(n11225) );
  XOR U1162 ( .A(n11377), .B(n11378), .Z(n11379) );
  XOR U1163 ( .A(n11371), .B(n11372), .Z(n11373) );
  XNOR U1164 ( .A(n11824), .B(n11825), .Z(n11827) );
  XNOR U1165 ( .A(n11818), .B(n11819), .Z(n11821) );
  XOR U1166 ( .A(n11812), .B(n11813), .Z(n11814) );
  XNOR U1167 ( .A(n11807), .B(n11806), .Z(n11808) );
  XNOR U1168 ( .A(n12119), .B(n12120), .Z(n12122) );
  XNOR U1169 ( .A(n12113), .B(n12114), .Z(n12116) );
  XOR U1170 ( .A(n12107), .B(n12108), .Z(n12109) );
  XOR U1171 ( .A(n12101), .B(n12102), .Z(n12103) );
  XOR U1172 ( .A(n12403), .B(n12404), .Z(n12405) );
  XNOR U1173 ( .A(n12398), .B(n12397), .Z(n12399) );
  XOR U1174 ( .A(n12569), .B(n12570), .Z(n12571) );
  XNOR U1175 ( .A(n12994), .B(n12995), .Z(n12997) );
  XNOR U1176 ( .A(n12988), .B(n12989), .Z(n12991) );
  XOR U1177 ( .A(n12982), .B(n12983), .Z(n12984) );
  XNOR U1178 ( .A(n12977), .B(n12976), .Z(n12978) );
  XNOR U1179 ( .A(n13291), .B(n13292), .Z(n13294) );
  XNOR U1180 ( .A(n13285), .B(n13286), .Z(n13288) );
  XOR U1181 ( .A(n13279), .B(n13280), .Z(n13281) );
  XOR U1182 ( .A(n13273), .B(n13274), .Z(n13275) );
  XNOR U1183 ( .A(n13468), .B(n13469), .Z(n13471) );
  XNOR U1184 ( .A(n13734), .B(n13735), .Z(n13737) );
  XNOR U1185 ( .A(n13728), .B(n13729), .Z(n13731) );
  XOR U1186 ( .A(n13722), .B(n13723), .Z(n13724) );
  XNOR U1187 ( .A(n13717), .B(n13716), .Z(n13718) );
  XNOR U1188 ( .A(n13899), .B(n13900), .Z(n13902) );
  XNOR U1189 ( .A(n14354), .B(n14355), .Z(n14357) );
  XNOR U1190 ( .A(n14475), .B(n14476), .Z(n14478) );
  XNOR U1191 ( .A(n14469), .B(n14470), .Z(n14472) );
  XOR U1192 ( .A(n14463), .B(n14464), .Z(n14465) );
  XNOR U1193 ( .A(n14458), .B(n14457), .Z(n14459) );
  XNOR U1194 ( .A(n14921), .B(n14920), .Z(n14922) );
  XNOR U1195 ( .A(n15126), .B(n15127), .Z(n15129) );
  XNOR U1196 ( .A(n15199), .B(n15200), .Z(n15202) );
  XNOR U1197 ( .A(n15193), .B(n15194), .Z(n15196) );
  XOR U1198 ( .A(n15187), .B(n15188), .Z(n15189) );
  XOR U1199 ( .A(n15181), .B(n15182), .Z(n15183) );
  XNOR U1200 ( .A(n15484), .B(n15485), .Z(n15487) );
  XNOR U1201 ( .A(n15478), .B(n15479), .Z(n15481) );
  XNOR U1202 ( .A(n15632), .B(n15633), .Z(n15635) );
  XNOR U1203 ( .A(n15626), .B(n15627), .Z(n15629) );
  XOR U1204 ( .A(n15620), .B(n15621), .Z(n15622) );
  XOR U1205 ( .A(n15614), .B(n15615), .Z(n15616) );
  XOR U1206 ( .A(n15926), .B(n15927), .Z(n15928) );
  XNOR U1207 ( .A(n15921), .B(n15920), .Z(n15922) );
  XNOR U1208 ( .A(n16232), .B(n16233), .Z(n16235) );
  XNOR U1209 ( .A(n16226), .B(n16227), .Z(n16229) );
  XOR U1210 ( .A(n16220), .B(n16221), .Z(n16222) );
  XNOR U1211 ( .A(n16215), .B(n16214), .Z(n16216) );
  XNOR U1212 ( .A(n16678), .B(n16677), .Z(n16679) );
  XNOR U1213 ( .A(n16820), .B(n16821), .Z(n16823) );
  XOR U1214 ( .A(n17075), .B(n17076), .Z(n17124) );
  XNOR U1215 ( .A(n17268), .B(n17269), .Z(n17271) );
  XNOR U1216 ( .A(n17391), .B(n17392), .Z(n17394) );
  XNOR U1217 ( .A(n17385), .B(n17386), .Z(n17388) );
  XNOR U1218 ( .A(n17535), .B(n17534), .Z(n17536) );
  XNOR U1219 ( .A(n17736), .B(n17735), .Z(n17737) );
  XNOR U1220 ( .A(n17953), .B(n17954), .Z(n17956) );
  XNOR U1221 ( .A(n17947), .B(n17948), .Z(n17950) );
  XOR U1222 ( .A(n18098), .B(n18099), .Z(n18100) );
  XNOR U1223 ( .A(n18093), .B(n18092), .Z(n18094) );
  XNOR U1224 ( .A(n18409), .B(n18408), .Z(n18410) );
  XNOR U1225 ( .A(n18830), .B(n18829), .Z(n18831) );
  XNOR U1226 ( .A(n19035), .B(n19036), .Z(n19038) );
  XNOR U1227 ( .A(n19108), .B(n19109), .Z(n19111) );
  XNOR U1228 ( .A(n19102), .B(n19103), .Z(n19105) );
  XOR U1229 ( .A(n19096), .B(n19097), .Z(n19098) );
  XOR U1230 ( .A(n19090), .B(n19091), .Z(n19092) );
  XOR U1231 ( .A(n19380), .B(n19381), .Z(n19382) );
  XNOR U1232 ( .A(n19375), .B(n19374), .Z(n19376) );
  XNOR U1233 ( .A(n19546), .B(n19545), .Z(n19547) );
  XOR U1234 ( .A(n19955), .B(n19956), .Z(n19957) );
  XOR U1235 ( .A(n19949), .B(n19950), .Z(n19951) );
  XNOR U1236 ( .A(n20290), .B(n20291), .Z(n20293) );
  XNOR U1237 ( .A(n20435), .B(n20436), .Z(n20438) );
  XNOR U1238 ( .A(n20872), .B(n20873), .Z(n20875) );
  XNOR U1239 ( .A(n21017), .B(n21018), .Z(n21020) );
  XNOR U1240 ( .A(n21454), .B(n21455), .Z(n21457) );
  XNOR U1241 ( .A(n21878), .B(n21877), .Z(n21879) );
  XNOR U1242 ( .A(n22020), .B(n22021), .Z(n22023) );
  XNOR U1243 ( .A(n22303), .B(n22304), .Z(n22306) );
  XNOR U1244 ( .A(n22297), .B(n22298), .Z(n22300) );
  XOR U1245 ( .A(n22428), .B(n22429), .Z(n22430) );
  XNOR U1246 ( .A(n22423), .B(n22422), .Z(n22424) );
  XNOR U1247 ( .A(n22598), .B(n22599), .Z(n22601) );
  XNOR U1248 ( .A(n22592), .B(n22593), .Z(n22595) );
  XOR U1249 ( .A(n22586), .B(n22587), .Z(n22588) );
  XOR U1250 ( .A(n22580), .B(n22581), .Z(n22582) );
  XNOR U1251 ( .A(n23046), .B(n23045), .Z(n23047) );
  XNOR U1252 ( .A(n23328), .B(n23327), .Z(n23329) );
  XOR U1253 ( .A(n23513), .B(n23514), .Z(n23515) );
  XNOR U1254 ( .A(n23746), .B(n23747), .Z(n23749) );
  XNOR U1255 ( .A(n23740), .B(n23741), .Z(n23743) );
  XOR U1256 ( .A(n23734), .B(n23735), .Z(n23736) );
  XOR U1257 ( .A(n23728), .B(n23729), .Z(n23730) );
  XOR U1258 ( .A(n24033), .B(n24034), .Z(n24035) );
  XOR U1259 ( .A(n24027), .B(n24028), .Z(n24029) );
  XOR U1260 ( .A(n24189), .B(n24190), .Z(n24191) );
  XNOR U1261 ( .A(n24507), .B(n24508), .Z(n24510) );
  XNOR U1262 ( .A(n24627), .B(n24628), .Z(n24630) );
  XNOR U1263 ( .A(n24621), .B(n24622), .Z(n24624) );
  XNOR U1264 ( .A(n24764), .B(n24765), .Z(n24767) );
  XNOR U1265 ( .A(n24758), .B(n24759), .Z(n24761) );
  XOR U1266 ( .A(n24752), .B(n24753), .Z(n24754) );
  XNOR U1267 ( .A(n24747), .B(n24746), .Z(n24748) );
  XNOR U1268 ( .A(n25232), .B(n25233), .Z(n25235) );
  XOR U1269 ( .A(n25495), .B(n25496), .Z(n25497) );
  XOR U1270 ( .A(n25489), .B(n25490), .Z(n25491) );
  XNOR U1271 ( .A(n25663), .B(n25662), .Z(n25664) );
  XNOR U1272 ( .A(n25943), .B(n25944), .Z(n25946) );
  XNOR U1273 ( .A(n25937), .B(n25938), .Z(n25940) );
  XOR U1274 ( .A(n26068), .B(n26069), .Z(n26070) );
  XNOR U1275 ( .A(n26063), .B(n26062), .Z(n26064) );
  XNOR U1276 ( .A(n26389), .B(n26388), .Z(n26390) );
  XNOR U1277 ( .A(n26672), .B(n26673), .Z(n26675) );
  XNOR U1278 ( .A(n26951), .B(n26952), .Z(n26954) );
  XNOR U1279 ( .A(n26945), .B(n26946), .Z(n26948) );
  XOR U1280 ( .A(n26939), .B(n26940), .Z(n26941) );
  XOR U1281 ( .A(n26933), .B(n26934), .Z(n26935) );
  XNOR U1282 ( .A(n27238), .B(n27239), .Z(n27241) );
  XNOR U1283 ( .A(n27232), .B(n27233), .Z(n27235) );
  XOR U1284 ( .A(n27226), .B(n27227), .Z(n27228) );
  XNOR U1285 ( .A(n27403), .B(n27404), .Z(n27406) );
  XOR U1286 ( .A(n27669), .B(n27670), .Z(n27671) );
  XNOR U1287 ( .A(n27664), .B(n27663), .Z(n27665) );
  XOR U1288 ( .A(n28118), .B(n28119), .Z(n28120) );
  XNOR U1289 ( .A(n28113), .B(n28112), .Z(n28114) );
  XNOR U1290 ( .A(n28279), .B(n28280), .Z(n28282) );
  XNOR U1291 ( .A(n28273), .B(n28274), .Z(n28276) );
  XOR U1292 ( .A(n28267), .B(n28268), .Z(n28269) );
  XNOR U1293 ( .A(n28262), .B(n28261), .Z(n28263) );
  XNOR U1294 ( .A(n28446), .B(n28447), .Z(n28449) );
  XNOR U1295 ( .A(n28937), .B(n28938), .Z(n28940) );
  XNOR U1296 ( .A(n29008), .B(n29009), .Z(n29011) );
  XNOR U1297 ( .A(n29002), .B(n29003), .Z(n29005) );
  XNOR U1298 ( .A(n29305), .B(n29304), .Z(n29306) );
  XNOR U1299 ( .A(n30161), .B(n30160), .Z(n30162) );
  XNOR U1300 ( .A(n30444), .B(n30445), .Z(n30447) );
  XOR U1301 ( .A(n30987), .B(n30988), .Z(n30989) );
  XOR U1302 ( .A(n30981), .B(n30982), .Z(n30983) );
  XNOR U1303 ( .A(n31311), .B(n31312), .Z(n31314) );
  XNOR U1304 ( .A(n31581), .B(n31582), .Z(n31584) );
  XNOR U1305 ( .A(n31575), .B(n31576), .Z(n31578) );
  XOR U1306 ( .A(n31717), .B(n31718), .Z(n31719) );
  XOR U1307 ( .A(n31711), .B(n31712), .Z(n31713) );
  XNOR U1308 ( .A(n32306), .B(n32307), .Z(n32309) );
  XNOR U1309 ( .A(n32300), .B(n32301), .Z(n32303) );
  XOR U1310 ( .A(n32294), .B(n32295), .Z(n32296) );
  XOR U1311 ( .A(n32288), .B(n32289), .Z(n32290) );
  XNOR U1312 ( .A(n32471), .B(n32472), .Z(n32474) );
  XOR U1313 ( .A(n32756), .B(n32757), .Z(n32758) );
  XNOR U1314 ( .A(n32895), .B(n32896), .Z(n32898) );
  XNOR U1315 ( .A(n32889), .B(n32890), .Z(n32892) );
  XOR U1316 ( .A(n32883), .B(n32884), .Z(n32885) );
  XNOR U1317 ( .A(n32878), .B(n32877), .Z(n32879) );
  XNOR U1318 ( .A(n33188), .B(n33189), .Z(n33191) );
  XNOR U1319 ( .A(n33182), .B(n33183), .Z(n33185) );
  XOR U1320 ( .A(n33176), .B(n33177), .Z(n33178) );
  XOR U1321 ( .A(n33170), .B(n33171), .Z(n33172) );
  XNOR U1322 ( .A(n33491), .B(n33490), .Z(n33492) );
  XNOR U1323 ( .A(n33785), .B(n33784), .Z(n33786) );
  XNOR U1324 ( .A(n33925), .B(n33926), .Z(n33928) );
  XNOR U1325 ( .A(n34078), .B(n34079), .Z(n34081) );
  XNOR U1326 ( .A(n34354), .B(n34355), .Z(n34357) );
  XNOR U1327 ( .A(n34348), .B(n34349), .Z(n34351) );
  XOR U1328 ( .A(n34342), .B(n34343), .Z(n34344) );
  XNOR U1329 ( .A(n34337), .B(n34336), .Z(n34338) );
  XOR U1330 ( .A(n34636), .B(n34637), .Z(n34686) );
  XOR U1331 ( .A(n35065), .B(n35066), .Z(n35067) );
  XNOR U1332 ( .A(n35060), .B(n35059), .Z(n35061) );
  NAND U1333 ( .A(a[255]), .B(n1049), .Z(n547) );
  AND U1334 ( .A(b[1]), .B(n547), .Z(n36122) );
  ANDN U1335 ( .B(n3393), .A(n1057), .Z(n548) );
  ANDN U1336 ( .B(n548), .A(n38268), .Z(n549) );
  NOR U1337 ( .A(n1057), .B(b[22]), .Z(n550) );
  NAND U1338 ( .A(n550), .B(n1056), .Z(n551) );
  NANDN U1339 ( .A(n549), .B(n551), .Z(n2402) );
  NAND U1340 ( .A(n3192), .B(n3193), .Z(n552) );
  NANDN U1341 ( .A(n3191), .B(n3190), .Z(n553) );
  NAND U1342 ( .A(n552), .B(n553), .Z(n3223) );
  NAND U1343 ( .A(n3268), .B(n3267), .Z(n554) );
  NANDN U1344 ( .A(n3266), .B(n3265), .Z(n555) );
  NAND U1345 ( .A(n554), .B(n555), .Z(n3363) );
  NAND U1346 ( .A(n3611), .B(n3610), .Z(n556) );
  NANDN U1347 ( .A(n3609), .B(n3608), .Z(n557) );
  AND U1348 ( .A(n556), .B(n557), .Z(n3764) );
  NAND U1349 ( .A(n3534), .B(n3533), .Z(n558) );
  NANDN U1350 ( .A(n3532), .B(n3531), .Z(n559) );
  NAND U1351 ( .A(n558), .B(n559), .Z(n3757) );
  XOR U1352 ( .A(n4259), .B(n4260), .Z(n4261) );
  NAND U1353 ( .A(n4141), .B(n4140), .Z(n560) );
  NANDN U1354 ( .A(n4139), .B(n4138), .Z(n561) );
  NAND U1355 ( .A(n560), .B(n561), .Z(n4325) );
  NAND U1356 ( .A(n4274), .B(n4273), .Z(n562) );
  NANDN U1357 ( .A(n4272), .B(n4271), .Z(n563) );
  NAND U1358 ( .A(n562), .B(n563), .Z(n4360) );
  NAND U1359 ( .A(n4849), .B(n4848), .Z(n564) );
  NANDN U1360 ( .A(n4847), .B(n4846), .Z(n565) );
  NAND U1361 ( .A(n564), .B(n565), .Z(n4920) );
  NAND U1362 ( .A(n5276), .B(n5275), .Z(n566) );
  NANDN U1363 ( .A(n5274), .B(n5273), .Z(n567) );
  NAND U1364 ( .A(n566), .B(n567), .Z(n5461) );
  XOR U1365 ( .A(n5543), .B(n5544), .Z(n5545) );
  NAND U1366 ( .A(n5411), .B(n5410), .Z(n568) );
  NANDN U1367 ( .A(n5409), .B(n5408), .Z(n569) );
  NAND U1368 ( .A(n568), .B(n569), .Z(n5610) );
  XNOR U1369 ( .A(n5690), .B(n5691), .Z(n5693) );
  XNOR U1370 ( .A(n5837), .B(n5838), .Z(n5840) );
  XNOR U1371 ( .A(n5982), .B(n5983), .Z(n5985) );
  XNOR U1372 ( .A(n6274), .B(n6275), .Z(n6277) );
  XOR U1373 ( .A(n6725), .B(n6726), .Z(n6727) );
  NAND U1374 ( .A(n6593), .B(n6592), .Z(n570) );
  NANDN U1375 ( .A(n6591), .B(n6590), .Z(n571) );
  NAND U1376 ( .A(n570), .B(n571), .Z(n6792) );
  XOR U1377 ( .A(n7157), .B(n7158), .Z(n7159) );
  NAND U1378 ( .A(n7038), .B(n7037), .Z(n572) );
  NANDN U1379 ( .A(n7036), .B(n7035), .Z(n573) );
  NAND U1380 ( .A(n572), .B(n573), .Z(n7225) );
  XOR U1381 ( .A(n7761), .B(n7762), .Z(n7763) );
  NAND U1382 ( .A(n7629), .B(n7628), .Z(n574) );
  NANDN U1383 ( .A(n7627), .B(n7626), .Z(n575) );
  NAND U1384 ( .A(n574), .B(n575), .Z(n7828) );
  XNOR U1385 ( .A(n7910), .B(n7911), .Z(n7913) );
  XNOR U1386 ( .A(n8205), .B(n8206), .Z(n8208) );
  NAND U1387 ( .A(n8510), .B(n8509), .Z(n576) );
  NANDN U1388 ( .A(n8508), .B(n8507), .Z(n577) );
  NAND U1389 ( .A(n576), .B(n577), .Z(n8707) );
  NAND U1390 ( .A(n8657), .B(n8656), .Z(n578) );
  NANDN U1391 ( .A(n8655), .B(n8654), .Z(n579) );
  NAND U1392 ( .A(n578), .B(n579), .Z(n8855) );
  XOR U1393 ( .A(n8937), .B(n8938), .Z(n8939) );
  NAND U1394 ( .A(n8804), .B(n8803), .Z(n580) );
  NANDN U1395 ( .A(n8802), .B(n8801), .Z(n581) );
  NAND U1396 ( .A(n580), .B(n581), .Z(n9004) );
  XOR U1397 ( .A(n9380), .B(n9381), .Z(n9382) );
  NAND U1398 ( .A(n9250), .B(n9249), .Z(n582) );
  NANDN U1399 ( .A(n9248), .B(n9247), .Z(n583) );
  NAND U1400 ( .A(n582), .B(n583), .Z(n9447) );
  XNOR U1401 ( .A(n9517), .B(n9518), .Z(n9520) );
  XOR U1402 ( .A(n9973), .B(n9974), .Z(n9975) );
  XNOR U1403 ( .A(n10120), .B(n10121), .Z(n10123) );
  XOR U1404 ( .A(n10541), .B(n10542), .Z(n10543) );
  NAND U1405 ( .A(n10556), .B(n10555), .Z(n584) );
  NANDN U1406 ( .A(n10554), .B(n10553), .Z(n585) );
  NAND U1407 ( .A(n584), .B(n585), .Z(n10748) );
  XOR U1408 ( .A(n11271), .B(n11272), .Z(n11273) );
  NAND U1409 ( .A(n11151), .B(n11150), .Z(n586) );
  NANDN U1410 ( .A(n11149), .B(n11148), .Z(n587) );
  NAND U1411 ( .A(n586), .B(n587), .Z(n11339) );
  XNOR U1412 ( .A(n11419), .B(n11420), .Z(n11422) );
  XNOR U1413 ( .A(n11564), .B(n11565), .Z(n11567) );
  XOR U1414 ( .A(n11854), .B(n11855), .Z(n11856) );
  XOR U1415 ( .A(n12149), .B(n12150), .Z(n12151) );
  XOR U1416 ( .A(n12445), .B(n12446), .Z(n12447) );
  XNOR U1417 ( .A(n12591), .B(n12592), .Z(n12594) );
  XOR U1418 ( .A(n13024), .B(n13025), .Z(n13026) );
  NAND U1419 ( .A(n12906), .B(n12905), .Z(n588) );
  NANDN U1420 ( .A(n12904), .B(n12903), .Z(n589) );
  NAND U1421 ( .A(n588), .B(n589), .Z(n13091) );
  XOR U1422 ( .A(n13321), .B(n13322), .Z(n13323) );
  XOR U1423 ( .A(n13764), .B(n13765), .Z(n13766) );
  NAND U1424 ( .A(n13632), .B(n13631), .Z(n590) );
  NANDN U1425 ( .A(n13630), .B(n13629), .Z(n591) );
  NAND U1426 ( .A(n590), .B(n591), .Z(n13831) );
  XOR U1427 ( .A(n14203), .B(n14204), .Z(n14205) );
  NAND U1428 ( .A(n14075), .B(n14074), .Z(n592) );
  NANDN U1429 ( .A(n14073), .B(n14072), .Z(n593) );
  NAND U1430 ( .A(n592), .B(n593), .Z(n14268) );
  NAND U1431 ( .A(n14218), .B(n14217), .Z(n594) );
  NANDN U1432 ( .A(n14216), .B(n14215), .Z(n595) );
  NAND U1433 ( .A(n594), .B(n595), .Z(n14303) );
  XOR U1434 ( .A(n14799), .B(n14800), .Z(n14801) );
  NAND U1435 ( .A(n14814), .B(n14813), .Z(n596) );
  NANDN U1436 ( .A(n14812), .B(n14811), .Z(n597) );
  NAND U1437 ( .A(n596), .B(n597), .Z(n14887) );
  XOR U1438 ( .A(n15514), .B(n15515), .Z(n15516) );
  XOR U1439 ( .A(n15968), .B(n15969), .Z(n15970) );
  XNOR U1440 ( .A(n16103), .B(n16104), .Z(n16106) );
  XOR U1441 ( .A(n16556), .B(n16557), .Z(n16558) );
  NAND U1442 ( .A(n16571), .B(n16570), .Z(n598) );
  NANDN U1443 ( .A(n16569), .B(n16568), .Z(n599) );
  NAND U1444 ( .A(n598), .B(n599), .Z(n16644) );
  NAND U1445 ( .A(n16845), .B(n16844), .Z(n600) );
  NANDN U1446 ( .A(n16843), .B(n16842), .Z(n601) );
  NAND U1447 ( .A(n600), .B(n601), .Z(n17050) );
  XOR U1448 ( .A(n17115), .B(n17116), .Z(n17117) );
  NAND U1449 ( .A(n17000), .B(n16999), .Z(n602) );
  NANDN U1450 ( .A(n16998), .B(n16997), .Z(n603) );
  NAND U1451 ( .A(n602), .B(n603), .Z(n17182) );
  NAND U1452 ( .A(n17668), .B(n17667), .Z(n604) );
  NANDN U1453 ( .A(n17666), .B(n17665), .Z(n605) );
  NAND U1454 ( .A(n604), .B(n605), .Z(n17900) );
  XOR U1455 ( .A(n17983), .B(n17984), .Z(n17985) );
  NAND U1456 ( .A(n17856), .B(n17855), .Z(n606) );
  NANDN U1457 ( .A(n17854), .B(n17853), .Z(n607) );
  NAND U1458 ( .A(n606), .B(n607), .Z(n18050) );
  XNOR U1459 ( .A(n18273), .B(n18274), .Z(n18276) );
  NAND U1460 ( .A(n18725), .B(n18724), .Z(n608) );
  NANDN U1461 ( .A(n18723), .B(n18722), .Z(n609) );
  NAND U1462 ( .A(n608), .B(n609), .Z(n18796) );
  XOR U1463 ( .A(n19422), .B(n19423), .Z(n19424) );
  XNOR U1464 ( .A(n19567), .B(n19568), .Z(n19570) );
  NAND U1465 ( .A(n19727), .B(n19726), .Z(n610) );
  NANDN U1466 ( .A(n19725), .B(n19724), .Z(n611) );
  NAND U1467 ( .A(n610), .B(n611), .Z(n19807) );
  XOR U1468 ( .A(n20051), .B(n20052), .Z(n20053) );
  XNOR U1469 ( .A(n20154), .B(n20155), .Z(n20157) );
  NAND U1470 ( .A(n20462), .B(n20461), .Z(n612) );
  NANDN U1471 ( .A(n20460), .B(n20459), .Z(n613) );
  NAND U1472 ( .A(n612), .B(n613), .Z(n20659) );
  XOR U1473 ( .A(n20727), .B(n20728), .Z(n20729) );
  NAND U1474 ( .A(n20609), .B(n20608), .Z(n614) );
  NANDN U1475 ( .A(n20607), .B(n20606), .Z(n615) );
  NAND U1476 ( .A(n614), .B(n615), .Z(n20792) );
  NAND U1477 ( .A(n20742), .B(n20741), .Z(n616) );
  NANDN U1478 ( .A(n20740), .B(n20739), .Z(n617) );
  NAND U1479 ( .A(n616), .B(n617), .Z(n20827) );
  NAND U1480 ( .A(n21044), .B(n21043), .Z(n618) );
  NANDN U1481 ( .A(n21042), .B(n21041), .Z(n619) );
  NAND U1482 ( .A(n618), .B(n619), .Z(n21229) );
  XOR U1483 ( .A(n21309), .B(n21310), .Z(n21311) );
  NAND U1484 ( .A(n21179), .B(n21178), .Z(n620) );
  NANDN U1485 ( .A(n21177), .B(n21176), .Z(n621) );
  NAND U1486 ( .A(n620), .B(n621), .Z(n21374) );
  NAND U1487 ( .A(n21324), .B(n21323), .Z(n622) );
  NANDN U1488 ( .A(n21322), .B(n21321), .Z(n623) );
  NAND U1489 ( .A(n622), .B(n623), .Z(n21409) );
  XOR U1490 ( .A(n21744), .B(n21745), .Z(n21746) );
  NAND U1491 ( .A(n21626), .B(n21625), .Z(n624) );
  NANDN U1492 ( .A(n21624), .B(n21623), .Z(n625) );
  NAND U1493 ( .A(n624), .B(n625), .Z(n21809) );
  NAND U1494 ( .A(n21759), .B(n21758), .Z(n626) );
  NANDN U1495 ( .A(n21757), .B(n21756), .Z(n627) );
  NAND U1496 ( .A(n626), .B(n627), .Z(n21844) );
  XOR U1497 ( .A(n22333), .B(n22334), .Z(n22335) );
  NAND U1498 ( .A(n22190), .B(n22189), .Z(n628) );
  NANDN U1499 ( .A(n22188), .B(n22187), .Z(n629) );
  NAND U1500 ( .A(n628), .B(n629), .Z(n22400) );
  XNOR U1501 ( .A(n22628), .B(n22629), .Z(n22631) );
  XOR U1502 ( .A(n22924), .B(n22925), .Z(n22926) );
  NAND U1503 ( .A(n22939), .B(n22938), .Z(n630) );
  NANDN U1504 ( .A(n22937), .B(n22936), .Z(n631) );
  NAND U1505 ( .A(n630), .B(n631), .Z(n23012) );
  NAND U1506 ( .A(n23362), .B(n23361), .Z(n632) );
  NANDN U1507 ( .A(n23360), .B(n23359), .Z(n633) );
  NAND U1508 ( .A(n632), .B(n633), .Z(n23536) );
  NAND U1509 ( .A(n23446), .B(n23445), .Z(n634) );
  NANDN U1510 ( .A(n23444), .B(n23443), .Z(n635) );
  NAND U1511 ( .A(n634), .B(n635), .Z(n23681) );
  XOR U1512 ( .A(n23776), .B(n23777), .Z(n23778) );
  XOR U1513 ( .A(n24075), .B(n24076), .Z(n24077) );
  XNOR U1514 ( .A(n24211), .B(n24212), .Z(n24214) );
  NAND U1515 ( .A(n24526), .B(n24525), .Z(n636) );
  NANDN U1516 ( .A(n24524), .B(n24523), .Z(n637) );
  NAND U1517 ( .A(n636), .B(n637), .Z(n24604) );
  XOR U1518 ( .A(n25086), .B(n25087), .Z(n25088) );
  NAND U1519 ( .A(n25101), .B(n25100), .Z(n638) );
  NANDN U1520 ( .A(n25099), .B(n25098), .Z(n639) );
  NAND U1521 ( .A(n638), .B(n639), .Z(n25186) );
  XOR U1522 ( .A(n25537), .B(n25538), .Z(n25539) );
  NAND U1523 ( .A(n25404), .B(n25403), .Z(n640) );
  NANDN U1524 ( .A(n25402), .B(n25401), .Z(n641) );
  NAND U1525 ( .A(n640), .B(n641), .Z(n25604) );
  XNOR U1526 ( .A(n25684), .B(n25685), .Z(n25687) );
  XOR U1527 ( .A(n25973), .B(n25974), .Z(n25975) );
  NAND U1528 ( .A(n25834), .B(n25833), .Z(n642) );
  NANDN U1529 ( .A(n25832), .B(n25831), .Z(n643) );
  NAND U1530 ( .A(n642), .B(n643), .Z(n26040) );
  XNOR U1531 ( .A(n26265), .B(n26266), .Z(n26268) );
  NAND U1532 ( .A(n26508), .B(n26507), .Z(n644) );
  NANDN U1533 ( .A(n26506), .B(n26505), .Z(n645) );
  NAND U1534 ( .A(n644), .B(n645), .Z(n26740) );
  XOR U1535 ( .A(n26981), .B(n26982), .Z(n26983) );
  NAND U1536 ( .A(n26838), .B(n26837), .Z(n646) );
  NANDN U1537 ( .A(n26836), .B(n26835), .Z(n647) );
  NAND U1538 ( .A(n646), .B(n647), .Z(n27048) );
  XOR U1539 ( .A(n27268), .B(n27269), .Z(n27270) );
  XOR U1540 ( .A(n27711), .B(n27712), .Z(n27713) );
  NAND U1541 ( .A(n27591), .B(n27590), .Z(n648) );
  NANDN U1542 ( .A(n27589), .B(n27588), .Z(n649) );
  NAND U1543 ( .A(n648), .B(n649), .Z(n27777) );
  XNOR U1544 ( .A(n27856), .B(n27857), .Z(n27859) );
  XOR U1545 ( .A(n28160), .B(n28161), .Z(n28162) );
  XNOR U1546 ( .A(n28309), .B(n28310), .Z(n28312) );
  XOR U1547 ( .A(n28752), .B(n28753), .Z(n28754) );
  NAND U1548 ( .A(n28610), .B(n28609), .Z(n650) );
  NANDN U1549 ( .A(n28608), .B(n28607), .Z(n651) );
  NAND U1550 ( .A(n650), .B(n651), .Z(n28817) );
  NAND U1551 ( .A(n28767), .B(n28766), .Z(n652) );
  NANDN U1552 ( .A(n28765), .B(n28764), .Z(n653) );
  NAND U1553 ( .A(n652), .B(n653), .Z(n28944) );
  XOR U1554 ( .A(n29751), .B(n29752), .Z(n29753) );
  NAND U1555 ( .A(n29623), .B(n29622), .Z(n654) );
  NANDN U1556 ( .A(n29621), .B(n29620), .Z(n655) );
  NAND U1557 ( .A(n654), .B(n655), .Z(n29816) );
  NAND U1558 ( .A(n29766), .B(n29765), .Z(n656) );
  NANDN U1559 ( .A(n29764), .B(n29763), .Z(n657) );
  NAND U1560 ( .A(n656), .B(n657), .Z(n29839) );
  XOR U1561 ( .A(n30027), .B(n30028), .Z(n30029) );
  NAND U1562 ( .A(n30042), .B(n30041), .Z(n658) );
  NANDN U1563 ( .A(n30040), .B(n30039), .Z(n659) );
  NAND U1564 ( .A(n658), .B(n659), .Z(n30127) );
  NAND U1565 ( .A(n30280), .B(n30279), .Z(n660) );
  NANDN U1566 ( .A(n30278), .B(n30277), .Z(n661) );
  NAND U1567 ( .A(n660), .B(n661), .Z(n30512) );
  XOR U1568 ( .A(n30750), .B(n30751), .Z(n30752) );
  NAND U1569 ( .A(n30620), .B(n30619), .Z(n662) );
  NANDN U1570 ( .A(n30618), .B(n30617), .Z(n663) );
  NAND U1571 ( .A(n662), .B(n663), .Z(n30815) );
  NAND U1572 ( .A(n30765), .B(n30764), .Z(n664) );
  NANDN U1573 ( .A(n30763), .B(n30762), .Z(n665) );
  NAND U1574 ( .A(n664), .B(n665), .Z(n30838) );
  XOR U1575 ( .A(n31029), .B(n31030), .Z(n31031) );
  XNOR U1576 ( .A(n31186), .B(n31187), .Z(n31189) );
  XOR U1577 ( .A(n31611), .B(n31612), .Z(n31613) );
  NAND U1578 ( .A(n31480), .B(n31479), .Z(n666) );
  NANDN U1579 ( .A(n31478), .B(n31477), .Z(n667) );
  NAND U1580 ( .A(n666), .B(n667), .Z(n31679) );
  XNOR U1581 ( .A(n31914), .B(n31915), .Z(n31917) );
  XOR U1582 ( .A(n32336), .B(n32337), .Z(n32338) );
  XOR U1583 ( .A(n32778), .B(n32779), .Z(n32780) );
  NAND U1584 ( .A(n32659), .B(n32658), .Z(n668) );
  NANDN U1585 ( .A(n32657), .B(n32656), .Z(n669) );
  NAND U1586 ( .A(n668), .B(n669), .Z(n32843) );
  NAND U1587 ( .A(n32793), .B(n32792), .Z(n670) );
  NANDN U1588 ( .A(n32791), .B(n32790), .Z(n671) );
  NAND U1589 ( .A(n670), .B(n671), .Z(n32984) );
  XOR U1590 ( .A(n33218), .B(n33219), .Z(n33220) );
  XOR U1591 ( .A(n33512), .B(n33513), .Z(n33514) );
  NAND U1592 ( .A(n33527), .B(n33526), .Z(n672) );
  NANDN U1593 ( .A(n33525), .B(n33524), .Z(n673) );
  NAND U1594 ( .A(n672), .B(n673), .Z(n33714) );
  NAND U1595 ( .A(n33670), .B(n33669), .Z(n674) );
  NANDN U1596 ( .A(n33668), .B(n33667), .Z(n675) );
  NAND U1597 ( .A(n674), .B(n675), .Z(n33751) );
  NAND U1598 ( .A(n34105), .B(n34104), .Z(n676) );
  NANDN U1599 ( .A(n34103), .B(n34102), .Z(n677) );
  NAND U1600 ( .A(n676), .B(n677), .Z(n34290) );
  XOR U1601 ( .A(n34384), .B(n34385), .Z(n34386) );
  NAND U1602 ( .A(n34240), .B(n34239), .Z(n678) );
  NANDN U1603 ( .A(n34238), .B(n34237), .Z(n679) );
  NAND U1604 ( .A(n678), .B(n679), .Z(n34451) );
  XOR U1605 ( .A(n34677), .B(n34678), .Z(n34679) );
  NAND U1606 ( .A(n34809), .B(n34810), .Z(n680) );
  NANDN U1607 ( .A(n34808), .B(n34807), .Z(n681) );
  NAND U1608 ( .A(n680), .B(n681), .Z(n35027) );
  OR U1609 ( .A(n34804), .B(n34803), .Z(n682) );
  NANDN U1610 ( .A(n34806), .B(n34805), .Z(n683) );
  NAND U1611 ( .A(n682), .B(n683), .Z(n35031) );
  XOR U1612 ( .A(n35107), .B(n35108), .Z(n35109) );
  XNOR U1613 ( .A(n35264), .B(n35265), .Z(n35267) );
  OR U1614 ( .A(b[11]), .B(b[12]), .Z(n684) );
  NANDN U1615 ( .A(a[0]), .B(n37424), .Z(n685) );
  NAND U1616 ( .A(n684), .B(n685), .Z(n686) );
  NANDN U1617 ( .A(n1053), .B(n686), .Z(n1524) );
  NAND U1618 ( .A(n2135), .B(n2134), .Z(n687) );
  NANDN U1619 ( .A(n2133), .B(n2132), .Z(n688) );
  AND U1620 ( .A(n687), .B(n688), .Z(n2218) );
  NAND U1621 ( .A(n2010), .B(n2009), .Z(n689) );
  NANDN U1622 ( .A(n2008), .B(n2007), .Z(n690) );
  NAND U1623 ( .A(n689), .B(n690), .Z(n2085) );
  XNOR U1624 ( .A(n2072), .B(n2073), .Z(n2065) );
  NAND U1625 ( .A(n2548), .B(n2549), .Z(n691) );
  NANDN U1626 ( .A(n2547), .B(n2546), .Z(n692) );
  NAND U1627 ( .A(n691), .B(n692), .Z(n2678) );
  NAND U1628 ( .A(n2422), .B(n2421), .Z(n693) );
  NANDN U1629 ( .A(n2420), .B(n2419), .Z(n694) );
  AND U1630 ( .A(n693), .B(n694), .Z(n2556) );
  NAND U1631 ( .A(n2722), .B(n2721), .Z(n695) );
  NANDN U1632 ( .A(n2720), .B(n2719), .Z(n696) );
  NAND U1633 ( .A(n695), .B(n696), .Z(n2919) );
  XNOR U1634 ( .A(n3152), .B(n3153), .Z(n3157) );
  NANDN U1635 ( .A(n3593), .B(n3592), .Z(n697) );
  NANDN U1636 ( .A(n3595), .B(n3594), .Z(n698) );
  NAND U1637 ( .A(n697), .B(n698), .Z(n3640) );
  XOR U1638 ( .A(n3900), .B(n3901), .Z(n3902) );
  NAND U1639 ( .A(n3792), .B(n3793), .Z(n699) );
  NANDN U1640 ( .A(n3791), .B(n3790), .Z(n700) );
  NAND U1641 ( .A(n699), .B(n700), .Z(n4038) );
  NAND U1642 ( .A(n3932), .B(n3931), .Z(n701) );
  NAND U1643 ( .A(n3929), .B(n3930), .Z(n702) );
  AND U1644 ( .A(n701), .B(n702), .Z(n4066) );
  XNOR U1645 ( .A(n4338), .B(n4339), .Z(n4333) );
  NAND U1646 ( .A(n4365), .B(n4366), .Z(n703) );
  NANDN U1647 ( .A(n4368), .B(n4367), .Z(n704) );
  NAND U1648 ( .A(n703), .B(n704), .Z(n4617) );
  OR U1649 ( .A(n4502), .B(n4503), .Z(n705) );
  NAND U1650 ( .A(n4501), .B(n4500), .Z(n706) );
  NAND U1651 ( .A(n705), .B(n706), .Z(n4755) );
  NAND U1652 ( .A(n4754), .B(n4753), .Z(n707) );
  NANDN U1653 ( .A(n4752), .B(n4751), .Z(n708) );
  NAND U1654 ( .A(n707), .B(n708), .Z(n4897) );
  NAND U1655 ( .A(n4838), .B(n4839), .Z(n709) );
  NANDN U1656 ( .A(n4837), .B(n4836), .Z(n710) );
  NAND U1657 ( .A(n709), .B(n710), .Z(n5038) );
  NAND U1658 ( .A(n4928), .B(n4927), .Z(n711) );
  NAND U1659 ( .A(n4925), .B(n4926), .Z(n712) );
  NAND U1660 ( .A(n711), .B(n712), .Z(n5177) );
  XNOR U1661 ( .A(n5474), .B(n5475), .Z(n5469) );
  XNOR U1662 ( .A(n5623), .B(n5624), .Z(n5618) );
  NAND U1663 ( .A(n6089), .B(n6090), .Z(n713) );
  NANDN U1664 ( .A(n6092), .B(n6091), .Z(n714) );
  NAND U1665 ( .A(n713), .B(n714), .Z(n6347) );
  NAND U1666 ( .A(n6381), .B(n6382), .Z(n715) );
  NANDN U1667 ( .A(n6384), .B(n6383), .Z(n716) );
  NAND U1668 ( .A(n715), .B(n716), .Z(n6519) );
  XNOR U1669 ( .A(n6673), .B(n6674), .Z(n6668) );
  XNOR U1670 ( .A(n6971), .B(n6972), .Z(n6966) );
  XNOR U1671 ( .A(n7238), .B(n7239), .Z(n7233) );
  NAND U1672 ( .A(n7380), .B(n7379), .Z(n717) );
  NAND U1673 ( .A(n7377), .B(n7378), .Z(n718) );
  NAND U1674 ( .A(n717), .B(n718), .Z(n7405) );
  XNOR U1675 ( .A(n7562), .B(n7563), .Z(n7557) );
  XNOR U1676 ( .A(n7709), .B(n7710), .Z(n7704) );
  NANDN U1677 ( .A(n8003), .B(n8002), .Z(n719) );
  NANDN U1678 ( .A(n8001), .B(n8000), .Z(n720) );
  NAND U1679 ( .A(n719), .B(n720), .Z(n8153) );
  NAND U1680 ( .A(n8300), .B(n8301), .Z(n721) );
  NANDN U1681 ( .A(n8303), .B(n8302), .Z(n722) );
  NAND U1682 ( .A(n721), .B(n722), .Z(n8438) );
  XNOR U1683 ( .A(n8590), .B(n8591), .Z(n8585) );
  XNOR U1684 ( .A(n8737), .B(n8738), .Z(n8732) );
  XNOR U1685 ( .A(n8885), .B(n8886), .Z(n8880) );
  XNOR U1686 ( .A(n9183), .B(n9184), .Z(n9178) );
  XNOR U1687 ( .A(n9328), .B(n9329), .Z(n9323) );
  NANDN U1688 ( .A(n9621), .B(n9620), .Z(n723) );
  NANDN U1689 ( .A(n9619), .B(n9618), .Z(n724) );
  NAND U1690 ( .A(n723), .B(n724), .Z(n9771) );
  XNOR U1691 ( .A(n9921), .B(n9922), .Z(n9916) );
  NAND U1692 ( .A(n10215), .B(n10216), .Z(n725) );
  NANDN U1693 ( .A(n10218), .B(n10217), .Z(n726) );
  NAND U1694 ( .A(n725), .B(n726), .Z(n10467) );
  NANDN U1695 ( .A(n10746), .B(n10745), .Z(n727) );
  NANDN U1696 ( .A(n10744), .B(n10743), .Z(n728) );
  NAND U1697 ( .A(n727), .B(n728), .Z(n10898) );
  NAND U1698 ( .A(n10788), .B(n10789), .Z(n729) );
  NANDN U1699 ( .A(n10791), .B(n10790), .Z(n730) );
  NAND U1700 ( .A(n729), .B(n730), .Z(n11048) );
  XNOR U1701 ( .A(n11084), .B(n11085), .Z(n11079) );
  XNOR U1702 ( .A(n11352), .B(n11353), .Z(n11347) );
  NAND U1703 ( .A(n11778), .B(n11777), .Z(n731) );
  NANDN U1704 ( .A(n11776), .B(n11775), .Z(n732) );
  NAND U1705 ( .A(n731), .B(n732), .Z(n11931) );
  XNOR U1706 ( .A(n12229), .B(n12230), .Z(n12224) );
  XNOR U1707 ( .A(n12526), .B(n12527), .Z(n12521) );
  NAND U1708 ( .A(n12895), .B(n12896), .Z(n733) );
  NANDN U1709 ( .A(n12894), .B(n12893), .Z(n734) );
  NAND U1710 ( .A(n733), .B(n734), .Z(n13103) );
  XNOR U1711 ( .A(n13401), .B(n13402), .Z(n13396) );
  XNOR U1712 ( .A(n13695), .B(n13696), .Z(n13690) );
  XNOR U1713 ( .A(n13844), .B(n13845), .Z(n13839) );
  XNOR U1714 ( .A(n14136), .B(n14137), .Z(n14131) );
  XNOR U1715 ( .A(n14281), .B(n14282), .Z(n14276) );
  NAND U1716 ( .A(n14308), .B(n14309), .Z(n735) );
  NANDN U1717 ( .A(n14311), .B(n14310), .Z(n736) );
  NAND U1718 ( .A(n735), .B(n736), .Z(n14566) );
  XNOR U1719 ( .A(n14749), .B(n14750), .Z(n14744) );
  NAND U1720 ( .A(n14892), .B(n14893), .Z(n737) );
  NANDN U1721 ( .A(n14895), .B(n14894), .Z(n738) );
  NAND U1722 ( .A(n737), .B(n738), .Z(n15145) );
  XNOR U1723 ( .A(n15595), .B(n15596), .Z(n15590) );
  NAND U1724 ( .A(n15725), .B(n15724), .Z(n739) );
  NAND U1725 ( .A(n15722), .B(n15723), .Z(n740) );
  NAND U1726 ( .A(n739), .B(n740), .Z(n15760) );
  XNOR U1727 ( .A(n15916), .B(n15917), .Z(n15911) );
  NAND U1728 ( .A(n16210), .B(n16211), .Z(n741) );
  NANDN U1729 ( .A(n16213), .B(n16212), .Z(n742) );
  NAND U1730 ( .A(n741), .B(n742), .Z(n16350) );
  XNOR U1731 ( .A(n16506), .B(n16507), .Z(n16501) );
  NAND U1732 ( .A(n16649), .B(n16650), .Z(n743) );
  NANDN U1733 ( .A(n16652), .B(n16651), .Z(n744) );
  NAND U1734 ( .A(n743), .B(n744), .Z(n16901) );
  OR U1735 ( .A(n16834), .B(n16835), .Z(n745) );
  NAND U1736 ( .A(n16833), .B(n16832), .Z(n746) );
  NAND U1737 ( .A(n745), .B(n746), .Z(n16927) );
  XNOR U1738 ( .A(n17195), .B(n17196), .Z(n17190) );
  OR U1739 ( .A(n17275), .B(n17274), .Z(n747) );
  NANDN U1740 ( .A(n17277), .B(n17276), .Z(n748) );
  NAND U1741 ( .A(n747), .B(n748), .Z(n17488) );
  NAND U1742 ( .A(n17619), .B(n17618), .Z(n749) );
  NANDN U1743 ( .A(n17617), .B(n17616), .Z(n750) );
  NAND U1744 ( .A(n749), .B(n750), .Z(n17768) );
  OR U1745 ( .A(n17657), .B(n17658), .Z(n751) );
  NAND U1746 ( .A(n17656), .B(n17655), .Z(n752) );
  NAND U1747 ( .A(n751), .B(n752), .Z(n17910) );
  OR U1748 ( .A(n17845), .B(n17846), .Z(n753) );
  NAND U1749 ( .A(n17844), .B(n17843), .Z(n754) );
  NAND U1750 ( .A(n753), .B(n754), .Z(n18055) );
  NAND U1751 ( .A(n18203), .B(n18202), .Z(n755) );
  NAND U1752 ( .A(n18200), .B(n18201), .Z(n756) );
  NAND U1753 ( .A(n755), .B(n756), .Z(n18346) );
  NAND U1754 ( .A(n18380), .B(n18381), .Z(n757) );
  NANDN U1755 ( .A(n18383), .B(n18382), .Z(n758) );
  NAND U1756 ( .A(n757), .B(n758), .Z(n18630) );
  NAND U1757 ( .A(n18714), .B(n18715), .Z(n759) );
  NANDN U1758 ( .A(n18713), .B(n18712), .Z(n760) );
  NAND U1759 ( .A(n759), .B(n760), .Z(n18914) );
  NAND U1760 ( .A(n18804), .B(n18803), .Z(n761) );
  NAND U1761 ( .A(n18801), .B(n18802), .Z(n762) );
  NAND U1762 ( .A(n761), .B(n762), .Z(n19054) );
  XNOR U1763 ( .A(n19502), .B(n19503), .Z(n19497) );
  OR U1764 ( .A(n19716), .B(n19717), .Z(n763) );
  NAND U1765 ( .A(n19715), .B(n19714), .Z(n764) );
  NAND U1766 ( .A(n763), .B(n764), .Z(n19922) );
  NAND U1767 ( .A(n19816), .B(n19815), .Z(n765) );
  NAND U1768 ( .A(n19813), .B(n19814), .Z(n766) );
  NAND U1769 ( .A(n765), .B(n766), .Z(n20070) );
  NAND U1770 ( .A(n20249), .B(n20250), .Z(n767) );
  NANDN U1771 ( .A(n20252), .B(n20251), .Z(n768) );
  NAND U1772 ( .A(n767), .B(n768), .Z(n20388) );
  XNOR U1773 ( .A(n20542), .B(n20543), .Z(n20537) );
  XNOR U1774 ( .A(n20805), .B(n20806), .Z(n20800) );
  NAND U1775 ( .A(n20832), .B(n20833), .Z(n769) );
  NANDN U1776 ( .A(n20835), .B(n20834), .Z(n770) );
  NAND U1777 ( .A(n769), .B(n770), .Z(n20970) );
  XNOR U1778 ( .A(n21242), .B(n21243), .Z(n21237) );
  XNOR U1779 ( .A(n21387), .B(n21388), .Z(n21382) );
  NAND U1780 ( .A(n21414), .B(n21415), .Z(n771) );
  NANDN U1781 ( .A(n21417), .B(n21416), .Z(n772) );
  NAND U1782 ( .A(n771), .B(n772), .Z(n21552) );
  XNOR U1783 ( .A(n21822), .B(n21823), .Z(n21817) );
  NAND U1784 ( .A(n21849), .B(n21850), .Z(n773) );
  NANDN U1785 ( .A(n21852), .B(n21851), .Z(n774) );
  NAND U1786 ( .A(n773), .B(n774), .Z(n22101) );
  XNOR U1787 ( .A(n22281), .B(n22282), .Z(n22276) );
  NAND U1788 ( .A(n22534), .B(n22533), .Z(n775) );
  NAND U1789 ( .A(n22531), .B(n22532), .Z(n776) );
  NAND U1790 ( .A(n775), .B(n776), .Z(n22569) );
  XNOR U1791 ( .A(n22874), .B(n22875), .Z(n22869) );
  NAND U1792 ( .A(n23017), .B(n23018), .Z(n777) );
  NANDN U1793 ( .A(n23020), .B(n23019), .Z(n778) );
  NAND U1794 ( .A(n777), .B(n778), .Z(n23267) );
  NAND U1795 ( .A(n23351), .B(n23352), .Z(n779) );
  NANDN U1796 ( .A(n23350), .B(n23349), .Z(n780) );
  NAND U1797 ( .A(n779), .B(n780), .Z(n23554) );
  OR U1798 ( .A(n23435), .B(n23436), .Z(n781) );
  NAND U1799 ( .A(n23434), .B(n23433), .Z(n782) );
  NAND U1800 ( .A(n781), .B(n782), .Z(n23693) );
  XNOR U1801 ( .A(n24023), .B(n24024), .Z(n24018) );
  NAND U1802 ( .A(n24515), .B(n24516), .Z(n783) );
  NANDN U1803 ( .A(n24514), .B(n24513), .Z(n784) );
  NAND U1804 ( .A(n783), .B(n784), .Z(n24724) );
  NAND U1805 ( .A(n24857), .B(n24856), .Z(n785) );
  NAND U1806 ( .A(n24854), .B(n24855), .Z(n786) );
  NAND U1807 ( .A(n785), .B(n786), .Z(n25012) );
  XNOR U1808 ( .A(n25164), .B(n25165), .Z(n25159) );
  NAND U1809 ( .A(n25191), .B(n25192), .Z(n787) );
  NANDN U1810 ( .A(n25194), .B(n25193), .Z(n788) );
  NAND U1811 ( .A(n787), .B(n788), .Z(n25330) );
  XNOR U1812 ( .A(n25485), .B(n25486), .Z(n25480) );
  OR U1813 ( .A(n25823), .B(n25824), .Z(n789) );
  NAND U1814 ( .A(n25822), .B(n25821), .Z(n790) );
  NAND U1815 ( .A(n789), .B(n790), .Z(n25915) );
  NAND U1816 ( .A(n26173), .B(n26172), .Z(n791) );
  NAND U1817 ( .A(n26170), .B(n26171), .Z(n792) );
  NAND U1818 ( .A(n791), .B(n792), .Z(n26208) );
  NAND U1819 ( .A(n26360), .B(n26361), .Z(n793) );
  NANDN U1820 ( .A(n26363), .B(n26362), .Z(n794) );
  NAND U1821 ( .A(n793), .B(n794), .Z(n26610) );
  OR U1822 ( .A(n26497), .B(n26498), .Z(n795) );
  NAND U1823 ( .A(n26496), .B(n26495), .Z(n796) );
  NAND U1824 ( .A(n795), .B(n796), .Z(n26750) );
  NAND U1825 ( .A(n26749), .B(n26748), .Z(n797) );
  NANDN U1826 ( .A(n26747), .B(n26746), .Z(n798) );
  NAND U1827 ( .A(n797), .B(n798), .Z(n26899) );
  XNOR U1828 ( .A(n26929), .B(n26930), .Z(n26924) );
  XNOR U1829 ( .A(n27348), .B(n27349), .Z(n27343) );
  XNOR U1830 ( .A(n27524), .B(n27525), .Z(n27519) );
  XNOR U1831 ( .A(n27791), .B(n27792), .Z(n27786) );
  NAND U1832 ( .A(n27963), .B(n27964), .Z(n799) );
  NANDN U1833 ( .A(n27966), .B(n27965), .Z(n800) );
  NAND U1834 ( .A(n799), .B(n800), .Z(n28101) );
  XNOR U1835 ( .A(n28673), .B(n28674), .Z(n28668) );
  XNOR U1836 ( .A(n28702), .B(n28703), .Z(n28697) );
  NAND U1837 ( .A(n28952), .B(n28951), .Z(n801) );
  NANDN U1838 ( .A(n28950), .B(n28949), .Z(n802) );
  NAND U1839 ( .A(n801), .B(n802), .Z(n29103) );
  NAND U1840 ( .A(n29234), .B(n29233), .Z(n803) );
  NANDN U1841 ( .A(n29232), .B(n29231), .Z(n804) );
  NAND U1842 ( .A(n803), .B(n804), .Z(n29383) );
  NAND U1843 ( .A(n29276), .B(n29277), .Z(n805) );
  NANDN U1844 ( .A(n29279), .B(n29278), .Z(n806) );
  NAND U1845 ( .A(n805), .B(n806), .Z(n29526) );
  NAND U1846 ( .A(n29612), .B(n29613), .Z(n807) );
  NANDN U1847 ( .A(n29611), .B(n29610), .Z(n808) );
  NAND U1848 ( .A(n807), .B(n808), .Z(n29700) );
  NAND U1849 ( .A(n29844), .B(n29845), .Z(n809) );
  NANDN U1850 ( .A(n29847), .B(n29846), .Z(n810) );
  NAND U1851 ( .A(n809), .B(n810), .Z(n30098) );
  NAND U1852 ( .A(n30132), .B(n30133), .Z(n811) );
  NANDN U1853 ( .A(n30135), .B(n30134), .Z(n812) );
  NAND U1854 ( .A(n811), .B(n812), .Z(n30382) );
  OR U1855 ( .A(n30269), .B(n30270), .Z(n813) );
  NAND U1856 ( .A(n30268), .B(n30267), .Z(n814) );
  NAND U1857 ( .A(n813), .B(n814), .Z(n30522) );
  NAND U1858 ( .A(n30521), .B(n30520), .Z(n815) );
  NANDN U1859 ( .A(n30519), .B(n30518), .Z(n816) );
  NAND U1860 ( .A(n815), .B(n816), .Z(n30552) );
  XNOR U1861 ( .A(n30700), .B(n30701), .Z(n30695) );
  NAND U1862 ( .A(n30843), .B(n30844), .Z(n817) );
  NANDN U1863 ( .A(n30846), .B(n30845), .Z(n818) );
  NAND U1864 ( .A(n817), .B(n818), .Z(n31102) );
  NAND U1865 ( .A(n31388), .B(n31387), .Z(n819) );
  NANDN U1866 ( .A(n31386), .B(n31385), .Z(n820) );
  NAND U1867 ( .A(n819), .B(n820), .Z(n31541) );
  XNOR U1868 ( .A(n31692), .B(n31693), .Z(n31687) );
  NAND U1869 ( .A(n31822), .B(n31821), .Z(n821) );
  NAND U1870 ( .A(n31819), .B(n31820), .Z(n822) );
  NAND U1871 ( .A(n821), .B(n822), .Z(n31857) );
  NAND U1872 ( .A(n32009), .B(n32010), .Z(n823) );
  NANDN U1873 ( .A(n32012), .B(n32011), .Z(n824) );
  NAND U1874 ( .A(n823), .B(n824), .Z(n32260) );
  NAND U1875 ( .A(n32153), .B(n32152), .Z(n825) );
  NAND U1876 ( .A(n32150), .B(n32151), .Z(n826) );
  NAND U1877 ( .A(n825), .B(n826), .Z(n32409) );
  XNOR U1878 ( .A(n32592), .B(n32593), .Z(n32587) );
  XNOR U1879 ( .A(n32856), .B(n32857), .Z(n32851) );
  OR U1880 ( .A(n32927), .B(n32928), .Z(n827) );
  NAND U1881 ( .A(n32926), .B(n32925), .Z(n828) );
  NAND U1882 ( .A(n827), .B(n828), .Z(n33022) );
  XNOR U1883 ( .A(n33298), .B(n33299), .Z(n33293) );
  XNOR U1884 ( .A(n33590), .B(n33591), .Z(n33585) );
  OR U1885 ( .A(n33659), .B(n33660), .Z(n829) );
  NAND U1886 ( .A(n33658), .B(n33657), .Z(n830) );
  NAND U1887 ( .A(n829), .B(n830), .Z(n33862) );
  NAND U1888 ( .A(n33759), .B(n33758), .Z(n831) );
  NAND U1889 ( .A(n33756), .B(n33757), .Z(n832) );
  NAND U1890 ( .A(n831), .B(n832), .Z(n34006) );
  XNOR U1891 ( .A(n34303), .B(n34304), .Z(n34298) );
  XNOR U1892 ( .A(n34332), .B(n34333), .Z(n34327) );
  XNOR U1893 ( .A(n34630), .B(n34631), .Z(n34625) );
  OR U1894 ( .A(n34824), .B(n34823), .Z(n833) );
  NANDN U1895 ( .A(n34826), .B(n34825), .Z(n834) );
  NAND U1896 ( .A(n833), .B(n834), .Z(n34917) );
  NAND U1897 ( .A(n35359), .B(n35360), .Z(n835) );
  NANDN U1898 ( .A(n35362), .B(n35361), .Z(n836) );
  NAND U1899 ( .A(n835), .B(n836), .Z(n35610) );
  XNOR U1900 ( .A(n36717), .B(n36718), .Z(n36736) );
  XOR U1901 ( .A(n37597), .B(n37598), .Z(n37599) );
  NANDN U1902 ( .A(n1051), .B(a[0]), .Z(n837) );
  AND U1903 ( .A(b[7]), .B(n837), .Z(n838) );
  XNOR U1904 ( .A(a[0]), .B(n1051), .Z(n839) );
  NAND U1905 ( .A(n839), .B(b[6]), .Z(n840) );
  NAND U1906 ( .A(n838), .B(n840), .Z(n1214) );
  NANDN U1907 ( .A(n3393), .B(b[10]), .Z(n841) );
  AND U1908 ( .A(b[11]), .B(n841), .Z(n842) );
  XNOR U1909 ( .A(b[10]), .B(n3393), .Z(n843) );
  NAND U1910 ( .A(n843), .B(b[9]), .Z(n844) );
  NAND U1911 ( .A(n842), .B(n844), .Z(n1396) );
  NAND U1912 ( .A(n1721), .B(n1720), .Z(n845) );
  NANDN U1913 ( .A(n1719), .B(n1718), .Z(n846) );
  NAND U1914 ( .A(n845), .B(n846), .Z(n1848) );
  NANDN U1915 ( .A(n2929), .B(n2928), .Z(n847) );
  NANDN U1916 ( .A(n2931), .B(n2930), .Z(n848) );
  AND U1917 ( .A(n847), .B(n848), .Z(n2950) );
  NANDN U1918 ( .A(n4893), .B(n4892), .Z(n849) );
  NANDN U1919 ( .A(n4895), .B(n4894), .Z(n850) );
  NAND U1920 ( .A(n849), .B(n850), .Z(n4913) );
  NANDN U1921 ( .A(n5204), .B(n5203), .Z(n851) );
  NANDN U1922 ( .A(n5206), .B(n5205), .Z(n852) );
  NAND U1923 ( .A(n851), .B(n852), .Z(n5342) );
  NANDN U1924 ( .A(n8444), .B(n8443), .Z(n853) );
  NANDN U1925 ( .A(n8446), .B(n8445), .Z(n854) );
  AND U1926 ( .A(n853), .B(n854), .Z(n8576) );
  NANDN U1927 ( .A(n10612), .B(n10611), .Z(n855) );
  NANDN U1928 ( .A(n10614), .B(n10613), .Z(n856) );
  NAND U1929 ( .A(n855), .B(n856), .Z(n10632) );
  NANDN U1930 ( .A(n11927), .B(n11926), .Z(n857) );
  NANDN U1931 ( .A(n11929), .B(n11928), .Z(n858) );
  NAND U1932 ( .A(n857), .B(n858), .Z(n11945) );
  NANDN U1933 ( .A(n12950), .B(n12949), .Z(n859) );
  NANDN U1934 ( .A(n12952), .B(n12951), .Z(n860) );
  NAND U1935 ( .A(n859), .B(n860), .Z(n12970) );
  NAND U1936 ( .A(n15291), .B(n15292), .Z(n861) );
  NANDN U1937 ( .A(n15290), .B(n15289), .Z(n862) );
  NAND U1938 ( .A(n861), .B(n862), .Z(n15310) );
  NANDN U1939 ( .A(n18769), .B(n18768), .Z(n863) );
  NANDN U1940 ( .A(n18771), .B(n18770), .Z(n864) );
  NAND U1941 ( .A(n863), .B(n864), .Z(n18789) );
  NAND U1942 ( .A(n19200), .B(n19201), .Z(n865) );
  NANDN U1943 ( .A(n19199), .B(n19198), .Z(n866) );
  NAND U1944 ( .A(n865), .B(n866), .Z(n19219) );
  NANDN U1945 ( .A(n22247), .B(n22246), .Z(n867) );
  NANDN U1946 ( .A(n22249), .B(n22248), .Z(n868) );
  NAND U1947 ( .A(n867), .B(n868), .Z(n22267) );
  NANDN U1948 ( .A(n23407), .B(n23406), .Z(n869) );
  NANDN U1949 ( .A(n23409), .B(n23408), .Z(n870) );
  NAND U1950 ( .A(n869), .B(n870), .Z(n23427) );
  NANDN U1951 ( .A(n23719), .B(n23718), .Z(n871) );
  NANDN U1952 ( .A(n23721), .B(n23720), .Z(n872) );
  NAND U1953 ( .A(n871), .B(n872), .Z(n23859) );
  NANDN U1954 ( .A(n24571), .B(n24570), .Z(n873) );
  NANDN U1955 ( .A(n24573), .B(n24572), .Z(n874) );
  NAND U1956 ( .A(n873), .B(n874), .Z(n24591) );
  NANDN U1957 ( .A(n26895), .B(n26894), .Z(n875) );
  NANDN U1958 ( .A(n26897), .B(n26896), .Z(n876) );
  NAND U1959 ( .A(n875), .B(n876), .Z(n26915) );
  NAND U1960 ( .A(n29100), .B(n29101), .Z(n877) );
  NANDN U1961 ( .A(n29099), .B(n29098), .Z(n878) );
  NAND U1962 ( .A(n877), .B(n878), .Z(n29119) );
  NANDN U1963 ( .A(n29667), .B(n29666), .Z(n879) );
  NANDN U1964 ( .A(n29669), .B(n29668), .Z(n880) );
  NAND U1965 ( .A(n879), .B(n880), .Z(n29687) );
  NANDN U1966 ( .A(n30548), .B(n30547), .Z(n881) );
  NANDN U1967 ( .A(n30550), .B(n30549), .Z(n882) );
  NAND U1968 ( .A(n881), .B(n882), .Z(n30686) );
  NANDN U1969 ( .A(n31537), .B(n31536), .Z(n883) );
  NANDN U1970 ( .A(n31539), .B(n31538), .Z(n884) );
  NAND U1971 ( .A(n883), .B(n884), .Z(n31557) );
  NANDN U1972 ( .A(n34033), .B(n34032), .Z(n885) );
  NANDN U1973 ( .A(n34035), .B(n34034), .Z(n886) );
  NAND U1974 ( .A(n885), .B(n886), .Z(n34171) );
  NAND U1975 ( .A(n35504), .B(n35503), .Z(n887) );
  NAND U1976 ( .A(n35501), .B(n35502), .Z(n888) );
  NAND U1977 ( .A(n887), .B(n888), .Z(n35759) );
  NAND U1978 ( .A(n36538), .B(n36537), .Z(n889) );
  NANDN U1979 ( .A(n36536), .B(n36535), .Z(n890) );
  NAND U1980 ( .A(n889), .B(n890), .Z(n36748) );
  NAND U1981 ( .A(n37032), .B(n37033), .Z(n891) );
  NANDN U1982 ( .A(n37035), .B(n37034), .Z(n892) );
  NAND U1983 ( .A(n891), .B(n892), .Z(n37225) );
  NAND U1984 ( .A(n37167), .B(n37166), .Z(n893) );
  NANDN U1985 ( .A(n37165), .B(n37164), .Z(n894) );
  NAND U1986 ( .A(n893), .B(n894), .Z(n37260) );
  NAND U1987 ( .A(n37338), .B(n37337), .Z(n895) );
  NANDN U1988 ( .A(n37336), .B(n37335), .Z(n896) );
  AND U1989 ( .A(n895), .B(n896), .Z(n37370) );
  NAND U1990 ( .A(n37282), .B(n37281), .Z(n897) );
  NANDN U1991 ( .A(n37280), .B(n37279), .Z(n898) );
  NAND U1992 ( .A(n897), .B(n898), .Z(n37361) );
  NAND U1993 ( .A(n37380), .B(n37379), .Z(n899) );
  NANDN U1994 ( .A(n37378), .B(n37377), .Z(n900) );
  NAND U1995 ( .A(n899), .B(n900), .Z(n37526) );
  NAND U1996 ( .A(n37457), .B(n37458), .Z(n901) );
  NANDN U1997 ( .A(n37456), .B(n37455), .Z(n902) );
  NAND U1998 ( .A(n901), .B(n902), .Z(n37554) );
  NAND U1999 ( .A(n1171), .B(n1170), .Z(n903) );
  NANDN U2000 ( .A(n1169), .B(n1168), .Z(n904) );
  NAND U2001 ( .A(n903), .B(n904), .Z(n1211) );
  NAND U2002 ( .A(n2959), .B(n2958), .Z(n905) );
  NANDN U2003 ( .A(n2957), .B(n2956), .Z(n906) );
  NAND U2004 ( .A(n905), .B(n906), .Z(n3198) );
  NAND U2005 ( .A(n35790), .B(n35789), .Z(n907) );
  NANDN U2006 ( .A(n35788), .B(n35787), .Z(n908) );
  NAND U2007 ( .A(n907), .B(n908), .Z(n36055) );
  NAND U2008 ( .A(n36476), .B(n36475), .Z(n909) );
  NAND U2009 ( .A(n36473), .B(n36474), .Z(n910) );
  NAND U2010 ( .A(n909), .B(n910), .Z(n36497) );
  NAND U2011 ( .A(n36516), .B(n36515), .Z(n911) );
  NAND U2012 ( .A(n36513), .B(n36514), .Z(n912) );
  NAND U2013 ( .A(n911), .B(n912), .Z(n36632) );
  NANDN U2014 ( .A(n36782), .B(n36781), .Z(n913) );
  NANDN U2015 ( .A(n36780), .B(n36779), .Z(n914) );
  NAND U2016 ( .A(n913), .B(n914), .Z(n36893) );
  NAND U2017 ( .A(n36901), .B(n36900), .Z(n915) );
  NANDN U2018 ( .A(n36899), .B(n36898), .Z(n916) );
  NAND U2019 ( .A(n915), .B(n916), .Z(n37008) );
  OR U2020 ( .A(n37264), .B(n37263), .Z(n917) );
  NAND U2021 ( .A(n37266), .B(n37265), .Z(n918) );
  NAND U2022 ( .A(n917), .B(n918), .Z(n37439) );
  NAND U2023 ( .A(n37376), .B(n37375), .Z(n919) );
  NANDN U2024 ( .A(n37374), .B(n37373), .Z(n920) );
  AND U2025 ( .A(n919), .B(n920), .Z(n37529) );
  NANDN U2026 ( .A(n37737), .B(n37736), .Z(n921) );
  NANDN U2027 ( .A(n37735), .B(n37734), .Z(n922) );
  NAND U2028 ( .A(n921), .B(n922), .Z(n37878) );
  NANDN U2029 ( .A(n38226), .B(n38225), .Z(n923) );
  NANDN U2030 ( .A(n38224), .B(n38223), .Z(n924) );
  AND U2031 ( .A(n923), .B(n924), .Z(n38250) );
  NAND U2032 ( .A(n38387), .B(n38386), .Z(n925) );
  NANDN U2033 ( .A(n38385), .B(n38384), .Z(n926) );
  NAND U2034 ( .A(n925), .B(n926), .Z(n38403) );
  NANDN U2035 ( .A(a[0]), .B(n36107), .Z(n927) );
  OR U2036 ( .A(b[1]), .B(b[2]), .Z(n928) );
  NAND U2037 ( .A(n928), .B(n927), .Z(n929) );
  NANDN U2038 ( .A(n1050), .B(n929), .Z(n1104) );
  NAND U2039 ( .A(n1335), .B(n1334), .Z(n930) );
  NANDN U2040 ( .A(n1333), .B(n1332), .Z(n931) );
  NAND U2041 ( .A(n930), .B(n931), .Z(n1384) );
  NAND U2042 ( .A(n1774), .B(n1773), .Z(n932) );
  NANDN U2043 ( .A(n1772), .B(n1771), .Z(n933) );
  AND U2044 ( .A(n932), .B(n933), .Z(n1786) );
  NAND U2045 ( .A(n3777), .B(n3776), .Z(n934) );
  NANDN U2046 ( .A(n3775), .B(n3774), .Z(n935) );
  NAND U2047 ( .A(n934), .B(n935), .Z(n3914) );
  NAND U2048 ( .A(n4773), .B(n4772), .Z(n936) );
  NAND U2049 ( .A(n4770), .B(n4771), .Z(n937) );
  NAND U2050 ( .A(n936), .B(n937), .Z(n4910) );
  NAND U2051 ( .A(n5196), .B(n5195), .Z(n938) );
  NAND U2052 ( .A(n5193), .B(n5194), .Z(n939) );
  NAND U2053 ( .A(n938), .B(n939), .Z(n5339) );
  NAND U2054 ( .A(n5929), .B(n5928), .Z(n940) );
  NAND U2055 ( .A(n5926), .B(n5927), .Z(n941) );
  NAND U2056 ( .A(n940), .B(n941), .Z(n6074) );
  NAND U2057 ( .A(n7250), .B(n7249), .Z(n942) );
  NAND U2058 ( .A(n7247), .B(n7248), .Z(n943) );
  NAND U2059 ( .A(n942), .B(n943), .Z(n7395) );
  NAND U2060 ( .A(n10486), .B(n10485), .Z(n944) );
  NAND U2061 ( .A(n10483), .B(n10484), .Z(n945) );
  NAND U2062 ( .A(n944), .B(n945), .Z(n10629) );
  NAND U2063 ( .A(n11364), .B(n11363), .Z(n946) );
  NAND U2064 ( .A(n11361), .B(n11362), .Z(n947) );
  NAND U2065 ( .A(n946), .B(n947), .Z(n11511) );
  NAND U2066 ( .A(n11799), .B(n11798), .Z(n948) );
  NAND U2067 ( .A(n11796), .B(n11797), .Z(n949) );
  NAND U2068 ( .A(n948), .B(n949), .Z(n11944) );
  NAND U2069 ( .A(n12241), .B(n12240), .Z(n950) );
  NAND U2070 ( .A(n12238), .B(n12239), .Z(n951) );
  NAND U2071 ( .A(n950), .B(n951), .Z(n12388) );
  NAND U2072 ( .A(n12828), .B(n12827), .Z(n952) );
  NAND U2073 ( .A(n12825), .B(n12826), .Z(n953) );
  NAND U2074 ( .A(n952), .B(n953), .Z(n12967) );
  NAND U2075 ( .A(n13413), .B(n13412), .Z(n954) );
  NAND U2076 ( .A(n13410), .B(n13411), .Z(n955) );
  NAND U2077 ( .A(n954), .B(n955), .Z(n13560) );
  NAND U2078 ( .A(n13856), .B(n13855), .Z(n956) );
  NAND U2079 ( .A(n13853), .B(n13854), .Z(n957) );
  NAND U2080 ( .A(n956), .B(n957), .Z(n14003) );
  NAND U2081 ( .A(n15164), .B(n15163), .Z(n958) );
  NAND U2082 ( .A(n15161), .B(n15162), .Z(n959) );
  NAND U2083 ( .A(n958), .B(n959), .Z(n15307) );
  NAND U2084 ( .A(n15752), .B(n15751), .Z(n960) );
  NAND U2085 ( .A(n15749), .B(n15750), .Z(n961) );
  NAND U2086 ( .A(n960), .B(n961), .Z(n15899) );
  NAND U2087 ( .A(n17207), .B(n17206), .Z(n962) );
  NAND U2088 ( .A(n17204), .B(n17205), .Z(n963) );
  NAND U2089 ( .A(n962), .B(n963), .Z(n17352) );
  NAND U2090 ( .A(n18073), .B(n18072), .Z(n964) );
  NAND U2091 ( .A(n18070), .B(n18071), .Z(n965) );
  NAND U2092 ( .A(n964), .B(n965), .Z(n18218) );
  NAND U2093 ( .A(n18649), .B(n18648), .Z(n966) );
  NAND U2094 ( .A(n18646), .B(n18647), .Z(n967) );
  NAND U2095 ( .A(n966), .B(n967), .Z(n18786) );
  NAND U2096 ( .A(n19073), .B(n19072), .Z(n968) );
  NAND U2097 ( .A(n19070), .B(n19071), .Z(n969) );
  NAND U2098 ( .A(n968), .B(n969), .Z(n19216) );
  NAND U2099 ( .A(n19514), .B(n19513), .Z(n970) );
  NAND U2100 ( .A(n19511), .B(n19512), .Z(n971) );
  NAND U2101 ( .A(n970), .B(n971), .Z(n19659) );
  NAND U2102 ( .A(n20089), .B(n20088), .Z(n972) );
  NAND U2103 ( .A(n20086), .B(n20087), .Z(n973) );
  NAND U2104 ( .A(n972), .B(n973), .Z(n20234) );
  NAND U2105 ( .A(n22120), .B(n22119), .Z(n974) );
  NAND U2106 ( .A(n22117), .B(n22118), .Z(n975) );
  NAND U2107 ( .A(n974), .B(n975), .Z(n22264) );
  NAND U2108 ( .A(n22561), .B(n22560), .Z(n976) );
  NAND U2109 ( .A(n22558), .B(n22559), .Z(n977) );
  NAND U2110 ( .A(n976), .B(n977), .Z(n22708) );
  NAND U2111 ( .A(n23286), .B(n23285), .Z(n978) );
  NAND U2112 ( .A(n23283), .B(n23284), .Z(n979) );
  NAND U2113 ( .A(n978), .B(n979), .Z(n23424) );
  NAND U2114 ( .A(n23711), .B(n23710), .Z(n980) );
  NAND U2115 ( .A(n23708), .B(n23709), .Z(n981) );
  NAND U2116 ( .A(n980), .B(n981), .Z(n23856) );
  NAND U2117 ( .A(n24448), .B(n24447), .Z(n982) );
  NAND U2118 ( .A(n24445), .B(n24446), .Z(n983) );
  NAND U2119 ( .A(n982), .B(n983), .Z(n24588) );
  NAND U2120 ( .A(n24884), .B(n24883), .Z(n984) );
  NAND U2121 ( .A(n24881), .B(n24882), .Z(n985) );
  NAND U2122 ( .A(n984), .B(n985), .Z(n25031) );
  NAND U2123 ( .A(n26200), .B(n26199), .Z(n986) );
  NAND U2124 ( .A(n26197), .B(n26198), .Z(n987) );
  NAND U2125 ( .A(n986), .B(n987), .Z(n26345) );
  NAND U2126 ( .A(n26768), .B(n26767), .Z(n988) );
  NAND U2127 ( .A(n26765), .B(n26766), .Z(n989) );
  NAND U2128 ( .A(n988), .B(n989), .Z(n26912) );
  NAND U2129 ( .A(n27360), .B(n27359), .Z(n990) );
  NAND U2130 ( .A(n27357), .B(n27358), .Z(n991) );
  NAND U2131 ( .A(n990), .B(n991), .Z(n27507) );
  NAND U2132 ( .A(n27803), .B(n27802), .Z(n992) );
  NAND U2133 ( .A(n27800), .B(n27801), .Z(n993) );
  NAND U2134 ( .A(n992), .B(n993), .Z(n27948) );
  NAND U2135 ( .A(n28973), .B(n28972), .Z(n994) );
  NAND U2136 ( .A(n28970), .B(n28971), .Z(n995) );
  NAND U2137 ( .A(n994), .B(n995), .Z(n29116) );
  NAND U2138 ( .A(n29545), .B(n29544), .Z(n996) );
  NAND U2139 ( .A(n29542), .B(n29543), .Z(n997) );
  NAND U2140 ( .A(n996), .B(n997), .Z(n29684) );
  NAND U2141 ( .A(n30540), .B(n30539), .Z(n998) );
  NAND U2142 ( .A(n30537), .B(n30538), .Z(n999) );
  NAND U2143 ( .A(n998), .B(n999), .Z(n30683) );
  NAND U2144 ( .A(n31409), .B(n31408), .Z(n1000) );
  NAND U2145 ( .A(n31406), .B(n31407), .Z(n1001) );
  NAND U2146 ( .A(n1000), .B(n1001), .Z(n31554) );
  NAND U2147 ( .A(n31849), .B(n31848), .Z(n1002) );
  NAND U2148 ( .A(n31846), .B(n31847), .Z(n1003) );
  NAND U2149 ( .A(n1002), .B(n1003), .Z(n31994) );
  NAND U2150 ( .A(n32428), .B(n32427), .Z(n1004) );
  NAND U2151 ( .A(n32425), .B(n32426), .Z(n1005) );
  NAND U2152 ( .A(n1004), .B(n1005), .Z(n32575) );
  NAND U2153 ( .A(n33310), .B(n33309), .Z(n1006) );
  NAND U2154 ( .A(n33307), .B(n33308), .Z(n1007) );
  NAND U2155 ( .A(n1006), .B(n1007), .Z(n33457) );
  NAND U2156 ( .A(n34025), .B(n34024), .Z(n1008) );
  NAND U2157 ( .A(n34022), .B(n34023), .Z(n1009) );
  NAND U2158 ( .A(n1008), .B(n1009), .Z(n34168) );
  NAND U2159 ( .A(n35199), .B(n35198), .Z(n1010) );
  NAND U2160 ( .A(n35196), .B(n35197), .Z(n1011) );
  NAND U2161 ( .A(n1010), .B(n1011), .Z(n35344) );
  NAND U2162 ( .A(n36218), .B(n36219), .Z(n1012) );
  NANDN U2163 ( .A(n36217), .B(n36216), .Z(n1013) );
  NAND U2164 ( .A(n1012), .B(n1013), .Z(n36355) );
  OR U2165 ( .A(n38469), .B(n38470), .Z(n1014) );
  NAND U2166 ( .A(n38468), .B(n38467), .Z(n1015) );
  NAND U2167 ( .A(n1014), .B(n1015), .Z(n38501) );
  ANDN U2168 ( .B(n1103), .A(n1102), .Z(n1109) );
  NAND U2169 ( .A(n1639), .B(n1638), .Z(n1016) );
  NANDN U2170 ( .A(n1637), .B(n1636), .Z(n1017) );
  NAND U2171 ( .A(n1016), .B(n1017), .Z(n1703) );
  NAND U2172 ( .A(n1961), .B(n1960), .Z(n1018) );
  NANDN U2173 ( .A(n1959), .B(n1958), .Z(n1019) );
  NAND U2174 ( .A(n1018), .B(n1019), .Z(n2043) );
  NAND U2175 ( .A(n2358), .B(n2357), .Z(n1020) );
  NANDN U2176 ( .A(n2356), .B(n2355), .Z(n1021) );
  NAND U2177 ( .A(n1020), .B(n1021), .Z(n2458) );
  NAND U2178 ( .A(n3350), .B(n3349), .Z(n1022) );
  NAND U2179 ( .A(n3347), .B(n3348), .Z(n1023) );
  NAND U2180 ( .A(n1022), .B(n1023), .Z(n3489) );
  NAND U2181 ( .A(n37003), .B(n37002), .Z(n1024) );
  XOR U2182 ( .A(n37002), .B(n37003), .Z(n1025) );
  NAND U2183 ( .A(n1025), .B(n37001), .Z(n1026) );
  NAND U2184 ( .A(n1024), .B(n1026), .Z(n37007) );
  NAND U2185 ( .A(n37238), .B(n37236), .Z(n1027) );
  XOR U2186 ( .A(n37236), .B(n37238), .Z(n1028) );
  NANDN U2187 ( .A(n37237), .B(n1028), .Z(n1029) );
  NAND U2188 ( .A(n1027), .B(n1029), .Z(n37345) );
  XOR U2189 ( .A(n37718), .B(n37717), .Z(n1030) );
  NANDN U2190 ( .A(n37716), .B(n1030), .Z(n1031) );
  NAND U2191 ( .A(n37718), .B(n37717), .Z(n1032) );
  AND U2192 ( .A(n1031), .B(n1032), .Z(n37802) );
  NAND U2193 ( .A(n37726), .B(n37727), .Z(n1033) );
  NANDN U2194 ( .A(n37725), .B(n37724), .Z(n1034) );
  NAND U2195 ( .A(n1033), .B(n1034), .Z(n37805) );
  NAND U2196 ( .A(n37966), .B(n37964), .Z(n1035) );
  XOR U2197 ( .A(n37964), .B(n37966), .Z(n1036) );
  NANDN U2198 ( .A(n37965), .B(n1036), .Z(n1037) );
  NAND U2199 ( .A(n1035), .B(n1037), .Z(n38045) );
  NAND U2200 ( .A(n38183), .B(n38181), .Z(n1038) );
  XOR U2201 ( .A(n38181), .B(n38183), .Z(n1039) );
  NANDN U2202 ( .A(n38182), .B(n1039), .Z(n1040) );
  NAND U2203 ( .A(n1038), .B(n1040), .Z(n38237) );
  XOR U2204 ( .A(n38349), .B(n38348), .Z(n1041) );
  NANDN U2205 ( .A(n38347), .B(n1041), .Z(n1042) );
  NAND U2206 ( .A(n38349), .B(n38348), .Z(n1043) );
  AND U2207 ( .A(n1042), .B(n1043), .Z(n38396) );
  NAND U2208 ( .A(n38545), .B(n38543), .Z(n1044) );
  XOR U2209 ( .A(n38543), .B(n38545), .Z(n1045) );
  NANDN U2210 ( .A(n38544), .B(n1045), .Z(n1046) );
  NAND U2211 ( .A(n1044), .B(n1046), .Z(n38581) );
  XOR U2212 ( .A(b[27]), .B(b[28]), .Z(n1047) );
  IV U2213 ( .A(n1047), .Z(n1048) );
  IV U2214 ( .A(b[0]), .Z(n1049) );
  IV U2215 ( .A(b[3]), .Z(n1050) );
  IV U2216 ( .A(b[5]), .Z(n1051) );
  IV U2217 ( .A(b[9]), .Z(n1052) );
  IV U2218 ( .A(b[13]), .Z(n1053) );
  IV U2219 ( .A(b[15]), .Z(n1054) );
  IV U2220 ( .A(b[19]), .Z(n1055) );
  IV U2221 ( .A(b[21]), .Z(n1056) );
  IV U2222 ( .A(b[23]), .Z(n1057) );
  IV U2223 ( .A(b[29]), .Z(n1058) );
  IV U2224 ( .A(b[31]), .Z(n1059) );
  NANDN U2225 ( .A(n1049), .B(a[0]), .Z(n1061) );
  XNOR U2226 ( .A(n1061), .B(sreg[224]), .Z(c[224]) );
  IV U2227 ( .A(a[0]), .Z(n3393) );
  ANDN U2228 ( .B(b[1]), .A(n3393), .Z(n1060) );
  NANDN U2229 ( .A(n1049), .B(a[1]), .Z(n1066) );
  XNOR U2230 ( .A(n1060), .B(n1066), .Z(n1069) );
  XNOR U2231 ( .A(sreg[225]), .B(n1069), .Z(n1071) );
  NANDN U2232 ( .A(n1061), .B(sreg[224]), .Z(n1070) );
  XOR U2233 ( .A(n1071), .B(n1070), .Z(c[225]) );
  NANDN U2234 ( .A(n1049), .B(a[2]), .Z(n1062) );
  XNOR U2235 ( .A(b[1]), .B(n1062), .Z(n1064) );
  NANDN U2236 ( .A(b[0]), .B(a[1]), .Z(n1063) );
  AND U2237 ( .A(n1064), .B(n1063), .Z(n1074) );
  NANDN U2238 ( .A(n3393), .B(b[2]), .Z(n1065) );
  XNOR U2239 ( .A(b[1]), .B(n1065), .Z(n1068) );
  OR U2240 ( .A(n1066), .B(a[0]), .Z(n1067) );
  AND U2241 ( .A(n1068), .B(n1067), .Z(n1075) );
  XOR U2242 ( .A(n1074), .B(n1075), .Z(n1085) );
  NAND U2243 ( .A(sreg[225]), .B(n1069), .Z(n1073) );
  OR U2244 ( .A(n1071), .B(n1070), .Z(n1072) );
  NAND U2245 ( .A(n1073), .B(n1072), .Z(n1084) );
  XNOR U2246 ( .A(n1084), .B(sreg[226]), .Z(n1086) );
  XNOR U2247 ( .A(n1085), .B(n1086), .Z(c[226]) );
  NAND U2248 ( .A(n1075), .B(n1074), .Z(n1106) );
  XOR U2249 ( .A(b[1]), .B(b[2]), .Z(n36107) );
  XNOR U2250 ( .A(n1050), .B(a[0]), .Z(n1077) );
  XNOR U2251 ( .A(n1050), .B(b[1]), .Z(n1095) );
  XNOR U2252 ( .A(n1050), .B(b[2]), .Z(n1094) );
  AND U2253 ( .A(n1095), .B(n1094), .Z(n1076) );
  NAND U2254 ( .A(n1077), .B(n1076), .Z(n1079) );
  XNOR U2255 ( .A(b[3]), .B(a[1]), .Z(n1096) );
  NANDN U2256 ( .A(n1096), .B(n36107), .Z(n1078) );
  AND U2257 ( .A(n1079), .B(n1078), .Z(n1102) );
  NANDN U2258 ( .A(n1049), .B(a[3]), .Z(n1080) );
  XNOR U2259 ( .A(b[1]), .B(n1080), .Z(n1082) );
  NANDN U2260 ( .A(b[0]), .B(a[2]), .Z(n1081) );
  AND U2261 ( .A(n1082), .B(n1081), .Z(n1103) );
  XOR U2262 ( .A(n1102), .B(n1103), .Z(n1105) );
  XOR U2263 ( .A(n1104), .B(n1105), .Z(n1083) );
  XNOR U2264 ( .A(n1106), .B(n1083), .Z(n1089) );
  XNOR U2265 ( .A(sreg[227]), .B(n1089), .Z(n1091) );
  NAND U2266 ( .A(n1084), .B(sreg[226]), .Z(n1088) );
  NANDN U2267 ( .A(n1086), .B(n1085), .Z(n1087) );
  AND U2268 ( .A(n1088), .B(n1087), .Z(n1090) );
  XOR U2269 ( .A(n1091), .B(n1090), .Z(c[227]) );
  NAND U2270 ( .A(sreg[227]), .B(n1089), .Z(n1093) );
  OR U2271 ( .A(n1091), .B(n1090), .Z(n1092) );
  NAND U2272 ( .A(n1093), .B(n1092), .Z(n1129) );
  XNOR U2273 ( .A(n1129), .B(sreg[228]), .Z(n1131) );
  NAND U2274 ( .A(n1095), .B(n1094), .Z(n36105) );
  OR U2275 ( .A(n1096), .B(n36105), .Z(n1098) );
  XNOR U2276 ( .A(b[3]), .B(a[2]), .Z(n1120) );
  NANDN U2277 ( .A(n1120), .B(n36107), .Z(n1097) );
  AND U2278 ( .A(n1098), .B(n1097), .Z(n1124) );
  NANDN U2279 ( .A(n1049), .B(a[4]), .Z(n1099) );
  XNOR U2280 ( .A(b[1]), .B(n1099), .Z(n1101) );
  NANDN U2281 ( .A(b[0]), .B(a[3]), .Z(n1100) );
  AND U2282 ( .A(n1101), .B(n1100), .Z(n1123) );
  XOR U2283 ( .A(n1124), .B(n1123), .Z(n1126) );
  XNOR U2284 ( .A(b[4]), .B(n1050), .Z(n36587) );
  NANDN U2285 ( .A(n3393), .B(n36587), .Z(n1125) );
  XNOR U2286 ( .A(n1126), .B(n1125), .Z(n1108) );
  XOR U2287 ( .A(n1109), .B(n1110), .Z(n1107) );
  XNOR U2288 ( .A(n1108), .B(n1107), .Z(n1130) );
  XNOR U2289 ( .A(n1131), .B(n1130), .Z(c[228]) );
  NANDN U2290 ( .A(n1049), .B(a[5]), .Z(n1111) );
  XNOR U2291 ( .A(b[1]), .B(n1111), .Z(n1113) );
  NANDN U2292 ( .A(b[0]), .B(a[4]), .Z(n1112) );
  AND U2293 ( .A(n1113), .B(n1112), .Z(n1140) );
  XNOR U2294 ( .A(n1051), .B(a[1]), .Z(n1148) );
  AND U2295 ( .A(n36587), .B(n1148), .Z(n1118) );
  XNOR U2296 ( .A(n1051), .B(a[0]), .Z(n1116) );
  XNOR U2297 ( .A(n1051), .B(b[3]), .Z(n1115) );
  XNOR U2298 ( .A(n1051), .B(b[4]), .Z(n1114) );
  AND U2299 ( .A(n1115), .B(n1114), .Z(n36588) );
  NAND U2300 ( .A(n1116), .B(n36588), .Z(n1117) );
  NANDN U2301 ( .A(n1118), .B(n1117), .Z(n1141) );
  XNOR U2302 ( .A(n1140), .B(n1141), .Z(n1154) );
  NANDN U2303 ( .A(n1050), .B(b[4]), .Z(n1119) );
  ANDN U2304 ( .B(n1119), .A(n1051), .Z(n36861) );
  AND U2305 ( .A(n36861), .B(n1125), .Z(n1152) );
  XNOR U2306 ( .A(b[3]), .B(a[3]), .Z(n1142) );
  NANDN U2307 ( .A(n1142), .B(n36107), .Z(n1122) );
  OR U2308 ( .A(n1120), .B(n36105), .Z(n1121) );
  AND U2309 ( .A(n1122), .B(n1121), .Z(n1151) );
  XNOR U2310 ( .A(n1152), .B(n1151), .Z(n1153) );
  XOR U2311 ( .A(n1154), .B(n1153), .Z(n1135) );
  NANDN U2312 ( .A(n1124), .B(n1123), .Z(n1128) );
  OR U2313 ( .A(n1126), .B(n1125), .Z(n1127) );
  AND U2314 ( .A(n1128), .B(n1127), .Z(n1134) );
  XOR U2315 ( .A(n1135), .B(n1134), .Z(n1136) );
  XNOR U2316 ( .A(n1137), .B(n1136), .Z(n1157) );
  XNOR U2317 ( .A(sreg[229]), .B(n1157), .Z(n1159) );
  NAND U2318 ( .A(n1129), .B(sreg[228]), .Z(n1133) );
  NANDN U2319 ( .A(n1131), .B(n1130), .Z(n1132) );
  AND U2320 ( .A(n1133), .B(n1132), .Z(n1158) );
  XOR U2321 ( .A(n1159), .B(n1158), .Z(c[229]) );
  OR U2322 ( .A(n1135), .B(n1134), .Z(n1139) );
  NANDN U2323 ( .A(n1137), .B(n1136), .Z(n1138) );
  NAND U2324 ( .A(n1139), .B(n1138), .Z(n1165) );
  AND U2325 ( .A(n1141), .B(n1140), .Z(n1189) );
  OR U2326 ( .A(n1142), .B(n36105), .Z(n1144) );
  XNOR U2327 ( .A(b[3]), .B(a[4]), .Z(n1183) );
  NANDN U2328 ( .A(n1183), .B(n36107), .Z(n1143) );
  NAND U2329 ( .A(n1144), .B(n1143), .Z(n1171) );
  NANDN U2330 ( .A(n1049), .B(a[6]), .Z(n1145) );
  XNOR U2331 ( .A(b[1]), .B(n1145), .Z(n1147) );
  NANDN U2332 ( .A(b[0]), .B(a[5]), .Z(n1146) );
  AND U2333 ( .A(n1147), .B(n1146), .Z(n1168) );
  XNOR U2334 ( .A(n1051), .B(b[6]), .Z(n36701) );
  NANDN U2335 ( .A(n3393), .B(n36701), .Z(n1169) );
  XNOR U2336 ( .A(n1168), .B(n1169), .Z(n1170) );
  XNOR U2337 ( .A(n1171), .B(n1170), .Z(n1186) );
  XNOR U2338 ( .A(b[5]), .B(a[2]), .Z(n1172) );
  NANDN U2339 ( .A(n1172), .B(n36587), .Z(n1150) );
  NAND U2340 ( .A(n36588), .B(n1148), .Z(n1149) );
  NAND U2341 ( .A(n1150), .B(n1149), .Z(n1187) );
  XNOR U2342 ( .A(n1186), .B(n1187), .Z(n1188) );
  XOR U2343 ( .A(n1189), .B(n1188), .Z(n1162) );
  NANDN U2344 ( .A(n1152), .B(n1151), .Z(n1156) );
  NAND U2345 ( .A(n1154), .B(n1153), .Z(n1155) );
  NAND U2346 ( .A(n1156), .B(n1155), .Z(n1163) );
  XNOR U2347 ( .A(n1162), .B(n1163), .Z(n1164) );
  XNOR U2348 ( .A(n1165), .B(n1164), .Z(n1194) );
  NAND U2349 ( .A(sreg[229]), .B(n1157), .Z(n1161) );
  OR U2350 ( .A(n1159), .B(n1158), .Z(n1160) );
  NAND U2351 ( .A(n1161), .B(n1160), .Z(n1192) );
  XNOR U2352 ( .A(n1192), .B(sreg[230]), .Z(n1193) );
  XOR U2353 ( .A(n1194), .B(n1193), .Z(c[230]) );
  NANDN U2354 ( .A(n1163), .B(n1162), .Z(n1167) );
  NAND U2355 ( .A(n1165), .B(n1164), .Z(n1166) );
  NAND U2356 ( .A(n1167), .B(n1166), .Z(n1205) );
  XNOR U2357 ( .A(n1051), .B(a[3]), .Z(n1231) );
  NAND U2358 ( .A(n1231), .B(n36587), .Z(n1174) );
  NANDN U2359 ( .A(n1172), .B(n36588), .Z(n1173) );
  NAND U2360 ( .A(n1174), .B(n1173), .Z(n1226) );
  XNOR U2361 ( .A(b[7]), .B(n3393), .Z(n1177) );
  XNOR U2362 ( .A(b[7]), .B(n1051), .Z(n1176) );
  XOR U2363 ( .A(b[7]), .B(b[6]), .Z(n1175) );
  AND U2364 ( .A(n1176), .B(n1175), .Z(n36702) );
  NAND U2365 ( .A(n1177), .B(n36702), .Z(n1179) );
  XOR U2366 ( .A(b[7]), .B(a[1]), .Z(n1220) );
  NAND U2367 ( .A(n1220), .B(n36701), .Z(n1178) );
  NAND U2368 ( .A(n1179), .B(n1178), .Z(n1227) );
  XNOR U2369 ( .A(n1226), .B(n1227), .Z(n1217) );
  NANDN U2370 ( .A(n1049), .B(a[7]), .Z(n1180) );
  XNOR U2371 ( .A(b[1]), .B(n1180), .Z(n1182) );
  IV U2372 ( .A(a[6]), .Z(n4305) );
  NANDN U2373 ( .A(n4305), .B(n1049), .Z(n1181) );
  AND U2374 ( .A(n1182), .B(n1181), .Z(n1215) );
  XNOR U2375 ( .A(n1214), .B(n1215), .Z(n1216) );
  XOR U2376 ( .A(n1217), .B(n1216), .Z(n1208) );
  XNOR U2377 ( .A(b[3]), .B(a[5]), .Z(n1223) );
  NANDN U2378 ( .A(n1223), .B(n36107), .Z(n1185) );
  OR U2379 ( .A(n1183), .B(n36105), .Z(n1184) );
  AND U2380 ( .A(n1185), .B(n1184), .Z(n1209) );
  XNOR U2381 ( .A(n1208), .B(n1209), .Z(n1210) );
  XNOR U2382 ( .A(n1211), .B(n1210), .Z(n1202) );
  NANDN U2383 ( .A(n1187), .B(n1186), .Z(n1191) );
  NANDN U2384 ( .A(n1189), .B(n1188), .Z(n1190) );
  NAND U2385 ( .A(n1191), .B(n1190), .Z(n1203) );
  XNOR U2386 ( .A(n1202), .B(n1203), .Z(n1204) );
  XOR U2387 ( .A(n1205), .B(n1204), .Z(n1197) );
  XNOR U2388 ( .A(sreg[231]), .B(n1197), .Z(n1199) );
  NAND U2389 ( .A(n1192), .B(sreg[230]), .Z(n1196) );
  OR U2390 ( .A(n1194), .B(n1193), .Z(n1195) );
  AND U2391 ( .A(n1196), .B(n1195), .Z(n1198) );
  XOR U2392 ( .A(n1199), .B(n1198), .Z(c[231]) );
  NAND U2393 ( .A(sreg[231]), .B(n1197), .Z(n1201) );
  OR U2394 ( .A(n1199), .B(n1198), .Z(n1200) );
  NAND U2395 ( .A(n1201), .B(n1200), .Z(n1277) );
  XNOR U2396 ( .A(n1277), .B(sreg[232]), .Z(n1279) );
  NANDN U2397 ( .A(n1203), .B(n1202), .Z(n1207) );
  NAND U2398 ( .A(n1205), .B(n1204), .Z(n1206) );
  NAND U2399 ( .A(n1207), .B(n1206), .Z(n1237) );
  NAND U2400 ( .A(n1209), .B(n1208), .Z(n1213) );
  OR U2401 ( .A(n1211), .B(n1210), .Z(n1212) );
  NAND U2402 ( .A(n1213), .B(n1212), .Z(n1234) );
  NANDN U2403 ( .A(n1215), .B(n1214), .Z(n1219) );
  NAND U2404 ( .A(n1217), .B(n1216), .Z(n1218) );
  NAND U2405 ( .A(n1219), .B(n1218), .Z(n1243) );
  XOR U2406 ( .A(b[7]), .B(a[2]), .Z(n1252) );
  NAND U2407 ( .A(n1252), .B(n36701), .Z(n1222) );
  NAND U2408 ( .A(n1220), .B(n36702), .Z(n1221) );
  NAND U2409 ( .A(n1222), .B(n1221), .Z(n1246) );
  OR U2410 ( .A(n1223), .B(n36105), .Z(n1225) );
  XOR U2411 ( .A(b[3]), .B(n4305), .Z(n1268) );
  NANDN U2412 ( .A(n1268), .B(n36107), .Z(n1224) );
  AND U2413 ( .A(n1225), .B(n1224), .Z(n1247) );
  XNOR U2414 ( .A(n1246), .B(n1247), .Z(n1248) );
  NAND U2415 ( .A(n1227), .B(n1226), .Z(n1249) );
  XOR U2416 ( .A(n1248), .B(n1249), .Z(n1240) );
  XOR U2417 ( .A(b[8]), .B(b[7]), .Z(n36925) );
  NAND U2418 ( .A(a[0]), .B(n36925), .Z(n1274) );
  NANDN U2419 ( .A(n1049), .B(a[8]), .Z(n1228) );
  XNOR U2420 ( .A(b[1]), .B(n1228), .Z(n1230) );
  NANDN U2421 ( .A(b[0]), .B(a[7]), .Z(n1229) );
  AND U2422 ( .A(n1230), .B(n1229), .Z(n1272) );
  XNOR U2423 ( .A(b[5]), .B(a[4]), .Z(n1262) );
  NANDN U2424 ( .A(n1262), .B(n36587), .Z(n1233) );
  NAND U2425 ( .A(n36588), .B(n1231), .Z(n1232) );
  AND U2426 ( .A(n1233), .B(n1232), .Z(n1271) );
  XNOR U2427 ( .A(n1272), .B(n1271), .Z(n1273) );
  XNOR U2428 ( .A(n1274), .B(n1273), .Z(n1241) );
  XNOR U2429 ( .A(n1240), .B(n1241), .Z(n1242) );
  XNOR U2430 ( .A(n1243), .B(n1242), .Z(n1235) );
  XNOR U2431 ( .A(n1234), .B(n1235), .Z(n1236) );
  XNOR U2432 ( .A(n1237), .B(n1236), .Z(n1278) );
  XOR U2433 ( .A(n1279), .B(n1278), .Z(c[232]) );
  NANDN U2434 ( .A(n1235), .B(n1234), .Z(n1239) );
  NANDN U2435 ( .A(n1237), .B(n1236), .Z(n1238) );
  NAND U2436 ( .A(n1239), .B(n1238), .Z(n1290) );
  NANDN U2437 ( .A(n1241), .B(n1240), .Z(n1245) );
  NAND U2438 ( .A(n1243), .B(n1242), .Z(n1244) );
  NAND U2439 ( .A(n1245), .B(n1244), .Z(n1287) );
  NANDN U2440 ( .A(n1247), .B(n1246), .Z(n1251) );
  NANDN U2441 ( .A(n1249), .B(n1248), .Z(n1250) );
  NAND U2442 ( .A(n1251), .B(n1250), .Z(n1296) );
  XOR U2443 ( .A(b[7]), .B(a[3]), .Z(n1323) );
  NAND U2444 ( .A(n1323), .B(n36701), .Z(n1254) );
  NAND U2445 ( .A(n1252), .B(n36702), .Z(n1253) );
  NAND U2446 ( .A(n1254), .B(n1253), .Z(n1315) );
  XNOR U2447 ( .A(n1052), .B(a[0]), .Z(n1257) );
  XNOR U2448 ( .A(n1052), .B(b[7]), .Z(n1256) );
  XNOR U2449 ( .A(n1052), .B(b[8]), .Z(n1255) );
  AND U2450 ( .A(n1256), .B(n1255), .Z(n36926) );
  NAND U2451 ( .A(n1257), .B(n36926), .Z(n1259) );
  XNOR U2452 ( .A(b[9]), .B(a[1]), .Z(n1312) );
  ANDN U2453 ( .B(n36925), .A(n1312), .Z(n1258) );
  ANDN U2454 ( .B(n1259), .A(n1258), .Z(n1316) );
  XOR U2455 ( .A(n1315), .B(n1316), .Z(n1301) );
  NAND U2456 ( .A(b[8]), .B(b[7]), .Z(n37183) );
  ANDN U2457 ( .B(n37183), .A(n1052), .Z(n1261) );
  NANDN U2458 ( .A(n3393), .B(n36925), .Z(n1260) );
  AND U2459 ( .A(n1261), .B(n1260), .Z(n1299) );
  XNOR U2460 ( .A(b[5]), .B(a[5]), .Z(n1309) );
  NANDN U2461 ( .A(n1309), .B(n36587), .Z(n1264) );
  NANDN U2462 ( .A(n1262), .B(n36588), .Z(n1263) );
  NAND U2463 ( .A(n1264), .B(n1263), .Z(n1300) );
  XNOR U2464 ( .A(n1299), .B(n1300), .Z(n1302) );
  XNOR U2465 ( .A(n1301), .B(n1302), .Z(n1308) );
  NANDN U2466 ( .A(n1049), .B(a[9]), .Z(n1265) );
  XNOR U2467 ( .A(b[1]), .B(n1265), .Z(n1267) );
  NANDN U2468 ( .A(b[0]), .B(a[8]), .Z(n1266) );
  AND U2469 ( .A(n1267), .B(n1266), .Z(n1305) );
  OR U2470 ( .A(n1268), .B(n36105), .Z(n1270) );
  XNOR U2471 ( .A(b[3]), .B(a[7]), .Z(n1317) );
  NANDN U2472 ( .A(n1317), .B(n36107), .Z(n1269) );
  AND U2473 ( .A(n1270), .B(n1269), .Z(n1306) );
  XNOR U2474 ( .A(n1305), .B(n1306), .Z(n1307) );
  XNOR U2475 ( .A(n1308), .B(n1307), .Z(n1293) );
  NANDN U2476 ( .A(n1272), .B(n1271), .Z(n1276) );
  NAND U2477 ( .A(n1274), .B(n1273), .Z(n1275) );
  AND U2478 ( .A(n1276), .B(n1275), .Z(n1294) );
  XOR U2479 ( .A(n1293), .B(n1294), .Z(n1295) );
  XOR U2480 ( .A(n1296), .B(n1295), .Z(n1288) );
  XNOR U2481 ( .A(n1287), .B(n1288), .Z(n1289) );
  XNOR U2482 ( .A(n1290), .B(n1289), .Z(n1282) );
  XNOR U2483 ( .A(n1282), .B(sreg[233]), .Z(n1284) );
  NAND U2484 ( .A(n1277), .B(sreg[232]), .Z(n1281) );
  OR U2485 ( .A(n1279), .B(n1278), .Z(n1280) );
  AND U2486 ( .A(n1281), .B(n1280), .Z(n1283) );
  XOR U2487 ( .A(n1284), .B(n1283), .Z(c[233]) );
  NAND U2488 ( .A(n1282), .B(sreg[233]), .Z(n1286) );
  OR U2489 ( .A(n1284), .B(n1283), .Z(n1285) );
  NAND U2490 ( .A(n1286), .B(n1285), .Z(n1374) );
  XNOR U2491 ( .A(n1374), .B(sreg[234]), .Z(n1376) );
  NANDN U2492 ( .A(n1288), .B(n1287), .Z(n1292) );
  NAND U2493 ( .A(n1290), .B(n1289), .Z(n1291) );
  NAND U2494 ( .A(n1292), .B(n1291), .Z(n1329) );
  NAND U2495 ( .A(n1294), .B(n1293), .Z(n1298) );
  NAND U2496 ( .A(n1296), .B(n1295), .Z(n1297) );
  NAND U2497 ( .A(n1298), .B(n1297), .Z(n1326) );
  OR U2498 ( .A(n1300), .B(n1299), .Z(n1304) );
  NANDN U2499 ( .A(n1302), .B(n1301), .Z(n1303) );
  NAND U2500 ( .A(n1304), .B(n1303), .Z(n1335) );
  XOR U2501 ( .A(n1051), .B(n4305), .Z(n1371) );
  NAND U2502 ( .A(n1371), .B(n36587), .Z(n1311) );
  NANDN U2503 ( .A(n1309), .B(n36588), .Z(n1310) );
  NAND U2504 ( .A(n1311), .B(n1310), .Z(n1348) );
  XNOR U2505 ( .A(b[9]), .B(a[2]), .Z(n1360) );
  NANDN U2506 ( .A(n1360), .B(n36925), .Z(n1314) );
  NANDN U2507 ( .A(n1312), .B(n36926), .Z(n1313) );
  AND U2508 ( .A(n1314), .B(n1313), .Z(n1349) );
  XNOR U2509 ( .A(n1348), .B(n1349), .Z(n1350) );
  NANDN U2510 ( .A(n1316), .B(n1315), .Z(n1351) );
  XOR U2511 ( .A(n1350), .B(n1351), .Z(n1336) );
  XNOR U2512 ( .A(b[3]), .B(a[8]), .Z(n1354) );
  NANDN U2513 ( .A(n1354), .B(n36107), .Z(n1319) );
  OR U2514 ( .A(n1317), .B(n36105), .Z(n1318) );
  NAND U2515 ( .A(n1319), .B(n1318), .Z(n1337) );
  XNOR U2516 ( .A(n1336), .B(n1337), .Z(n1338) );
  XOR U2517 ( .A(n1052), .B(b[10]), .Z(n37311) );
  NOR U2518 ( .A(n3393), .B(n37311), .Z(n1345) );
  NANDN U2519 ( .A(n1049), .B(a[10]), .Z(n1320) );
  XNOR U2520 ( .A(b[1]), .B(n1320), .Z(n1322) );
  NANDN U2521 ( .A(b[0]), .B(a[9]), .Z(n1321) );
  AND U2522 ( .A(n1322), .B(n1321), .Z(n1343) );
  XNOR U2523 ( .A(b[7]), .B(a[4]), .Z(n1357) );
  NANDN U2524 ( .A(n1357), .B(n36701), .Z(n1325) );
  NAND U2525 ( .A(n36702), .B(n1323), .Z(n1324) );
  AND U2526 ( .A(n1325), .B(n1324), .Z(n1342) );
  XNOR U2527 ( .A(n1343), .B(n1342), .Z(n1344) );
  XOR U2528 ( .A(n1345), .B(n1344), .Z(n1339) );
  XNOR U2529 ( .A(n1338), .B(n1339), .Z(n1332) );
  XNOR U2530 ( .A(n1333), .B(n1332), .Z(n1334) );
  XNOR U2531 ( .A(n1335), .B(n1334), .Z(n1327) );
  XOR U2532 ( .A(n1326), .B(n1327), .Z(n1328) );
  XOR U2533 ( .A(n1329), .B(n1328), .Z(n1375) );
  XOR U2534 ( .A(n1376), .B(n1375), .Z(c[234]) );
  OR U2535 ( .A(n1327), .B(n1326), .Z(n1331) );
  NAND U2536 ( .A(n1329), .B(n1328), .Z(n1330) );
  NAND U2537 ( .A(n1331), .B(n1330), .Z(n1387) );
  NANDN U2538 ( .A(n1337), .B(n1336), .Z(n1341) );
  NANDN U2539 ( .A(n1339), .B(n1338), .Z(n1340) );
  NAND U2540 ( .A(n1341), .B(n1340), .Z(n1393) );
  NANDN U2541 ( .A(n1343), .B(n1342), .Z(n1347) );
  NANDN U2542 ( .A(n1345), .B(n1344), .Z(n1346) );
  NAND U2543 ( .A(n1347), .B(n1346), .Z(n1390) );
  NANDN U2544 ( .A(n1349), .B(n1348), .Z(n1353) );
  NANDN U2545 ( .A(n1351), .B(n1350), .Z(n1352) );
  NAND U2546 ( .A(n1353), .B(n1352), .Z(n1431) );
  XNOR U2547 ( .A(b[3]), .B(a[9]), .Z(n1413) );
  NANDN U2548 ( .A(n1413), .B(n36107), .Z(n1356) );
  OR U2549 ( .A(n1354), .B(n36105), .Z(n1355) );
  NAND U2550 ( .A(n1356), .B(n1355), .Z(n1397) );
  XOR U2551 ( .A(n1396), .B(n1397), .Z(n1399) );
  XNOR U2552 ( .A(b[7]), .B(a[5]), .Z(n1410) );
  NANDN U2553 ( .A(n1410), .B(n36701), .Z(n1359) );
  NANDN U2554 ( .A(n1357), .B(n36702), .Z(n1358) );
  NAND U2555 ( .A(n1359), .B(n1358), .Z(n1398) );
  XNOR U2556 ( .A(n1399), .B(n1398), .Z(n1428) );
  XNOR U2557 ( .A(n1052), .B(a[3]), .Z(n1419) );
  NAND U2558 ( .A(n36925), .B(n1419), .Z(n1362) );
  NANDN U2559 ( .A(n1360), .B(n36926), .Z(n1361) );
  NAND U2560 ( .A(n1362), .B(n1361), .Z(n1409) );
  XOR U2561 ( .A(b[11]), .B(a[1]), .Z(n1405) );
  ANDN U2562 ( .B(n1405), .A(n37311), .Z(n1367) );
  XNOR U2563 ( .A(b[11]), .B(n3393), .Z(n1365) );
  XNOR U2564 ( .A(b[11]), .B(n1052), .Z(n1364) );
  XOR U2565 ( .A(b[11]), .B(b[10]), .Z(n1363) );
  AND U2566 ( .A(n1364), .B(n1363), .Z(n37218) );
  NAND U2567 ( .A(n1365), .B(n37218), .Z(n1366) );
  NANDN U2568 ( .A(n1367), .B(n1366), .Z(n1408) );
  XNOR U2569 ( .A(n1409), .B(n1408), .Z(n1425) );
  NANDN U2570 ( .A(n1049), .B(a[11]), .Z(n1368) );
  XNOR U2571 ( .A(b[1]), .B(n1368), .Z(n1370) );
  NANDN U2572 ( .A(b[0]), .B(a[10]), .Z(n1369) );
  AND U2573 ( .A(n1370), .B(n1369), .Z(n1423) );
  XOR U2574 ( .A(n1051), .B(a[7]), .Z(n1402) );
  NANDN U2575 ( .A(n1402), .B(n36587), .Z(n1373) );
  NAND U2576 ( .A(n36588), .B(n1371), .Z(n1372) );
  AND U2577 ( .A(n1373), .B(n1372), .Z(n1422) );
  XNOR U2578 ( .A(n1423), .B(n1422), .Z(n1424) );
  XOR U2579 ( .A(n1425), .B(n1424), .Z(n1429) );
  XNOR U2580 ( .A(n1428), .B(n1429), .Z(n1430) );
  XOR U2581 ( .A(n1431), .B(n1430), .Z(n1391) );
  XNOR U2582 ( .A(n1390), .B(n1391), .Z(n1392) );
  XNOR U2583 ( .A(n1393), .B(n1392), .Z(n1385) );
  XNOR U2584 ( .A(n1384), .B(n1385), .Z(n1386) );
  XNOR U2585 ( .A(n1387), .B(n1386), .Z(n1379) );
  XNOR U2586 ( .A(n1379), .B(sreg[235]), .Z(n1381) );
  NAND U2587 ( .A(n1374), .B(sreg[234]), .Z(n1378) );
  OR U2588 ( .A(n1376), .B(n1375), .Z(n1377) );
  AND U2589 ( .A(n1378), .B(n1377), .Z(n1380) );
  XOR U2590 ( .A(n1381), .B(n1380), .Z(c[235]) );
  NAND U2591 ( .A(n1379), .B(sreg[235]), .Z(n1383) );
  OR U2592 ( .A(n1381), .B(n1380), .Z(n1382) );
  NAND U2593 ( .A(n1383), .B(n1382), .Z(n1493) );
  XNOR U2594 ( .A(n1493), .B(sreg[236]), .Z(n1495) );
  NANDN U2595 ( .A(n1385), .B(n1384), .Z(n1389) );
  NAND U2596 ( .A(n1387), .B(n1386), .Z(n1388) );
  NAND U2597 ( .A(n1389), .B(n1388), .Z(n1437) );
  NANDN U2598 ( .A(n1391), .B(n1390), .Z(n1395) );
  NAND U2599 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U2600 ( .A(n1395), .B(n1394), .Z(n1434) );
  NANDN U2601 ( .A(n1397), .B(n1396), .Z(n1401) );
  OR U2602 ( .A(n1399), .B(n1398), .Z(n1400) );
  NAND U2603 ( .A(n1401), .B(n1400), .Z(n1443) );
  XOR U2604 ( .A(n1051), .B(a[8]), .Z(n1476) );
  NANDN U2605 ( .A(n1476), .B(n36587), .Z(n1404) );
  NANDN U2606 ( .A(n1402), .B(n36588), .Z(n1403) );
  NAND U2607 ( .A(n1404), .B(n1403), .Z(n1453) );
  XOR U2608 ( .A(b[11]), .B(a[2]), .Z(n1479) );
  NANDN U2609 ( .A(n37311), .B(n1479), .Z(n1407) );
  NAND U2610 ( .A(n37218), .B(n1405), .Z(n1406) );
  AND U2611 ( .A(n1407), .B(n1406), .Z(n1452) );
  XNOR U2612 ( .A(n1453), .B(n1452), .Z(n1454) );
  NAND U2613 ( .A(n1409), .B(n1408), .Z(n1461) );
  XOR U2614 ( .A(b[7]), .B(n4305), .Z(n1490) );
  NANDN U2615 ( .A(n1490), .B(n36701), .Z(n1412) );
  NANDN U2616 ( .A(n1410), .B(n36702), .Z(n1411) );
  NAND U2617 ( .A(n1412), .B(n1411), .Z(n1459) );
  XNOR U2618 ( .A(b[3]), .B(a[10]), .Z(n1470) );
  NANDN U2619 ( .A(n1470), .B(n36107), .Z(n1415) );
  OR U2620 ( .A(n1413), .B(n36105), .Z(n1414) );
  AND U2621 ( .A(n1415), .B(n1414), .Z(n1458) );
  XNOR U2622 ( .A(n1459), .B(n1458), .Z(n1460) );
  XNOR U2623 ( .A(n1461), .B(n1460), .Z(n1455) );
  XOR U2624 ( .A(n1454), .B(n1455), .Z(n1449) );
  NANDN U2625 ( .A(n1049), .B(a[12]), .Z(n1416) );
  XNOR U2626 ( .A(b[1]), .B(n1416), .Z(n1418) );
  NANDN U2627 ( .A(b[0]), .B(a[11]), .Z(n1417) );
  AND U2628 ( .A(n1418), .B(n1417), .Z(n1464) );
  XNOR U2629 ( .A(b[9]), .B(a[4]), .Z(n1473) );
  NANDN U2630 ( .A(n1473), .B(n36925), .Z(n1421) );
  NAND U2631 ( .A(n1419), .B(n36926), .Z(n1420) );
  AND U2632 ( .A(n1421), .B(n1420), .Z(n1465) );
  XOR U2633 ( .A(n1464), .B(n1465), .Z(n1467) );
  XOR U2634 ( .A(b[11]), .B(b[12]), .Z(n37424) );
  NANDN U2635 ( .A(n3393), .B(n37424), .Z(n1466) );
  XOR U2636 ( .A(n1467), .B(n1466), .Z(n1446) );
  NANDN U2637 ( .A(n1423), .B(n1422), .Z(n1427) );
  NAND U2638 ( .A(n1425), .B(n1424), .Z(n1426) );
  AND U2639 ( .A(n1427), .B(n1426), .Z(n1447) );
  XOR U2640 ( .A(n1446), .B(n1447), .Z(n1448) );
  XNOR U2641 ( .A(n1449), .B(n1448), .Z(n1440) );
  NANDN U2642 ( .A(n1429), .B(n1428), .Z(n1433) );
  NAND U2643 ( .A(n1431), .B(n1430), .Z(n1432) );
  NAND U2644 ( .A(n1433), .B(n1432), .Z(n1441) );
  XNOR U2645 ( .A(n1440), .B(n1441), .Z(n1442) );
  XNOR U2646 ( .A(n1443), .B(n1442), .Z(n1435) );
  XNOR U2647 ( .A(n1434), .B(n1435), .Z(n1436) );
  XOR U2648 ( .A(n1437), .B(n1436), .Z(n1494) );
  XOR U2649 ( .A(n1495), .B(n1494), .Z(c[236]) );
  NANDN U2650 ( .A(n1435), .B(n1434), .Z(n1439) );
  NAND U2651 ( .A(n1437), .B(n1436), .Z(n1438) );
  NAND U2652 ( .A(n1439), .B(n1438), .Z(n1506) );
  NANDN U2653 ( .A(n1441), .B(n1440), .Z(n1445) );
  NAND U2654 ( .A(n1443), .B(n1442), .Z(n1444) );
  NAND U2655 ( .A(n1445), .B(n1444), .Z(n1504) );
  NAND U2656 ( .A(n1447), .B(n1446), .Z(n1451) );
  NAND U2657 ( .A(n1449), .B(n1448), .Z(n1450) );
  NAND U2658 ( .A(n1451), .B(n1450), .Z(n1510) );
  NANDN U2659 ( .A(n1453), .B(n1452), .Z(n1457) );
  NANDN U2660 ( .A(n1455), .B(n1454), .Z(n1456) );
  NAND U2661 ( .A(n1457), .B(n1456), .Z(n1508) );
  NANDN U2662 ( .A(n1459), .B(n1458), .Z(n1463) );
  NAND U2663 ( .A(n1461), .B(n1460), .Z(n1462) );
  NAND U2664 ( .A(n1463), .B(n1462), .Z(n1548) );
  NANDN U2665 ( .A(n1465), .B(n1464), .Z(n1469) );
  OR U2666 ( .A(n1467), .B(n1466), .Z(n1468) );
  NAND U2667 ( .A(n1469), .B(n1468), .Z(n1549) );
  XNOR U2668 ( .A(n1548), .B(n1549), .Z(n1550) );
  OR U2669 ( .A(n1470), .B(n36105), .Z(n1472) );
  XNOR U2670 ( .A(b[3]), .B(a[11]), .Z(n1539) );
  NANDN U2671 ( .A(n1539), .B(n36107), .Z(n1471) );
  NAND U2672 ( .A(n1472), .B(n1471), .Z(n1521) );
  XNOR U2673 ( .A(b[9]), .B(a[5]), .Z(n1516) );
  NANDN U2674 ( .A(n1516), .B(n36925), .Z(n1475) );
  NANDN U2675 ( .A(n1473), .B(n36926), .Z(n1474) );
  AND U2676 ( .A(n1475), .B(n1474), .Z(n1522) );
  XNOR U2677 ( .A(n1521), .B(n1522), .Z(n1523) );
  XNOR U2678 ( .A(n1524), .B(n1523), .Z(n1554) );
  XNOR U2679 ( .A(b[5]), .B(a[9]), .Z(n1533) );
  NANDN U2680 ( .A(n1533), .B(n36587), .Z(n1478) );
  NANDN U2681 ( .A(n1476), .B(n36588), .Z(n1477) );
  NAND U2682 ( .A(n1478), .B(n1477), .Z(n1555) );
  XNOR U2683 ( .A(n1554), .B(n1555), .Z(n1557) );
  XOR U2684 ( .A(b[11]), .B(a[3]), .Z(n1530) );
  NANDN U2685 ( .A(n37311), .B(n1530), .Z(n1481) );
  NAND U2686 ( .A(n1479), .B(n37218), .Z(n1480) );
  NAND U2687 ( .A(n1481), .B(n1480), .Z(n1519) );
  XNOR U2688 ( .A(n1053), .B(a[0]), .Z(n1484) );
  XNOR U2689 ( .A(n1053), .B(b[11]), .Z(n1483) );
  XNOR U2690 ( .A(n1053), .B(b[12]), .Z(n1482) );
  AND U2691 ( .A(n1483), .B(n1482), .Z(n37425) );
  NAND U2692 ( .A(n1484), .B(n37425), .Z(n1486) );
  XNOR U2693 ( .A(n1053), .B(a[1]), .Z(n1513) );
  NAND U2694 ( .A(n1513), .B(n37424), .Z(n1485) );
  NAND U2695 ( .A(n1486), .B(n1485), .Z(n1520) );
  XNOR U2696 ( .A(n1519), .B(n1520), .Z(n1545) );
  NANDN U2697 ( .A(n1049), .B(a[13]), .Z(n1487) );
  XNOR U2698 ( .A(b[1]), .B(n1487), .Z(n1489) );
  NANDN U2699 ( .A(b[0]), .B(a[12]), .Z(n1488) );
  AND U2700 ( .A(n1489), .B(n1488), .Z(n1543) );
  XOR U2701 ( .A(b[7]), .B(a[7]), .Z(n1536) );
  NAND U2702 ( .A(n36701), .B(n1536), .Z(n1492) );
  NANDN U2703 ( .A(n1490), .B(n36702), .Z(n1491) );
  AND U2704 ( .A(n1492), .B(n1491), .Z(n1542) );
  XNOR U2705 ( .A(n1543), .B(n1542), .Z(n1544) );
  XOR U2706 ( .A(n1545), .B(n1544), .Z(n1556) );
  XNOR U2707 ( .A(n1557), .B(n1556), .Z(n1551) );
  XOR U2708 ( .A(n1550), .B(n1551), .Z(n1507) );
  XOR U2709 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U2710 ( .A(n1510), .B(n1509), .Z(n1503) );
  XOR U2711 ( .A(n1504), .B(n1503), .Z(n1505) );
  XNOR U2712 ( .A(n1506), .B(n1505), .Z(n1498) );
  XNOR U2713 ( .A(n1498), .B(sreg[237]), .Z(n1500) );
  NAND U2714 ( .A(n1493), .B(sreg[236]), .Z(n1497) );
  OR U2715 ( .A(n1495), .B(n1494), .Z(n1496) );
  AND U2716 ( .A(n1497), .B(n1496), .Z(n1499) );
  XOR U2717 ( .A(n1500), .B(n1499), .Z(c[237]) );
  NAND U2718 ( .A(n1498), .B(sreg[237]), .Z(n1502) );
  OR U2719 ( .A(n1500), .B(n1499), .Z(n1501) );
  NAND U2720 ( .A(n1502), .B(n1501), .Z(n1626) );
  XNOR U2721 ( .A(n1626), .B(sreg[238]), .Z(n1628) );
  NAND U2722 ( .A(n1508), .B(n1507), .Z(n1512) );
  NANDN U2723 ( .A(n1510), .B(n1509), .Z(n1511) );
  NAND U2724 ( .A(n1512), .B(n1511), .Z(n1560) );
  XNOR U2725 ( .A(b[13]), .B(a[2]), .Z(n1582) );
  NANDN U2726 ( .A(n1582), .B(n37424), .Z(n1515) );
  NAND U2727 ( .A(n1513), .B(n37425), .Z(n1514) );
  NAND U2728 ( .A(n1515), .B(n1514), .Z(n1620) );
  XOR U2729 ( .A(b[9]), .B(n4305), .Z(n1579) );
  NANDN U2730 ( .A(n1579), .B(n36925), .Z(n1518) );
  NANDN U2731 ( .A(n1516), .B(n36926), .Z(n1517) );
  AND U2732 ( .A(n1518), .B(n1517), .Z(n1621) );
  XNOR U2733 ( .A(n1620), .B(n1621), .Z(n1622) );
  NAND U2734 ( .A(n1520), .B(n1519), .Z(n1623) );
  XOR U2735 ( .A(n1622), .B(n1623), .Z(n1575) );
  NANDN U2736 ( .A(n1522), .B(n1521), .Z(n1526) );
  NANDN U2737 ( .A(n1524), .B(n1523), .Z(n1525) );
  NAND U2738 ( .A(n1526), .B(n1525), .Z(n1613) );
  XOR U2739 ( .A(n1053), .B(b[14]), .Z(n37665) );
  NOR U2740 ( .A(n3393), .B(n37665), .Z(n1617) );
  NANDN U2741 ( .A(n1049), .B(a[14]), .Z(n1527) );
  XNOR U2742 ( .A(b[1]), .B(n1527), .Z(n1529) );
  NANDN U2743 ( .A(b[0]), .B(a[13]), .Z(n1528) );
  AND U2744 ( .A(n1529), .B(n1528), .Z(n1615) );
  XOR U2745 ( .A(b[11]), .B(a[4]), .Z(n1596) );
  NANDN U2746 ( .A(n37311), .B(n1596), .Z(n1532) );
  NAND U2747 ( .A(n37218), .B(n1530), .Z(n1531) );
  AND U2748 ( .A(n1532), .B(n1531), .Z(n1614) );
  XNOR U2749 ( .A(n1615), .B(n1614), .Z(n1616) );
  XOR U2750 ( .A(n1617), .B(n1616), .Z(n1610) );
  XNOR U2751 ( .A(b[5]), .B(a[10]), .Z(n1599) );
  NANDN U2752 ( .A(n1599), .B(n36587), .Z(n1535) );
  NANDN U2753 ( .A(n1533), .B(n36588), .Z(n1534) );
  NAND U2754 ( .A(n1535), .B(n1534), .Z(n1593) );
  XOR U2755 ( .A(b[7]), .B(a[8]), .Z(n1607) );
  NAND U2756 ( .A(n1607), .B(n36701), .Z(n1538) );
  NAND U2757 ( .A(n1536), .B(n36702), .Z(n1537) );
  NAND U2758 ( .A(n1538), .B(n1537), .Z(n1590) );
  OR U2759 ( .A(n1539), .B(n36105), .Z(n1541) );
  XNOR U2760 ( .A(b[3]), .B(a[12]), .Z(n1602) );
  NANDN U2761 ( .A(n1602), .B(n36107), .Z(n1540) );
  AND U2762 ( .A(n1541), .B(n1540), .Z(n1591) );
  XNOR U2763 ( .A(n1590), .B(n1591), .Z(n1592) );
  XNOR U2764 ( .A(n1593), .B(n1592), .Z(n1611) );
  XNOR U2765 ( .A(n1610), .B(n1611), .Z(n1612) );
  XNOR U2766 ( .A(n1613), .B(n1612), .Z(n1572) );
  NANDN U2767 ( .A(n1543), .B(n1542), .Z(n1547) );
  NAND U2768 ( .A(n1545), .B(n1544), .Z(n1546) );
  AND U2769 ( .A(n1547), .B(n1546), .Z(n1573) );
  XNOR U2770 ( .A(n1572), .B(n1573), .Z(n1574) );
  XNOR U2771 ( .A(n1575), .B(n1574), .Z(n1569) );
  NANDN U2772 ( .A(n1549), .B(n1548), .Z(n1553) );
  NAND U2773 ( .A(n1551), .B(n1550), .Z(n1552) );
  NAND U2774 ( .A(n1553), .B(n1552), .Z(n1567) );
  OR U2775 ( .A(n1555), .B(n1554), .Z(n1559) );
  NANDN U2776 ( .A(n1557), .B(n1556), .Z(n1558) );
  AND U2777 ( .A(n1559), .B(n1558), .Z(n1566) );
  XNOR U2778 ( .A(n1567), .B(n1566), .Z(n1568) );
  XOR U2779 ( .A(n1569), .B(n1568), .Z(n1561) );
  XNOR U2780 ( .A(n1560), .B(n1561), .Z(n1562) );
  XOR U2781 ( .A(n1563), .B(n1562), .Z(n1627) );
  XOR U2782 ( .A(n1628), .B(n1627), .Z(c[238]) );
  NANDN U2783 ( .A(n1561), .B(n1560), .Z(n1565) );
  NAND U2784 ( .A(n1563), .B(n1562), .Z(n1564) );
  NAND U2785 ( .A(n1565), .B(n1564), .Z(n1639) );
  NANDN U2786 ( .A(n1567), .B(n1566), .Z(n1571) );
  NAND U2787 ( .A(n1569), .B(n1568), .Z(n1570) );
  NAND U2788 ( .A(n1571), .B(n1570), .Z(n1637) );
  NANDN U2789 ( .A(n1049), .B(a[15]), .Z(n1576) );
  XNOR U2790 ( .A(b[1]), .B(n1576), .Z(n1578) );
  NANDN U2791 ( .A(b[0]), .B(a[14]), .Z(n1577) );
  AND U2792 ( .A(n1578), .B(n1577), .Z(n1664) );
  XNOR U2793 ( .A(n1052), .B(a[7]), .Z(n1676) );
  NAND U2794 ( .A(n36925), .B(n1676), .Z(n1581) );
  NANDN U2795 ( .A(n1579), .B(n36926), .Z(n1580) );
  AND U2796 ( .A(n1581), .B(n1580), .Z(n1665) );
  XNOR U2797 ( .A(n1664), .B(n1665), .Z(n1666) );
  XNOR U2798 ( .A(b[13]), .B(a[3]), .Z(n1661) );
  NANDN U2799 ( .A(n1661), .B(n37424), .Z(n1584) );
  NANDN U2800 ( .A(n1582), .B(n37425), .Z(n1583) );
  NAND U2801 ( .A(n1584), .B(n1583), .Z(n1674) );
  XOR U2802 ( .A(b[15]), .B(a[0]), .Z(n1587) );
  XNOR U2803 ( .A(n1054), .B(b[13]), .Z(n1586) );
  XNOR U2804 ( .A(n1054), .B(b[14]), .Z(n1585) );
  AND U2805 ( .A(n1586), .B(n1585), .Z(n37604) );
  NAND U2806 ( .A(n1587), .B(n37604), .Z(n1589) );
  XNOR U2807 ( .A(n1054), .B(a[1]), .Z(n1688) );
  ANDN U2808 ( .B(n1688), .A(n37665), .Z(n1588) );
  ANDN U2809 ( .B(n1589), .A(n1588), .Z(n1675) );
  XNOR U2810 ( .A(n1674), .B(n1675), .Z(n1667) );
  XOR U2811 ( .A(n1666), .B(n1667), .Z(n1694) );
  NANDN U2812 ( .A(n1591), .B(n1590), .Z(n1595) );
  NAND U2813 ( .A(n1593), .B(n1592), .Z(n1594) );
  NAND U2814 ( .A(n1595), .B(n1594), .Z(n1695) );
  XOR U2815 ( .A(n1694), .B(n1695), .Z(n1696) );
  XOR U2816 ( .A(b[11]), .B(a[5]), .Z(n1685) );
  NANDN U2817 ( .A(n37311), .B(n1685), .Z(n1598) );
  NAND U2818 ( .A(n1596), .B(n37218), .Z(n1597) );
  NAND U2819 ( .A(n1598), .B(n1597), .Z(n1655) );
  XNOR U2820 ( .A(b[5]), .B(a[11]), .Z(n1691) );
  NANDN U2821 ( .A(n1691), .B(n36587), .Z(n1601) );
  NANDN U2822 ( .A(n1599), .B(n36588), .Z(n1600) );
  NAND U2823 ( .A(n1601), .B(n1600), .Z(n1652) );
  OR U2824 ( .A(n1602), .B(n36105), .Z(n1604) );
  XNOR U2825 ( .A(b[3]), .B(a[13]), .Z(n1679) );
  NANDN U2826 ( .A(n1679), .B(n36107), .Z(n1603) );
  AND U2827 ( .A(n1604), .B(n1603), .Z(n1653) );
  XNOR U2828 ( .A(n1652), .B(n1653), .Z(n1654) );
  XNOR U2829 ( .A(n1655), .B(n1654), .Z(n1671) );
  NOR U2830 ( .A(b[13]), .B(b[14]), .Z(n1605) );
  OR U2831 ( .A(n1605), .B(n3393), .Z(n1606) );
  NANDN U2832 ( .A(n1053), .B(b[14]), .Z(n37663) );
  AND U2833 ( .A(n37663), .B(b[15]), .Z(n37851) );
  AND U2834 ( .A(n1606), .B(n37851), .Z(n1669) );
  XOR U2835 ( .A(b[7]), .B(a[9]), .Z(n1682) );
  NAND U2836 ( .A(n36701), .B(n1682), .Z(n1609) );
  NAND U2837 ( .A(n36702), .B(n1607), .Z(n1608) );
  NAND U2838 ( .A(n1609), .B(n1608), .Z(n1668) );
  XOR U2839 ( .A(n1669), .B(n1668), .Z(n1670) );
  XOR U2840 ( .A(n1671), .B(n1670), .Z(n1697) );
  XOR U2841 ( .A(n1696), .B(n1697), .Z(n1640) );
  XNOR U2842 ( .A(n1641), .B(n1640), .Z(n1642) );
  NANDN U2843 ( .A(n1615), .B(n1614), .Z(n1619) );
  NANDN U2844 ( .A(n1617), .B(n1616), .Z(n1618) );
  NAND U2845 ( .A(n1619), .B(n1618), .Z(n1646) );
  NANDN U2846 ( .A(n1621), .B(n1620), .Z(n1625) );
  NANDN U2847 ( .A(n1623), .B(n1622), .Z(n1624) );
  NAND U2848 ( .A(n1625), .B(n1624), .Z(n1647) );
  XNOR U2849 ( .A(n1646), .B(n1647), .Z(n1648) );
  XOR U2850 ( .A(n1649), .B(n1648), .Z(n1643) );
  XOR U2851 ( .A(n1642), .B(n1643), .Z(n1636) );
  XNOR U2852 ( .A(n1637), .B(n1636), .Z(n1638) );
  XNOR U2853 ( .A(n1639), .B(n1638), .Z(n1631) );
  XNOR U2854 ( .A(n1631), .B(sreg[239]), .Z(n1633) );
  NAND U2855 ( .A(n1626), .B(sreg[238]), .Z(n1630) );
  OR U2856 ( .A(n1628), .B(n1627), .Z(n1629) );
  AND U2857 ( .A(n1630), .B(n1629), .Z(n1632) );
  XOR U2858 ( .A(n1633), .B(n1632), .Z(c[239]) );
  NAND U2859 ( .A(n1631), .B(sreg[239]), .Z(n1635) );
  OR U2860 ( .A(n1633), .B(n1632), .Z(n1634) );
  NAND U2861 ( .A(n1635), .B(n1634), .Z(n1775) );
  XNOR U2862 ( .A(n1775), .B(sreg[240]), .Z(n1777) );
  NAND U2863 ( .A(n1641), .B(n1640), .Z(n1645) );
  OR U2864 ( .A(n1643), .B(n1642), .Z(n1644) );
  NAND U2865 ( .A(n1645), .B(n1644), .Z(n1700) );
  NANDN U2866 ( .A(n1647), .B(n1646), .Z(n1651) );
  NANDN U2867 ( .A(n1649), .B(n1648), .Z(n1650) );
  NAND U2868 ( .A(n1651), .B(n1650), .Z(n1774) );
  NANDN U2869 ( .A(n1653), .B(n1652), .Z(n1657) );
  NAND U2870 ( .A(n1655), .B(n1654), .Z(n1656) );
  NAND U2871 ( .A(n1657), .B(n1656), .Z(n1715) );
  NANDN U2872 ( .A(n1049), .B(a[16]), .Z(n1658) );
  XNOR U2873 ( .A(b[1]), .B(n1658), .Z(n1660) );
  NANDN U2874 ( .A(b[0]), .B(a[15]), .Z(n1659) );
  AND U2875 ( .A(n1660), .B(n1659), .Z(n1745) );
  XNOR U2876 ( .A(b[13]), .B(a[4]), .Z(n1728) );
  NANDN U2877 ( .A(n1728), .B(n37424), .Z(n1663) );
  NANDN U2878 ( .A(n1661), .B(n37425), .Z(n1662) );
  NAND U2879 ( .A(n1663), .B(n1662), .Z(n1743) );
  XOR U2880 ( .A(b[15]), .B(b[16]), .Z(n37764) );
  NANDN U2881 ( .A(n3393), .B(n37764), .Z(n1744) );
  XNOR U2882 ( .A(n1743), .B(n1744), .Z(n1746) );
  XOR U2883 ( .A(n1745), .B(n1746), .Z(n1712) );
  XOR U2884 ( .A(n1712), .B(n1713), .Z(n1714) );
  XOR U2885 ( .A(n1715), .B(n1714), .Z(n1706) );
  OR U2886 ( .A(n1669), .B(n1668), .Z(n1673) );
  NAND U2887 ( .A(n1671), .B(n1670), .Z(n1672) );
  NAND U2888 ( .A(n1673), .B(n1672), .Z(n1707) );
  XNOR U2889 ( .A(n1706), .B(n1707), .Z(n1708) );
  NANDN U2890 ( .A(n1675), .B(n1674), .Z(n1720) );
  XOR U2891 ( .A(n1052), .B(a[8]), .Z(n1759) );
  NANDN U2892 ( .A(n1759), .B(n36925), .Z(n1678) );
  NAND U2893 ( .A(n36926), .B(n1676), .Z(n1677) );
  NAND U2894 ( .A(n1678), .B(n1677), .Z(n1719) );
  XNOR U2895 ( .A(b[3]), .B(a[14]), .Z(n1765) );
  NANDN U2896 ( .A(n1765), .B(n36107), .Z(n1681) );
  OR U2897 ( .A(n1679), .B(n36105), .Z(n1680) );
  AND U2898 ( .A(n1681), .B(n1680), .Z(n1718) );
  XNOR U2899 ( .A(n1719), .B(n1718), .Z(n1721) );
  XNOR U2900 ( .A(n1720), .B(n1721), .Z(n1740) );
  XOR U2901 ( .A(b[7]), .B(a[10]), .Z(n1722) );
  NAND U2902 ( .A(n1722), .B(n36701), .Z(n1684) );
  NAND U2903 ( .A(n1682), .B(n36702), .Z(n1683) );
  NAND U2904 ( .A(n1684), .B(n1683), .Z(n1737) );
  XNOR U2905 ( .A(b[11]), .B(a[6]), .Z(n1725) );
  OR U2906 ( .A(n1725), .B(n37311), .Z(n1687) );
  NAND U2907 ( .A(n1685), .B(n37218), .Z(n1686) );
  NAND U2908 ( .A(n1687), .B(n1686), .Z(n1734) );
  XNOR U2909 ( .A(b[15]), .B(a[2]), .Z(n1749) );
  OR U2910 ( .A(n1749), .B(n37665), .Z(n1690) );
  NAND U2911 ( .A(n1688), .B(n37604), .Z(n1689) );
  NAND U2912 ( .A(n1690), .B(n1689), .Z(n1731) );
  XNOR U2913 ( .A(b[5]), .B(a[12]), .Z(n1768) );
  NANDN U2914 ( .A(n1768), .B(n36587), .Z(n1693) );
  NANDN U2915 ( .A(n1691), .B(n36588), .Z(n1692) );
  AND U2916 ( .A(n1693), .B(n1692), .Z(n1732) );
  XNOR U2917 ( .A(n1731), .B(n1732), .Z(n1733) );
  XNOR U2918 ( .A(n1734), .B(n1733), .Z(n1738) );
  XNOR U2919 ( .A(n1737), .B(n1738), .Z(n1739) );
  XOR U2920 ( .A(n1740), .B(n1739), .Z(n1709) );
  XNOR U2921 ( .A(n1708), .B(n1709), .Z(n1771) );
  OR U2922 ( .A(n1695), .B(n1694), .Z(n1699) );
  NAND U2923 ( .A(n1697), .B(n1696), .Z(n1698) );
  AND U2924 ( .A(n1699), .B(n1698), .Z(n1772) );
  XNOR U2925 ( .A(n1771), .B(n1772), .Z(n1773) );
  XNOR U2926 ( .A(n1774), .B(n1773), .Z(n1701) );
  XNOR U2927 ( .A(n1700), .B(n1701), .Z(n1702) );
  XOR U2928 ( .A(n1703), .B(n1702), .Z(n1776) );
  XOR U2929 ( .A(n1777), .B(n1776), .Z(c[240]) );
  NANDN U2930 ( .A(n1701), .B(n1700), .Z(n1705) );
  NAND U2931 ( .A(n1703), .B(n1702), .Z(n1704) );
  NAND U2932 ( .A(n1705), .B(n1704), .Z(n1788) );
  NANDN U2933 ( .A(n1707), .B(n1706), .Z(n1711) );
  NAND U2934 ( .A(n1709), .B(n1708), .Z(n1710) );
  NAND U2935 ( .A(n1711), .B(n1710), .Z(n1854) );
  OR U2936 ( .A(n1713), .B(n1712), .Z(n1717) );
  NANDN U2937 ( .A(n1715), .B(n1714), .Z(n1716) );
  NAND U2938 ( .A(n1717), .B(n1716), .Z(n1855) );
  XNOR U2939 ( .A(n1854), .B(n1855), .Z(n1856) );
  XOR U2940 ( .A(b[7]), .B(a[11]), .Z(n1835) );
  NAND U2941 ( .A(n1835), .B(n36701), .Z(n1724) );
  NAND U2942 ( .A(n1722), .B(n36702), .Z(n1723) );
  NAND U2943 ( .A(n1724), .B(n1723), .Z(n1820) );
  XOR U2944 ( .A(b[11]), .B(a[7]), .Z(n1814) );
  NANDN U2945 ( .A(n37311), .B(n1814), .Z(n1727) );
  NANDN U2946 ( .A(n1725), .B(n37218), .Z(n1726) );
  NAND U2947 ( .A(n1727), .B(n1726), .Z(n1817) );
  XNOR U2948 ( .A(b[13]), .B(a[5]), .Z(n1829) );
  NANDN U2949 ( .A(n1829), .B(n37424), .Z(n1730) );
  NANDN U2950 ( .A(n1728), .B(n37425), .Z(n1729) );
  AND U2951 ( .A(n1730), .B(n1729), .Z(n1818) );
  XNOR U2952 ( .A(n1817), .B(n1818), .Z(n1819) );
  XOR U2953 ( .A(n1820), .B(n1819), .Z(n1849) );
  XNOR U2954 ( .A(n1848), .B(n1849), .Z(n1850) );
  NANDN U2955 ( .A(n1732), .B(n1731), .Z(n1736) );
  NAND U2956 ( .A(n1734), .B(n1733), .Z(n1735) );
  NAND U2957 ( .A(n1736), .B(n1735), .Z(n1851) );
  XOR U2958 ( .A(n1850), .B(n1851), .Z(n1794) );
  NANDN U2959 ( .A(n1738), .B(n1737), .Z(n1742) );
  NAND U2960 ( .A(n1740), .B(n1739), .Z(n1741) );
  NAND U2961 ( .A(n1742), .B(n1741), .Z(n1791) );
  NANDN U2962 ( .A(n1744), .B(n1743), .Z(n1748) );
  NAND U2963 ( .A(n1746), .B(n1745), .Z(n1747) );
  NAND U2964 ( .A(n1748), .B(n1747), .Z(n1841) );
  XNOR U2965 ( .A(n1054), .B(a[3]), .Z(n1806) );
  NANDN U2966 ( .A(n37665), .B(n1806), .Z(n1751) );
  NANDN U2967 ( .A(n1749), .B(n37604), .Z(n1750) );
  NAND U2968 ( .A(n1751), .B(n1750), .Z(n1810) );
  XOR U2969 ( .A(b[17]), .B(a[1]), .Z(n1811) );
  AND U2970 ( .A(n37764), .B(n1811), .Z(n1756) );
  XNOR U2971 ( .A(b[17]), .B(n3393), .Z(n1754) );
  XNOR U2972 ( .A(b[17]), .B(n1054), .Z(n1753) );
  XOR U2973 ( .A(b[17]), .B(b[16]), .Z(n1752) );
  AND U2974 ( .A(n1753), .B(n1752), .Z(n37762) );
  NAND U2975 ( .A(n1754), .B(n37762), .Z(n1755) );
  NANDN U2976 ( .A(n1756), .B(n1755), .Z(n1809) );
  XNOR U2977 ( .A(n1810), .B(n1809), .Z(n1800) );
  NANDN U2978 ( .A(b[16]), .B(n1054), .Z(n1757) );
  NANDN U2979 ( .A(n3393), .B(n1757), .Z(n1758) );
  NANDN U2980 ( .A(n1054), .B(b[16]), .Z(n37822) );
  AND U2981 ( .A(n37822), .B(b[17]), .Z(n38025) );
  NAND U2982 ( .A(n1758), .B(n38025), .Z(n1797) );
  XNOR U2983 ( .A(b[9]), .B(a[9]), .Z(n1826) );
  NANDN U2984 ( .A(n1826), .B(n36925), .Z(n1761) );
  NANDN U2985 ( .A(n1759), .B(n36926), .Z(n1760) );
  NAND U2986 ( .A(n1761), .B(n1760), .Z(n1798) );
  XNOR U2987 ( .A(n1797), .B(n1798), .Z(n1799) );
  XOR U2988 ( .A(n1800), .B(n1799), .Z(n1838) );
  NANDN U2989 ( .A(n1049), .B(a[17]), .Z(n1762) );
  XNOR U2990 ( .A(b[1]), .B(n1762), .Z(n1764) );
  NANDN U2991 ( .A(b[0]), .B(a[16]), .Z(n1763) );
  AND U2992 ( .A(n1764), .B(n1763), .Z(n1846) );
  XNOR U2993 ( .A(b[3]), .B(a[15]), .Z(n1823) );
  NANDN U2994 ( .A(n1823), .B(n36107), .Z(n1767) );
  OR U2995 ( .A(n1765), .B(n36105), .Z(n1766) );
  NAND U2996 ( .A(n1767), .B(n1766), .Z(n1844) );
  XNOR U2997 ( .A(n1051), .B(a[13]), .Z(n1832) );
  NAND U2998 ( .A(n1832), .B(n36587), .Z(n1770) );
  NANDN U2999 ( .A(n1768), .B(n36588), .Z(n1769) );
  AND U3000 ( .A(n1770), .B(n1769), .Z(n1845) );
  XNOR U3001 ( .A(n1844), .B(n1845), .Z(n1847) );
  XNOR U3002 ( .A(n1846), .B(n1847), .Z(n1839) );
  XOR U3003 ( .A(n1838), .B(n1839), .Z(n1840) );
  XNOR U3004 ( .A(n1841), .B(n1840), .Z(n1792) );
  XNOR U3005 ( .A(n1791), .B(n1792), .Z(n1793) );
  XNOR U3006 ( .A(n1794), .B(n1793), .Z(n1857) );
  XOR U3007 ( .A(n1856), .B(n1857), .Z(n1785) );
  XNOR U3008 ( .A(n1785), .B(n1786), .Z(n1787) );
  XNOR U3009 ( .A(n1788), .B(n1787), .Z(n1780) );
  XNOR U3010 ( .A(n1780), .B(sreg[241]), .Z(n1782) );
  NAND U3011 ( .A(n1775), .B(sreg[240]), .Z(n1779) );
  OR U3012 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U3013 ( .A(n1779), .B(n1778), .Z(n1781) );
  XOR U3014 ( .A(n1782), .B(n1781), .Z(c[241]) );
  NAND U3015 ( .A(n1780), .B(sreg[241]), .Z(n1784) );
  OR U3016 ( .A(n1782), .B(n1781), .Z(n1783) );
  NAND U3017 ( .A(n1784), .B(n1783), .Z(n1948) );
  XNOR U3018 ( .A(n1948), .B(sreg[242]), .Z(n1950) );
  NANDN U3019 ( .A(n1786), .B(n1785), .Z(n1790) );
  NAND U3020 ( .A(n1788), .B(n1787), .Z(n1789) );
  NAND U3021 ( .A(n1790), .B(n1789), .Z(n1863) );
  NANDN U3022 ( .A(n1792), .B(n1791), .Z(n1796) );
  NAND U3023 ( .A(n1794), .B(n1793), .Z(n1795) );
  NAND U3024 ( .A(n1796), .B(n1795), .Z(n1869) );
  NANDN U3025 ( .A(n1798), .B(n1797), .Z(n1802) );
  NAND U3026 ( .A(n1800), .B(n1799), .Z(n1801) );
  NAND U3027 ( .A(n1802), .B(n1801), .Z(n1945) );
  NANDN U3028 ( .A(n1049), .B(a[18]), .Z(n1803) );
  XNOR U3029 ( .A(b[1]), .B(n1803), .Z(n1805) );
  NANDN U3030 ( .A(b[0]), .B(a[17]), .Z(n1804) );
  AND U3031 ( .A(n1805), .B(n1804), .Z(n1909) );
  XNOR U3032 ( .A(b[15]), .B(a[4]), .Z(n1891) );
  OR U3033 ( .A(n1891), .B(n37665), .Z(n1808) );
  NAND U3034 ( .A(n1806), .B(n37604), .Z(n1807) );
  AND U3035 ( .A(n1808), .B(n1807), .Z(n1910) );
  XOR U3036 ( .A(n1909), .B(n1910), .Z(n1912) );
  XOR U3037 ( .A(b[17]), .B(b[18]), .Z(n37934) );
  NANDN U3038 ( .A(n3393), .B(n37934), .Z(n1911) );
  XNOR U3039 ( .A(n1912), .B(n1911), .Z(n1942) );
  NAND U3040 ( .A(n1810), .B(n1809), .Z(n1939) );
  XNOR U3041 ( .A(b[17]), .B(a[2]), .Z(n1915) );
  NANDN U3042 ( .A(n1915), .B(n37764), .Z(n1813) );
  NAND U3043 ( .A(n1811), .B(n37762), .Z(n1812) );
  NAND U3044 ( .A(n1813), .B(n1812), .Z(n1937) );
  XOR U3045 ( .A(b[11]), .B(a[8]), .Z(n1903) );
  NANDN U3046 ( .A(n37311), .B(n1903), .Z(n1816) );
  NAND U3047 ( .A(n37218), .B(n1814), .Z(n1815) );
  AND U3048 ( .A(n1816), .B(n1815), .Z(n1936) );
  XNOR U3049 ( .A(n1937), .B(n1936), .Z(n1938) );
  XNOR U3050 ( .A(n1939), .B(n1938), .Z(n1943) );
  XNOR U3051 ( .A(n1942), .B(n1943), .Z(n1944) );
  XNOR U3052 ( .A(n1945), .B(n1944), .Z(n1877) );
  NANDN U3053 ( .A(n1818), .B(n1817), .Z(n1822) );
  NAND U3054 ( .A(n1820), .B(n1819), .Z(n1821) );
  AND U3055 ( .A(n1822), .B(n1821), .Z(n1876) );
  XNOR U3056 ( .A(n1877), .B(n1876), .Z(n1878) );
  OR U3057 ( .A(n1823), .B(n36105), .Z(n1825) );
  XNOR U3058 ( .A(b[3]), .B(a[16]), .Z(n1897) );
  NANDN U3059 ( .A(n1897), .B(n36107), .Z(n1824) );
  NAND U3060 ( .A(n1825), .B(n1824), .Z(n1933) );
  XNOR U3061 ( .A(n1052), .B(a[10]), .Z(n1927) );
  NAND U3062 ( .A(n36925), .B(n1927), .Z(n1828) );
  NANDN U3063 ( .A(n1826), .B(n36926), .Z(n1827) );
  NAND U3064 ( .A(n1828), .B(n1827), .Z(n1930) );
  XOR U3065 ( .A(b[13]), .B(n4305), .Z(n1888) );
  NANDN U3066 ( .A(n1888), .B(n37424), .Z(n1831) );
  NANDN U3067 ( .A(n1829), .B(n37425), .Z(n1830) );
  AND U3068 ( .A(n1831), .B(n1830), .Z(n1931) );
  XNOR U3069 ( .A(n1930), .B(n1931), .Z(n1932) );
  XNOR U3070 ( .A(n1933), .B(n1932), .Z(n1885) );
  XNOR U3071 ( .A(b[5]), .B(a[14]), .Z(n1894) );
  NANDN U3072 ( .A(n1894), .B(n36587), .Z(n1834) );
  NAND U3073 ( .A(n36588), .B(n1832), .Z(n1833) );
  NAND U3074 ( .A(n1834), .B(n1833), .Z(n1883) );
  XNOR U3075 ( .A(b[7]), .B(a[12]), .Z(n1906) );
  NANDN U3076 ( .A(n1906), .B(n36701), .Z(n1837) );
  NAND U3077 ( .A(n36702), .B(n1835), .Z(n1836) );
  AND U3078 ( .A(n1837), .B(n1836), .Z(n1882) );
  XNOR U3079 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U3080 ( .A(n1885), .B(n1884), .Z(n1879) );
  XOR U3081 ( .A(n1878), .B(n1879), .Z(n1872) );
  OR U3082 ( .A(n1839), .B(n1838), .Z(n1843) );
  NAND U3083 ( .A(n1841), .B(n1840), .Z(n1842) );
  NAND U3084 ( .A(n1843), .B(n1842), .Z(n1871) );
  XNOR U3085 ( .A(n1871), .B(n1870), .Z(n1873) );
  XNOR U3086 ( .A(n1872), .B(n1873), .Z(n1866) );
  NANDN U3087 ( .A(n1849), .B(n1848), .Z(n1853) );
  NANDN U3088 ( .A(n1851), .B(n1850), .Z(n1852) );
  NAND U3089 ( .A(n1853), .B(n1852), .Z(n1867) );
  XNOR U3090 ( .A(n1866), .B(n1867), .Z(n1868) );
  XNOR U3091 ( .A(n1869), .B(n1868), .Z(n1860) );
  NANDN U3092 ( .A(n1855), .B(n1854), .Z(n1859) );
  NANDN U3093 ( .A(n1857), .B(n1856), .Z(n1858) );
  NAND U3094 ( .A(n1859), .B(n1858), .Z(n1861) );
  XNOR U3095 ( .A(n1860), .B(n1861), .Z(n1862) );
  XOR U3096 ( .A(n1863), .B(n1862), .Z(n1949) );
  XOR U3097 ( .A(n1950), .B(n1949), .Z(c[242]) );
  NANDN U3098 ( .A(n1861), .B(n1860), .Z(n1865) );
  NAND U3099 ( .A(n1863), .B(n1862), .Z(n1864) );
  NAND U3100 ( .A(n1865), .B(n1864), .Z(n1961) );
  NANDN U3101 ( .A(n1871), .B(n1870), .Z(n1875) );
  NAND U3102 ( .A(n1873), .B(n1872), .Z(n1874) );
  NAND U3103 ( .A(n1875), .B(n1874), .Z(n1964) );
  NANDN U3104 ( .A(n1877), .B(n1876), .Z(n1881) );
  NAND U3105 ( .A(n1879), .B(n1878), .Z(n1880) );
  NAND U3106 ( .A(n1881), .B(n1880), .Z(n1963) );
  NANDN U3107 ( .A(n1883), .B(n1882), .Z(n1887) );
  NAND U3108 ( .A(n1885), .B(n1884), .Z(n1886) );
  NAND U3109 ( .A(n1887), .B(n1886), .Z(n1969) );
  XNOR U3110 ( .A(b[13]), .B(a[7]), .Z(n2022) );
  NANDN U3111 ( .A(n2022), .B(n37424), .Z(n1890) );
  NANDN U3112 ( .A(n1888), .B(n37425), .Z(n1889) );
  NAND U3113 ( .A(n1890), .B(n1889), .Z(n1983) );
  XNOR U3114 ( .A(b[15]), .B(a[5]), .Z(n2019) );
  OR U3115 ( .A(n2019), .B(n37665), .Z(n1893) );
  NANDN U3116 ( .A(n1891), .B(n37604), .Z(n1892) );
  NAND U3117 ( .A(n1893), .B(n1892), .Z(n1980) );
  XNOR U3118 ( .A(n1051), .B(a[15]), .Z(n1995) );
  NAND U3119 ( .A(n1995), .B(n36587), .Z(n1896) );
  NANDN U3120 ( .A(n1894), .B(n36588), .Z(n1895) );
  AND U3121 ( .A(n1896), .B(n1895), .Z(n1981) );
  XNOR U3122 ( .A(n1980), .B(n1981), .Z(n1982) );
  XNOR U3123 ( .A(n1983), .B(n1982), .Z(n2031) );
  OR U3124 ( .A(n1897), .B(n36105), .Z(n1899) );
  XNOR U3125 ( .A(n1050), .B(a[17]), .Z(n1992) );
  NAND U3126 ( .A(n1992), .B(n36107), .Z(n1898) );
  NAND U3127 ( .A(n1899), .B(n1898), .Z(n2010) );
  NANDN U3128 ( .A(n1049), .B(a[19]), .Z(n1900) );
  XNOR U3129 ( .A(b[1]), .B(n1900), .Z(n1902) );
  NANDN U3130 ( .A(b[0]), .B(a[18]), .Z(n1901) );
  AND U3131 ( .A(n1902), .B(n1901), .Z(n2007) );
  XOR U3132 ( .A(b[11]), .B(a[9]), .Z(n2016) );
  NANDN U3133 ( .A(n37311), .B(n2016), .Z(n1905) );
  NAND U3134 ( .A(n1903), .B(n37218), .Z(n1904) );
  AND U3135 ( .A(n1905), .B(n1904), .Z(n2008) );
  XNOR U3136 ( .A(n2007), .B(n2008), .Z(n2009) );
  XNOR U3137 ( .A(n2010), .B(n2009), .Z(n2028) );
  XOR U3138 ( .A(b[7]), .B(a[13]), .Z(n1998) );
  NAND U3139 ( .A(n36701), .B(n1998), .Z(n1908) );
  NANDN U3140 ( .A(n1906), .B(n36702), .Z(n1907) );
  NAND U3141 ( .A(n1908), .B(n1907), .Z(n2029) );
  XNOR U3142 ( .A(n2028), .B(n2029), .Z(n2030) );
  XOR U3143 ( .A(n2031), .B(n2030), .Z(n1968) );
  XNOR U3144 ( .A(n1969), .B(n1968), .Z(n1971) );
  NANDN U3145 ( .A(n1910), .B(n1909), .Z(n1914) );
  OR U3146 ( .A(n1912), .B(n1911), .Z(n1913) );
  AND U3147 ( .A(n1914), .B(n1913), .Z(n1970) );
  XNOR U3148 ( .A(n1971), .B(n1970), .Z(n1977) );
  NANDN U3149 ( .A(n1915), .B(n37762), .Z(n1917) );
  XOR U3150 ( .A(b[17]), .B(a[3]), .Z(n1989) );
  NAND U3151 ( .A(n1989), .B(n37764), .Z(n1916) );
  NAND U3152 ( .A(n1917), .B(n1916), .Z(n2012) );
  XNOR U3153 ( .A(n1055), .B(a[0]), .Z(n1920) );
  XNOR U3154 ( .A(n1055), .B(b[17]), .Z(n1919) );
  XNOR U3155 ( .A(n1055), .B(b[18]), .Z(n1918) );
  AND U3156 ( .A(n1919), .B(n1918), .Z(n37935) );
  NAND U3157 ( .A(n1920), .B(n37935), .Z(n1922) );
  XNOR U3158 ( .A(n1055), .B(a[1]), .Z(n2013) );
  NAND U3159 ( .A(n2013), .B(n37934), .Z(n1921) );
  NAND U3160 ( .A(n1922), .B(n1921), .Z(n2011) );
  XNOR U3161 ( .A(n2012), .B(n2011), .Z(n2004) );
  ANDN U3162 ( .B(b[17]), .A(n3393), .Z(n1923) );
  OR U3163 ( .A(n1923), .B(b[18]), .Z(n1925) );
  OR U3164 ( .A(b[17]), .B(a[0]), .Z(n1924) );
  NAND U3165 ( .A(n1925), .B(n1924), .Z(n1926) );
  AND U3166 ( .A(n1926), .B(b[19]), .Z(n2001) );
  XOR U3167 ( .A(n1052), .B(a[11]), .Z(n2025) );
  NANDN U3168 ( .A(n2025), .B(n36925), .Z(n1929) );
  NAND U3169 ( .A(n36926), .B(n1927), .Z(n1928) );
  NAND U3170 ( .A(n1929), .B(n1928), .Z(n2002) );
  XOR U3171 ( .A(n2001), .B(n2002), .Z(n2003) );
  XOR U3172 ( .A(n2004), .B(n2003), .Z(n2035) );
  NANDN U3173 ( .A(n1931), .B(n1930), .Z(n1935) );
  NAND U3174 ( .A(n1933), .B(n1932), .Z(n1934) );
  AND U3175 ( .A(n1935), .B(n1934), .Z(n2034) );
  XOR U3176 ( .A(n2035), .B(n2034), .Z(n2036) );
  NANDN U3177 ( .A(n1937), .B(n1936), .Z(n1941) );
  NAND U3178 ( .A(n1939), .B(n1938), .Z(n1940) );
  NAND U3179 ( .A(n1941), .B(n1940), .Z(n2037) );
  XOR U3180 ( .A(n2036), .B(n2037), .Z(n1974) );
  NANDN U3181 ( .A(n1943), .B(n1942), .Z(n1947) );
  NAND U3182 ( .A(n1945), .B(n1944), .Z(n1946) );
  AND U3183 ( .A(n1947), .B(n1946), .Z(n1975) );
  XNOR U3184 ( .A(n1974), .B(n1975), .Z(n1976) );
  XOR U3185 ( .A(n1977), .B(n1976), .Z(n1962) );
  XNOR U3186 ( .A(n1963), .B(n1962), .Z(n1965) );
  XNOR U3187 ( .A(n1964), .B(n1965), .Z(n1958) );
  XNOR U3188 ( .A(n1959), .B(n1958), .Z(n1960) );
  XNOR U3189 ( .A(n1961), .B(n1960), .Z(n1953) );
  XNOR U3190 ( .A(n1953), .B(sreg[243]), .Z(n1955) );
  NAND U3191 ( .A(n1948), .B(sreg[242]), .Z(n1952) );
  OR U3192 ( .A(n1950), .B(n1949), .Z(n1951) );
  AND U3193 ( .A(n1952), .B(n1951), .Z(n1954) );
  XOR U3194 ( .A(n1955), .B(n1954), .Z(c[243]) );
  NAND U3195 ( .A(n1953), .B(sreg[243]), .Z(n1957) );
  OR U3196 ( .A(n1955), .B(n1954), .Z(n1956) );
  NAND U3197 ( .A(n1957), .B(n1956), .Z(n2136) );
  XNOR U3198 ( .A(n2136), .B(sreg[244]), .Z(n2138) );
  NAND U3199 ( .A(n1963), .B(n1962), .Z(n1967) );
  NANDN U3200 ( .A(n1965), .B(n1964), .Z(n1966) );
  NAND U3201 ( .A(n1967), .B(n1966), .Z(n2040) );
  OR U3202 ( .A(n1969), .B(n1968), .Z(n1973) );
  OR U3203 ( .A(n1971), .B(n1970), .Z(n1972) );
  NAND U3204 ( .A(n1973), .B(n1972), .Z(n2049) );
  NANDN U3205 ( .A(n1975), .B(n1974), .Z(n1979) );
  NAND U3206 ( .A(n1977), .B(n1976), .Z(n1978) );
  NAND U3207 ( .A(n1979), .B(n1978), .Z(n2046) );
  NANDN U3208 ( .A(n1981), .B(n1980), .Z(n1985) );
  NAND U3209 ( .A(n1983), .B(n1982), .Z(n1984) );
  NAND U3210 ( .A(n1985), .B(n1984), .Z(n2067) );
  NANDN U3211 ( .A(n1049), .B(a[20]), .Z(n1986) );
  XNOR U3212 ( .A(b[1]), .B(n1986), .Z(n1988) );
  NANDN U3213 ( .A(b[0]), .B(a[19]), .Z(n1987) );
  AND U3214 ( .A(n1988), .B(n1987), .Z(n2102) );
  NAND U3215 ( .A(n1989), .B(n37762), .Z(n1991) );
  XOR U3216 ( .A(b[17]), .B(a[4]), .Z(n2126) );
  NAND U3217 ( .A(n2126), .B(n37764), .Z(n1990) );
  AND U3218 ( .A(n1991), .B(n1990), .Z(n2103) );
  XOR U3219 ( .A(n2102), .B(n2103), .Z(n2105) );
  IV U3220 ( .A(b[20]), .Z(n38141) );
  XOR U3221 ( .A(n1055), .B(n38141), .Z(n38101) );
  NANDN U3222 ( .A(n3393), .B(n38101), .Z(n2104) );
  XOR U3223 ( .A(n2105), .B(n2104), .Z(n2064) );
  XNOR U3224 ( .A(b[3]), .B(a[18]), .Z(n2111) );
  NANDN U3225 ( .A(n2111), .B(n36107), .Z(n1994) );
  NANDN U3226 ( .A(n36105), .B(n1992), .Z(n1993) );
  AND U3227 ( .A(n1994), .B(n1993), .Z(n2073) );
  XNOR U3228 ( .A(b[5]), .B(a[16]), .Z(n2120) );
  NANDN U3229 ( .A(n2120), .B(n36587), .Z(n1997) );
  NAND U3230 ( .A(n36588), .B(n1995), .Z(n1996) );
  AND U3231 ( .A(n1997), .B(n1996), .Z(n2070) );
  XOR U3232 ( .A(b[7]), .B(a[14]), .Z(n2117) );
  NAND U3233 ( .A(n2117), .B(n36701), .Z(n2000) );
  NAND U3234 ( .A(n1998), .B(n36702), .Z(n1999) );
  AND U3235 ( .A(n2000), .B(n1999), .Z(n2071) );
  XNOR U3236 ( .A(n2070), .B(n2071), .Z(n2072) );
  XNOR U3237 ( .A(n2064), .B(n2065), .Z(n2066) );
  XNOR U3238 ( .A(n2067), .B(n2066), .Z(n2059) );
  OR U3239 ( .A(n2002), .B(n2001), .Z(n2006) );
  NAND U3240 ( .A(n2004), .B(n2003), .Z(n2005) );
  AND U3241 ( .A(n2006), .B(n2005), .Z(n2058) );
  XNOR U3242 ( .A(n2059), .B(n2058), .Z(n2060) );
  NAND U3243 ( .A(n2012), .B(n2011), .Z(n2134) );
  XNOR U3244 ( .A(b[19]), .B(a[2]), .Z(n2088) );
  NANDN U3245 ( .A(n2088), .B(n37934), .Z(n2015) );
  NAND U3246 ( .A(n37935), .B(n2013), .Z(n2014) );
  NAND U3247 ( .A(n2015), .B(n2014), .Z(n2133) );
  XNOR U3248 ( .A(b[11]), .B(a[10]), .Z(n2099) );
  OR U3249 ( .A(n2099), .B(n37311), .Z(n2018) );
  NAND U3250 ( .A(n37218), .B(n2016), .Z(n2017) );
  AND U3251 ( .A(n2018), .B(n2017), .Z(n2132) );
  XNOR U3252 ( .A(n2133), .B(n2132), .Z(n2135) );
  XNOR U3253 ( .A(n2134), .B(n2135), .Z(n2082) );
  XNOR U3254 ( .A(n1054), .B(a[6]), .Z(n2129) );
  NANDN U3255 ( .A(n37665), .B(n2129), .Z(n2021) );
  NANDN U3256 ( .A(n2019), .B(n37604), .Z(n2020) );
  AND U3257 ( .A(n2021), .B(n2020), .Z(n2076) );
  XNOR U3258 ( .A(b[13]), .B(a[8]), .Z(n2123) );
  NANDN U3259 ( .A(n2123), .B(n37424), .Z(n2024) );
  NANDN U3260 ( .A(n2022), .B(n37425), .Z(n2023) );
  AND U3261 ( .A(n2024), .B(n2023), .Z(n2077) );
  XNOR U3262 ( .A(n2076), .B(n2077), .Z(n2078) );
  XOR U3263 ( .A(n1052), .B(a[12]), .Z(n2114) );
  NANDN U3264 ( .A(n2114), .B(n36925), .Z(n2027) );
  NANDN U3265 ( .A(n2025), .B(n36926), .Z(n2026) );
  AND U3266 ( .A(n2027), .B(n2026), .Z(n2079) );
  XNOR U3267 ( .A(n2082), .B(n2083), .Z(n2084) );
  XNOR U3268 ( .A(n2085), .B(n2084), .Z(n2061) );
  XOR U3269 ( .A(n2060), .B(n2061), .Z(n2055) );
  NANDN U3270 ( .A(n2029), .B(n2028), .Z(n2033) );
  NAND U3271 ( .A(n2031), .B(n2030), .Z(n2032) );
  NAND U3272 ( .A(n2033), .B(n2032), .Z(n2052) );
  OR U3273 ( .A(n2035), .B(n2034), .Z(n2039) );
  NANDN U3274 ( .A(n2037), .B(n2036), .Z(n2038) );
  NAND U3275 ( .A(n2039), .B(n2038), .Z(n2053) );
  XNOR U3276 ( .A(n2052), .B(n2053), .Z(n2054) );
  XNOR U3277 ( .A(n2055), .B(n2054), .Z(n2047) );
  XNOR U3278 ( .A(n2046), .B(n2047), .Z(n2048) );
  XOR U3279 ( .A(n2049), .B(n2048), .Z(n2041) );
  XNOR U3280 ( .A(n2040), .B(n2041), .Z(n2042) );
  XOR U3281 ( .A(n2043), .B(n2042), .Z(n2137) );
  XOR U3282 ( .A(n2138), .B(n2137), .Z(c[244]) );
  NANDN U3283 ( .A(n2041), .B(n2040), .Z(n2045) );
  NAND U3284 ( .A(n2043), .B(n2042), .Z(n2044) );
  NAND U3285 ( .A(n2045), .B(n2044), .Z(n2149) );
  NANDN U3286 ( .A(n2047), .B(n2046), .Z(n2051) );
  NANDN U3287 ( .A(n2049), .B(n2048), .Z(n2050) );
  NAND U3288 ( .A(n2051), .B(n2050), .Z(n2146) );
  NANDN U3289 ( .A(n2053), .B(n2052), .Z(n2057) );
  NAND U3290 ( .A(n2055), .B(n2054), .Z(n2056) );
  NAND U3291 ( .A(n2057), .B(n2056), .Z(n2238) );
  NANDN U3292 ( .A(n2059), .B(n2058), .Z(n2063) );
  NANDN U3293 ( .A(n2061), .B(n2060), .Z(n2062) );
  NAND U3294 ( .A(n2063), .B(n2062), .Z(n2236) );
  NANDN U3295 ( .A(n2065), .B(n2064), .Z(n2069) );
  NAND U3296 ( .A(n2067), .B(n2066), .Z(n2068) );
  NAND U3297 ( .A(n2069), .B(n2068), .Z(n2230) );
  OR U3298 ( .A(n2071), .B(n2070), .Z(n2075) );
  OR U3299 ( .A(n2073), .B(n2072), .Z(n2074) );
  NAND U3300 ( .A(n2075), .B(n2074), .Z(n2229) );
  XOR U3301 ( .A(n2230), .B(n2229), .Z(n2231) );
  OR U3302 ( .A(n2077), .B(n2076), .Z(n2081) );
  OR U3303 ( .A(n2079), .B(n2078), .Z(n2080) );
  NAND U3304 ( .A(n2081), .B(n2080), .Z(n2232) );
  XNOR U3305 ( .A(n2231), .B(n2232), .Z(n2225) );
  NANDN U3306 ( .A(n2083), .B(n2082), .Z(n2087) );
  NAND U3307 ( .A(n2085), .B(n2084), .Z(n2086) );
  NAND U3308 ( .A(n2087), .B(n2086), .Z(n2224) );
  XNOR U3309 ( .A(b[19]), .B(a[3]), .Z(n2214) );
  NANDN U3310 ( .A(n2214), .B(n37934), .Z(n2090) );
  NANDN U3311 ( .A(n2088), .B(n37935), .Z(n2089) );
  NAND U3312 ( .A(n2090), .B(n2089), .Z(n2204) );
  XNOR U3313 ( .A(b[21]), .B(a[1]), .Z(n2173) );
  ANDN U3314 ( .B(n38101), .A(n2173), .Z(n2095) );
  XNOR U3315 ( .A(n1056), .B(a[0]), .Z(n2093) );
  XNOR U3316 ( .A(n1056), .B(b[19]), .Z(n2092) );
  XNOR U3317 ( .A(n1056), .B(b[20]), .Z(n2091) );
  AND U3318 ( .A(n2092), .B(n2091), .Z(n38102) );
  NAND U3319 ( .A(n2093), .B(n38102), .Z(n2094) );
  NANDN U3320 ( .A(n2095), .B(n2094), .Z(n2203) );
  XNOR U3321 ( .A(n2204), .B(n2203), .Z(n2200) );
  NANDN U3322 ( .A(n1055), .B(b[20]), .Z(n38212) );
  ANDN U3323 ( .B(n38212), .A(n1056), .Z(n2098) );
  XNOR U3324 ( .A(n38141), .B(b[19]), .Z(n2096) );
  NANDN U3325 ( .A(n3393), .B(n2096), .Z(n2097) );
  AND U3326 ( .A(n2098), .B(n2097), .Z(n2198) );
  XNOR U3327 ( .A(b[11]), .B(a[11]), .Z(n2176) );
  OR U3328 ( .A(n2176), .B(n37311), .Z(n2101) );
  NANDN U3329 ( .A(n2099), .B(n37218), .Z(n2100) );
  AND U3330 ( .A(n2101), .B(n2100), .Z(n2197) );
  XNOR U3331 ( .A(n2198), .B(n2197), .Z(n2199) );
  XOR U3332 ( .A(n2200), .B(n2199), .Z(n2155) );
  NANDN U3333 ( .A(n2103), .B(n2102), .Z(n2107) );
  OR U3334 ( .A(n2105), .B(n2104), .Z(n2106) );
  NAND U3335 ( .A(n2107), .B(n2106), .Z(n2153) );
  NANDN U3336 ( .A(n1049), .B(a[21]), .Z(n2108) );
  XNOR U3337 ( .A(b[1]), .B(n2108), .Z(n2110) );
  NANDN U3338 ( .A(b[0]), .B(a[20]), .Z(n2109) );
  AND U3339 ( .A(n2110), .B(n2109), .Z(n2186) );
  XNOR U3340 ( .A(b[3]), .B(a[19]), .Z(n2208) );
  NANDN U3341 ( .A(n2208), .B(n36107), .Z(n2113) );
  OR U3342 ( .A(n2111), .B(n36105), .Z(n2112) );
  AND U3343 ( .A(n2113), .B(n2112), .Z(n2185) );
  XNOR U3344 ( .A(n2186), .B(n2185), .Z(n2187) );
  XNOR U3345 ( .A(b[9]), .B(a[13]), .Z(n2167) );
  NANDN U3346 ( .A(n2167), .B(n36925), .Z(n2116) );
  NANDN U3347 ( .A(n2114), .B(n36926), .Z(n2115) );
  NAND U3348 ( .A(n2116), .B(n2115), .Z(n2188) );
  XOR U3349 ( .A(n2187), .B(n2188), .Z(n2152) );
  XOR U3350 ( .A(n2153), .B(n2152), .Z(n2154) );
  XOR U3351 ( .A(n2155), .B(n2154), .Z(n2219) );
  XOR U3352 ( .A(b[7]), .B(a[15]), .Z(n2158) );
  NAND U3353 ( .A(n2158), .B(n36701), .Z(n2119) );
  NAND U3354 ( .A(n2117), .B(n36702), .Z(n2118) );
  NAND U3355 ( .A(n2119), .B(n2118), .Z(n2191) );
  XNOR U3356 ( .A(b[5]), .B(a[17]), .Z(n2161) );
  NANDN U3357 ( .A(n2161), .B(n36587), .Z(n2122) );
  NANDN U3358 ( .A(n2120), .B(n36588), .Z(n2121) );
  AND U3359 ( .A(n2122), .B(n2121), .Z(n2192) );
  XNOR U3360 ( .A(n2191), .B(n2192), .Z(n2193) );
  XNOR U3361 ( .A(n1053), .B(a[9]), .Z(n2205) );
  NAND U3362 ( .A(n2205), .B(n37424), .Z(n2125) );
  NANDN U3363 ( .A(n2123), .B(n37425), .Z(n2124) );
  NAND U3364 ( .A(n2125), .B(n2124), .Z(n2182) );
  NAND U3365 ( .A(n2126), .B(n37762), .Z(n2128) );
  XOR U3366 ( .A(b[17]), .B(a[5]), .Z(n2170) );
  NAND U3367 ( .A(n2170), .B(n37764), .Z(n2127) );
  NAND U3368 ( .A(n2128), .B(n2127), .Z(n2179) );
  XNOR U3369 ( .A(b[15]), .B(a[7]), .Z(n2164) );
  OR U3370 ( .A(n2164), .B(n37665), .Z(n2131) );
  NAND U3371 ( .A(n2129), .B(n37604), .Z(n2130) );
  AND U3372 ( .A(n2131), .B(n2130), .Z(n2180) );
  XNOR U3373 ( .A(n2179), .B(n2180), .Z(n2181) );
  XOR U3374 ( .A(n2182), .B(n2181), .Z(n2194) );
  XOR U3375 ( .A(n2193), .B(n2194), .Z(n2217) );
  XNOR U3376 ( .A(n2217), .B(n2218), .Z(n2220) );
  XOR U3377 ( .A(n2219), .B(n2220), .Z(n2223) );
  XNOR U3378 ( .A(n2224), .B(n2223), .Z(n2226) );
  XOR U3379 ( .A(n2225), .B(n2226), .Z(n2235) );
  XNOR U3380 ( .A(n2236), .B(n2235), .Z(n2237) );
  XOR U3381 ( .A(n2238), .B(n2237), .Z(n2147) );
  XNOR U3382 ( .A(n2146), .B(n2147), .Z(n2148) );
  XNOR U3383 ( .A(n2149), .B(n2148), .Z(n2141) );
  XNOR U3384 ( .A(n2141), .B(sreg[245]), .Z(n2143) );
  NAND U3385 ( .A(n2136), .B(sreg[244]), .Z(n2140) );
  OR U3386 ( .A(n2138), .B(n2137), .Z(n2139) );
  AND U3387 ( .A(n2140), .B(n2139), .Z(n2142) );
  XOR U3388 ( .A(n2143), .B(n2142), .Z(c[245]) );
  NAND U3389 ( .A(n2141), .B(sreg[245]), .Z(n2145) );
  OR U3390 ( .A(n2143), .B(n2142), .Z(n2144) );
  NAND U3391 ( .A(n2145), .B(n2144), .Z(n2345) );
  XNOR U3392 ( .A(n2345), .B(sreg[246]), .Z(n2347) );
  NANDN U3393 ( .A(n2147), .B(n2146), .Z(n2151) );
  NAND U3394 ( .A(n2149), .B(n2148), .Z(n2150) );
  NAND U3395 ( .A(n2151), .B(n2150), .Z(n2244) );
  OR U3396 ( .A(n2153), .B(n2152), .Z(n2157) );
  NAND U3397 ( .A(n2155), .B(n2154), .Z(n2156) );
  NAND U3398 ( .A(n2157), .B(n2156), .Z(n2256) );
  XOR U3399 ( .A(b[7]), .B(a[16]), .Z(n2265) );
  NAND U3400 ( .A(n2265), .B(n36701), .Z(n2160) );
  NAND U3401 ( .A(n2158), .B(n36702), .Z(n2159) );
  NAND U3402 ( .A(n2160), .B(n2159), .Z(n2291) );
  XNOR U3403 ( .A(b[5]), .B(a[18]), .Z(n2271) );
  NANDN U3404 ( .A(n2271), .B(n36587), .Z(n2163) );
  NANDN U3405 ( .A(n2161), .B(n36588), .Z(n2162) );
  NAND U3406 ( .A(n2163), .B(n2162), .Z(n2288) );
  XNOR U3407 ( .A(b[15]), .B(a[8]), .Z(n2318) );
  OR U3408 ( .A(n2318), .B(n37665), .Z(n2166) );
  NANDN U3409 ( .A(n2164), .B(n37604), .Z(n2165) );
  AND U3410 ( .A(n2166), .B(n2165), .Z(n2289) );
  XNOR U3411 ( .A(n2288), .B(n2289), .Z(n2290) );
  XNOR U3412 ( .A(n2291), .B(n2290), .Z(n2323) );
  XNOR U3413 ( .A(b[9]), .B(a[14]), .Z(n2268) );
  NANDN U3414 ( .A(n2268), .B(n36925), .Z(n2169) );
  NANDN U3415 ( .A(n2167), .B(n36926), .Z(n2168) );
  NAND U3416 ( .A(n2169), .B(n2168), .Z(n2297) );
  NAND U3417 ( .A(n2170), .B(n37762), .Z(n2172) );
  XNOR U3418 ( .A(b[17]), .B(a[6]), .Z(n2306) );
  NANDN U3419 ( .A(n2306), .B(n37764), .Z(n2171) );
  NAND U3420 ( .A(n2172), .B(n2171), .Z(n2294) );
  XNOR U3421 ( .A(b[21]), .B(a[2]), .Z(n2280) );
  NANDN U3422 ( .A(n2280), .B(n38101), .Z(n2175) );
  NANDN U3423 ( .A(n2173), .B(n38102), .Z(n2174) );
  AND U3424 ( .A(n2175), .B(n2174), .Z(n2295) );
  XNOR U3425 ( .A(n2294), .B(n2295), .Z(n2296) );
  XNOR U3426 ( .A(n2297), .B(n2296), .Z(n2321) );
  XOR U3427 ( .A(b[11]), .B(a[12]), .Z(n2277) );
  NANDN U3428 ( .A(n37311), .B(n2277), .Z(n2178) );
  NANDN U3429 ( .A(n2176), .B(n37218), .Z(n2177) );
  NAND U3430 ( .A(n2178), .B(n2177), .Z(n2322) );
  XOR U3431 ( .A(n2321), .B(n2322), .Z(n2324) );
  XNOR U3432 ( .A(n2323), .B(n2324), .Z(n2342) );
  NANDN U3433 ( .A(n2180), .B(n2179), .Z(n2184) );
  NAND U3434 ( .A(n2182), .B(n2181), .Z(n2183) );
  NAND U3435 ( .A(n2184), .B(n2183), .Z(n2339) );
  NANDN U3436 ( .A(n2186), .B(n2185), .Z(n2190) );
  NANDN U3437 ( .A(n2188), .B(n2187), .Z(n2189) );
  NAND U3438 ( .A(n2190), .B(n2189), .Z(n2340) );
  XNOR U3439 ( .A(n2339), .B(n2340), .Z(n2341) );
  XNOR U3440 ( .A(n2342), .B(n2341), .Z(n2329) );
  NANDN U3441 ( .A(n2192), .B(n2191), .Z(n2196) );
  NAND U3442 ( .A(n2194), .B(n2193), .Z(n2195) );
  NAND U3443 ( .A(n2196), .B(n2195), .Z(n2328) );
  NANDN U3444 ( .A(n2198), .B(n2197), .Z(n2202) );
  NAND U3445 ( .A(n2200), .B(n2199), .Z(n2201) );
  NAND U3446 ( .A(n2202), .B(n2201), .Z(n2333) );
  NAND U3447 ( .A(n2204), .B(n2203), .Z(n2262) );
  XNOR U3448 ( .A(b[13]), .B(a[10]), .Z(n2312) );
  NANDN U3449 ( .A(n2312), .B(n37424), .Z(n2207) );
  NAND U3450 ( .A(n37425), .B(n2205), .Z(n2206) );
  NAND U3451 ( .A(n2207), .B(n2206), .Z(n2260) );
  XNOR U3452 ( .A(b[3]), .B(a[20]), .Z(n2315) );
  NANDN U3453 ( .A(n2315), .B(n36107), .Z(n2210) );
  OR U3454 ( .A(n2208), .B(n36105), .Z(n2209) );
  AND U3455 ( .A(n2210), .B(n2209), .Z(n2259) );
  XNOR U3456 ( .A(n2260), .B(n2259), .Z(n2261) );
  XNOR U3457 ( .A(n2262), .B(n2261), .Z(n2334) );
  XNOR U3458 ( .A(n2333), .B(n2334), .Z(n2335) );
  XOR U3459 ( .A(n1056), .B(b[22]), .Z(n38268) );
  NOR U3460 ( .A(n3393), .B(n38268), .Z(n2303) );
  NANDN U3461 ( .A(n1049), .B(a[22]), .Z(n2211) );
  XNOR U3462 ( .A(b[1]), .B(n2211), .Z(n2213) );
  NANDN U3463 ( .A(b[0]), .B(a[21]), .Z(n2212) );
  AND U3464 ( .A(n2213), .B(n2212), .Z(n2301) );
  XNOR U3465 ( .A(b[19]), .B(a[4]), .Z(n2309) );
  NANDN U3466 ( .A(n2309), .B(n37934), .Z(n2216) );
  NANDN U3467 ( .A(n2214), .B(n37935), .Z(n2215) );
  AND U3468 ( .A(n2216), .B(n2215), .Z(n2300) );
  XNOR U3469 ( .A(n2301), .B(n2300), .Z(n2302) );
  XOR U3470 ( .A(n2303), .B(n2302), .Z(n2336) );
  XNOR U3471 ( .A(n2335), .B(n2336), .Z(n2327) );
  XOR U3472 ( .A(n2328), .B(n2327), .Z(n2330) );
  XOR U3473 ( .A(n2329), .B(n2330), .Z(n2253) );
  NAND U3474 ( .A(n2218), .B(n2217), .Z(n2222) );
  OR U3475 ( .A(n2220), .B(n2219), .Z(n2221) );
  AND U3476 ( .A(n2222), .B(n2221), .Z(n2254) );
  XOR U3477 ( .A(n2253), .B(n2254), .Z(n2255) );
  XNOR U3478 ( .A(n2256), .B(n2255), .Z(n2247) );
  NAND U3479 ( .A(n2224), .B(n2223), .Z(n2228) );
  OR U3480 ( .A(n2226), .B(n2225), .Z(n2227) );
  AND U3481 ( .A(n2228), .B(n2227), .Z(n2248) );
  XOR U3482 ( .A(n2247), .B(n2248), .Z(n2250) );
  OR U3483 ( .A(n2230), .B(n2229), .Z(n2234) );
  NANDN U3484 ( .A(n2232), .B(n2231), .Z(n2233) );
  NAND U3485 ( .A(n2234), .B(n2233), .Z(n2249) );
  XNOR U3486 ( .A(n2250), .B(n2249), .Z(n2241) );
  NAND U3487 ( .A(n2236), .B(n2235), .Z(n2240) );
  OR U3488 ( .A(n2238), .B(n2237), .Z(n2239) );
  NAND U3489 ( .A(n2240), .B(n2239), .Z(n2242) );
  XNOR U3490 ( .A(n2241), .B(n2242), .Z(n2243) );
  XOR U3491 ( .A(n2244), .B(n2243), .Z(n2346) );
  XOR U3492 ( .A(n2347), .B(n2346), .Z(c[246]) );
  NANDN U3493 ( .A(n2242), .B(n2241), .Z(n2246) );
  NAND U3494 ( .A(n2244), .B(n2243), .Z(n2245) );
  NAND U3495 ( .A(n2246), .B(n2245), .Z(n2358) );
  NANDN U3496 ( .A(n2248), .B(n2247), .Z(n2252) );
  OR U3497 ( .A(n2250), .B(n2249), .Z(n2251) );
  NAND U3498 ( .A(n2252), .B(n2251), .Z(n2356) );
  NAND U3499 ( .A(n2254), .B(n2253), .Z(n2258) );
  NAND U3500 ( .A(n2256), .B(n2255), .Z(n2257) );
  NAND U3501 ( .A(n2258), .B(n2257), .Z(n2362) );
  NANDN U3502 ( .A(n2260), .B(n2259), .Z(n2264) );
  NAND U3503 ( .A(n2262), .B(n2261), .Z(n2263) );
  NAND U3504 ( .A(n2264), .B(n2263), .Z(n2440) );
  XOR U3505 ( .A(b[7]), .B(a[17]), .Z(n2392) );
  NAND U3506 ( .A(n2392), .B(n36701), .Z(n2267) );
  NAND U3507 ( .A(n2265), .B(n36702), .Z(n2266) );
  NAND U3508 ( .A(n2267), .B(n2266), .Z(n2410) );
  XNOR U3509 ( .A(n1052), .B(a[15]), .Z(n2383) );
  NAND U3510 ( .A(n36925), .B(n2383), .Z(n2270) );
  NANDN U3511 ( .A(n2268), .B(n36926), .Z(n2269) );
  NAND U3512 ( .A(n2270), .B(n2269), .Z(n2407) );
  XNOR U3513 ( .A(b[5]), .B(a[19]), .Z(n2395) );
  NANDN U3514 ( .A(n2395), .B(n36587), .Z(n2273) );
  NANDN U3515 ( .A(n2271), .B(n36588), .Z(n2272) );
  AND U3516 ( .A(n2273), .B(n2272), .Z(n2408) );
  XNOR U3517 ( .A(n2407), .B(n2408), .Z(n2409) );
  XNOR U3518 ( .A(n2410), .B(n2409), .Z(n2438) );
  NANDN U3519 ( .A(n1049), .B(a[23]), .Z(n2274) );
  XNOR U3520 ( .A(b[1]), .B(n2274), .Z(n2276) );
  NANDN U3521 ( .A(b[0]), .B(a[22]), .Z(n2275) );
  AND U3522 ( .A(n2276), .B(n2275), .Z(n2419) );
  XOR U3523 ( .A(b[11]), .B(a[13]), .Z(n2377) );
  NANDN U3524 ( .A(n37311), .B(n2377), .Z(n2279) );
  NAND U3525 ( .A(n2277), .B(n37218), .Z(n2278) );
  AND U3526 ( .A(n2279), .B(n2278), .Z(n2420) );
  XNOR U3527 ( .A(n2419), .B(n2420), .Z(n2421) );
  XNOR U3528 ( .A(b[21]), .B(a[3]), .Z(n2374) );
  NANDN U3529 ( .A(n2374), .B(n38101), .Z(n2282) );
  NANDN U3530 ( .A(n2280), .B(n38102), .Z(n2281) );
  NAND U3531 ( .A(n2282), .B(n2281), .Z(n2423) );
  XNOR U3532 ( .A(n1057), .B(a[0]), .Z(n2285) );
  XNOR U3533 ( .A(n1057), .B(b[21]), .Z(n2284) );
  XNOR U3534 ( .A(n1057), .B(b[22]), .Z(n2283) );
  AND U3535 ( .A(n2284), .B(n2283), .Z(n38205) );
  NAND U3536 ( .A(n2285), .B(n38205), .Z(n2287) );
  XNOR U3537 ( .A(n1057), .B(a[1]), .Z(n2389) );
  ANDN U3538 ( .B(n2389), .A(n38268), .Z(n2286) );
  ANDN U3539 ( .B(n2287), .A(n2286), .Z(n2424) );
  XNOR U3540 ( .A(n2423), .B(n2424), .Z(n2422) );
  XOR U3541 ( .A(n2421), .B(n2422), .Z(n2437) );
  XNOR U3542 ( .A(n2438), .B(n2437), .Z(n2439) );
  XNOR U3543 ( .A(n2440), .B(n2439), .Z(n2434) );
  NANDN U3544 ( .A(n2289), .B(n2288), .Z(n2293) );
  NAND U3545 ( .A(n2291), .B(n2290), .Z(n2292) );
  NAND U3546 ( .A(n2293), .B(n2292), .Z(n2432) );
  NANDN U3547 ( .A(n2295), .B(n2294), .Z(n2299) );
  NAND U3548 ( .A(n2297), .B(n2296), .Z(n2298) );
  AND U3549 ( .A(n2299), .B(n2298), .Z(n2431) );
  XNOR U3550 ( .A(n2432), .B(n2431), .Z(n2433) );
  XNOR U3551 ( .A(n2434), .B(n2433), .Z(n2452) );
  NANDN U3552 ( .A(n2301), .B(n2300), .Z(n2305) );
  NANDN U3553 ( .A(n2303), .B(n2302), .Z(n2304) );
  NAND U3554 ( .A(n2305), .B(n2304), .Z(n2365) );
  NANDN U3555 ( .A(n2306), .B(n37762), .Z(n2308) );
  XOR U3556 ( .A(b[17]), .B(a[7]), .Z(n2398) );
  NAND U3557 ( .A(n2398), .B(n37764), .Z(n2307) );
  NAND U3558 ( .A(n2308), .B(n2307), .Z(n2416) );
  XNOR U3559 ( .A(n1055), .B(a[5]), .Z(n2386) );
  NAND U3560 ( .A(n2386), .B(n37934), .Z(n2311) );
  NANDN U3561 ( .A(n2309), .B(n37935), .Z(n2310) );
  NAND U3562 ( .A(n2311), .B(n2310), .Z(n2413) );
  XNOR U3563 ( .A(n1053), .B(a[11]), .Z(n2428) );
  NAND U3564 ( .A(n2428), .B(n37424), .Z(n2314) );
  NANDN U3565 ( .A(n2312), .B(n37425), .Z(n2313) );
  AND U3566 ( .A(n2314), .B(n2313), .Z(n2414) );
  XNOR U3567 ( .A(n2413), .B(n2414), .Z(n2415) );
  XOR U3568 ( .A(n2416), .B(n2415), .Z(n2366) );
  XNOR U3569 ( .A(n2365), .B(n2366), .Z(n2367) );
  XNOR U3570 ( .A(b[3]), .B(a[21]), .Z(n2425) );
  NANDN U3571 ( .A(n2425), .B(n36107), .Z(n2317) );
  OR U3572 ( .A(n2315), .B(n36105), .Z(n2316) );
  AND U3573 ( .A(n2317), .B(n2316), .Z(n2401) );
  XNOR U3574 ( .A(n2402), .B(n2401), .Z(n2403) );
  XNOR U3575 ( .A(n1054), .B(a[9]), .Z(n2380) );
  NANDN U3576 ( .A(n37665), .B(n2380), .Z(n2320) );
  NANDN U3577 ( .A(n2318), .B(n37604), .Z(n2319) );
  AND U3578 ( .A(n2320), .B(n2319), .Z(n2404) );
  XNOR U3579 ( .A(n2403), .B(n2404), .Z(n2368) );
  XOR U3580 ( .A(n2367), .B(n2368), .Z(n2449) );
  NANDN U3581 ( .A(n2322), .B(n2321), .Z(n2326) );
  NANDN U3582 ( .A(n2324), .B(n2323), .Z(n2325) );
  NAND U3583 ( .A(n2326), .B(n2325), .Z(n2450) );
  XNOR U3584 ( .A(n2449), .B(n2450), .Z(n2451) );
  XNOR U3585 ( .A(n2452), .B(n2451), .Z(n2359) );
  NANDN U3586 ( .A(n2328), .B(n2327), .Z(n2332) );
  OR U3587 ( .A(n2330), .B(n2329), .Z(n2331) );
  NAND U3588 ( .A(n2332), .B(n2331), .Z(n2446) );
  NANDN U3589 ( .A(n2334), .B(n2333), .Z(n2338) );
  NANDN U3590 ( .A(n2336), .B(n2335), .Z(n2337) );
  NAND U3591 ( .A(n2338), .B(n2337), .Z(n2443) );
  NANDN U3592 ( .A(n2340), .B(n2339), .Z(n2344) );
  NANDN U3593 ( .A(n2342), .B(n2341), .Z(n2343) );
  NAND U3594 ( .A(n2344), .B(n2343), .Z(n2444) );
  XNOR U3595 ( .A(n2443), .B(n2444), .Z(n2445) );
  XNOR U3596 ( .A(n2446), .B(n2445), .Z(n2360) );
  XOR U3597 ( .A(n2359), .B(n2360), .Z(n2361) );
  XOR U3598 ( .A(n2362), .B(n2361), .Z(n2355) );
  XNOR U3599 ( .A(n2356), .B(n2355), .Z(n2357) );
  XNOR U3600 ( .A(n2358), .B(n2357), .Z(n2350) );
  XNOR U3601 ( .A(n2350), .B(sreg[247]), .Z(n2352) );
  NAND U3602 ( .A(n2345), .B(sreg[246]), .Z(n2349) );
  OR U3603 ( .A(n2347), .B(n2346), .Z(n2348) );
  AND U3604 ( .A(n2349), .B(n2348), .Z(n2351) );
  XOR U3605 ( .A(n2352), .B(n2351), .Z(c[247]) );
  NAND U3606 ( .A(n2350), .B(sreg[247]), .Z(n2354) );
  OR U3607 ( .A(n2352), .B(n2351), .Z(n2353) );
  NAND U3608 ( .A(n2354), .B(n2353), .Z(n2568) );
  XNOR U3609 ( .A(n2568), .B(sreg[248]), .Z(n2570) );
  OR U3610 ( .A(n2360), .B(n2359), .Z(n2364) );
  NAND U3611 ( .A(n2362), .B(n2361), .Z(n2363) );
  NAND U3612 ( .A(n2364), .B(n2363), .Z(n2455) );
  NANDN U3613 ( .A(n2366), .B(n2365), .Z(n2370) );
  NANDN U3614 ( .A(n2368), .B(n2367), .Z(n2369) );
  NAND U3615 ( .A(n2370), .B(n2369), .Z(n2565) );
  NANDN U3616 ( .A(n1049), .B(a[24]), .Z(n2371) );
  XNOR U3617 ( .A(b[1]), .B(n2371), .Z(n2373) );
  NANDN U3618 ( .A(b[0]), .B(a[23]), .Z(n2372) );
  AND U3619 ( .A(n2373), .B(n2372), .Z(n2514) );
  XNOR U3620 ( .A(b[21]), .B(a[4]), .Z(n2488) );
  NANDN U3621 ( .A(n2488), .B(n38101), .Z(n2376) );
  NANDN U3622 ( .A(n2374), .B(n38102), .Z(n2375) );
  NAND U3623 ( .A(n2376), .B(n2375), .Z(n2512) );
  IV U3624 ( .A(b[24]), .Z(n38351) );
  XOR U3625 ( .A(n1057), .B(n38351), .Z(n38325) );
  NANDN U3626 ( .A(n3393), .B(n38325), .Z(n2513) );
  XNOR U3627 ( .A(n2512), .B(n2513), .Z(n2515) );
  XOR U3628 ( .A(n2514), .B(n2515), .Z(n2475) );
  XOR U3629 ( .A(b[11]), .B(a[14]), .Z(n2503) );
  NANDN U3630 ( .A(n37311), .B(n2503), .Z(n2379) );
  NAND U3631 ( .A(n2377), .B(n37218), .Z(n2378) );
  NAND U3632 ( .A(n2379), .B(n2378), .Z(n2479) );
  XNOR U3633 ( .A(b[15]), .B(a[10]), .Z(n2523) );
  OR U3634 ( .A(n2523), .B(n37665), .Z(n2382) );
  NAND U3635 ( .A(n2380), .B(n37604), .Z(n2381) );
  AND U3636 ( .A(n2382), .B(n2381), .Z(n2480) );
  XNOR U3637 ( .A(n2479), .B(n2480), .Z(n2481) );
  XNOR U3638 ( .A(b[9]), .B(a[16]), .Z(n2491) );
  NANDN U3639 ( .A(n2491), .B(n36925), .Z(n2385) );
  NAND U3640 ( .A(n36926), .B(n2383), .Z(n2384) );
  NAND U3641 ( .A(n2385), .B(n2384), .Z(n2548) );
  XOR U3642 ( .A(b[19]), .B(n4305), .Z(n2485) );
  NANDN U3643 ( .A(n2485), .B(n37934), .Z(n2388) );
  NAND U3644 ( .A(n37935), .B(n2386), .Z(n2387) );
  NAND U3645 ( .A(n2388), .B(n2387), .Z(n2546) );
  NAND U3646 ( .A(n2389), .B(n38205), .Z(n2391) );
  XNOR U3647 ( .A(b[23]), .B(a[2]), .Z(n2532) );
  OR U3648 ( .A(n2532), .B(n38268), .Z(n2390) );
  AND U3649 ( .A(n2391), .B(n2390), .Z(n2547) );
  XNOR U3650 ( .A(n2546), .B(n2547), .Z(n2549) );
  XNOR U3651 ( .A(n2548), .B(n2549), .Z(n2482) );
  XNOR U3652 ( .A(n2481), .B(n2482), .Z(n2473) );
  XOR U3653 ( .A(b[7]), .B(a[18]), .Z(n2494) );
  NAND U3654 ( .A(n2494), .B(n36701), .Z(n2394) );
  NAND U3655 ( .A(n2392), .B(n36702), .Z(n2393) );
  NAND U3656 ( .A(n2394), .B(n2393), .Z(n2509) );
  XNOR U3657 ( .A(b[5]), .B(a[20]), .Z(n2497) );
  NANDN U3658 ( .A(n2497), .B(n36587), .Z(n2397) );
  NANDN U3659 ( .A(n2395), .B(n36588), .Z(n2396) );
  NAND U3660 ( .A(n2397), .B(n2396), .Z(n2506) );
  NAND U3661 ( .A(n2398), .B(n37762), .Z(n2400) );
  XOR U3662 ( .A(b[17]), .B(a[8]), .Z(n2500) );
  NAND U3663 ( .A(n2500), .B(n37764), .Z(n2399) );
  AND U3664 ( .A(n2400), .B(n2399), .Z(n2507) );
  XNOR U3665 ( .A(n2506), .B(n2507), .Z(n2508) );
  XOR U3666 ( .A(n2509), .B(n2508), .Z(n2474) );
  XNOR U3667 ( .A(n2473), .B(n2474), .Z(n2476) );
  XNOR U3668 ( .A(n2475), .B(n2476), .Z(n2553) );
  NANDN U3669 ( .A(n2402), .B(n2401), .Z(n2406) );
  NAND U3670 ( .A(n2404), .B(n2403), .Z(n2405) );
  NAND U3671 ( .A(n2406), .B(n2405), .Z(n2550) );
  NANDN U3672 ( .A(n2408), .B(n2407), .Z(n2412) );
  NAND U3673 ( .A(n2410), .B(n2409), .Z(n2411) );
  NAND U3674 ( .A(n2412), .B(n2411), .Z(n2551) );
  XNOR U3675 ( .A(n2550), .B(n2551), .Z(n2552) );
  XOR U3676 ( .A(n2553), .B(n2552), .Z(n2470) );
  NANDN U3677 ( .A(n2414), .B(n2413), .Z(n2418) );
  NAND U3678 ( .A(n2416), .B(n2415), .Z(n2417) );
  NAND U3679 ( .A(n2418), .B(n2417), .Z(n2557) );
  XNOR U3680 ( .A(n2557), .B(n2556), .Z(n2558) );
  NANDN U3681 ( .A(n2424), .B(n2423), .Z(n2543) );
  XNOR U3682 ( .A(b[3]), .B(a[22]), .Z(n2520) );
  NANDN U3683 ( .A(n2520), .B(n36107), .Z(n2427) );
  OR U3684 ( .A(n2425), .B(n36105), .Z(n2426) );
  NAND U3685 ( .A(n2427), .B(n2426), .Z(n2541) );
  XNOR U3686 ( .A(b[13]), .B(a[12]), .Z(n2529) );
  NANDN U3687 ( .A(n2529), .B(n37424), .Z(n2430) );
  NAND U3688 ( .A(n37425), .B(n2428), .Z(n2429) );
  AND U3689 ( .A(n2430), .B(n2429), .Z(n2540) );
  XNOR U3690 ( .A(n2541), .B(n2540), .Z(n2542) );
  XNOR U3691 ( .A(n2543), .B(n2542), .Z(n2559) );
  XOR U3692 ( .A(n2558), .B(n2559), .Z(n2467) );
  NANDN U3693 ( .A(n2432), .B(n2431), .Z(n2436) );
  NANDN U3694 ( .A(n2434), .B(n2433), .Z(n2435) );
  NAND U3695 ( .A(n2436), .B(n2435), .Z(n2468) );
  XNOR U3696 ( .A(n2467), .B(n2468), .Z(n2469) );
  XNOR U3697 ( .A(n2470), .B(n2469), .Z(n2562) );
  NANDN U3698 ( .A(n2438), .B(n2437), .Z(n2442) );
  NANDN U3699 ( .A(n2440), .B(n2439), .Z(n2441) );
  NAND U3700 ( .A(n2442), .B(n2441), .Z(n2563) );
  XNOR U3701 ( .A(n2562), .B(n2563), .Z(n2564) );
  XNOR U3702 ( .A(n2565), .B(n2564), .Z(n2464) );
  NANDN U3703 ( .A(n2444), .B(n2443), .Z(n2448) );
  NAND U3704 ( .A(n2446), .B(n2445), .Z(n2447) );
  NAND U3705 ( .A(n2448), .B(n2447), .Z(n2461) );
  NANDN U3706 ( .A(n2450), .B(n2449), .Z(n2454) );
  NANDN U3707 ( .A(n2452), .B(n2451), .Z(n2453) );
  NAND U3708 ( .A(n2454), .B(n2453), .Z(n2462) );
  XNOR U3709 ( .A(n2461), .B(n2462), .Z(n2463) );
  XOR U3710 ( .A(n2464), .B(n2463), .Z(n2456) );
  XNOR U3711 ( .A(n2455), .B(n2456), .Z(n2457) );
  XOR U3712 ( .A(n2458), .B(n2457), .Z(n2569) );
  XOR U3713 ( .A(n2570), .B(n2569), .Z(c[248]) );
  NANDN U3714 ( .A(n2456), .B(n2455), .Z(n2460) );
  NAND U3715 ( .A(n2458), .B(n2457), .Z(n2459) );
  NAND U3716 ( .A(n2460), .B(n2459), .Z(n2581) );
  NANDN U3717 ( .A(n2462), .B(n2461), .Z(n2466) );
  NANDN U3718 ( .A(n2464), .B(n2463), .Z(n2465) );
  NAND U3719 ( .A(n2466), .B(n2465), .Z(n2578) );
  NANDN U3720 ( .A(n2468), .B(n2467), .Z(n2472) );
  NAND U3721 ( .A(n2470), .B(n2469), .Z(n2471) );
  NAND U3722 ( .A(n2472), .B(n2471), .Z(n2585) );
  OR U3723 ( .A(n2474), .B(n2473), .Z(n2478) );
  OR U3724 ( .A(n2476), .B(n2475), .Z(n2477) );
  AND U3725 ( .A(n2478), .B(n2477), .Z(n2590) );
  NANDN U3726 ( .A(n2480), .B(n2479), .Z(n2484) );
  NANDN U3727 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U3728 ( .A(n2484), .B(n2483), .Z(n2686) );
  XNOR U3729 ( .A(b[19]), .B(a[7]), .Z(n2628) );
  NANDN U3730 ( .A(n2628), .B(n37934), .Z(n2487) );
  NANDN U3731 ( .A(n2485), .B(n37935), .Z(n2486) );
  NAND U3732 ( .A(n2487), .B(n2486), .Z(n2634) );
  XNOR U3733 ( .A(b[21]), .B(a[5]), .Z(n2661) );
  NANDN U3734 ( .A(n2661), .B(n38101), .Z(n2490) );
  NANDN U3735 ( .A(n2488), .B(n38102), .Z(n2489) );
  NAND U3736 ( .A(n2490), .B(n2489), .Z(n2631) );
  XNOR U3737 ( .A(b[9]), .B(a[17]), .Z(n2640) );
  NANDN U3738 ( .A(n2640), .B(n36925), .Z(n2493) );
  NANDN U3739 ( .A(n2491), .B(n36926), .Z(n2492) );
  AND U3740 ( .A(n2493), .B(n2492), .Z(n2632) );
  XNOR U3741 ( .A(n2631), .B(n2632), .Z(n2633) );
  XNOR U3742 ( .A(n2634), .B(n2633), .Z(n2605) );
  XOR U3743 ( .A(b[7]), .B(a[19]), .Z(n2637) );
  NAND U3744 ( .A(n2637), .B(n36701), .Z(n2496) );
  NAND U3745 ( .A(n2494), .B(n36702), .Z(n2495) );
  NAND U3746 ( .A(n2496), .B(n2495), .Z(n2611) );
  XNOR U3747 ( .A(b[5]), .B(a[21]), .Z(n2622) );
  NANDN U3748 ( .A(n2622), .B(n36587), .Z(n2499) );
  NANDN U3749 ( .A(n2497), .B(n36588), .Z(n2498) );
  NAND U3750 ( .A(n2499), .B(n2498), .Z(n2608) );
  NAND U3751 ( .A(n2500), .B(n37762), .Z(n2502) );
  XOR U3752 ( .A(b[17]), .B(a[9]), .Z(n2658) );
  NAND U3753 ( .A(n2658), .B(n37764), .Z(n2501) );
  AND U3754 ( .A(n2502), .B(n2501), .Z(n2609) );
  XNOR U3755 ( .A(n2608), .B(n2609), .Z(n2610) );
  XNOR U3756 ( .A(n2611), .B(n2610), .Z(n2602) );
  XOR U3757 ( .A(b[11]), .B(a[15]), .Z(n2643) );
  NANDN U3758 ( .A(n37311), .B(n2643), .Z(n2505) );
  NAND U3759 ( .A(n37218), .B(n2503), .Z(n2504) );
  NAND U3760 ( .A(n2505), .B(n2504), .Z(n2603) );
  XNOR U3761 ( .A(n2602), .B(n2603), .Z(n2604) );
  XOR U3762 ( .A(n2605), .B(n2604), .Z(n2684) );
  NANDN U3763 ( .A(n2507), .B(n2506), .Z(n2511) );
  NAND U3764 ( .A(n2509), .B(n2508), .Z(n2510) );
  AND U3765 ( .A(n2511), .B(n2510), .Z(n2683) );
  XOR U3766 ( .A(n2684), .B(n2683), .Z(n2685) );
  XOR U3767 ( .A(n2686), .B(n2685), .Z(n2591) );
  XOR U3768 ( .A(n2590), .B(n2591), .Z(n2593) );
  NANDN U3769 ( .A(n2513), .B(n2512), .Z(n2517) );
  NAND U3770 ( .A(n2515), .B(n2514), .Z(n2516) );
  NAND U3771 ( .A(n2517), .B(n2516), .Z(n2674) );
  NANDN U3772 ( .A(n1057), .B(b[24]), .Z(n38350) );
  AND U3773 ( .A(n38350), .B(b[25]), .Z(n38456) );
  XNOR U3774 ( .A(n38351), .B(b[23]), .Z(n2518) );
  NANDN U3775 ( .A(n3393), .B(n2518), .Z(n2519) );
  AND U3776 ( .A(n38456), .B(n2519), .Z(n2653) );
  XNOR U3777 ( .A(b[3]), .B(a[23]), .Z(n2619) );
  NANDN U3778 ( .A(n2619), .B(n36107), .Z(n2522) );
  OR U3779 ( .A(n2520), .B(n36105), .Z(n2521) );
  AND U3780 ( .A(n2522), .B(n2521), .Z(n2652) );
  XNOR U3781 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3782 ( .A(b[15]), .B(a[11]), .Z(n2616) );
  OR U3783 ( .A(n2616), .B(n37665), .Z(n2525) );
  NANDN U3784 ( .A(n2523), .B(n37604), .Z(n2524) );
  NAND U3785 ( .A(n2525), .B(n2524), .Z(n2655) );
  XOR U3786 ( .A(n2654), .B(n2655), .Z(n2672) );
  NANDN U3787 ( .A(n1049), .B(a[25]), .Z(n2526) );
  XNOR U3788 ( .A(b[1]), .B(n2526), .Z(n2528) );
  NANDN U3789 ( .A(b[0]), .B(a[24]), .Z(n2527) );
  AND U3790 ( .A(n2528), .B(n2527), .Z(n2667) );
  XNOR U3791 ( .A(b[13]), .B(a[13]), .Z(n2625) );
  NANDN U3792 ( .A(n2625), .B(n37424), .Z(n2531) );
  NANDN U3793 ( .A(n2529), .B(n37425), .Z(n2530) );
  AND U3794 ( .A(n2531), .B(n2530), .Z(n2668) );
  XNOR U3795 ( .A(n2667), .B(n2668), .Z(n2669) );
  NANDN U3796 ( .A(n2532), .B(n38205), .Z(n2534) );
  XNOR U3797 ( .A(b[23]), .B(a[3]), .Z(n2649) );
  OR U3798 ( .A(n2649), .B(n38268), .Z(n2533) );
  NAND U3799 ( .A(n2534), .B(n2533), .Z(n2614) );
  XNOR U3800 ( .A(b[25]), .B(n3393), .Z(n2537) );
  XNOR U3801 ( .A(b[25]), .B(n1057), .Z(n2536) );
  XNOR U3802 ( .A(b[25]), .B(n38351), .Z(n2535) );
  AND U3803 ( .A(n2536), .B(n2535), .Z(n38326) );
  NAND U3804 ( .A(n2537), .B(n38326), .Z(n2539) );
  XOR U3805 ( .A(b[25]), .B(a[1]), .Z(n2664) );
  AND U3806 ( .A(n38325), .B(n2664), .Z(n2538) );
  ANDN U3807 ( .B(n2539), .A(n2538), .Z(n2615) );
  XNOR U3808 ( .A(n2614), .B(n2615), .Z(n2670) );
  XOR U3809 ( .A(n2669), .B(n2670), .Z(n2671) );
  XOR U3810 ( .A(n2672), .B(n2671), .Z(n2673) );
  XNOR U3811 ( .A(n2674), .B(n2673), .Z(n2680) );
  NANDN U3812 ( .A(n2541), .B(n2540), .Z(n2545) );
  NAND U3813 ( .A(n2543), .B(n2542), .Z(n2544) );
  NAND U3814 ( .A(n2545), .B(n2544), .Z(n2677) );
  XNOR U3815 ( .A(n2677), .B(n2678), .Z(n2679) );
  XOR U3816 ( .A(n2680), .B(n2679), .Z(n2592) );
  XOR U3817 ( .A(n2593), .B(n2592), .Z(n2599) );
  NANDN U3818 ( .A(n2551), .B(n2550), .Z(n2555) );
  NANDN U3819 ( .A(n2553), .B(n2552), .Z(n2554) );
  NAND U3820 ( .A(n2555), .B(n2554), .Z(n2597) );
  NANDN U3821 ( .A(n2557), .B(n2556), .Z(n2561) );
  NANDN U3822 ( .A(n2559), .B(n2558), .Z(n2560) );
  AND U3823 ( .A(n2561), .B(n2560), .Z(n2596) );
  XNOR U3824 ( .A(n2597), .B(n2596), .Z(n2598) );
  XNOR U3825 ( .A(n2599), .B(n2598), .Z(n2584) );
  XNOR U3826 ( .A(n2585), .B(n2584), .Z(n2587) );
  NANDN U3827 ( .A(n2563), .B(n2562), .Z(n2567) );
  NAND U3828 ( .A(n2565), .B(n2564), .Z(n2566) );
  NAND U3829 ( .A(n2567), .B(n2566), .Z(n2586) );
  XOR U3830 ( .A(n2587), .B(n2586), .Z(n2579) );
  XNOR U3831 ( .A(n2578), .B(n2579), .Z(n2580) );
  XNOR U3832 ( .A(n2581), .B(n2580), .Z(n2573) );
  XNOR U3833 ( .A(n2573), .B(sreg[249]), .Z(n2575) );
  NAND U3834 ( .A(n2568), .B(sreg[248]), .Z(n2572) );
  OR U3835 ( .A(n2570), .B(n2569), .Z(n2571) );
  AND U3836 ( .A(n2572), .B(n2571), .Z(n2574) );
  XOR U3837 ( .A(n2575), .B(n2574), .Z(c[249]) );
  NAND U3838 ( .A(n2573), .B(sreg[249]), .Z(n2577) );
  OR U3839 ( .A(n2575), .B(n2574), .Z(n2576) );
  NAND U3840 ( .A(n2577), .B(n2576), .Z(n2808) );
  XNOR U3841 ( .A(n2808), .B(sreg[250]), .Z(n2810) );
  NANDN U3842 ( .A(n2579), .B(n2578), .Z(n2583) );
  NAND U3843 ( .A(n2581), .B(n2580), .Z(n2582) );
  NAND U3844 ( .A(n2583), .B(n2582), .Z(n2692) );
  NAND U3845 ( .A(n2585), .B(n2584), .Z(n2589) );
  OR U3846 ( .A(n2587), .B(n2586), .Z(n2588) );
  NAND U3847 ( .A(n2589), .B(n2588), .Z(n2690) );
  OR U3848 ( .A(n2591), .B(n2590), .Z(n2595) );
  NAND U3849 ( .A(n2593), .B(n2592), .Z(n2594) );
  NAND U3850 ( .A(n2595), .B(n2594), .Z(n2698) );
  NANDN U3851 ( .A(n2597), .B(n2596), .Z(n2601) );
  NANDN U3852 ( .A(n2599), .B(n2598), .Z(n2600) );
  NAND U3853 ( .A(n2601), .B(n2600), .Z(n2695) );
  NANDN U3854 ( .A(n2603), .B(n2602), .Z(n2607) );
  NAND U3855 ( .A(n2605), .B(n2604), .Z(n2606) );
  AND U3856 ( .A(n2607), .B(n2606), .Z(n2707) );
  NANDN U3857 ( .A(n2609), .B(n2608), .Z(n2613) );
  NAND U3858 ( .A(n2611), .B(n2610), .Z(n2612) );
  NAND U3859 ( .A(n2613), .B(n2612), .Z(n2732) );
  NANDN U3860 ( .A(n2615), .B(n2614), .Z(n2794) );
  XNOR U3861 ( .A(n1054), .B(a[12]), .Z(n2766) );
  NANDN U3862 ( .A(n37665), .B(n2766), .Z(n2618) );
  NANDN U3863 ( .A(n2616), .B(n37604), .Z(n2617) );
  NAND U3864 ( .A(n2618), .B(n2617), .Z(n2793) );
  XNOR U3865 ( .A(b[3]), .B(a[24]), .Z(n2763) );
  NANDN U3866 ( .A(n2763), .B(n36107), .Z(n2621) );
  OR U3867 ( .A(n2619), .B(n36105), .Z(n2620) );
  AND U3868 ( .A(n2621), .B(n2620), .Z(n2792) );
  XNOR U3869 ( .A(n2793), .B(n2792), .Z(n2795) );
  XNOR U3870 ( .A(n2794), .B(n2795), .Z(n2729) );
  XNOR U3871 ( .A(b[5]), .B(a[22]), .Z(n2786) );
  NANDN U3872 ( .A(n2786), .B(n36587), .Z(n2624) );
  NANDN U3873 ( .A(n2622), .B(n36588), .Z(n2623) );
  NAND U3874 ( .A(n2624), .B(n2623), .Z(n2738) );
  XNOR U3875 ( .A(n1053), .B(a[14]), .Z(n2780) );
  NAND U3876 ( .A(n2780), .B(n37424), .Z(n2627) );
  NANDN U3877 ( .A(n2625), .B(n37425), .Z(n2626) );
  NAND U3878 ( .A(n2627), .B(n2626), .Z(n2735) );
  XNOR U3879 ( .A(b[19]), .B(a[8]), .Z(n2789) );
  NANDN U3880 ( .A(n2789), .B(n37934), .Z(n2630) );
  NANDN U3881 ( .A(n2628), .B(n37935), .Z(n2629) );
  AND U3882 ( .A(n2630), .B(n2629), .Z(n2736) );
  XNOR U3883 ( .A(n2735), .B(n2736), .Z(n2737) );
  XNOR U3884 ( .A(n2738), .B(n2737), .Z(n2730) );
  XNOR U3885 ( .A(n2729), .B(n2730), .Z(n2731) );
  XOR U3886 ( .A(n2732), .B(n2731), .Z(n2708) );
  XOR U3887 ( .A(n2707), .B(n2708), .Z(n2710) );
  NANDN U3888 ( .A(n2632), .B(n2631), .Z(n2636) );
  NAND U3889 ( .A(n2634), .B(n2633), .Z(n2635) );
  NAND U3890 ( .A(n2636), .B(n2635), .Z(n2725) );
  XOR U3891 ( .A(b[7]), .B(a[20]), .Z(n2783) );
  NAND U3892 ( .A(n2783), .B(n36701), .Z(n2639) );
  NAND U3893 ( .A(n2637), .B(n36702), .Z(n2638) );
  NAND U3894 ( .A(n2639), .B(n2638), .Z(n2799) );
  XNOR U3895 ( .A(b[9]), .B(a[18]), .Z(n2747) );
  NANDN U3896 ( .A(n2747), .B(n36925), .Z(n2642) );
  NANDN U3897 ( .A(n2640), .B(n36926), .Z(n2641) );
  NAND U3898 ( .A(n2642), .B(n2641), .Z(n2796) );
  XOR U3899 ( .A(b[11]), .B(a[16]), .Z(n2744) );
  NANDN U3900 ( .A(n37311), .B(n2744), .Z(n2645) );
  NAND U3901 ( .A(n2643), .B(n37218), .Z(n2644) );
  AND U3902 ( .A(n2645), .B(n2644), .Z(n2797) );
  XNOR U3903 ( .A(n2796), .B(n2797), .Z(n2798) );
  XNOR U3904 ( .A(n2799), .B(n2798), .Z(n2723) );
  XOR U3905 ( .A(b[26]), .B(b[25]), .Z(n38423) );
  NAND U3906 ( .A(a[0]), .B(n38423), .Z(n2759) );
  NANDN U3907 ( .A(n1049), .B(a[26]), .Z(n2646) );
  XNOR U3908 ( .A(b[1]), .B(n2646), .Z(n2648) );
  IV U3909 ( .A(a[25]), .Z(n7069) );
  NANDN U3910 ( .A(n7069), .B(n1049), .Z(n2647) );
  AND U3911 ( .A(n2648), .B(n2647), .Z(n2757) );
  XNOR U3912 ( .A(b[23]), .B(a[4]), .Z(n2753) );
  OR U3913 ( .A(n2753), .B(n38268), .Z(n2651) );
  NANDN U3914 ( .A(n2649), .B(n38205), .Z(n2650) );
  AND U3915 ( .A(n2651), .B(n2650), .Z(n2756) );
  XNOR U3916 ( .A(n2757), .B(n2756), .Z(n2758) );
  XNOR U3917 ( .A(n2759), .B(n2758), .Z(n2724) );
  XOR U3918 ( .A(n2723), .B(n2724), .Z(n2726) );
  XOR U3919 ( .A(n2725), .B(n2726), .Z(n2709) );
  XOR U3920 ( .A(n2710), .B(n2709), .Z(n2715) );
  NANDN U3921 ( .A(n2653), .B(n2652), .Z(n2657) );
  NANDN U3922 ( .A(n2655), .B(n2654), .Z(n2656) );
  NAND U3923 ( .A(n2657), .B(n2656), .Z(n2722) );
  NAND U3924 ( .A(n2658), .B(n37762), .Z(n2660) );
  XOR U3925 ( .A(b[17]), .B(a[10]), .Z(n2741) );
  NAND U3926 ( .A(n2741), .B(n37764), .Z(n2659) );
  NAND U3927 ( .A(n2660), .B(n2659), .Z(n2805) );
  XOR U3928 ( .A(b[21]), .B(n4305), .Z(n2750) );
  NANDN U3929 ( .A(n2750), .B(n38101), .Z(n2663) );
  NANDN U3930 ( .A(n2661), .B(n38102), .Z(n2662) );
  NAND U3931 ( .A(n2663), .B(n2662), .Z(n2802) );
  XOR U3932 ( .A(b[25]), .B(a[2]), .Z(n2769) );
  NAND U3933 ( .A(n2769), .B(n38325), .Z(n2666) );
  NAND U3934 ( .A(n2664), .B(n38326), .Z(n2665) );
  AND U3935 ( .A(n2666), .B(n2665), .Z(n2803) );
  XNOR U3936 ( .A(n2802), .B(n2803), .Z(n2804) );
  XNOR U3937 ( .A(n2805), .B(n2804), .Z(n2719) );
  XNOR U3938 ( .A(n2719), .B(n2720), .Z(n2721) );
  XNOR U3939 ( .A(n2722), .B(n2721), .Z(n2713) );
  NAND U3940 ( .A(n2672), .B(n2671), .Z(n2676) );
  NAND U3941 ( .A(n2674), .B(n2673), .Z(n2675) );
  AND U3942 ( .A(n2676), .B(n2675), .Z(n2714) );
  XOR U3943 ( .A(n2713), .B(n2714), .Z(n2716) );
  XOR U3944 ( .A(n2715), .B(n2716), .Z(n2704) );
  NANDN U3945 ( .A(n2678), .B(n2677), .Z(n2682) );
  NAND U3946 ( .A(n2680), .B(n2679), .Z(n2681) );
  NAND U3947 ( .A(n2682), .B(n2681), .Z(n2701) );
  OR U3948 ( .A(n2684), .B(n2683), .Z(n2688) );
  NAND U3949 ( .A(n2686), .B(n2685), .Z(n2687) );
  NAND U3950 ( .A(n2688), .B(n2687), .Z(n2702) );
  XNOR U3951 ( .A(n2701), .B(n2702), .Z(n2703) );
  XOR U3952 ( .A(n2704), .B(n2703), .Z(n2696) );
  XOR U3953 ( .A(n2695), .B(n2696), .Z(n2697) );
  XOR U3954 ( .A(n2698), .B(n2697), .Z(n2689) );
  XNOR U3955 ( .A(n2690), .B(n2689), .Z(n2691) );
  XOR U3956 ( .A(n2692), .B(n2691), .Z(n2809) );
  XOR U3957 ( .A(n2810), .B(n2809), .Z(c[250]) );
  NANDN U3958 ( .A(n2690), .B(n2689), .Z(n2694) );
  NAND U3959 ( .A(n2692), .B(n2691), .Z(n2693) );
  NAND U3960 ( .A(n2694), .B(n2693), .Z(n2821) );
  OR U3961 ( .A(n2696), .B(n2695), .Z(n2700) );
  NAND U3962 ( .A(n2698), .B(n2697), .Z(n2699) );
  NAND U3963 ( .A(n2700), .B(n2699), .Z(n2818) );
  NANDN U3964 ( .A(n2702), .B(n2701), .Z(n2706) );
  NANDN U3965 ( .A(n2704), .B(n2703), .Z(n2705) );
  NAND U3966 ( .A(n2706), .B(n2705), .Z(n2827) );
  OR U3967 ( .A(n2708), .B(n2707), .Z(n2712) );
  NAND U3968 ( .A(n2710), .B(n2709), .Z(n2711) );
  NAND U3969 ( .A(n2712), .B(n2711), .Z(n2824) );
  NANDN U3970 ( .A(n2714), .B(n2713), .Z(n2718) );
  OR U3971 ( .A(n2716), .B(n2715), .Z(n2717) );
  NAND U3972 ( .A(n2718), .B(n2717), .Z(n2935) );
  NANDN U3973 ( .A(n2724), .B(n2723), .Z(n2728) );
  OR U3974 ( .A(n2726), .B(n2725), .Z(n2727) );
  NAND U3975 ( .A(n2728), .B(n2727), .Z(n2916) );
  NANDN U3976 ( .A(n2730), .B(n2729), .Z(n2734) );
  NAND U3977 ( .A(n2732), .B(n2731), .Z(n2733) );
  NAND U3978 ( .A(n2734), .B(n2733), .Z(n2917) );
  XNOR U3979 ( .A(n2916), .B(n2917), .Z(n2918) );
  XNOR U3980 ( .A(n2919), .B(n2918), .Z(n2932) );
  NANDN U3981 ( .A(n2736), .B(n2735), .Z(n2740) );
  NAND U3982 ( .A(n2738), .B(n2737), .Z(n2739) );
  NAND U3983 ( .A(n2740), .B(n2739), .Z(n2923) );
  NAND U3984 ( .A(n2741), .B(n37762), .Z(n2743) );
  XOR U3985 ( .A(b[17]), .B(a[11]), .Z(n2872) );
  NAND U3986 ( .A(n2872), .B(n37764), .Z(n2742) );
  NAND U3987 ( .A(n2743), .B(n2742), .Z(n2878) );
  XOR U3988 ( .A(b[11]), .B(a[17]), .Z(n2869) );
  NANDN U3989 ( .A(n37311), .B(n2869), .Z(n2746) );
  NAND U3990 ( .A(n2744), .B(n37218), .Z(n2745) );
  AND U3991 ( .A(n2746), .B(n2745), .Z(n2879) );
  XNOR U3992 ( .A(n2878), .B(n2879), .Z(n2880) );
  XNOR U3993 ( .A(b[9]), .B(a[19]), .Z(n2875) );
  NANDN U3994 ( .A(n2875), .B(n36925), .Z(n2749) );
  NANDN U3995 ( .A(n2747), .B(n36926), .Z(n2748) );
  NAND U3996 ( .A(n2749), .B(n2748), .Z(n2839) );
  XNOR U3997 ( .A(b[21]), .B(a[7]), .Z(n2863) );
  NANDN U3998 ( .A(n2863), .B(n38101), .Z(n2752) );
  NANDN U3999 ( .A(n2750), .B(n38102), .Z(n2751) );
  NAND U4000 ( .A(n2752), .B(n2751), .Z(n2836) );
  NANDN U4001 ( .A(n2753), .B(n38205), .Z(n2755) );
  XNOR U4002 ( .A(b[23]), .B(a[5]), .Z(n2854) );
  OR U4003 ( .A(n2854), .B(n38268), .Z(n2754) );
  AND U4004 ( .A(n2755), .B(n2754), .Z(n2837) );
  XNOR U4005 ( .A(n2836), .B(n2837), .Z(n2838) );
  XNOR U4006 ( .A(n2839), .B(n2838), .Z(n2881) );
  XOR U4007 ( .A(n2880), .B(n2881), .Z(n2913) );
  NANDN U4008 ( .A(n2757), .B(n2756), .Z(n2761) );
  NAND U4009 ( .A(n2759), .B(n2758), .Z(n2760) );
  NAND U4010 ( .A(n2761), .B(n2760), .Z(n2910) );
  NAND U4011 ( .A(b[26]), .B(b[25]), .Z(n38444) );
  AND U4012 ( .A(n38444), .B(b[27]), .Z(n38522) );
  NANDN U4013 ( .A(n3393), .B(n38423), .Z(n2762) );
  AND U4014 ( .A(n38522), .B(n2762), .Z(n2907) );
  OR U4015 ( .A(n2763), .B(n36105), .Z(n2765) );
  XOR U4016 ( .A(b[3]), .B(n7069), .Z(n2851) );
  NANDN U4017 ( .A(n2851), .B(n36107), .Z(n2764) );
  NAND U4018 ( .A(n2765), .B(n2764), .Z(n2904) );
  XNOR U4019 ( .A(b[15]), .B(a[13]), .Z(n2899) );
  OR U4020 ( .A(n2899), .B(n37665), .Z(n2768) );
  NAND U4021 ( .A(n2766), .B(n37604), .Z(n2767) );
  AND U4022 ( .A(n2768), .B(n2767), .Z(n2905) );
  XNOR U4023 ( .A(n2904), .B(n2905), .Z(n2906) );
  XOR U4024 ( .A(n2907), .B(n2906), .Z(n2911) );
  XNOR U4025 ( .A(n2910), .B(n2911), .Z(n2912) );
  XOR U4026 ( .A(n2913), .B(n2912), .Z(n2922) );
  XOR U4027 ( .A(n2923), .B(n2922), .Z(n2925) );
  XOR U4028 ( .A(b[25]), .B(a[3]), .Z(n2893) );
  NAND U4029 ( .A(n2893), .B(n38325), .Z(n2771) );
  NAND U4030 ( .A(n2769), .B(n38326), .Z(n2770) );
  NAND U4031 ( .A(n2771), .B(n2770), .Z(n2903) );
  XOR U4032 ( .A(b[27]), .B(a[1]), .Z(n2896) );
  AND U4033 ( .A(n2896), .B(n38423), .Z(n2776) );
  XNOR U4034 ( .A(b[27]), .B(n3393), .Z(n2774) );
  XOR U4035 ( .A(b[27]), .B(b[25]), .Z(n2773) );
  XOR U4036 ( .A(b[27]), .B(b[26]), .Z(n2772) );
  AND U4037 ( .A(n2773), .B(n2772), .Z(n38424) );
  NAND U4038 ( .A(n2774), .B(n38424), .Z(n2775) );
  NANDN U4039 ( .A(n2776), .B(n2775), .Z(n2902) );
  XNOR U4040 ( .A(n2903), .B(n2902), .Z(n2845) );
  NANDN U4041 ( .A(n1049), .B(a[27]), .Z(n2777) );
  XNOR U4042 ( .A(b[1]), .B(n2777), .Z(n2779) );
  IV U4043 ( .A(a[26]), .Z(n7202) );
  NANDN U4044 ( .A(n7202), .B(n1049), .Z(n2778) );
  AND U4045 ( .A(n2779), .B(n2778), .Z(n2843) );
  XNOR U4046 ( .A(b[13]), .B(a[15]), .Z(n2848) );
  NANDN U4047 ( .A(n2848), .B(n37424), .Z(n2782) );
  NAND U4048 ( .A(n37425), .B(n2780), .Z(n2781) );
  AND U4049 ( .A(n2782), .B(n2781), .Z(n2842) );
  XNOR U4050 ( .A(n2843), .B(n2842), .Z(n2844) );
  XOR U4051 ( .A(n2845), .B(n2844), .Z(n2830) );
  XOR U4052 ( .A(b[7]), .B(a[21]), .Z(n2866) );
  NAND U4053 ( .A(n2866), .B(n36701), .Z(n2785) );
  NAND U4054 ( .A(n2783), .B(n36702), .Z(n2784) );
  NAND U4055 ( .A(n2785), .B(n2784), .Z(n2887) );
  XNOR U4056 ( .A(b[5]), .B(a[23]), .Z(n2857) );
  NANDN U4057 ( .A(n2857), .B(n36587), .Z(n2788) );
  NANDN U4058 ( .A(n2786), .B(n36588), .Z(n2787) );
  NAND U4059 ( .A(n2788), .B(n2787), .Z(n2884) );
  XNOR U4060 ( .A(b[19]), .B(a[9]), .Z(n2860) );
  NANDN U4061 ( .A(n2860), .B(n37934), .Z(n2791) );
  NANDN U4062 ( .A(n2789), .B(n37935), .Z(n2790) );
  AND U4063 ( .A(n2791), .B(n2790), .Z(n2885) );
  XNOR U4064 ( .A(n2884), .B(n2885), .Z(n2886) );
  XNOR U4065 ( .A(n2887), .B(n2886), .Z(n2831) );
  XOR U4066 ( .A(n2830), .B(n2831), .Z(n2832) );
  XOR U4067 ( .A(n2832), .B(n2833), .Z(n2931) );
  NANDN U4068 ( .A(n2797), .B(n2796), .Z(n2801) );
  NAND U4069 ( .A(n2799), .B(n2798), .Z(n2800) );
  NAND U4070 ( .A(n2801), .B(n2800), .Z(n2929) );
  NANDN U4071 ( .A(n2803), .B(n2802), .Z(n2807) );
  NAND U4072 ( .A(n2805), .B(n2804), .Z(n2806) );
  AND U4073 ( .A(n2807), .B(n2806), .Z(n2928) );
  XNOR U4074 ( .A(n2929), .B(n2928), .Z(n2930) );
  XOR U4075 ( .A(n2931), .B(n2930), .Z(n2924) );
  XOR U4076 ( .A(n2925), .B(n2924), .Z(n2933) );
  XNOR U4077 ( .A(n2932), .B(n2933), .Z(n2934) );
  XOR U4078 ( .A(n2935), .B(n2934), .Z(n2825) );
  XNOR U4079 ( .A(n2824), .B(n2825), .Z(n2826) );
  XNOR U4080 ( .A(n2827), .B(n2826), .Z(n2819) );
  XNOR U4081 ( .A(n2818), .B(n2819), .Z(n2820) );
  XNOR U4082 ( .A(n2821), .B(n2820), .Z(n2813) );
  XNOR U4083 ( .A(n2813), .B(sreg[251]), .Z(n2815) );
  NAND U4084 ( .A(n2808), .B(sreg[250]), .Z(n2812) );
  OR U4085 ( .A(n2810), .B(n2809), .Z(n2811) );
  AND U4086 ( .A(n2812), .B(n2811), .Z(n2814) );
  XOR U4087 ( .A(n2815), .B(n2814), .Z(c[251]) );
  NAND U4088 ( .A(n2813), .B(sreg[251]), .Z(n2817) );
  OR U4089 ( .A(n2815), .B(n2814), .Z(n2816) );
  NAND U4090 ( .A(n2817), .B(n2816), .Z(n3066) );
  XNOR U4091 ( .A(n3066), .B(sreg[252]), .Z(n3068) );
  NANDN U4092 ( .A(n2819), .B(n2818), .Z(n2823) );
  NAND U4093 ( .A(n2821), .B(n2820), .Z(n2822) );
  NAND U4094 ( .A(n2823), .B(n2822), .Z(n2941) );
  NANDN U4095 ( .A(n2825), .B(n2824), .Z(n2829) );
  NAND U4096 ( .A(n2827), .B(n2826), .Z(n2828) );
  NAND U4097 ( .A(n2829), .B(n2828), .Z(n2939) );
  OR U4098 ( .A(n2831), .B(n2830), .Z(n2835) );
  NAND U4099 ( .A(n2833), .B(n2832), .Z(n2834) );
  NAND U4100 ( .A(n2835), .B(n2834), .Z(n3063) );
  NANDN U4101 ( .A(n2837), .B(n2836), .Z(n2841) );
  NAND U4102 ( .A(n2839), .B(n2838), .Z(n2840) );
  NAND U4103 ( .A(n2841), .B(n2840), .Z(n3051) );
  NANDN U4104 ( .A(n2843), .B(n2842), .Z(n2847) );
  NAND U4105 ( .A(n2845), .B(n2844), .Z(n2846) );
  NAND U4106 ( .A(n2847), .B(n2846), .Z(n3048) );
  XNOR U4107 ( .A(b[13]), .B(a[16]), .Z(n2999) );
  NANDN U4108 ( .A(n2999), .B(n37424), .Z(n2850) );
  NANDN U4109 ( .A(n2848), .B(n37425), .Z(n2849) );
  NAND U4110 ( .A(n2850), .B(n2849), .Z(n3011) );
  OR U4111 ( .A(n2851), .B(n36105), .Z(n2853) );
  XOR U4112 ( .A(b[3]), .B(n7202), .Z(n3017) );
  NANDN U4113 ( .A(n3017), .B(n36107), .Z(n2852) );
  NAND U4114 ( .A(n2853), .B(n2852), .Z(n3008) );
  NANDN U4115 ( .A(n2854), .B(n38205), .Z(n2856) );
  XOR U4116 ( .A(b[23]), .B(n4305), .Z(n2960) );
  OR U4117 ( .A(n2960), .B(n38268), .Z(n2855) );
  AND U4118 ( .A(n2856), .B(n2855), .Z(n3009) );
  XNOR U4119 ( .A(n3008), .B(n3009), .Z(n3010) );
  XOR U4120 ( .A(n3011), .B(n3010), .Z(n3049) );
  XNOR U4121 ( .A(n3048), .B(n3049), .Z(n3050) );
  XOR U4122 ( .A(n3051), .B(n3050), .Z(n3060) );
  XNOR U4123 ( .A(b[5]), .B(a[24]), .Z(n3014) );
  NANDN U4124 ( .A(n3014), .B(n36587), .Z(n2859) );
  NANDN U4125 ( .A(n2857), .B(n36588), .Z(n2858) );
  NAND U4126 ( .A(n2859), .B(n2858), .Z(n3033) );
  XNOR U4127 ( .A(b[19]), .B(a[10]), .Z(n3002) );
  NANDN U4128 ( .A(n3002), .B(n37934), .Z(n2862) );
  NANDN U4129 ( .A(n2860), .B(n37935), .Z(n2861) );
  NAND U4130 ( .A(n2862), .B(n2861), .Z(n3030) );
  XNOR U4131 ( .A(n1056), .B(a[8]), .Z(n3027) );
  NAND U4132 ( .A(n3027), .B(n38101), .Z(n2865) );
  NANDN U4133 ( .A(n2863), .B(n38102), .Z(n2864) );
  AND U4134 ( .A(n2865), .B(n2864), .Z(n3031) );
  XNOR U4135 ( .A(n3030), .B(n3031), .Z(n3032) );
  XNOR U4136 ( .A(n3033), .B(n3032), .Z(n3045) );
  XOR U4137 ( .A(b[7]), .B(a[22]), .Z(n3024) );
  NAND U4138 ( .A(n3024), .B(n36701), .Z(n2868) );
  NAND U4139 ( .A(n2866), .B(n36702), .Z(n2867) );
  NAND U4140 ( .A(n2868), .B(n2867), .Z(n2977) );
  XOR U4141 ( .A(b[11]), .B(a[18]), .Z(n3005) );
  NANDN U4142 ( .A(n37311), .B(n3005), .Z(n2871) );
  NAND U4143 ( .A(n2869), .B(n37218), .Z(n2870) );
  NAND U4144 ( .A(n2871), .B(n2870), .Z(n2974) );
  NAND U4145 ( .A(n2872), .B(n37762), .Z(n2874) );
  XOR U4146 ( .A(b[17]), .B(a[12]), .Z(n3020) );
  NAND U4147 ( .A(n3020), .B(n37764), .Z(n2873) );
  AND U4148 ( .A(n2874), .B(n2873), .Z(n2975) );
  XNOR U4149 ( .A(n2974), .B(n2975), .Z(n2976) );
  XNOR U4150 ( .A(n2977), .B(n2976), .Z(n3042) );
  XNOR U4151 ( .A(b[9]), .B(a[20]), .Z(n2966) );
  NANDN U4152 ( .A(n2966), .B(n36925), .Z(n2877) );
  NANDN U4153 ( .A(n2875), .B(n36926), .Z(n2876) );
  NAND U4154 ( .A(n2877), .B(n2876), .Z(n3043) );
  XNOR U4155 ( .A(n3042), .B(n3043), .Z(n3044) );
  XOR U4156 ( .A(n3045), .B(n3044), .Z(n3061) );
  XNOR U4157 ( .A(n3060), .B(n3061), .Z(n3062) );
  XNOR U4158 ( .A(n3063), .B(n3062), .Z(n2959) );
  NANDN U4159 ( .A(n2879), .B(n2878), .Z(n2883) );
  NANDN U4160 ( .A(n2881), .B(n2880), .Z(n2882) );
  NAND U4161 ( .A(n2883), .B(n2882), .Z(n3039) );
  NANDN U4162 ( .A(n2885), .B(n2884), .Z(n2889) );
  NAND U4163 ( .A(n2887), .B(n2886), .Z(n2888) );
  NAND U4164 ( .A(n2889), .B(n2888), .Z(n3057) );
  NANDN U4165 ( .A(n1049), .B(a[28]), .Z(n2890) );
  XNOR U4166 ( .A(b[1]), .B(n2890), .Z(n2892) );
  NANDN U4167 ( .A(b[0]), .B(a[27]), .Z(n2891) );
  AND U4168 ( .A(n2892), .B(n2891), .Z(n2970) );
  AND U4169 ( .A(a[0]), .B(n1047), .Z(n3023) );
  XOR U4170 ( .A(b[25]), .B(a[4]), .Z(n2963) );
  NAND U4171 ( .A(n2963), .B(n38325), .Z(n2895) );
  NAND U4172 ( .A(n2893), .B(n38326), .Z(n2894) );
  NAND U4173 ( .A(n2895), .B(n2894), .Z(n2969) );
  XNOR U4174 ( .A(n3023), .B(n2969), .Z(n2971) );
  XNOR U4175 ( .A(n2970), .B(n2971), .Z(n3055) );
  XOR U4176 ( .A(b[27]), .B(a[2]), .Z(n2986) );
  NAND U4177 ( .A(n38423), .B(n2986), .Z(n2898) );
  NAND U4178 ( .A(n2896), .B(n38424), .Z(n2897) );
  NAND U4179 ( .A(n2898), .B(n2897), .Z(n2980) );
  XNOR U4180 ( .A(b[15]), .B(a[14]), .Z(n2996) );
  OR U4181 ( .A(n2996), .B(n37665), .Z(n2901) );
  NANDN U4182 ( .A(n2899), .B(n37604), .Z(n2900) );
  AND U4183 ( .A(n2901), .B(n2900), .Z(n2981) );
  XNOR U4184 ( .A(n2980), .B(n2981), .Z(n2982) );
  NAND U4185 ( .A(n2903), .B(n2902), .Z(n2983) );
  XNOR U4186 ( .A(n2982), .B(n2983), .Z(n3054) );
  XOR U4187 ( .A(n3055), .B(n3054), .Z(n3056) );
  XOR U4188 ( .A(n3057), .B(n3056), .Z(n3036) );
  NANDN U4189 ( .A(n2905), .B(n2904), .Z(n2909) );
  NAND U4190 ( .A(n2907), .B(n2906), .Z(n2908) );
  AND U4191 ( .A(n2909), .B(n2908), .Z(n3037) );
  XNOR U4192 ( .A(n3036), .B(n3037), .Z(n3038) );
  XNOR U4193 ( .A(n3039), .B(n3038), .Z(n2956) );
  NANDN U4194 ( .A(n2911), .B(n2910), .Z(n2915) );
  NAND U4195 ( .A(n2913), .B(n2912), .Z(n2914) );
  AND U4196 ( .A(n2915), .B(n2914), .Z(n2957) );
  XNOR U4197 ( .A(n2956), .B(n2957), .Z(n2958) );
  XOR U4198 ( .A(n2959), .B(n2958), .Z(n2946) );
  NANDN U4199 ( .A(n2917), .B(n2916), .Z(n2921) );
  NAND U4200 ( .A(n2919), .B(n2918), .Z(n2920) );
  NAND U4201 ( .A(n2921), .B(n2920), .Z(n2953) );
  NANDN U4202 ( .A(n2923), .B(n2922), .Z(n2927) );
  OR U4203 ( .A(n2925), .B(n2924), .Z(n2926) );
  NAND U4204 ( .A(n2927), .B(n2926), .Z(n2951) );
  XNOR U4205 ( .A(n2951), .B(n2950), .Z(n2952) );
  XOR U4206 ( .A(n2953), .B(n2952), .Z(n2944) );
  NANDN U4207 ( .A(n2933), .B(n2932), .Z(n2937) );
  NAND U4208 ( .A(n2935), .B(n2934), .Z(n2936) );
  NAND U4209 ( .A(n2937), .B(n2936), .Z(n2945) );
  XNOR U4210 ( .A(n2944), .B(n2945), .Z(n2947) );
  XOR U4211 ( .A(n2946), .B(n2947), .Z(n2938) );
  XOR U4212 ( .A(n2939), .B(n2938), .Z(n2940) );
  XOR U4213 ( .A(n2941), .B(n2940), .Z(n3067) );
  XOR U4214 ( .A(n3068), .B(n3067), .Z(c[252]) );
  NAND U4215 ( .A(n2939), .B(n2938), .Z(n2943) );
  NAND U4216 ( .A(n2941), .B(n2940), .Z(n2942) );
  NAND U4217 ( .A(n2943), .B(n2942), .Z(n3079) );
  NANDN U4218 ( .A(n2945), .B(n2944), .Z(n2949) );
  NAND U4219 ( .A(n2947), .B(n2946), .Z(n2948) );
  NAND U4220 ( .A(n2949), .B(n2948), .Z(n3076) );
  NANDN U4221 ( .A(n2951), .B(n2950), .Z(n2955) );
  NANDN U4222 ( .A(n2953), .B(n2952), .Z(n2954) );
  NAND U4223 ( .A(n2955), .B(n2954), .Z(n3201) );
  NANDN U4224 ( .A(n2960), .B(n38205), .Z(n2962) );
  XNOR U4225 ( .A(b[23]), .B(a[7]), .Z(n3169) );
  OR U4226 ( .A(n3169), .B(n38268), .Z(n2961) );
  NAND U4227 ( .A(n2962), .B(n2961), .Z(n3187) );
  XOR U4228 ( .A(b[25]), .B(a[5]), .Z(n3172) );
  NAND U4229 ( .A(n3172), .B(n38325), .Z(n2965) );
  NAND U4230 ( .A(n2963), .B(n38326), .Z(n2964) );
  NAND U4231 ( .A(n2965), .B(n2964), .Z(n3184) );
  XNOR U4232 ( .A(b[9]), .B(a[21]), .Z(n3117) );
  NANDN U4233 ( .A(n3117), .B(n36925), .Z(n2968) );
  NANDN U4234 ( .A(n2966), .B(n36926), .Z(n2967) );
  AND U4235 ( .A(n2968), .B(n2967), .Z(n3185) );
  XNOR U4236 ( .A(n3184), .B(n3185), .Z(n3186) );
  XNOR U4237 ( .A(n3187), .B(n3186), .Z(n3088) );
  NAND U4238 ( .A(n2969), .B(n3023), .Z(n2973) );
  NANDN U4239 ( .A(n2971), .B(n2970), .Z(n2972) );
  NAND U4240 ( .A(n2973), .B(n2972), .Z(n3089) );
  XNOR U4241 ( .A(n3088), .B(n3089), .Z(n3090) );
  NANDN U4242 ( .A(n2975), .B(n2974), .Z(n2979) );
  NAND U4243 ( .A(n2977), .B(n2976), .Z(n2978) );
  AND U4244 ( .A(n2979), .B(n2978), .Z(n3091) );
  XNOR U4245 ( .A(n3090), .B(n3091), .Z(n3083) );
  NANDN U4246 ( .A(n2981), .B(n2980), .Z(n2985) );
  NANDN U4247 ( .A(n2983), .B(n2982), .Z(n2984) );
  NAND U4248 ( .A(n2985), .B(n2984), .Z(n3097) );
  XOR U4249 ( .A(b[27]), .B(a[3]), .Z(n3166) );
  NAND U4250 ( .A(n38423), .B(n3166), .Z(n2988) );
  NAND U4251 ( .A(n2986), .B(n38424), .Z(n2987) );
  NAND U4252 ( .A(n2988), .B(n2987), .Z(n3101) );
  XNOR U4253 ( .A(b[29]), .B(a[1]), .Z(n3105) );
  NOR U4254 ( .A(n1048), .B(n3105), .Z(n2992) );
  XNOR U4255 ( .A(n3393), .B(b[29]), .Z(n2990) );
  XNOR U4256 ( .A(n1058), .B(b[28]), .Z(n2989) );
  ANDN U4257 ( .B(n2989), .A(n1047), .Z(n38490) );
  NAND U4258 ( .A(n2990), .B(n38490), .Z(n2991) );
  NANDN U4259 ( .A(n2992), .B(n2991), .Z(n3100) );
  XNOR U4260 ( .A(n3101), .B(n3100), .Z(n3135) );
  NANDN U4261 ( .A(n1049), .B(a[29]), .Z(n2993) );
  XNOR U4262 ( .A(b[1]), .B(n2993), .Z(n2995) );
  NANDN U4263 ( .A(b[0]), .B(a[28]), .Z(n2994) );
  AND U4264 ( .A(n2995), .B(n2994), .Z(n3133) );
  XNOR U4265 ( .A(n1054), .B(a[15]), .Z(n3108) );
  NANDN U4266 ( .A(n37665), .B(n3108), .Z(n2998) );
  NANDN U4267 ( .A(n2996), .B(n37604), .Z(n2997) );
  AND U4268 ( .A(n2998), .B(n2997), .Z(n3132) );
  XNOR U4269 ( .A(n3133), .B(n3132), .Z(n3134) );
  XOR U4270 ( .A(n3135), .B(n3134), .Z(n3094) );
  XNOR U4271 ( .A(b[13]), .B(a[17]), .Z(n3123) );
  NANDN U4272 ( .A(n3123), .B(n37424), .Z(n3001) );
  NANDN U4273 ( .A(n2999), .B(n37425), .Z(n3000) );
  NAND U4274 ( .A(n3001), .B(n3000), .Z(n3141) );
  XNOR U4275 ( .A(b[19]), .B(a[11]), .Z(n3126) );
  NANDN U4276 ( .A(n3126), .B(n37934), .Z(n3004) );
  NANDN U4277 ( .A(n3002), .B(n37935), .Z(n3003) );
  NAND U4278 ( .A(n3004), .B(n3003), .Z(n3138) );
  XOR U4279 ( .A(b[11]), .B(a[19]), .Z(n3120) );
  NANDN U4280 ( .A(n37311), .B(n3120), .Z(n3007) );
  NAND U4281 ( .A(n3005), .B(n37218), .Z(n3006) );
  AND U4282 ( .A(n3007), .B(n3006), .Z(n3139) );
  XNOR U4283 ( .A(n3138), .B(n3139), .Z(n3140) );
  XNOR U4284 ( .A(n3141), .B(n3140), .Z(n3095) );
  XOR U4285 ( .A(n3094), .B(n3095), .Z(n3096) );
  XNOR U4286 ( .A(n3097), .B(n3096), .Z(n3159) );
  NANDN U4287 ( .A(n3009), .B(n3008), .Z(n3013) );
  NAND U4288 ( .A(n3011), .B(n3010), .Z(n3012) );
  NAND U4289 ( .A(n3013), .B(n3012), .Z(n3156) );
  XOR U4290 ( .A(b[5]), .B(n7069), .Z(n3111) );
  NANDN U4291 ( .A(n3111), .B(n36587), .Z(n3016) );
  NANDN U4292 ( .A(n3014), .B(n36588), .Z(n3015) );
  NAND U4293 ( .A(n3016), .B(n3015), .Z(n3181) );
  OR U4294 ( .A(n3017), .B(n36105), .Z(n3019) );
  XNOR U4295 ( .A(b[3]), .B(a[27]), .Z(n3114) );
  NANDN U4296 ( .A(n3114), .B(n36107), .Z(n3018) );
  NAND U4297 ( .A(n3019), .B(n3018), .Z(n3178) );
  NAND U4298 ( .A(n3020), .B(n37762), .Z(n3022) );
  XOR U4299 ( .A(b[17]), .B(a[13]), .Z(n3102) );
  NAND U4300 ( .A(n3102), .B(n37764), .Z(n3021) );
  AND U4301 ( .A(n3022), .B(n3021), .Z(n3179) );
  XNOR U4302 ( .A(n3178), .B(n3179), .Z(n3180) );
  XNOR U4303 ( .A(n3181), .B(n3180), .Z(n3150) );
  NAND U4304 ( .A(b[28]), .B(b[27]), .Z(n38527) );
  AND U4305 ( .A(n38527), .B(b[29]), .Z(n38567) );
  NANDN U4306 ( .A(n3023), .B(n38567), .Z(n3190) );
  XOR U4307 ( .A(b[7]), .B(a[23]), .Z(n3129) );
  NAND U4308 ( .A(n36701), .B(n3129), .Z(n3026) );
  NAND U4309 ( .A(n36702), .B(n3024), .Z(n3025) );
  NAND U4310 ( .A(n3026), .B(n3025), .Z(n3191) );
  XNOR U4311 ( .A(n3190), .B(n3191), .Z(n3192) );
  XNOR U4312 ( .A(b[21]), .B(a[9]), .Z(n3175) );
  NANDN U4313 ( .A(n3175), .B(n38101), .Z(n3029) );
  NAND U4314 ( .A(n38102), .B(n3027), .Z(n3028) );
  AND U4315 ( .A(n3029), .B(n3028), .Z(n3193) );
  XNOR U4316 ( .A(n3192), .B(n3193), .Z(n3151) );
  XOR U4317 ( .A(n3150), .B(n3151), .Z(n3153) );
  NANDN U4318 ( .A(n3031), .B(n3030), .Z(n3035) );
  NAND U4319 ( .A(n3033), .B(n3032), .Z(n3034) );
  NAND U4320 ( .A(n3035), .B(n3034), .Z(n3152) );
  XOR U4321 ( .A(n3156), .B(n3157), .Z(n3158) );
  XOR U4322 ( .A(n3159), .B(n3158), .Z(n3082) );
  XOR U4323 ( .A(n3083), .B(n3082), .Z(n3085) );
  NANDN U4324 ( .A(n3037), .B(n3036), .Z(n3041) );
  NAND U4325 ( .A(n3039), .B(n3038), .Z(n3040) );
  NAND U4326 ( .A(n3041), .B(n3040), .Z(n3084) );
  XNOR U4327 ( .A(n3085), .B(n3084), .Z(n3197) );
  NANDN U4328 ( .A(n3043), .B(n3042), .Z(n3047) );
  NAND U4329 ( .A(n3045), .B(n3044), .Z(n3046) );
  NAND U4330 ( .A(n3047), .B(n3046), .Z(n3147) );
  NANDN U4331 ( .A(n3049), .B(n3048), .Z(n3053) );
  NANDN U4332 ( .A(n3051), .B(n3050), .Z(n3052) );
  NAND U4333 ( .A(n3053), .B(n3052), .Z(n3144) );
  OR U4334 ( .A(n3055), .B(n3054), .Z(n3059) );
  NANDN U4335 ( .A(n3057), .B(n3056), .Z(n3058) );
  AND U4336 ( .A(n3059), .B(n3058), .Z(n3145) );
  XNOR U4337 ( .A(n3144), .B(n3145), .Z(n3146) );
  XNOR U4338 ( .A(n3147), .B(n3146), .Z(n3194) );
  NANDN U4339 ( .A(n3061), .B(n3060), .Z(n3065) );
  NAND U4340 ( .A(n3063), .B(n3062), .Z(n3064) );
  AND U4341 ( .A(n3065), .B(n3064), .Z(n3195) );
  XNOR U4342 ( .A(n3194), .B(n3195), .Z(n3196) );
  XNOR U4343 ( .A(n3197), .B(n3196), .Z(n3199) );
  XOR U4344 ( .A(n3198), .B(n3199), .Z(n3200) );
  XOR U4345 ( .A(n3201), .B(n3200), .Z(n3077) );
  XNOR U4346 ( .A(n3076), .B(n3077), .Z(n3078) );
  XNOR U4347 ( .A(n3079), .B(n3078), .Z(n3071) );
  XNOR U4348 ( .A(n3071), .B(sreg[253]), .Z(n3073) );
  NAND U4349 ( .A(n3066), .B(sreg[252]), .Z(n3070) );
  OR U4350 ( .A(n3068), .B(n3067), .Z(n3069) );
  AND U4351 ( .A(n3070), .B(n3069), .Z(n3072) );
  XOR U4352 ( .A(n3073), .B(n3072), .Z(c[253]) );
  NAND U4353 ( .A(n3071), .B(sreg[253]), .Z(n3075) );
  OR U4354 ( .A(n3073), .B(n3072), .Z(n3074) );
  NAND U4355 ( .A(n3075), .B(n3074), .Z(n3337) );
  XNOR U4356 ( .A(n3337), .B(sreg[254]), .Z(n3339) );
  NANDN U4357 ( .A(n3077), .B(n3076), .Z(n3081) );
  NAND U4358 ( .A(n3079), .B(n3078), .Z(n3080) );
  NAND U4359 ( .A(n3081), .B(n3080), .Z(n3207) );
  NANDN U4360 ( .A(n3083), .B(n3082), .Z(n3087) );
  OR U4361 ( .A(n3085), .B(n3084), .Z(n3086) );
  NAND U4362 ( .A(n3087), .B(n3086), .Z(n3210) );
  NANDN U4363 ( .A(n3089), .B(n3088), .Z(n3093) );
  NAND U4364 ( .A(n3091), .B(n3090), .Z(n3092) );
  NAND U4365 ( .A(n3093), .B(n3092), .Z(n3262) );
  OR U4366 ( .A(n3095), .B(n3094), .Z(n3099) );
  NAND U4367 ( .A(n3097), .B(n3096), .Z(n3098) );
  NAND U4368 ( .A(n3099), .B(n3098), .Z(n3259) );
  NAND U4369 ( .A(n3101), .B(n3100), .Z(n3290) );
  XNOR U4370 ( .A(b[17]), .B(a[14]), .Z(n3285) );
  NANDN U4371 ( .A(n3285), .B(n37764), .Z(n3104) );
  NAND U4372 ( .A(n3102), .B(n37762), .Z(n3103) );
  NAND U4373 ( .A(n3104), .B(n3103), .Z(n3289) );
  NANDN U4374 ( .A(n3105), .B(n38490), .Z(n3107) );
  XNOR U4375 ( .A(n1058), .B(a[2]), .Z(n3240) );
  NANDN U4376 ( .A(n1048), .B(n3240), .Z(n3106) );
  AND U4377 ( .A(n3107), .B(n3106), .Z(n3288) );
  XNOR U4378 ( .A(n3289), .B(n3288), .Z(n3291) );
  XNOR U4379 ( .A(n3290), .B(n3291), .Z(n3265) );
  XNOR U4380 ( .A(b[15]), .B(a[16]), .Z(n3250) );
  OR U4381 ( .A(n3250), .B(n37665), .Z(n3110) );
  NAND U4382 ( .A(n3108), .B(n37604), .Z(n3109) );
  NAND U4383 ( .A(n3110), .B(n3109), .Z(n3307) );
  XOR U4384 ( .A(b[5]), .B(n7202), .Z(n3276) );
  NANDN U4385 ( .A(n3276), .B(n36587), .Z(n3113) );
  NANDN U4386 ( .A(n3111), .B(n36588), .Z(n3112) );
  NAND U4387 ( .A(n3113), .B(n3112), .Z(n3304) );
  OR U4388 ( .A(n3114), .B(n36105), .Z(n3116) );
  XNOR U4389 ( .A(b[3]), .B(a[28]), .Z(n3282) );
  NANDN U4390 ( .A(n3282), .B(n36107), .Z(n3115) );
  AND U4391 ( .A(n3116), .B(n3115), .Z(n3305) );
  XNOR U4392 ( .A(n3304), .B(n3305), .Z(n3306) );
  XNOR U4393 ( .A(n3307), .B(n3306), .Z(n3266) );
  XNOR U4394 ( .A(n3265), .B(n3266), .Z(n3267) );
  XNOR U4395 ( .A(b[9]), .B(a[22]), .Z(n3310) );
  NANDN U4396 ( .A(n3310), .B(n36925), .Z(n3119) );
  NANDN U4397 ( .A(n3117), .B(n36926), .Z(n3118) );
  NAND U4398 ( .A(n3119), .B(n3118), .Z(n3292) );
  XOR U4399 ( .A(b[11]), .B(a[20]), .Z(n3328) );
  NANDN U4400 ( .A(n37311), .B(n3328), .Z(n3122) );
  NAND U4401 ( .A(n3120), .B(n37218), .Z(n3121) );
  AND U4402 ( .A(n3122), .B(n3121), .Z(n3293) );
  XNOR U4403 ( .A(n3292), .B(n3293), .Z(n3294) );
  XNOR U4404 ( .A(b[13]), .B(a[18]), .Z(n3313) );
  NANDN U4405 ( .A(n3313), .B(n37424), .Z(n3125) );
  NANDN U4406 ( .A(n3123), .B(n37425), .Z(n3124) );
  NAND U4407 ( .A(n3125), .B(n3124), .Z(n3237) );
  XNOR U4408 ( .A(b[19]), .B(a[12]), .Z(n3279) );
  NANDN U4409 ( .A(n3279), .B(n37934), .Z(n3128) );
  NANDN U4410 ( .A(n3126), .B(n37935), .Z(n3127) );
  NAND U4411 ( .A(n3128), .B(n3127), .Z(n3234) );
  XOR U4412 ( .A(b[7]), .B(a[24]), .Z(n3273) );
  NAND U4413 ( .A(n3273), .B(n36701), .Z(n3131) );
  NAND U4414 ( .A(n3129), .B(n36702), .Z(n3130) );
  AND U4415 ( .A(n3131), .B(n3130), .Z(n3235) );
  XNOR U4416 ( .A(n3234), .B(n3235), .Z(n3236) );
  XOR U4417 ( .A(n3237), .B(n3236), .Z(n3295) );
  XOR U4418 ( .A(n3294), .B(n3295), .Z(n3268) );
  XOR U4419 ( .A(n3267), .B(n3268), .Z(n3231) );
  NANDN U4420 ( .A(n3133), .B(n3132), .Z(n3137) );
  NAND U4421 ( .A(n3135), .B(n3134), .Z(n3136) );
  NAND U4422 ( .A(n3137), .B(n3136), .Z(n3228) );
  NANDN U4423 ( .A(n3139), .B(n3138), .Z(n3143) );
  NAND U4424 ( .A(n3141), .B(n3140), .Z(n3142) );
  NAND U4425 ( .A(n3143), .B(n3142), .Z(n3229) );
  XNOR U4426 ( .A(n3228), .B(n3229), .Z(n3230) );
  XOR U4427 ( .A(n3231), .B(n3230), .Z(n3260) );
  XOR U4428 ( .A(n3259), .B(n3260), .Z(n3261) );
  XNOR U4429 ( .A(n3262), .B(n3261), .Z(n3216) );
  NANDN U4430 ( .A(n3145), .B(n3144), .Z(n3149) );
  NAND U4431 ( .A(n3147), .B(n3146), .Z(n3148) );
  NAND U4432 ( .A(n3149), .B(n3148), .Z(n3217) );
  XNOR U4433 ( .A(n3216), .B(n3217), .Z(n3218) );
  NANDN U4434 ( .A(n3151), .B(n3150), .Z(n3155) );
  OR U4435 ( .A(n3153), .B(n3152), .Z(n3154) );
  NAND U4436 ( .A(n3155), .B(n3154), .Z(n3332) );
  OR U4437 ( .A(n3157), .B(n3156), .Z(n3161) );
  NAND U4438 ( .A(n3159), .B(n3158), .Z(n3160) );
  AND U4439 ( .A(n3161), .B(n3160), .Z(n3331) );
  XNOR U4440 ( .A(n3332), .B(n3331), .Z(n3333) );
  ANDN U4441 ( .B(a[30]), .A(n1049), .Z(n3162) );
  XOR U4442 ( .A(b[1]), .B(n3162), .Z(n3165) );
  NANDN U4443 ( .A(b[0]), .B(b[1]), .Z(n3163) );
  NANDN U4444 ( .A(n3163), .B(a[29]), .Z(n3164) );
  NAND U4445 ( .A(n3165), .B(n3164), .Z(n3256) );
  XOR U4446 ( .A(b[27]), .B(a[4]), .Z(n3325) );
  NAND U4447 ( .A(n38423), .B(n3325), .Z(n3168) );
  NAND U4448 ( .A(n3166), .B(n38424), .Z(n3167) );
  NAND U4449 ( .A(n3168), .B(n3167), .Z(n3253) );
  XNOR U4450 ( .A(n1058), .B(b[30]), .Z(n38552) );
  NANDN U4451 ( .A(n3393), .B(n38552), .Z(n3254) );
  XNOR U4452 ( .A(n3253), .B(n3254), .Z(n3255) );
  XOR U4453 ( .A(n3256), .B(n3255), .Z(n3272) );
  NANDN U4454 ( .A(n3169), .B(n38205), .Z(n3171) );
  XNOR U4455 ( .A(b[23]), .B(a[8]), .Z(n3319) );
  OR U4456 ( .A(n3319), .B(n38268), .Z(n3170) );
  NAND U4457 ( .A(n3171), .B(n3170), .Z(n3301) );
  XNOR U4458 ( .A(b[25]), .B(a[6]), .Z(n3322) );
  NANDN U4459 ( .A(n3322), .B(n38325), .Z(n3174) );
  NAND U4460 ( .A(n3172), .B(n38326), .Z(n3173) );
  NAND U4461 ( .A(n3174), .B(n3173), .Z(n3298) );
  XNOR U4462 ( .A(b[21]), .B(a[10]), .Z(n3316) );
  NANDN U4463 ( .A(n3316), .B(n38101), .Z(n3177) );
  NANDN U4464 ( .A(n3175), .B(n38102), .Z(n3176) );
  AND U4465 ( .A(n3177), .B(n3176), .Z(n3299) );
  XNOR U4466 ( .A(n3298), .B(n3299), .Z(n3300) );
  XNOR U4467 ( .A(n3301), .B(n3300), .Z(n3269) );
  NANDN U4468 ( .A(n3179), .B(n3178), .Z(n3183) );
  NAND U4469 ( .A(n3181), .B(n3180), .Z(n3182) );
  NAND U4470 ( .A(n3183), .B(n3182), .Z(n3270) );
  XNOR U4471 ( .A(n3269), .B(n3270), .Z(n3271) );
  XNOR U4472 ( .A(n3272), .B(n3271), .Z(n3225) );
  NANDN U4473 ( .A(n3185), .B(n3184), .Z(n3189) );
  NAND U4474 ( .A(n3187), .B(n3186), .Z(n3188) );
  NAND U4475 ( .A(n3189), .B(n3188), .Z(n3222) );
  XNOR U4476 ( .A(n3222), .B(n3223), .Z(n3224) );
  XOR U4477 ( .A(n3225), .B(n3224), .Z(n3334) );
  XOR U4478 ( .A(n3333), .B(n3334), .Z(n3219) );
  XOR U4479 ( .A(n3218), .B(n3219), .Z(n3211) );
  XNOR U4480 ( .A(n3210), .B(n3211), .Z(n3212) );
  XNOR U4481 ( .A(n3212), .B(n3213), .Z(n3205) );
  OR U4482 ( .A(n3199), .B(n3198), .Z(n3203) );
  NAND U4483 ( .A(n3201), .B(n3200), .Z(n3202) );
  AND U4484 ( .A(n3203), .B(n3202), .Z(n3204) );
  XNOR U4485 ( .A(n3205), .B(n3204), .Z(n3206) );
  XOR U4486 ( .A(n3207), .B(n3206), .Z(n3338) );
  XOR U4487 ( .A(n3339), .B(n3338), .Z(c[254]) );
  NANDN U4488 ( .A(n3205), .B(n3204), .Z(n3209) );
  NAND U4489 ( .A(n3207), .B(n3206), .Z(n3208) );
  NAND U4490 ( .A(n3209), .B(n3208), .Z(n3350) );
  NANDN U4491 ( .A(n3211), .B(n3210), .Z(n3215) );
  NAND U4492 ( .A(n3213), .B(n3212), .Z(n3214) );
  NAND U4493 ( .A(n3215), .B(n3214), .Z(n3348) );
  NANDN U4494 ( .A(n3217), .B(n3216), .Z(n3221) );
  NAND U4495 ( .A(n3219), .B(n3218), .Z(n3220) );
  NAND U4496 ( .A(n3221), .B(n3220), .Z(n3483) );
  NANDN U4497 ( .A(n3223), .B(n3222), .Z(n3227) );
  NAND U4498 ( .A(n3225), .B(n3224), .Z(n3226) );
  NAND U4499 ( .A(n3227), .B(n3226), .Z(n3360) );
  NANDN U4500 ( .A(n3229), .B(n3228), .Z(n3233) );
  NANDN U4501 ( .A(n3231), .B(n3230), .Z(n3232) );
  NAND U4502 ( .A(n3233), .B(n3232), .Z(n3358) );
  NANDN U4503 ( .A(n3235), .B(n3234), .Z(n3239) );
  NAND U4504 ( .A(n3237), .B(n3236), .Z(n3238) );
  NAND U4505 ( .A(n3239), .B(n3238), .Z(n3418) );
  NAND U4506 ( .A(n3240), .B(n38490), .Z(n3242) );
  XNOR U4507 ( .A(n1058), .B(a[3]), .Z(n3387) );
  NANDN U4508 ( .A(n1048), .B(n3387), .Z(n3241) );
  NAND U4509 ( .A(n3242), .B(n3241), .Z(n3449) );
  XNOR U4510 ( .A(b[31]), .B(a[1]), .Z(n3436) );
  ANDN U4511 ( .B(n38552), .A(n3436), .Z(n3246) );
  XNOR U4512 ( .A(n1059), .B(a[0]), .Z(n3244) );
  XOR U4513 ( .A(b[31]), .B(b[29]), .Z(n3243) );
  XOR U4514 ( .A(n1058), .B(b[30]), .Z(n38574) );
  AND U4515 ( .A(n3243), .B(n38574), .Z(n38553) );
  NAND U4516 ( .A(n3244), .B(n38553), .Z(n3245) );
  NANDN U4517 ( .A(n3246), .B(n3245), .Z(n3448) );
  XNOR U4518 ( .A(n3449), .B(n3448), .Z(n3384) );
  NANDN U4519 ( .A(n1049), .B(a[31]), .Z(n3247) );
  XNOR U4520 ( .A(b[1]), .B(n3247), .Z(n3249) );
  IV U4521 ( .A(a[30]), .Z(n7434) );
  NANDN U4522 ( .A(n7434), .B(n1049), .Z(n3248) );
  AND U4523 ( .A(n3249), .B(n3248), .Z(n3382) );
  XNOR U4524 ( .A(n1054), .B(a[17]), .Z(n3400) );
  NANDN U4525 ( .A(n37665), .B(n3400), .Z(n3252) );
  NANDN U4526 ( .A(n3250), .B(n37604), .Z(n3251) );
  AND U4527 ( .A(n3252), .B(n3251), .Z(n3381) );
  XNOR U4528 ( .A(n3382), .B(n3381), .Z(n3383) );
  XOR U4529 ( .A(n3384), .B(n3383), .Z(n3416) );
  NANDN U4530 ( .A(n3254), .B(n3253), .Z(n3258) );
  NANDN U4531 ( .A(n3256), .B(n3255), .Z(n3257) );
  AND U4532 ( .A(n3258), .B(n3257), .Z(n3415) );
  XOR U4533 ( .A(n3416), .B(n3415), .Z(n3417) );
  XOR U4534 ( .A(n3418), .B(n3417), .Z(n3357) );
  XNOR U4535 ( .A(n3358), .B(n3357), .Z(n3359) );
  XNOR U4536 ( .A(n3360), .B(n3359), .Z(n3354) );
  OR U4537 ( .A(n3260), .B(n3259), .Z(n3264) );
  NAND U4538 ( .A(n3262), .B(n3261), .Z(n3263) );
  NAND U4539 ( .A(n3264), .B(n3263), .Z(n3351) );
  XNOR U4540 ( .A(n3363), .B(n3364), .Z(n3365) );
  XNOR U4541 ( .A(b[7]), .B(a[25]), .Z(n3465) );
  NANDN U4542 ( .A(n3465), .B(n36701), .Z(n3275) );
  NAND U4543 ( .A(n3273), .B(n36702), .Z(n3274) );
  NAND U4544 ( .A(n3275), .B(n3274), .Z(n3445) );
  XNOR U4545 ( .A(b[5]), .B(a[27]), .Z(n3468) );
  NANDN U4546 ( .A(n3468), .B(n36587), .Z(n3278) );
  NANDN U4547 ( .A(n3276), .B(n36588), .Z(n3277) );
  NAND U4548 ( .A(n3278), .B(n3277), .Z(n3442) );
  XNOR U4549 ( .A(b[19]), .B(a[13]), .Z(n3471) );
  NANDN U4550 ( .A(n3471), .B(n37934), .Z(n3281) );
  NANDN U4551 ( .A(n3279), .B(n37935), .Z(n3280) );
  AND U4552 ( .A(n3281), .B(n3280), .Z(n3443) );
  XNOR U4553 ( .A(n3442), .B(n3443), .Z(n3444) );
  XNOR U4554 ( .A(n3445), .B(n3444), .Z(n3410) );
  OR U4555 ( .A(n3282), .B(n36105), .Z(n3284) );
  XNOR U4556 ( .A(b[3]), .B(a[29]), .Z(n3453) );
  NANDN U4557 ( .A(n3453), .B(n36107), .Z(n3283) );
  NAND U4558 ( .A(n3284), .B(n3283), .Z(n3378) );
  NANDN U4559 ( .A(n3285), .B(n37762), .Z(n3287) );
  XOR U4560 ( .A(b[17]), .B(a[15]), .Z(n3450) );
  NAND U4561 ( .A(n3450), .B(n37764), .Z(n3286) );
  NAND U4562 ( .A(n3287), .B(n3286), .Z(n3375) );
  XNOR U4563 ( .A(n3375), .B(n3376), .Z(n3377) );
  XOR U4564 ( .A(n3378), .B(n3377), .Z(n3409) );
  XNOR U4565 ( .A(n3410), .B(n3409), .Z(n3411) );
  XNOR U4566 ( .A(n3411), .B(n3412), .Z(n3370) );
  NANDN U4567 ( .A(n3293), .B(n3292), .Z(n3297) );
  NAND U4568 ( .A(n3295), .B(n3294), .Z(n3296) );
  NAND U4569 ( .A(n3297), .B(n3296), .Z(n3424) );
  NANDN U4570 ( .A(n3299), .B(n3298), .Z(n3303) );
  NAND U4571 ( .A(n3301), .B(n3300), .Z(n3302) );
  NAND U4572 ( .A(n3303), .B(n3302), .Z(n3421) );
  NANDN U4573 ( .A(n3305), .B(n3304), .Z(n3309) );
  NAND U4574 ( .A(n3307), .B(n3306), .Z(n3308) );
  AND U4575 ( .A(n3309), .B(n3308), .Z(n3422) );
  XNOR U4576 ( .A(n3421), .B(n3422), .Z(n3423) );
  XNOR U4577 ( .A(n3424), .B(n3423), .Z(n3369) );
  XNOR U4578 ( .A(n3370), .B(n3369), .Z(n3372) );
  XNOR U4579 ( .A(b[9]), .B(a[23]), .Z(n3433) );
  NANDN U4580 ( .A(n3433), .B(n36925), .Z(n3312) );
  NANDN U4581 ( .A(n3310), .B(n36926), .Z(n3311) );
  NAND U4582 ( .A(n3312), .B(n3311), .Z(n3406) );
  XNOR U4583 ( .A(b[13]), .B(a[19]), .Z(n3394) );
  NANDN U4584 ( .A(n3394), .B(n37424), .Z(n3315) );
  NANDN U4585 ( .A(n3313), .B(n37425), .Z(n3314) );
  NAND U4586 ( .A(n3315), .B(n3314), .Z(n3403) );
  XNOR U4587 ( .A(b[21]), .B(a[11]), .Z(n3397) );
  NANDN U4588 ( .A(n3397), .B(n38101), .Z(n3318) );
  NANDN U4589 ( .A(n3316), .B(n38102), .Z(n3317) );
  AND U4590 ( .A(n3318), .B(n3317), .Z(n3404) );
  XNOR U4591 ( .A(n3403), .B(n3404), .Z(n3405) );
  XNOR U4592 ( .A(n3406), .B(n3405), .Z(n3430) );
  NANDN U4593 ( .A(n3319), .B(n38205), .Z(n3321) );
  XNOR U4594 ( .A(b[23]), .B(a[9]), .Z(n3439) );
  OR U4595 ( .A(n3439), .B(n38268), .Z(n3320) );
  NAND U4596 ( .A(n3321), .B(n3320), .Z(n3477) );
  XOR U4597 ( .A(b[25]), .B(a[7]), .Z(n3459) );
  NAND U4598 ( .A(n3459), .B(n38325), .Z(n3324) );
  NANDN U4599 ( .A(n3322), .B(n38326), .Z(n3323) );
  NAND U4600 ( .A(n3324), .B(n3323), .Z(n3474) );
  XOR U4601 ( .A(b[27]), .B(a[5]), .Z(n3462) );
  NAND U4602 ( .A(n38423), .B(n3462), .Z(n3327) );
  NAND U4603 ( .A(n3325), .B(n38424), .Z(n3326) );
  AND U4604 ( .A(n3327), .B(n3326), .Z(n3475) );
  XNOR U4605 ( .A(n3474), .B(n3475), .Z(n3476) );
  XNOR U4606 ( .A(n3477), .B(n3476), .Z(n3427) );
  XOR U4607 ( .A(b[11]), .B(a[21]), .Z(n3456) );
  NANDN U4608 ( .A(n37311), .B(n3456), .Z(n3330) );
  NAND U4609 ( .A(n37218), .B(n3328), .Z(n3329) );
  NAND U4610 ( .A(n3330), .B(n3329), .Z(n3428) );
  XNOR U4611 ( .A(n3427), .B(n3428), .Z(n3429) );
  XOR U4612 ( .A(n3430), .B(n3429), .Z(n3371) );
  XNOR U4613 ( .A(n3372), .B(n3371), .Z(n3366) );
  XOR U4614 ( .A(n3365), .B(n3366), .Z(n3352) );
  XOR U4615 ( .A(n3351), .B(n3352), .Z(n3353) );
  XOR U4616 ( .A(n3354), .B(n3353), .Z(n3480) );
  NANDN U4617 ( .A(n3332), .B(n3331), .Z(n3336) );
  NAND U4618 ( .A(n3334), .B(n3333), .Z(n3335) );
  NAND U4619 ( .A(n3336), .B(n3335), .Z(n3481) );
  XNOR U4620 ( .A(n3480), .B(n3481), .Z(n3482) );
  XNOR U4621 ( .A(n3483), .B(n3482), .Z(n3347) );
  XOR U4622 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4623 ( .A(n3350), .B(n3349), .Z(n3342) );
  XNOR U4624 ( .A(n3342), .B(sreg[255]), .Z(n3344) );
  NAND U4625 ( .A(n3337), .B(sreg[254]), .Z(n3341) );
  OR U4626 ( .A(n3339), .B(n3338), .Z(n3340) );
  AND U4627 ( .A(n3341), .B(n3340), .Z(n3343) );
  XOR U4628 ( .A(n3344), .B(n3343), .Z(c[255]) );
  NAND U4629 ( .A(n3342), .B(sreg[255]), .Z(n3346) );
  OR U4630 ( .A(n3344), .B(n3343), .Z(n3345) );
  NAND U4631 ( .A(n3346), .B(n3345), .Z(n3624) );
  XNOR U4632 ( .A(n3624), .B(sreg[256]), .Z(n3626) );
  OR U4633 ( .A(n3352), .B(n3351), .Z(n3356) );
  NANDN U4634 ( .A(n3354), .B(n3353), .Z(n3355) );
  NAND U4635 ( .A(n3356), .B(n3355), .Z(n3621) );
  NANDN U4636 ( .A(n3358), .B(n3357), .Z(n3362) );
  NAND U4637 ( .A(n3360), .B(n3359), .Z(n3361) );
  NAND U4638 ( .A(n3362), .B(n3361), .Z(n3619) );
  NANDN U4639 ( .A(n3364), .B(n3363), .Z(n3368) );
  NANDN U4640 ( .A(n3366), .B(n3365), .Z(n3367) );
  NAND U4641 ( .A(n3368), .B(n3367), .Z(n3586) );
  OR U4642 ( .A(n3370), .B(n3369), .Z(n3374) );
  OR U4643 ( .A(n3372), .B(n3371), .Z(n3373) );
  AND U4644 ( .A(n3374), .B(n3373), .Z(n3587) );
  XNOR U4645 ( .A(n3586), .B(n3587), .Z(n3588) );
  NANDN U4646 ( .A(n3376), .B(n3375), .Z(n3380) );
  NAND U4647 ( .A(n3378), .B(n3377), .Z(n3379) );
  NAND U4648 ( .A(n3380), .B(n3379), .Z(n3596) );
  NANDN U4649 ( .A(n3382), .B(n3381), .Z(n3386) );
  NAND U4650 ( .A(n3384), .B(n3383), .Z(n3385) );
  NAND U4651 ( .A(n3386), .B(n3385), .Z(n3597) );
  XNOR U4652 ( .A(n3596), .B(n3597), .Z(n3598) );
  NAND U4653 ( .A(n38490), .B(n3387), .Z(n3389) );
  XNOR U4654 ( .A(n1058), .B(a[4]), .Z(n3510) );
  NANDN U4655 ( .A(n1048), .B(n3510), .Z(n3388) );
  AND U4656 ( .A(n3389), .B(n3388), .Z(n3526) );
  NANDN U4657 ( .A(n1049), .B(a[32]), .Z(n3390) );
  XNOR U4658 ( .A(b[1]), .B(n3390), .Z(n3392) );
  IV U4659 ( .A(a[31]), .Z(n7955) );
  NANDN U4660 ( .A(n7955), .B(n1049), .Z(n3391) );
  AND U4661 ( .A(n3392), .B(n3391), .Z(n3525) );
  XOR U4662 ( .A(n3526), .B(n3525), .Z(n3528) );
  NANDN U4663 ( .A(n3393), .B(b[31]), .Z(n3527) );
  XOR U4664 ( .A(n3528), .B(n3527), .Z(n3492) );
  XNOR U4665 ( .A(n1053), .B(a[20]), .Z(n3571) );
  NAND U4666 ( .A(n3571), .B(n37424), .Z(n3396) );
  NANDN U4667 ( .A(n3394), .B(n37425), .Z(n3395) );
  NAND U4668 ( .A(n3396), .B(n3395), .Z(n3538) );
  XNOR U4669 ( .A(b[21]), .B(a[12]), .Z(n3498) );
  NANDN U4670 ( .A(n3498), .B(n38101), .Z(n3399) );
  NANDN U4671 ( .A(n3397), .B(n38102), .Z(n3398) );
  NAND U4672 ( .A(n3399), .B(n3398), .Z(n3535) );
  XNOR U4673 ( .A(b[15]), .B(a[18]), .Z(n3507) );
  OR U4674 ( .A(n3507), .B(n37665), .Z(n3402) );
  NAND U4675 ( .A(n3400), .B(n37604), .Z(n3401) );
  AND U4676 ( .A(n3402), .B(n3401), .Z(n3536) );
  XNOR U4677 ( .A(n3535), .B(n3536), .Z(n3537) );
  XNOR U4678 ( .A(n3538), .B(n3537), .Z(n3493) );
  XOR U4679 ( .A(n3492), .B(n3493), .Z(n3495) );
  NANDN U4680 ( .A(n3404), .B(n3403), .Z(n3408) );
  NAND U4681 ( .A(n3406), .B(n3405), .Z(n3407) );
  AND U4682 ( .A(n3408), .B(n3407), .Z(n3494) );
  XOR U4683 ( .A(n3495), .B(n3494), .Z(n3599) );
  XNOR U4684 ( .A(n3598), .B(n3599), .Z(n3592) );
  NANDN U4685 ( .A(n3410), .B(n3409), .Z(n3414) );
  NAND U4686 ( .A(n3412), .B(n3411), .Z(n3413) );
  NAND U4687 ( .A(n3414), .B(n3413), .Z(n3593) );
  XNOR U4688 ( .A(n3592), .B(n3593), .Z(n3594) );
  OR U4689 ( .A(n3416), .B(n3415), .Z(n3420) );
  NAND U4690 ( .A(n3418), .B(n3417), .Z(n3419) );
  NAND U4691 ( .A(n3420), .B(n3419), .Z(n3595) );
  XOR U4692 ( .A(n3594), .B(n3595), .Z(n3615) );
  NANDN U4693 ( .A(n3422), .B(n3421), .Z(n3426) );
  NAND U4694 ( .A(n3424), .B(n3423), .Z(n3425) );
  NAND U4695 ( .A(n3426), .B(n3425), .Z(n3612) );
  NANDN U4696 ( .A(n3428), .B(n3427), .Z(n3432) );
  NAND U4697 ( .A(n3430), .B(n3429), .Z(n3431) );
  NAND U4698 ( .A(n3432), .B(n3431), .Z(n3583) );
  XNOR U4699 ( .A(n1052), .B(a[24]), .Z(n3544) );
  NAND U4700 ( .A(n36925), .B(n3544), .Z(n3435) );
  NANDN U4701 ( .A(n3433), .B(n36926), .Z(n3434) );
  NAND U4702 ( .A(n3435), .B(n3434), .Z(n3522) );
  XNOR U4703 ( .A(b[31]), .B(a[2]), .Z(n3562) );
  NANDN U4704 ( .A(n3562), .B(n38552), .Z(n3438) );
  NANDN U4705 ( .A(n3436), .B(n38553), .Z(n3437) );
  NAND U4706 ( .A(n3438), .B(n3437), .Z(n3519) );
  NANDN U4707 ( .A(n3439), .B(n38205), .Z(n3441) );
  XNOR U4708 ( .A(b[23]), .B(a[10]), .Z(n3501) );
  OR U4709 ( .A(n3501), .B(n38268), .Z(n3440) );
  AND U4710 ( .A(n3441), .B(n3440), .Z(n3520) );
  XNOR U4711 ( .A(n3519), .B(n3520), .Z(n3521) );
  XNOR U4712 ( .A(n3522), .B(n3521), .Z(n3602) );
  NANDN U4713 ( .A(n3443), .B(n3442), .Z(n3447) );
  NAND U4714 ( .A(n3445), .B(n3444), .Z(n3446) );
  NAND U4715 ( .A(n3447), .B(n3446), .Z(n3603) );
  XNOR U4716 ( .A(n3602), .B(n3603), .Z(n3604) );
  NAND U4717 ( .A(n3449), .B(n3448), .Z(n3533) );
  XNOR U4718 ( .A(b[17]), .B(a[16]), .Z(n3556) );
  NANDN U4719 ( .A(n3556), .B(n37764), .Z(n3452) );
  NAND U4720 ( .A(n3450), .B(n37762), .Z(n3451) );
  NAND U4721 ( .A(n3452), .B(n3451), .Z(n3532) );
  XOR U4722 ( .A(b[3]), .B(n7434), .Z(n3541) );
  NANDN U4723 ( .A(n3541), .B(n36107), .Z(n3455) );
  OR U4724 ( .A(n3453), .B(n36105), .Z(n3454) );
  AND U4725 ( .A(n3455), .B(n3454), .Z(n3531) );
  XNOR U4726 ( .A(n3532), .B(n3531), .Z(n3534) );
  XNOR U4727 ( .A(n3533), .B(n3534), .Z(n3605) );
  XNOR U4728 ( .A(n3604), .B(n3605), .Z(n3581) );
  XOR U4729 ( .A(b[11]), .B(a[22]), .Z(n3547) );
  NANDN U4730 ( .A(n37311), .B(n3547), .Z(n3458) );
  NAND U4731 ( .A(n3456), .B(n37218), .Z(n3457) );
  NAND U4732 ( .A(n3458), .B(n3457), .Z(n3577) );
  XOR U4733 ( .A(b[25]), .B(a[8]), .Z(n3568) );
  NAND U4734 ( .A(n3568), .B(n38325), .Z(n3461) );
  NAND U4735 ( .A(n3459), .B(n38326), .Z(n3460) );
  NAND U4736 ( .A(n3461), .B(n3460), .Z(n3574) );
  XNOR U4737 ( .A(b[27]), .B(a[6]), .Z(n3559) );
  NANDN U4738 ( .A(n3559), .B(n38423), .Z(n3464) );
  NAND U4739 ( .A(n3462), .B(n38424), .Z(n3463) );
  AND U4740 ( .A(n3464), .B(n3463), .Z(n3575) );
  XNOR U4741 ( .A(n3574), .B(n3575), .Z(n3576) );
  XNOR U4742 ( .A(n3577), .B(n3576), .Z(n3608) );
  XNOR U4743 ( .A(b[7]), .B(n7202), .Z(n3550) );
  NAND U4744 ( .A(n3550), .B(n36701), .Z(n3467) );
  NANDN U4745 ( .A(n3465), .B(n36702), .Z(n3466) );
  NAND U4746 ( .A(n3467), .B(n3466), .Z(n3516) );
  XNOR U4747 ( .A(n1051), .B(a[28]), .Z(n3553) );
  NAND U4748 ( .A(n3553), .B(n36587), .Z(n3470) );
  NANDN U4749 ( .A(n3468), .B(n36588), .Z(n3469) );
  NAND U4750 ( .A(n3470), .B(n3469), .Z(n3513) );
  XNOR U4751 ( .A(b[19]), .B(a[14]), .Z(n3504) );
  NANDN U4752 ( .A(n3504), .B(n37934), .Z(n3473) );
  NANDN U4753 ( .A(n3471), .B(n37935), .Z(n3472) );
  AND U4754 ( .A(n3473), .B(n3472), .Z(n3514) );
  XNOR U4755 ( .A(n3513), .B(n3514), .Z(n3515) );
  XOR U4756 ( .A(n3516), .B(n3515), .Z(n3609) );
  XNOR U4757 ( .A(n3608), .B(n3609), .Z(n3610) );
  NANDN U4758 ( .A(n3475), .B(n3474), .Z(n3479) );
  NAND U4759 ( .A(n3477), .B(n3476), .Z(n3478) );
  AND U4760 ( .A(n3479), .B(n3478), .Z(n3611) );
  XNOR U4761 ( .A(n3610), .B(n3611), .Z(n3580) );
  XOR U4762 ( .A(n3581), .B(n3580), .Z(n3582) );
  XNOR U4763 ( .A(n3583), .B(n3582), .Z(n3613) );
  XNOR U4764 ( .A(n3612), .B(n3613), .Z(n3614) );
  XOR U4765 ( .A(n3615), .B(n3614), .Z(n3589) );
  XOR U4766 ( .A(n3588), .B(n3589), .Z(n3618) );
  XOR U4767 ( .A(n3619), .B(n3618), .Z(n3620) );
  XNOR U4768 ( .A(n3621), .B(n3620), .Z(n3486) );
  NANDN U4769 ( .A(n3481), .B(n3480), .Z(n3485) );
  NANDN U4770 ( .A(n3483), .B(n3482), .Z(n3484) );
  AND U4771 ( .A(n3485), .B(n3484), .Z(n3487) );
  XNOR U4772 ( .A(n3486), .B(n3487), .Z(n3488) );
  XOR U4773 ( .A(n3489), .B(n3488), .Z(n3625) );
  XOR U4774 ( .A(n3626), .B(n3625), .Z(c[256]) );
  NANDN U4775 ( .A(n3487), .B(n3486), .Z(n3491) );
  NAND U4776 ( .A(n3489), .B(n3488), .Z(n3490) );
  NAND U4777 ( .A(n3491), .B(n3490), .Z(n3632) );
  NANDN U4778 ( .A(n3493), .B(n3492), .Z(n3497) );
  OR U4779 ( .A(n3495), .B(n3494), .Z(n3496) );
  NAND U4780 ( .A(n3497), .B(n3496), .Z(n3646) );
  XNOR U4781 ( .A(n1056), .B(a[13]), .Z(n3715) );
  NAND U4782 ( .A(n3715), .B(n38101), .Z(n3500) );
  NANDN U4783 ( .A(n3498), .B(n38102), .Z(n3499) );
  NAND U4784 ( .A(n3500), .B(n3499), .Z(n3748) );
  NANDN U4785 ( .A(n3501), .B(n38205), .Z(n3503) );
  XNOR U4786 ( .A(b[23]), .B(a[11]), .Z(n3730) );
  OR U4787 ( .A(n3730), .B(n38268), .Z(n3502) );
  NAND U4788 ( .A(n3503), .B(n3502), .Z(n3745) );
  XNOR U4789 ( .A(b[19]), .B(a[15]), .Z(n3688) );
  NANDN U4790 ( .A(n3688), .B(n37934), .Z(n3506) );
  NANDN U4791 ( .A(n3504), .B(n37935), .Z(n3505) );
  AND U4792 ( .A(n3506), .B(n3505), .Z(n3746) );
  XNOR U4793 ( .A(n3745), .B(n3746), .Z(n3747) );
  XNOR U4794 ( .A(n3748), .B(n3747), .Z(n3651) );
  XNOR U4795 ( .A(n1054), .B(a[19]), .Z(n3712) );
  NANDN U4796 ( .A(n37665), .B(n3712), .Z(n3509) );
  NANDN U4797 ( .A(n3507), .B(n37604), .Z(n3508) );
  NAND U4798 ( .A(n3509), .B(n3508), .Z(n3676) );
  NAND U4799 ( .A(n38490), .B(n3510), .Z(n3512) );
  XNOR U4800 ( .A(n1058), .B(a[5]), .Z(n3724) );
  NANDN U4801 ( .A(n1048), .B(n3724), .Z(n3511) );
  NAND U4802 ( .A(n3512), .B(n3511), .Z(n3673) );
  NANDN U4803 ( .A(n1059), .B(a[1]), .Z(n3674) );
  XNOR U4804 ( .A(n3673), .B(n3674), .Z(n3675) );
  XOR U4805 ( .A(n3676), .B(n3675), .Z(n3652) );
  XNOR U4806 ( .A(n3651), .B(n3652), .Z(n3653) );
  NANDN U4807 ( .A(n3514), .B(n3513), .Z(n3518) );
  NAND U4808 ( .A(n3516), .B(n3515), .Z(n3517) );
  NAND U4809 ( .A(n3518), .B(n3517), .Z(n3654) );
  XOR U4810 ( .A(n3653), .B(n3654), .Z(n3706) );
  NANDN U4811 ( .A(n3520), .B(n3519), .Z(n3524) );
  NAND U4812 ( .A(n3522), .B(n3521), .Z(n3523) );
  NAND U4813 ( .A(n3524), .B(n3523), .Z(n3703) );
  NANDN U4814 ( .A(n3526), .B(n3525), .Z(n3530) );
  OR U4815 ( .A(n3528), .B(n3527), .Z(n3529) );
  AND U4816 ( .A(n3530), .B(n3529), .Z(n3704) );
  XNOR U4817 ( .A(n3703), .B(n3704), .Z(n3705) );
  XNOR U4818 ( .A(n3706), .B(n3705), .Z(n3760) );
  NANDN U4819 ( .A(n3536), .B(n3535), .Z(n3540) );
  NAND U4820 ( .A(n3538), .B(n3537), .Z(n3539) );
  NAND U4821 ( .A(n3540), .B(n3539), .Z(n3700) );
  XOR U4822 ( .A(b[3]), .B(n7955), .Z(n3685) );
  NANDN U4823 ( .A(n3685), .B(n36107), .Z(n3543) );
  OR U4824 ( .A(n3541), .B(n36105), .Z(n3542) );
  NAND U4825 ( .A(n3543), .B(n3542), .Z(n3671) );
  XOR U4826 ( .A(n1052), .B(a[25]), .Z(n3709) );
  NANDN U4827 ( .A(n3709), .B(n36925), .Z(n3546) );
  NAND U4828 ( .A(n36926), .B(n3544), .Z(n3545) );
  NAND U4829 ( .A(n3546), .B(n3545), .Z(n3669) );
  XNOR U4830 ( .A(b[11]), .B(a[23]), .Z(n3718) );
  OR U4831 ( .A(n3718), .B(n37311), .Z(n3549) );
  NAND U4832 ( .A(n37218), .B(n3547), .Z(n3548) );
  NAND U4833 ( .A(n3549), .B(n3548), .Z(n3670) );
  XNOR U4834 ( .A(n3669), .B(n3670), .Z(n3672) );
  XOR U4835 ( .A(n3671), .B(n3672), .Z(n3660) );
  XOR U4836 ( .A(b[7]), .B(a[27]), .Z(n3733) );
  NAND U4837 ( .A(n36701), .B(n3733), .Z(n3552) );
  NAND U4838 ( .A(n36702), .B(n3550), .Z(n3551) );
  NAND U4839 ( .A(n3552), .B(n3551), .Z(n3658) );
  XNOR U4840 ( .A(b[5]), .B(a[29]), .Z(n3694) );
  NANDN U4841 ( .A(n3694), .B(n36587), .Z(n3555) );
  NAND U4842 ( .A(n36588), .B(n3553), .Z(n3554) );
  AND U4843 ( .A(n3555), .B(n3554), .Z(n3657) );
  XNOR U4844 ( .A(n3658), .B(n3657), .Z(n3659) );
  XNOR U4845 ( .A(n3660), .B(n3659), .Z(n3753) );
  NANDN U4846 ( .A(n3556), .B(n37762), .Z(n3558) );
  XOR U4847 ( .A(b[17]), .B(a[17]), .Z(n3679) );
  NAND U4848 ( .A(n3679), .B(n37764), .Z(n3557) );
  NAND U4849 ( .A(n3558), .B(n3557), .Z(n3666) );
  XOR U4850 ( .A(b[27]), .B(a[7]), .Z(n3691) );
  NAND U4851 ( .A(n38423), .B(n3691), .Z(n3561) );
  NANDN U4852 ( .A(n3559), .B(n38424), .Z(n3560) );
  NAND U4853 ( .A(n3561), .B(n3560), .Z(n3663) );
  XNOR U4854 ( .A(n1059), .B(a[3]), .Z(n3682) );
  NAND U4855 ( .A(n3682), .B(n38552), .Z(n3564) );
  NANDN U4856 ( .A(n3562), .B(n38553), .Z(n3563) );
  AND U4857 ( .A(n3564), .B(n3563), .Z(n3664) );
  XNOR U4858 ( .A(n3663), .B(n3664), .Z(n3665) );
  XNOR U4859 ( .A(n3666), .B(n3665), .Z(n3751) );
  NANDN U4860 ( .A(n1049), .B(a[33]), .Z(n3565) );
  XNOR U4861 ( .A(b[1]), .B(n3565), .Z(n3567) );
  NANDN U4862 ( .A(b[0]), .B(a[32]), .Z(n3566) );
  AND U4863 ( .A(n3567), .B(n3566), .Z(n3740) );
  XOR U4864 ( .A(b[25]), .B(a[9]), .Z(n3736) );
  NAND U4865 ( .A(n38325), .B(n3736), .Z(n3570) );
  NAND U4866 ( .A(n38326), .B(n3568), .Z(n3569) );
  AND U4867 ( .A(n3570), .B(n3569), .Z(n3739) );
  XNOR U4868 ( .A(n3740), .B(n3739), .Z(n3741) );
  XNOR U4869 ( .A(b[13]), .B(a[21]), .Z(n3721) );
  NANDN U4870 ( .A(n3721), .B(n37424), .Z(n3573) );
  NAND U4871 ( .A(n37425), .B(n3571), .Z(n3572) );
  AND U4872 ( .A(n3573), .B(n3572), .Z(n3742) );
  XNOR U4873 ( .A(n3741), .B(n3742), .Z(n3752) );
  XOR U4874 ( .A(n3751), .B(n3752), .Z(n3754) );
  XOR U4875 ( .A(n3753), .B(n3754), .Z(n3697) );
  NANDN U4876 ( .A(n3575), .B(n3574), .Z(n3579) );
  NAND U4877 ( .A(n3577), .B(n3576), .Z(n3578) );
  AND U4878 ( .A(n3579), .B(n3578), .Z(n3698) );
  XOR U4879 ( .A(n3700), .B(n3699), .Z(n3758) );
  XNOR U4880 ( .A(n3757), .B(n3758), .Z(n3759) );
  XOR U4881 ( .A(n3760), .B(n3759), .Z(n3645) );
  XOR U4882 ( .A(n3646), .B(n3645), .Z(n3648) );
  NANDN U4883 ( .A(n3581), .B(n3580), .Z(n3585) );
  OR U4884 ( .A(n3583), .B(n3582), .Z(n3584) );
  NAND U4885 ( .A(n3585), .B(n3584), .Z(n3647) );
  XNOR U4886 ( .A(n3648), .B(n3647), .Z(n3636) );
  NANDN U4887 ( .A(n3587), .B(n3586), .Z(n3591) );
  NAND U4888 ( .A(n3589), .B(n3588), .Z(n3590) );
  NAND U4889 ( .A(n3591), .B(n3590), .Z(n3633) );
  NANDN U4890 ( .A(n3597), .B(n3596), .Z(n3601) );
  NAND U4891 ( .A(n3599), .B(n3598), .Z(n3600) );
  NAND U4892 ( .A(n3601), .B(n3600), .Z(n3766) );
  NANDN U4893 ( .A(n3603), .B(n3602), .Z(n3607) );
  NANDN U4894 ( .A(n3605), .B(n3604), .Z(n3606) );
  NAND U4895 ( .A(n3607), .B(n3606), .Z(n3763) );
  XNOR U4896 ( .A(n3763), .B(n3764), .Z(n3765) );
  XNOR U4897 ( .A(n3766), .B(n3765), .Z(n3639) );
  XNOR U4898 ( .A(n3640), .B(n3639), .Z(n3642) );
  NANDN U4899 ( .A(n3613), .B(n3612), .Z(n3617) );
  NAND U4900 ( .A(n3615), .B(n3614), .Z(n3616) );
  NAND U4901 ( .A(n3617), .B(n3616), .Z(n3641) );
  XOR U4902 ( .A(n3642), .B(n3641), .Z(n3634) );
  XNOR U4903 ( .A(n3633), .B(n3634), .Z(n3635) );
  XNOR U4904 ( .A(n3636), .B(n3635), .Z(n3629) );
  NAND U4905 ( .A(n3619), .B(n3618), .Z(n3623) );
  NAND U4906 ( .A(n3621), .B(n3620), .Z(n3622) );
  NAND U4907 ( .A(n3623), .B(n3622), .Z(n3630) );
  XNOR U4908 ( .A(n3629), .B(n3630), .Z(n3631) );
  XNOR U4909 ( .A(n3632), .B(n3631), .Z(n3769) );
  XNOR U4910 ( .A(n3769), .B(sreg[257]), .Z(n3771) );
  NAND U4911 ( .A(n3624), .B(sreg[256]), .Z(n3628) );
  OR U4912 ( .A(n3626), .B(n3625), .Z(n3627) );
  AND U4913 ( .A(n3628), .B(n3627), .Z(n3770) );
  XOR U4914 ( .A(n3771), .B(n3770), .Z(c[257]) );
  NANDN U4915 ( .A(n3634), .B(n3633), .Z(n3638) );
  NAND U4916 ( .A(n3636), .B(n3635), .Z(n3637) );
  NAND U4917 ( .A(n3638), .B(n3637), .Z(n3775) );
  NAND U4918 ( .A(n3640), .B(n3639), .Z(n3644) );
  OR U4919 ( .A(n3642), .B(n3641), .Z(n3643) );
  NAND U4920 ( .A(n3644), .B(n3643), .Z(n3778) );
  NANDN U4921 ( .A(n3646), .B(n3645), .Z(n3650) );
  OR U4922 ( .A(n3648), .B(n3647), .Z(n3649) );
  AND U4923 ( .A(n3650), .B(n3649), .Z(n3779) );
  XNOR U4924 ( .A(n3778), .B(n3779), .Z(n3780) );
  NANDN U4925 ( .A(n3652), .B(n3651), .Z(n3656) );
  NANDN U4926 ( .A(n3654), .B(n3653), .Z(n3655) );
  NAND U4927 ( .A(n3656), .B(n3655), .Z(n3793) );
  NANDN U4928 ( .A(n3658), .B(n3657), .Z(n3662) );
  NAND U4929 ( .A(n3660), .B(n3659), .Z(n3661) );
  NAND U4930 ( .A(n3662), .B(n3661), .Z(n3892) );
  NANDN U4931 ( .A(n3664), .B(n3663), .Z(n3668) );
  NAND U4932 ( .A(n3666), .B(n3665), .Z(n3667) );
  NAND U4933 ( .A(n3668), .B(n3667), .Z(n3891) );
  XNOR U4934 ( .A(n3891), .B(n3890), .Z(n3893) );
  XOR U4935 ( .A(n3892), .B(n3893), .Z(n3790) );
  NANDN U4936 ( .A(n3674), .B(n3673), .Z(n3678) );
  NAND U4937 ( .A(n3676), .B(n3675), .Z(n3677) );
  NAND U4938 ( .A(n3678), .B(n3677), .Z(n3887) );
  XNOR U4939 ( .A(b[17]), .B(a[18]), .Z(n3809) );
  NANDN U4940 ( .A(n3809), .B(n37764), .Z(n3681) );
  NAND U4941 ( .A(n3679), .B(n37762), .Z(n3680) );
  NAND U4942 ( .A(n3681), .B(n3680), .Z(n3824) );
  XNOR U4943 ( .A(b[31]), .B(a[4]), .Z(n3812) );
  NANDN U4944 ( .A(n3812), .B(n38552), .Z(n3684) );
  NAND U4945 ( .A(n38553), .B(n3682), .Z(n3683) );
  NAND U4946 ( .A(n3684), .B(n3683), .Z(n3822) );
  XNOR U4947 ( .A(b[3]), .B(a[32]), .Z(n3815) );
  NANDN U4948 ( .A(n3815), .B(n36107), .Z(n3687) );
  OR U4949 ( .A(n3685), .B(n36105), .Z(n3686) );
  NAND U4950 ( .A(n3687), .B(n3686), .Z(n3823) );
  XNOR U4951 ( .A(n3822), .B(n3823), .Z(n3825) );
  XOR U4952 ( .A(n3824), .B(n3825), .Z(n3884) );
  XNOR U4953 ( .A(b[19]), .B(a[16]), .Z(n3800) );
  NANDN U4954 ( .A(n3800), .B(n37934), .Z(n3690) );
  NANDN U4955 ( .A(n3688), .B(n37935), .Z(n3689) );
  NAND U4956 ( .A(n3690), .B(n3689), .Z(n3851) );
  XOR U4957 ( .A(b[27]), .B(a[8]), .Z(n3803) );
  NAND U4958 ( .A(n38423), .B(n3803), .Z(n3693) );
  NAND U4959 ( .A(n3691), .B(n38424), .Z(n3692) );
  NAND U4960 ( .A(n3693), .B(n3692), .Z(n3848) );
  XOR U4961 ( .A(b[5]), .B(n7434), .Z(n3806) );
  NANDN U4962 ( .A(n3806), .B(n36587), .Z(n3696) );
  NANDN U4963 ( .A(n3694), .B(n36588), .Z(n3695) );
  AND U4964 ( .A(n3696), .B(n3695), .Z(n3849) );
  XNOR U4965 ( .A(n3848), .B(n3849), .Z(n3850) );
  XOR U4966 ( .A(n3851), .B(n3850), .Z(n3885) );
  XNOR U4967 ( .A(n3884), .B(n3885), .Z(n3886) );
  XOR U4968 ( .A(n3887), .B(n3886), .Z(n3791) );
  XNOR U4969 ( .A(n3790), .B(n3791), .Z(n3792) );
  XNOR U4970 ( .A(n3793), .B(n3792), .Z(n3903) );
  OR U4971 ( .A(n3698), .B(n3697), .Z(n3702) );
  NAND U4972 ( .A(n3700), .B(n3699), .Z(n3701) );
  AND U4973 ( .A(n3702), .B(n3701), .Z(n3900) );
  NANDN U4974 ( .A(n3704), .B(n3703), .Z(n3708) );
  NAND U4975 ( .A(n3706), .B(n3705), .Z(n3707) );
  NAND U4976 ( .A(n3708), .B(n3707), .Z(n3787) );
  XOR U4977 ( .A(b[9]), .B(n7202), .Z(n3854) );
  NANDN U4978 ( .A(n3854), .B(n36925), .Z(n3711) );
  NANDN U4979 ( .A(n3709), .B(n36926), .Z(n3710) );
  NAND U4980 ( .A(n3711), .B(n3710), .Z(n3828) );
  XNOR U4981 ( .A(n1054), .B(a[20]), .Z(n3857) );
  NANDN U4982 ( .A(n37665), .B(n3857), .Z(n3714) );
  NAND U4983 ( .A(n3712), .B(n37604), .Z(n3713) );
  NAND U4984 ( .A(n3714), .B(n3713), .Z(n3826) );
  XNOR U4985 ( .A(b[21]), .B(a[14]), .Z(n3860) );
  NANDN U4986 ( .A(n3860), .B(n38101), .Z(n3717) );
  NAND U4987 ( .A(n3715), .B(n38102), .Z(n3716) );
  AND U4988 ( .A(n3717), .B(n3716), .Z(n3827) );
  XNOR U4989 ( .A(n3826), .B(n3827), .Z(n3829) );
  XOR U4990 ( .A(n3828), .B(n3829), .Z(n3821) );
  XNOR U4991 ( .A(b[11]), .B(a[24]), .Z(n3863) );
  OR U4992 ( .A(n3863), .B(n37311), .Z(n3720) );
  NANDN U4993 ( .A(n3718), .B(n37218), .Z(n3719) );
  NAND U4994 ( .A(n3720), .B(n3719), .Z(n3819) );
  XNOR U4995 ( .A(n1053), .B(a[22]), .Z(n3866) );
  NAND U4996 ( .A(n3866), .B(n37424), .Z(n3723) );
  NANDN U4997 ( .A(n3721), .B(n37425), .Z(n3722) );
  AND U4998 ( .A(n3723), .B(n3722), .Z(n3818) );
  XNOR U4999 ( .A(n3819), .B(n3818), .Z(n3820) );
  XOR U5000 ( .A(n3821), .B(n3820), .Z(n3833) );
  NAND U5001 ( .A(n38490), .B(n3724), .Z(n3726) );
  XOR U5002 ( .A(n1058), .B(n4305), .Z(n3872) );
  NANDN U5003 ( .A(n1048), .B(n3872), .Z(n3725) );
  NAND U5004 ( .A(n3726), .B(n3725), .Z(n3794) );
  NANDN U5005 ( .A(n1059), .B(a[2]), .Z(n3795) );
  XNOR U5006 ( .A(n3794), .B(n3795), .Z(n3797) );
  NANDN U5007 ( .A(n1049), .B(a[34]), .Z(n3727) );
  XNOR U5008 ( .A(b[1]), .B(n3727), .Z(n3729) );
  NANDN U5009 ( .A(b[0]), .B(a[33]), .Z(n3728) );
  AND U5010 ( .A(n3729), .B(n3728), .Z(n3796) );
  XOR U5011 ( .A(n3797), .B(n3796), .Z(n3830) );
  NANDN U5012 ( .A(n3730), .B(n38205), .Z(n3732) );
  XNOR U5013 ( .A(b[23]), .B(a[12]), .Z(n3875) );
  OR U5014 ( .A(n3875), .B(n38268), .Z(n3731) );
  NAND U5015 ( .A(n3732), .B(n3731), .Z(n3845) );
  XOR U5016 ( .A(b[7]), .B(a[28]), .Z(n3878) );
  NAND U5017 ( .A(n3878), .B(n36701), .Z(n3735) );
  NAND U5018 ( .A(n3733), .B(n36702), .Z(n3734) );
  NAND U5019 ( .A(n3735), .B(n3734), .Z(n3842) );
  XOR U5020 ( .A(b[25]), .B(a[10]), .Z(n3881) );
  NAND U5021 ( .A(n3881), .B(n38325), .Z(n3738) );
  NAND U5022 ( .A(n3736), .B(n38326), .Z(n3737) );
  AND U5023 ( .A(n3738), .B(n3737), .Z(n3843) );
  XNOR U5024 ( .A(n3842), .B(n3843), .Z(n3844) );
  XNOR U5025 ( .A(n3845), .B(n3844), .Z(n3831) );
  XNOR U5026 ( .A(n3830), .B(n3831), .Z(n3832) );
  XNOR U5027 ( .A(n3833), .B(n3832), .Z(n3839) );
  NANDN U5028 ( .A(n3740), .B(n3739), .Z(n3744) );
  NAND U5029 ( .A(n3742), .B(n3741), .Z(n3743) );
  NAND U5030 ( .A(n3744), .B(n3743), .Z(n3836) );
  NANDN U5031 ( .A(n3746), .B(n3745), .Z(n3750) );
  NAND U5032 ( .A(n3748), .B(n3747), .Z(n3749) );
  NAND U5033 ( .A(n3750), .B(n3749), .Z(n3837) );
  XNOR U5034 ( .A(n3836), .B(n3837), .Z(n3838) );
  XOR U5035 ( .A(n3839), .B(n3838), .Z(n3784) );
  NANDN U5036 ( .A(n3752), .B(n3751), .Z(n3756) );
  OR U5037 ( .A(n3754), .B(n3753), .Z(n3755) );
  NAND U5038 ( .A(n3756), .B(n3755), .Z(n3785) );
  XOR U5039 ( .A(n3784), .B(n3785), .Z(n3786) );
  XNOR U5040 ( .A(n3787), .B(n3786), .Z(n3901) );
  XOR U5041 ( .A(n3903), .B(n3902), .Z(n3897) );
  NANDN U5042 ( .A(n3758), .B(n3757), .Z(n3762) );
  NAND U5043 ( .A(n3760), .B(n3759), .Z(n3761) );
  NAND U5044 ( .A(n3762), .B(n3761), .Z(n3894) );
  NANDN U5045 ( .A(n3764), .B(n3763), .Z(n3768) );
  NANDN U5046 ( .A(n3766), .B(n3765), .Z(n3767) );
  AND U5047 ( .A(n3768), .B(n3767), .Z(n3895) );
  XNOR U5048 ( .A(n3894), .B(n3895), .Z(n3896) );
  XOR U5049 ( .A(n3897), .B(n3896), .Z(n3781) );
  XNOR U5050 ( .A(n3780), .B(n3781), .Z(n3774) );
  XNOR U5051 ( .A(n3775), .B(n3774), .Z(n3776) );
  XNOR U5052 ( .A(n3777), .B(n3776), .Z(n3906) );
  XNOR U5053 ( .A(n3906), .B(sreg[258]), .Z(n3908) );
  NAND U5054 ( .A(n3769), .B(sreg[257]), .Z(n3773) );
  OR U5055 ( .A(n3771), .B(n3770), .Z(n3772) );
  AND U5056 ( .A(n3773), .B(n3772), .Z(n3907) );
  XOR U5057 ( .A(n3908), .B(n3907), .Z(c[258]) );
  NANDN U5058 ( .A(n3779), .B(n3778), .Z(n3783) );
  NANDN U5059 ( .A(n3781), .B(n3780), .Z(n3782) );
  NAND U5060 ( .A(n3783), .B(n3782), .Z(n3911) );
  OR U5061 ( .A(n3785), .B(n3784), .Z(n3789) );
  NAND U5062 ( .A(n3787), .B(n3786), .Z(n3788) );
  NAND U5063 ( .A(n3789), .B(n3788), .Z(n4037) );
  XNOR U5064 ( .A(n4037), .B(n4038), .Z(n4039) );
  NANDN U5065 ( .A(n3795), .B(n3794), .Z(n3799) );
  NAND U5066 ( .A(n3797), .B(n3796), .Z(n3798) );
  NAND U5067 ( .A(n3799), .B(n3798), .Z(n3994) );
  XNOR U5068 ( .A(b[19]), .B(a[17]), .Z(n3939) );
  NANDN U5069 ( .A(n3939), .B(n37934), .Z(n3802) );
  NANDN U5070 ( .A(n3800), .B(n37935), .Z(n3801) );
  NAND U5071 ( .A(n3802), .B(n3801), .Z(n4004) );
  XOR U5072 ( .A(b[27]), .B(a[9]), .Z(n3942) );
  NAND U5073 ( .A(n38423), .B(n3942), .Z(n3805) );
  NAND U5074 ( .A(n3803), .B(n38424), .Z(n3804) );
  NAND U5075 ( .A(n3805), .B(n3804), .Z(n4001) );
  XOR U5076 ( .A(b[5]), .B(n7955), .Z(n3945) );
  NANDN U5077 ( .A(n3945), .B(n36587), .Z(n3808) );
  NANDN U5078 ( .A(n3806), .B(n36588), .Z(n3807) );
  AND U5079 ( .A(n3808), .B(n3807), .Z(n4002) );
  XNOR U5080 ( .A(n4001), .B(n4002), .Z(n4003) );
  XNOR U5081 ( .A(n4004), .B(n4003), .Z(n3992) );
  NANDN U5082 ( .A(n3809), .B(n37762), .Z(n3811) );
  XOR U5083 ( .A(b[17]), .B(a[19]), .Z(n3948) );
  NAND U5084 ( .A(n3948), .B(n37764), .Z(n3810) );
  NAND U5085 ( .A(n3811), .B(n3810), .Z(n3966) );
  XNOR U5086 ( .A(b[31]), .B(a[5]), .Z(n3951) );
  NANDN U5087 ( .A(n3951), .B(n38552), .Z(n3814) );
  NANDN U5088 ( .A(n3812), .B(n38553), .Z(n3813) );
  NAND U5089 ( .A(n3814), .B(n3813), .Z(n3963) );
  OR U5090 ( .A(n3815), .B(n36105), .Z(n3817) );
  XNOR U5091 ( .A(b[3]), .B(a[33]), .Z(n3954) );
  NANDN U5092 ( .A(n3954), .B(n36107), .Z(n3816) );
  AND U5093 ( .A(n3817), .B(n3816), .Z(n3964) );
  XNOR U5094 ( .A(n3963), .B(n3964), .Z(n3965) );
  XOR U5095 ( .A(n3966), .B(n3965), .Z(n3991) );
  XNOR U5096 ( .A(n3992), .B(n3991), .Z(n3993) );
  XNOR U5097 ( .A(n3994), .B(n3993), .Z(n3930) );
  XNOR U5098 ( .A(n3982), .B(n3981), .Z(n3984) );
  XOR U5099 ( .A(n3983), .B(n3984), .Z(n3929) );
  XOR U5100 ( .A(n3930), .B(n3929), .Z(n3931) );
  NANDN U5101 ( .A(n3831), .B(n3830), .Z(n3835) );
  NAND U5102 ( .A(n3833), .B(n3832), .Z(n3834) );
  AND U5103 ( .A(n3835), .B(n3834), .Z(n3932) );
  XOR U5104 ( .A(n3931), .B(n3932), .Z(n4045) );
  NANDN U5105 ( .A(n3837), .B(n3836), .Z(n3841) );
  NAND U5106 ( .A(n3839), .B(n3838), .Z(n3840) );
  NAND U5107 ( .A(n3841), .B(n3840), .Z(n3926) );
  NANDN U5108 ( .A(n3843), .B(n3842), .Z(n3847) );
  NAND U5109 ( .A(n3845), .B(n3844), .Z(n3846) );
  NAND U5110 ( .A(n3847), .B(n3846), .Z(n3985) );
  NANDN U5111 ( .A(n3849), .B(n3848), .Z(n3853) );
  NAND U5112 ( .A(n3851), .B(n3850), .Z(n3852) );
  AND U5113 ( .A(n3853), .B(n3852), .Z(n3986) );
  XNOR U5114 ( .A(n3985), .B(n3986), .Z(n3987) );
  XNOR U5115 ( .A(b[9]), .B(a[27]), .Z(n4007) );
  NANDN U5116 ( .A(n4007), .B(n36925), .Z(n3856) );
  NANDN U5117 ( .A(n3854), .B(n36926), .Z(n3855) );
  NAND U5118 ( .A(n3856), .B(n3855), .Z(n3971) );
  XNOR U5119 ( .A(b[15]), .B(a[21]), .Z(n4010) );
  OR U5120 ( .A(n4010), .B(n37665), .Z(n3859) );
  NAND U5121 ( .A(n3857), .B(n37604), .Z(n3858) );
  AND U5122 ( .A(n3859), .B(n3858), .Z(n3969) );
  XNOR U5123 ( .A(b[21]), .B(a[15]), .Z(n4013) );
  NANDN U5124 ( .A(n4013), .B(n38101), .Z(n3862) );
  NANDN U5125 ( .A(n3860), .B(n38102), .Z(n3861) );
  AND U5126 ( .A(n3862), .B(n3861), .Z(n3970) );
  XOR U5127 ( .A(n3971), .B(n3972), .Z(n3960) );
  XOR U5128 ( .A(b[11]), .B(n7069), .Z(n4016) );
  OR U5129 ( .A(n4016), .B(n37311), .Z(n3865) );
  NANDN U5130 ( .A(n3863), .B(n37218), .Z(n3864) );
  NAND U5131 ( .A(n3865), .B(n3864), .Z(n3958) );
  XOR U5132 ( .A(n1053), .B(a[23]), .Z(n4019) );
  NANDN U5133 ( .A(n4019), .B(n37424), .Z(n3868) );
  NAND U5134 ( .A(n37425), .B(n3866), .Z(n3867) );
  AND U5135 ( .A(n3868), .B(n3867), .Z(n3957) );
  XNOR U5136 ( .A(n3958), .B(n3957), .Z(n3959) );
  XOR U5137 ( .A(n3960), .B(n3959), .Z(n3977) );
  NANDN U5138 ( .A(n1049), .B(a[35]), .Z(n3869) );
  XNOR U5139 ( .A(b[1]), .B(n3869), .Z(n3871) );
  NANDN U5140 ( .A(b[0]), .B(a[34]), .Z(n3870) );
  AND U5141 ( .A(n3871), .B(n3870), .Z(n3935) );
  NAND U5142 ( .A(n38490), .B(n3872), .Z(n3874) );
  XNOR U5143 ( .A(n1058), .B(a[7]), .Z(n4025) );
  NANDN U5144 ( .A(n1048), .B(n4025), .Z(n3873) );
  NAND U5145 ( .A(n3874), .B(n3873), .Z(n3933) );
  NANDN U5146 ( .A(n1059), .B(a[3]), .Z(n3934) );
  XNOR U5147 ( .A(n3933), .B(n3934), .Z(n3936) );
  XOR U5148 ( .A(n3935), .B(n3936), .Z(n3975) );
  NANDN U5149 ( .A(n3875), .B(n38205), .Z(n3877) );
  XNOR U5150 ( .A(b[23]), .B(a[13]), .Z(n4028) );
  OR U5151 ( .A(n4028), .B(n38268), .Z(n3876) );
  NAND U5152 ( .A(n3877), .B(n3876), .Z(n3998) );
  XOR U5153 ( .A(b[7]), .B(a[29]), .Z(n4031) );
  NAND U5154 ( .A(n4031), .B(n36701), .Z(n3880) );
  NAND U5155 ( .A(n3878), .B(n36702), .Z(n3879) );
  NAND U5156 ( .A(n3880), .B(n3879), .Z(n3995) );
  XOR U5157 ( .A(b[25]), .B(a[11]), .Z(n4034) );
  NAND U5158 ( .A(n4034), .B(n38325), .Z(n3883) );
  NAND U5159 ( .A(n3881), .B(n38326), .Z(n3882) );
  AND U5160 ( .A(n3883), .B(n3882), .Z(n3996) );
  XNOR U5161 ( .A(n3995), .B(n3996), .Z(n3997) );
  XNOR U5162 ( .A(n3998), .B(n3997), .Z(n3976) );
  XOR U5163 ( .A(n3975), .B(n3976), .Z(n3978) );
  XNOR U5164 ( .A(n3977), .B(n3978), .Z(n3988) );
  XOR U5165 ( .A(n3987), .B(n3988), .Z(n3923) );
  NANDN U5166 ( .A(n3885), .B(n3884), .Z(n3889) );
  NANDN U5167 ( .A(n3887), .B(n3886), .Z(n3888) );
  AND U5168 ( .A(n3889), .B(n3888), .Z(n3924) );
  XNOR U5169 ( .A(n3923), .B(n3924), .Z(n3925) );
  XOR U5170 ( .A(n3926), .B(n3925), .Z(n4043) );
  XNOR U5171 ( .A(n4043), .B(n4044), .Z(n4046) );
  XNOR U5172 ( .A(n4045), .B(n4046), .Z(n4040) );
  XOR U5173 ( .A(n4039), .B(n4040), .Z(n3920) );
  NANDN U5174 ( .A(n3895), .B(n3894), .Z(n3899) );
  NANDN U5175 ( .A(n3897), .B(n3896), .Z(n3898) );
  NAND U5176 ( .A(n3899), .B(n3898), .Z(n3917) );
  OR U5177 ( .A(n3901), .B(n3900), .Z(n3905) );
  NAND U5178 ( .A(n3903), .B(n3902), .Z(n3904) );
  NAND U5179 ( .A(n3905), .B(n3904), .Z(n3918) );
  XNOR U5180 ( .A(n3917), .B(n3918), .Z(n3919) );
  XNOR U5181 ( .A(n3920), .B(n3919), .Z(n3912) );
  XNOR U5182 ( .A(n3911), .B(n3912), .Z(n3913) );
  XNOR U5183 ( .A(n3914), .B(n3913), .Z(n4049) );
  XNOR U5184 ( .A(n4049), .B(sreg[259]), .Z(n4051) );
  NAND U5185 ( .A(n3906), .B(sreg[258]), .Z(n3910) );
  OR U5186 ( .A(n3908), .B(n3907), .Z(n3909) );
  AND U5187 ( .A(n3910), .B(n3909), .Z(n4050) );
  XOR U5188 ( .A(n4051), .B(n4050), .Z(c[259]) );
  NANDN U5189 ( .A(n3912), .B(n3911), .Z(n3916) );
  NAND U5190 ( .A(n3914), .B(n3913), .Z(n3915) );
  NAND U5191 ( .A(n3916), .B(n3915), .Z(n4057) );
  NANDN U5192 ( .A(n3918), .B(n3917), .Z(n3922) );
  NAND U5193 ( .A(n3920), .B(n3919), .Z(n3921) );
  NAND U5194 ( .A(n3922), .B(n3921), .Z(n4054) );
  NANDN U5195 ( .A(n3924), .B(n3923), .Z(n3928) );
  NAND U5196 ( .A(n3926), .B(n3925), .Z(n3927) );
  NAND U5197 ( .A(n3928), .B(n3927), .Z(n4067) );
  XNOR U5198 ( .A(n4067), .B(n4066), .Z(n4068) );
  NANDN U5199 ( .A(n3934), .B(n3933), .Z(n3938) );
  NAND U5200 ( .A(n3936), .B(n3935), .Z(n3937) );
  NAND U5201 ( .A(n3938), .B(n3937), .Z(n4141) );
  XNOR U5202 ( .A(b[19]), .B(a[18]), .Z(n4084) );
  NANDN U5203 ( .A(n4084), .B(n37934), .Z(n3941) );
  NANDN U5204 ( .A(n3939), .B(n37935), .Z(n3940) );
  NAND U5205 ( .A(n3941), .B(n3940), .Z(n4151) );
  XOR U5206 ( .A(b[27]), .B(a[10]), .Z(n4087) );
  NAND U5207 ( .A(n38423), .B(n4087), .Z(n3944) );
  NAND U5208 ( .A(n3942), .B(n38424), .Z(n3943) );
  NAND U5209 ( .A(n3944), .B(n3943), .Z(n4148) );
  XNOR U5210 ( .A(b[5]), .B(a[32]), .Z(n4090) );
  NANDN U5211 ( .A(n4090), .B(n36587), .Z(n3947) );
  NANDN U5212 ( .A(n3945), .B(n36588), .Z(n3946) );
  AND U5213 ( .A(n3947), .B(n3946), .Z(n4149) );
  XNOR U5214 ( .A(n4148), .B(n4149), .Z(n4150) );
  XNOR U5215 ( .A(n4151), .B(n4150), .Z(n4139) );
  NAND U5216 ( .A(n3948), .B(n37762), .Z(n3950) );
  XOR U5217 ( .A(b[17]), .B(a[20]), .Z(n4093) );
  NAND U5218 ( .A(n4093), .B(n37764), .Z(n3949) );
  NAND U5219 ( .A(n3950), .B(n3949), .Z(n4111) );
  XOR U5220 ( .A(b[31]), .B(n4305), .Z(n4096) );
  NANDN U5221 ( .A(n4096), .B(n38552), .Z(n3953) );
  NANDN U5222 ( .A(n3951), .B(n38553), .Z(n3952) );
  NAND U5223 ( .A(n3953), .B(n3952), .Z(n4108) );
  OR U5224 ( .A(n3954), .B(n36105), .Z(n3956) );
  XNOR U5225 ( .A(b[3]), .B(a[34]), .Z(n4099) );
  NANDN U5226 ( .A(n4099), .B(n36107), .Z(n3955) );
  AND U5227 ( .A(n3956), .B(n3955), .Z(n4109) );
  XNOR U5228 ( .A(n4108), .B(n4109), .Z(n4110) );
  XOR U5229 ( .A(n4111), .B(n4110), .Z(n4138) );
  XNOR U5230 ( .A(n4139), .B(n4138), .Z(n4140) );
  XNOR U5231 ( .A(n4141), .B(n4140), .Z(n4184) );
  NANDN U5232 ( .A(n3958), .B(n3957), .Z(n3962) );
  NAND U5233 ( .A(n3960), .B(n3959), .Z(n3961) );
  NAND U5234 ( .A(n3962), .B(n3961), .Z(n4129) );
  NANDN U5235 ( .A(n3964), .B(n3963), .Z(n3968) );
  NAND U5236 ( .A(n3966), .B(n3965), .Z(n3967) );
  NAND U5237 ( .A(n3968), .B(n3967), .Z(n4127) );
  OR U5238 ( .A(n3970), .B(n3969), .Z(n3974) );
  NANDN U5239 ( .A(n3972), .B(n3971), .Z(n3973) );
  NAND U5240 ( .A(n3974), .B(n3973), .Z(n4126) );
  XNOR U5241 ( .A(n4129), .B(n4128), .Z(n4185) );
  XNOR U5242 ( .A(n4184), .B(n4185), .Z(n4186) );
  NANDN U5243 ( .A(n3976), .B(n3975), .Z(n3980) );
  OR U5244 ( .A(n3978), .B(n3977), .Z(n3979) );
  AND U5245 ( .A(n3980), .B(n3979), .Z(n4187) );
  XOR U5246 ( .A(n4186), .B(n4187), .Z(n4074) );
  NANDN U5247 ( .A(n3986), .B(n3985), .Z(n3990) );
  NANDN U5248 ( .A(n3988), .B(n3987), .Z(n3989) );
  NAND U5249 ( .A(n3990), .B(n3989), .Z(n4193) );
  NANDN U5250 ( .A(n3996), .B(n3995), .Z(n4000) );
  NAND U5251 ( .A(n3998), .B(n3997), .Z(n3999) );
  NAND U5252 ( .A(n4000), .B(n3999), .Z(n4132) );
  NANDN U5253 ( .A(n4002), .B(n4001), .Z(n4006) );
  NAND U5254 ( .A(n4004), .B(n4003), .Z(n4005) );
  AND U5255 ( .A(n4006), .B(n4005), .Z(n4133) );
  XNOR U5256 ( .A(n4132), .B(n4133), .Z(n4134) );
  XNOR U5257 ( .A(n1052), .B(a[28]), .Z(n4154) );
  NAND U5258 ( .A(n36925), .B(n4154), .Z(n4009) );
  NANDN U5259 ( .A(n4007), .B(n36926), .Z(n4008) );
  NAND U5260 ( .A(n4009), .B(n4008), .Z(n4116) );
  XNOR U5261 ( .A(b[15]), .B(a[22]), .Z(n4157) );
  OR U5262 ( .A(n4157), .B(n37665), .Z(n4012) );
  NANDN U5263 ( .A(n4010), .B(n37604), .Z(n4011) );
  AND U5264 ( .A(n4012), .B(n4011), .Z(n4114) );
  XNOR U5265 ( .A(n1056), .B(a[16]), .Z(n4160) );
  NAND U5266 ( .A(n4160), .B(n38101), .Z(n4015) );
  NANDN U5267 ( .A(n4013), .B(n38102), .Z(n4014) );
  AND U5268 ( .A(n4015), .B(n4014), .Z(n4115) );
  XOR U5269 ( .A(n4116), .B(n4117), .Z(n4105) );
  XOR U5270 ( .A(b[11]), .B(n7202), .Z(n4163) );
  OR U5271 ( .A(n4163), .B(n37311), .Z(n4018) );
  NANDN U5272 ( .A(n4016), .B(n37218), .Z(n4017) );
  NAND U5273 ( .A(n4018), .B(n4017), .Z(n4103) );
  XOR U5274 ( .A(n1053), .B(a[24]), .Z(n4166) );
  NANDN U5275 ( .A(n4166), .B(n37424), .Z(n4021) );
  NANDN U5276 ( .A(n4019), .B(n37425), .Z(n4020) );
  AND U5277 ( .A(n4021), .B(n4020), .Z(n4102) );
  XNOR U5278 ( .A(n4103), .B(n4102), .Z(n4104) );
  XOR U5279 ( .A(n4105), .B(n4104), .Z(n4122) );
  NANDN U5280 ( .A(n1049), .B(a[36]), .Z(n4022) );
  XNOR U5281 ( .A(b[1]), .B(n4022), .Z(n4024) );
  NANDN U5282 ( .A(b[0]), .B(a[35]), .Z(n4023) );
  AND U5283 ( .A(n4024), .B(n4023), .Z(n4080) );
  NAND U5284 ( .A(n38490), .B(n4025), .Z(n4027) );
  XNOR U5285 ( .A(n1058), .B(a[8]), .Z(n4172) );
  NANDN U5286 ( .A(n1048), .B(n4172), .Z(n4026) );
  NAND U5287 ( .A(n4027), .B(n4026), .Z(n4078) );
  NANDN U5288 ( .A(n1059), .B(a[4]), .Z(n4079) );
  XNOR U5289 ( .A(n4078), .B(n4079), .Z(n4081) );
  XOR U5290 ( .A(n4080), .B(n4081), .Z(n4120) );
  NANDN U5291 ( .A(n4028), .B(n38205), .Z(n4030) );
  XNOR U5292 ( .A(b[23]), .B(a[14]), .Z(n4175) );
  OR U5293 ( .A(n4175), .B(n38268), .Z(n4029) );
  NAND U5294 ( .A(n4030), .B(n4029), .Z(n4145) );
  XNOR U5295 ( .A(b[7]), .B(a[30]), .Z(n4178) );
  NANDN U5296 ( .A(n4178), .B(n36701), .Z(n4033) );
  NAND U5297 ( .A(n4031), .B(n36702), .Z(n4032) );
  NAND U5298 ( .A(n4033), .B(n4032), .Z(n4142) );
  XOR U5299 ( .A(b[25]), .B(a[12]), .Z(n4181) );
  NAND U5300 ( .A(n4181), .B(n38325), .Z(n4036) );
  NAND U5301 ( .A(n4034), .B(n38326), .Z(n4035) );
  AND U5302 ( .A(n4036), .B(n4035), .Z(n4143) );
  XNOR U5303 ( .A(n4142), .B(n4143), .Z(n4144) );
  XNOR U5304 ( .A(n4145), .B(n4144), .Z(n4121) );
  XOR U5305 ( .A(n4120), .B(n4121), .Z(n4123) );
  XNOR U5306 ( .A(n4122), .B(n4123), .Z(n4135) );
  XOR U5307 ( .A(n4134), .B(n4135), .Z(n4191) );
  XNOR U5308 ( .A(n4190), .B(n4191), .Z(n4192) );
  XNOR U5309 ( .A(n4193), .B(n4192), .Z(n4072) );
  XNOR U5310 ( .A(n4073), .B(n4072), .Z(n4075) );
  XNOR U5311 ( .A(n4074), .B(n4075), .Z(n4069) );
  XOR U5312 ( .A(n4068), .B(n4069), .Z(n4063) );
  NANDN U5313 ( .A(n4038), .B(n4037), .Z(n4042) );
  NANDN U5314 ( .A(n4040), .B(n4039), .Z(n4041) );
  NAND U5315 ( .A(n4042), .B(n4041), .Z(n4061) );
  OR U5316 ( .A(n4044), .B(n4043), .Z(n4048) );
  OR U5317 ( .A(n4046), .B(n4045), .Z(n4047) );
  AND U5318 ( .A(n4048), .B(n4047), .Z(n4060) );
  XNOR U5319 ( .A(n4061), .B(n4060), .Z(n4062) );
  XNOR U5320 ( .A(n4063), .B(n4062), .Z(n4055) );
  XNOR U5321 ( .A(n4054), .B(n4055), .Z(n4056) );
  XNOR U5322 ( .A(n4057), .B(n4056), .Z(n4196) );
  XNOR U5323 ( .A(n4196), .B(sreg[260]), .Z(n4198) );
  NAND U5324 ( .A(n4049), .B(sreg[259]), .Z(n4053) );
  OR U5325 ( .A(n4051), .B(n4050), .Z(n4052) );
  AND U5326 ( .A(n4053), .B(n4052), .Z(n4197) );
  XOR U5327 ( .A(n4198), .B(n4197), .Z(c[260]) );
  NANDN U5328 ( .A(n4055), .B(n4054), .Z(n4059) );
  NAND U5329 ( .A(n4057), .B(n4056), .Z(n4058) );
  NAND U5330 ( .A(n4059), .B(n4058), .Z(n4204) );
  NANDN U5331 ( .A(n4061), .B(n4060), .Z(n4065) );
  NAND U5332 ( .A(n4063), .B(n4062), .Z(n4064) );
  NAND U5333 ( .A(n4065), .B(n4064), .Z(n4202) );
  NANDN U5334 ( .A(n4067), .B(n4066), .Z(n4071) );
  NANDN U5335 ( .A(n4069), .B(n4068), .Z(n4070) );
  NAND U5336 ( .A(n4071), .B(n4070), .Z(n4208) );
  OR U5337 ( .A(n4073), .B(n4072), .Z(n4077) );
  OR U5338 ( .A(n4075), .B(n4074), .Z(n4076) );
  AND U5339 ( .A(n4077), .B(n4076), .Z(n4207) );
  XNOR U5340 ( .A(n4208), .B(n4207), .Z(n4209) );
  NANDN U5341 ( .A(n4079), .B(n4078), .Z(n4083) );
  NAND U5342 ( .A(n4081), .B(n4080), .Z(n4082) );
  NAND U5343 ( .A(n4083), .B(n4082), .Z(n4274) );
  XNOR U5344 ( .A(b[19]), .B(a[19]), .Z(n4219) );
  NANDN U5345 ( .A(n4219), .B(n37934), .Z(n4086) );
  NANDN U5346 ( .A(n4084), .B(n37935), .Z(n4085) );
  NAND U5347 ( .A(n4086), .B(n4085), .Z(n4284) );
  XOR U5348 ( .A(b[27]), .B(a[11]), .Z(n4222) );
  NAND U5349 ( .A(n38423), .B(n4222), .Z(n4089) );
  NAND U5350 ( .A(n4087), .B(n38424), .Z(n4088) );
  NAND U5351 ( .A(n4089), .B(n4088), .Z(n4281) );
  XNOR U5352 ( .A(b[5]), .B(a[33]), .Z(n4225) );
  NANDN U5353 ( .A(n4225), .B(n36587), .Z(n4092) );
  NANDN U5354 ( .A(n4090), .B(n36588), .Z(n4091) );
  AND U5355 ( .A(n4092), .B(n4091), .Z(n4282) );
  XNOR U5356 ( .A(n4281), .B(n4282), .Z(n4283) );
  XNOR U5357 ( .A(n4284), .B(n4283), .Z(n4272) );
  NAND U5358 ( .A(n4093), .B(n37762), .Z(n4095) );
  XOR U5359 ( .A(b[17]), .B(a[21]), .Z(n4228) );
  NAND U5360 ( .A(n4228), .B(n37764), .Z(n4094) );
  NAND U5361 ( .A(n4095), .B(n4094), .Z(n4246) );
  XNOR U5362 ( .A(b[31]), .B(a[7]), .Z(n4231) );
  NANDN U5363 ( .A(n4231), .B(n38552), .Z(n4098) );
  NANDN U5364 ( .A(n4096), .B(n38553), .Z(n4097) );
  NAND U5365 ( .A(n4098), .B(n4097), .Z(n4243) );
  OR U5366 ( .A(n4099), .B(n36105), .Z(n4101) );
  XNOR U5367 ( .A(b[3]), .B(a[35]), .Z(n4234) );
  NANDN U5368 ( .A(n4234), .B(n36107), .Z(n4100) );
  AND U5369 ( .A(n4101), .B(n4100), .Z(n4244) );
  XNOR U5370 ( .A(n4243), .B(n4244), .Z(n4245) );
  XOR U5371 ( .A(n4246), .B(n4245), .Z(n4271) );
  XNOR U5372 ( .A(n4272), .B(n4271), .Z(n4273) );
  XNOR U5373 ( .A(n4274), .B(n4273), .Z(n4318) );
  NANDN U5374 ( .A(n4103), .B(n4102), .Z(n4107) );
  NAND U5375 ( .A(n4105), .B(n4104), .Z(n4106) );
  NAND U5376 ( .A(n4107), .B(n4106), .Z(n4262) );
  NANDN U5377 ( .A(n4109), .B(n4108), .Z(n4113) );
  NAND U5378 ( .A(n4111), .B(n4110), .Z(n4112) );
  NAND U5379 ( .A(n4113), .B(n4112), .Z(n4260) );
  OR U5380 ( .A(n4115), .B(n4114), .Z(n4119) );
  NANDN U5381 ( .A(n4117), .B(n4116), .Z(n4118) );
  NAND U5382 ( .A(n4119), .B(n4118), .Z(n4259) );
  XNOR U5383 ( .A(n4262), .B(n4261), .Z(n4319) );
  XOR U5384 ( .A(n4318), .B(n4319), .Z(n4321) );
  NANDN U5385 ( .A(n4121), .B(n4120), .Z(n4125) );
  OR U5386 ( .A(n4123), .B(n4122), .Z(n4124) );
  NAND U5387 ( .A(n4125), .B(n4124), .Z(n4320) );
  XOR U5388 ( .A(n4321), .B(n4320), .Z(n4338) );
  OR U5389 ( .A(n4127), .B(n4126), .Z(n4131) );
  NAND U5390 ( .A(n4129), .B(n4128), .Z(n4130) );
  NAND U5391 ( .A(n4131), .B(n4130), .Z(n4337) );
  NANDN U5392 ( .A(n4133), .B(n4132), .Z(n4137) );
  NANDN U5393 ( .A(n4135), .B(n4134), .Z(n4136) );
  NAND U5394 ( .A(n4137), .B(n4136), .Z(n4326) );
  NANDN U5395 ( .A(n4143), .B(n4142), .Z(n4147) );
  NAND U5396 ( .A(n4145), .B(n4144), .Z(n4146) );
  NAND U5397 ( .A(n4147), .B(n4146), .Z(n4265) );
  NANDN U5398 ( .A(n4149), .B(n4148), .Z(n4153) );
  NAND U5399 ( .A(n4151), .B(n4150), .Z(n4152) );
  AND U5400 ( .A(n4153), .B(n4152), .Z(n4266) );
  XNOR U5401 ( .A(n4265), .B(n4266), .Z(n4267) );
  XOR U5402 ( .A(n1052), .B(a[29]), .Z(n4293) );
  NANDN U5403 ( .A(n4293), .B(n36925), .Z(n4156) );
  NAND U5404 ( .A(n36926), .B(n4154), .Z(n4155) );
  NAND U5405 ( .A(n4156), .B(n4155), .Z(n4251) );
  XNOR U5406 ( .A(n1054), .B(a[23]), .Z(n4290) );
  NANDN U5407 ( .A(n37665), .B(n4290), .Z(n4159) );
  NANDN U5408 ( .A(n4157), .B(n37604), .Z(n4158) );
  NAND U5409 ( .A(n4159), .B(n4158), .Z(n4249) );
  XOR U5410 ( .A(n1056), .B(a[17]), .Z(n4287) );
  NANDN U5411 ( .A(n4287), .B(n38101), .Z(n4162) );
  NAND U5412 ( .A(n38102), .B(n4160), .Z(n4161) );
  NAND U5413 ( .A(n4162), .B(n4161), .Z(n4250) );
  XNOR U5414 ( .A(n4249), .B(n4250), .Z(n4252) );
  XOR U5415 ( .A(n4251), .B(n4252), .Z(n4240) );
  XNOR U5416 ( .A(b[11]), .B(a[27]), .Z(n4296) );
  OR U5417 ( .A(n4296), .B(n37311), .Z(n4165) );
  NANDN U5418 ( .A(n4163), .B(n37218), .Z(n4164) );
  NAND U5419 ( .A(n4165), .B(n4164), .Z(n4238) );
  XOR U5420 ( .A(n1053), .B(a[25]), .Z(n4299) );
  NANDN U5421 ( .A(n4299), .B(n37424), .Z(n4168) );
  NANDN U5422 ( .A(n4166), .B(n37425), .Z(n4167) );
  AND U5423 ( .A(n4168), .B(n4167), .Z(n4237) );
  XNOR U5424 ( .A(n4238), .B(n4237), .Z(n4239) );
  XNOR U5425 ( .A(n4240), .B(n4239), .Z(n4256) );
  NANDN U5426 ( .A(n1049), .B(a[37]), .Z(n4169) );
  XNOR U5427 ( .A(b[1]), .B(n4169), .Z(n4171) );
  NANDN U5428 ( .A(b[0]), .B(a[36]), .Z(n4170) );
  AND U5429 ( .A(n4171), .B(n4170), .Z(n4215) );
  NAND U5430 ( .A(n38490), .B(n4172), .Z(n4174) );
  XNOR U5431 ( .A(b[29]), .B(a[9]), .Z(n4306) );
  OR U5432 ( .A(n4306), .B(n1048), .Z(n4173) );
  NAND U5433 ( .A(n4174), .B(n4173), .Z(n4213) );
  NANDN U5434 ( .A(n1059), .B(a[5]), .Z(n4214) );
  XNOR U5435 ( .A(n4213), .B(n4214), .Z(n4216) );
  XNOR U5436 ( .A(n4215), .B(n4216), .Z(n4254) );
  NANDN U5437 ( .A(n4175), .B(n38205), .Z(n4177) );
  XNOR U5438 ( .A(b[23]), .B(a[15]), .Z(n4309) );
  OR U5439 ( .A(n4309), .B(n38268), .Z(n4176) );
  NAND U5440 ( .A(n4177), .B(n4176), .Z(n4278) );
  XNOR U5441 ( .A(b[7]), .B(a[31]), .Z(n4312) );
  NANDN U5442 ( .A(n4312), .B(n36701), .Z(n4180) );
  NANDN U5443 ( .A(n4178), .B(n36702), .Z(n4179) );
  NAND U5444 ( .A(n4180), .B(n4179), .Z(n4275) );
  XOR U5445 ( .A(b[25]), .B(a[13]), .Z(n4315) );
  NAND U5446 ( .A(n4315), .B(n38325), .Z(n4183) );
  NAND U5447 ( .A(n4181), .B(n38326), .Z(n4182) );
  AND U5448 ( .A(n4183), .B(n4182), .Z(n4276) );
  XNOR U5449 ( .A(n4275), .B(n4276), .Z(n4277) );
  XOR U5450 ( .A(n4278), .B(n4277), .Z(n4253) );
  XOR U5451 ( .A(n4256), .B(n4255), .Z(n4268) );
  XOR U5452 ( .A(n4267), .B(n4268), .Z(n4324) );
  XNOR U5453 ( .A(n4325), .B(n4324), .Z(n4327) );
  XNOR U5454 ( .A(n4326), .B(n4327), .Z(n4336) );
  XOR U5455 ( .A(n4337), .B(n4336), .Z(n4339) );
  NANDN U5456 ( .A(n4185), .B(n4184), .Z(n4189) );
  NAND U5457 ( .A(n4187), .B(n4186), .Z(n4188) );
  NAND U5458 ( .A(n4189), .B(n4188), .Z(n4330) );
  NANDN U5459 ( .A(n4191), .B(n4190), .Z(n4195) );
  NAND U5460 ( .A(n4193), .B(n4192), .Z(n4194) );
  NAND U5461 ( .A(n4195), .B(n4194), .Z(n4331) );
  XNOR U5462 ( .A(n4330), .B(n4331), .Z(n4332) );
  XOR U5463 ( .A(n4333), .B(n4332), .Z(n4210) );
  XOR U5464 ( .A(n4209), .B(n4210), .Z(n4201) );
  XOR U5465 ( .A(n4202), .B(n4201), .Z(n4203) );
  XNOR U5466 ( .A(n4204), .B(n4203), .Z(n4342) );
  XNOR U5467 ( .A(n4342), .B(sreg[261]), .Z(n4344) );
  NAND U5468 ( .A(n4196), .B(sreg[260]), .Z(n4200) );
  OR U5469 ( .A(n4198), .B(n4197), .Z(n4199) );
  AND U5470 ( .A(n4200), .B(n4199), .Z(n4343) );
  XOR U5471 ( .A(n4344), .B(n4343), .Z(c[261]) );
  NAND U5472 ( .A(n4202), .B(n4201), .Z(n4206) );
  NAND U5473 ( .A(n4204), .B(n4203), .Z(n4205) );
  NAND U5474 ( .A(n4206), .B(n4205), .Z(n4350) );
  NANDN U5475 ( .A(n4208), .B(n4207), .Z(n4212) );
  NAND U5476 ( .A(n4210), .B(n4209), .Z(n4211) );
  NAND U5477 ( .A(n4212), .B(n4211), .Z(n4348) );
  NANDN U5478 ( .A(n4214), .B(n4213), .Z(n4218) );
  NAND U5479 ( .A(n4216), .B(n4215), .Z(n4217) );
  NAND U5480 ( .A(n4218), .B(n4217), .Z(n4428) );
  XNOR U5481 ( .A(b[19]), .B(a[20]), .Z(n4375) );
  NANDN U5482 ( .A(n4375), .B(n37934), .Z(n4221) );
  NANDN U5483 ( .A(n4219), .B(n37935), .Z(n4220) );
  NAND U5484 ( .A(n4221), .B(n4220), .Z(n4462) );
  XOR U5485 ( .A(b[27]), .B(a[12]), .Z(n4378) );
  NAND U5486 ( .A(n38423), .B(n4378), .Z(n4224) );
  NAND U5487 ( .A(n4222), .B(n38424), .Z(n4223) );
  NAND U5488 ( .A(n4224), .B(n4223), .Z(n4459) );
  XNOR U5489 ( .A(b[5]), .B(a[34]), .Z(n4381) );
  NANDN U5490 ( .A(n4381), .B(n36587), .Z(n4227) );
  NANDN U5491 ( .A(n4225), .B(n36588), .Z(n4226) );
  AND U5492 ( .A(n4227), .B(n4226), .Z(n4460) );
  XNOR U5493 ( .A(n4459), .B(n4460), .Z(n4461) );
  XNOR U5494 ( .A(n4462), .B(n4461), .Z(n4426) );
  NAND U5495 ( .A(n4228), .B(n37762), .Z(n4230) );
  XOR U5496 ( .A(b[17]), .B(a[22]), .Z(n4384) );
  NAND U5497 ( .A(n4384), .B(n37764), .Z(n4229) );
  NAND U5498 ( .A(n4230), .B(n4229), .Z(n4402) );
  XNOR U5499 ( .A(b[31]), .B(a[8]), .Z(n4387) );
  NANDN U5500 ( .A(n4387), .B(n38552), .Z(n4233) );
  NANDN U5501 ( .A(n4231), .B(n38553), .Z(n4232) );
  NAND U5502 ( .A(n4233), .B(n4232), .Z(n4399) );
  OR U5503 ( .A(n4234), .B(n36105), .Z(n4236) );
  XNOR U5504 ( .A(b[3]), .B(a[36]), .Z(n4390) );
  NANDN U5505 ( .A(n4390), .B(n36107), .Z(n4235) );
  AND U5506 ( .A(n4236), .B(n4235), .Z(n4400) );
  XNOR U5507 ( .A(n4399), .B(n4400), .Z(n4401) );
  XOR U5508 ( .A(n4402), .B(n4401), .Z(n4425) );
  XNOR U5509 ( .A(n4426), .B(n4425), .Z(n4427) );
  XNOR U5510 ( .A(n4428), .B(n4427), .Z(n4366) );
  NANDN U5511 ( .A(n4238), .B(n4237), .Z(n4242) );
  NAND U5512 ( .A(n4240), .B(n4239), .Z(n4241) );
  NAND U5513 ( .A(n4242), .B(n4241), .Z(n4417) );
  NANDN U5514 ( .A(n4244), .B(n4243), .Z(n4248) );
  NAND U5515 ( .A(n4246), .B(n4245), .Z(n4247) );
  NAND U5516 ( .A(n4248), .B(n4247), .Z(n4416) );
  XNOR U5517 ( .A(n4416), .B(n4415), .Z(n4418) );
  XOR U5518 ( .A(n4417), .B(n4418), .Z(n4365) );
  XOR U5519 ( .A(n4366), .B(n4365), .Z(n4367) );
  NANDN U5520 ( .A(n4254), .B(n4253), .Z(n4258) );
  NAND U5521 ( .A(n4256), .B(n4255), .Z(n4257) );
  NAND U5522 ( .A(n4258), .B(n4257), .Z(n4368) );
  XNOR U5523 ( .A(n4367), .B(n4368), .Z(n4479) );
  OR U5524 ( .A(n4260), .B(n4259), .Z(n4264) );
  NAND U5525 ( .A(n4262), .B(n4261), .Z(n4263) );
  NAND U5526 ( .A(n4264), .B(n4263), .Z(n4478) );
  NANDN U5527 ( .A(n4266), .B(n4265), .Z(n4270) );
  NAND U5528 ( .A(n4268), .B(n4267), .Z(n4269) );
  NAND U5529 ( .A(n4270), .B(n4269), .Z(n4361) );
  NANDN U5530 ( .A(n4276), .B(n4275), .Z(n4280) );
  NAND U5531 ( .A(n4278), .B(n4277), .Z(n4279) );
  NAND U5532 ( .A(n4280), .B(n4279), .Z(n4419) );
  NANDN U5533 ( .A(n4282), .B(n4281), .Z(n4286) );
  NAND U5534 ( .A(n4284), .B(n4283), .Z(n4285) );
  AND U5535 ( .A(n4286), .B(n4285), .Z(n4420) );
  XNOR U5536 ( .A(n4419), .B(n4420), .Z(n4421) );
  XOR U5537 ( .A(n1056), .B(a[18]), .Z(n4429) );
  NANDN U5538 ( .A(n4429), .B(n38101), .Z(n4289) );
  NANDN U5539 ( .A(n4287), .B(n38102), .Z(n4288) );
  NAND U5540 ( .A(n4289), .B(n4288), .Z(n4411) );
  XNOR U5541 ( .A(b[15]), .B(a[24]), .Z(n4432) );
  OR U5542 ( .A(n4432), .B(n37665), .Z(n4292) );
  NAND U5543 ( .A(n4290), .B(n37604), .Z(n4291) );
  AND U5544 ( .A(n4292), .B(n4291), .Z(n4412) );
  XNOR U5545 ( .A(n4411), .B(n4412), .Z(n4414) );
  XOR U5546 ( .A(n1052), .B(a[30]), .Z(n4435) );
  NANDN U5547 ( .A(n4435), .B(n36925), .Z(n4295) );
  NANDN U5548 ( .A(n4293), .B(n36926), .Z(n4294) );
  NAND U5549 ( .A(n4295), .B(n4294), .Z(n4413) );
  XNOR U5550 ( .A(n4414), .B(n4413), .Z(n4407) );
  XNOR U5551 ( .A(b[11]), .B(a[28]), .Z(n4438) );
  OR U5552 ( .A(n4438), .B(n37311), .Z(n4298) );
  NANDN U5553 ( .A(n4296), .B(n37218), .Z(n4297) );
  NAND U5554 ( .A(n4298), .B(n4297), .Z(n4406) );
  XOR U5555 ( .A(n1053), .B(a[26]), .Z(n4441) );
  NANDN U5556 ( .A(n4441), .B(n37424), .Z(n4301) );
  NANDN U5557 ( .A(n4299), .B(n37425), .Z(n4300) );
  NAND U5558 ( .A(n4301), .B(n4300), .Z(n4405) );
  XNOR U5559 ( .A(n4406), .B(n4405), .Z(n4408) );
  XNOR U5560 ( .A(n4407), .B(n4408), .Z(n4396) );
  NANDN U5561 ( .A(n1049), .B(a[38]), .Z(n4302) );
  XNOR U5562 ( .A(b[1]), .B(n4302), .Z(n4304) );
  IV U5563 ( .A(a[37]), .Z(n8832) );
  NANDN U5564 ( .A(n8832), .B(n1049), .Z(n4303) );
  AND U5565 ( .A(n4304), .B(n4303), .Z(n4372) );
  ANDN U5566 ( .B(b[31]), .A(n4305), .Z(n4369) );
  NANDN U5567 ( .A(n4306), .B(n38490), .Z(n4308) );
  XNOR U5568 ( .A(n1058), .B(a[10]), .Z(n4444) );
  NANDN U5569 ( .A(n1048), .B(n4444), .Z(n4307) );
  NAND U5570 ( .A(n4308), .B(n4307), .Z(n4370) );
  XOR U5571 ( .A(n4369), .B(n4370), .Z(n4371) );
  XNOR U5572 ( .A(n4372), .B(n4371), .Z(n4393) );
  NANDN U5573 ( .A(n4309), .B(n38205), .Z(n4311) );
  XNOR U5574 ( .A(b[23]), .B(a[16]), .Z(n4450) );
  OR U5575 ( .A(n4450), .B(n38268), .Z(n4310) );
  NAND U5576 ( .A(n4311), .B(n4310), .Z(n4468) );
  XOR U5577 ( .A(b[7]), .B(a[32]), .Z(n4453) );
  NAND U5578 ( .A(n4453), .B(n36701), .Z(n4314) );
  NANDN U5579 ( .A(n4312), .B(n36702), .Z(n4313) );
  NAND U5580 ( .A(n4314), .B(n4313), .Z(n4465) );
  XOR U5581 ( .A(b[25]), .B(a[14]), .Z(n4456) );
  NAND U5582 ( .A(n4456), .B(n38325), .Z(n4317) );
  NAND U5583 ( .A(n4315), .B(n38326), .Z(n4316) );
  AND U5584 ( .A(n4317), .B(n4316), .Z(n4466) );
  XNOR U5585 ( .A(n4465), .B(n4466), .Z(n4467) );
  XNOR U5586 ( .A(n4468), .B(n4467), .Z(n4394) );
  XOR U5587 ( .A(n4396), .B(n4395), .Z(n4422) );
  XNOR U5588 ( .A(n4421), .B(n4422), .Z(n4359) );
  XNOR U5589 ( .A(n4360), .B(n4359), .Z(n4362) );
  XNOR U5590 ( .A(n4361), .B(n4362), .Z(n4477) );
  XOR U5591 ( .A(n4478), .B(n4477), .Z(n4480) );
  NANDN U5592 ( .A(n4319), .B(n4318), .Z(n4323) );
  OR U5593 ( .A(n4321), .B(n4320), .Z(n4322) );
  NAND U5594 ( .A(n4323), .B(n4322), .Z(n4471) );
  NAND U5595 ( .A(n4325), .B(n4324), .Z(n4329) );
  NANDN U5596 ( .A(n4327), .B(n4326), .Z(n4328) );
  NAND U5597 ( .A(n4329), .B(n4328), .Z(n4472) );
  XNOR U5598 ( .A(n4471), .B(n4472), .Z(n4473) );
  XOR U5599 ( .A(n4474), .B(n4473), .Z(n4355) );
  NANDN U5600 ( .A(n4331), .B(n4330), .Z(n4335) );
  NAND U5601 ( .A(n4333), .B(n4332), .Z(n4334) );
  NAND U5602 ( .A(n4335), .B(n4334), .Z(n4353) );
  NANDN U5603 ( .A(n4337), .B(n4336), .Z(n4341) );
  OR U5604 ( .A(n4339), .B(n4338), .Z(n4340) );
  NAND U5605 ( .A(n4341), .B(n4340), .Z(n4354) );
  XNOR U5606 ( .A(n4353), .B(n4354), .Z(n4356) );
  XOR U5607 ( .A(n4355), .B(n4356), .Z(n4347) );
  XOR U5608 ( .A(n4348), .B(n4347), .Z(n4349) );
  XNOR U5609 ( .A(n4350), .B(n4349), .Z(n4483) );
  XNOR U5610 ( .A(n4483), .B(sreg[262]), .Z(n4485) );
  NAND U5611 ( .A(n4342), .B(sreg[261]), .Z(n4346) );
  OR U5612 ( .A(n4344), .B(n4343), .Z(n4345) );
  AND U5613 ( .A(n4346), .B(n4345), .Z(n4484) );
  XOR U5614 ( .A(n4485), .B(n4484), .Z(c[262]) );
  NAND U5615 ( .A(n4348), .B(n4347), .Z(n4352) );
  NAND U5616 ( .A(n4350), .B(n4349), .Z(n4351) );
  NAND U5617 ( .A(n4352), .B(n4351), .Z(n4491) );
  NANDN U5618 ( .A(n4354), .B(n4353), .Z(n4358) );
  NAND U5619 ( .A(n4356), .B(n4355), .Z(n4357) );
  NAND U5620 ( .A(n4358), .B(n4357), .Z(n4488) );
  NAND U5621 ( .A(n4360), .B(n4359), .Z(n4364) );
  NANDN U5622 ( .A(n4362), .B(n4361), .Z(n4363) );
  NAND U5623 ( .A(n4364), .B(n4363), .Z(n4616) );
  XNOR U5624 ( .A(n4616), .B(n4617), .Z(n4618) );
  OR U5625 ( .A(n4370), .B(n4369), .Z(n4374) );
  NANDN U5626 ( .A(n4372), .B(n4371), .Z(n4373) );
  NAND U5627 ( .A(n4374), .B(n4373), .Z(n4512) );
  XNOR U5628 ( .A(b[19]), .B(a[21]), .Z(n4564) );
  NANDN U5629 ( .A(n4564), .B(n37934), .Z(n4377) );
  NANDN U5630 ( .A(n4375), .B(n37935), .Z(n4376) );
  NAND U5631 ( .A(n4377), .B(n4376), .Z(n4549) );
  XOR U5632 ( .A(b[27]), .B(a[13]), .Z(n4567) );
  NAND U5633 ( .A(n38423), .B(n4567), .Z(n4380) );
  NAND U5634 ( .A(n4378), .B(n38424), .Z(n4379) );
  NAND U5635 ( .A(n4380), .B(n4379), .Z(n4546) );
  XNOR U5636 ( .A(b[5]), .B(a[35]), .Z(n4570) );
  NANDN U5637 ( .A(n4570), .B(n36587), .Z(n4383) );
  NANDN U5638 ( .A(n4381), .B(n36588), .Z(n4382) );
  AND U5639 ( .A(n4383), .B(n4382), .Z(n4547) );
  XNOR U5640 ( .A(n4546), .B(n4547), .Z(n4548) );
  XNOR U5641 ( .A(n4549), .B(n4548), .Z(n4511) );
  NAND U5642 ( .A(n4384), .B(n37762), .Z(n4386) );
  XOR U5643 ( .A(b[17]), .B(a[23]), .Z(n4573) );
  NAND U5644 ( .A(n4573), .B(n37764), .Z(n4385) );
  NAND U5645 ( .A(n4386), .B(n4385), .Z(n4591) );
  XNOR U5646 ( .A(b[31]), .B(a[9]), .Z(n4576) );
  NANDN U5647 ( .A(n4576), .B(n38552), .Z(n4389) );
  NANDN U5648 ( .A(n4387), .B(n38553), .Z(n4388) );
  NAND U5649 ( .A(n4389), .B(n4388), .Z(n4588) );
  OR U5650 ( .A(n4390), .B(n36105), .Z(n4392) );
  XOR U5651 ( .A(b[3]), .B(n8832), .Z(n4579) );
  NANDN U5652 ( .A(n4579), .B(n36107), .Z(n4391) );
  AND U5653 ( .A(n4392), .B(n4391), .Z(n4589) );
  XNOR U5654 ( .A(n4588), .B(n4589), .Z(n4590) );
  XOR U5655 ( .A(n4591), .B(n4590), .Z(n4510) );
  XOR U5656 ( .A(n4511), .B(n4510), .Z(n4513) );
  XNOR U5657 ( .A(n4512), .B(n4513), .Z(n4610) );
  OR U5658 ( .A(n4394), .B(n4393), .Z(n4398) );
  NANDN U5659 ( .A(n4396), .B(n4395), .Z(n4397) );
  NAND U5660 ( .A(n4398), .B(n4397), .Z(n4611) );
  XNOR U5661 ( .A(n4610), .B(n4611), .Z(n4612) );
  NANDN U5662 ( .A(n4400), .B(n4399), .Z(n4404) );
  NAND U5663 ( .A(n4402), .B(n4401), .Z(n4403) );
  NAND U5664 ( .A(n4404), .B(n4403), .Z(n4503) );
  OR U5665 ( .A(n4406), .B(n4405), .Z(n4410) );
  NANDN U5666 ( .A(n4408), .B(n4407), .Z(n4409) );
  NAND U5667 ( .A(n4410), .B(n4409), .Z(n4501) );
  XNOR U5668 ( .A(n4501), .B(n4500), .Z(n4502) );
  XOR U5669 ( .A(n4503), .B(n4502), .Z(n4613) );
  XOR U5670 ( .A(n4612), .B(n4613), .Z(n4624) );
  NANDN U5671 ( .A(n4420), .B(n4419), .Z(n4424) );
  NANDN U5672 ( .A(n4422), .B(n4421), .Z(n4423) );
  NAND U5673 ( .A(n4424), .B(n4423), .Z(n4607) );
  XOR U5674 ( .A(n1056), .B(a[19]), .Z(n4522) );
  NANDN U5675 ( .A(n4522), .B(n38101), .Z(n4431) );
  NANDN U5676 ( .A(n4429), .B(n38102), .Z(n4430) );
  NAND U5677 ( .A(n4431), .B(n4430), .Z(n4600) );
  XOR U5678 ( .A(b[15]), .B(n7069), .Z(n4519) );
  OR U5679 ( .A(n4519), .B(n37665), .Z(n4434) );
  NANDN U5680 ( .A(n4432), .B(n37604), .Z(n4433) );
  AND U5681 ( .A(n4434), .B(n4433), .Z(n4601) );
  XNOR U5682 ( .A(n4600), .B(n4601), .Z(n4603) );
  XOR U5683 ( .A(n1052), .B(a[31]), .Z(n4516) );
  NANDN U5684 ( .A(n4516), .B(n36925), .Z(n4437) );
  NANDN U5685 ( .A(n4435), .B(n36926), .Z(n4436) );
  NAND U5686 ( .A(n4437), .B(n4436), .Z(n4602) );
  XNOR U5687 ( .A(n4603), .B(n4602), .Z(n4596) );
  XNOR U5688 ( .A(b[11]), .B(a[29]), .Z(n4525) );
  OR U5689 ( .A(n4525), .B(n37311), .Z(n4440) );
  NANDN U5690 ( .A(n4438), .B(n37218), .Z(n4439) );
  NAND U5691 ( .A(n4440), .B(n4439), .Z(n4595) );
  XOR U5692 ( .A(n1053), .B(a[27]), .Z(n4528) );
  NANDN U5693 ( .A(n4528), .B(n37424), .Z(n4443) );
  NANDN U5694 ( .A(n4441), .B(n37425), .Z(n4442) );
  NAND U5695 ( .A(n4443), .B(n4442), .Z(n4594) );
  XNOR U5696 ( .A(n4595), .B(n4594), .Z(n4597) );
  XNOR U5697 ( .A(n4596), .B(n4597), .Z(n4585) );
  NAND U5698 ( .A(n4444), .B(n38490), .Z(n4446) );
  XNOR U5699 ( .A(n1058), .B(a[11]), .Z(n4534) );
  NANDN U5700 ( .A(n1048), .B(n4534), .Z(n4445) );
  NAND U5701 ( .A(n4446), .B(n4445), .Z(n4558) );
  NANDN U5702 ( .A(n1059), .B(a[7]), .Z(n4559) );
  XNOR U5703 ( .A(n4558), .B(n4559), .Z(n4561) );
  NANDN U5704 ( .A(n1049), .B(a[39]), .Z(n4447) );
  XNOR U5705 ( .A(b[1]), .B(n4447), .Z(n4449) );
  NANDN U5706 ( .A(b[0]), .B(a[38]), .Z(n4448) );
  AND U5707 ( .A(n4449), .B(n4448), .Z(n4560) );
  XNOR U5708 ( .A(n4561), .B(n4560), .Z(n4583) );
  NANDN U5709 ( .A(n4450), .B(n38205), .Z(n4452) );
  XNOR U5710 ( .A(b[23]), .B(a[17]), .Z(n4537) );
  OR U5711 ( .A(n4537), .B(n38268), .Z(n4451) );
  NAND U5712 ( .A(n4452), .B(n4451), .Z(n4555) );
  XOR U5713 ( .A(b[7]), .B(a[33]), .Z(n4540) );
  NAND U5714 ( .A(n4540), .B(n36701), .Z(n4455) );
  NAND U5715 ( .A(n4453), .B(n36702), .Z(n4454) );
  NAND U5716 ( .A(n4455), .B(n4454), .Z(n4552) );
  XOR U5717 ( .A(b[25]), .B(a[15]), .Z(n4543) );
  NAND U5718 ( .A(n4543), .B(n38325), .Z(n4458) );
  NAND U5719 ( .A(n4456), .B(n38326), .Z(n4457) );
  AND U5720 ( .A(n4458), .B(n4457), .Z(n4553) );
  XNOR U5721 ( .A(n4552), .B(n4553), .Z(n4554) );
  XOR U5722 ( .A(n4555), .B(n4554), .Z(n4582) );
  XNOR U5723 ( .A(n4585), .B(n4584), .Z(n4507) );
  NANDN U5724 ( .A(n4460), .B(n4459), .Z(n4464) );
  NAND U5725 ( .A(n4462), .B(n4461), .Z(n4463) );
  NAND U5726 ( .A(n4464), .B(n4463), .Z(n4505) );
  NANDN U5727 ( .A(n4466), .B(n4465), .Z(n4470) );
  NAND U5728 ( .A(n4468), .B(n4467), .Z(n4469) );
  AND U5729 ( .A(n4470), .B(n4469), .Z(n4504) );
  XNOR U5730 ( .A(n4505), .B(n4504), .Z(n4506) );
  XNOR U5731 ( .A(n4507), .B(n4506), .Z(n4605) );
  XNOR U5732 ( .A(n4604), .B(n4605), .Z(n4606) );
  XNOR U5733 ( .A(n4607), .B(n4606), .Z(n4622) );
  XNOR U5734 ( .A(n4623), .B(n4622), .Z(n4625) );
  XNOR U5735 ( .A(n4624), .B(n4625), .Z(n4619) );
  XOR U5736 ( .A(n4618), .B(n4619), .Z(n4497) );
  NANDN U5737 ( .A(n4472), .B(n4471), .Z(n4476) );
  NAND U5738 ( .A(n4474), .B(n4473), .Z(n4475) );
  NAND U5739 ( .A(n4476), .B(n4475), .Z(n4494) );
  NANDN U5740 ( .A(n4478), .B(n4477), .Z(n4482) );
  OR U5741 ( .A(n4480), .B(n4479), .Z(n4481) );
  NAND U5742 ( .A(n4482), .B(n4481), .Z(n4495) );
  XNOR U5743 ( .A(n4494), .B(n4495), .Z(n4496) );
  XNOR U5744 ( .A(n4497), .B(n4496), .Z(n4489) );
  XNOR U5745 ( .A(n4488), .B(n4489), .Z(n4490) );
  XNOR U5746 ( .A(n4491), .B(n4490), .Z(n4628) );
  XNOR U5747 ( .A(n4628), .B(sreg[263]), .Z(n4630) );
  NAND U5748 ( .A(n4483), .B(sreg[262]), .Z(n4487) );
  OR U5749 ( .A(n4485), .B(n4484), .Z(n4486) );
  AND U5750 ( .A(n4487), .B(n4486), .Z(n4629) );
  XOR U5751 ( .A(n4630), .B(n4629), .Z(c[263]) );
  NANDN U5752 ( .A(n4489), .B(n4488), .Z(n4493) );
  NAND U5753 ( .A(n4491), .B(n4490), .Z(n4492) );
  NAND U5754 ( .A(n4493), .B(n4492), .Z(n4636) );
  NANDN U5755 ( .A(n4495), .B(n4494), .Z(n4499) );
  NAND U5756 ( .A(n4497), .B(n4496), .Z(n4498) );
  NAND U5757 ( .A(n4499), .B(n4498), .Z(n4634) );
  NANDN U5758 ( .A(n4505), .B(n4504), .Z(n4509) );
  NANDN U5759 ( .A(n4507), .B(n4506), .Z(n4508) );
  NAND U5760 ( .A(n4509), .B(n4508), .Z(n4748) );
  NANDN U5761 ( .A(n4511), .B(n4510), .Z(n4515) );
  OR U5762 ( .A(n4513), .B(n4512), .Z(n4514) );
  NAND U5763 ( .A(n4515), .B(n4514), .Z(n4745) );
  XOR U5764 ( .A(n1052), .B(a[32]), .Z(n4715) );
  NANDN U5765 ( .A(n4715), .B(n36925), .Z(n4518) );
  NANDN U5766 ( .A(n4516), .B(n36926), .Z(n4517) );
  NAND U5767 ( .A(n4518), .B(n4517), .Z(n4681) );
  XOR U5768 ( .A(b[15]), .B(n7202), .Z(n4718) );
  OR U5769 ( .A(n4718), .B(n37665), .Z(n4521) );
  NANDN U5770 ( .A(n4519), .B(n37604), .Z(n4520) );
  NAND U5771 ( .A(n4521), .B(n4520), .Z(n4679) );
  XOR U5772 ( .A(n1056), .B(a[20]), .Z(n4721) );
  NANDN U5773 ( .A(n4721), .B(n38101), .Z(n4524) );
  NANDN U5774 ( .A(n4522), .B(n38102), .Z(n4523) );
  NAND U5775 ( .A(n4524), .B(n4523), .Z(n4680) );
  XNOR U5776 ( .A(n4679), .B(n4680), .Z(n4682) );
  XOR U5777 ( .A(n4681), .B(n4682), .Z(n4670) );
  XOR U5778 ( .A(b[11]), .B(n7434), .Z(n4724) );
  OR U5779 ( .A(n4724), .B(n37311), .Z(n4527) );
  NANDN U5780 ( .A(n4525), .B(n37218), .Z(n4526) );
  NAND U5781 ( .A(n4527), .B(n4526), .Z(n4668) );
  XOR U5782 ( .A(n1053), .B(a[28]), .Z(n4727) );
  NANDN U5783 ( .A(n4727), .B(n37424), .Z(n4530) );
  NANDN U5784 ( .A(n4528), .B(n37425), .Z(n4529) );
  AND U5785 ( .A(n4530), .B(n4529), .Z(n4667) );
  XNOR U5786 ( .A(n4668), .B(n4667), .Z(n4669) );
  XNOR U5787 ( .A(n4670), .B(n4669), .Z(n4686) );
  NANDN U5788 ( .A(n1049), .B(a[40]), .Z(n4531) );
  XNOR U5789 ( .A(b[1]), .B(n4531), .Z(n4533) );
  NANDN U5790 ( .A(b[0]), .B(a[39]), .Z(n4532) );
  AND U5791 ( .A(n4533), .B(n4532), .Z(n4645) );
  NAND U5792 ( .A(n38490), .B(n4534), .Z(n4536) );
  XNOR U5793 ( .A(n1058), .B(a[12]), .Z(n4733) );
  NANDN U5794 ( .A(n1048), .B(n4733), .Z(n4535) );
  NAND U5795 ( .A(n4536), .B(n4535), .Z(n4643) );
  NANDN U5796 ( .A(n1059), .B(a[8]), .Z(n4644) );
  XNOR U5797 ( .A(n4643), .B(n4644), .Z(n4646) );
  XNOR U5798 ( .A(n4645), .B(n4646), .Z(n4684) );
  NANDN U5799 ( .A(n4537), .B(n38205), .Z(n4539) );
  XNOR U5800 ( .A(b[23]), .B(a[18]), .Z(n4736) );
  OR U5801 ( .A(n4736), .B(n38268), .Z(n4538) );
  NAND U5802 ( .A(n4539), .B(n4538), .Z(n4706) );
  XOR U5803 ( .A(b[7]), .B(a[34]), .Z(n4739) );
  NAND U5804 ( .A(n4739), .B(n36701), .Z(n4542) );
  NAND U5805 ( .A(n4540), .B(n36702), .Z(n4541) );
  NAND U5806 ( .A(n4542), .B(n4541), .Z(n4703) );
  XOR U5807 ( .A(b[25]), .B(a[16]), .Z(n4742) );
  NAND U5808 ( .A(n4742), .B(n38325), .Z(n4545) );
  NAND U5809 ( .A(n4543), .B(n38326), .Z(n4544) );
  AND U5810 ( .A(n4545), .B(n4544), .Z(n4704) );
  XNOR U5811 ( .A(n4703), .B(n4704), .Z(n4705) );
  XOR U5812 ( .A(n4706), .B(n4705), .Z(n4683) );
  XOR U5813 ( .A(n4686), .B(n4685), .Z(n4696) );
  NANDN U5814 ( .A(n4547), .B(n4546), .Z(n4551) );
  NAND U5815 ( .A(n4549), .B(n4548), .Z(n4550) );
  NAND U5816 ( .A(n4551), .B(n4550), .Z(n4694) );
  NANDN U5817 ( .A(n4553), .B(n4552), .Z(n4557) );
  NAND U5818 ( .A(n4555), .B(n4554), .Z(n4556) );
  AND U5819 ( .A(n4557), .B(n4556), .Z(n4693) );
  XNOR U5820 ( .A(n4694), .B(n4693), .Z(n4695) );
  XNOR U5821 ( .A(n4696), .B(n4695), .Z(n4746) );
  XNOR U5822 ( .A(n4745), .B(n4746), .Z(n4747) );
  XNOR U5823 ( .A(n4748), .B(n4747), .Z(n4756) );
  XNOR U5824 ( .A(n4755), .B(n4756), .Z(n4758) );
  NANDN U5825 ( .A(n4559), .B(n4558), .Z(n4563) );
  NAND U5826 ( .A(n4561), .B(n4560), .Z(n4562) );
  NAND U5827 ( .A(n4563), .B(n4562), .Z(n4702) );
  XNOR U5828 ( .A(b[19]), .B(a[22]), .Z(n4649) );
  NANDN U5829 ( .A(n4649), .B(n37934), .Z(n4566) );
  NANDN U5830 ( .A(n4564), .B(n37935), .Z(n4565) );
  NAND U5831 ( .A(n4566), .B(n4565), .Z(n4712) );
  XOR U5832 ( .A(b[27]), .B(a[14]), .Z(n4652) );
  NAND U5833 ( .A(n38423), .B(n4652), .Z(n4569) );
  NAND U5834 ( .A(n4567), .B(n38424), .Z(n4568) );
  NAND U5835 ( .A(n4569), .B(n4568), .Z(n4709) );
  XNOR U5836 ( .A(b[5]), .B(a[36]), .Z(n4655) );
  NANDN U5837 ( .A(n4655), .B(n36587), .Z(n4572) );
  NANDN U5838 ( .A(n4570), .B(n36588), .Z(n4571) );
  AND U5839 ( .A(n4572), .B(n4571), .Z(n4710) );
  XNOR U5840 ( .A(n4709), .B(n4710), .Z(n4711) );
  XNOR U5841 ( .A(n4712), .B(n4711), .Z(n4700) );
  NAND U5842 ( .A(n4573), .B(n37762), .Z(n4575) );
  XOR U5843 ( .A(b[17]), .B(a[24]), .Z(n4658) );
  NAND U5844 ( .A(n4658), .B(n37764), .Z(n4574) );
  NAND U5845 ( .A(n4575), .B(n4574), .Z(n4676) );
  XNOR U5846 ( .A(b[31]), .B(a[10]), .Z(n4661) );
  NANDN U5847 ( .A(n4661), .B(n38552), .Z(n4578) );
  NANDN U5848 ( .A(n4576), .B(n38553), .Z(n4577) );
  NAND U5849 ( .A(n4578), .B(n4577), .Z(n4673) );
  OR U5850 ( .A(n4579), .B(n36105), .Z(n4581) );
  XNOR U5851 ( .A(b[3]), .B(a[38]), .Z(n4664) );
  NANDN U5852 ( .A(n4664), .B(n36107), .Z(n4580) );
  AND U5853 ( .A(n4581), .B(n4580), .Z(n4674) );
  XNOR U5854 ( .A(n4673), .B(n4674), .Z(n4675) );
  XOR U5855 ( .A(n4676), .B(n4675), .Z(n4699) );
  XNOR U5856 ( .A(n4700), .B(n4699), .Z(n4701) );
  XNOR U5857 ( .A(n4702), .B(n4701), .Z(n4751) );
  NANDN U5858 ( .A(n4583), .B(n4582), .Z(n4587) );
  NANDN U5859 ( .A(n4585), .B(n4584), .Z(n4586) );
  NAND U5860 ( .A(n4587), .B(n4586), .Z(n4752) );
  XNOR U5861 ( .A(n4751), .B(n4752), .Z(n4753) );
  NANDN U5862 ( .A(n4589), .B(n4588), .Z(n4593) );
  NAND U5863 ( .A(n4591), .B(n4590), .Z(n4592) );
  NAND U5864 ( .A(n4593), .B(n4592), .Z(n4692) );
  OR U5865 ( .A(n4595), .B(n4594), .Z(n4599) );
  NANDN U5866 ( .A(n4597), .B(n4596), .Z(n4598) );
  NAND U5867 ( .A(n4599), .B(n4598), .Z(n4690) );
  XNOR U5868 ( .A(n4690), .B(n4689), .Z(n4691) );
  XOR U5869 ( .A(n4692), .B(n4691), .Z(n4754) );
  XOR U5870 ( .A(n4753), .B(n4754), .Z(n4757) );
  XOR U5871 ( .A(n4758), .B(n4757), .Z(n4762) );
  NANDN U5872 ( .A(n4605), .B(n4604), .Z(n4609) );
  NAND U5873 ( .A(n4607), .B(n4606), .Z(n4608) );
  NAND U5874 ( .A(n4609), .B(n4608), .Z(n4759) );
  NANDN U5875 ( .A(n4611), .B(n4610), .Z(n4615) );
  NAND U5876 ( .A(n4613), .B(n4612), .Z(n4614) );
  NAND U5877 ( .A(n4615), .B(n4614), .Z(n4760) );
  XNOR U5878 ( .A(n4759), .B(n4760), .Z(n4761) );
  XNOR U5879 ( .A(n4762), .B(n4761), .Z(n4640) );
  NANDN U5880 ( .A(n4617), .B(n4616), .Z(n4621) );
  NANDN U5881 ( .A(n4619), .B(n4618), .Z(n4620) );
  NAND U5882 ( .A(n4621), .B(n4620), .Z(n4638) );
  OR U5883 ( .A(n4623), .B(n4622), .Z(n4627) );
  OR U5884 ( .A(n4625), .B(n4624), .Z(n4626) );
  AND U5885 ( .A(n4627), .B(n4626), .Z(n4637) );
  XNOR U5886 ( .A(n4638), .B(n4637), .Z(n4639) );
  XNOR U5887 ( .A(n4640), .B(n4639), .Z(n4633) );
  XOR U5888 ( .A(n4634), .B(n4633), .Z(n4635) );
  XNOR U5889 ( .A(n4636), .B(n4635), .Z(n4765) );
  XNOR U5890 ( .A(n4765), .B(sreg[264]), .Z(n4767) );
  NAND U5891 ( .A(n4628), .B(sreg[263]), .Z(n4632) );
  OR U5892 ( .A(n4630), .B(n4629), .Z(n4631) );
  AND U5893 ( .A(n4632), .B(n4631), .Z(n4766) );
  XOR U5894 ( .A(n4767), .B(n4766), .Z(c[264]) );
  NANDN U5895 ( .A(n4638), .B(n4637), .Z(n4642) );
  NANDN U5896 ( .A(n4640), .B(n4639), .Z(n4641) );
  NAND U5897 ( .A(n4642), .B(n4641), .Z(n4771) );
  NANDN U5898 ( .A(n4644), .B(n4643), .Z(n4648) );
  NAND U5899 ( .A(n4646), .B(n4645), .Z(n4647) );
  NAND U5900 ( .A(n4648), .B(n4647), .Z(n4849) );
  XNOR U5901 ( .A(b[19]), .B(a[23]), .Z(n4796) );
  NANDN U5902 ( .A(n4796), .B(n37934), .Z(n4651) );
  NANDN U5903 ( .A(n4649), .B(n37935), .Z(n4650) );
  NAND U5904 ( .A(n4651), .B(n4650), .Z(n4859) );
  XOR U5905 ( .A(b[27]), .B(a[15]), .Z(n4799) );
  NAND U5906 ( .A(n38423), .B(n4799), .Z(n4654) );
  NAND U5907 ( .A(n4652), .B(n38424), .Z(n4653) );
  NAND U5908 ( .A(n4654), .B(n4653), .Z(n4856) );
  XOR U5909 ( .A(b[5]), .B(n8832), .Z(n4802) );
  NANDN U5910 ( .A(n4802), .B(n36587), .Z(n4657) );
  NANDN U5911 ( .A(n4655), .B(n36588), .Z(n4656) );
  AND U5912 ( .A(n4657), .B(n4656), .Z(n4857) );
  XNOR U5913 ( .A(n4856), .B(n4857), .Z(n4858) );
  XNOR U5914 ( .A(n4859), .B(n4858), .Z(n4847) );
  NAND U5915 ( .A(n4658), .B(n37762), .Z(n4660) );
  XNOR U5916 ( .A(b[17]), .B(a[25]), .Z(n4805) );
  NANDN U5917 ( .A(n4805), .B(n37764), .Z(n4659) );
  NAND U5918 ( .A(n4660), .B(n4659), .Z(n4823) );
  XNOR U5919 ( .A(b[31]), .B(a[11]), .Z(n4808) );
  NANDN U5920 ( .A(n4808), .B(n38552), .Z(n4663) );
  NANDN U5921 ( .A(n4661), .B(n38553), .Z(n4662) );
  NAND U5922 ( .A(n4663), .B(n4662), .Z(n4820) );
  OR U5923 ( .A(n4664), .B(n36105), .Z(n4666) );
  XNOR U5924 ( .A(b[3]), .B(a[39]), .Z(n4811) );
  NANDN U5925 ( .A(n4811), .B(n36107), .Z(n4665) );
  AND U5926 ( .A(n4666), .B(n4665), .Z(n4821) );
  XNOR U5927 ( .A(n4820), .B(n4821), .Z(n4822) );
  XOR U5928 ( .A(n4823), .B(n4822), .Z(n4846) );
  XNOR U5929 ( .A(n4847), .B(n4846), .Z(n4848) );
  XNOR U5930 ( .A(n4849), .B(n4848), .Z(n4787) );
  NANDN U5931 ( .A(n4668), .B(n4667), .Z(n4672) );
  NAND U5932 ( .A(n4670), .B(n4669), .Z(n4671) );
  NAND U5933 ( .A(n4672), .B(n4671), .Z(n4838) );
  NANDN U5934 ( .A(n4674), .B(n4673), .Z(n4678) );
  NAND U5935 ( .A(n4676), .B(n4675), .Z(n4677) );
  NAND U5936 ( .A(n4678), .B(n4677), .Z(n4837) );
  XNOR U5937 ( .A(n4837), .B(n4836), .Z(n4839) );
  XOR U5938 ( .A(n4838), .B(n4839), .Z(n4786) );
  XOR U5939 ( .A(n4787), .B(n4786), .Z(n4788) );
  NANDN U5940 ( .A(n4684), .B(n4683), .Z(n4688) );
  NAND U5941 ( .A(n4686), .B(n4685), .Z(n4687) );
  AND U5942 ( .A(n4688), .B(n4687), .Z(n4789) );
  XNOR U5943 ( .A(n4788), .B(n4789), .Z(n4895) );
  NANDN U5944 ( .A(n4694), .B(n4693), .Z(n4698) );
  NANDN U5945 ( .A(n4696), .B(n4695), .Z(n4697) );
  NAND U5946 ( .A(n4698), .B(n4697), .Z(n4783) );
  NANDN U5947 ( .A(n4704), .B(n4703), .Z(n4708) );
  NAND U5948 ( .A(n4706), .B(n4705), .Z(n4707) );
  NAND U5949 ( .A(n4708), .B(n4707), .Z(n4840) );
  NANDN U5950 ( .A(n4710), .B(n4709), .Z(n4714) );
  NAND U5951 ( .A(n4712), .B(n4711), .Z(n4713) );
  AND U5952 ( .A(n4714), .B(n4713), .Z(n4841) );
  XNOR U5953 ( .A(n4840), .B(n4841), .Z(n4842) );
  XOR U5954 ( .A(n1052), .B(a[33]), .Z(n4868) );
  NANDN U5955 ( .A(n4868), .B(n36925), .Z(n4717) );
  NANDN U5956 ( .A(n4715), .B(n36926), .Z(n4716) );
  NAND U5957 ( .A(n4717), .B(n4716), .Z(n4828) );
  XNOR U5958 ( .A(n1054), .B(a[27]), .Z(n4865) );
  NANDN U5959 ( .A(n37665), .B(n4865), .Z(n4720) );
  NANDN U5960 ( .A(n4718), .B(n37604), .Z(n4719) );
  NAND U5961 ( .A(n4720), .B(n4719), .Z(n4826) );
  XOR U5962 ( .A(n1056), .B(a[21]), .Z(n4862) );
  NANDN U5963 ( .A(n4862), .B(n38101), .Z(n4723) );
  NANDN U5964 ( .A(n4721), .B(n38102), .Z(n4722) );
  NAND U5965 ( .A(n4723), .B(n4722), .Z(n4827) );
  XNOR U5966 ( .A(n4826), .B(n4827), .Z(n4829) );
  XOR U5967 ( .A(n4828), .B(n4829), .Z(n4817) );
  XOR U5968 ( .A(b[11]), .B(n7955), .Z(n4871) );
  OR U5969 ( .A(n4871), .B(n37311), .Z(n4726) );
  NANDN U5970 ( .A(n4724), .B(n37218), .Z(n4725) );
  NAND U5971 ( .A(n4726), .B(n4725), .Z(n4815) );
  XOR U5972 ( .A(n1053), .B(a[29]), .Z(n4874) );
  NANDN U5973 ( .A(n4874), .B(n37424), .Z(n4729) );
  NANDN U5974 ( .A(n4727), .B(n37425), .Z(n4728) );
  AND U5975 ( .A(n4729), .B(n4728), .Z(n4814) );
  XNOR U5976 ( .A(n4815), .B(n4814), .Z(n4816) );
  XNOR U5977 ( .A(n4817), .B(n4816), .Z(n4833) );
  NANDN U5978 ( .A(n1049), .B(a[41]), .Z(n4730) );
  XNOR U5979 ( .A(b[1]), .B(n4730), .Z(n4732) );
  NANDN U5980 ( .A(b[0]), .B(a[40]), .Z(n4731) );
  AND U5981 ( .A(n4732), .B(n4731), .Z(n4792) );
  NAND U5982 ( .A(n38490), .B(n4733), .Z(n4735) );
  XNOR U5983 ( .A(n1058), .B(a[13]), .Z(n4880) );
  NANDN U5984 ( .A(n1048), .B(n4880), .Z(n4734) );
  NAND U5985 ( .A(n4735), .B(n4734), .Z(n4790) );
  NANDN U5986 ( .A(n1059), .B(a[9]), .Z(n4791) );
  XNOR U5987 ( .A(n4790), .B(n4791), .Z(n4793) );
  XNOR U5988 ( .A(n4792), .B(n4793), .Z(n4831) );
  NANDN U5989 ( .A(n4736), .B(n38205), .Z(n4738) );
  XNOR U5990 ( .A(b[23]), .B(a[19]), .Z(n4883) );
  OR U5991 ( .A(n4883), .B(n38268), .Z(n4737) );
  NAND U5992 ( .A(n4738), .B(n4737), .Z(n4853) );
  XOR U5993 ( .A(b[7]), .B(a[35]), .Z(n4886) );
  NAND U5994 ( .A(n4886), .B(n36701), .Z(n4741) );
  NAND U5995 ( .A(n4739), .B(n36702), .Z(n4740) );
  NAND U5996 ( .A(n4741), .B(n4740), .Z(n4850) );
  XOR U5997 ( .A(b[25]), .B(a[17]), .Z(n4889) );
  NAND U5998 ( .A(n4889), .B(n38325), .Z(n4744) );
  NAND U5999 ( .A(n4742), .B(n38326), .Z(n4743) );
  AND U6000 ( .A(n4744), .B(n4743), .Z(n4851) );
  XNOR U6001 ( .A(n4850), .B(n4851), .Z(n4852) );
  XOR U6002 ( .A(n4853), .B(n4852), .Z(n4830) );
  XOR U6003 ( .A(n4833), .B(n4832), .Z(n4843) );
  XOR U6004 ( .A(n4842), .B(n4843), .Z(n4780) );
  XNOR U6005 ( .A(n4781), .B(n4780), .Z(n4782) );
  XOR U6006 ( .A(n4783), .B(n4782), .Z(n4893) );
  XNOR U6007 ( .A(n4892), .B(n4893), .Z(n4894) );
  XNOR U6008 ( .A(n4895), .B(n4894), .Z(n4899) );
  NANDN U6009 ( .A(n4746), .B(n4745), .Z(n4750) );
  NANDN U6010 ( .A(n4748), .B(n4747), .Z(n4749) );
  NAND U6011 ( .A(n4750), .B(n4749), .Z(n4896) );
  XNOR U6012 ( .A(n4896), .B(n4897), .Z(n4898) );
  XNOR U6013 ( .A(n4899), .B(n4898), .Z(n4777) );
  NANDN U6014 ( .A(n4760), .B(n4759), .Z(n4764) );
  NANDN U6015 ( .A(n4762), .B(n4761), .Z(n4763) );
  NAND U6016 ( .A(n4764), .B(n4763), .Z(n4775) );
  XNOR U6017 ( .A(n4774), .B(n4775), .Z(n4776) );
  XNOR U6018 ( .A(n4777), .B(n4776), .Z(n4770) );
  XOR U6019 ( .A(n4771), .B(n4770), .Z(n4772) );
  XNOR U6020 ( .A(n4773), .B(n4772), .Z(n4902) );
  XNOR U6021 ( .A(n4902), .B(sreg[265]), .Z(n4904) );
  NAND U6022 ( .A(n4765), .B(sreg[264]), .Z(n4769) );
  OR U6023 ( .A(n4767), .B(n4766), .Z(n4768) );
  AND U6024 ( .A(n4769), .B(n4768), .Z(n4903) );
  XOR U6025 ( .A(n4904), .B(n4903), .Z(c[265]) );
  NANDN U6026 ( .A(n4775), .B(n4774), .Z(n4779) );
  NANDN U6027 ( .A(n4777), .B(n4776), .Z(n4778) );
  NAND U6028 ( .A(n4779), .B(n4778), .Z(n4907) );
  NAND U6029 ( .A(n4781), .B(n4780), .Z(n4785) );
  OR U6030 ( .A(n4783), .B(n4782), .Z(n4784) );
  NAND U6031 ( .A(n4785), .B(n4784), .Z(n5031) );
  XNOR U6032 ( .A(n5031), .B(n5032), .Z(n5033) );
  NANDN U6033 ( .A(n4791), .B(n4790), .Z(n4795) );
  NAND U6034 ( .A(n4793), .B(n4792), .Z(n4794) );
  NAND U6035 ( .A(n4795), .B(n4794), .Z(n4988) );
  XNOR U6036 ( .A(b[19]), .B(a[24]), .Z(n4935) );
  NANDN U6037 ( .A(n4935), .B(n37934), .Z(n4798) );
  NANDN U6038 ( .A(n4796), .B(n37935), .Z(n4797) );
  NAND U6039 ( .A(n4798), .B(n4797), .Z(n4998) );
  XOR U6040 ( .A(b[27]), .B(a[16]), .Z(n4938) );
  NAND U6041 ( .A(n38423), .B(n4938), .Z(n4801) );
  NAND U6042 ( .A(n4799), .B(n38424), .Z(n4800) );
  NAND U6043 ( .A(n4801), .B(n4800), .Z(n4995) );
  XNOR U6044 ( .A(b[5]), .B(a[38]), .Z(n4941) );
  NANDN U6045 ( .A(n4941), .B(n36587), .Z(n4804) );
  NANDN U6046 ( .A(n4802), .B(n36588), .Z(n4803) );
  AND U6047 ( .A(n4804), .B(n4803), .Z(n4996) );
  XNOR U6048 ( .A(n4995), .B(n4996), .Z(n4997) );
  XNOR U6049 ( .A(n4998), .B(n4997), .Z(n4986) );
  NANDN U6050 ( .A(n4805), .B(n37762), .Z(n4807) );
  XNOR U6051 ( .A(b[17]), .B(a[26]), .Z(n4944) );
  NANDN U6052 ( .A(n4944), .B(n37764), .Z(n4806) );
  NAND U6053 ( .A(n4807), .B(n4806), .Z(n4962) );
  XNOR U6054 ( .A(b[31]), .B(a[12]), .Z(n4947) );
  NANDN U6055 ( .A(n4947), .B(n38552), .Z(n4810) );
  NANDN U6056 ( .A(n4808), .B(n38553), .Z(n4809) );
  NAND U6057 ( .A(n4810), .B(n4809), .Z(n4959) );
  OR U6058 ( .A(n4811), .B(n36105), .Z(n4813) );
  XNOR U6059 ( .A(b[3]), .B(a[40]), .Z(n4950) );
  NANDN U6060 ( .A(n4950), .B(n36107), .Z(n4812) );
  AND U6061 ( .A(n4813), .B(n4812), .Z(n4960) );
  XNOR U6062 ( .A(n4959), .B(n4960), .Z(n4961) );
  XOR U6063 ( .A(n4962), .B(n4961), .Z(n4985) );
  XNOR U6064 ( .A(n4986), .B(n4985), .Z(n4987) );
  XNOR U6065 ( .A(n4988), .B(n4987), .Z(n4926) );
  NANDN U6066 ( .A(n4815), .B(n4814), .Z(n4819) );
  NAND U6067 ( .A(n4817), .B(n4816), .Z(n4818) );
  NAND U6068 ( .A(n4819), .B(n4818), .Z(n4977) );
  NANDN U6069 ( .A(n4821), .B(n4820), .Z(n4825) );
  NAND U6070 ( .A(n4823), .B(n4822), .Z(n4824) );
  NAND U6071 ( .A(n4825), .B(n4824), .Z(n4976) );
  XNOR U6072 ( .A(n4976), .B(n4975), .Z(n4978) );
  XOR U6073 ( .A(n4977), .B(n4978), .Z(n4925) );
  XOR U6074 ( .A(n4926), .B(n4925), .Z(n4927) );
  NANDN U6075 ( .A(n4831), .B(n4830), .Z(n4835) );
  NAND U6076 ( .A(n4833), .B(n4832), .Z(n4834) );
  AND U6077 ( .A(n4835), .B(n4834), .Z(n4928) );
  XOR U6078 ( .A(n4927), .B(n4928), .Z(n5039) );
  NANDN U6079 ( .A(n4841), .B(n4840), .Z(n4845) );
  NAND U6080 ( .A(n4843), .B(n4842), .Z(n4844) );
  NAND U6081 ( .A(n4845), .B(n4844), .Z(n4922) );
  NANDN U6082 ( .A(n4851), .B(n4850), .Z(n4855) );
  NAND U6083 ( .A(n4853), .B(n4852), .Z(n4854) );
  NAND U6084 ( .A(n4855), .B(n4854), .Z(n4979) );
  NANDN U6085 ( .A(n4857), .B(n4856), .Z(n4861) );
  NAND U6086 ( .A(n4859), .B(n4858), .Z(n4860) );
  AND U6087 ( .A(n4861), .B(n4860), .Z(n4980) );
  XNOR U6088 ( .A(n4979), .B(n4980), .Z(n4981) );
  XNOR U6089 ( .A(b[21]), .B(a[22]), .Z(n5007) );
  NANDN U6090 ( .A(n5007), .B(n38101), .Z(n4864) );
  NANDN U6091 ( .A(n4862), .B(n38102), .Z(n4863) );
  NAND U6092 ( .A(n4864), .B(n4863), .Z(n4971) );
  XNOR U6093 ( .A(b[15]), .B(a[28]), .Z(n5004) );
  OR U6094 ( .A(n5004), .B(n37665), .Z(n4867) );
  NAND U6095 ( .A(n4865), .B(n37604), .Z(n4866) );
  AND U6096 ( .A(n4867), .B(n4866), .Z(n4972) );
  XNOR U6097 ( .A(n4971), .B(n4972), .Z(n4974) );
  XNOR U6098 ( .A(b[9]), .B(a[34]), .Z(n5001) );
  NANDN U6099 ( .A(n5001), .B(n36925), .Z(n4870) );
  NANDN U6100 ( .A(n4868), .B(n36926), .Z(n4869) );
  NAND U6101 ( .A(n4870), .B(n4869), .Z(n4973) );
  XNOR U6102 ( .A(n4974), .B(n4973), .Z(n4967) );
  XNOR U6103 ( .A(b[11]), .B(a[32]), .Z(n5010) );
  OR U6104 ( .A(n5010), .B(n37311), .Z(n4873) );
  NANDN U6105 ( .A(n4871), .B(n37218), .Z(n4872) );
  NAND U6106 ( .A(n4873), .B(n4872), .Z(n4966) );
  XOR U6107 ( .A(n1053), .B(a[30]), .Z(n5013) );
  NANDN U6108 ( .A(n5013), .B(n37424), .Z(n4876) );
  NANDN U6109 ( .A(n4874), .B(n37425), .Z(n4875) );
  NAND U6110 ( .A(n4876), .B(n4875), .Z(n4965) );
  XNOR U6111 ( .A(n4966), .B(n4965), .Z(n4968) );
  XNOR U6112 ( .A(n4967), .B(n4968), .Z(n4956) );
  NANDN U6113 ( .A(n1049), .B(a[42]), .Z(n4877) );
  XNOR U6114 ( .A(b[1]), .B(n4877), .Z(n4879) );
  NANDN U6115 ( .A(b[0]), .B(a[41]), .Z(n4878) );
  AND U6116 ( .A(n4879), .B(n4878), .Z(n4931) );
  NAND U6117 ( .A(n38490), .B(n4880), .Z(n4882) );
  XNOR U6118 ( .A(n1058), .B(a[14]), .Z(n5019) );
  NANDN U6119 ( .A(n1048), .B(n5019), .Z(n4881) );
  NAND U6120 ( .A(n4882), .B(n4881), .Z(n4929) );
  NANDN U6121 ( .A(n1059), .B(a[10]), .Z(n4930) );
  XNOR U6122 ( .A(n4929), .B(n4930), .Z(n4932) );
  XNOR U6123 ( .A(n4931), .B(n4932), .Z(n4954) );
  NANDN U6124 ( .A(n4883), .B(n38205), .Z(n4885) );
  XNOR U6125 ( .A(b[23]), .B(a[20]), .Z(n5022) );
  OR U6126 ( .A(n5022), .B(n38268), .Z(n4884) );
  NAND U6127 ( .A(n4885), .B(n4884), .Z(n4992) );
  XOR U6128 ( .A(b[7]), .B(a[36]), .Z(n5025) );
  NAND U6129 ( .A(n5025), .B(n36701), .Z(n4888) );
  NAND U6130 ( .A(n4886), .B(n36702), .Z(n4887) );
  NAND U6131 ( .A(n4888), .B(n4887), .Z(n4989) );
  XOR U6132 ( .A(b[25]), .B(a[18]), .Z(n5028) );
  NAND U6133 ( .A(n5028), .B(n38325), .Z(n4891) );
  NAND U6134 ( .A(n4889), .B(n38326), .Z(n4890) );
  AND U6135 ( .A(n4891), .B(n4890), .Z(n4990) );
  XNOR U6136 ( .A(n4989), .B(n4990), .Z(n4991) );
  XOR U6137 ( .A(n4992), .B(n4991), .Z(n4953) );
  XOR U6138 ( .A(n4956), .B(n4955), .Z(n4982) );
  XNOR U6139 ( .A(n4981), .B(n4982), .Z(n4919) );
  XOR U6140 ( .A(n4920), .B(n4919), .Z(n4921) );
  XNOR U6141 ( .A(n4922), .B(n4921), .Z(n5037) );
  XNOR U6142 ( .A(n5038), .B(n5037), .Z(n5040) );
  XNOR U6143 ( .A(n5039), .B(n5040), .Z(n5034) );
  XOR U6144 ( .A(n5033), .B(n5034), .Z(n4916) );
  NANDN U6145 ( .A(n4897), .B(n4896), .Z(n4901) );
  NANDN U6146 ( .A(n4899), .B(n4898), .Z(n4900) );
  NAND U6147 ( .A(n4901), .B(n4900), .Z(n4914) );
  XNOR U6148 ( .A(n4913), .B(n4914), .Z(n4915) );
  XNOR U6149 ( .A(n4916), .B(n4915), .Z(n4908) );
  XNOR U6150 ( .A(n4907), .B(n4908), .Z(n4909) );
  XNOR U6151 ( .A(n4910), .B(n4909), .Z(n5043) );
  XNOR U6152 ( .A(n5043), .B(sreg[266]), .Z(n5045) );
  NAND U6153 ( .A(n4902), .B(sreg[265]), .Z(n4906) );
  OR U6154 ( .A(n4904), .B(n4903), .Z(n4905) );
  AND U6155 ( .A(n4906), .B(n4905), .Z(n5044) );
  XOR U6156 ( .A(n5045), .B(n5044), .Z(c[266]) );
  NANDN U6157 ( .A(n4908), .B(n4907), .Z(n4912) );
  NAND U6158 ( .A(n4910), .B(n4909), .Z(n4911) );
  NAND U6159 ( .A(n4912), .B(n4911), .Z(n5051) );
  NANDN U6160 ( .A(n4914), .B(n4913), .Z(n4918) );
  NAND U6161 ( .A(n4916), .B(n4915), .Z(n4917) );
  NAND U6162 ( .A(n4918), .B(n4917), .Z(n5048) );
  NAND U6163 ( .A(n4920), .B(n4919), .Z(n4924) );
  NAND U6164 ( .A(n4922), .B(n4921), .Z(n4923) );
  NAND U6165 ( .A(n4924), .B(n4923), .Z(n5176) );
  XNOR U6166 ( .A(n5176), .B(n5177), .Z(n5178) );
  NANDN U6167 ( .A(n4930), .B(n4929), .Z(n4934) );
  NAND U6168 ( .A(n4932), .B(n4931), .Z(n4933) );
  NAND U6169 ( .A(n4934), .B(n4933), .Z(n5121) );
  XOR U6170 ( .A(b[19]), .B(n7069), .Z(n5066) );
  NANDN U6171 ( .A(n5066), .B(n37934), .Z(n4937) );
  NANDN U6172 ( .A(n4935), .B(n37935), .Z(n4936) );
  NAND U6173 ( .A(n4937), .B(n4936), .Z(n5131) );
  XOR U6174 ( .A(b[27]), .B(a[17]), .Z(n5069) );
  NAND U6175 ( .A(n38423), .B(n5069), .Z(n4940) );
  NAND U6176 ( .A(n4938), .B(n38424), .Z(n4939) );
  NAND U6177 ( .A(n4940), .B(n4939), .Z(n5128) );
  XNOR U6178 ( .A(b[5]), .B(a[39]), .Z(n5072) );
  NANDN U6179 ( .A(n5072), .B(n36587), .Z(n4943) );
  NANDN U6180 ( .A(n4941), .B(n36588), .Z(n4942) );
  AND U6181 ( .A(n4943), .B(n4942), .Z(n5129) );
  XNOR U6182 ( .A(n5128), .B(n5129), .Z(n5130) );
  XNOR U6183 ( .A(n5131), .B(n5130), .Z(n5119) );
  NANDN U6184 ( .A(n4944), .B(n37762), .Z(n4946) );
  XOR U6185 ( .A(b[17]), .B(a[27]), .Z(n5075) );
  NAND U6186 ( .A(n5075), .B(n37764), .Z(n4945) );
  NAND U6187 ( .A(n4946), .B(n4945), .Z(n5093) );
  XNOR U6188 ( .A(b[31]), .B(a[13]), .Z(n5078) );
  NANDN U6189 ( .A(n5078), .B(n38552), .Z(n4949) );
  NANDN U6190 ( .A(n4947), .B(n38553), .Z(n4948) );
  NAND U6191 ( .A(n4949), .B(n4948), .Z(n5090) );
  OR U6192 ( .A(n4950), .B(n36105), .Z(n4952) );
  XNOR U6193 ( .A(b[3]), .B(a[41]), .Z(n5081) );
  NANDN U6194 ( .A(n5081), .B(n36107), .Z(n4951) );
  AND U6195 ( .A(n4952), .B(n4951), .Z(n5091) );
  XNOR U6196 ( .A(n5090), .B(n5091), .Z(n5092) );
  XOR U6197 ( .A(n5093), .B(n5092), .Z(n5118) );
  XNOR U6198 ( .A(n5119), .B(n5118), .Z(n5120) );
  XNOR U6199 ( .A(n5121), .B(n5120), .Z(n5170) );
  NANDN U6200 ( .A(n4954), .B(n4953), .Z(n4958) );
  NANDN U6201 ( .A(n4956), .B(n4955), .Z(n4957) );
  NAND U6202 ( .A(n4958), .B(n4957), .Z(n5171) );
  XNOR U6203 ( .A(n5170), .B(n5171), .Z(n5172) );
  NANDN U6204 ( .A(n4960), .B(n4959), .Z(n4964) );
  NAND U6205 ( .A(n4962), .B(n4961), .Z(n4963) );
  NAND U6206 ( .A(n4964), .B(n4963), .Z(n5111) );
  OR U6207 ( .A(n4966), .B(n4965), .Z(n4970) );
  NANDN U6208 ( .A(n4968), .B(n4967), .Z(n4969) );
  NAND U6209 ( .A(n4970), .B(n4969), .Z(n5109) );
  XNOR U6210 ( .A(n5109), .B(n5108), .Z(n5110) );
  XOR U6211 ( .A(n5111), .B(n5110), .Z(n5173) );
  XOR U6212 ( .A(n5172), .B(n5173), .Z(n5184) );
  NANDN U6213 ( .A(n4980), .B(n4979), .Z(n4984) );
  NANDN U6214 ( .A(n4982), .B(n4981), .Z(n4983) );
  NAND U6215 ( .A(n4984), .B(n4983), .Z(n5167) );
  NANDN U6216 ( .A(n4990), .B(n4989), .Z(n4994) );
  NAND U6217 ( .A(n4992), .B(n4991), .Z(n4993) );
  NAND U6218 ( .A(n4994), .B(n4993), .Z(n5112) );
  NANDN U6219 ( .A(n4996), .B(n4995), .Z(n5000) );
  NAND U6220 ( .A(n4998), .B(n4997), .Z(n4999) );
  AND U6221 ( .A(n5000), .B(n4999), .Z(n5113) );
  XNOR U6222 ( .A(n5112), .B(n5113), .Z(n5114) );
  XNOR U6223 ( .A(b[9]), .B(a[35]), .Z(n5134) );
  NANDN U6224 ( .A(n5134), .B(n36925), .Z(n5003) );
  NANDN U6225 ( .A(n5001), .B(n36926), .Z(n5002) );
  NAND U6226 ( .A(n5003), .B(n5002), .Z(n5098) );
  XNOR U6227 ( .A(b[15]), .B(a[29]), .Z(n5137) );
  OR U6228 ( .A(n5137), .B(n37665), .Z(n5006) );
  NANDN U6229 ( .A(n5004), .B(n37604), .Z(n5005) );
  AND U6230 ( .A(n5006), .B(n5005), .Z(n5096) );
  XNOR U6231 ( .A(b[21]), .B(a[23]), .Z(n5140) );
  NANDN U6232 ( .A(n5140), .B(n38101), .Z(n5009) );
  NANDN U6233 ( .A(n5007), .B(n38102), .Z(n5008) );
  AND U6234 ( .A(n5009), .B(n5008), .Z(n5097) );
  XOR U6235 ( .A(n5098), .B(n5099), .Z(n5087) );
  XNOR U6236 ( .A(b[11]), .B(a[33]), .Z(n5143) );
  OR U6237 ( .A(n5143), .B(n37311), .Z(n5012) );
  NANDN U6238 ( .A(n5010), .B(n37218), .Z(n5011) );
  NAND U6239 ( .A(n5012), .B(n5011), .Z(n5085) );
  XOR U6240 ( .A(n1053), .B(a[31]), .Z(n5146) );
  NANDN U6241 ( .A(n5146), .B(n37424), .Z(n5015) );
  NANDN U6242 ( .A(n5013), .B(n37425), .Z(n5014) );
  AND U6243 ( .A(n5015), .B(n5014), .Z(n5084) );
  XNOR U6244 ( .A(n5085), .B(n5084), .Z(n5086) );
  XOR U6245 ( .A(n5087), .B(n5086), .Z(n5104) );
  NANDN U6246 ( .A(n1049), .B(a[43]), .Z(n5016) );
  XNOR U6247 ( .A(b[1]), .B(n5016), .Z(n5018) );
  NANDN U6248 ( .A(b[0]), .B(a[42]), .Z(n5017) );
  AND U6249 ( .A(n5018), .B(n5017), .Z(n5062) );
  NAND U6250 ( .A(n38490), .B(n5019), .Z(n5021) );
  XNOR U6251 ( .A(n1058), .B(a[15]), .Z(n5152) );
  NANDN U6252 ( .A(n1048), .B(n5152), .Z(n5020) );
  NAND U6253 ( .A(n5021), .B(n5020), .Z(n5060) );
  NANDN U6254 ( .A(n1059), .B(a[11]), .Z(n5061) );
  XNOR U6255 ( .A(n5060), .B(n5061), .Z(n5063) );
  XOR U6256 ( .A(n5062), .B(n5063), .Z(n5102) );
  NANDN U6257 ( .A(n5022), .B(n38205), .Z(n5024) );
  XNOR U6258 ( .A(b[23]), .B(a[21]), .Z(n5155) );
  OR U6259 ( .A(n5155), .B(n38268), .Z(n5023) );
  NAND U6260 ( .A(n5024), .B(n5023), .Z(n5125) );
  XNOR U6261 ( .A(b[7]), .B(a[37]), .Z(n5158) );
  NANDN U6262 ( .A(n5158), .B(n36701), .Z(n5027) );
  NAND U6263 ( .A(n5025), .B(n36702), .Z(n5026) );
  NAND U6264 ( .A(n5027), .B(n5026), .Z(n5122) );
  XOR U6265 ( .A(b[25]), .B(a[19]), .Z(n5161) );
  NAND U6266 ( .A(n5161), .B(n38325), .Z(n5030) );
  NAND U6267 ( .A(n5028), .B(n38326), .Z(n5029) );
  AND U6268 ( .A(n5030), .B(n5029), .Z(n5123) );
  XNOR U6269 ( .A(n5122), .B(n5123), .Z(n5124) );
  XNOR U6270 ( .A(n5125), .B(n5124), .Z(n5103) );
  XOR U6271 ( .A(n5102), .B(n5103), .Z(n5105) );
  XNOR U6272 ( .A(n5104), .B(n5105), .Z(n5115) );
  XOR U6273 ( .A(n5114), .B(n5115), .Z(n5165) );
  XNOR U6274 ( .A(n5164), .B(n5165), .Z(n5166) );
  XNOR U6275 ( .A(n5167), .B(n5166), .Z(n5182) );
  XNOR U6276 ( .A(n5183), .B(n5182), .Z(n5185) );
  XNOR U6277 ( .A(n5184), .B(n5185), .Z(n5179) );
  XOR U6278 ( .A(n5178), .B(n5179), .Z(n5057) );
  NANDN U6279 ( .A(n5032), .B(n5031), .Z(n5036) );
  NANDN U6280 ( .A(n5034), .B(n5033), .Z(n5035) );
  NAND U6281 ( .A(n5036), .B(n5035), .Z(n5055) );
  OR U6282 ( .A(n5038), .B(n5037), .Z(n5042) );
  OR U6283 ( .A(n5040), .B(n5039), .Z(n5041) );
  AND U6284 ( .A(n5042), .B(n5041), .Z(n5054) );
  XNOR U6285 ( .A(n5055), .B(n5054), .Z(n5056) );
  XNOR U6286 ( .A(n5057), .B(n5056), .Z(n5049) );
  XNOR U6287 ( .A(n5048), .B(n5049), .Z(n5050) );
  XNOR U6288 ( .A(n5051), .B(n5050), .Z(n5188) );
  XNOR U6289 ( .A(n5188), .B(sreg[267]), .Z(n5190) );
  NAND U6290 ( .A(n5043), .B(sreg[266]), .Z(n5047) );
  OR U6291 ( .A(n5045), .B(n5044), .Z(n5046) );
  AND U6292 ( .A(n5047), .B(n5046), .Z(n5189) );
  XOR U6293 ( .A(n5190), .B(n5189), .Z(c[267]) );
  NANDN U6294 ( .A(n5049), .B(n5048), .Z(n5053) );
  NAND U6295 ( .A(n5051), .B(n5050), .Z(n5052) );
  NAND U6296 ( .A(n5053), .B(n5052), .Z(n5196) );
  NANDN U6297 ( .A(n5055), .B(n5054), .Z(n5059) );
  NAND U6298 ( .A(n5057), .B(n5056), .Z(n5058) );
  NAND U6299 ( .A(n5059), .B(n5058), .Z(n5194) );
  NANDN U6300 ( .A(n5061), .B(n5060), .Z(n5065) );
  NAND U6301 ( .A(n5063), .B(n5062), .Z(n5064) );
  NAND U6302 ( .A(n5065), .B(n5064), .Z(n5276) );
  XOR U6303 ( .A(b[19]), .B(n7202), .Z(n5219) );
  NANDN U6304 ( .A(n5219), .B(n37934), .Z(n5068) );
  NANDN U6305 ( .A(n5066), .B(n37935), .Z(n5067) );
  NAND U6306 ( .A(n5068), .B(n5067), .Z(n5286) );
  XOR U6307 ( .A(b[27]), .B(a[18]), .Z(n5222) );
  NAND U6308 ( .A(n38423), .B(n5222), .Z(n5071) );
  NAND U6309 ( .A(n5069), .B(n38424), .Z(n5070) );
  NAND U6310 ( .A(n5071), .B(n5070), .Z(n5283) );
  XNOR U6311 ( .A(b[5]), .B(a[40]), .Z(n5225) );
  NANDN U6312 ( .A(n5225), .B(n36587), .Z(n5074) );
  NANDN U6313 ( .A(n5072), .B(n36588), .Z(n5073) );
  AND U6314 ( .A(n5074), .B(n5073), .Z(n5284) );
  XNOR U6315 ( .A(n5283), .B(n5284), .Z(n5285) );
  XNOR U6316 ( .A(n5286), .B(n5285), .Z(n5274) );
  NAND U6317 ( .A(n5075), .B(n37762), .Z(n5077) );
  XOR U6318 ( .A(b[17]), .B(a[28]), .Z(n5228) );
  NAND U6319 ( .A(n5228), .B(n37764), .Z(n5076) );
  NAND U6320 ( .A(n5077), .B(n5076), .Z(n5246) );
  XNOR U6321 ( .A(b[31]), .B(a[14]), .Z(n5231) );
  NANDN U6322 ( .A(n5231), .B(n38552), .Z(n5080) );
  NANDN U6323 ( .A(n5078), .B(n38553), .Z(n5079) );
  NAND U6324 ( .A(n5080), .B(n5079), .Z(n5243) );
  OR U6325 ( .A(n5081), .B(n36105), .Z(n5083) );
  XNOR U6326 ( .A(b[3]), .B(a[42]), .Z(n5234) );
  NANDN U6327 ( .A(n5234), .B(n36107), .Z(n5082) );
  AND U6328 ( .A(n5083), .B(n5082), .Z(n5244) );
  XNOR U6329 ( .A(n5243), .B(n5244), .Z(n5245) );
  XOR U6330 ( .A(n5246), .B(n5245), .Z(n5273) );
  XNOR U6331 ( .A(n5274), .B(n5273), .Z(n5275) );
  XNOR U6332 ( .A(n5276), .B(n5275), .Z(n5319) );
  NANDN U6333 ( .A(n5085), .B(n5084), .Z(n5089) );
  NAND U6334 ( .A(n5087), .B(n5086), .Z(n5088) );
  NAND U6335 ( .A(n5089), .B(n5088), .Z(n5264) );
  NANDN U6336 ( .A(n5091), .B(n5090), .Z(n5095) );
  NAND U6337 ( .A(n5093), .B(n5092), .Z(n5094) );
  NAND U6338 ( .A(n5095), .B(n5094), .Z(n5262) );
  OR U6339 ( .A(n5097), .B(n5096), .Z(n5101) );
  NANDN U6340 ( .A(n5099), .B(n5098), .Z(n5100) );
  NAND U6341 ( .A(n5101), .B(n5100), .Z(n5261) );
  XNOR U6342 ( .A(n5264), .B(n5263), .Z(n5320) );
  XNOR U6343 ( .A(n5319), .B(n5320), .Z(n5321) );
  NANDN U6344 ( .A(n5103), .B(n5102), .Z(n5107) );
  OR U6345 ( .A(n5105), .B(n5104), .Z(n5106) );
  AND U6346 ( .A(n5107), .B(n5106), .Z(n5322) );
  XNOR U6347 ( .A(n5321), .B(n5322), .Z(n5206) );
  NANDN U6348 ( .A(n5113), .B(n5112), .Z(n5117) );
  NANDN U6349 ( .A(n5115), .B(n5114), .Z(n5116) );
  NAND U6350 ( .A(n5117), .B(n5116), .Z(n5328) );
  NANDN U6351 ( .A(n5123), .B(n5122), .Z(n5127) );
  NAND U6352 ( .A(n5125), .B(n5124), .Z(n5126) );
  NAND U6353 ( .A(n5127), .B(n5126), .Z(n5267) );
  NANDN U6354 ( .A(n5129), .B(n5128), .Z(n5133) );
  NAND U6355 ( .A(n5131), .B(n5130), .Z(n5132) );
  AND U6356 ( .A(n5133), .B(n5132), .Z(n5268) );
  XNOR U6357 ( .A(n5267), .B(n5268), .Z(n5269) );
  XNOR U6358 ( .A(b[9]), .B(a[36]), .Z(n5289) );
  NANDN U6359 ( .A(n5289), .B(n36925), .Z(n5136) );
  NANDN U6360 ( .A(n5134), .B(n36926), .Z(n5135) );
  NAND U6361 ( .A(n5136), .B(n5135), .Z(n5251) );
  XOR U6362 ( .A(b[15]), .B(n7434), .Z(n5292) );
  OR U6363 ( .A(n5292), .B(n37665), .Z(n5139) );
  NANDN U6364 ( .A(n5137), .B(n37604), .Z(n5138) );
  AND U6365 ( .A(n5139), .B(n5138), .Z(n5249) );
  XNOR U6366 ( .A(b[21]), .B(a[24]), .Z(n5295) );
  NANDN U6367 ( .A(n5295), .B(n38101), .Z(n5142) );
  NANDN U6368 ( .A(n5140), .B(n38102), .Z(n5141) );
  AND U6369 ( .A(n5142), .B(n5141), .Z(n5250) );
  XOR U6370 ( .A(n5251), .B(n5252), .Z(n5240) );
  XNOR U6371 ( .A(b[11]), .B(a[34]), .Z(n5298) );
  OR U6372 ( .A(n5298), .B(n37311), .Z(n5145) );
  NANDN U6373 ( .A(n5143), .B(n37218), .Z(n5144) );
  NAND U6374 ( .A(n5145), .B(n5144), .Z(n5238) );
  XOR U6375 ( .A(n1053), .B(a[32]), .Z(n5301) );
  NANDN U6376 ( .A(n5301), .B(n37424), .Z(n5148) );
  NANDN U6377 ( .A(n5146), .B(n37425), .Z(n5147) );
  AND U6378 ( .A(n5148), .B(n5147), .Z(n5237) );
  XNOR U6379 ( .A(n5238), .B(n5237), .Z(n5239) );
  XOR U6380 ( .A(n5240), .B(n5239), .Z(n5257) );
  NANDN U6381 ( .A(n1049), .B(a[44]), .Z(n5149) );
  XNOR U6382 ( .A(b[1]), .B(n5149), .Z(n5151) );
  NANDN U6383 ( .A(b[0]), .B(a[43]), .Z(n5150) );
  AND U6384 ( .A(n5151), .B(n5150), .Z(n5215) );
  NAND U6385 ( .A(n38490), .B(n5152), .Z(n5154) );
  XNOR U6386 ( .A(n1058), .B(a[16]), .Z(n5307) );
  NANDN U6387 ( .A(n1048), .B(n5307), .Z(n5153) );
  NAND U6388 ( .A(n5154), .B(n5153), .Z(n5213) );
  NANDN U6389 ( .A(n1059), .B(a[12]), .Z(n5214) );
  XNOR U6390 ( .A(n5213), .B(n5214), .Z(n5216) );
  XOR U6391 ( .A(n5215), .B(n5216), .Z(n5255) );
  NANDN U6392 ( .A(n5155), .B(n38205), .Z(n5157) );
  XNOR U6393 ( .A(b[23]), .B(a[22]), .Z(n5310) );
  OR U6394 ( .A(n5310), .B(n38268), .Z(n5156) );
  NAND U6395 ( .A(n5157), .B(n5156), .Z(n5280) );
  XOR U6396 ( .A(b[7]), .B(a[38]), .Z(n5313) );
  NAND U6397 ( .A(n5313), .B(n36701), .Z(n5160) );
  NANDN U6398 ( .A(n5158), .B(n36702), .Z(n5159) );
  NAND U6399 ( .A(n5160), .B(n5159), .Z(n5277) );
  XOR U6400 ( .A(b[25]), .B(a[20]), .Z(n5316) );
  NAND U6401 ( .A(n5316), .B(n38325), .Z(n5163) );
  NAND U6402 ( .A(n5161), .B(n38326), .Z(n5162) );
  AND U6403 ( .A(n5163), .B(n5162), .Z(n5278) );
  XNOR U6404 ( .A(n5277), .B(n5278), .Z(n5279) );
  XNOR U6405 ( .A(n5280), .B(n5279), .Z(n5256) );
  XOR U6406 ( .A(n5255), .B(n5256), .Z(n5258) );
  XNOR U6407 ( .A(n5257), .B(n5258), .Z(n5270) );
  XOR U6408 ( .A(n5269), .B(n5270), .Z(n5326) );
  XNOR U6409 ( .A(n5325), .B(n5326), .Z(n5327) );
  XOR U6410 ( .A(n5328), .B(n5327), .Z(n5204) );
  XNOR U6411 ( .A(n5203), .B(n5204), .Z(n5205) );
  XNOR U6412 ( .A(n5206), .B(n5205), .Z(n5210) );
  NANDN U6413 ( .A(n5165), .B(n5164), .Z(n5169) );
  NAND U6414 ( .A(n5167), .B(n5166), .Z(n5168) );
  NAND U6415 ( .A(n5169), .B(n5168), .Z(n5207) );
  NANDN U6416 ( .A(n5171), .B(n5170), .Z(n5175) );
  NAND U6417 ( .A(n5173), .B(n5172), .Z(n5174) );
  NAND U6418 ( .A(n5175), .B(n5174), .Z(n5208) );
  XNOR U6419 ( .A(n5207), .B(n5208), .Z(n5209) );
  XNOR U6420 ( .A(n5210), .B(n5209), .Z(n5200) );
  NANDN U6421 ( .A(n5177), .B(n5176), .Z(n5181) );
  NANDN U6422 ( .A(n5179), .B(n5178), .Z(n5180) );
  NAND U6423 ( .A(n5181), .B(n5180), .Z(n5198) );
  OR U6424 ( .A(n5183), .B(n5182), .Z(n5187) );
  OR U6425 ( .A(n5185), .B(n5184), .Z(n5186) );
  AND U6426 ( .A(n5187), .B(n5186), .Z(n5197) );
  XNOR U6427 ( .A(n5198), .B(n5197), .Z(n5199) );
  XNOR U6428 ( .A(n5200), .B(n5199), .Z(n5193) );
  XOR U6429 ( .A(n5194), .B(n5193), .Z(n5195) );
  XNOR U6430 ( .A(n5196), .B(n5195), .Z(n5331) );
  XNOR U6431 ( .A(n5331), .B(sreg[268]), .Z(n5333) );
  NAND U6432 ( .A(n5188), .B(sreg[267]), .Z(n5192) );
  OR U6433 ( .A(n5190), .B(n5189), .Z(n5191) );
  AND U6434 ( .A(n5192), .B(n5191), .Z(n5332) );
  XOR U6435 ( .A(n5333), .B(n5332), .Z(c[268]) );
  NANDN U6436 ( .A(n5198), .B(n5197), .Z(n5202) );
  NANDN U6437 ( .A(n5200), .B(n5199), .Z(n5201) );
  NAND U6438 ( .A(n5202), .B(n5201), .Z(n5337) );
  NANDN U6439 ( .A(n5208), .B(n5207), .Z(n5212) );
  NANDN U6440 ( .A(n5210), .B(n5209), .Z(n5211) );
  NAND U6441 ( .A(n5212), .B(n5211), .Z(n5343) );
  XNOR U6442 ( .A(n5342), .B(n5343), .Z(n5344) );
  NANDN U6443 ( .A(n5214), .B(n5213), .Z(n5218) );
  NAND U6444 ( .A(n5216), .B(n5215), .Z(n5217) );
  NAND U6445 ( .A(n5218), .B(n5217), .Z(n5411) );
  XNOR U6446 ( .A(b[19]), .B(a[27]), .Z(n5354) );
  NANDN U6447 ( .A(n5354), .B(n37934), .Z(n5221) );
  NANDN U6448 ( .A(n5219), .B(n37935), .Z(n5220) );
  NAND U6449 ( .A(n5221), .B(n5220), .Z(n5421) );
  XOR U6450 ( .A(b[27]), .B(a[19]), .Z(n5357) );
  NAND U6451 ( .A(n38423), .B(n5357), .Z(n5224) );
  NAND U6452 ( .A(n5222), .B(n38424), .Z(n5223) );
  NAND U6453 ( .A(n5224), .B(n5223), .Z(n5418) );
  XNOR U6454 ( .A(b[5]), .B(a[41]), .Z(n5360) );
  NANDN U6455 ( .A(n5360), .B(n36587), .Z(n5227) );
  NANDN U6456 ( .A(n5225), .B(n36588), .Z(n5226) );
  AND U6457 ( .A(n5227), .B(n5226), .Z(n5419) );
  XNOR U6458 ( .A(n5418), .B(n5419), .Z(n5420) );
  XNOR U6459 ( .A(n5421), .B(n5420), .Z(n5409) );
  NAND U6460 ( .A(n5228), .B(n37762), .Z(n5230) );
  XOR U6461 ( .A(b[17]), .B(a[29]), .Z(n5363) );
  NAND U6462 ( .A(n5363), .B(n37764), .Z(n5229) );
  NAND U6463 ( .A(n5230), .B(n5229), .Z(n5381) );
  XNOR U6464 ( .A(b[31]), .B(a[15]), .Z(n5366) );
  NANDN U6465 ( .A(n5366), .B(n38552), .Z(n5233) );
  NANDN U6466 ( .A(n5231), .B(n38553), .Z(n5232) );
  NAND U6467 ( .A(n5233), .B(n5232), .Z(n5378) );
  OR U6468 ( .A(n5234), .B(n36105), .Z(n5236) );
  XNOR U6469 ( .A(b[3]), .B(a[43]), .Z(n5369) );
  NANDN U6470 ( .A(n5369), .B(n36107), .Z(n5235) );
  AND U6471 ( .A(n5236), .B(n5235), .Z(n5379) );
  XNOR U6472 ( .A(n5378), .B(n5379), .Z(n5380) );
  XOR U6473 ( .A(n5381), .B(n5380), .Z(n5408) );
  XNOR U6474 ( .A(n5409), .B(n5408), .Z(n5410) );
  XNOR U6475 ( .A(n5411), .B(n5410), .Z(n5454) );
  NANDN U6476 ( .A(n5238), .B(n5237), .Z(n5242) );
  NAND U6477 ( .A(n5240), .B(n5239), .Z(n5241) );
  NAND U6478 ( .A(n5242), .B(n5241), .Z(n5399) );
  NANDN U6479 ( .A(n5244), .B(n5243), .Z(n5248) );
  NAND U6480 ( .A(n5246), .B(n5245), .Z(n5247) );
  NAND U6481 ( .A(n5248), .B(n5247), .Z(n5397) );
  OR U6482 ( .A(n5250), .B(n5249), .Z(n5254) );
  NANDN U6483 ( .A(n5252), .B(n5251), .Z(n5253) );
  NAND U6484 ( .A(n5254), .B(n5253), .Z(n5396) );
  XNOR U6485 ( .A(n5399), .B(n5398), .Z(n5455) );
  XOR U6486 ( .A(n5454), .B(n5455), .Z(n5457) );
  NANDN U6487 ( .A(n5256), .B(n5255), .Z(n5260) );
  OR U6488 ( .A(n5258), .B(n5257), .Z(n5259) );
  NAND U6489 ( .A(n5260), .B(n5259), .Z(n5456) );
  XOR U6490 ( .A(n5457), .B(n5456), .Z(n5474) );
  OR U6491 ( .A(n5262), .B(n5261), .Z(n5266) );
  NAND U6492 ( .A(n5264), .B(n5263), .Z(n5265) );
  NAND U6493 ( .A(n5266), .B(n5265), .Z(n5473) );
  NANDN U6494 ( .A(n5268), .B(n5267), .Z(n5272) );
  NANDN U6495 ( .A(n5270), .B(n5269), .Z(n5271) );
  NAND U6496 ( .A(n5272), .B(n5271), .Z(n5462) );
  NANDN U6497 ( .A(n5278), .B(n5277), .Z(n5282) );
  NAND U6498 ( .A(n5280), .B(n5279), .Z(n5281) );
  NAND U6499 ( .A(n5282), .B(n5281), .Z(n5402) );
  NANDN U6500 ( .A(n5284), .B(n5283), .Z(n5288) );
  NAND U6501 ( .A(n5286), .B(n5285), .Z(n5287) );
  AND U6502 ( .A(n5288), .B(n5287), .Z(n5403) );
  XNOR U6503 ( .A(n5402), .B(n5403), .Z(n5404) );
  XOR U6504 ( .A(b[9]), .B(n8832), .Z(n5424) );
  NANDN U6505 ( .A(n5424), .B(n36925), .Z(n5291) );
  NANDN U6506 ( .A(n5289), .B(n36926), .Z(n5290) );
  NAND U6507 ( .A(n5291), .B(n5290), .Z(n5386) );
  XOR U6508 ( .A(b[15]), .B(n7955), .Z(n5427) );
  OR U6509 ( .A(n5427), .B(n37665), .Z(n5294) );
  NANDN U6510 ( .A(n5292), .B(n37604), .Z(n5293) );
  AND U6511 ( .A(n5294), .B(n5293), .Z(n5384) );
  XOR U6512 ( .A(b[21]), .B(n7069), .Z(n5430) );
  NANDN U6513 ( .A(n5430), .B(n38101), .Z(n5297) );
  NANDN U6514 ( .A(n5295), .B(n38102), .Z(n5296) );
  AND U6515 ( .A(n5297), .B(n5296), .Z(n5385) );
  XOR U6516 ( .A(n5386), .B(n5387), .Z(n5375) );
  XNOR U6517 ( .A(b[11]), .B(a[35]), .Z(n5433) );
  OR U6518 ( .A(n5433), .B(n37311), .Z(n5300) );
  NANDN U6519 ( .A(n5298), .B(n37218), .Z(n5299) );
  NAND U6520 ( .A(n5300), .B(n5299), .Z(n5373) );
  XOR U6521 ( .A(n1053), .B(a[33]), .Z(n5436) );
  NANDN U6522 ( .A(n5436), .B(n37424), .Z(n5303) );
  NANDN U6523 ( .A(n5301), .B(n37425), .Z(n5302) );
  AND U6524 ( .A(n5303), .B(n5302), .Z(n5372) );
  XNOR U6525 ( .A(n5373), .B(n5372), .Z(n5374) );
  XOR U6526 ( .A(n5375), .B(n5374), .Z(n5392) );
  NANDN U6527 ( .A(n1049), .B(a[45]), .Z(n5304) );
  XNOR U6528 ( .A(b[1]), .B(n5304), .Z(n5306) );
  IV U6529 ( .A(a[44]), .Z(n9873) );
  NANDN U6530 ( .A(n9873), .B(n1049), .Z(n5305) );
  AND U6531 ( .A(n5306), .B(n5305), .Z(n5350) );
  NAND U6532 ( .A(n38490), .B(n5307), .Z(n5309) );
  XNOR U6533 ( .A(n1058), .B(a[17]), .Z(n5442) );
  NANDN U6534 ( .A(n1048), .B(n5442), .Z(n5308) );
  NAND U6535 ( .A(n5309), .B(n5308), .Z(n5348) );
  NANDN U6536 ( .A(n1059), .B(a[13]), .Z(n5349) );
  XNOR U6537 ( .A(n5348), .B(n5349), .Z(n5351) );
  XOR U6538 ( .A(n5350), .B(n5351), .Z(n5390) );
  NANDN U6539 ( .A(n5310), .B(n38205), .Z(n5312) );
  XNOR U6540 ( .A(b[23]), .B(a[23]), .Z(n5445) );
  OR U6541 ( .A(n5445), .B(n38268), .Z(n5311) );
  NAND U6542 ( .A(n5312), .B(n5311), .Z(n5415) );
  XOR U6543 ( .A(b[7]), .B(a[39]), .Z(n5448) );
  NAND U6544 ( .A(n5448), .B(n36701), .Z(n5315) );
  NAND U6545 ( .A(n5313), .B(n36702), .Z(n5314) );
  NAND U6546 ( .A(n5315), .B(n5314), .Z(n5412) );
  XOR U6547 ( .A(b[25]), .B(a[21]), .Z(n5451) );
  NAND U6548 ( .A(n5451), .B(n38325), .Z(n5318) );
  NAND U6549 ( .A(n5316), .B(n38326), .Z(n5317) );
  AND U6550 ( .A(n5318), .B(n5317), .Z(n5413) );
  XNOR U6551 ( .A(n5412), .B(n5413), .Z(n5414) );
  XNOR U6552 ( .A(n5415), .B(n5414), .Z(n5391) );
  XOR U6553 ( .A(n5390), .B(n5391), .Z(n5393) );
  XNOR U6554 ( .A(n5392), .B(n5393), .Z(n5405) );
  XNOR U6555 ( .A(n5404), .B(n5405), .Z(n5460) );
  XNOR U6556 ( .A(n5461), .B(n5460), .Z(n5463) );
  XNOR U6557 ( .A(n5462), .B(n5463), .Z(n5472) );
  XOR U6558 ( .A(n5473), .B(n5472), .Z(n5475) );
  NANDN U6559 ( .A(n5320), .B(n5319), .Z(n5324) );
  NAND U6560 ( .A(n5322), .B(n5321), .Z(n5323) );
  NAND U6561 ( .A(n5324), .B(n5323), .Z(n5466) );
  NANDN U6562 ( .A(n5326), .B(n5325), .Z(n5330) );
  NAND U6563 ( .A(n5328), .B(n5327), .Z(n5329) );
  NAND U6564 ( .A(n5330), .B(n5329), .Z(n5467) );
  XNOR U6565 ( .A(n5466), .B(n5467), .Z(n5468) );
  XOR U6566 ( .A(n5469), .B(n5468), .Z(n5345) );
  XOR U6567 ( .A(n5344), .B(n5345), .Z(n5336) );
  XOR U6568 ( .A(n5337), .B(n5336), .Z(n5338) );
  XNOR U6569 ( .A(n5339), .B(n5338), .Z(n5478) );
  XNOR U6570 ( .A(n5478), .B(sreg[269]), .Z(n5480) );
  NAND U6571 ( .A(n5331), .B(sreg[268]), .Z(n5335) );
  OR U6572 ( .A(n5333), .B(n5332), .Z(n5334) );
  AND U6573 ( .A(n5335), .B(n5334), .Z(n5479) );
  XOR U6574 ( .A(n5480), .B(n5479), .Z(c[269]) );
  NAND U6575 ( .A(n5337), .B(n5336), .Z(n5341) );
  NAND U6576 ( .A(n5339), .B(n5338), .Z(n5340) );
  NAND U6577 ( .A(n5341), .B(n5340), .Z(n5486) );
  NANDN U6578 ( .A(n5343), .B(n5342), .Z(n5347) );
  NAND U6579 ( .A(n5345), .B(n5344), .Z(n5346) );
  NAND U6580 ( .A(n5347), .B(n5346), .Z(n5484) );
  NANDN U6581 ( .A(n5349), .B(n5348), .Z(n5353) );
  NAND U6582 ( .A(n5351), .B(n5350), .Z(n5352) );
  NAND U6583 ( .A(n5353), .B(n5352), .Z(n5558) );
  XNOR U6584 ( .A(b[19]), .B(a[28]), .Z(n5525) );
  NANDN U6585 ( .A(n5525), .B(n37934), .Z(n5356) );
  NANDN U6586 ( .A(n5354), .B(n37935), .Z(n5355) );
  NAND U6587 ( .A(n5356), .B(n5355), .Z(n5570) );
  XOR U6588 ( .A(b[27]), .B(a[20]), .Z(n5528) );
  NAND U6589 ( .A(n38423), .B(n5528), .Z(n5359) );
  NAND U6590 ( .A(n5357), .B(n38424), .Z(n5358) );
  NAND U6591 ( .A(n5359), .B(n5358), .Z(n5567) );
  XNOR U6592 ( .A(b[5]), .B(a[42]), .Z(n5531) );
  NANDN U6593 ( .A(n5531), .B(n36587), .Z(n5362) );
  NANDN U6594 ( .A(n5360), .B(n36588), .Z(n5361) );
  AND U6595 ( .A(n5362), .B(n5361), .Z(n5568) );
  XNOR U6596 ( .A(n5567), .B(n5568), .Z(n5569) );
  XNOR U6597 ( .A(n5570), .B(n5569), .Z(n5555) );
  NAND U6598 ( .A(n5363), .B(n37762), .Z(n5365) );
  XNOR U6599 ( .A(b[17]), .B(a[30]), .Z(n5534) );
  NANDN U6600 ( .A(n5534), .B(n37764), .Z(n5364) );
  NAND U6601 ( .A(n5365), .B(n5364), .Z(n5509) );
  XNOR U6602 ( .A(b[31]), .B(a[16]), .Z(n5537) );
  NANDN U6603 ( .A(n5537), .B(n38552), .Z(n5368) );
  NANDN U6604 ( .A(n5366), .B(n38553), .Z(n5367) );
  AND U6605 ( .A(n5368), .B(n5367), .Z(n5507) );
  OR U6606 ( .A(n5369), .B(n36105), .Z(n5371) );
  XOR U6607 ( .A(b[3]), .B(n9873), .Z(n5540) );
  NANDN U6608 ( .A(n5540), .B(n36107), .Z(n5370) );
  AND U6609 ( .A(n5371), .B(n5370), .Z(n5508) );
  XOR U6610 ( .A(n5509), .B(n5510), .Z(n5556) );
  XOR U6611 ( .A(n5555), .B(n5556), .Z(n5557) );
  XNOR U6612 ( .A(n5558), .B(n5557), .Z(n5603) );
  NANDN U6613 ( .A(n5373), .B(n5372), .Z(n5377) );
  NAND U6614 ( .A(n5375), .B(n5374), .Z(n5376) );
  NAND U6615 ( .A(n5377), .B(n5376), .Z(n5546) );
  NANDN U6616 ( .A(n5379), .B(n5378), .Z(n5383) );
  NAND U6617 ( .A(n5381), .B(n5380), .Z(n5382) );
  NAND U6618 ( .A(n5383), .B(n5382), .Z(n5544) );
  OR U6619 ( .A(n5385), .B(n5384), .Z(n5389) );
  NANDN U6620 ( .A(n5387), .B(n5386), .Z(n5388) );
  NAND U6621 ( .A(n5389), .B(n5388), .Z(n5543) );
  XNOR U6622 ( .A(n5546), .B(n5545), .Z(n5604) );
  XOR U6623 ( .A(n5603), .B(n5604), .Z(n5606) );
  NANDN U6624 ( .A(n5391), .B(n5390), .Z(n5395) );
  OR U6625 ( .A(n5393), .B(n5392), .Z(n5394) );
  NAND U6626 ( .A(n5395), .B(n5394), .Z(n5605) );
  XOR U6627 ( .A(n5606), .B(n5605), .Z(n5623) );
  OR U6628 ( .A(n5397), .B(n5396), .Z(n5401) );
  NAND U6629 ( .A(n5399), .B(n5398), .Z(n5400) );
  NAND U6630 ( .A(n5401), .B(n5400), .Z(n5622) );
  NANDN U6631 ( .A(n5403), .B(n5402), .Z(n5407) );
  NANDN U6632 ( .A(n5405), .B(n5404), .Z(n5406) );
  NAND U6633 ( .A(n5407), .B(n5406), .Z(n5611) );
  NANDN U6634 ( .A(n5413), .B(n5412), .Z(n5417) );
  NAND U6635 ( .A(n5415), .B(n5414), .Z(n5416) );
  NAND U6636 ( .A(n5417), .B(n5416), .Z(n5549) );
  NANDN U6637 ( .A(n5419), .B(n5418), .Z(n5423) );
  NAND U6638 ( .A(n5421), .B(n5420), .Z(n5422) );
  AND U6639 ( .A(n5423), .B(n5422), .Z(n5550) );
  XNOR U6640 ( .A(n5549), .B(n5550), .Z(n5551) );
  XNOR U6641 ( .A(b[9]), .B(a[38]), .Z(n5573) );
  NANDN U6642 ( .A(n5573), .B(n36925), .Z(n5426) );
  NANDN U6643 ( .A(n5424), .B(n36926), .Z(n5425) );
  NAND U6644 ( .A(n5426), .B(n5425), .Z(n5515) );
  XNOR U6645 ( .A(b[15]), .B(a[32]), .Z(n5576) );
  OR U6646 ( .A(n5576), .B(n37665), .Z(n5429) );
  NANDN U6647 ( .A(n5427), .B(n37604), .Z(n5428) );
  AND U6648 ( .A(n5429), .B(n5428), .Z(n5513) );
  XOR U6649 ( .A(b[21]), .B(n7202), .Z(n5579) );
  NANDN U6650 ( .A(n5579), .B(n38101), .Z(n5432) );
  NANDN U6651 ( .A(n5430), .B(n38102), .Z(n5431) );
  AND U6652 ( .A(n5432), .B(n5431), .Z(n5514) );
  XOR U6653 ( .A(n5515), .B(n5516), .Z(n5504) );
  XNOR U6654 ( .A(b[11]), .B(a[36]), .Z(n5582) );
  OR U6655 ( .A(n5582), .B(n37311), .Z(n5435) );
  NANDN U6656 ( .A(n5433), .B(n37218), .Z(n5434) );
  NAND U6657 ( .A(n5435), .B(n5434), .Z(n5502) );
  XOR U6658 ( .A(n1053), .B(a[34]), .Z(n5585) );
  NANDN U6659 ( .A(n5585), .B(n37424), .Z(n5438) );
  NANDN U6660 ( .A(n5436), .B(n37425), .Z(n5437) );
  NAND U6661 ( .A(n5438), .B(n5437), .Z(n5501) );
  XOR U6662 ( .A(n5504), .B(n5503), .Z(n5498) );
  NANDN U6663 ( .A(n1049), .B(a[46]), .Z(n5439) );
  XNOR U6664 ( .A(b[1]), .B(n5439), .Z(n5441) );
  NANDN U6665 ( .A(b[0]), .B(a[45]), .Z(n5440) );
  AND U6666 ( .A(n5441), .B(n5440), .Z(n5521) );
  NAND U6667 ( .A(n38490), .B(n5442), .Z(n5444) );
  XNOR U6668 ( .A(n1058), .B(a[18]), .Z(n5591) );
  NANDN U6669 ( .A(n1048), .B(n5591), .Z(n5443) );
  NAND U6670 ( .A(n5444), .B(n5443), .Z(n5519) );
  NANDN U6671 ( .A(n1059), .B(a[14]), .Z(n5520) );
  XNOR U6672 ( .A(n5519), .B(n5520), .Z(n5522) );
  XNOR U6673 ( .A(n5521), .B(n5522), .Z(n5496) );
  NANDN U6674 ( .A(n5445), .B(n38205), .Z(n5447) );
  XNOR U6675 ( .A(b[23]), .B(a[24]), .Z(n5594) );
  OR U6676 ( .A(n5594), .B(n38268), .Z(n5446) );
  NAND U6677 ( .A(n5447), .B(n5446), .Z(n5564) );
  XOR U6678 ( .A(b[7]), .B(a[40]), .Z(n5597) );
  NAND U6679 ( .A(n5597), .B(n36701), .Z(n5450) );
  NAND U6680 ( .A(n5448), .B(n36702), .Z(n5449) );
  NAND U6681 ( .A(n5450), .B(n5449), .Z(n5561) );
  XOR U6682 ( .A(b[25]), .B(a[22]), .Z(n5600) );
  NAND U6683 ( .A(n5600), .B(n38325), .Z(n5453) );
  NAND U6684 ( .A(n5451), .B(n38326), .Z(n5452) );
  AND U6685 ( .A(n5453), .B(n5452), .Z(n5562) );
  XNOR U6686 ( .A(n5561), .B(n5562), .Z(n5563) );
  XOR U6687 ( .A(n5564), .B(n5563), .Z(n5495) );
  XOR U6688 ( .A(n5498), .B(n5497), .Z(n5552) );
  XNOR U6689 ( .A(n5551), .B(n5552), .Z(n5609) );
  XNOR U6690 ( .A(n5610), .B(n5609), .Z(n5612) );
  XNOR U6691 ( .A(n5611), .B(n5612), .Z(n5621) );
  XOR U6692 ( .A(n5622), .B(n5621), .Z(n5624) );
  NANDN U6693 ( .A(n5455), .B(n5454), .Z(n5459) );
  OR U6694 ( .A(n5457), .B(n5456), .Z(n5458) );
  NAND U6695 ( .A(n5459), .B(n5458), .Z(n5615) );
  NAND U6696 ( .A(n5461), .B(n5460), .Z(n5465) );
  NANDN U6697 ( .A(n5463), .B(n5462), .Z(n5464) );
  NAND U6698 ( .A(n5465), .B(n5464), .Z(n5616) );
  XNOR U6699 ( .A(n5615), .B(n5616), .Z(n5617) );
  XOR U6700 ( .A(n5618), .B(n5617), .Z(n5491) );
  NANDN U6701 ( .A(n5467), .B(n5466), .Z(n5471) );
  NAND U6702 ( .A(n5469), .B(n5468), .Z(n5470) );
  NAND U6703 ( .A(n5471), .B(n5470), .Z(n5489) );
  NANDN U6704 ( .A(n5473), .B(n5472), .Z(n5477) );
  OR U6705 ( .A(n5475), .B(n5474), .Z(n5476) );
  NAND U6706 ( .A(n5477), .B(n5476), .Z(n5490) );
  XNOR U6707 ( .A(n5489), .B(n5490), .Z(n5492) );
  XOR U6708 ( .A(n5491), .B(n5492), .Z(n5483) );
  XOR U6709 ( .A(n5484), .B(n5483), .Z(n5485) );
  XNOR U6710 ( .A(n5486), .B(n5485), .Z(n5627) );
  XNOR U6711 ( .A(n5627), .B(sreg[270]), .Z(n5629) );
  NAND U6712 ( .A(n5478), .B(sreg[269]), .Z(n5482) );
  OR U6713 ( .A(n5480), .B(n5479), .Z(n5481) );
  AND U6714 ( .A(n5482), .B(n5481), .Z(n5628) );
  XOR U6715 ( .A(n5629), .B(n5628), .Z(c[270]) );
  NAND U6716 ( .A(n5484), .B(n5483), .Z(n5488) );
  NAND U6717 ( .A(n5486), .B(n5485), .Z(n5487) );
  NAND U6718 ( .A(n5488), .B(n5487), .Z(n5635) );
  NANDN U6719 ( .A(n5490), .B(n5489), .Z(n5494) );
  NAND U6720 ( .A(n5492), .B(n5491), .Z(n5493) );
  NAND U6721 ( .A(n5494), .B(n5493), .Z(n5633) );
  NANDN U6722 ( .A(n5496), .B(n5495), .Z(n5500) );
  NANDN U6723 ( .A(n5498), .B(n5497), .Z(n5499) );
  NAND U6724 ( .A(n5500), .B(n5499), .Z(n5753) );
  OR U6725 ( .A(n5502), .B(n5501), .Z(n5506) );
  NAND U6726 ( .A(n5504), .B(n5503), .Z(n5505) );
  NAND U6727 ( .A(n5506), .B(n5505), .Z(n5692) );
  OR U6728 ( .A(n5508), .B(n5507), .Z(n5512) );
  NANDN U6729 ( .A(n5510), .B(n5509), .Z(n5511) );
  NAND U6730 ( .A(n5512), .B(n5511), .Z(n5691) );
  OR U6731 ( .A(n5514), .B(n5513), .Z(n5518) );
  NANDN U6732 ( .A(n5516), .B(n5515), .Z(n5517) );
  NAND U6733 ( .A(n5518), .B(n5517), .Z(n5690) );
  XOR U6734 ( .A(n5692), .B(n5693), .Z(n5750) );
  NANDN U6735 ( .A(n5520), .B(n5519), .Z(n5524) );
  NAND U6736 ( .A(n5522), .B(n5521), .Z(n5523) );
  NAND U6737 ( .A(n5524), .B(n5523), .Z(n5705) );
  XNOR U6738 ( .A(b[19]), .B(a[29]), .Z(n5672) );
  NANDN U6739 ( .A(n5672), .B(n37934), .Z(n5527) );
  NANDN U6740 ( .A(n5525), .B(n37935), .Z(n5526) );
  NAND U6741 ( .A(n5527), .B(n5526), .Z(n5717) );
  XOR U6742 ( .A(b[27]), .B(a[21]), .Z(n5675) );
  NAND U6743 ( .A(n38423), .B(n5675), .Z(n5530) );
  NAND U6744 ( .A(n5528), .B(n38424), .Z(n5529) );
  NAND U6745 ( .A(n5530), .B(n5529), .Z(n5714) );
  XNOR U6746 ( .A(b[5]), .B(a[43]), .Z(n5678) );
  NANDN U6747 ( .A(n5678), .B(n36587), .Z(n5533) );
  NANDN U6748 ( .A(n5531), .B(n36588), .Z(n5532) );
  AND U6749 ( .A(n5533), .B(n5532), .Z(n5715) );
  XNOR U6750 ( .A(n5714), .B(n5715), .Z(n5716) );
  XNOR U6751 ( .A(n5717), .B(n5716), .Z(n5702) );
  NANDN U6752 ( .A(n5534), .B(n37762), .Z(n5536) );
  XNOR U6753 ( .A(b[17]), .B(a[31]), .Z(n5681) );
  NANDN U6754 ( .A(n5681), .B(n37764), .Z(n5535) );
  NAND U6755 ( .A(n5536), .B(n5535), .Z(n5656) );
  XNOR U6756 ( .A(b[31]), .B(a[17]), .Z(n5684) );
  NANDN U6757 ( .A(n5684), .B(n38552), .Z(n5539) );
  NANDN U6758 ( .A(n5537), .B(n38553), .Z(n5538) );
  AND U6759 ( .A(n5539), .B(n5538), .Z(n5654) );
  OR U6760 ( .A(n5540), .B(n36105), .Z(n5542) );
  XNOR U6761 ( .A(b[3]), .B(a[45]), .Z(n5687) );
  NANDN U6762 ( .A(n5687), .B(n36107), .Z(n5541) );
  AND U6763 ( .A(n5542), .B(n5541), .Z(n5655) );
  XOR U6764 ( .A(n5656), .B(n5657), .Z(n5703) );
  XOR U6765 ( .A(n5702), .B(n5703), .Z(n5704) );
  XNOR U6766 ( .A(n5705), .B(n5704), .Z(n5751) );
  XNOR U6767 ( .A(n5750), .B(n5751), .Z(n5752) );
  XNOR U6768 ( .A(n5753), .B(n5752), .Z(n5771) );
  OR U6769 ( .A(n5544), .B(n5543), .Z(n5548) );
  NAND U6770 ( .A(n5546), .B(n5545), .Z(n5547) );
  NAND U6771 ( .A(n5548), .B(n5547), .Z(n5769) );
  NANDN U6772 ( .A(n5550), .B(n5549), .Z(n5554) );
  NANDN U6773 ( .A(n5552), .B(n5551), .Z(n5553) );
  NAND U6774 ( .A(n5554), .B(n5553), .Z(n5758) );
  OR U6775 ( .A(n5556), .B(n5555), .Z(n5560) );
  NAND U6776 ( .A(n5558), .B(n5557), .Z(n5559) );
  NAND U6777 ( .A(n5560), .B(n5559), .Z(n5757) );
  NANDN U6778 ( .A(n5562), .B(n5561), .Z(n5566) );
  NAND U6779 ( .A(n5564), .B(n5563), .Z(n5565) );
  NAND U6780 ( .A(n5566), .B(n5565), .Z(n5696) );
  NANDN U6781 ( .A(n5568), .B(n5567), .Z(n5572) );
  NAND U6782 ( .A(n5570), .B(n5569), .Z(n5571) );
  AND U6783 ( .A(n5572), .B(n5571), .Z(n5697) );
  XNOR U6784 ( .A(n5696), .B(n5697), .Z(n5698) );
  XNOR U6785 ( .A(b[9]), .B(a[39]), .Z(n5720) );
  NANDN U6786 ( .A(n5720), .B(n36925), .Z(n5575) );
  NANDN U6787 ( .A(n5573), .B(n36926), .Z(n5574) );
  NAND U6788 ( .A(n5575), .B(n5574), .Z(n5662) );
  XNOR U6789 ( .A(b[15]), .B(a[33]), .Z(n5723) );
  OR U6790 ( .A(n5723), .B(n37665), .Z(n5578) );
  NANDN U6791 ( .A(n5576), .B(n37604), .Z(n5577) );
  AND U6792 ( .A(n5578), .B(n5577), .Z(n5660) );
  XNOR U6793 ( .A(b[21]), .B(a[27]), .Z(n5726) );
  NANDN U6794 ( .A(n5726), .B(n38101), .Z(n5581) );
  NANDN U6795 ( .A(n5579), .B(n38102), .Z(n5580) );
  AND U6796 ( .A(n5581), .B(n5580), .Z(n5661) );
  XOR U6797 ( .A(n5662), .B(n5663), .Z(n5651) );
  XOR U6798 ( .A(b[11]), .B(n8832), .Z(n5729) );
  OR U6799 ( .A(n5729), .B(n37311), .Z(n5584) );
  NANDN U6800 ( .A(n5582), .B(n37218), .Z(n5583) );
  NAND U6801 ( .A(n5584), .B(n5583), .Z(n5649) );
  XOR U6802 ( .A(n1053), .B(a[35]), .Z(n5732) );
  NANDN U6803 ( .A(n5732), .B(n37424), .Z(n5587) );
  NANDN U6804 ( .A(n5585), .B(n37425), .Z(n5586) );
  NAND U6805 ( .A(n5587), .B(n5586), .Z(n5648) );
  XOR U6806 ( .A(n5651), .B(n5650), .Z(n5645) );
  NANDN U6807 ( .A(n1049), .B(a[47]), .Z(n5588) );
  XNOR U6808 ( .A(b[1]), .B(n5588), .Z(n5590) );
  NANDN U6809 ( .A(b[0]), .B(a[46]), .Z(n5589) );
  AND U6810 ( .A(n5590), .B(n5589), .Z(n5668) );
  NAND U6811 ( .A(n38490), .B(n5591), .Z(n5593) );
  XNOR U6812 ( .A(n1058), .B(a[19]), .Z(n5735) );
  NANDN U6813 ( .A(n1048), .B(n5735), .Z(n5592) );
  NAND U6814 ( .A(n5593), .B(n5592), .Z(n5666) );
  NANDN U6815 ( .A(n1059), .B(a[15]), .Z(n5667) );
  XNOR U6816 ( .A(n5666), .B(n5667), .Z(n5669) );
  XNOR U6817 ( .A(n5668), .B(n5669), .Z(n5643) );
  NANDN U6818 ( .A(n5594), .B(n38205), .Z(n5596) );
  XOR U6819 ( .A(b[23]), .B(n7069), .Z(n5741) );
  OR U6820 ( .A(n5741), .B(n38268), .Z(n5595) );
  NAND U6821 ( .A(n5596), .B(n5595), .Z(n5711) );
  XOR U6822 ( .A(b[7]), .B(a[41]), .Z(n5744) );
  NAND U6823 ( .A(n5744), .B(n36701), .Z(n5599) );
  NAND U6824 ( .A(n5597), .B(n36702), .Z(n5598) );
  NAND U6825 ( .A(n5599), .B(n5598), .Z(n5708) );
  XOR U6826 ( .A(b[25]), .B(a[23]), .Z(n5747) );
  NAND U6827 ( .A(n5747), .B(n38325), .Z(n5602) );
  NAND U6828 ( .A(n5600), .B(n38326), .Z(n5601) );
  AND U6829 ( .A(n5602), .B(n5601), .Z(n5709) );
  XNOR U6830 ( .A(n5708), .B(n5709), .Z(n5710) );
  XOR U6831 ( .A(n5711), .B(n5710), .Z(n5642) );
  XOR U6832 ( .A(n5645), .B(n5644), .Z(n5699) );
  XNOR U6833 ( .A(n5698), .B(n5699), .Z(n5756) );
  XNOR U6834 ( .A(n5757), .B(n5756), .Z(n5759) );
  XNOR U6835 ( .A(n5758), .B(n5759), .Z(n5768) );
  XNOR U6836 ( .A(n5769), .B(n5768), .Z(n5770) );
  XOR U6837 ( .A(n5771), .B(n5770), .Z(n5765) );
  NANDN U6838 ( .A(n5604), .B(n5603), .Z(n5608) );
  OR U6839 ( .A(n5606), .B(n5605), .Z(n5607) );
  NAND U6840 ( .A(n5608), .B(n5607), .Z(n5762) );
  NAND U6841 ( .A(n5610), .B(n5609), .Z(n5614) );
  NANDN U6842 ( .A(n5612), .B(n5611), .Z(n5613) );
  NAND U6843 ( .A(n5614), .B(n5613), .Z(n5763) );
  XNOR U6844 ( .A(n5762), .B(n5763), .Z(n5764) );
  XNOR U6845 ( .A(n5765), .B(n5764), .Z(n5639) );
  NANDN U6846 ( .A(n5616), .B(n5615), .Z(n5620) );
  NAND U6847 ( .A(n5618), .B(n5617), .Z(n5619) );
  NAND U6848 ( .A(n5620), .B(n5619), .Z(n5636) );
  NANDN U6849 ( .A(n5622), .B(n5621), .Z(n5626) );
  OR U6850 ( .A(n5624), .B(n5623), .Z(n5625) );
  NAND U6851 ( .A(n5626), .B(n5625), .Z(n5637) );
  XNOR U6852 ( .A(n5636), .B(n5637), .Z(n5638) );
  XNOR U6853 ( .A(n5639), .B(n5638), .Z(n5632) );
  XOR U6854 ( .A(n5633), .B(n5632), .Z(n5634) );
  XNOR U6855 ( .A(n5635), .B(n5634), .Z(n5774) );
  XNOR U6856 ( .A(n5774), .B(sreg[271]), .Z(n5776) );
  NAND U6857 ( .A(n5627), .B(sreg[270]), .Z(n5631) );
  OR U6858 ( .A(n5629), .B(n5628), .Z(n5630) );
  AND U6859 ( .A(n5631), .B(n5630), .Z(n5775) );
  XOR U6860 ( .A(n5776), .B(n5775), .Z(c[271]) );
  NANDN U6861 ( .A(n5637), .B(n5636), .Z(n5641) );
  NANDN U6862 ( .A(n5639), .B(n5638), .Z(n5640) );
  NAND U6863 ( .A(n5641), .B(n5640), .Z(n5780) );
  NANDN U6864 ( .A(n5643), .B(n5642), .Z(n5647) );
  NANDN U6865 ( .A(n5645), .B(n5644), .Z(n5646) );
  NAND U6866 ( .A(n5647), .B(n5646), .Z(n5900) );
  OR U6867 ( .A(n5649), .B(n5648), .Z(n5653) );
  NAND U6868 ( .A(n5651), .B(n5650), .Z(n5652) );
  NAND U6869 ( .A(n5653), .B(n5652), .Z(n5839) );
  OR U6870 ( .A(n5655), .B(n5654), .Z(n5659) );
  NANDN U6871 ( .A(n5657), .B(n5656), .Z(n5658) );
  NAND U6872 ( .A(n5659), .B(n5658), .Z(n5838) );
  OR U6873 ( .A(n5661), .B(n5660), .Z(n5665) );
  NANDN U6874 ( .A(n5663), .B(n5662), .Z(n5664) );
  NAND U6875 ( .A(n5665), .B(n5664), .Z(n5837) );
  XOR U6876 ( .A(n5839), .B(n5840), .Z(n5897) );
  NANDN U6877 ( .A(n5667), .B(n5666), .Z(n5671) );
  NAND U6878 ( .A(n5669), .B(n5668), .Z(n5670) );
  NAND U6879 ( .A(n5671), .B(n5670), .Z(n5852) );
  XOR U6880 ( .A(b[19]), .B(n7434), .Z(n5819) );
  NANDN U6881 ( .A(n5819), .B(n37934), .Z(n5674) );
  NANDN U6882 ( .A(n5672), .B(n37935), .Z(n5673) );
  NAND U6883 ( .A(n5674), .B(n5673), .Z(n5888) );
  XOR U6884 ( .A(b[27]), .B(a[22]), .Z(n5822) );
  NAND U6885 ( .A(n38423), .B(n5822), .Z(n5677) );
  NAND U6886 ( .A(n5675), .B(n38424), .Z(n5676) );
  NAND U6887 ( .A(n5677), .B(n5676), .Z(n5885) );
  XOR U6888 ( .A(b[5]), .B(n9873), .Z(n5825) );
  NANDN U6889 ( .A(n5825), .B(n36587), .Z(n5680) );
  NANDN U6890 ( .A(n5678), .B(n36588), .Z(n5679) );
  AND U6891 ( .A(n5680), .B(n5679), .Z(n5886) );
  XNOR U6892 ( .A(n5885), .B(n5886), .Z(n5887) );
  XNOR U6893 ( .A(n5888), .B(n5887), .Z(n5849) );
  NANDN U6894 ( .A(n5681), .B(n37762), .Z(n5683) );
  XOR U6895 ( .A(b[17]), .B(a[32]), .Z(n5828) );
  NAND U6896 ( .A(n5828), .B(n37764), .Z(n5682) );
  NAND U6897 ( .A(n5683), .B(n5682), .Z(n5803) );
  XNOR U6898 ( .A(b[31]), .B(a[18]), .Z(n5831) );
  NANDN U6899 ( .A(n5831), .B(n38552), .Z(n5686) );
  NANDN U6900 ( .A(n5684), .B(n38553), .Z(n5685) );
  AND U6901 ( .A(n5686), .B(n5685), .Z(n5801) );
  OR U6902 ( .A(n5687), .B(n36105), .Z(n5689) );
  XNOR U6903 ( .A(b[3]), .B(a[46]), .Z(n5834) );
  NANDN U6904 ( .A(n5834), .B(n36107), .Z(n5688) );
  AND U6905 ( .A(n5689), .B(n5688), .Z(n5802) );
  XOR U6906 ( .A(n5803), .B(n5804), .Z(n5850) );
  XOR U6907 ( .A(n5849), .B(n5850), .Z(n5851) );
  XNOR U6908 ( .A(n5852), .B(n5851), .Z(n5898) );
  XNOR U6909 ( .A(n5897), .B(n5898), .Z(n5899) );
  XNOR U6910 ( .A(n5900), .B(n5899), .Z(n5918) );
  OR U6911 ( .A(n5691), .B(n5690), .Z(n5695) );
  NANDN U6912 ( .A(n5693), .B(n5692), .Z(n5694) );
  NAND U6913 ( .A(n5695), .B(n5694), .Z(n5916) );
  NANDN U6914 ( .A(n5697), .B(n5696), .Z(n5701) );
  NANDN U6915 ( .A(n5699), .B(n5698), .Z(n5700) );
  NAND U6916 ( .A(n5701), .B(n5700), .Z(n5905) );
  OR U6917 ( .A(n5703), .B(n5702), .Z(n5707) );
  NAND U6918 ( .A(n5705), .B(n5704), .Z(n5706) );
  NAND U6919 ( .A(n5707), .B(n5706), .Z(n5904) );
  NANDN U6920 ( .A(n5709), .B(n5708), .Z(n5713) );
  NAND U6921 ( .A(n5711), .B(n5710), .Z(n5712) );
  NAND U6922 ( .A(n5713), .B(n5712), .Z(n5843) );
  NANDN U6923 ( .A(n5715), .B(n5714), .Z(n5719) );
  NAND U6924 ( .A(n5717), .B(n5716), .Z(n5718) );
  AND U6925 ( .A(n5719), .B(n5718), .Z(n5844) );
  XNOR U6926 ( .A(n5843), .B(n5844), .Z(n5845) );
  XNOR U6927 ( .A(n1052), .B(a[40]), .Z(n5855) );
  NAND U6928 ( .A(n36925), .B(n5855), .Z(n5722) );
  NANDN U6929 ( .A(n5720), .B(n36926), .Z(n5721) );
  NAND U6930 ( .A(n5722), .B(n5721), .Z(n5809) );
  XNOR U6931 ( .A(b[15]), .B(a[34]), .Z(n5858) );
  OR U6932 ( .A(n5858), .B(n37665), .Z(n5725) );
  NANDN U6933 ( .A(n5723), .B(n37604), .Z(n5724) );
  AND U6934 ( .A(n5725), .B(n5724), .Z(n5807) );
  XNOR U6935 ( .A(n1056), .B(a[28]), .Z(n5861) );
  NAND U6936 ( .A(n5861), .B(n38101), .Z(n5728) );
  NANDN U6937 ( .A(n5726), .B(n38102), .Z(n5727) );
  AND U6938 ( .A(n5728), .B(n5727), .Z(n5808) );
  XOR U6939 ( .A(n5809), .B(n5810), .Z(n5798) );
  XNOR U6940 ( .A(b[11]), .B(a[38]), .Z(n5864) );
  OR U6941 ( .A(n5864), .B(n37311), .Z(n5731) );
  NANDN U6942 ( .A(n5729), .B(n37218), .Z(n5730) );
  NAND U6943 ( .A(n5731), .B(n5730), .Z(n5796) );
  XOR U6944 ( .A(n1053), .B(a[36]), .Z(n5867) );
  NANDN U6945 ( .A(n5867), .B(n37424), .Z(n5734) );
  NANDN U6946 ( .A(n5732), .B(n37425), .Z(n5733) );
  NAND U6947 ( .A(n5734), .B(n5733), .Z(n5795) );
  XOR U6948 ( .A(n5798), .B(n5797), .Z(n5792) );
  NAND U6949 ( .A(n38490), .B(n5735), .Z(n5737) );
  XNOR U6950 ( .A(n1058), .B(a[20]), .Z(n5873) );
  NANDN U6951 ( .A(n1048), .B(n5873), .Z(n5736) );
  NAND U6952 ( .A(n5737), .B(n5736), .Z(n5813) );
  NANDN U6953 ( .A(n1059), .B(a[16]), .Z(n5814) );
  XNOR U6954 ( .A(n5813), .B(n5814), .Z(n5816) );
  NANDN U6955 ( .A(n1049), .B(a[48]), .Z(n5738) );
  XNOR U6956 ( .A(b[1]), .B(n5738), .Z(n5740) );
  NANDN U6957 ( .A(b[0]), .B(a[47]), .Z(n5739) );
  AND U6958 ( .A(n5740), .B(n5739), .Z(n5815) );
  XNOR U6959 ( .A(n5816), .B(n5815), .Z(n5790) );
  NANDN U6960 ( .A(n5741), .B(n38205), .Z(n5743) );
  XOR U6961 ( .A(b[23]), .B(n7202), .Z(n5876) );
  OR U6962 ( .A(n5876), .B(n38268), .Z(n5742) );
  NAND U6963 ( .A(n5743), .B(n5742), .Z(n5894) );
  XOR U6964 ( .A(b[7]), .B(a[42]), .Z(n5879) );
  NAND U6965 ( .A(n5879), .B(n36701), .Z(n5746) );
  NAND U6966 ( .A(n5744), .B(n36702), .Z(n5745) );
  NAND U6967 ( .A(n5746), .B(n5745), .Z(n5891) );
  XOR U6968 ( .A(b[25]), .B(a[24]), .Z(n5882) );
  NAND U6969 ( .A(n5882), .B(n38325), .Z(n5749) );
  NAND U6970 ( .A(n5747), .B(n38326), .Z(n5748) );
  AND U6971 ( .A(n5749), .B(n5748), .Z(n5892) );
  XNOR U6972 ( .A(n5891), .B(n5892), .Z(n5893) );
  XOR U6973 ( .A(n5894), .B(n5893), .Z(n5789) );
  XOR U6974 ( .A(n5792), .B(n5791), .Z(n5846) );
  XNOR U6975 ( .A(n5845), .B(n5846), .Z(n5903) );
  XNOR U6976 ( .A(n5904), .B(n5903), .Z(n5906) );
  XNOR U6977 ( .A(n5905), .B(n5906), .Z(n5915) );
  XNOR U6978 ( .A(n5916), .B(n5915), .Z(n5917) );
  XOR U6979 ( .A(n5918), .B(n5917), .Z(n5912) );
  NANDN U6980 ( .A(n5751), .B(n5750), .Z(n5755) );
  NAND U6981 ( .A(n5753), .B(n5752), .Z(n5754) );
  NAND U6982 ( .A(n5755), .B(n5754), .Z(n5910) );
  NAND U6983 ( .A(n5757), .B(n5756), .Z(n5761) );
  NANDN U6984 ( .A(n5759), .B(n5758), .Z(n5760) );
  AND U6985 ( .A(n5761), .B(n5760), .Z(n5909) );
  XNOR U6986 ( .A(n5910), .B(n5909), .Z(n5911) );
  XNOR U6987 ( .A(n5912), .B(n5911), .Z(n5786) );
  NANDN U6988 ( .A(n5763), .B(n5762), .Z(n5767) );
  NAND U6989 ( .A(n5765), .B(n5764), .Z(n5766) );
  NAND U6990 ( .A(n5767), .B(n5766), .Z(n5783) );
  NANDN U6991 ( .A(n5769), .B(n5768), .Z(n5773) );
  NANDN U6992 ( .A(n5771), .B(n5770), .Z(n5772) );
  NAND U6993 ( .A(n5773), .B(n5772), .Z(n5784) );
  XNOR U6994 ( .A(n5783), .B(n5784), .Z(n5785) );
  XNOR U6995 ( .A(n5786), .B(n5785), .Z(n5779) );
  XOR U6996 ( .A(n5780), .B(n5779), .Z(n5781) );
  XNOR U6997 ( .A(n5782), .B(n5781), .Z(n5921) );
  XNOR U6998 ( .A(n5921), .B(sreg[272]), .Z(n5923) );
  NAND U6999 ( .A(n5774), .B(sreg[271]), .Z(n5778) );
  OR U7000 ( .A(n5776), .B(n5775), .Z(n5777) );
  AND U7001 ( .A(n5778), .B(n5777), .Z(n5922) );
  XOR U7002 ( .A(n5923), .B(n5922), .Z(c[272]) );
  NANDN U7003 ( .A(n5784), .B(n5783), .Z(n5788) );
  NANDN U7004 ( .A(n5786), .B(n5785), .Z(n5787) );
  NAND U7005 ( .A(n5788), .B(n5787), .Z(n5927) );
  NANDN U7006 ( .A(n5790), .B(n5789), .Z(n5794) );
  NANDN U7007 ( .A(n5792), .B(n5791), .Z(n5793) );
  NAND U7008 ( .A(n5794), .B(n5793), .Z(n6045) );
  OR U7009 ( .A(n5796), .B(n5795), .Z(n5800) );
  NAND U7010 ( .A(n5798), .B(n5797), .Z(n5799) );
  NAND U7011 ( .A(n5800), .B(n5799), .Z(n5984) );
  OR U7012 ( .A(n5802), .B(n5801), .Z(n5806) );
  NANDN U7013 ( .A(n5804), .B(n5803), .Z(n5805) );
  NAND U7014 ( .A(n5806), .B(n5805), .Z(n5983) );
  OR U7015 ( .A(n5808), .B(n5807), .Z(n5812) );
  NANDN U7016 ( .A(n5810), .B(n5809), .Z(n5811) );
  NAND U7017 ( .A(n5812), .B(n5811), .Z(n5982) );
  XOR U7018 ( .A(n5984), .B(n5985), .Z(n6042) );
  NANDN U7019 ( .A(n5814), .B(n5813), .Z(n5818) );
  NAND U7020 ( .A(n5816), .B(n5815), .Z(n5817) );
  NAND U7021 ( .A(n5818), .B(n5817), .Z(n5997) );
  XOR U7022 ( .A(b[19]), .B(n7955), .Z(n5942) );
  NANDN U7023 ( .A(n5942), .B(n37934), .Z(n5821) );
  NANDN U7024 ( .A(n5819), .B(n37935), .Z(n5820) );
  NAND U7025 ( .A(n5821), .B(n5820), .Z(n6009) );
  XOR U7026 ( .A(b[27]), .B(a[23]), .Z(n5945) );
  NAND U7027 ( .A(n38423), .B(n5945), .Z(n5824) );
  NAND U7028 ( .A(n5822), .B(n38424), .Z(n5823) );
  NAND U7029 ( .A(n5824), .B(n5823), .Z(n6006) );
  XNOR U7030 ( .A(b[5]), .B(a[45]), .Z(n5948) );
  NANDN U7031 ( .A(n5948), .B(n36587), .Z(n5827) );
  NANDN U7032 ( .A(n5825), .B(n36588), .Z(n5826) );
  AND U7033 ( .A(n5827), .B(n5826), .Z(n6007) );
  XNOR U7034 ( .A(n6006), .B(n6007), .Z(n6008) );
  XNOR U7035 ( .A(n6009), .B(n6008), .Z(n5995) );
  NAND U7036 ( .A(n5828), .B(n37762), .Z(n5830) );
  XOR U7037 ( .A(b[17]), .B(a[33]), .Z(n5951) );
  NAND U7038 ( .A(n5951), .B(n37764), .Z(n5829) );
  NAND U7039 ( .A(n5830), .B(n5829), .Z(n5969) );
  XNOR U7040 ( .A(b[31]), .B(a[19]), .Z(n5954) );
  NANDN U7041 ( .A(n5954), .B(n38552), .Z(n5833) );
  NANDN U7042 ( .A(n5831), .B(n38553), .Z(n5832) );
  NAND U7043 ( .A(n5833), .B(n5832), .Z(n5966) );
  OR U7044 ( .A(n5834), .B(n36105), .Z(n5836) );
  XNOR U7045 ( .A(b[3]), .B(a[47]), .Z(n5957) );
  NANDN U7046 ( .A(n5957), .B(n36107), .Z(n5835) );
  AND U7047 ( .A(n5836), .B(n5835), .Z(n5967) );
  XNOR U7048 ( .A(n5966), .B(n5967), .Z(n5968) );
  XOR U7049 ( .A(n5969), .B(n5968), .Z(n5994) );
  XNOR U7050 ( .A(n5995), .B(n5994), .Z(n5996) );
  XNOR U7051 ( .A(n5997), .B(n5996), .Z(n6043) );
  XNOR U7052 ( .A(n6042), .B(n6043), .Z(n6044) );
  XNOR U7053 ( .A(n6045), .B(n6044), .Z(n6063) );
  OR U7054 ( .A(n5838), .B(n5837), .Z(n5842) );
  NANDN U7055 ( .A(n5840), .B(n5839), .Z(n5841) );
  NAND U7056 ( .A(n5842), .B(n5841), .Z(n6061) );
  NANDN U7057 ( .A(n5844), .B(n5843), .Z(n5848) );
  NANDN U7058 ( .A(n5846), .B(n5845), .Z(n5847) );
  NAND U7059 ( .A(n5848), .B(n5847), .Z(n6051) );
  OR U7060 ( .A(n5850), .B(n5849), .Z(n5854) );
  NAND U7061 ( .A(n5852), .B(n5851), .Z(n5853) );
  NAND U7062 ( .A(n5854), .B(n5853), .Z(n6048) );
  XNOR U7063 ( .A(b[9]), .B(a[41]), .Z(n6012) );
  NANDN U7064 ( .A(n6012), .B(n36925), .Z(n5857) );
  NAND U7065 ( .A(n36926), .B(n5855), .Z(n5856) );
  NAND U7066 ( .A(n5857), .B(n5856), .Z(n5974) );
  XNOR U7067 ( .A(n1054), .B(a[35]), .Z(n6015) );
  NANDN U7068 ( .A(n37665), .B(n6015), .Z(n5860) );
  NANDN U7069 ( .A(n5858), .B(n37604), .Z(n5859) );
  NAND U7070 ( .A(n5860), .B(n5859), .Z(n5972) );
  XNOR U7071 ( .A(b[21]), .B(a[29]), .Z(n6018) );
  NANDN U7072 ( .A(n6018), .B(n38101), .Z(n5863) );
  NAND U7073 ( .A(n38102), .B(n5861), .Z(n5862) );
  NAND U7074 ( .A(n5863), .B(n5862), .Z(n5973) );
  XNOR U7075 ( .A(n5972), .B(n5973), .Z(n5975) );
  XOR U7076 ( .A(n5974), .B(n5975), .Z(n5963) );
  XNOR U7077 ( .A(b[11]), .B(a[39]), .Z(n6021) );
  OR U7078 ( .A(n6021), .B(n37311), .Z(n5866) );
  NANDN U7079 ( .A(n5864), .B(n37218), .Z(n5865) );
  NAND U7080 ( .A(n5866), .B(n5865), .Z(n5961) );
  XOR U7081 ( .A(n1053), .B(a[37]), .Z(n6024) );
  NANDN U7082 ( .A(n6024), .B(n37424), .Z(n5869) );
  NANDN U7083 ( .A(n5867), .B(n37425), .Z(n5868) );
  AND U7084 ( .A(n5869), .B(n5868), .Z(n5960) );
  XNOR U7085 ( .A(n5961), .B(n5960), .Z(n5962) );
  XNOR U7086 ( .A(n5963), .B(n5962), .Z(n5979) );
  NANDN U7087 ( .A(n1049), .B(a[49]), .Z(n5870) );
  XNOR U7088 ( .A(b[1]), .B(n5870), .Z(n5872) );
  NANDN U7089 ( .A(b[0]), .B(a[48]), .Z(n5871) );
  AND U7090 ( .A(n5872), .B(n5871), .Z(n5938) );
  NAND U7091 ( .A(n38490), .B(n5873), .Z(n5875) );
  XNOR U7092 ( .A(n1058), .B(a[21]), .Z(n6030) );
  NANDN U7093 ( .A(n1048), .B(n6030), .Z(n5874) );
  NAND U7094 ( .A(n5875), .B(n5874), .Z(n5936) );
  NANDN U7095 ( .A(n1059), .B(a[17]), .Z(n5937) );
  XNOR U7096 ( .A(n5936), .B(n5937), .Z(n5939) );
  XNOR U7097 ( .A(n5938), .B(n5939), .Z(n5977) );
  NANDN U7098 ( .A(n5876), .B(n38205), .Z(n5878) );
  XNOR U7099 ( .A(b[23]), .B(a[27]), .Z(n6033) );
  OR U7100 ( .A(n6033), .B(n38268), .Z(n5877) );
  NAND U7101 ( .A(n5878), .B(n5877), .Z(n6003) );
  XOR U7102 ( .A(b[7]), .B(a[43]), .Z(n6036) );
  NAND U7103 ( .A(n6036), .B(n36701), .Z(n5881) );
  NAND U7104 ( .A(n5879), .B(n36702), .Z(n5880) );
  NAND U7105 ( .A(n5881), .B(n5880), .Z(n6000) );
  XNOR U7106 ( .A(b[25]), .B(a[25]), .Z(n6039) );
  NANDN U7107 ( .A(n6039), .B(n38325), .Z(n5884) );
  NAND U7108 ( .A(n5882), .B(n38326), .Z(n5883) );
  AND U7109 ( .A(n5884), .B(n5883), .Z(n6001) );
  XNOR U7110 ( .A(n6000), .B(n6001), .Z(n6002) );
  XOR U7111 ( .A(n6003), .B(n6002), .Z(n5976) );
  XOR U7112 ( .A(n5979), .B(n5978), .Z(n5991) );
  NANDN U7113 ( .A(n5886), .B(n5885), .Z(n5890) );
  NAND U7114 ( .A(n5888), .B(n5887), .Z(n5889) );
  NAND U7115 ( .A(n5890), .B(n5889), .Z(n5989) );
  NANDN U7116 ( .A(n5892), .B(n5891), .Z(n5896) );
  NAND U7117 ( .A(n5894), .B(n5893), .Z(n5895) );
  AND U7118 ( .A(n5896), .B(n5895), .Z(n5988) );
  XNOR U7119 ( .A(n5989), .B(n5988), .Z(n5990) );
  XNOR U7120 ( .A(n5991), .B(n5990), .Z(n6049) );
  XNOR U7121 ( .A(n6048), .B(n6049), .Z(n6050) );
  XOR U7122 ( .A(n6051), .B(n6050), .Z(n6060) );
  XNOR U7123 ( .A(n6061), .B(n6060), .Z(n6062) );
  XOR U7124 ( .A(n6063), .B(n6062), .Z(n6057) );
  NANDN U7125 ( .A(n5898), .B(n5897), .Z(n5902) );
  NAND U7126 ( .A(n5900), .B(n5899), .Z(n5901) );
  NAND U7127 ( .A(n5902), .B(n5901), .Z(n6055) );
  NAND U7128 ( .A(n5904), .B(n5903), .Z(n5908) );
  NANDN U7129 ( .A(n5906), .B(n5905), .Z(n5907) );
  AND U7130 ( .A(n5908), .B(n5907), .Z(n6054) );
  XNOR U7131 ( .A(n6055), .B(n6054), .Z(n6056) );
  XNOR U7132 ( .A(n6057), .B(n6056), .Z(n5933) );
  NANDN U7133 ( .A(n5910), .B(n5909), .Z(n5914) );
  NAND U7134 ( .A(n5912), .B(n5911), .Z(n5913) );
  NAND U7135 ( .A(n5914), .B(n5913), .Z(n5930) );
  NANDN U7136 ( .A(n5916), .B(n5915), .Z(n5920) );
  NANDN U7137 ( .A(n5918), .B(n5917), .Z(n5919) );
  NAND U7138 ( .A(n5920), .B(n5919), .Z(n5931) );
  XNOR U7139 ( .A(n5930), .B(n5931), .Z(n5932) );
  XNOR U7140 ( .A(n5933), .B(n5932), .Z(n5926) );
  XOR U7141 ( .A(n5927), .B(n5926), .Z(n5928) );
  XNOR U7142 ( .A(n5929), .B(n5928), .Z(n6066) );
  XNOR U7143 ( .A(n6066), .B(sreg[273]), .Z(n6068) );
  NAND U7144 ( .A(n5921), .B(sreg[272]), .Z(n5925) );
  OR U7145 ( .A(n5923), .B(n5922), .Z(n5924) );
  AND U7146 ( .A(n5925), .B(n5924), .Z(n6067) );
  XOR U7147 ( .A(n6068), .B(n6067), .Z(c[273]) );
  NANDN U7148 ( .A(n5931), .B(n5930), .Z(n5935) );
  NANDN U7149 ( .A(n5933), .B(n5932), .Z(n5934) );
  NAND U7150 ( .A(n5935), .B(n5934), .Z(n6072) );
  NANDN U7151 ( .A(n5937), .B(n5936), .Z(n5941) );
  NAND U7152 ( .A(n5939), .B(n5938), .Z(n5940) );
  NAND U7153 ( .A(n5941), .B(n5940), .Z(n6154) );
  XNOR U7154 ( .A(b[19]), .B(a[32]), .Z(n6123) );
  NANDN U7155 ( .A(n6123), .B(n37934), .Z(n5944) );
  NANDN U7156 ( .A(n5942), .B(n37935), .Z(n5943) );
  NAND U7157 ( .A(n5944), .B(n5943), .Z(n6166) );
  XOR U7158 ( .A(b[27]), .B(a[24]), .Z(n6126) );
  NAND U7159 ( .A(n38423), .B(n6126), .Z(n5947) );
  NAND U7160 ( .A(n5945), .B(n38424), .Z(n5946) );
  NAND U7161 ( .A(n5947), .B(n5946), .Z(n6163) );
  XNOR U7162 ( .A(b[5]), .B(a[46]), .Z(n6129) );
  NANDN U7163 ( .A(n6129), .B(n36587), .Z(n5950) );
  NANDN U7164 ( .A(n5948), .B(n36588), .Z(n5949) );
  AND U7165 ( .A(n5950), .B(n5949), .Z(n6164) );
  XNOR U7166 ( .A(n6163), .B(n6164), .Z(n6165) );
  XNOR U7167 ( .A(n6166), .B(n6165), .Z(n6151) );
  NAND U7168 ( .A(n5951), .B(n37762), .Z(n5953) );
  XOR U7169 ( .A(b[17]), .B(a[34]), .Z(n6132) );
  NAND U7170 ( .A(n6132), .B(n37764), .Z(n5952) );
  NAND U7171 ( .A(n5953), .B(n5952), .Z(n6107) );
  XNOR U7172 ( .A(b[31]), .B(a[20]), .Z(n6135) );
  NANDN U7173 ( .A(n6135), .B(n38552), .Z(n5956) );
  NANDN U7174 ( .A(n5954), .B(n38553), .Z(n5955) );
  AND U7175 ( .A(n5956), .B(n5955), .Z(n6105) );
  OR U7176 ( .A(n5957), .B(n36105), .Z(n5959) );
  XNOR U7177 ( .A(b[3]), .B(a[48]), .Z(n6138) );
  NANDN U7178 ( .A(n6138), .B(n36107), .Z(n5958) );
  AND U7179 ( .A(n5959), .B(n5958), .Z(n6106) );
  XOR U7180 ( .A(n6107), .B(n6108), .Z(n6152) );
  XOR U7181 ( .A(n6151), .B(n6152), .Z(n6153) );
  XNOR U7182 ( .A(n6154), .B(n6153), .Z(n6090) );
  NANDN U7183 ( .A(n5961), .B(n5960), .Z(n5965) );
  NAND U7184 ( .A(n5963), .B(n5962), .Z(n5964) );
  NAND U7185 ( .A(n5965), .B(n5964), .Z(n6143) );
  NANDN U7186 ( .A(n5967), .B(n5966), .Z(n5971) );
  NAND U7187 ( .A(n5969), .B(n5968), .Z(n5970) );
  NAND U7188 ( .A(n5971), .B(n5970), .Z(n6142) );
  XNOR U7189 ( .A(n6142), .B(n6141), .Z(n6144) );
  XOR U7190 ( .A(n6143), .B(n6144), .Z(n6089) );
  XOR U7191 ( .A(n6090), .B(n6089), .Z(n6091) );
  NANDN U7192 ( .A(n5977), .B(n5976), .Z(n5981) );
  NAND U7193 ( .A(n5979), .B(n5978), .Z(n5980) );
  NAND U7194 ( .A(n5981), .B(n5980), .Z(n6092) );
  XNOR U7195 ( .A(n6091), .B(n6092), .Z(n6207) );
  OR U7196 ( .A(n5983), .B(n5982), .Z(n5987) );
  NANDN U7197 ( .A(n5985), .B(n5984), .Z(n5986) );
  NAND U7198 ( .A(n5987), .B(n5986), .Z(n6206) );
  NANDN U7199 ( .A(n5989), .B(n5988), .Z(n5993) );
  NANDN U7200 ( .A(n5991), .B(n5990), .Z(n5992) );
  NAND U7201 ( .A(n5993), .B(n5992), .Z(n6086) );
  NANDN U7202 ( .A(n5995), .B(n5994), .Z(n5999) );
  NAND U7203 ( .A(n5997), .B(n5996), .Z(n5998) );
  NAND U7204 ( .A(n5999), .B(n5998), .Z(n6084) );
  NANDN U7205 ( .A(n6001), .B(n6000), .Z(n6005) );
  NAND U7206 ( .A(n6003), .B(n6002), .Z(n6004) );
  NAND U7207 ( .A(n6005), .B(n6004), .Z(n6145) );
  NANDN U7208 ( .A(n6007), .B(n6006), .Z(n6011) );
  NAND U7209 ( .A(n6009), .B(n6008), .Z(n6010) );
  AND U7210 ( .A(n6011), .B(n6010), .Z(n6146) );
  XNOR U7211 ( .A(n6145), .B(n6146), .Z(n6147) );
  XNOR U7212 ( .A(n1052), .B(a[42]), .Z(n6169) );
  NAND U7213 ( .A(n36925), .B(n6169), .Z(n6014) );
  NANDN U7214 ( .A(n6012), .B(n36926), .Z(n6013) );
  NAND U7215 ( .A(n6014), .B(n6013), .Z(n6113) );
  XNOR U7216 ( .A(b[15]), .B(a[36]), .Z(n6172) );
  OR U7217 ( .A(n6172), .B(n37665), .Z(n6017) );
  NAND U7218 ( .A(n6015), .B(n37604), .Z(n6016) );
  AND U7219 ( .A(n6017), .B(n6016), .Z(n6111) );
  XOR U7220 ( .A(n1056), .B(n7434), .Z(n6175) );
  NAND U7221 ( .A(n6175), .B(n38101), .Z(n6020) );
  NANDN U7222 ( .A(n6018), .B(n38102), .Z(n6019) );
  AND U7223 ( .A(n6020), .B(n6019), .Z(n6112) );
  XOR U7224 ( .A(n6113), .B(n6114), .Z(n6102) );
  XNOR U7225 ( .A(b[11]), .B(a[40]), .Z(n6178) );
  OR U7226 ( .A(n6178), .B(n37311), .Z(n6023) );
  NANDN U7227 ( .A(n6021), .B(n37218), .Z(n6022) );
  NAND U7228 ( .A(n6023), .B(n6022), .Z(n6100) );
  XOR U7229 ( .A(n1053), .B(a[38]), .Z(n6181) );
  NANDN U7230 ( .A(n6181), .B(n37424), .Z(n6026) );
  NANDN U7231 ( .A(n6024), .B(n37425), .Z(n6025) );
  NAND U7232 ( .A(n6026), .B(n6025), .Z(n6099) );
  XOR U7233 ( .A(n6102), .B(n6101), .Z(n6096) );
  NANDN U7234 ( .A(n1049), .B(a[50]), .Z(n6027) );
  XNOR U7235 ( .A(b[1]), .B(n6027), .Z(n6029) );
  NANDN U7236 ( .A(b[0]), .B(a[49]), .Z(n6028) );
  AND U7237 ( .A(n6029), .B(n6028), .Z(n6119) );
  NAND U7238 ( .A(n38490), .B(n6030), .Z(n6032) );
  XNOR U7239 ( .A(n1058), .B(a[22]), .Z(n6187) );
  NANDN U7240 ( .A(n1048), .B(n6187), .Z(n6031) );
  NAND U7241 ( .A(n6032), .B(n6031), .Z(n6117) );
  NANDN U7242 ( .A(n1059), .B(a[18]), .Z(n6118) );
  XNOR U7243 ( .A(n6117), .B(n6118), .Z(n6120) );
  XNOR U7244 ( .A(n6119), .B(n6120), .Z(n6094) );
  NANDN U7245 ( .A(n6033), .B(n38205), .Z(n6035) );
  XNOR U7246 ( .A(b[23]), .B(a[28]), .Z(n6190) );
  OR U7247 ( .A(n6190), .B(n38268), .Z(n6034) );
  NAND U7248 ( .A(n6035), .B(n6034), .Z(n6160) );
  XNOR U7249 ( .A(b[7]), .B(a[44]), .Z(n6193) );
  NANDN U7250 ( .A(n6193), .B(n36701), .Z(n6038) );
  NAND U7251 ( .A(n6036), .B(n36702), .Z(n6037) );
  NAND U7252 ( .A(n6038), .B(n6037), .Z(n6157) );
  XNOR U7253 ( .A(b[25]), .B(a[26]), .Z(n6196) );
  NANDN U7254 ( .A(n6196), .B(n38325), .Z(n6041) );
  NANDN U7255 ( .A(n6039), .B(n38326), .Z(n6040) );
  AND U7256 ( .A(n6041), .B(n6040), .Z(n6158) );
  XNOR U7257 ( .A(n6157), .B(n6158), .Z(n6159) );
  XOR U7258 ( .A(n6160), .B(n6159), .Z(n6093) );
  XOR U7259 ( .A(n6096), .B(n6095), .Z(n6148) );
  XNOR U7260 ( .A(n6147), .B(n6148), .Z(n6083) );
  XOR U7261 ( .A(n6084), .B(n6083), .Z(n6085) );
  XNOR U7262 ( .A(n6086), .B(n6085), .Z(n6205) );
  XOR U7263 ( .A(n6206), .B(n6205), .Z(n6208) );
  NANDN U7264 ( .A(n6043), .B(n6042), .Z(n6047) );
  NAND U7265 ( .A(n6045), .B(n6044), .Z(n6046) );
  NAND U7266 ( .A(n6047), .B(n6046), .Z(n6200) );
  NANDN U7267 ( .A(n6049), .B(n6048), .Z(n6053) );
  NAND U7268 ( .A(n6051), .B(n6050), .Z(n6052) );
  AND U7269 ( .A(n6053), .B(n6052), .Z(n6199) );
  XNOR U7270 ( .A(n6200), .B(n6199), .Z(n6201) );
  XOR U7271 ( .A(n6202), .B(n6201), .Z(n6079) );
  NANDN U7272 ( .A(n6055), .B(n6054), .Z(n6059) );
  NAND U7273 ( .A(n6057), .B(n6056), .Z(n6058) );
  NAND U7274 ( .A(n6059), .B(n6058), .Z(n6077) );
  NANDN U7275 ( .A(n6061), .B(n6060), .Z(n6065) );
  NANDN U7276 ( .A(n6063), .B(n6062), .Z(n6064) );
  NAND U7277 ( .A(n6065), .B(n6064), .Z(n6078) );
  XNOR U7278 ( .A(n6077), .B(n6078), .Z(n6080) );
  XOR U7279 ( .A(n6079), .B(n6080), .Z(n6071) );
  XOR U7280 ( .A(n6072), .B(n6071), .Z(n6073) );
  XNOR U7281 ( .A(n6074), .B(n6073), .Z(n6211) );
  XNOR U7282 ( .A(n6211), .B(sreg[274]), .Z(n6213) );
  NAND U7283 ( .A(n6066), .B(sreg[273]), .Z(n6070) );
  OR U7284 ( .A(n6068), .B(n6067), .Z(n6069) );
  AND U7285 ( .A(n6070), .B(n6069), .Z(n6212) );
  XOR U7286 ( .A(n6213), .B(n6212), .Z(c[274]) );
  NAND U7287 ( .A(n6072), .B(n6071), .Z(n6076) );
  NAND U7288 ( .A(n6074), .B(n6073), .Z(n6075) );
  NAND U7289 ( .A(n6076), .B(n6075), .Z(n6219) );
  NANDN U7290 ( .A(n6078), .B(n6077), .Z(n6082) );
  NAND U7291 ( .A(n6080), .B(n6079), .Z(n6081) );
  NAND U7292 ( .A(n6082), .B(n6081), .Z(n6216) );
  NAND U7293 ( .A(n6084), .B(n6083), .Z(n6088) );
  NANDN U7294 ( .A(n6086), .B(n6085), .Z(n6087) );
  NAND U7295 ( .A(n6088), .B(n6087), .Z(n6346) );
  XNOR U7296 ( .A(n6346), .B(n6347), .Z(n6348) );
  NANDN U7297 ( .A(n6094), .B(n6093), .Z(n6098) );
  NANDN U7298 ( .A(n6096), .B(n6095), .Z(n6097) );
  NAND U7299 ( .A(n6098), .B(n6097), .Z(n6337) );
  OR U7300 ( .A(n6100), .B(n6099), .Z(n6104) );
  NAND U7301 ( .A(n6102), .B(n6101), .Z(n6103) );
  NAND U7302 ( .A(n6104), .B(n6103), .Z(n6276) );
  OR U7303 ( .A(n6106), .B(n6105), .Z(n6110) );
  NANDN U7304 ( .A(n6108), .B(n6107), .Z(n6109) );
  NAND U7305 ( .A(n6110), .B(n6109), .Z(n6275) );
  OR U7306 ( .A(n6112), .B(n6111), .Z(n6116) );
  NANDN U7307 ( .A(n6114), .B(n6113), .Z(n6115) );
  NAND U7308 ( .A(n6116), .B(n6115), .Z(n6274) );
  XOR U7309 ( .A(n6276), .B(n6277), .Z(n6334) );
  NANDN U7310 ( .A(n6118), .B(n6117), .Z(n6122) );
  NAND U7311 ( .A(n6120), .B(n6119), .Z(n6121) );
  NAND U7312 ( .A(n6122), .B(n6121), .Z(n6289) );
  XNOR U7313 ( .A(b[19]), .B(a[33]), .Z(n6234) );
  NANDN U7314 ( .A(n6234), .B(n37934), .Z(n6125) );
  NANDN U7315 ( .A(n6123), .B(n37935), .Z(n6124) );
  NAND U7316 ( .A(n6125), .B(n6124), .Z(n6301) );
  XNOR U7317 ( .A(b[27]), .B(a[25]), .Z(n6237) );
  NANDN U7318 ( .A(n6237), .B(n38423), .Z(n6128) );
  NAND U7319 ( .A(n6126), .B(n38424), .Z(n6127) );
  NAND U7320 ( .A(n6128), .B(n6127), .Z(n6298) );
  XNOR U7321 ( .A(b[5]), .B(a[47]), .Z(n6240) );
  NANDN U7322 ( .A(n6240), .B(n36587), .Z(n6131) );
  NANDN U7323 ( .A(n6129), .B(n36588), .Z(n6130) );
  AND U7324 ( .A(n6131), .B(n6130), .Z(n6299) );
  XNOR U7325 ( .A(n6298), .B(n6299), .Z(n6300) );
  XNOR U7326 ( .A(n6301), .B(n6300), .Z(n6287) );
  NAND U7327 ( .A(n6132), .B(n37762), .Z(n6134) );
  XOR U7328 ( .A(b[17]), .B(a[35]), .Z(n6243) );
  NAND U7329 ( .A(n6243), .B(n37764), .Z(n6133) );
  NAND U7330 ( .A(n6134), .B(n6133), .Z(n6261) );
  XNOR U7331 ( .A(b[31]), .B(a[21]), .Z(n6246) );
  NANDN U7332 ( .A(n6246), .B(n38552), .Z(n6137) );
  NANDN U7333 ( .A(n6135), .B(n38553), .Z(n6136) );
  NAND U7334 ( .A(n6137), .B(n6136), .Z(n6258) );
  OR U7335 ( .A(n6138), .B(n36105), .Z(n6140) );
  XNOR U7336 ( .A(b[3]), .B(a[49]), .Z(n6249) );
  NANDN U7337 ( .A(n6249), .B(n36107), .Z(n6139) );
  AND U7338 ( .A(n6140), .B(n6139), .Z(n6259) );
  XNOR U7339 ( .A(n6258), .B(n6259), .Z(n6260) );
  XOR U7340 ( .A(n6261), .B(n6260), .Z(n6286) );
  XNOR U7341 ( .A(n6287), .B(n6286), .Z(n6288) );
  XNOR U7342 ( .A(n6289), .B(n6288), .Z(n6335) );
  XNOR U7343 ( .A(n6334), .B(n6335), .Z(n6336) );
  XNOR U7344 ( .A(n6337), .B(n6336), .Z(n6355) );
  NANDN U7345 ( .A(n6146), .B(n6145), .Z(n6150) );
  NANDN U7346 ( .A(n6148), .B(n6147), .Z(n6149) );
  NAND U7347 ( .A(n6150), .B(n6149), .Z(n6342) );
  OR U7348 ( .A(n6152), .B(n6151), .Z(n6156) );
  NAND U7349 ( .A(n6154), .B(n6153), .Z(n6155) );
  NAND U7350 ( .A(n6156), .B(n6155), .Z(n6341) );
  NANDN U7351 ( .A(n6158), .B(n6157), .Z(n6162) );
  NAND U7352 ( .A(n6160), .B(n6159), .Z(n6161) );
  NAND U7353 ( .A(n6162), .B(n6161), .Z(n6280) );
  NANDN U7354 ( .A(n6164), .B(n6163), .Z(n6168) );
  NAND U7355 ( .A(n6166), .B(n6165), .Z(n6167) );
  AND U7356 ( .A(n6168), .B(n6167), .Z(n6281) );
  XNOR U7357 ( .A(n6280), .B(n6281), .Z(n6282) );
  XNOR U7358 ( .A(b[9]), .B(a[43]), .Z(n6304) );
  NANDN U7359 ( .A(n6304), .B(n36925), .Z(n6171) );
  NAND U7360 ( .A(n36926), .B(n6169), .Z(n6170) );
  NAND U7361 ( .A(n6171), .B(n6170), .Z(n6266) );
  XNOR U7362 ( .A(n1054), .B(a[37]), .Z(n6307) );
  NANDN U7363 ( .A(n37665), .B(n6307), .Z(n6174) );
  NANDN U7364 ( .A(n6172), .B(n37604), .Z(n6173) );
  NAND U7365 ( .A(n6174), .B(n6173), .Z(n6264) );
  XOR U7366 ( .A(b[21]), .B(n7955), .Z(n6310) );
  NANDN U7367 ( .A(n6310), .B(n38101), .Z(n6177) );
  NAND U7368 ( .A(n38102), .B(n6175), .Z(n6176) );
  NAND U7369 ( .A(n6177), .B(n6176), .Z(n6265) );
  XNOR U7370 ( .A(n6264), .B(n6265), .Z(n6267) );
  XOR U7371 ( .A(n6266), .B(n6267), .Z(n6255) );
  XNOR U7372 ( .A(b[11]), .B(a[41]), .Z(n6313) );
  OR U7373 ( .A(n6313), .B(n37311), .Z(n6180) );
  NANDN U7374 ( .A(n6178), .B(n37218), .Z(n6179) );
  NAND U7375 ( .A(n6180), .B(n6179), .Z(n6253) );
  XOR U7376 ( .A(n1053), .B(a[39]), .Z(n6316) );
  NANDN U7377 ( .A(n6316), .B(n37424), .Z(n6183) );
  NANDN U7378 ( .A(n6181), .B(n37425), .Z(n6182) );
  AND U7379 ( .A(n6183), .B(n6182), .Z(n6252) );
  XNOR U7380 ( .A(n6253), .B(n6252), .Z(n6254) );
  XNOR U7381 ( .A(n6255), .B(n6254), .Z(n6271) );
  NANDN U7382 ( .A(n1049), .B(a[51]), .Z(n6184) );
  XNOR U7383 ( .A(b[1]), .B(n6184), .Z(n6186) );
  IV U7384 ( .A(a[50]), .Z(n10724) );
  NANDN U7385 ( .A(n10724), .B(n1049), .Z(n6185) );
  AND U7386 ( .A(n6186), .B(n6185), .Z(n6230) );
  NAND U7387 ( .A(n38490), .B(n6187), .Z(n6189) );
  XNOR U7388 ( .A(n1058), .B(a[23]), .Z(n6322) );
  NANDN U7389 ( .A(n1048), .B(n6322), .Z(n6188) );
  NAND U7390 ( .A(n6189), .B(n6188), .Z(n6228) );
  NANDN U7391 ( .A(n1059), .B(a[19]), .Z(n6229) );
  XNOR U7392 ( .A(n6228), .B(n6229), .Z(n6231) );
  XNOR U7393 ( .A(n6230), .B(n6231), .Z(n6269) );
  NANDN U7394 ( .A(n6190), .B(n38205), .Z(n6192) );
  XNOR U7395 ( .A(b[23]), .B(a[29]), .Z(n6325) );
  OR U7396 ( .A(n6325), .B(n38268), .Z(n6191) );
  NAND U7397 ( .A(n6192), .B(n6191), .Z(n6295) );
  XOR U7398 ( .A(b[7]), .B(a[45]), .Z(n6328) );
  NAND U7399 ( .A(n6328), .B(n36701), .Z(n6195) );
  NANDN U7400 ( .A(n6193), .B(n36702), .Z(n6194) );
  NAND U7401 ( .A(n6195), .B(n6194), .Z(n6292) );
  XOR U7402 ( .A(b[25]), .B(a[27]), .Z(n6331) );
  NAND U7403 ( .A(n6331), .B(n38325), .Z(n6198) );
  NANDN U7404 ( .A(n6196), .B(n38326), .Z(n6197) );
  AND U7405 ( .A(n6198), .B(n6197), .Z(n6293) );
  XNOR U7406 ( .A(n6292), .B(n6293), .Z(n6294) );
  XOR U7407 ( .A(n6295), .B(n6294), .Z(n6268) );
  XOR U7408 ( .A(n6271), .B(n6270), .Z(n6283) );
  XOR U7409 ( .A(n6282), .B(n6283), .Z(n6340) );
  XNOR U7410 ( .A(n6341), .B(n6340), .Z(n6343) );
  XNOR U7411 ( .A(n6342), .B(n6343), .Z(n6352) );
  XNOR U7412 ( .A(n6353), .B(n6352), .Z(n6354) );
  XOR U7413 ( .A(n6355), .B(n6354), .Z(n6349) );
  XOR U7414 ( .A(n6348), .B(n6349), .Z(n6225) );
  NANDN U7415 ( .A(n6200), .B(n6199), .Z(n6204) );
  NAND U7416 ( .A(n6202), .B(n6201), .Z(n6203) );
  NAND U7417 ( .A(n6204), .B(n6203), .Z(n6222) );
  NANDN U7418 ( .A(n6206), .B(n6205), .Z(n6210) );
  OR U7419 ( .A(n6208), .B(n6207), .Z(n6209) );
  NAND U7420 ( .A(n6210), .B(n6209), .Z(n6223) );
  XNOR U7421 ( .A(n6222), .B(n6223), .Z(n6224) );
  XNOR U7422 ( .A(n6225), .B(n6224), .Z(n6217) );
  XNOR U7423 ( .A(n6216), .B(n6217), .Z(n6218) );
  XNOR U7424 ( .A(n6219), .B(n6218), .Z(n6358) );
  XNOR U7425 ( .A(n6358), .B(sreg[275]), .Z(n6360) );
  NAND U7426 ( .A(n6211), .B(sreg[274]), .Z(n6215) );
  OR U7427 ( .A(n6213), .B(n6212), .Z(n6214) );
  AND U7428 ( .A(n6215), .B(n6214), .Z(n6359) );
  XOR U7429 ( .A(n6360), .B(n6359), .Z(c[275]) );
  NANDN U7430 ( .A(n6217), .B(n6216), .Z(n6221) );
  NAND U7431 ( .A(n6219), .B(n6218), .Z(n6220) );
  NAND U7432 ( .A(n6221), .B(n6220), .Z(n6366) );
  NANDN U7433 ( .A(n6223), .B(n6222), .Z(n6227) );
  NAND U7434 ( .A(n6225), .B(n6224), .Z(n6226) );
  NAND U7435 ( .A(n6227), .B(n6226), .Z(n6364) );
  NANDN U7436 ( .A(n6229), .B(n6228), .Z(n6233) );
  NAND U7437 ( .A(n6231), .B(n6230), .Z(n6232) );
  NAND U7438 ( .A(n6233), .B(n6232), .Z(n6446) );
  XNOR U7439 ( .A(b[19]), .B(a[34]), .Z(n6391) );
  NANDN U7440 ( .A(n6391), .B(n37934), .Z(n6236) );
  NANDN U7441 ( .A(n6234), .B(n37935), .Z(n6235) );
  NAND U7442 ( .A(n6236), .B(n6235), .Z(n6456) );
  XNOR U7443 ( .A(b[27]), .B(a[26]), .Z(n6394) );
  NANDN U7444 ( .A(n6394), .B(n38423), .Z(n6239) );
  NANDN U7445 ( .A(n6237), .B(n38424), .Z(n6238) );
  NAND U7446 ( .A(n6239), .B(n6238), .Z(n6453) );
  XNOR U7447 ( .A(b[5]), .B(a[48]), .Z(n6397) );
  NANDN U7448 ( .A(n6397), .B(n36587), .Z(n6242) );
  NANDN U7449 ( .A(n6240), .B(n36588), .Z(n6241) );
  AND U7450 ( .A(n6242), .B(n6241), .Z(n6454) );
  XNOR U7451 ( .A(n6453), .B(n6454), .Z(n6455) );
  XNOR U7452 ( .A(n6456), .B(n6455), .Z(n6444) );
  NAND U7453 ( .A(n6243), .B(n37762), .Z(n6245) );
  XOR U7454 ( .A(b[17]), .B(a[36]), .Z(n6400) );
  NAND U7455 ( .A(n6400), .B(n37764), .Z(n6244) );
  NAND U7456 ( .A(n6245), .B(n6244), .Z(n6418) );
  XNOR U7457 ( .A(b[31]), .B(a[22]), .Z(n6403) );
  NANDN U7458 ( .A(n6403), .B(n38552), .Z(n6248) );
  NANDN U7459 ( .A(n6246), .B(n38553), .Z(n6247) );
  NAND U7460 ( .A(n6248), .B(n6247), .Z(n6415) );
  OR U7461 ( .A(n6249), .B(n36105), .Z(n6251) );
  XOR U7462 ( .A(b[3]), .B(n10724), .Z(n6406) );
  NANDN U7463 ( .A(n6406), .B(n36107), .Z(n6250) );
  AND U7464 ( .A(n6251), .B(n6250), .Z(n6416) );
  XNOR U7465 ( .A(n6415), .B(n6416), .Z(n6417) );
  XOR U7466 ( .A(n6418), .B(n6417), .Z(n6443) );
  XNOR U7467 ( .A(n6444), .B(n6443), .Z(n6445) );
  XNOR U7468 ( .A(n6446), .B(n6445), .Z(n6382) );
  NANDN U7469 ( .A(n6253), .B(n6252), .Z(n6257) );
  NAND U7470 ( .A(n6255), .B(n6254), .Z(n6256) );
  NAND U7471 ( .A(n6257), .B(n6256), .Z(n6435) );
  NANDN U7472 ( .A(n6259), .B(n6258), .Z(n6263) );
  NAND U7473 ( .A(n6261), .B(n6260), .Z(n6262) );
  NAND U7474 ( .A(n6263), .B(n6262), .Z(n6434) );
  XNOR U7475 ( .A(n6434), .B(n6433), .Z(n6436) );
  XOR U7476 ( .A(n6435), .B(n6436), .Z(n6381) );
  XOR U7477 ( .A(n6382), .B(n6381), .Z(n6383) );
  NANDN U7478 ( .A(n6269), .B(n6268), .Z(n6273) );
  NAND U7479 ( .A(n6271), .B(n6270), .Z(n6272) );
  NAND U7480 ( .A(n6273), .B(n6272), .Z(n6384) );
  XNOR U7481 ( .A(n6383), .B(n6384), .Z(n6497) );
  OR U7482 ( .A(n6275), .B(n6274), .Z(n6279) );
  NANDN U7483 ( .A(n6277), .B(n6276), .Z(n6278) );
  NAND U7484 ( .A(n6279), .B(n6278), .Z(n6496) );
  NANDN U7485 ( .A(n6281), .B(n6280), .Z(n6285) );
  NAND U7486 ( .A(n6283), .B(n6282), .Z(n6284) );
  NAND U7487 ( .A(n6285), .B(n6284), .Z(n6377) );
  NANDN U7488 ( .A(n6287), .B(n6286), .Z(n6291) );
  NAND U7489 ( .A(n6289), .B(n6288), .Z(n6290) );
  NAND U7490 ( .A(n6291), .B(n6290), .Z(n6376) );
  NANDN U7491 ( .A(n6293), .B(n6292), .Z(n6297) );
  NAND U7492 ( .A(n6295), .B(n6294), .Z(n6296) );
  NAND U7493 ( .A(n6297), .B(n6296), .Z(n6437) );
  NANDN U7494 ( .A(n6299), .B(n6298), .Z(n6303) );
  NAND U7495 ( .A(n6301), .B(n6300), .Z(n6302) );
  AND U7496 ( .A(n6303), .B(n6302), .Z(n6438) );
  XNOR U7497 ( .A(n6437), .B(n6438), .Z(n6439) );
  XOR U7498 ( .A(b[9]), .B(n9873), .Z(n6459) );
  NANDN U7499 ( .A(n6459), .B(n36925), .Z(n6306) );
  NANDN U7500 ( .A(n6304), .B(n36926), .Z(n6305) );
  NAND U7501 ( .A(n6306), .B(n6305), .Z(n6423) );
  XNOR U7502 ( .A(b[15]), .B(a[38]), .Z(n6462) );
  OR U7503 ( .A(n6462), .B(n37665), .Z(n6309) );
  NAND U7504 ( .A(n6307), .B(n37604), .Z(n6308) );
  AND U7505 ( .A(n6309), .B(n6308), .Z(n6421) );
  XNOR U7506 ( .A(b[21]), .B(a[32]), .Z(n6465) );
  NANDN U7507 ( .A(n6465), .B(n38101), .Z(n6312) );
  NANDN U7508 ( .A(n6310), .B(n38102), .Z(n6311) );
  AND U7509 ( .A(n6312), .B(n6311), .Z(n6422) );
  XOR U7510 ( .A(n6423), .B(n6424), .Z(n6412) );
  XNOR U7511 ( .A(b[11]), .B(a[42]), .Z(n6468) );
  OR U7512 ( .A(n6468), .B(n37311), .Z(n6315) );
  NANDN U7513 ( .A(n6313), .B(n37218), .Z(n6314) );
  NAND U7514 ( .A(n6315), .B(n6314), .Z(n6410) );
  XOR U7515 ( .A(n1053), .B(a[40]), .Z(n6471) );
  NANDN U7516 ( .A(n6471), .B(n37424), .Z(n6318) );
  NANDN U7517 ( .A(n6316), .B(n37425), .Z(n6317) );
  AND U7518 ( .A(n6318), .B(n6317), .Z(n6409) );
  XNOR U7519 ( .A(n6410), .B(n6409), .Z(n6411) );
  XOR U7520 ( .A(n6412), .B(n6411), .Z(n6429) );
  NANDN U7521 ( .A(n1049), .B(a[52]), .Z(n6319) );
  XNOR U7522 ( .A(b[1]), .B(n6319), .Z(n6321) );
  NANDN U7523 ( .A(b[0]), .B(a[51]), .Z(n6320) );
  AND U7524 ( .A(n6321), .B(n6320), .Z(n6387) );
  NAND U7525 ( .A(n38490), .B(n6322), .Z(n6324) );
  XNOR U7526 ( .A(n1058), .B(a[24]), .Z(n6477) );
  NANDN U7527 ( .A(n1048), .B(n6477), .Z(n6323) );
  NAND U7528 ( .A(n6324), .B(n6323), .Z(n6385) );
  NANDN U7529 ( .A(n1059), .B(a[20]), .Z(n6386) );
  XNOR U7530 ( .A(n6385), .B(n6386), .Z(n6388) );
  XOR U7531 ( .A(n6387), .B(n6388), .Z(n6427) );
  NANDN U7532 ( .A(n6325), .B(n38205), .Z(n6327) );
  XOR U7533 ( .A(b[23]), .B(n7434), .Z(n6480) );
  OR U7534 ( .A(n6480), .B(n38268), .Z(n6326) );
  NAND U7535 ( .A(n6327), .B(n6326), .Z(n6450) );
  XOR U7536 ( .A(b[7]), .B(a[46]), .Z(n6483) );
  NAND U7537 ( .A(n6483), .B(n36701), .Z(n6330) );
  NAND U7538 ( .A(n6328), .B(n36702), .Z(n6329) );
  NAND U7539 ( .A(n6330), .B(n6329), .Z(n6447) );
  XOR U7540 ( .A(b[25]), .B(a[28]), .Z(n6486) );
  NAND U7541 ( .A(n6486), .B(n38325), .Z(n6333) );
  NAND U7542 ( .A(n6331), .B(n38326), .Z(n6332) );
  AND U7543 ( .A(n6333), .B(n6332), .Z(n6448) );
  XNOR U7544 ( .A(n6447), .B(n6448), .Z(n6449) );
  XNOR U7545 ( .A(n6450), .B(n6449), .Z(n6428) );
  XOR U7546 ( .A(n6427), .B(n6428), .Z(n6430) );
  XNOR U7547 ( .A(n6429), .B(n6430), .Z(n6440) );
  XNOR U7548 ( .A(n6439), .B(n6440), .Z(n6375) );
  XNOR U7549 ( .A(n6376), .B(n6375), .Z(n6378) );
  XNOR U7550 ( .A(n6377), .B(n6378), .Z(n6495) );
  XOR U7551 ( .A(n6496), .B(n6495), .Z(n6498) );
  NANDN U7552 ( .A(n6335), .B(n6334), .Z(n6339) );
  NAND U7553 ( .A(n6337), .B(n6336), .Z(n6338) );
  NAND U7554 ( .A(n6339), .B(n6338), .Z(n6490) );
  NAND U7555 ( .A(n6341), .B(n6340), .Z(n6345) );
  NANDN U7556 ( .A(n6343), .B(n6342), .Z(n6344) );
  AND U7557 ( .A(n6345), .B(n6344), .Z(n6489) );
  XNOR U7558 ( .A(n6490), .B(n6489), .Z(n6491) );
  XOR U7559 ( .A(n6492), .B(n6491), .Z(n6371) );
  NANDN U7560 ( .A(n6347), .B(n6346), .Z(n6351) );
  NANDN U7561 ( .A(n6349), .B(n6348), .Z(n6350) );
  NAND U7562 ( .A(n6351), .B(n6350), .Z(n6370) );
  NANDN U7563 ( .A(n6353), .B(n6352), .Z(n6357) );
  NANDN U7564 ( .A(n6355), .B(n6354), .Z(n6356) );
  AND U7565 ( .A(n6357), .B(n6356), .Z(n6369) );
  XNOR U7566 ( .A(n6370), .B(n6369), .Z(n6372) );
  XOR U7567 ( .A(n6371), .B(n6372), .Z(n6363) );
  XOR U7568 ( .A(n6364), .B(n6363), .Z(n6365) );
  XNOR U7569 ( .A(n6366), .B(n6365), .Z(n6501) );
  XNOR U7570 ( .A(n6501), .B(sreg[276]), .Z(n6503) );
  NAND U7571 ( .A(n6358), .B(sreg[275]), .Z(n6362) );
  OR U7572 ( .A(n6360), .B(n6359), .Z(n6361) );
  AND U7573 ( .A(n6362), .B(n6361), .Z(n6502) );
  XOR U7574 ( .A(n6503), .B(n6502), .Z(c[276]) );
  NAND U7575 ( .A(n6364), .B(n6363), .Z(n6368) );
  NAND U7576 ( .A(n6366), .B(n6365), .Z(n6367) );
  NAND U7577 ( .A(n6368), .B(n6367), .Z(n6509) );
  NANDN U7578 ( .A(n6370), .B(n6369), .Z(n6374) );
  NAND U7579 ( .A(n6372), .B(n6371), .Z(n6373) );
  NAND U7580 ( .A(n6374), .B(n6373), .Z(n6506) );
  NAND U7581 ( .A(n6376), .B(n6375), .Z(n6380) );
  NANDN U7582 ( .A(n6378), .B(n6377), .Z(n6379) );
  NAND U7583 ( .A(n6380), .B(n6379), .Z(n6518) );
  XNOR U7584 ( .A(n6518), .B(n6519), .Z(n6520) );
  NANDN U7585 ( .A(n6386), .B(n6385), .Z(n6390) );
  NAND U7586 ( .A(n6388), .B(n6387), .Z(n6389) );
  NAND U7587 ( .A(n6390), .B(n6389), .Z(n6593) );
  XNOR U7588 ( .A(b[19]), .B(a[35]), .Z(n6536) );
  NANDN U7589 ( .A(n6536), .B(n37934), .Z(n6393) );
  NANDN U7590 ( .A(n6391), .B(n37935), .Z(n6392) );
  NAND U7591 ( .A(n6393), .B(n6392), .Z(n6603) );
  XOR U7592 ( .A(b[27]), .B(a[27]), .Z(n6539) );
  NAND U7593 ( .A(n38423), .B(n6539), .Z(n6396) );
  NANDN U7594 ( .A(n6394), .B(n38424), .Z(n6395) );
  NAND U7595 ( .A(n6396), .B(n6395), .Z(n6600) );
  XNOR U7596 ( .A(b[5]), .B(a[49]), .Z(n6542) );
  NANDN U7597 ( .A(n6542), .B(n36587), .Z(n6399) );
  NANDN U7598 ( .A(n6397), .B(n36588), .Z(n6398) );
  AND U7599 ( .A(n6399), .B(n6398), .Z(n6601) );
  XNOR U7600 ( .A(n6600), .B(n6601), .Z(n6602) );
  XNOR U7601 ( .A(n6603), .B(n6602), .Z(n6591) );
  NAND U7602 ( .A(n6400), .B(n37762), .Z(n6402) );
  XNOR U7603 ( .A(b[17]), .B(a[37]), .Z(n6545) );
  NANDN U7604 ( .A(n6545), .B(n37764), .Z(n6401) );
  NAND U7605 ( .A(n6402), .B(n6401), .Z(n6563) );
  XNOR U7606 ( .A(b[31]), .B(a[23]), .Z(n6548) );
  NANDN U7607 ( .A(n6548), .B(n38552), .Z(n6405) );
  NANDN U7608 ( .A(n6403), .B(n38553), .Z(n6404) );
  NAND U7609 ( .A(n6405), .B(n6404), .Z(n6560) );
  OR U7610 ( .A(n6406), .B(n36105), .Z(n6408) );
  XNOR U7611 ( .A(b[3]), .B(a[51]), .Z(n6551) );
  NANDN U7612 ( .A(n6551), .B(n36107), .Z(n6407) );
  AND U7613 ( .A(n6408), .B(n6407), .Z(n6561) );
  XNOR U7614 ( .A(n6560), .B(n6561), .Z(n6562) );
  XOR U7615 ( .A(n6563), .B(n6562), .Z(n6590) );
  XNOR U7616 ( .A(n6591), .B(n6590), .Z(n6592) );
  XNOR U7617 ( .A(n6593), .B(n6592), .Z(n6636) );
  NANDN U7618 ( .A(n6410), .B(n6409), .Z(n6414) );
  NAND U7619 ( .A(n6412), .B(n6411), .Z(n6413) );
  NAND U7620 ( .A(n6414), .B(n6413), .Z(n6581) );
  NANDN U7621 ( .A(n6416), .B(n6415), .Z(n6420) );
  NAND U7622 ( .A(n6418), .B(n6417), .Z(n6419) );
  NAND U7623 ( .A(n6420), .B(n6419), .Z(n6579) );
  OR U7624 ( .A(n6422), .B(n6421), .Z(n6426) );
  NANDN U7625 ( .A(n6424), .B(n6423), .Z(n6425) );
  NAND U7626 ( .A(n6426), .B(n6425), .Z(n6578) );
  XNOR U7627 ( .A(n6581), .B(n6580), .Z(n6637) );
  XNOR U7628 ( .A(n6636), .B(n6637), .Z(n6638) );
  NANDN U7629 ( .A(n6428), .B(n6427), .Z(n6432) );
  OR U7630 ( .A(n6430), .B(n6429), .Z(n6431) );
  AND U7631 ( .A(n6432), .B(n6431), .Z(n6639) );
  XOR U7632 ( .A(n6638), .B(n6639), .Z(n6526) );
  NANDN U7633 ( .A(n6438), .B(n6437), .Z(n6442) );
  NANDN U7634 ( .A(n6440), .B(n6439), .Z(n6441) );
  NAND U7635 ( .A(n6442), .B(n6441), .Z(n6645) );
  NANDN U7636 ( .A(n6448), .B(n6447), .Z(n6452) );
  NAND U7637 ( .A(n6450), .B(n6449), .Z(n6451) );
  NAND U7638 ( .A(n6452), .B(n6451), .Z(n6584) );
  NANDN U7639 ( .A(n6454), .B(n6453), .Z(n6458) );
  NAND U7640 ( .A(n6456), .B(n6455), .Z(n6457) );
  AND U7641 ( .A(n6458), .B(n6457), .Z(n6585) );
  XNOR U7642 ( .A(n6584), .B(n6585), .Z(n6586) );
  XNOR U7643 ( .A(b[9]), .B(a[45]), .Z(n6606) );
  NANDN U7644 ( .A(n6606), .B(n36925), .Z(n6461) );
  NANDN U7645 ( .A(n6459), .B(n36926), .Z(n6460) );
  NAND U7646 ( .A(n6461), .B(n6460), .Z(n6568) );
  XNOR U7647 ( .A(b[15]), .B(a[39]), .Z(n6609) );
  OR U7648 ( .A(n6609), .B(n37665), .Z(n6464) );
  NANDN U7649 ( .A(n6462), .B(n37604), .Z(n6463) );
  AND U7650 ( .A(n6464), .B(n6463), .Z(n6566) );
  XNOR U7651 ( .A(b[21]), .B(a[33]), .Z(n6612) );
  NANDN U7652 ( .A(n6612), .B(n38101), .Z(n6467) );
  NANDN U7653 ( .A(n6465), .B(n38102), .Z(n6466) );
  AND U7654 ( .A(n6467), .B(n6466), .Z(n6567) );
  XOR U7655 ( .A(n6568), .B(n6569), .Z(n6557) );
  XNOR U7656 ( .A(b[11]), .B(a[43]), .Z(n6615) );
  OR U7657 ( .A(n6615), .B(n37311), .Z(n6470) );
  NANDN U7658 ( .A(n6468), .B(n37218), .Z(n6469) );
  NAND U7659 ( .A(n6470), .B(n6469), .Z(n6555) );
  XOR U7660 ( .A(n1053), .B(a[41]), .Z(n6618) );
  NANDN U7661 ( .A(n6618), .B(n37424), .Z(n6473) );
  NANDN U7662 ( .A(n6471), .B(n37425), .Z(n6472) );
  AND U7663 ( .A(n6473), .B(n6472), .Z(n6554) );
  XNOR U7664 ( .A(n6555), .B(n6554), .Z(n6556) );
  XOR U7665 ( .A(n6557), .B(n6556), .Z(n6574) );
  NANDN U7666 ( .A(n1049), .B(a[53]), .Z(n6474) );
  XNOR U7667 ( .A(b[1]), .B(n6474), .Z(n6476) );
  NANDN U7668 ( .A(b[0]), .B(a[52]), .Z(n6475) );
  AND U7669 ( .A(n6476), .B(n6475), .Z(n6532) );
  NAND U7670 ( .A(n38490), .B(n6477), .Z(n6479) );
  XOR U7671 ( .A(n1058), .B(n7069), .Z(n6621) );
  NANDN U7672 ( .A(n1048), .B(n6621), .Z(n6478) );
  NAND U7673 ( .A(n6479), .B(n6478), .Z(n6530) );
  NANDN U7674 ( .A(n1059), .B(a[21]), .Z(n6531) );
  XNOR U7675 ( .A(n6530), .B(n6531), .Z(n6533) );
  XOR U7676 ( .A(n6532), .B(n6533), .Z(n6572) );
  NANDN U7677 ( .A(n6480), .B(n38205), .Z(n6482) );
  XOR U7678 ( .A(b[23]), .B(n7955), .Z(n6627) );
  OR U7679 ( .A(n6627), .B(n38268), .Z(n6481) );
  NAND U7680 ( .A(n6482), .B(n6481), .Z(n6597) );
  XOR U7681 ( .A(b[7]), .B(a[47]), .Z(n6630) );
  NAND U7682 ( .A(n6630), .B(n36701), .Z(n6485) );
  NAND U7683 ( .A(n6483), .B(n36702), .Z(n6484) );
  NAND U7684 ( .A(n6485), .B(n6484), .Z(n6594) );
  XOR U7685 ( .A(b[25]), .B(a[29]), .Z(n6633) );
  NAND U7686 ( .A(n6633), .B(n38325), .Z(n6488) );
  NAND U7687 ( .A(n6486), .B(n38326), .Z(n6487) );
  AND U7688 ( .A(n6488), .B(n6487), .Z(n6595) );
  XNOR U7689 ( .A(n6594), .B(n6595), .Z(n6596) );
  XNOR U7690 ( .A(n6597), .B(n6596), .Z(n6573) );
  XOR U7691 ( .A(n6572), .B(n6573), .Z(n6575) );
  XNOR U7692 ( .A(n6574), .B(n6575), .Z(n6587) );
  XOR U7693 ( .A(n6586), .B(n6587), .Z(n6643) );
  XNOR U7694 ( .A(n6642), .B(n6643), .Z(n6644) );
  XNOR U7695 ( .A(n6645), .B(n6644), .Z(n6524) );
  XNOR U7696 ( .A(n6525), .B(n6524), .Z(n6527) );
  XNOR U7697 ( .A(n6526), .B(n6527), .Z(n6521) );
  XOR U7698 ( .A(n6520), .B(n6521), .Z(n6515) );
  NANDN U7699 ( .A(n6490), .B(n6489), .Z(n6494) );
  NAND U7700 ( .A(n6492), .B(n6491), .Z(n6493) );
  NAND U7701 ( .A(n6494), .B(n6493), .Z(n6512) );
  NANDN U7702 ( .A(n6496), .B(n6495), .Z(n6500) );
  OR U7703 ( .A(n6498), .B(n6497), .Z(n6499) );
  NAND U7704 ( .A(n6500), .B(n6499), .Z(n6513) );
  XNOR U7705 ( .A(n6512), .B(n6513), .Z(n6514) );
  XNOR U7706 ( .A(n6515), .B(n6514), .Z(n6507) );
  XNOR U7707 ( .A(n6506), .B(n6507), .Z(n6508) );
  XNOR U7708 ( .A(n6509), .B(n6508), .Z(n6648) );
  XNOR U7709 ( .A(n6648), .B(sreg[277]), .Z(n6650) );
  NAND U7710 ( .A(n6501), .B(sreg[276]), .Z(n6505) );
  OR U7711 ( .A(n6503), .B(n6502), .Z(n6504) );
  AND U7712 ( .A(n6505), .B(n6504), .Z(n6649) );
  XOR U7713 ( .A(n6650), .B(n6649), .Z(c[277]) );
  NANDN U7714 ( .A(n6507), .B(n6506), .Z(n6511) );
  NAND U7715 ( .A(n6509), .B(n6508), .Z(n6510) );
  NAND U7716 ( .A(n6511), .B(n6510), .Z(n6656) );
  NANDN U7717 ( .A(n6513), .B(n6512), .Z(n6517) );
  NAND U7718 ( .A(n6515), .B(n6514), .Z(n6516) );
  NAND U7719 ( .A(n6517), .B(n6516), .Z(n6654) );
  NANDN U7720 ( .A(n6519), .B(n6518), .Z(n6523) );
  NANDN U7721 ( .A(n6521), .B(n6520), .Z(n6522) );
  NAND U7722 ( .A(n6523), .B(n6522), .Z(n6660) );
  OR U7723 ( .A(n6525), .B(n6524), .Z(n6529) );
  OR U7724 ( .A(n6527), .B(n6526), .Z(n6528) );
  AND U7725 ( .A(n6529), .B(n6528), .Z(n6659) );
  XNOR U7726 ( .A(n6660), .B(n6659), .Z(n6661) );
  NANDN U7727 ( .A(n6531), .B(n6530), .Z(n6535) );
  NAND U7728 ( .A(n6533), .B(n6532), .Z(n6534) );
  NAND U7729 ( .A(n6535), .B(n6534), .Z(n6740) );
  XNOR U7730 ( .A(b[19]), .B(a[36]), .Z(n6707) );
  NANDN U7731 ( .A(n6707), .B(n37934), .Z(n6538) );
  NANDN U7732 ( .A(n6536), .B(n37935), .Z(n6537) );
  NAND U7733 ( .A(n6538), .B(n6537), .Z(n6776) );
  XOR U7734 ( .A(b[27]), .B(a[28]), .Z(n6710) );
  NAND U7735 ( .A(n38423), .B(n6710), .Z(n6541) );
  NAND U7736 ( .A(n6539), .B(n38424), .Z(n6540) );
  NAND U7737 ( .A(n6541), .B(n6540), .Z(n6773) );
  XOR U7738 ( .A(b[5]), .B(n10724), .Z(n6713) );
  NANDN U7739 ( .A(n6713), .B(n36587), .Z(n6544) );
  NANDN U7740 ( .A(n6542), .B(n36588), .Z(n6543) );
  AND U7741 ( .A(n6544), .B(n6543), .Z(n6774) );
  XNOR U7742 ( .A(n6773), .B(n6774), .Z(n6775) );
  XNOR U7743 ( .A(n6776), .B(n6775), .Z(n6737) );
  NANDN U7744 ( .A(n6545), .B(n37762), .Z(n6547) );
  XOR U7745 ( .A(b[17]), .B(a[38]), .Z(n6716) );
  NAND U7746 ( .A(n6716), .B(n37764), .Z(n6546) );
  NAND U7747 ( .A(n6547), .B(n6546), .Z(n6691) );
  XNOR U7748 ( .A(b[31]), .B(a[24]), .Z(n6719) );
  NANDN U7749 ( .A(n6719), .B(n38552), .Z(n6550) );
  NANDN U7750 ( .A(n6548), .B(n38553), .Z(n6549) );
  AND U7751 ( .A(n6550), .B(n6549), .Z(n6689) );
  OR U7752 ( .A(n6551), .B(n36105), .Z(n6553) );
  XNOR U7753 ( .A(b[3]), .B(a[52]), .Z(n6722) );
  NANDN U7754 ( .A(n6722), .B(n36107), .Z(n6552) );
  AND U7755 ( .A(n6553), .B(n6552), .Z(n6690) );
  XOR U7756 ( .A(n6691), .B(n6692), .Z(n6738) );
  XOR U7757 ( .A(n6737), .B(n6738), .Z(n6739) );
  XNOR U7758 ( .A(n6740), .B(n6739), .Z(n6785) );
  NANDN U7759 ( .A(n6555), .B(n6554), .Z(n6559) );
  NAND U7760 ( .A(n6557), .B(n6556), .Z(n6558) );
  NAND U7761 ( .A(n6559), .B(n6558), .Z(n6728) );
  NANDN U7762 ( .A(n6561), .B(n6560), .Z(n6565) );
  NAND U7763 ( .A(n6563), .B(n6562), .Z(n6564) );
  NAND U7764 ( .A(n6565), .B(n6564), .Z(n6726) );
  OR U7765 ( .A(n6567), .B(n6566), .Z(n6571) );
  NANDN U7766 ( .A(n6569), .B(n6568), .Z(n6570) );
  NAND U7767 ( .A(n6571), .B(n6570), .Z(n6725) );
  XNOR U7768 ( .A(n6728), .B(n6727), .Z(n6786) );
  XOR U7769 ( .A(n6785), .B(n6786), .Z(n6788) );
  NANDN U7770 ( .A(n6573), .B(n6572), .Z(n6577) );
  OR U7771 ( .A(n6575), .B(n6574), .Z(n6576) );
  NAND U7772 ( .A(n6577), .B(n6576), .Z(n6787) );
  XOR U7773 ( .A(n6788), .B(n6787), .Z(n6673) );
  OR U7774 ( .A(n6579), .B(n6578), .Z(n6583) );
  NAND U7775 ( .A(n6581), .B(n6580), .Z(n6582) );
  NAND U7776 ( .A(n6583), .B(n6582), .Z(n6672) );
  NANDN U7777 ( .A(n6585), .B(n6584), .Z(n6589) );
  NANDN U7778 ( .A(n6587), .B(n6586), .Z(n6588) );
  NAND U7779 ( .A(n6589), .B(n6588), .Z(n6793) );
  NANDN U7780 ( .A(n6595), .B(n6594), .Z(n6599) );
  NAND U7781 ( .A(n6597), .B(n6596), .Z(n6598) );
  NAND U7782 ( .A(n6599), .B(n6598), .Z(n6731) );
  NANDN U7783 ( .A(n6601), .B(n6600), .Z(n6605) );
  NAND U7784 ( .A(n6603), .B(n6602), .Z(n6604) );
  AND U7785 ( .A(n6605), .B(n6604), .Z(n6732) );
  XNOR U7786 ( .A(n6731), .B(n6732), .Z(n6733) );
  XNOR U7787 ( .A(b[9]), .B(a[46]), .Z(n6743) );
  NANDN U7788 ( .A(n6743), .B(n36925), .Z(n6608) );
  NANDN U7789 ( .A(n6606), .B(n36926), .Z(n6607) );
  NAND U7790 ( .A(n6608), .B(n6607), .Z(n6697) );
  XNOR U7791 ( .A(b[15]), .B(a[40]), .Z(n6746) );
  OR U7792 ( .A(n6746), .B(n37665), .Z(n6611) );
  NANDN U7793 ( .A(n6609), .B(n37604), .Z(n6610) );
  AND U7794 ( .A(n6611), .B(n6610), .Z(n6695) );
  XNOR U7795 ( .A(b[21]), .B(a[34]), .Z(n6749) );
  NANDN U7796 ( .A(n6749), .B(n38101), .Z(n6614) );
  NANDN U7797 ( .A(n6612), .B(n38102), .Z(n6613) );
  AND U7798 ( .A(n6614), .B(n6613), .Z(n6696) );
  XOR U7799 ( .A(n6697), .B(n6698), .Z(n6686) );
  XOR U7800 ( .A(b[11]), .B(n9873), .Z(n6752) );
  OR U7801 ( .A(n6752), .B(n37311), .Z(n6617) );
  NANDN U7802 ( .A(n6615), .B(n37218), .Z(n6616) );
  NAND U7803 ( .A(n6617), .B(n6616), .Z(n6684) );
  XOR U7804 ( .A(n1053), .B(a[42]), .Z(n6755) );
  NANDN U7805 ( .A(n6755), .B(n37424), .Z(n6620) );
  NANDN U7806 ( .A(n6618), .B(n37425), .Z(n6619) );
  NAND U7807 ( .A(n6620), .B(n6619), .Z(n6683) );
  XOR U7808 ( .A(n6686), .B(n6685), .Z(n6680) );
  NAND U7809 ( .A(n38490), .B(n6621), .Z(n6623) );
  XOR U7810 ( .A(n1058), .B(n7202), .Z(n6761) );
  NANDN U7811 ( .A(n1048), .B(n6761), .Z(n6622) );
  NAND U7812 ( .A(n6623), .B(n6622), .Z(n6701) );
  NANDN U7813 ( .A(n1059), .B(a[22]), .Z(n6702) );
  XNOR U7814 ( .A(n6701), .B(n6702), .Z(n6704) );
  NANDN U7815 ( .A(n1049), .B(a[54]), .Z(n6624) );
  XNOR U7816 ( .A(b[1]), .B(n6624), .Z(n6626) );
  NANDN U7817 ( .A(b[0]), .B(a[53]), .Z(n6625) );
  AND U7818 ( .A(n6626), .B(n6625), .Z(n6703) );
  XNOR U7819 ( .A(n6704), .B(n6703), .Z(n6678) );
  NANDN U7820 ( .A(n6627), .B(n38205), .Z(n6629) );
  XNOR U7821 ( .A(b[23]), .B(a[32]), .Z(n6764) );
  OR U7822 ( .A(n6764), .B(n38268), .Z(n6628) );
  NAND U7823 ( .A(n6629), .B(n6628), .Z(n6782) );
  XOR U7824 ( .A(b[7]), .B(a[48]), .Z(n6767) );
  NAND U7825 ( .A(n6767), .B(n36701), .Z(n6632) );
  NAND U7826 ( .A(n6630), .B(n36702), .Z(n6631) );
  NAND U7827 ( .A(n6632), .B(n6631), .Z(n6779) );
  XNOR U7828 ( .A(b[25]), .B(a[30]), .Z(n6770) );
  NANDN U7829 ( .A(n6770), .B(n38325), .Z(n6635) );
  NAND U7830 ( .A(n6633), .B(n38326), .Z(n6634) );
  AND U7831 ( .A(n6635), .B(n6634), .Z(n6780) );
  XNOR U7832 ( .A(n6779), .B(n6780), .Z(n6781) );
  XOR U7833 ( .A(n6782), .B(n6781), .Z(n6677) );
  XOR U7834 ( .A(n6680), .B(n6679), .Z(n6734) );
  XNOR U7835 ( .A(n6733), .B(n6734), .Z(n6791) );
  XNOR U7836 ( .A(n6792), .B(n6791), .Z(n6794) );
  XNOR U7837 ( .A(n6793), .B(n6794), .Z(n6671) );
  XOR U7838 ( .A(n6672), .B(n6671), .Z(n6674) );
  NANDN U7839 ( .A(n6637), .B(n6636), .Z(n6641) );
  NAND U7840 ( .A(n6639), .B(n6638), .Z(n6640) );
  NAND U7841 ( .A(n6641), .B(n6640), .Z(n6665) );
  NANDN U7842 ( .A(n6643), .B(n6642), .Z(n6647) );
  NAND U7843 ( .A(n6645), .B(n6644), .Z(n6646) );
  NAND U7844 ( .A(n6647), .B(n6646), .Z(n6666) );
  XNOR U7845 ( .A(n6665), .B(n6666), .Z(n6667) );
  XOR U7846 ( .A(n6668), .B(n6667), .Z(n6662) );
  XOR U7847 ( .A(n6661), .B(n6662), .Z(n6653) );
  XOR U7848 ( .A(n6654), .B(n6653), .Z(n6655) );
  XNOR U7849 ( .A(n6656), .B(n6655), .Z(n6797) );
  XNOR U7850 ( .A(n6797), .B(sreg[278]), .Z(n6799) );
  NAND U7851 ( .A(n6648), .B(sreg[277]), .Z(n6652) );
  OR U7852 ( .A(n6650), .B(n6649), .Z(n6651) );
  AND U7853 ( .A(n6652), .B(n6651), .Z(n6798) );
  XOR U7854 ( .A(n6799), .B(n6798), .Z(c[278]) );
  NAND U7855 ( .A(n6654), .B(n6653), .Z(n6658) );
  NAND U7856 ( .A(n6656), .B(n6655), .Z(n6657) );
  NAND U7857 ( .A(n6658), .B(n6657), .Z(n6805) );
  NANDN U7858 ( .A(n6660), .B(n6659), .Z(n6664) );
  NAND U7859 ( .A(n6662), .B(n6661), .Z(n6663) );
  NAND U7860 ( .A(n6664), .B(n6663), .Z(n6803) );
  NANDN U7861 ( .A(n6666), .B(n6665), .Z(n6670) );
  NAND U7862 ( .A(n6668), .B(n6667), .Z(n6669) );
  NAND U7863 ( .A(n6670), .B(n6669), .Z(n6808) );
  NANDN U7864 ( .A(n6672), .B(n6671), .Z(n6676) );
  OR U7865 ( .A(n6674), .B(n6673), .Z(n6675) );
  NAND U7866 ( .A(n6676), .B(n6675), .Z(n6809) );
  XNOR U7867 ( .A(n6808), .B(n6809), .Z(n6810) );
  NANDN U7868 ( .A(n6678), .B(n6677), .Z(n6682) );
  NANDN U7869 ( .A(n6680), .B(n6679), .Z(n6681) );
  NAND U7870 ( .A(n6682), .B(n6681), .Z(n6925) );
  OR U7871 ( .A(n6684), .B(n6683), .Z(n6688) );
  NAND U7872 ( .A(n6686), .B(n6685), .Z(n6687) );
  NAND U7873 ( .A(n6688), .B(n6687), .Z(n6864) );
  OR U7874 ( .A(n6690), .B(n6689), .Z(n6694) );
  NANDN U7875 ( .A(n6692), .B(n6691), .Z(n6693) );
  NAND U7876 ( .A(n6694), .B(n6693), .Z(n6863) );
  OR U7877 ( .A(n6696), .B(n6695), .Z(n6700) );
  NANDN U7878 ( .A(n6698), .B(n6697), .Z(n6699) );
  NAND U7879 ( .A(n6700), .B(n6699), .Z(n6862) );
  XOR U7880 ( .A(n6864), .B(n6865), .Z(n6922) );
  NANDN U7881 ( .A(n6702), .B(n6701), .Z(n6706) );
  NAND U7882 ( .A(n6704), .B(n6703), .Z(n6705) );
  NAND U7883 ( .A(n6706), .B(n6705), .Z(n6877) );
  XOR U7884 ( .A(b[19]), .B(n8832), .Z(n6820) );
  NANDN U7885 ( .A(n6820), .B(n37934), .Z(n6709) );
  NANDN U7886 ( .A(n6707), .B(n37935), .Z(n6708) );
  NAND U7887 ( .A(n6709), .B(n6708), .Z(n6889) );
  XOR U7888 ( .A(b[27]), .B(a[29]), .Z(n6823) );
  NAND U7889 ( .A(n38423), .B(n6823), .Z(n6712) );
  NAND U7890 ( .A(n6710), .B(n38424), .Z(n6711) );
  NAND U7891 ( .A(n6712), .B(n6711), .Z(n6886) );
  XNOR U7892 ( .A(b[5]), .B(a[51]), .Z(n6826) );
  NANDN U7893 ( .A(n6826), .B(n36587), .Z(n6715) );
  NANDN U7894 ( .A(n6713), .B(n36588), .Z(n6714) );
  AND U7895 ( .A(n6715), .B(n6714), .Z(n6887) );
  XNOR U7896 ( .A(n6886), .B(n6887), .Z(n6888) );
  XNOR U7897 ( .A(n6889), .B(n6888), .Z(n6875) );
  NAND U7898 ( .A(n6716), .B(n37762), .Z(n6718) );
  XOR U7899 ( .A(b[17]), .B(a[39]), .Z(n6829) );
  NAND U7900 ( .A(n6829), .B(n37764), .Z(n6717) );
  NAND U7901 ( .A(n6718), .B(n6717), .Z(n6847) );
  XOR U7902 ( .A(b[31]), .B(n7069), .Z(n6832) );
  NANDN U7903 ( .A(n6832), .B(n38552), .Z(n6721) );
  NANDN U7904 ( .A(n6719), .B(n38553), .Z(n6720) );
  NAND U7905 ( .A(n6721), .B(n6720), .Z(n6844) );
  OR U7906 ( .A(n6722), .B(n36105), .Z(n6724) );
  XNOR U7907 ( .A(b[3]), .B(a[53]), .Z(n6835) );
  NANDN U7908 ( .A(n6835), .B(n36107), .Z(n6723) );
  AND U7909 ( .A(n6724), .B(n6723), .Z(n6845) );
  XNOR U7910 ( .A(n6844), .B(n6845), .Z(n6846) );
  XOR U7911 ( .A(n6847), .B(n6846), .Z(n6874) );
  XNOR U7912 ( .A(n6875), .B(n6874), .Z(n6876) );
  XNOR U7913 ( .A(n6877), .B(n6876), .Z(n6923) );
  XNOR U7914 ( .A(n6922), .B(n6923), .Z(n6924) );
  XNOR U7915 ( .A(n6925), .B(n6924), .Z(n6943) );
  OR U7916 ( .A(n6726), .B(n6725), .Z(n6730) );
  NAND U7917 ( .A(n6728), .B(n6727), .Z(n6729) );
  NAND U7918 ( .A(n6730), .B(n6729), .Z(n6941) );
  NANDN U7919 ( .A(n6732), .B(n6731), .Z(n6736) );
  NANDN U7920 ( .A(n6734), .B(n6733), .Z(n6735) );
  NAND U7921 ( .A(n6736), .B(n6735), .Z(n6931) );
  OR U7922 ( .A(n6738), .B(n6737), .Z(n6742) );
  NAND U7923 ( .A(n6740), .B(n6739), .Z(n6741) );
  NAND U7924 ( .A(n6742), .B(n6741), .Z(n6928) );
  XNOR U7925 ( .A(b[9]), .B(a[47]), .Z(n6892) );
  NANDN U7926 ( .A(n6892), .B(n36925), .Z(n6745) );
  NANDN U7927 ( .A(n6743), .B(n36926), .Z(n6744) );
  NAND U7928 ( .A(n6745), .B(n6744), .Z(n6852) );
  XNOR U7929 ( .A(b[15]), .B(a[41]), .Z(n6895) );
  OR U7930 ( .A(n6895), .B(n37665), .Z(n6748) );
  NANDN U7931 ( .A(n6746), .B(n37604), .Z(n6747) );
  AND U7932 ( .A(n6748), .B(n6747), .Z(n6850) );
  XNOR U7933 ( .A(b[21]), .B(a[35]), .Z(n6898) );
  NANDN U7934 ( .A(n6898), .B(n38101), .Z(n6751) );
  NANDN U7935 ( .A(n6749), .B(n38102), .Z(n6750) );
  AND U7936 ( .A(n6751), .B(n6750), .Z(n6851) );
  XOR U7937 ( .A(n6852), .B(n6853), .Z(n6841) );
  XNOR U7938 ( .A(b[11]), .B(a[45]), .Z(n6901) );
  OR U7939 ( .A(n6901), .B(n37311), .Z(n6754) );
  NANDN U7940 ( .A(n6752), .B(n37218), .Z(n6753) );
  NAND U7941 ( .A(n6754), .B(n6753), .Z(n6839) );
  XOR U7942 ( .A(n1053), .B(a[43]), .Z(n6904) );
  NANDN U7943 ( .A(n6904), .B(n37424), .Z(n6757) );
  NANDN U7944 ( .A(n6755), .B(n37425), .Z(n6756) );
  AND U7945 ( .A(n6757), .B(n6756), .Z(n6838) );
  XNOR U7946 ( .A(n6839), .B(n6838), .Z(n6840) );
  XOR U7947 ( .A(n6841), .B(n6840), .Z(n6859) );
  NANDN U7948 ( .A(n1049), .B(a[55]), .Z(n6758) );
  XNOR U7949 ( .A(b[1]), .B(n6758), .Z(n6760) );
  IV U7950 ( .A(a[54]), .Z(n11319) );
  NANDN U7951 ( .A(n11319), .B(n1049), .Z(n6759) );
  AND U7952 ( .A(n6760), .B(n6759), .Z(n6816) );
  NAND U7953 ( .A(n38490), .B(n6761), .Z(n6763) );
  XNOR U7954 ( .A(n1058), .B(a[27]), .Z(n6910) );
  NANDN U7955 ( .A(n1048), .B(n6910), .Z(n6762) );
  NAND U7956 ( .A(n6763), .B(n6762), .Z(n6814) );
  NANDN U7957 ( .A(n1059), .B(a[23]), .Z(n6815) );
  XNOR U7958 ( .A(n6814), .B(n6815), .Z(n6817) );
  XOR U7959 ( .A(n6816), .B(n6817), .Z(n6856) );
  NANDN U7960 ( .A(n6764), .B(n38205), .Z(n6766) );
  XNOR U7961 ( .A(b[23]), .B(a[33]), .Z(n6913) );
  OR U7962 ( .A(n6913), .B(n38268), .Z(n6765) );
  NAND U7963 ( .A(n6766), .B(n6765), .Z(n6883) );
  XOR U7964 ( .A(b[7]), .B(a[49]), .Z(n6916) );
  NAND U7965 ( .A(n6916), .B(n36701), .Z(n6769) );
  NAND U7966 ( .A(n6767), .B(n36702), .Z(n6768) );
  NAND U7967 ( .A(n6769), .B(n6768), .Z(n6880) );
  XNOR U7968 ( .A(b[25]), .B(a[31]), .Z(n6919) );
  NANDN U7969 ( .A(n6919), .B(n38325), .Z(n6772) );
  NANDN U7970 ( .A(n6770), .B(n38326), .Z(n6771) );
  AND U7971 ( .A(n6772), .B(n6771), .Z(n6881) );
  XNOR U7972 ( .A(n6880), .B(n6881), .Z(n6882) );
  XNOR U7973 ( .A(n6883), .B(n6882), .Z(n6857) );
  XNOR U7974 ( .A(n6856), .B(n6857), .Z(n6858) );
  XNOR U7975 ( .A(n6859), .B(n6858), .Z(n6871) );
  NANDN U7976 ( .A(n6774), .B(n6773), .Z(n6778) );
  NAND U7977 ( .A(n6776), .B(n6775), .Z(n6777) );
  NAND U7978 ( .A(n6778), .B(n6777), .Z(n6869) );
  NANDN U7979 ( .A(n6780), .B(n6779), .Z(n6784) );
  NAND U7980 ( .A(n6782), .B(n6781), .Z(n6783) );
  AND U7981 ( .A(n6784), .B(n6783), .Z(n6868) );
  XNOR U7982 ( .A(n6869), .B(n6868), .Z(n6870) );
  XNOR U7983 ( .A(n6871), .B(n6870), .Z(n6929) );
  XNOR U7984 ( .A(n6928), .B(n6929), .Z(n6930) );
  XOR U7985 ( .A(n6931), .B(n6930), .Z(n6940) );
  XNOR U7986 ( .A(n6941), .B(n6940), .Z(n6942) );
  XOR U7987 ( .A(n6943), .B(n6942), .Z(n6937) );
  NANDN U7988 ( .A(n6786), .B(n6785), .Z(n6790) );
  OR U7989 ( .A(n6788), .B(n6787), .Z(n6789) );
  NAND U7990 ( .A(n6790), .B(n6789), .Z(n6934) );
  NAND U7991 ( .A(n6792), .B(n6791), .Z(n6796) );
  NANDN U7992 ( .A(n6794), .B(n6793), .Z(n6795) );
  NAND U7993 ( .A(n6796), .B(n6795), .Z(n6935) );
  XNOR U7994 ( .A(n6934), .B(n6935), .Z(n6936) );
  XOR U7995 ( .A(n6937), .B(n6936), .Z(n6811) );
  XOR U7996 ( .A(n6810), .B(n6811), .Z(n6802) );
  XOR U7997 ( .A(n6803), .B(n6802), .Z(n6804) );
  XNOR U7998 ( .A(n6805), .B(n6804), .Z(n6946) );
  XNOR U7999 ( .A(n6946), .B(sreg[279]), .Z(n6948) );
  NAND U8000 ( .A(n6797), .B(sreg[278]), .Z(n6801) );
  OR U8001 ( .A(n6799), .B(n6798), .Z(n6800) );
  AND U8002 ( .A(n6801), .B(n6800), .Z(n6947) );
  XOR U8003 ( .A(n6948), .B(n6947), .Z(c[279]) );
  NAND U8004 ( .A(n6803), .B(n6802), .Z(n6807) );
  NAND U8005 ( .A(n6805), .B(n6804), .Z(n6806) );
  NAND U8006 ( .A(n6807), .B(n6806), .Z(n6954) );
  NANDN U8007 ( .A(n6809), .B(n6808), .Z(n6813) );
  NAND U8008 ( .A(n6811), .B(n6810), .Z(n6812) );
  NAND U8009 ( .A(n6813), .B(n6812), .Z(n6952) );
  NANDN U8010 ( .A(n6815), .B(n6814), .Z(n6819) );
  NAND U8011 ( .A(n6817), .B(n6816), .Z(n6818) );
  NAND U8012 ( .A(n6819), .B(n6818), .Z(n7038) );
  XNOR U8013 ( .A(b[19]), .B(a[38]), .Z(n6981) );
  NANDN U8014 ( .A(n6981), .B(n37934), .Z(n6822) );
  NANDN U8015 ( .A(n6820), .B(n37935), .Z(n6821) );
  NAND U8016 ( .A(n6822), .B(n6821), .Z(n7048) );
  XNOR U8017 ( .A(b[27]), .B(a[30]), .Z(n6984) );
  NANDN U8018 ( .A(n6984), .B(n38423), .Z(n6825) );
  NAND U8019 ( .A(n6823), .B(n38424), .Z(n6824) );
  NAND U8020 ( .A(n6825), .B(n6824), .Z(n7045) );
  XNOR U8021 ( .A(b[5]), .B(a[52]), .Z(n6987) );
  NANDN U8022 ( .A(n6987), .B(n36587), .Z(n6828) );
  NANDN U8023 ( .A(n6826), .B(n36588), .Z(n6827) );
  AND U8024 ( .A(n6828), .B(n6827), .Z(n7046) );
  XNOR U8025 ( .A(n7045), .B(n7046), .Z(n7047) );
  XNOR U8026 ( .A(n7048), .B(n7047), .Z(n7036) );
  NAND U8027 ( .A(n6829), .B(n37762), .Z(n6831) );
  XOR U8028 ( .A(b[17]), .B(a[40]), .Z(n6990) );
  NAND U8029 ( .A(n6990), .B(n37764), .Z(n6830) );
  NAND U8030 ( .A(n6831), .B(n6830), .Z(n7008) );
  XOR U8031 ( .A(b[31]), .B(n7202), .Z(n6993) );
  NANDN U8032 ( .A(n6993), .B(n38552), .Z(n6834) );
  NANDN U8033 ( .A(n6832), .B(n38553), .Z(n6833) );
  NAND U8034 ( .A(n6834), .B(n6833), .Z(n7005) );
  OR U8035 ( .A(n6835), .B(n36105), .Z(n6837) );
  XOR U8036 ( .A(b[3]), .B(n11319), .Z(n6996) );
  NANDN U8037 ( .A(n6996), .B(n36107), .Z(n6836) );
  AND U8038 ( .A(n6837), .B(n6836), .Z(n7006) );
  XNOR U8039 ( .A(n7005), .B(n7006), .Z(n7007) );
  XOR U8040 ( .A(n7008), .B(n7007), .Z(n7035) );
  XNOR U8041 ( .A(n7036), .B(n7035), .Z(n7037) );
  XNOR U8042 ( .A(n7038), .B(n7037), .Z(n7082) );
  NANDN U8043 ( .A(n6839), .B(n6838), .Z(n6843) );
  NAND U8044 ( .A(n6841), .B(n6840), .Z(n6842) );
  NAND U8045 ( .A(n6843), .B(n6842), .Z(n7026) );
  NANDN U8046 ( .A(n6845), .B(n6844), .Z(n6849) );
  NAND U8047 ( .A(n6847), .B(n6846), .Z(n6848) );
  NAND U8048 ( .A(n6849), .B(n6848), .Z(n7024) );
  OR U8049 ( .A(n6851), .B(n6850), .Z(n6855) );
  NANDN U8050 ( .A(n6853), .B(n6852), .Z(n6854) );
  NAND U8051 ( .A(n6855), .B(n6854), .Z(n7023) );
  XNOR U8052 ( .A(n7026), .B(n7025), .Z(n7083) );
  XOR U8053 ( .A(n7082), .B(n7083), .Z(n7085) );
  NANDN U8054 ( .A(n6857), .B(n6856), .Z(n6861) );
  NANDN U8055 ( .A(n6859), .B(n6858), .Z(n6860) );
  NAND U8056 ( .A(n6861), .B(n6860), .Z(n7084) );
  XOR U8057 ( .A(n7085), .B(n7084), .Z(n6971) );
  OR U8058 ( .A(n6863), .B(n6862), .Z(n6867) );
  NANDN U8059 ( .A(n6865), .B(n6864), .Z(n6866) );
  NAND U8060 ( .A(n6867), .B(n6866), .Z(n6970) );
  NANDN U8061 ( .A(n6869), .B(n6868), .Z(n6873) );
  NANDN U8062 ( .A(n6871), .B(n6870), .Z(n6872) );
  NAND U8063 ( .A(n6873), .B(n6872), .Z(n7090) );
  NANDN U8064 ( .A(n6875), .B(n6874), .Z(n6879) );
  NAND U8065 ( .A(n6877), .B(n6876), .Z(n6878) );
  NAND U8066 ( .A(n6879), .B(n6878), .Z(n7089) );
  NANDN U8067 ( .A(n6881), .B(n6880), .Z(n6885) );
  NAND U8068 ( .A(n6883), .B(n6882), .Z(n6884) );
  NAND U8069 ( .A(n6885), .B(n6884), .Z(n7029) );
  NANDN U8070 ( .A(n6887), .B(n6886), .Z(n6891) );
  NAND U8071 ( .A(n6889), .B(n6888), .Z(n6890) );
  AND U8072 ( .A(n6891), .B(n6890), .Z(n7030) );
  XNOR U8073 ( .A(n7029), .B(n7030), .Z(n7031) );
  XNOR U8074 ( .A(b[9]), .B(a[48]), .Z(n7051) );
  NANDN U8075 ( .A(n7051), .B(n36925), .Z(n6894) );
  NANDN U8076 ( .A(n6892), .B(n36926), .Z(n6893) );
  NAND U8077 ( .A(n6894), .B(n6893), .Z(n7013) );
  XNOR U8078 ( .A(b[15]), .B(a[42]), .Z(n7054) );
  OR U8079 ( .A(n7054), .B(n37665), .Z(n6897) );
  NANDN U8080 ( .A(n6895), .B(n37604), .Z(n6896) );
  AND U8081 ( .A(n6897), .B(n6896), .Z(n7011) );
  XNOR U8082 ( .A(b[21]), .B(a[36]), .Z(n7057) );
  NANDN U8083 ( .A(n7057), .B(n38101), .Z(n6900) );
  NANDN U8084 ( .A(n6898), .B(n38102), .Z(n6899) );
  AND U8085 ( .A(n6900), .B(n6899), .Z(n7012) );
  XOR U8086 ( .A(n7013), .B(n7014), .Z(n7002) );
  XNOR U8087 ( .A(b[11]), .B(a[46]), .Z(n7060) );
  OR U8088 ( .A(n7060), .B(n37311), .Z(n6903) );
  NANDN U8089 ( .A(n6901), .B(n37218), .Z(n6902) );
  NAND U8090 ( .A(n6903), .B(n6902), .Z(n7000) );
  XOR U8091 ( .A(n1053), .B(a[44]), .Z(n7063) );
  NANDN U8092 ( .A(n7063), .B(n37424), .Z(n6906) );
  NANDN U8093 ( .A(n6904), .B(n37425), .Z(n6905) );
  AND U8094 ( .A(n6906), .B(n6905), .Z(n6999) );
  XNOR U8095 ( .A(n7000), .B(n6999), .Z(n7001) );
  XOR U8096 ( .A(n7002), .B(n7001), .Z(n7019) );
  NANDN U8097 ( .A(n1049), .B(a[56]), .Z(n6907) );
  XNOR U8098 ( .A(b[1]), .B(n6907), .Z(n6909) );
  NANDN U8099 ( .A(b[0]), .B(a[55]), .Z(n6908) );
  AND U8100 ( .A(n6909), .B(n6908), .Z(n6977) );
  NAND U8101 ( .A(n38490), .B(n6910), .Z(n6912) );
  XNOR U8102 ( .A(b[29]), .B(a[28]), .Z(n7070) );
  OR U8103 ( .A(n7070), .B(n1048), .Z(n6911) );
  NAND U8104 ( .A(n6912), .B(n6911), .Z(n6975) );
  NANDN U8105 ( .A(n1059), .B(a[24]), .Z(n6976) );
  XNOR U8106 ( .A(n6975), .B(n6976), .Z(n6978) );
  XOR U8107 ( .A(n6977), .B(n6978), .Z(n7017) );
  NANDN U8108 ( .A(n6913), .B(n38205), .Z(n6915) );
  XNOR U8109 ( .A(b[23]), .B(a[34]), .Z(n7073) );
  OR U8110 ( .A(n7073), .B(n38268), .Z(n6914) );
  NAND U8111 ( .A(n6915), .B(n6914), .Z(n7042) );
  XNOR U8112 ( .A(b[7]), .B(a[50]), .Z(n7076) );
  NANDN U8113 ( .A(n7076), .B(n36701), .Z(n6918) );
  NAND U8114 ( .A(n6916), .B(n36702), .Z(n6917) );
  NAND U8115 ( .A(n6918), .B(n6917), .Z(n7039) );
  XOR U8116 ( .A(b[25]), .B(a[32]), .Z(n7079) );
  NAND U8117 ( .A(n7079), .B(n38325), .Z(n6921) );
  NANDN U8118 ( .A(n6919), .B(n38326), .Z(n6920) );
  AND U8119 ( .A(n6921), .B(n6920), .Z(n7040) );
  XNOR U8120 ( .A(n7039), .B(n7040), .Z(n7041) );
  XNOR U8121 ( .A(n7042), .B(n7041), .Z(n7018) );
  XOR U8122 ( .A(n7017), .B(n7018), .Z(n7020) );
  XNOR U8123 ( .A(n7019), .B(n7020), .Z(n7032) );
  XNOR U8124 ( .A(n7031), .B(n7032), .Z(n7088) );
  XNOR U8125 ( .A(n7089), .B(n7088), .Z(n7091) );
  XOR U8126 ( .A(n7090), .B(n7091), .Z(n6969) );
  XOR U8127 ( .A(n6970), .B(n6969), .Z(n6972) );
  NANDN U8128 ( .A(n6923), .B(n6922), .Z(n6927) );
  NAND U8129 ( .A(n6925), .B(n6924), .Z(n6926) );
  NAND U8130 ( .A(n6927), .B(n6926), .Z(n6964) );
  NANDN U8131 ( .A(n6929), .B(n6928), .Z(n6933) );
  NAND U8132 ( .A(n6931), .B(n6930), .Z(n6932) );
  AND U8133 ( .A(n6933), .B(n6932), .Z(n6963) );
  XNOR U8134 ( .A(n6964), .B(n6963), .Z(n6965) );
  XOR U8135 ( .A(n6966), .B(n6965), .Z(n6959) );
  NANDN U8136 ( .A(n6935), .B(n6934), .Z(n6939) );
  NAND U8137 ( .A(n6937), .B(n6936), .Z(n6938) );
  NAND U8138 ( .A(n6939), .B(n6938), .Z(n6957) );
  NANDN U8139 ( .A(n6941), .B(n6940), .Z(n6945) );
  NANDN U8140 ( .A(n6943), .B(n6942), .Z(n6944) );
  NAND U8141 ( .A(n6945), .B(n6944), .Z(n6958) );
  XNOR U8142 ( .A(n6957), .B(n6958), .Z(n6960) );
  XOR U8143 ( .A(n6959), .B(n6960), .Z(n6951) );
  XOR U8144 ( .A(n6952), .B(n6951), .Z(n6953) );
  XNOR U8145 ( .A(n6954), .B(n6953), .Z(n7092) );
  XNOR U8146 ( .A(n7092), .B(sreg[280]), .Z(n7094) );
  NAND U8147 ( .A(n6946), .B(sreg[279]), .Z(n6950) );
  OR U8148 ( .A(n6948), .B(n6947), .Z(n6949) );
  AND U8149 ( .A(n6950), .B(n6949), .Z(n7093) );
  XOR U8150 ( .A(n7094), .B(n7093), .Z(c[280]) );
  NAND U8151 ( .A(n6952), .B(n6951), .Z(n6956) );
  NAND U8152 ( .A(n6954), .B(n6953), .Z(n6955) );
  NAND U8153 ( .A(n6956), .B(n6955), .Z(n7100) );
  NANDN U8154 ( .A(n6958), .B(n6957), .Z(n6962) );
  NAND U8155 ( .A(n6960), .B(n6959), .Z(n6961) );
  NAND U8156 ( .A(n6962), .B(n6961), .Z(n7098) );
  NANDN U8157 ( .A(n6964), .B(n6963), .Z(n6968) );
  NAND U8158 ( .A(n6966), .B(n6965), .Z(n6967) );
  NAND U8159 ( .A(n6968), .B(n6967), .Z(n7103) );
  NANDN U8160 ( .A(n6970), .B(n6969), .Z(n6974) );
  OR U8161 ( .A(n6972), .B(n6971), .Z(n6973) );
  NAND U8162 ( .A(n6974), .B(n6973), .Z(n7104) );
  XNOR U8163 ( .A(n7103), .B(n7104), .Z(n7105) );
  NANDN U8164 ( .A(n6976), .B(n6975), .Z(n6980) );
  NAND U8165 ( .A(n6978), .B(n6977), .Z(n6979) );
  NAND U8166 ( .A(n6980), .B(n6979), .Z(n7172) );
  XNOR U8167 ( .A(b[19]), .B(a[39]), .Z(n7139) );
  NANDN U8168 ( .A(n7139), .B(n37934), .Z(n6983) );
  NANDN U8169 ( .A(n6981), .B(n37935), .Z(n6982) );
  NAND U8170 ( .A(n6983), .B(n6982), .Z(n7184) );
  XNOR U8171 ( .A(b[27]), .B(a[31]), .Z(n7142) );
  NANDN U8172 ( .A(n7142), .B(n38423), .Z(n6986) );
  NANDN U8173 ( .A(n6984), .B(n38424), .Z(n6985) );
  NAND U8174 ( .A(n6986), .B(n6985), .Z(n7181) );
  XNOR U8175 ( .A(b[5]), .B(a[53]), .Z(n7145) );
  NANDN U8176 ( .A(n7145), .B(n36587), .Z(n6989) );
  NANDN U8177 ( .A(n6987), .B(n36588), .Z(n6988) );
  AND U8178 ( .A(n6989), .B(n6988), .Z(n7182) );
  XNOR U8179 ( .A(n7181), .B(n7182), .Z(n7183) );
  XNOR U8180 ( .A(n7184), .B(n7183), .Z(n7169) );
  NAND U8181 ( .A(n6990), .B(n37762), .Z(n6992) );
  XOR U8182 ( .A(b[17]), .B(a[41]), .Z(n7148) );
  NAND U8183 ( .A(n7148), .B(n37764), .Z(n6991) );
  NAND U8184 ( .A(n6992), .B(n6991), .Z(n7123) );
  XNOR U8185 ( .A(b[31]), .B(a[27]), .Z(n7151) );
  NANDN U8186 ( .A(n7151), .B(n38552), .Z(n6995) );
  NANDN U8187 ( .A(n6993), .B(n38553), .Z(n6994) );
  AND U8188 ( .A(n6995), .B(n6994), .Z(n7121) );
  OR U8189 ( .A(n6996), .B(n36105), .Z(n6998) );
  XNOR U8190 ( .A(b[3]), .B(a[55]), .Z(n7154) );
  NANDN U8191 ( .A(n7154), .B(n36107), .Z(n6997) );
  AND U8192 ( .A(n6998), .B(n6997), .Z(n7122) );
  XOR U8193 ( .A(n7123), .B(n7124), .Z(n7170) );
  XOR U8194 ( .A(n7169), .B(n7170), .Z(n7171) );
  XNOR U8195 ( .A(n7172), .B(n7171), .Z(n7218) );
  NANDN U8196 ( .A(n7000), .B(n6999), .Z(n7004) );
  NAND U8197 ( .A(n7002), .B(n7001), .Z(n7003) );
  NAND U8198 ( .A(n7004), .B(n7003), .Z(n7160) );
  NANDN U8199 ( .A(n7006), .B(n7005), .Z(n7010) );
  NAND U8200 ( .A(n7008), .B(n7007), .Z(n7009) );
  NAND U8201 ( .A(n7010), .B(n7009), .Z(n7158) );
  OR U8202 ( .A(n7012), .B(n7011), .Z(n7016) );
  NANDN U8203 ( .A(n7014), .B(n7013), .Z(n7015) );
  NAND U8204 ( .A(n7016), .B(n7015), .Z(n7157) );
  XNOR U8205 ( .A(n7160), .B(n7159), .Z(n7219) );
  XOR U8206 ( .A(n7218), .B(n7219), .Z(n7221) );
  NANDN U8207 ( .A(n7018), .B(n7017), .Z(n7022) );
  OR U8208 ( .A(n7020), .B(n7019), .Z(n7021) );
  NAND U8209 ( .A(n7022), .B(n7021), .Z(n7220) );
  XOR U8210 ( .A(n7221), .B(n7220), .Z(n7238) );
  OR U8211 ( .A(n7024), .B(n7023), .Z(n7028) );
  NAND U8212 ( .A(n7026), .B(n7025), .Z(n7027) );
  NAND U8213 ( .A(n7028), .B(n7027), .Z(n7237) );
  NANDN U8214 ( .A(n7030), .B(n7029), .Z(n7034) );
  NANDN U8215 ( .A(n7032), .B(n7031), .Z(n7033) );
  NAND U8216 ( .A(n7034), .B(n7033), .Z(n7226) );
  NANDN U8217 ( .A(n7040), .B(n7039), .Z(n7044) );
  NAND U8218 ( .A(n7042), .B(n7041), .Z(n7043) );
  NAND U8219 ( .A(n7044), .B(n7043), .Z(n7163) );
  NANDN U8220 ( .A(n7046), .B(n7045), .Z(n7050) );
  NAND U8221 ( .A(n7048), .B(n7047), .Z(n7049) );
  AND U8222 ( .A(n7050), .B(n7049), .Z(n7164) );
  XNOR U8223 ( .A(n7163), .B(n7164), .Z(n7165) );
  XNOR U8224 ( .A(b[9]), .B(a[49]), .Z(n7187) );
  NANDN U8225 ( .A(n7187), .B(n36925), .Z(n7053) );
  NANDN U8226 ( .A(n7051), .B(n36926), .Z(n7052) );
  NAND U8227 ( .A(n7053), .B(n7052), .Z(n7129) );
  XNOR U8228 ( .A(b[15]), .B(a[43]), .Z(n7190) );
  OR U8229 ( .A(n7190), .B(n37665), .Z(n7056) );
  NANDN U8230 ( .A(n7054), .B(n37604), .Z(n7055) );
  AND U8231 ( .A(n7056), .B(n7055), .Z(n7127) );
  XOR U8232 ( .A(b[21]), .B(n8832), .Z(n7193) );
  NANDN U8233 ( .A(n7193), .B(n38101), .Z(n7059) );
  NANDN U8234 ( .A(n7057), .B(n38102), .Z(n7058) );
  AND U8235 ( .A(n7059), .B(n7058), .Z(n7128) );
  XOR U8236 ( .A(n7129), .B(n7130), .Z(n7118) );
  XNOR U8237 ( .A(b[11]), .B(a[47]), .Z(n7196) );
  OR U8238 ( .A(n7196), .B(n37311), .Z(n7062) );
  NANDN U8239 ( .A(n7060), .B(n37218), .Z(n7061) );
  NAND U8240 ( .A(n7062), .B(n7061), .Z(n7116) );
  XOR U8241 ( .A(n1053), .B(a[45]), .Z(n7199) );
  NANDN U8242 ( .A(n7199), .B(n37424), .Z(n7065) );
  NANDN U8243 ( .A(n7063), .B(n37425), .Z(n7064) );
  NAND U8244 ( .A(n7065), .B(n7064), .Z(n7115) );
  XOR U8245 ( .A(n7118), .B(n7117), .Z(n7112) );
  NANDN U8246 ( .A(n1049), .B(a[57]), .Z(n7066) );
  XNOR U8247 ( .A(b[1]), .B(n7066), .Z(n7068) );
  NANDN U8248 ( .A(b[0]), .B(a[56]), .Z(n7067) );
  AND U8249 ( .A(n7068), .B(n7067), .Z(n7136) );
  ANDN U8250 ( .B(b[31]), .A(n7069), .Z(n7133) );
  NANDN U8251 ( .A(n7070), .B(n38490), .Z(n7072) );
  XNOR U8252 ( .A(b[29]), .B(a[29]), .Z(n7203) );
  OR U8253 ( .A(n7203), .B(n1048), .Z(n7071) );
  NAND U8254 ( .A(n7072), .B(n7071), .Z(n7134) );
  XOR U8255 ( .A(n7133), .B(n7134), .Z(n7135) );
  XNOR U8256 ( .A(n7136), .B(n7135), .Z(n7109) );
  NANDN U8257 ( .A(n7073), .B(n38205), .Z(n7075) );
  XNOR U8258 ( .A(b[23]), .B(a[35]), .Z(n7209) );
  OR U8259 ( .A(n7209), .B(n38268), .Z(n7074) );
  NAND U8260 ( .A(n7075), .B(n7074), .Z(n7178) );
  XOR U8261 ( .A(b[7]), .B(a[51]), .Z(n7212) );
  NAND U8262 ( .A(n7212), .B(n36701), .Z(n7078) );
  NANDN U8263 ( .A(n7076), .B(n36702), .Z(n7077) );
  NAND U8264 ( .A(n7078), .B(n7077), .Z(n7175) );
  XOR U8265 ( .A(b[25]), .B(a[33]), .Z(n7215) );
  NAND U8266 ( .A(n7215), .B(n38325), .Z(n7081) );
  NAND U8267 ( .A(n7079), .B(n38326), .Z(n7080) );
  AND U8268 ( .A(n7081), .B(n7080), .Z(n7176) );
  XNOR U8269 ( .A(n7175), .B(n7176), .Z(n7177) );
  XNOR U8270 ( .A(n7178), .B(n7177), .Z(n7110) );
  XOR U8271 ( .A(n7112), .B(n7111), .Z(n7166) );
  XNOR U8272 ( .A(n7165), .B(n7166), .Z(n7224) );
  XNOR U8273 ( .A(n7225), .B(n7224), .Z(n7227) );
  XNOR U8274 ( .A(n7226), .B(n7227), .Z(n7236) );
  XOR U8275 ( .A(n7237), .B(n7236), .Z(n7239) );
  NANDN U8276 ( .A(n7083), .B(n7082), .Z(n7087) );
  OR U8277 ( .A(n7085), .B(n7084), .Z(n7086) );
  NAND U8278 ( .A(n7087), .B(n7086), .Z(n7230) );
  XNOR U8279 ( .A(n7230), .B(n7231), .Z(n7232) );
  XOR U8280 ( .A(n7233), .B(n7232), .Z(n7106) );
  XOR U8281 ( .A(n7105), .B(n7106), .Z(n7097) );
  XOR U8282 ( .A(n7098), .B(n7097), .Z(n7099) );
  XNOR U8283 ( .A(n7100), .B(n7099), .Z(n7242) );
  XNOR U8284 ( .A(n7242), .B(sreg[281]), .Z(n7244) );
  NAND U8285 ( .A(n7092), .B(sreg[280]), .Z(n7096) );
  OR U8286 ( .A(n7094), .B(n7093), .Z(n7095) );
  AND U8287 ( .A(n7096), .B(n7095), .Z(n7243) );
  XOR U8288 ( .A(n7244), .B(n7243), .Z(c[281]) );
  NAND U8289 ( .A(n7098), .B(n7097), .Z(n7102) );
  NAND U8290 ( .A(n7100), .B(n7099), .Z(n7101) );
  NAND U8291 ( .A(n7102), .B(n7101), .Z(n7250) );
  NANDN U8292 ( .A(n7104), .B(n7103), .Z(n7108) );
  NAND U8293 ( .A(n7106), .B(n7105), .Z(n7107) );
  NAND U8294 ( .A(n7108), .B(n7107), .Z(n7248) );
  OR U8295 ( .A(n7110), .B(n7109), .Z(n7114) );
  NANDN U8296 ( .A(n7112), .B(n7111), .Z(n7113) );
  NAND U8297 ( .A(n7114), .B(n7113), .Z(n7380) );
  OR U8298 ( .A(n7116), .B(n7115), .Z(n7120) );
  NAND U8299 ( .A(n7118), .B(n7117), .Z(n7119) );
  NAND U8300 ( .A(n7120), .B(n7119), .Z(n7319) );
  OR U8301 ( .A(n7122), .B(n7121), .Z(n7126) );
  NANDN U8302 ( .A(n7124), .B(n7123), .Z(n7125) );
  NAND U8303 ( .A(n7126), .B(n7125), .Z(n7318) );
  OR U8304 ( .A(n7128), .B(n7127), .Z(n7132) );
  NANDN U8305 ( .A(n7130), .B(n7129), .Z(n7131) );
  NAND U8306 ( .A(n7132), .B(n7131), .Z(n7317) );
  XOR U8307 ( .A(n7319), .B(n7320), .Z(n7378) );
  OR U8308 ( .A(n7134), .B(n7133), .Z(n7138) );
  NANDN U8309 ( .A(n7136), .B(n7135), .Z(n7137) );
  NAND U8310 ( .A(n7138), .B(n7137), .Z(n7332) );
  XNOR U8311 ( .A(b[19]), .B(a[40]), .Z(n7299) );
  NANDN U8312 ( .A(n7299), .B(n37934), .Z(n7141) );
  NANDN U8313 ( .A(n7139), .B(n37935), .Z(n7140) );
  NAND U8314 ( .A(n7141), .B(n7140), .Z(n7344) );
  XOR U8315 ( .A(b[27]), .B(a[32]), .Z(n7302) );
  NAND U8316 ( .A(n38423), .B(n7302), .Z(n7144) );
  NANDN U8317 ( .A(n7142), .B(n38424), .Z(n7143) );
  NAND U8318 ( .A(n7144), .B(n7143), .Z(n7341) );
  XOR U8319 ( .A(b[5]), .B(n11319), .Z(n7305) );
  NANDN U8320 ( .A(n7305), .B(n36587), .Z(n7147) );
  NANDN U8321 ( .A(n7145), .B(n36588), .Z(n7146) );
  AND U8322 ( .A(n7147), .B(n7146), .Z(n7342) );
  XNOR U8323 ( .A(n7341), .B(n7342), .Z(n7343) );
  XNOR U8324 ( .A(n7344), .B(n7343), .Z(n7329) );
  NAND U8325 ( .A(n7148), .B(n37762), .Z(n7150) );
  XOR U8326 ( .A(b[17]), .B(a[42]), .Z(n7308) );
  NAND U8327 ( .A(n7308), .B(n37764), .Z(n7149) );
  NAND U8328 ( .A(n7150), .B(n7149), .Z(n7283) );
  XNOR U8329 ( .A(b[31]), .B(a[28]), .Z(n7311) );
  NANDN U8330 ( .A(n7311), .B(n38552), .Z(n7153) );
  NANDN U8331 ( .A(n7151), .B(n38553), .Z(n7152) );
  AND U8332 ( .A(n7153), .B(n7152), .Z(n7281) );
  OR U8333 ( .A(n7154), .B(n36105), .Z(n7156) );
  XNOR U8334 ( .A(b[3]), .B(a[56]), .Z(n7314) );
  NANDN U8335 ( .A(n7314), .B(n36107), .Z(n7155) );
  AND U8336 ( .A(n7156), .B(n7155), .Z(n7282) );
  XOR U8337 ( .A(n7283), .B(n7284), .Z(n7330) );
  XOR U8338 ( .A(n7329), .B(n7330), .Z(n7331) );
  XNOR U8339 ( .A(n7332), .B(n7331), .Z(n7377) );
  XOR U8340 ( .A(n7378), .B(n7377), .Z(n7379) );
  XNOR U8341 ( .A(n7380), .B(n7379), .Z(n7266) );
  OR U8342 ( .A(n7158), .B(n7157), .Z(n7162) );
  NAND U8343 ( .A(n7160), .B(n7159), .Z(n7161) );
  NAND U8344 ( .A(n7162), .B(n7161), .Z(n7264) );
  NANDN U8345 ( .A(n7164), .B(n7163), .Z(n7168) );
  NANDN U8346 ( .A(n7166), .B(n7165), .Z(n7167) );
  NAND U8347 ( .A(n7168), .B(n7167), .Z(n7383) );
  OR U8348 ( .A(n7170), .B(n7169), .Z(n7174) );
  NAND U8349 ( .A(n7172), .B(n7171), .Z(n7173) );
  NAND U8350 ( .A(n7174), .B(n7173), .Z(n7382) );
  NANDN U8351 ( .A(n7176), .B(n7175), .Z(n7180) );
  NAND U8352 ( .A(n7178), .B(n7177), .Z(n7179) );
  NAND U8353 ( .A(n7180), .B(n7179), .Z(n7323) );
  NANDN U8354 ( .A(n7182), .B(n7181), .Z(n7186) );
  NAND U8355 ( .A(n7184), .B(n7183), .Z(n7185) );
  AND U8356 ( .A(n7186), .B(n7185), .Z(n7324) );
  XNOR U8357 ( .A(n7323), .B(n7324), .Z(n7325) );
  XOR U8358 ( .A(b[9]), .B(n10724), .Z(n7347) );
  NANDN U8359 ( .A(n7347), .B(n36925), .Z(n7189) );
  NANDN U8360 ( .A(n7187), .B(n36926), .Z(n7188) );
  NAND U8361 ( .A(n7189), .B(n7188), .Z(n7289) );
  XOR U8362 ( .A(b[15]), .B(n9873), .Z(n7350) );
  OR U8363 ( .A(n7350), .B(n37665), .Z(n7192) );
  NANDN U8364 ( .A(n7190), .B(n37604), .Z(n7191) );
  AND U8365 ( .A(n7192), .B(n7191), .Z(n7287) );
  XNOR U8366 ( .A(b[21]), .B(a[38]), .Z(n7353) );
  NANDN U8367 ( .A(n7353), .B(n38101), .Z(n7195) );
  NANDN U8368 ( .A(n7193), .B(n38102), .Z(n7194) );
  AND U8369 ( .A(n7195), .B(n7194), .Z(n7288) );
  XOR U8370 ( .A(n7289), .B(n7290), .Z(n7278) );
  XNOR U8371 ( .A(b[11]), .B(a[48]), .Z(n7356) );
  OR U8372 ( .A(n7356), .B(n37311), .Z(n7198) );
  NANDN U8373 ( .A(n7196), .B(n37218), .Z(n7197) );
  NAND U8374 ( .A(n7198), .B(n7197), .Z(n7276) );
  XOR U8375 ( .A(n1053), .B(a[46]), .Z(n7359) );
  NANDN U8376 ( .A(n7359), .B(n37424), .Z(n7201) );
  NANDN U8377 ( .A(n7199), .B(n37425), .Z(n7200) );
  NAND U8378 ( .A(n7201), .B(n7200), .Z(n7275) );
  XOR U8379 ( .A(n7278), .B(n7277), .Z(n7272) );
  ANDN U8380 ( .B(b[31]), .A(n7202), .Z(n7293) );
  NANDN U8381 ( .A(n7203), .B(n38490), .Z(n7205) );
  XNOR U8382 ( .A(n1058), .B(a[30]), .Z(n7365) );
  NANDN U8383 ( .A(n1048), .B(n7365), .Z(n7204) );
  NAND U8384 ( .A(n7205), .B(n7204), .Z(n7294) );
  XOR U8385 ( .A(n7293), .B(n7294), .Z(n7295) );
  NANDN U8386 ( .A(n1049), .B(a[58]), .Z(n7206) );
  XNOR U8387 ( .A(b[1]), .B(n7206), .Z(n7208) );
  NANDN U8388 ( .A(b[0]), .B(a[57]), .Z(n7207) );
  AND U8389 ( .A(n7208), .B(n7207), .Z(n7296) );
  XNOR U8390 ( .A(n7295), .B(n7296), .Z(n7269) );
  NANDN U8391 ( .A(n7209), .B(n38205), .Z(n7211) );
  XNOR U8392 ( .A(b[23]), .B(a[36]), .Z(n7368) );
  OR U8393 ( .A(n7368), .B(n38268), .Z(n7210) );
  NAND U8394 ( .A(n7211), .B(n7210), .Z(n7338) );
  XOR U8395 ( .A(b[7]), .B(a[52]), .Z(n7371) );
  NAND U8396 ( .A(n7371), .B(n36701), .Z(n7214) );
  NAND U8397 ( .A(n7212), .B(n36702), .Z(n7213) );
  NAND U8398 ( .A(n7214), .B(n7213), .Z(n7335) );
  XOR U8399 ( .A(b[25]), .B(a[34]), .Z(n7374) );
  NAND U8400 ( .A(n7374), .B(n38325), .Z(n7217) );
  NAND U8401 ( .A(n7215), .B(n38326), .Z(n7216) );
  AND U8402 ( .A(n7217), .B(n7216), .Z(n7336) );
  XNOR U8403 ( .A(n7335), .B(n7336), .Z(n7337) );
  XNOR U8404 ( .A(n7338), .B(n7337), .Z(n7270) );
  XOR U8405 ( .A(n7272), .B(n7271), .Z(n7326) );
  XNOR U8406 ( .A(n7325), .B(n7326), .Z(n7381) );
  XNOR U8407 ( .A(n7382), .B(n7381), .Z(n7384) );
  XNOR U8408 ( .A(n7383), .B(n7384), .Z(n7263) );
  XNOR U8409 ( .A(n7264), .B(n7263), .Z(n7265) );
  XOR U8410 ( .A(n7266), .B(n7265), .Z(n7260) );
  NANDN U8411 ( .A(n7219), .B(n7218), .Z(n7223) );
  OR U8412 ( .A(n7221), .B(n7220), .Z(n7222) );
  NAND U8413 ( .A(n7223), .B(n7222), .Z(n7257) );
  NAND U8414 ( .A(n7225), .B(n7224), .Z(n7229) );
  NANDN U8415 ( .A(n7227), .B(n7226), .Z(n7228) );
  NAND U8416 ( .A(n7229), .B(n7228), .Z(n7258) );
  XNOR U8417 ( .A(n7257), .B(n7258), .Z(n7259) );
  XNOR U8418 ( .A(n7260), .B(n7259), .Z(n7254) );
  NANDN U8419 ( .A(n7231), .B(n7230), .Z(n7235) );
  NAND U8420 ( .A(n7233), .B(n7232), .Z(n7234) );
  NAND U8421 ( .A(n7235), .B(n7234), .Z(n7251) );
  NANDN U8422 ( .A(n7237), .B(n7236), .Z(n7241) );
  OR U8423 ( .A(n7239), .B(n7238), .Z(n7240) );
  NAND U8424 ( .A(n7241), .B(n7240), .Z(n7252) );
  XNOR U8425 ( .A(n7251), .B(n7252), .Z(n7253) );
  XNOR U8426 ( .A(n7254), .B(n7253), .Z(n7247) );
  XOR U8427 ( .A(n7248), .B(n7247), .Z(n7249) );
  XNOR U8428 ( .A(n7250), .B(n7249), .Z(n7387) );
  XNOR U8429 ( .A(n7387), .B(sreg[282]), .Z(n7389) );
  NAND U8430 ( .A(n7242), .B(sreg[281]), .Z(n7246) );
  OR U8431 ( .A(n7244), .B(n7243), .Z(n7245) );
  AND U8432 ( .A(n7246), .B(n7245), .Z(n7388) );
  XOR U8433 ( .A(n7389), .B(n7388), .Z(c[282]) );
  NANDN U8434 ( .A(n7252), .B(n7251), .Z(n7256) );
  NANDN U8435 ( .A(n7254), .B(n7253), .Z(n7255) );
  NAND U8436 ( .A(n7256), .B(n7255), .Z(n7393) );
  NANDN U8437 ( .A(n7258), .B(n7257), .Z(n7262) );
  NAND U8438 ( .A(n7260), .B(n7259), .Z(n7261) );
  NAND U8439 ( .A(n7262), .B(n7261), .Z(n7398) );
  NANDN U8440 ( .A(n7264), .B(n7263), .Z(n7268) );
  NANDN U8441 ( .A(n7266), .B(n7265), .Z(n7267) );
  NAND U8442 ( .A(n7268), .B(n7267), .Z(n7399) );
  XNOR U8443 ( .A(n7398), .B(n7399), .Z(n7400) );
  OR U8444 ( .A(n7270), .B(n7269), .Z(n7274) );
  NANDN U8445 ( .A(n7272), .B(n7271), .Z(n7273) );
  NAND U8446 ( .A(n7274), .B(n7273), .Z(n7528) );
  OR U8447 ( .A(n7276), .B(n7275), .Z(n7280) );
  NAND U8448 ( .A(n7278), .B(n7277), .Z(n7279) );
  NAND U8449 ( .A(n7280), .B(n7279), .Z(n7467) );
  OR U8450 ( .A(n7282), .B(n7281), .Z(n7286) );
  NANDN U8451 ( .A(n7284), .B(n7283), .Z(n7285) );
  NAND U8452 ( .A(n7286), .B(n7285), .Z(n7466) );
  OR U8453 ( .A(n7288), .B(n7287), .Z(n7292) );
  NANDN U8454 ( .A(n7290), .B(n7289), .Z(n7291) );
  NAND U8455 ( .A(n7292), .B(n7291), .Z(n7465) );
  XOR U8456 ( .A(n7467), .B(n7468), .Z(n7526) );
  OR U8457 ( .A(n7294), .B(n7293), .Z(n7298) );
  NANDN U8458 ( .A(n7296), .B(n7295), .Z(n7297) );
  NAND U8459 ( .A(n7298), .B(n7297), .Z(n7479) );
  XNOR U8460 ( .A(b[19]), .B(a[41]), .Z(n7422) );
  NANDN U8461 ( .A(n7422), .B(n37934), .Z(n7301) );
  NANDN U8462 ( .A(n7299), .B(n37935), .Z(n7300) );
  NAND U8463 ( .A(n7301), .B(n7300), .Z(n7492) );
  XOR U8464 ( .A(b[27]), .B(a[33]), .Z(n7425) );
  NAND U8465 ( .A(n38423), .B(n7425), .Z(n7304) );
  NAND U8466 ( .A(n7302), .B(n38424), .Z(n7303) );
  NAND U8467 ( .A(n7304), .B(n7303), .Z(n7489) );
  XNOR U8468 ( .A(b[5]), .B(a[55]), .Z(n7428) );
  NANDN U8469 ( .A(n7428), .B(n36587), .Z(n7307) );
  NANDN U8470 ( .A(n7305), .B(n36588), .Z(n7306) );
  AND U8471 ( .A(n7307), .B(n7306), .Z(n7490) );
  XNOR U8472 ( .A(n7489), .B(n7490), .Z(n7491) );
  XNOR U8473 ( .A(n7492), .B(n7491), .Z(n7478) );
  NAND U8474 ( .A(n7308), .B(n37762), .Z(n7310) );
  XOR U8475 ( .A(b[17]), .B(a[43]), .Z(n7431) );
  NAND U8476 ( .A(n7431), .B(n37764), .Z(n7309) );
  NAND U8477 ( .A(n7310), .B(n7309), .Z(n7450) );
  XNOR U8478 ( .A(b[31]), .B(a[29]), .Z(n7435) );
  NANDN U8479 ( .A(n7435), .B(n38552), .Z(n7313) );
  NANDN U8480 ( .A(n7311), .B(n38553), .Z(n7312) );
  NAND U8481 ( .A(n7313), .B(n7312), .Z(n7447) );
  OR U8482 ( .A(n7314), .B(n36105), .Z(n7316) );
  XNOR U8483 ( .A(b[3]), .B(a[57]), .Z(n7438) );
  NANDN U8484 ( .A(n7438), .B(n36107), .Z(n7315) );
  AND U8485 ( .A(n7316), .B(n7315), .Z(n7448) );
  XNOR U8486 ( .A(n7447), .B(n7448), .Z(n7449) );
  XOR U8487 ( .A(n7450), .B(n7449), .Z(n7477) );
  XOR U8488 ( .A(n7478), .B(n7477), .Z(n7480) );
  XOR U8489 ( .A(n7479), .B(n7480), .Z(n7525) );
  XOR U8490 ( .A(n7526), .B(n7525), .Z(n7527) );
  XNOR U8491 ( .A(n7528), .B(n7527), .Z(n7413) );
  OR U8492 ( .A(n7318), .B(n7317), .Z(n7322) );
  NANDN U8493 ( .A(n7320), .B(n7319), .Z(n7321) );
  NAND U8494 ( .A(n7322), .B(n7321), .Z(n7411) );
  NANDN U8495 ( .A(n7324), .B(n7323), .Z(n7328) );
  NANDN U8496 ( .A(n7326), .B(n7325), .Z(n7327) );
  NAND U8497 ( .A(n7328), .B(n7327), .Z(n7533) );
  OR U8498 ( .A(n7330), .B(n7329), .Z(n7334) );
  NANDN U8499 ( .A(n7332), .B(n7331), .Z(n7333) );
  NAND U8500 ( .A(n7334), .B(n7333), .Z(n7532) );
  NANDN U8501 ( .A(n7336), .B(n7335), .Z(n7340) );
  NAND U8502 ( .A(n7338), .B(n7337), .Z(n7339) );
  NAND U8503 ( .A(n7340), .B(n7339), .Z(n7471) );
  NANDN U8504 ( .A(n7342), .B(n7341), .Z(n7346) );
  NAND U8505 ( .A(n7344), .B(n7343), .Z(n7345) );
  AND U8506 ( .A(n7346), .B(n7345), .Z(n7472) );
  XNOR U8507 ( .A(n7471), .B(n7472), .Z(n7473) );
  XNOR U8508 ( .A(b[9]), .B(a[51]), .Z(n7495) );
  NANDN U8509 ( .A(n7495), .B(n36925), .Z(n7349) );
  NANDN U8510 ( .A(n7347), .B(n36926), .Z(n7348) );
  NAND U8511 ( .A(n7349), .B(n7348), .Z(n7455) );
  XNOR U8512 ( .A(b[15]), .B(a[45]), .Z(n7498) );
  OR U8513 ( .A(n7498), .B(n37665), .Z(n7352) );
  NANDN U8514 ( .A(n7350), .B(n37604), .Z(n7351) );
  AND U8515 ( .A(n7352), .B(n7351), .Z(n7453) );
  XNOR U8516 ( .A(b[21]), .B(a[39]), .Z(n7501) );
  NANDN U8517 ( .A(n7501), .B(n38101), .Z(n7355) );
  NANDN U8518 ( .A(n7353), .B(n38102), .Z(n7354) );
  AND U8519 ( .A(n7355), .B(n7354), .Z(n7454) );
  XOR U8520 ( .A(n7455), .B(n7456), .Z(n7444) );
  XNOR U8521 ( .A(b[11]), .B(a[49]), .Z(n7504) );
  OR U8522 ( .A(n7504), .B(n37311), .Z(n7358) );
  NANDN U8523 ( .A(n7356), .B(n37218), .Z(n7357) );
  NAND U8524 ( .A(n7358), .B(n7357), .Z(n7442) );
  XOR U8525 ( .A(n1053), .B(a[47]), .Z(n7507) );
  NANDN U8526 ( .A(n7507), .B(n37424), .Z(n7361) );
  NANDN U8527 ( .A(n7359), .B(n37425), .Z(n7360) );
  AND U8528 ( .A(n7361), .B(n7360), .Z(n7441) );
  XNOR U8529 ( .A(n7442), .B(n7441), .Z(n7443) );
  XOR U8530 ( .A(n7444), .B(n7443), .Z(n7461) );
  NANDN U8531 ( .A(n1049), .B(a[59]), .Z(n7362) );
  XNOR U8532 ( .A(b[1]), .B(n7362), .Z(n7364) );
  NANDN U8533 ( .A(b[0]), .B(a[58]), .Z(n7363) );
  AND U8534 ( .A(n7364), .B(n7363), .Z(n7418) );
  NAND U8535 ( .A(n7365), .B(n38490), .Z(n7367) );
  XOR U8536 ( .A(n1058), .B(n7955), .Z(n7513) );
  NANDN U8537 ( .A(n1048), .B(n7513), .Z(n7366) );
  NAND U8538 ( .A(n7367), .B(n7366), .Z(n7416) );
  NANDN U8539 ( .A(n1059), .B(a[27]), .Z(n7417) );
  XNOR U8540 ( .A(n7416), .B(n7417), .Z(n7419) );
  XOR U8541 ( .A(n7418), .B(n7419), .Z(n7459) );
  NANDN U8542 ( .A(n7368), .B(n38205), .Z(n7370) );
  XOR U8543 ( .A(b[23]), .B(n8832), .Z(n7516) );
  OR U8544 ( .A(n7516), .B(n38268), .Z(n7369) );
  NAND U8545 ( .A(n7370), .B(n7369), .Z(n7486) );
  XOR U8546 ( .A(b[7]), .B(a[53]), .Z(n7519) );
  NAND U8547 ( .A(n7519), .B(n36701), .Z(n7373) );
  NAND U8548 ( .A(n7371), .B(n36702), .Z(n7372) );
  NAND U8549 ( .A(n7373), .B(n7372), .Z(n7483) );
  XOR U8550 ( .A(b[25]), .B(a[35]), .Z(n7522) );
  NAND U8551 ( .A(n7522), .B(n38325), .Z(n7376) );
  NAND U8552 ( .A(n7374), .B(n38326), .Z(n7375) );
  AND U8553 ( .A(n7376), .B(n7375), .Z(n7484) );
  XNOR U8554 ( .A(n7483), .B(n7484), .Z(n7485) );
  XNOR U8555 ( .A(n7486), .B(n7485), .Z(n7460) );
  XOR U8556 ( .A(n7459), .B(n7460), .Z(n7462) );
  XNOR U8557 ( .A(n7461), .B(n7462), .Z(n7474) );
  XNOR U8558 ( .A(n7473), .B(n7474), .Z(n7531) );
  XNOR U8559 ( .A(n7532), .B(n7531), .Z(n7534) );
  XNOR U8560 ( .A(n7533), .B(n7534), .Z(n7410) );
  XNOR U8561 ( .A(n7411), .B(n7410), .Z(n7412) );
  XOR U8562 ( .A(n7413), .B(n7412), .Z(n7407) );
  NAND U8563 ( .A(n7382), .B(n7381), .Z(n7386) );
  NANDN U8564 ( .A(n7384), .B(n7383), .Z(n7385) );
  AND U8565 ( .A(n7386), .B(n7385), .Z(n7404) );
  XNOR U8566 ( .A(n7405), .B(n7404), .Z(n7406) );
  XOR U8567 ( .A(n7407), .B(n7406), .Z(n7401) );
  XOR U8568 ( .A(n7400), .B(n7401), .Z(n7392) );
  XOR U8569 ( .A(n7393), .B(n7392), .Z(n7394) );
  XNOR U8570 ( .A(n7395), .B(n7394), .Z(n7537) );
  XNOR U8571 ( .A(n7537), .B(sreg[283]), .Z(n7539) );
  NAND U8572 ( .A(n7387), .B(sreg[282]), .Z(n7391) );
  OR U8573 ( .A(n7389), .B(n7388), .Z(n7390) );
  AND U8574 ( .A(n7391), .B(n7390), .Z(n7538) );
  XOR U8575 ( .A(n7539), .B(n7538), .Z(c[283]) );
  NAND U8576 ( .A(n7393), .B(n7392), .Z(n7397) );
  NAND U8577 ( .A(n7395), .B(n7394), .Z(n7396) );
  NAND U8578 ( .A(n7397), .B(n7396), .Z(n7545) );
  NANDN U8579 ( .A(n7399), .B(n7398), .Z(n7403) );
  NAND U8580 ( .A(n7401), .B(n7400), .Z(n7402) );
  NAND U8581 ( .A(n7403), .B(n7402), .Z(n7543) );
  NANDN U8582 ( .A(n7405), .B(n7404), .Z(n7409) );
  NAND U8583 ( .A(n7407), .B(n7406), .Z(n7408) );
  NAND U8584 ( .A(n7409), .B(n7408), .Z(n7548) );
  NANDN U8585 ( .A(n7411), .B(n7410), .Z(n7415) );
  NANDN U8586 ( .A(n7413), .B(n7412), .Z(n7414) );
  NAND U8587 ( .A(n7415), .B(n7414), .Z(n7549) );
  XNOR U8588 ( .A(n7548), .B(n7549), .Z(n7550) );
  NANDN U8589 ( .A(n7417), .B(n7416), .Z(n7421) );
  NAND U8590 ( .A(n7419), .B(n7418), .Z(n7420) );
  NAND U8591 ( .A(n7421), .B(n7420), .Z(n7629) );
  XNOR U8592 ( .A(b[19]), .B(a[42]), .Z(n7572) );
  NANDN U8593 ( .A(n7572), .B(n37934), .Z(n7424) );
  NANDN U8594 ( .A(n7422), .B(n37935), .Z(n7423) );
  NAND U8595 ( .A(n7424), .B(n7423), .Z(n7639) );
  XOR U8596 ( .A(b[27]), .B(a[34]), .Z(n7575) );
  NAND U8597 ( .A(n38423), .B(n7575), .Z(n7427) );
  NAND U8598 ( .A(n7425), .B(n38424), .Z(n7426) );
  NAND U8599 ( .A(n7427), .B(n7426), .Z(n7636) );
  XNOR U8600 ( .A(b[5]), .B(a[56]), .Z(n7578) );
  NANDN U8601 ( .A(n7578), .B(n36587), .Z(n7430) );
  NANDN U8602 ( .A(n7428), .B(n36588), .Z(n7429) );
  AND U8603 ( .A(n7430), .B(n7429), .Z(n7637) );
  XNOR U8604 ( .A(n7636), .B(n7637), .Z(n7638) );
  XNOR U8605 ( .A(n7639), .B(n7638), .Z(n7627) );
  NAND U8606 ( .A(n7431), .B(n37762), .Z(n7433) );
  XNOR U8607 ( .A(b[17]), .B(a[44]), .Z(n7581) );
  NANDN U8608 ( .A(n7581), .B(n37764), .Z(n7432) );
  NAND U8609 ( .A(n7433), .B(n7432), .Z(n7599) );
  XOR U8610 ( .A(b[31]), .B(n7434), .Z(n7584) );
  NANDN U8611 ( .A(n7584), .B(n38552), .Z(n7437) );
  NANDN U8612 ( .A(n7435), .B(n38553), .Z(n7436) );
  NAND U8613 ( .A(n7437), .B(n7436), .Z(n7596) );
  OR U8614 ( .A(n7438), .B(n36105), .Z(n7440) );
  XNOR U8615 ( .A(b[3]), .B(a[58]), .Z(n7587) );
  NANDN U8616 ( .A(n7587), .B(n36107), .Z(n7439) );
  AND U8617 ( .A(n7440), .B(n7439), .Z(n7597) );
  XNOR U8618 ( .A(n7596), .B(n7597), .Z(n7598) );
  XOR U8619 ( .A(n7599), .B(n7598), .Z(n7626) );
  XNOR U8620 ( .A(n7627), .B(n7626), .Z(n7628) );
  XNOR U8621 ( .A(n7629), .B(n7628), .Z(n7672) );
  NANDN U8622 ( .A(n7442), .B(n7441), .Z(n7446) );
  NAND U8623 ( .A(n7444), .B(n7443), .Z(n7445) );
  NAND U8624 ( .A(n7446), .B(n7445), .Z(n7617) );
  NANDN U8625 ( .A(n7448), .B(n7447), .Z(n7452) );
  NAND U8626 ( .A(n7450), .B(n7449), .Z(n7451) );
  NAND U8627 ( .A(n7452), .B(n7451), .Z(n7615) );
  OR U8628 ( .A(n7454), .B(n7453), .Z(n7458) );
  NANDN U8629 ( .A(n7456), .B(n7455), .Z(n7457) );
  NAND U8630 ( .A(n7458), .B(n7457), .Z(n7614) );
  XNOR U8631 ( .A(n7617), .B(n7616), .Z(n7673) );
  XOR U8632 ( .A(n7672), .B(n7673), .Z(n7675) );
  NANDN U8633 ( .A(n7460), .B(n7459), .Z(n7464) );
  OR U8634 ( .A(n7462), .B(n7461), .Z(n7463) );
  NAND U8635 ( .A(n7464), .B(n7463), .Z(n7674) );
  XOR U8636 ( .A(n7675), .B(n7674), .Z(n7562) );
  OR U8637 ( .A(n7466), .B(n7465), .Z(n7470) );
  NANDN U8638 ( .A(n7468), .B(n7467), .Z(n7469) );
  NAND U8639 ( .A(n7470), .B(n7469), .Z(n7561) );
  NANDN U8640 ( .A(n7472), .B(n7471), .Z(n7476) );
  NANDN U8641 ( .A(n7474), .B(n7473), .Z(n7475) );
  NAND U8642 ( .A(n7476), .B(n7475), .Z(n7680) );
  NANDN U8643 ( .A(n7478), .B(n7477), .Z(n7482) );
  OR U8644 ( .A(n7480), .B(n7479), .Z(n7481) );
  NAND U8645 ( .A(n7482), .B(n7481), .Z(n7679) );
  NANDN U8646 ( .A(n7484), .B(n7483), .Z(n7488) );
  NAND U8647 ( .A(n7486), .B(n7485), .Z(n7487) );
  NAND U8648 ( .A(n7488), .B(n7487), .Z(n7620) );
  NANDN U8649 ( .A(n7490), .B(n7489), .Z(n7494) );
  NAND U8650 ( .A(n7492), .B(n7491), .Z(n7493) );
  AND U8651 ( .A(n7494), .B(n7493), .Z(n7621) );
  XNOR U8652 ( .A(n7620), .B(n7621), .Z(n7622) );
  XNOR U8653 ( .A(b[9]), .B(a[52]), .Z(n7642) );
  NANDN U8654 ( .A(n7642), .B(n36925), .Z(n7497) );
  NANDN U8655 ( .A(n7495), .B(n36926), .Z(n7496) );
  NAND U8656 ( .A(n7497), .B(n7496), .Z(n7604) );
  XNOR U8657 ( .A(b[15]), .B(a[46]), .Z(n7645) );
  OR U8658 ( .A(n7645), .B(n37665), .Z(n7500) );
  NANDN U8659 ( .A(n7498), .B(n37604), .Z(n7499) );
  AND U8660 ( .A(n7500), .B(n7499), .Z(n7602) );
  XNOR U8661 ( .A(b[21]), .B(a[40]), .Z(n7648) );
  NANDN U8662 ( .A(n7648), .B(n38101), .Z(n7503) );
  NANDN U8663 ( .A(n7501), .B(n38102), .Z(n7502) );
  AND U8664 ( .A(n7503), .B(n7502), .Z(n7603) );
  XOR U8665 ( .A(n7604), .B(n7605), .Z(n7593) );
  XOR U8666 ( .A(b[11]), .B(n10724), .Z(n7651) );
  OR U8667 ( .A(n7651), .B(n37311), .Z(n7506) );
  NANDN U8668 ( .A(n7504), .B(n37218), .Z(n7505) );
  NAND U8669 ( .A(n7506), .B(n7505), .Z(n7591) );
  XOR U8670 ( .A(n1053), .B(a[48]), .Z(n7654) );
  NANDN U8671 ( .A(n7654), .B(n37424), .Z(n7509) );
  NANDN U8672 ( .A(n7507), .B(n37425), .Z(n7508) );
  AND U8673 ( .A(n7509), .B(n7508), .Z(n7590) );
  XNOR U8674 ( .A(n7591), .B(n7590), .Z(n7592) );
  XOR U8675 ( .A(n7593), .B(n7592), .Z(n7610) );
  NANDN U8676 ( .A(n1049), .B(a[60]), .Z(n7510) );
  XNOR U8677 ( .A(b[1]), .B(n7510), .Z(n7512) );
  IV U8678 ( .A(a[59]), .Z(n12056) );
  NANDN U8679 ( .A(n12056), .B(n1049), .Z(n7511) );
  AND U8680 ( .A(n7512), .B(n7511), .Z(n7568) );
  NAND U8681 ( .A(n38490), .B(n7513), .Z(n7515) );
  XNOR U8682 ( .A(n1058), .B(a[32]), .Z(n7657) );
  NANDN U8683 ( .A(n1048), .B(n7657), .Z(n7514) );
  NAND U8684 ( .A(n7515), .B(n7514), .Z(n7566) );
  NANDN U8685 ( .A(n1059), .B(a[28]), .Z(n7567) );
  XNOR U8686 ( .A(n7566), .B(n7567), .Z(n7569) );
  XOR U8687 ( .A(n7568), .B(n7569), .Z(n7608) );
  NANDN U8688 ( .A(n7516), .B(n38205), .Z(n7518) );
  XNOR U8689 ( .A(b[23]), .B(a[38]), .Z(n7663) );
  OR U8690 ( .A(n7663), .B(n38268), .Z(n7517) );
  NAND U8691 ( .A(n7518), .B(n7517), .Z(n7633) );
  XNOR U8692 ( .A(b[7]), .B(a[54]), .Z(n7666) );
  NANDN U8693 ( .A(n7666), .B(n36701), .Z(n7521) );
  NAND U8694 ( .A(n7519), .B(n36702), .Z(n7520) );
  NAND U8695 ( .A(n7521), .B(n7520), .Z(n7630) );
  XOR U8696 ( .A(b[25]), .B(a[36]), .Z(n7669) );
  NAND U8697 ( .A(n7669), .B(n38325), .Z(n7524) );
  NAND U8698 ( .A(n7522), .B(n38326), .Z(n7523) );
  AND U8699 ( .A(n7524), .B(n7523), .Z(n7631) );
  XNOR U8700 ( .A(n7630), .B(n7631), .Z(n7632) );
  XNOR U8701 ( .A(n7633), .B(n7632), .Z(n7609) );
  XOR U8702 ( .A(n7608), .B(n7609), .Z(n7611) );
  XNOR U8703 ( .A(n7610), .B(n7611), .Z(n7623) );
  XNOR U8704 ( .A(n7622), .B(n7623), .Z(n7678) );
  XNOR U8705 ( .A(n7679), .B(n7678), .Z(n7681) );
  XNOR U8706 ( .A(n7680), .B(n7681), .Z(n7560) );
  XOR U8707 ( .A(n7561), .B(n7560), .Z(n7563) );
  NAND U8708 ( .A(n7526), .B(n7525), .Z(n7530) );
  NAND U8709 ( .A(n7528), .B(n7527), .Z(n7529) );
  NAND U8710 ( .A(n7530), .B(n7529), .Z(n7555) );
  NAND U8711 ( .A(n7532), .B(n7531), .Z(n7536) );
  NANDN U8712 ( .A(n7534), .B(n7533), .Z(n7535) );
  AND U8713 ( .A(n7536), .B(n7535), .Z(n7554) );
  XNOR U8714 ( .A(n7555), .B(n7554), .Z(n7556) );
  XOR U8715 ( .A(n7557), .B(n7556), .Z(n7551) );
  XOR U8716 ( .A(n7550), .B(n7551), .Z(n7542) );
  XOR U8717 ( .A(n7543), .B(n7542), .Z(n7544) );
  XNOR U8718 ( .A(n7545), .B(n7544), .Z(n7684) );
  XNOR U8719 ( .A(n7684), .B(sreg[284]), .Z(n7686) );
  NAND U8720 ( .A(n7537), .B(sreg[283]), .Z(n7541) );
  OR U8721 ( .A(n7539), .B(n7538), .Z(n7540) );
  AND U8722 ( .A(n7541), .B(n7540), .Z(n7685) );
  XOR U8723 ( .A(n7686), .B(n7685), .Z(c[284]) );
  NAND U8724 ( .A(n7543), .B(n7542), .Z(n7547) );
  NAND U8725 ( .A(n7545), .B(n7544), .Z(n7546) );
  NAND U8726 ( .A(n7547), .B(n7546), .Z(n7692) );
  NANDN U8727 ( .A(n7549), .B(n7548), .Z(n7553) );
  NAND U8728 ( .A(n7551), .B(n7550), .Z(n7552) );
  NAND U8729 ( .A(n7553), .B(n7552), .Z(n7690) );
  NANDN U8730 ( .A(n7555), .B(n7554), .Z(n7559) );
  NAND U8731 ( .A(n7557), .B(n7556), .Z(n7558) );
  NAND U8732 ( .A(n7559), .B(n7558), .Z(n7695) );
  NANDN U8733 ( .A(n7561), .B(n7560), .Z(n7565) );
  OR U8734 ( .A(n7563), .B(n7562), .Z(n7564) );
  NAND U8735 ( .A(n7565), .B(n7564), .Z(n7696) );
  XNOR U8736 ( .A(n7695), .B(n7696), .Z(n7697) );
  NANDN U8737 ( .A(n7567), .B(n7566), .Z(n7571) );
  NAND U8738 ( .A(n7569), .B(n7568), .Z(n7570) );
  NAND U8739 ( .A(n7571), .B(n7570), .Z(n7776) );
  XNOR U8740 ( .A(b[19]), .B(a[43]), .Z(n7743) );
  NANDN U8741 ( .A(n7743), .B(n37934), .Z(n7574) );
  NANDN U8742 ( .A(n7572), .B(n37935), .Z(n7573) );
  NAND U8743 ( .A(n7574), .B(n7573), .Z(n7788) );
  XOR U8744 ( .A(b[27]), .B(a[35]), .Z(n7746) );
  NAND U8745 ( .A(n38423), .B(n7746), .Z(n7577) );
  NAND U8746 ( .A(n7575), .B(n38424), .Z(n7576) );
  NAND U8747 ( .A(n7577), .B(n7576), .Z(n7785) );
  XNOR U8748 ( .A(b[5]), .B(a[57]), .Z(n7749) );
  NANDN U8749 ( .A(n7749), .B(n36587), .Z(n7580) );
  NANDN U8750 ( .A(n7578), .B(n36588), .Z(n7579) );
  AND U8751 ( .A(n7580), .B(n7579), .Z(n7786) );
  XNOR U8752 ( .A(n7785), .B(n7786), .Z(n7787) );
  XNOR U8753 ( .A(n7788), .B(n7787), .Z(n7773) );
  NANDN U8754 ( .A(n7581), .B(n37762), .Z(n7583) );
  XOR U8755 ( .A(b[17]), .B(a[45]), .Z(n7752) );
  NAND U8756 ( .A(n7752), .B(n37764), .Z(n7582) );
  NAND U8757 ( .A(n7583), .B(n7582), .Z(n7727) );
  XOR U8758 ( .A(b[31]), .B(n7955), .Z(n7755) );
  NANDN U8759 ( .A(n7755), .B(n38552), .Z(n7586) );
  NANDN U8760 ( .A(n7584), .B(n38553), .Z(n7585) );
  AND U8761 ( .A(n7586), .B(n7585), .Z(n7725) );
  OR U8762 ( .A(n7587), .B(n36105), .Z(n7589) );
  XOR U8763 ( .A(b[3]), .B(n12056), .Z(n7758) );
  NANDN U8764 ( .A(n7758), .B(n36107), .Z(n7588) );
  AND U8765 ( .A(n7589), .B(n7588), .Z(n7726) );
  XOR U8766 ( .A(n7727), .B(n7728), .Z(n7774) );
  XOR U8767 ( .A(n7773), .B(n7774), .Z(n7775) );
  XNOR U8768 ( .A(n7776), .B(n7775), .Z(n7821) );
  NANDN U8769 ( .A(n7591), .B(n7590), .Z(n7595) );
  NAND U8770 ( .A(n7593), .B(n7592), .Z(n7594) );
  NAND U8771 ( .A(n7595), .B(n7594), .Z(n7764) );
  NANDN U8772 ( .A(n7597), .B(n7596), .Z(n7601) );
  NAND U8773 ( .A(n7599), .B(n7598), .Z(n7600) );
  NAND U8774 ( .A(n7601), .B(n7600), .Z(n7762) );
  OR U8775 ( .A(n7603), .B(n7602), .Z(n7607) );
  NANDN U8776 ( .A(n7605), .B(n7604), .Z(n7606) );
  NAND U8777 ( .A(n7607), .B(n7606), .Z(n7761) );
  XNOR U8778 ( .A(n7764), .B(n7763), .Z(n7822) );
  XOR U8779 ( .A(n7821), .B(n7822), .Z(n7824) );
  NANDN U8780 ( .A(n7609), .B(n7608), .Z(n7613) );
  OR U8781 ( .A(n7611), .B(n7610), .Z(n7612) );
  NAND U8782 ( .A(n7613), .B(n7612), .Z(n7823) );
  XOR U8783 ( .A(n7824), .B(n7823), .Z(n7709) );
  OR U8784 ( .A(n7615), .B(n7614), .Z(n7619) );
  NAND U8785 ( .A(n7617), .B(n7616), .Z(n7618) );
  NAND U8786 ( .A(n7619), .B(n7618), .Z(n7708) );
  NANDN U8787 ( .A(n7621), .B(n7620), .Z(n7625) );
  NANDN U8788 ( .A(n7623), .B(n7622), .Z(n7624) );
  NAND U8789 ( .A(n7625), .B(n7624), .Z(n7829) );
  NANDN U8790 ( .A(n7631), .B(n7630), .Z(n7635) );
  NAND U8791 ( .A(n7633), .B(n7632), .Z(n7634) );
  NAND U8792 ( .A(n7635), .B(n7634), .Z(n7767) );
  NANDN U8793 ( .A(n7637), .B(n7636), .Z(n7641) );
  NAND U8794 ( .A(n7639), .B(n7638), .Z(n7640) );
  AND U8795 ( .A(n7641), .B(n7640), .Z(n7768) );
  XNOR U8796 ( .A(n7767), .B(n7768), .Z(n7769) );
  XNOR U8797 ( .A(b[9]), .B(a[53]), .Z(n7791) );
  NANDN U8798 ( .A(n7791), .B(n36925), .Z(n7644) );
  NANDN U8799 ( .A(n7642), .B(n36926), .Z(n7643) );
  NAND U8800 ( .A(n7644), .B(n7643), .Z(n7733) );
  XNOR U8801 ( .A(b[15]), .B(a[47]), .Z(n7794) );
  OR U8802 ( .A(n7794), .B(n37665), .Z(n7647) );
  NANDN U8803 ( .A(n7645), .B(n37604), .Z(n7646) );
  AND U8804 ( .A(n7647), .B(n7646), .Z(n7731) );
  XNOR U8805 ( .A(b[21]), .B(a[41]), .Z(n7797) );
  NANDN U8806 ( .A(n7797), .B(n38101), .Z(n7650) );
  NANDN U8807 ( .A(n7648), .B(n38102), .Z(n7649) );
  AND U8808 ( .A(n7650), .B(n7649), .Z(n7732) );
  XOR U8809 ( .A(n7733), .B(n7734), .Z(n7722) );
  XNOR U8810 ( .A(b[11]), .B(a[51]), .Z(n7800) );
  OR U8811 ( .A(n7800), .B(n37311), .Z(n7653) );
  NANDN U8812 ( .A(n7651), .B(n37218), .Z(n7652) );
  NAND U8813 ( .A(n7653), .B(n7652), .Z(n7720) );
  XOR U8814 ( .A(n1053), .B(a[49]), .Z(n7803) );
  NANDN U8815 ( .A(n7803), .B(n37424), .Z(n7656) );
  NANDN U8816 ( .A(n7654), .B(n37425), .Z(n7655) );
  NAND U8817 ( .A(n7656), .B(n7655), .Z(n7719) );
  XOR U8818 ( .A(n7722), .B(n7721), .Z(n7716) );
  NAND U8819 ( .A(n38490), .B(n7657), .Z(n7659) );
  XNOR U8820 ( .A(n1058), .B(a[33]), .Z(n7809) );
  NANDN U8821 ( .A(n1048), .B(n7809), .Z(n7658) );
  NAND U8822 ( .A(n7659), .B(n7658), .Z(n7737) );
  NANDN U8823 ( .A(n1059), .B(a[29]), .Z(n7738) );
  XNOR U8824 ( .A(n7737), .B(n7738), .Z(n7740) );
  NANDN U8825 ( .A(n1049), .B(a[61]), .Z(n7660) );
  XNOR U8826 ( .A(b[1]), .B(n7660), .Z(n7662) );
  NANDN U8827 ( .A(b[0]), .B(a[60]), .Z(n7661) );
  AND U8828 ( .A(n7662), .B(n7661), .Z(n7739) );
  XNOR U8829 ( .A(n7740), .B(n7739), .Z(n7714) );
  NANDN U8830 ( .A(n7663), .B(n38205), .Z(n7665) );
  XNOR U8831 ( .A(b[23]), .B(a[39]), .Z(n7812) );
  OR U8832 ( .A(n7812), .B(n38268), .Z(n7664) );
  NAND U8833 ( .A(n7665), .B(n7664), .Z(n7782) );
  XOR U8834 ( .A(b[7]), .B(a[55]), .Z(n7815) );
  NAND U8835 ( .A(n7815), .B(n36701), .Z(n7668) );
  NANDN U8836 ( .A(n7666), .B(n36702), .Z(n7667) );
  NAND U8837 ( .A(n7668), .B(n7667), .Z(n7779) );
  XNOR U8838 ( .A(b[25]), .B(a[37]), .Z(n7818) );
  NANDN U8839 ( .A(n7818), .B(n38325), .Z(n7671) );
  NAND U8840 ( .A(n7669), .B(n38326), .Z(n7670) );
  AND U8841 ( .A(n7671), .B(n7670), .Z(n7780) );
  XNOR U8842 ( .A(n7779), .B(n7780), .Z(n7781) );
  XOR U8843 ( .A(n7782), .B(n7781), .Z(n7713) );
  XOR U8844 ( .A(n7716), .B(n7715), .Z(n7770) );
  XNOR U8845 ( .A(n7769), .B(n7770), .Z(n7827) );
  XNOR U8846 ( .A(n7828), .B(n7827), .Z(n7830) );
  XNOR U8847 ( .A(n7829), .B(n7830), .Z(n7707) );
  XOR U8848 ( .A(n7708), .B(n7707), .Z(n7710) );
  NANDN U8849 ( .A(n7673), .B(n7672), .Z(n7677) );
  OR U8850 ( .A(n7675), .B(n7674), .Z(n7676) );
  NAND U8851 ( .A(n7677), .B(n7676), .Z(n7701) );
  NAND U8852 ( .A(n7679), .B(n7678), .Z(n7683) );
  NANDN U8853 ( .A(n7681), .B(n7680), .Z(n7682) );
  NAND U8854 ( .A(n7683), .B(n7682), .Z(n7702) );
  XNOR U8855 ( .A(n7701), .B(n7702), .Z(n7703) );
  XOR U8856 ( .A(n7704), .B(n7703), .Z(n7698) );
  XOR U8857 ( .A(n7697), .B(n7698), .Z(n7689) );
  XOR U8858 ( .A(n7690), .B(n7689), .Z(n7691) );
  XNOR U8859 ( .A(n7692), .B(n7691), .Z(n7833) );
  XNOR U8860 ( .A(n7833), .B(sreg[285]), .Z(n7835) );
  NAND U8861 ( .A(n7684), .B(sreg[284]), .Z(n7688) );
  OR U8862 ( .A(n7686), .B(n7685), .Z(n7687) );
  AND U8863 ( .A(n7688), .B(n7687), .Z(n7834) );
  XOR U8864 ( .A(n7835), .B(n7834), .Z(c[285]) );
  NAND U8865 ( .A(n7690), .B(n7689), .Z(n7694) );
  NAND U8866 ( .A(n7692), .B(n7691), .Z(n7693) );
  NAND U8867 ( .A(n7694), .B(n7693), .Z(n7841) );
  NANDN U8868 ( .A(n7696), .B(n7695), .Z(n7700) );
  NAND U8869 ( .A(n7698), .B(n7697), .Z(n7699) );
  NAND U8870 ( .A(n7700), .B(n7699), .Z(n7839) );
  NANDN U8871 ( .A(n7702), .B(n7701), .Z(n7706) );
  NAND U8872 ( .A(n7704), .B(n7703), .Z(n7705) );
  NAND U8873 ( .A(n7706), .B(n7705), .Z(n7844) );
  NANDN U8874 ( .A(n7708), .B(n7707), .Z(n7712) );
  OR U8875 ( .A(n7710), .B(n7709), .Z(n7711) );
  NAND U8876 ( .A(n7712), .B(n7711), .Z(n7845) );
  XNOR U8877 ( .A(n7844), .B(n7845), .Z(n7846) );
  NANDN U8878 ( .A(n7714), .B(n7713), .Z(n7718) );
  NANDN U8879 ( .A(n7716), .B(n7715), .Z(n7717) );
  NAND U8880 ( .A(n7718), .B(n7717), .Z(n7974) );
  OR U8881 ( .A(n7720), .B(n7719), .Z(n7724) );
  NAND U8882 ( .A(n7722), .B(n7721), .Z(n7723) );
  NAND U8883 ( .A(n7724), .B(n7723), .Z(n7912) );
  OR U8884 ( .A(n7726), .B(n7725), .Z(n7730) );
  NANDN U8885 ( .A(n7728), .B(n7727), .Z(n7729) );
  NAND U8886 ( .A(n7730), .B(n7729), .Z(n7911) );
  OR U8887 ( .A(n7732), .B(n7731), .Z(n7736) );
  NANDN U8888 ( .A(n7734), .B(n7733), .Z(n7735) );
  NAND U8889 ( .A(n7736), .B(n7735), .Z(n7910) );
  XOR U8890 ( .A(n7912), .B(n7913), .Z(n7971) );
  NANDN U8891 ( .A(n7738), .B(n7737), .Z(n7742) );
  NAND U8892 ( .A(n7740), .B(n7739), .Z(n7741) );
  NAND U8893 ( .A(n7742), .B(n7741), .Z(n7925) );
  XOR U8894 ( .A(b[19]), .B(n9873), .Z(n7868) );
  NANDN U8895 ( .A(n7868), .B(n37934), .Z(n7745) );
  NANDN U8896 ( .A(n7743), .B(n37935), .Z(n7744) );
  NAND U8897 ( .A(n7745), .B(n7744), .Z(n7937) );
  XOR U8898 ( .A(b[27]), .B(a[36]), .Z(n7871) );
  NAND U8899 ( .A(n38423), .B(n7871), .Z(n7748) );
  NAND U8900 ( .A(n7746), .B(n38424), .Z(n7747) );
  NAND U8901 ( .A(n7748), .B(n7747), .Z(n7934) );
  XNOR U8902 ( .A(b[5]), .B(a[58]), .Z(n7874) );
  NANDN U8903 ( .A(n7874), .B(n36587), .Z(n7751) );
  NANDN U8904 ( .A(n7749), .B(n36588), .Z(n7750) );
  AND U8905 ( .A(n7751), .B(n7750), .Z(n7935) );
  XNOR U8906 ( .A(n7934), .B(n7935), .Z(n7936) );
  XNOR U8907 ( .A(n7937), .B(n7936), .Z(n7923) );
  NAND U8908 ( .A(n7752), .B(n37762), .Z(n7754) );
  XOR U8909 ( .A(b[17]), .B(a[46]), .Z(n7877) );
  NAND U8910 ( .A(n7877), .B(n37764), .Z(n7753) );
  NAND U8911 ( .A(n7754), .B(n7753), .Z(n7895) );
  XNOR U8912 ( .A(b[31]), .B(a[32]), .Z(n7880) );
  NANDN U8913 ( .A(n7880), .B(n38552), .Z(n7757) );
  NANDN U8914 ( .A(n7755), .B(n38553), .Z(n7756) );
  NAND U8915 ( .A(n7757), .B(n7756), .Z(n7892) );
  OR U8916 ( .A(n7758), .B(n36105), .Z(n7760) );
  XNOR U8917 ( .A(b[3]), .B(a[60]), .Z(n7883) );
  NANDN U8918 ( .A(n7883), .B(n36107), .Z(n7759) );
  AND U8919 ( .A(n7760), .B(n7759), .Z(n7893) );
  XNOR U8920 ( .A(n7892), .B(n7893), .Z(n7894) );
  XOR U8921 ( .A(n7895), .B(n7894), .Z(n7922) );
  XNOR U8922 ( .A(n7923), .B(n7922), .Z(n7924) );
  XNOR U8923 ( .A(n7925), .B(n7924), .Z(n7972) );
  XNOR U8924 ( .A(n7971), .B(n7972), .Z(n7973) );
  XNOR U8925 ( .A(n7974), .B(n7973), .Z(n7859) );
  OR U8926 ( .A(n7762), .B(n7761), .Z(n7766) );
  NAND U8927 ( .A(n7764), .B(n7763), .Z(n7765) );
  NAND U8928 ( .A(n7766), .B(n7765), .Z(n7857) );
  NANDN U8929 ( .A(n7768), .B(n7767), .Z(n7772) );
  NANDN U8930 ( .A(n7770), .B(n7769), .Z(n7771) );
  NAND U8931 ( .A(n7772), .B(n7771), .Z(n7979) );
  OR U8932 ( .A(n7774), .B(n7773), .Z(n7778) );
  NAND U8933 ( .A(n7776), .B(n7775), .Z(n7777) );
  NAND U8934 ( .A(n7778), .B(n7777), .Z(n7978) );
  NANDN U8935 ( .A(n7780), .B(n7779), .Z(n7784) );
  NAND U8936 ( .A(n7782), .B(n7781), .Z(n7783) );
  NAND U8937 ( .A(n7784), .B(n7783), .Z(n7916) );
  NANDN U8938 ( .A(n7786), .B(n7785), .Z(n7790) );
  NAND U8939 ( .A(n7788), .B(n7787), .Z(n7789) );
  AND U8940 ( .A(n7790), .B(n7789), .Z(n7917) );
  XNOR U8941 ( .A(n7916), .B(n7917), .Z(n7918) );
  XOR U8942 ( .A(b[9]), .B(n11319), .Z(n7940) );
  NANDN U8943 ( .A(n7940), .B(n36925), .Z(n7793) );
  NANDN U8944 ( .A(n7791), .B(n36926), .Z(n7792) );
  NAND U8945 ( .A(n7793), .B(n7792), .Z(n7906) );
  XNOR U8946 ( .A(b[15]), .B(a[48]), .Z(n7943) );
  OR U8947 ( .A(n7943), .B(n37665), .Z(n7796) );
  NANDN U8948 ( .A(n7794), .B(n37604), .Z(n7795) );
  AND U8949 ( .A(n7796), .B(n7795), .Z(n7904) );
  XNOR U8950 ( .A(b[21]), .B(a[42]), .Z(n7946) );
  NANDN U8951 ( .A(n7946), .B(n38101), .Z(n7799) );
  NANDN U8952 ( .A(n7797), .B(n38102), .Z(n7798) );
  AND U8953 ( .A(n7799), .B(n7798), .Z(n7905) );
  XOR U8954 ( .A(n7906), .B(n7907), .Z(n7901) );
  XNOR U8955 ( .A(b[11]), .B(a[52]), .Z(n7949) );
  OR U8956 ( .A(n7949), .B(n37311), .Z(n7802) );
  NANDN U8957 ( .A(n7800), .B(n37218), .Z(n7801) );
  NAND U8958 ( .A(n7802), .B(n7801), .Z(n7899) );
  XOR U8959 ( .A(n1053), .B(a[50]), .Z(n7952) );
  NANDN U8960 ( .A(n7952), .B(n37424), .Z(n7805) );
  NANDN U8961 ( .A(n7803), .B(n37425), .Z(n7804) );
  AND U8962 ( .A(n7805), .B(n7804), .Z(n7898) );
  XNOR U8963 ( .A(n7899), .B(n7898), .Z(n7900) );
  XOR U8964 ( .A(n7901), .B(n7900), .Z(n7888) );
  NANDN U8965 ( .A(n1049), .B(a[62]), .Z(n7806) );
  XNOR U8966 ( .A(b[1]), .B(n7806), .Z(n7808) );
  NANDN U8967 ( .A(b[0]), .B(a[61]), .Z(n7807) );
  AND U8968 ( .A(n7808), .B(n7807), .Z(n7864) );
  NAND U8969 ( .A(n38490), .B(n7809), .Z(n7811) );
  XNOR U8970 ( .A(b[29]), .B(a[34]), .Z(n7956) );
  OR U8971 ( .A(n7956), .B(n1048), .Z(n7810) );
  NAND U8972 ( .A(n7811), .B(n7810), .Z(n7862) );
  NANDN U8973 ( .A(n1059), .B(a[30]), .Z(n7863) );
  XNOR U8974 ( .A(n7862), .B(n7863), .Z(n7865) );
  XOR U8975 ( .A(n7864), .B(n7865), .Z(n7886) );
  NANDN U8976 ( .A(n7812), .B(n38205), .Z(n7814) );
  XNOR U8977 ( .A(b[23]), .B(a[40]), .Z(n7962) );
  OR U8978 ( .A(n7962), .B(n38268), .Z(n7813) );
  NAND U8979 ( .A(n7814), .B(n7813), .Z(n7931) );
  XOR U8980 ( .A(b[7]), .B(a[56]), .Z(n7965) );
  NAND U8981 ( .A(n7965), .B(n36701), .Z(n7817) );
  NAND U8982 ( .A(n7815), .B(n36702), .Z(n7816) );
  NAND U8983 ( .A(n7817), .B(n7816), .Z(n7928) );
  XOR U8984 ( .A(b[25]), .B(a[38]), .Z(n7968) );
  NAND U8985 ( .A(n7968), .B(n38325), .Z(n7820) );
  NANDN U8986 ( .A(n7818), .B(n38326), .Z(n7819) );
  AND U8987 ( .A(n7820), .B(n7819), .Z(n7929) );
  XNOR U8988 ( .A(n7928), .B(n7929), .Z(n7930) );
  XNOR U8989 ( .A(n7931), .B(n7930), .Z(n7887) );
  XOR U8990 ( .A(n7886), .B(n7887), .Z(n7889) );
  XNOR U8991 ( .A(n7888), .B(n7889), .Z(n7919) );
  XNOR U8992 ( .A(n7918), .B(n7919), .Z(n7977) );
  XNOR U8993 ( .A(n7978), .B(n7977), .Z(n7980) );
  XNOR U8994 ( .A(n7979), .B(n7980), .Z(n7856) );
  XNOR U8995 ( .A(n7857), .B(n7856), .Z(n7858) );
  XOR U8996 ( .A(n7859), .B(n7858), .Z(n7853) );
  NANDN U8997 ( .A(n7822), .B(n7821), .Z(n7826) );
  OR U8998 ( .A(n7824), .B(n7823), .Z(n7825) );
  NAND U8999 ( .A(n7826), .B(n7825), .Z(n7850) );
  NAND U9000 ( .A(n7828), .B(n7827), .Z(n7832) );
  NANDN U9001 ( .A(n7830), .B(n7829), .Z(n7831) );
  NAND U9002 ( .A(n7832), .B(n7831), .Z(n7851) );
  XNOR U9003 ( .A(n7850), .B(n7851), .Z(n7852) );
  XOR U9004 ( .A(n7853), .B(n7852), .Z(n7847) );
  XOR U9005 ( .A(n7846), .B(n7847), .Z(n7838) );
  XOR U9006 ( .A(n7839), .B(n7838), .Z(n7840) );
  XNOR U9007 ( .A(n7841), .B(n7840), .Z(n7983) );
  XNOR U9008 ( .A(n7983), .B(sreg[286]), .Z(n7985) );
  NAND U9009 ( .A(n7833), .B(sreg[285]), .Z(n7837) );
  OR U9010 ( .A(n7835), .B(n7834), .Z(n7836) );
  AND U9011 ( .A(n7837), .B(n7836), .Z(n7984) );
  XOR U9012 ( .A(n7985), .B(n7984), .Z(c[286]) );
  NAND U9013 ( .A(n7839), .B(n7838), .Z(n7843) );
  NAND U9014 ( .A(n7841), .B(n7840), .Z(n7842) );
  NAND U9015 ( .A(n7843), .B(n7842), .Z(n7991) );
  NANDN U9016 ( .A(n7845), .B(n7844), .Z(n7849) );
  NAND U9017 ( .A(n7847), .B(n7846), .Z(n7848) );
  NAND U9018 ( .A(n7849), .B(n7848), .Z(n7989) );
  NANDN U9019 ( .A(n7851), .B(n7850), .Z(n7855) );
  NAND U9020 ( .A(n7853), .B(n7852), .Z(n7854) );
  NAND U9021 ( .A(n7855), .B(n7854), .Z(n7994) );
  NANDN U9022 ( .A(n7857), .B(n7856), .Z(n7861) );
  NANDN U9023 ( .A(n7859), .B(n7858), .Z(n7860) );
  NAND U9024 ( .A(n7861), .B(n7860), .Z(n7995) );
  XNOR U9025 ( .A(n7994), .B(n7995), .Z(n7996) );
  NANDN U9026 ( .A(n7863), .B(n7862), .Z(n7867) );
  NAND U9027 ( .A(n7865), .B(n7864), .Z(n7866) );
  NAND U9028 ( .A(n7867), .B(n7866), .Z(n8073) );
  XNOR U9029 ( .A(b[19]), .B(a[45]), .Z(n8040) );
  NANDN U9030 ( .A(n8040), .B(n37934), .Z(n7870) );
  NANDN U9031 ( .A(n7868), .B(n37935), .Z(n7869) );
  NAND U9032 ( .A(n7870), .B(n7869), .Z(n8085) );
  XNOR U9033 ( .A(b[27]), .B(a[37]), .Z(n8043) );
  NANDN U9034 ( .A(n8043), .B(n38423), .Z(n7873) );
  NAND U9035 ( .A(n7871), .B(n38424), .Z(n7872) );
  NAND U9036 ( .A(n7873), .B(n7872), .Z(n8082) );
  XOR U9037 ( .A(b[5]), .B(n12056), .Z(n8046) );
  NANDN U9038 ( .A(n8046), .B(n36587), .Z(n7876) );
  NANDN U9039 ( .A(n7874), .B(n36588), .Z(n7875) );
  AND U9040 ( .A(n7876), .B(n7875), .Z(n8083) );
  XNOR U9041 ( .A(n8082), .B(n8083), .Z(n8084) );
  XNOR U9042 ( .A(n8085), .B(n8084), .Z(n8070) );
  NAND U9043 ( .A(n7877), .B(n37762), .Z(n7879) );
  XOR U9044 ( .A(b[17]), .B(a[47]), .Z(n8049) );
  NAND U9045 ( .A(n8049), .B(n37764), .Z(n7878) );
  NAND U9046 ( .A(n7879), .B(n7878), .Z(n8024) );
  XNOR U9047 ( .A(b[31]), .B(a[33]), .Z(n8052) );
  NANDN U9048 ( .A(n8052), .B(n38552), .Z(n7882) );
  NANDN U9049 ( .A(n7880), .B(n38553), .Z(n7881) );
  AND U9050 ( .A(n7882), .B(n7881), .Z(n8022) );
  OR U9051 ( .A(n7883), .B(n36105), .Z(n7885) );
  XNOR U9052 ( .A(b[3]), .B(a[61]), .Z(n8055) );
  NANDN U9053 ( .A(n8055), .B(n36107), .Z(n7884) );
  AND U9054 ( .A(n7885), .B(n7884), .Z(n8023) );
  XOR U9055 ( .A(n8024), .B(n8025), .Z(n8071) );
  XOR U9056 ( .A(n8070), .B(n8071), .Z(n8072) );
  XNOR U9057 ( .A(n8073), .B(n8072), .Z(n8000) );
  NANDN U9058 ( .A(n7887), .B(n7886), .Z(n7891) );
  OR U9059 ( .A(n7889), .B(n7888), .Z(n7890) );
  NAND U9060 ( .A(n7891), .B(n7890), .Z(n8001) );
  XNOR U9061 ( .A(n8000), .B(n8001), .Z(n8002) );
  NANDN U9062 ( .A(n7893), .B(n7892), .Z(n7897) );
  NAND U9063 ( .A(n7895), .B(n7894), .Z(n7896) );
  NAND U9064 ( .A(n7897), .B(n7896), .Z(n8061) );
  NANDN U9065 ( .A(n7899), .B(n7898), .Z(n7903) );
  NAND U9066 ( .A(n7901), .B(n7900), .Z(n7902) );
  NAND U9067 ( .A(n7903), .B(n7902), .Z(n8058) );
  OR U9068 ( .A(n7905), .B(n7904), .Z(n7909) );
  NANDN U9069 ( .A(n7907), .B(n7906), .Z(n7908) );
  NAND U9070 ( .A(n7909), .B(n7908), .Z(n8059) );
  XNOR U9071 ( .A(n8058), .B(n8059), .Z(n8060) );
  XOR U9072 ( .A(n8061), .B(n8060), .Z(n8003) );
  XNOR U9073 ( .A(n8002), .B(n8003), .Z(n8127) );
  OR U9074 ( .A(n7911), .B(n7910), .Z(n7915) );
  NANDN U9075 ( .A(n7913), .B(n7912), .Z(n7914) );
  NAND U9076 ( .A(n7915), .B(n7914), .Z(n8125) );
  NANDN U9077 ( .A(n7917), .B(n7916), .Z(n7921) );
  NANDN U9078 ( .A(n7919), .B(n7918), .Z(n7920) );
  NAND U9079 ( .A(n7921), .B(n7920), .Z(n8006) );
  NANDN U9080 ( .A(n7923), .B(n7922), .Z(n7927) );
  NAND U9081 ( .A(n7925), .B(n7924), .Z(n7926) );
  NAND U9082 ( .A(n7927), .B(n7926), .Z(n8005) );
  NANDN U9083 ( .A(n7929), .B(n7928), .Z(n7933) );
  NAND U9084 ( .A(n7931), .B(n7930), .Z(n7932) );
  NAND U9085 ( .A(n7933), .B(n7932), .Z(n8064) );
  NANDN U9086 ( .A(n7935), .B(n7934), .Z(n7939) );
  NAND U9087 ( .A(n7937), .B(n7936), .Z(n7938) );
  AND U9088 ( .A(n7939), .B(n7938), .Z(n8065) );
  XNOR U9089 ( .A(n8064), .B(n8065), .Z(n8066) );
  XNOR U9090 ( .A(n1052), .B(a[55]), .Z(n8088) );
  NAND U9091 ( .A(n36925), .B(n8088), .Z(n7942) );
  NANDN U9092 ( .A(n7940), .B(n36926), .Z(n7941) );
  NAND U9093 ( .A(n7942), .B(n7941), .Z(n8030) );
  XNOR U9094 ( .A(b[15]), .B(a[49]), .Z(n8091) );
  OR U9095 ( .A(n8091), .B(n37665), .Z(n7945) );
  NANDN U9096 ( .A(n7943), .B(n37604), .Z(n7944) );
  AND U9097 ( .A(n7945), .B(n7944), .Z(n8028) );
  XNOR U9098 ( .A(n1056), .B(a[43]), .Z(n8094) );
  NAND U9099 ( .A(n8094), .B(n38101), .Z(n7948) );
  NANDN U9100 ( .A(n7946), .B(n38102), .Z(n7947) );
  AND U9101 ( .A(n7948), .B(n7947), .Z(n8029) );
  XOR U9102 ( .A(n8030), .B(n8031), .Z(n8019) );
  XNOR U9103 ( .A(b[11]), .B(a[53]), .Z(n8097) );
  OR U9104 ( .A(n8097), .B(n37311), .Z(n7951) );
  NANDN U9105 ( .A(n7949), .B(n37218), .Z(n7950) );
  NAND U9106 ( .A(n7951), .B(n7950), .Z(n8017) );
  XOR U9107 ( .A(n1053), .B(a[51]), .Z(n8100) );
  NANDN U9108 ( .A(n8100), .B(n37424), .Z(n7954) );
  NANDN U9109 ( .A(n7952), .B(n37425), .Z(n7953) );
  NAND U9110 ( .A(n7954), .B(n7953), .Z(n8016) );
  XOR U9111 ( .A(n8019), .B(n8018), .Z(n8013) );
  ANDN U9112 ( .B(b[31]), .A(n7955), .Z(n8034) );
  NANDN U9113 ( .A(n7956), .B(n38490), .Z(n7958) );
  XNOR U9114 ( .A(n1058), .B(a[35]), .Z(n8106) );
  NANDN U9115 ( .A(n1048), .B(n8106), .Z(n7957) );
  NAND U9116 ( .A(n7958), .B(n7957), .Z(n8035) );
  XOR U9117 ( .A(n8034), .B(n8035), .Z(n8036) );
  NANDN U9118 ( .A(n1049), .B(a[63]), .Z(n7959) );
  XNOR U9119 ( .A(b[1]), .B(n7959), .Z(n7961) );
  IV U9120 ( .A(a[62]), .Z(n12493) );
  NANDN U9121 ( .A(n12493), .B(n1049), .Z(n7960) );
  AND U9122 ( .A(n7961), .B(n7960), .Z(n8037) );
  XNOR U9123 ( .A(n8036), .B(n8037), .Z(n8010) );
  NANDN U9124 ( .A(n7962), .B(n38205), .Z(n7964) );
  XNOR U9125 ( .A(b[23]), .B(a[41]), .Z(n8109) );
  OR U9126 ( .A(n8109), .B(n38268), .Z(n7963) );
  NAND U9127 ( .A(n7964), .B(n7963), .Z(n8079) );
  XOR U9128 ( .A(b[7]), .B(a[57]), .Z(n8112) );
  NAND U9129 ( .A(n8112), .B(n36701), .Z(n7967) );
  NAND U9130 ( .A(n7965), .B(n36702), .Z(n7966) );
  NAND U9131 ( .A(n7967), .B(n7966), .Z(n8076) );
  XOR U9132 ( .A(b[25]), .B(a[39]), .Z(n8115) );
  NAND U9133 ( .A(n8115), .B(n38325), .Z(n7970) );
  NAND U9134 ( .A(n7968), .B(n38326), .Z(n7969) );
  AND U9135 ( .A(n7970), .B(n7969), .Z(n8077) );
  XNOR U9136 ( .A(n8076), .B(n8077), .Z(n8078) );
  XNOR U9137 ( .A(n8079), .B(n8078), .Z(n8011) );
  XOR U9138 ( .A(n8013), .B(n8012), .Z(n8067) );
  XNOR U9139 ( .A(n8066), .B(n8067), .Z(n8004) );
  XNOR U9140 ( .A(n8005), .B(n8004), .Z(n8007) );
  XNOR U9141 ( .A(n8006), .B(n8007), .Z(n8124) );
  XOR U9142 ( .A(n8125), .B(n8124), .Z(n8126) );
  XNOR U9143 ( .A(n8127), .B(n8126), .Z(n8121) );
  NANDN U9144 ( .A(n7972), .B(n7971), .Z(n7976) );
  NAND U9145 ( .A(n7974), .B(n7973), .Z(n7975) );
  NAND U9146 ( .A(n7976), .B(n7975), .Z(n8119) );
  NAND U9147 ( .A(n7978), .B(n7977), .Z(n7982) );
  NANDN U9148 ( .A(n7980), .B(n7979), .Z(n7981) );
  AND U9149 ( .A(n7982), .B(n7981), .Z(n8118) );
  XNOR U9150 ( .A(n8119), .B(n8118), .Z(n8120) );
  XOR U9151 ( .A(n8121), .B(n8120), .Z(n7997) );
  XOR U9152 ( .A(n7996), .B(n7997), .Z(n7988) );
  XOR U9153 ( .A(n7989), .B(n7988), .Z(n7990) );
  XNOR U9154 ( .A(n7991), .B(n7990), .Z(n8130) );
  XNOR U9155 ( .A(n8130), .B(sreg[287]), .Z(n8132) );
  NAND U9156 ( .A(n7983), .B(sreg[286]), .Z(n7987) );
  OR U9157 ( .A(n7985), .B(n7984), .Z(n7986) );
  AND U9158 ( .A(n7987), .B(n7986), .Z(n8131) );
  XOR U9159 ( .A(n8132), .B(n8131), .Z(c[287]) );
  NAND U9160 ( .A(n7989), .B(n7988), .Z(n7993) );
  NAND U9161 ( .A(n7991), .B(n7990), .Z(n7992) );
  NAND U9162 ( .A(n7993), .B(n7992), .Z(n8138) );
  NANDN U9163 ( .A(n7995), .B(n7994), .Z(n7999) );
  NAND U9164 ( .A(n7997), .B(n7996), .Z(n7998) );
  NAND U9165 ( .A(n7999), .B(n7998), .Z(n8136) );
  NAND U9166 ( .A(n8005), .B(n8004), .Z(n8009) );
  NANDN U9167 ( .A(n8007), .B(n8006), .Z(n8008) );
  NAND U9168 ( .A(n8009), .B(n8008), .Z(n8154) );
  XNOR U9169 ( .A(n8153), .B(n8154), .Z(n8155) );
  OR U9170 ( .A(n8011), .B(n8010), .Z(n8015) );
  NANDN U9171 ( .A(n8013), .B(n8012), .Z(n8014) );
  NAND U9172 ( .A(n8015), .B(n8014), .Z(n8268) );
  OR U9173 ( .A(n8017), .B(n8016), .Z(n8021) );
  NAND U9174 ( .A(n8019), .B(n8018), .Z(n8020) );
  NAND U9175 ( .A(n8021), .B(n8020), .Z(n8207) );
  OR U9176 ( .A(n8023), .B(n8022), .Z(n8027) );
  NANDN U9177 ( .A(n8025), .B(n8024), .Z(n8026) );
  NAND U9178 ( .A(n8027), .B(n8026), .Z(n8206) );
  OR U9179 ( .A(n8029), .B(n8028), .Z(n8033) );
  NANDN U9180 ( .A(n8031), .B(n8030), .Z(n8032) );
  NAND U9181 ( .A(n8033), .B(n8032), .Z(n8205) );
  XOR U9182 ( .A(n8207), .B(n8208), .Z(n8266) );
  OR U9183 ( .A(n8035), .B(n8034), .Z(n8039) );
  NANDN U9184 ( .A(n8037), .B(n8036), .Z(n8038) );
  NAND U9185 ( .A(n8039), .B(n8038), .Z(n8219) );
  XNOR U9186 ( .A(b[19]), .B(a[46]), .Z(n8165) );
  NANDN U9187 ( .A(n8165), .B(n37934), .Z(n8042) );
  NANDN U9188 ( .A(n8040), .B(n37935), .Z(n8041) );
  NAND U9189 ( .A(n8042), .B(n8041), .Z(n8256) );
  XOR U9190 ( .A(b[27]), .B(a[38]), .Z(n8168) );
  NAND U9191 ( .A(n38423), .B(n8168), .Z(n8045) );
  NANDN U9192 ( .A(n8043), .B(n38424), .Z(n8044) );
  NAND U9193 ( .A(n8045), .B(n8044), .Z(n8253) );
  XNOR U9194 ( .A(b[5]), .B(a[60]), .Z(n8171) );
  NANDN U9195 ( .A(n8171), .B(n36587), .Z(n8048) );
  NANDN U9196 ( .A(n8046), .B(n36588), .Z(n8047) );
  AND U9197 ( .A(n8048), .B(n8047), .Z(n8254) );
  XNOR U9198 ( .A(n8253), .B(n8254), .Z(n8255) );
  XNOR U9199 ( .A(n8256), .B(n8255), .Z(n8218) );
  NAND U9200 ( .A(n8049), .B(n37762), .Z(n8051) );
  XOR U9201 ( .A(b[17]), .B(a[48]), .Z(n8174) );
  NAND U9202 ( .A(n8174), .B(n37764), .Z(n8050) );
  NAND U9203 ( .A(n8051), .B(n8050), .Z(n8192) );
  XNOR U9204 ( .A(b[31]), .B(a[34]), .Z(n8177) );
  NANDN U9205 ( .A(n8177), .B(n38552), .Z(n8054) );
  NANDN U9206 ( .A(n8052), .B(n38553), .Z(n8053) );
  NAND U9207 ( .A(n8054), .B(n8053), .Z(n8189) );
  OR U9208 ( .A(n8055), .B(n36105), .Z(n8057) );
  XOR U9209 ( .A(b[3]), .B(n12493), .Z(n8180) );
  NANDN U9210 ( .A(n8180), .B(n36107), .Z(n8056) );
  AND U9211 ( .A(n8057), .B(n8056), .Z(n8190) );
  XNOR U9212 ( .A(n8189), .B(n8190), .Z(n8191) );
  XOR U9213 ( .A(n8192), .B(n8191), .Z(n8217) );
  XOR U9214 ( .A(n8218), .B(n8217), .Z(n8220) );
  XOR U9215 ( .A(n8219), .B(n8220), .Z(n8265) );
  XOR U9216 ( .A(n8266), .B(n8265), .Z(n8267) );
  XNOR U9217 ( .A(n8268), .B(n8267), .Z(n8150) );
  NANDN U9218 ( .A(n8059), .B(n8058), .Z(n8063) );
  NANDN U9219 ( .A(n8061), .B(n8060), .Z(n8062) );
  NAND U9220 ( .A(n8063), .B(n8062), .Z(n8147) );
  NANDN U9221 ( .A(n8065), .B(n8064), .Z(n8069) );
  NANDN U9222 ( .A(n8067), .B(n8066), .Z(n8068) );
  NAND U9223 ( .A(n8069), .B(n8068), .Z(n8274) );
  OR U9224 ( .A(n8071), .B(n8070), .Z(n8075) );
  NAND U9225 ( .A(n8073), .B(n8072), .Z(n8074) );
  NAND U9226 ( .A(n8075), .B(n8074), .Z(n8272) );
  NANDN U9227 ( .A(n8077), .B(n8076), .Z(n8081) );
  NAND U9228 ( .A(n8079), .B(n8078), .Z(n8080) );
  NAND U9229 ( .A(n8081), .B(n8080), .Z(n8211) );
  NANDN U9230 ( .A(n8083), .B(n8082), .Z(n8087) );
  NAND U9231 ( .A(n8085), .B(n8084), .Z(n8086) );
  AND U9232 ( .A(n8087), .B(n8086), .Z(n8212) );
  XNOR U9233 ( .A(n8211), .B(n8212), .Z(n8213) );
  XNOR U9234 ( .A(b[9]), .B(a[56]), .Z(n8223) );
  NANDN U9235 ( .A(n8223), .B(n36925), .Z(n8090) );
  NAND U9236 ( .A(n36926), .B(n8088), .Z(n8089) );
  NAND U9237 ( .A(n8090), .B(n8089), .Z(n8197) );
  XNOR U9238 ( .A(n1054), .B(a[50]), .Z(n8226) );
  NANDN U9239 ( .A(n37665), .B(n8226), .Z(n8093) );
  NANDN U9240 ( .A(n8091), .B(n37604), .Z(n8092) );
  NAND U9241 ( .A(n8093), .B(n8092), .Z(n8195) );
  XOR U9242 ( .A(b[21]), .B(n9873), .Z(n8229) );
  NANDN U9243 ( .A(n8229), .B(n38101), .Z(n8096) );
  NAND U9244 ( .A(n38102), .B(n8094), .Z(n8095) );
  NAND U9245 ( .A(n8096), .B(n8095), .Z(n8196) );
  XNOR U9246 ( .A(n8195), .B(n8196), .Z(n8198) );
  XOR U9247 ( .A(n8197), .B(n8198), .Z(n8186) );
  XOR U9248 ( .A(b[11]), .B(n11319), .Z(n8232) );
  OR U9249 ( .A(n8232), .B(n37311), .Z(n8099) );
  NANDN U9250 ( .A(n8097), .B(n37218), .Z(n8098) );
  NAND U9251 ( .A(n8099), .B(n8098), .Z(n8184) );
  XOR U9252 ( .A(n1053), .B(a[52]), .Z(n8235) );
  NANDN U9253 ( .A(n8235), .B(n37424), .Z(n8102) );
  NANDN U9254 ( .A(n8100), .B(n37425), .Z(n8101) );
  AND U9255 ( .A(n8102), .B(n8101), .Z(n8183) );
  XNOR U9256 ( .A(n8184), .B(n8183), .Z(n8185) );
  XNOR U9257 ( .A(n8186), .B(n8185), .Z(n8202) );
  NANDN U9258 ( .A(n1049), .B(a[64]), .Z(n8103) );
  XNOR U9259 ( .A(b[1]), .B(n8103), .Z(n8105) );
  NANDN U9260 ( .A(b[0]), .B(a[63]), .Z(n8104) );
  AND U9261 ( .A(n8105), .B(n8104), .Z(n8161) );
  NAND U9262 ( .A(n8106), .B(n38490), .Z(n8108) );
  XNOR U9263 ( .A(n1058), .B(a[36]), .Z(n8241) );
  NANDN U9264 ( .A(n1048), .B(n8241), .Z(n8107) );
  NAND U9265 ( .A(n8108), .B(n8107), .Z(n8159) );
  NANDN U9266 ( .A(n1059), .B(a[32]), .Z(n8160) );
  XNOR U9267 ( .A(n8159), .B(n8160), .Z(n8162) );
  XNOR U9268 ( .A(n8161), .B(n8162), .Z(n8200) );
  NANDN U9269 ( .A(n8109), .B(n38205), .Z(n8111) );
  XNOR U9270 ( .A(b[23]), .B(a[42]), .Z(n8244) );
  OR U9271 ( .A(n8244), .B(n38268), .Z(n8110) );
  NAND U9272 ( .A(n8111), .B(n8110), .Z(n8262) );
  XOR U9273 ( .A(b[7]), .B(a[58]), .Z(n8247) );
  NAND U9274 ( .A(n8247), .B(n36701), .Z(n8114) );
  NAND U9275 ( .A(n8112), .B(n36702), .Z(n8113) );
  NAND U9276 ( .A(n8114), .B(n8113), .Z(n8259) );
  XOR U9277 ( .A(b[25]), .B(a[40]), .Z(n8250) );
  NAND U9278 ( .A(n8250), .B(n38325), .Z(n8117) );
  NAND U9279 ( .A(n8115), .B(n38326), .Z(n8116) );
  AND U9280 ( .A(n8117), .B(n8116), .Z(n8260) );
  XNOR U9281 ( .A(n8259), .B(n8260), .Z(n8261) );
  XOR U9282 ( .A(n8262), .B(n8261), .Z(n8199) );
  XOR U9283 ( .A(n8202), .B(n8201), .Z(n8214) );
  XOR U9284 ( .A(n8213), .B(n8214), .Z(n8271) );
  XOR U9285 ( .A(n8272), .B(n8271), .Z(n8273) );
  XOR U9286 ( .A(n8274), .B(n8273), .Z(n8148) );
  XNOR U9287 ( .A(n8147), .B(n8148), .Z(n8149) );
  XOR U9288 ( .A(n8150), .B(n8149), .Z(n8156) );
  XOR U9289 ( .A(n8155), .B(n8156), .Z(n8143) );
  NANDN U9290 ( .A(n8119), .B(n8118), .Z(n8123) );
  NAND U9291 ( .A(n8121), .B(n8120), .Z(n8122) );
  NAND U9292 ( .A(n8123), .B(n8122), .Z(n8141) );
  NANDN U9293 ( .A(n8125), .B(n8124), .Z(n8129) );
  OR U9294 ( .A(n8127), .B(n8126), .Z(n8128) );
  NAND U9295 ( .A(n8129), .B(n8128), .Z(n8142) );
  XNOR U9296 ( .A(n8141), .B(n8142), .Z(n8144) );
  XOR U9297 ( .A(n8143), .B(n8144), .Z(n8135) );
  XOR U9298 ( .A(n8136), .B(n8135), .Z(n8137) );
  XNOR U9299 ( .A(n8138), .B(n8137), .Z(n8277) );
  XNOR U9300 ( .A(n8277), .B(sreg[288]), .Z(n8279) );
  NAND U9301 ( .A(n8130), .B(sreg[287]), .Z(n8134) );
  OR U9302 ( .A(n8132), .B(n8131), .Z(n8133) );
  AND U9303 ( .A(n8134), .B(n8133), .Z(n8278) );
  XOR U9304 ( .A(n8279), .B(n8278), .Z(c[288]) );
  NAND U9305 ( .A(n8136), .B(n8135), .Z(n8140) );
  NAND U9306 ( .A(n8138), .B(n8137), .Z(n8139) );
  NAND U9307 ( .A(n8140), .B(n8139), .Z(n8285) );
  NANDN U9308 ( .A(n8142), .B(n8141), .Z(n8146) );
  NAND U9309 ( .A(n8144), .B(n8143), .Z(n8145) );
  NAND U9310 ( .A(n8146), .B(n8145), .Z(n8283) );
  NANDN U9311 ( .A(n8148), .B(n8147), .Z(n8152) );
  NAND U9312 ( .A(n8150), .B(n8149), .Z(n8151) );
  NAND U9313 ( .A(n8152), .B(n8151), .Z(n8288) );
  NANDN U9314 ( .A(n8154), .B(n8153), .Z(n8158) );
  NAND U9315 ( .A(n8156), .B(n8155), .Z(n8157) );
  AND U9316 ( .A(n8158), .B(n8157), .Z(n8289) );
  XNOR U9317 ( .A(n8288), .B(n8289), .Z(n8290) );
  NANDN U9318 ( .A(n8160), .B(n8159), .Z(n8164) );
  NAND U9319 ( .A(n8162), .B(n8161), .Z(n8163) );
  NAND U9320 ( .A(n8164), .B(n8163), .Z(n8365) );
  XNOR U9321 ( .A(b[19]), .B(a[47]), .Z(n8310) );
  NANDN U9322 ( .A(n8310), .B(n37934), .Z(n8167) );
  NANDN U9323 ( .A(n8165), .B(n37935), .Z(n8166) );
  NAND U9324 ( .A(n8167), .B(n8166), .Z(n8375) );
  XOR U9325 ( .A(b[27]), .B(a[39]), .Z(n8313) );
  NAND U9326 ( .A(n38423), .B(n8313), .Z(n8170) );
  NAND U9327 ( .A(n8168), .B(n38424), .Z(n8169) );
  NAND U9328 ( .A(n8170), .B(n8169), .Z(n8372) );
  XNOR U9329 ( .A(b[5]), .B(a[61]), .Z(n8316) );
  NANDN U9330 ( .A(n8316), .B(n36587), .Z(n8173) );
  NANDN U9331 ( .A(n8171), .B(n36588), .Z(n8172) );
  AND U9332 ( .A(n8173), .B(n8172), .Z(n8373) );
  XNOR U9333 ( .A(n8372), .B(n8373), .Z(n8374) );
  XNOR U9334 ( .A(n8375), .B(n8374), .Z(n8363) );
  NAND U9335 ( .A(n8174), .B(n37762), .Z(n8176) );
  XOR U9336 ( .A(b[17]), .B(a[49]), .Z(n8319) );
  NAND U9337 ( .A(n8319), .B(n37764), .Z(n8175) );
  NAND U9338 ( .A(n8176), .B(n8175), .Z(n8337) );
  XNOR U9339 ( .A(b[31]), .B(a[35]), .Z(n8322) );
  NANDN U9340 ( .A(n8322), .B(n38552), .Z(n8179) );
  NANDN U9341 ( .A(n8177), .B(n38553), .Z(n8178) );
  NAND U9342 ( .A(n8179), .B(n8178), .Z(n8334) );
  OR U9343 ( .A(n8180), .B(n36105), .Z(n8182) );
  XNOR U9344 ( .A(b[3]), .B(a[63]), .Z(n8325) );
  NANDN U9345 ( .A(n8325), .B(n36107), .Z(n8181) );
  AND U9346 ( .A(n8182), .B(n8181), .Z(n8335) );
  XNOR U9347 ( .A(n8334), .B(n8335), .Z(n8336) );
  XOR U9348 ( .A(n8337), .B(n8336), .Z(n8362) );
  XNOR U9349 ( .A(n8363), .B(n8362), .Z(n8364) );
  XNOR U9350 ( .A(n8365), .B(n8364), .Z(n8301) );
  NANDN U9351 ( .A(n8184), .B(n8183), .Z(n8188) );
  NAND U9352 ( .A(n8186), .B(n8185), .Z(n8187) );
  NAND U9353 ( .A(n8188), .B(n8187), .Z(n8354) );
  NANDN U9354 ( .A(n8190), .B(n8189), .Z(n8194) );
  NAND U9355 ( .A(n8192), .B(n8191), .Z(n8193) );
  NAND U9356 ( .A(n8194), .B(n8193), .Z(n8353) );
  XNOR U9357 ( .A(n8353), .B(n8352), .Z(n8355) );
  XOR U9358 ( .A(n8354), .B(n8355), .Z(n8300) );
  XOR U9359 ( .A(n8301), .B(n8300), .Z(n8302) );
  NANDN U9360 ( .A(n8200), .B(n8199), .Z(n8204) );
  NAND U9361 ( .A(n8202), .B(n8201), .Z(n8203) );
  NAND U9362 ( .A(n8204), .B(n8203), .Z(n8303) );
  XNOR U9363 ( .A(n8302), .B(n8303), .Z(n8416) );
  OR U9364 ( .A(n8206), .B(n8205), .Z(n8210) );
  NANDN U9365 ( .A(n8208), .B(n8207), .Z(n8209) );
  NAND U9366 ( .A(n8210), .B(n8209), .Z(n8415) );
  NANDN U9367 ( .A(n8212), .B(n8211), .Z(n8216) );
  NAND U9368 ( .A(n8214), .B(n8213), .Z(n8215) );
  NAND U9369 ( .A(n8216), .B(n8215), .Z(n8297) );
  NANDN U9370 ( .A(n8218), .B(n8217), .Z(n8222) );
  OR U9371 ( .A(n8220), .B(n8219), .Z(n8221) );
  NAND U9372 ( .A(n8222), .B(n8221), .Z(n8294) );
  XNOR U9373 ( .A(b[9]), .B(a[57]), .Z(n8378) );
  NANDN U9374 ( .A(n8378), .B(n36925), .Z(n8225) );
  NANDN U9375 ( .A(n8223), .B(n36926), .Z(n8224) );
  NAND U9376 ( .A(n8225), .B(n8224), .Z(n8342) );
  XNOR U9377 ( .A(b[15]), .B(a[51]), .Z(n8381) );
  OR U9378 ( .A(n8381), .B(n37665), .Z(n8228) );
  NAND U9379 ( .A(n8226), .B(n37604), .Z(n8227) );
  AND U9380 ( .A(n8228), .B(n8227), .Z(n8340) );
  XNOR U9381 ( .A(b[21]), .B(a[45]), .Z(n8384) );
  NANDN U9382 ( .A(n8384), .B(n38101), .Z(n8231) );
  NANDN U9383 ( .A(n8229), .B(n38102), .Z(n8230) );
  AND U9384 ( .A(n8231), .B(n8230), .Z(n8341) );
  XOR U9385 ( .A(n8342), .B(n8343), .Z(n8331) );
  XNOR U9386 ( .A(b[11]), .B(a[55]), .Z(n8387) );
  OR U9387 ( .A(n8387), .B(n37311), .Z(n8234) );
  NANDN U9388 ( .A(n8232), .B(n37218), .Z(n8233) );
  NAND U9389 ( .A(n8234), .B(n8233), .Z(n8329) );
  XOR U9390 ( .A(n1053), .B(a[53]), .Z(n8390) );
  NANDN U9391 ( .A(n8390), .B(n37424), .Z(n8237) );
  NANDN U9392 ( .A(n8235), .B(n37425), .Z(n8236) );
  AND U9393 ( .A(n8237), .B(n8236), .Z(n8328) );
  XNOR U9394 ( .A(n8329), .B(n8328), .Z(n8330) );
  XOR U9395 ( .A(n8331), .B(n8330), .Z(n8349) );
  NANDN U9396 ( .A(n1049), .B(a[65]), .Z(n8238) );
  XNOR U9397 ( .A(b[1]), .B(n8238), .Z(n8240) );
  NANDN U9398 ( .A(b[0]), .B(a[64]), .Z(n8239) );
  AND U9399 ( .A(n8240), .B(n8239), .Z(n8306) );
  NAND U9400 ( .A(n38490), .B(n8241), .Z(n8243) );
  XOR U9401 ( .A(n1058), .B(n8832), .Z(n8396) );
  NANDN U9402 ( .A(n1048), .B(n8396), .Z(n8242) );
  NAND U9403 ( .A(n8243), .B(n8242), .Z(n8304) );
  NANDN U9404 ( .A(n1059), .B(a[33]), .Z(n8305) );
  XNOR U9405 ( .A(n8304), .B(n8305), .Z(n8307) );
  XOR U9406 ( .A(n8306), .B(n8307), .Z(n8346) );
  NANDN U9407 ( .A(n8244), .B(n38205), .Z(n8246) );
  XNOR U9408 ( .A(b[23]), .B(a[43]), .Z(n8399) );
  OR U9409 ( .A(n8399), .B(n38268), .Z(n8245) );
  NAND U9410 ( .A(n8246), .B(n8245), .Z(n8369) );
  XNOR U9411 ( .A(b[7]), .B(a[59]), .Z(n8402) );
  NANDN U9412 ( .A(n8402), .B(n36701), .Z(n8249) );
  NAND U9413 ( .A(n8247), .B(n36702), .Z(n8248) );
  NAND U9414 ( .A(n8249), .B(n8248), .Z(n8366) );
  XOR U9415 ( .A(b[25]), .B(a[41]), .Z(n8405) );
  NAND U9416 ( .A(n8405), .B(n38325), .Z(n8252) );
  NAND U9417 ( .A(n8250), .B(n38326), .Z(n8251) );
  AND U9418 ( .A(n8252), .B(n8251), .Z(n8367) );
  XNOR U9419 ( .A(n8366), .B(n8367), .Z(n8368) );
  XNOR U9420 ( .A(n8369), .B(n8368), .Z(n8347) );
  XNOR U9421 ( .A(n8346), .B(n8347), .Z(n8348) );
  XNOR U9422 ( .A(n8349), .B(n8348), .Z(n8359) );
  NANDN U9423 ( .A(n8254), .B(n8253), .Z(n8258) );
  NAND U9424 ( .A(n8256), .B(n8255), .Z(n8257) );
  NAND U9425 ( .A(n8258), .B(n8257), .Z(n8357) );
  NANDN U9426 ( .A(n8260), .B(n8259), .Z(n8264) );
  NAND U9427 ( .A(n8262), .B(n8261), .Z(n8263) );
  AND U9428 ( .A(n8264), .B(n8263), .Z(n8356) );
  XNOR U9429 ( .A(n8357), .B(n8356), .Z(n8358) );
  XNOR U9430 ( .A(n8359), .B(n8358), .Z(n8295) );
  XNOR U9431 ( .A(n8294), .B(n8295), .Z(n8296) );
  XOR U9432 ( .A(n8297), .B(n8296), .Z(n8414) );
  XOR U9433 ( .A(n8415), .B(n8414), .Z(n8417) );
  NAND U9434 ( .A(n8266), .B(n8265), .Z(n8270) );
  NAND U9435 ( .A(n8268), .B(n8267), .Z(n8269) );
  NAND U9436 ( .A(n8270), .B(n8269), .Z(n8409) );
  NAND U9437 ( .A(n8272), .B(n8271), .Z(n8276) );
  NAND U9438 ( .A(n8274), .B(n8273), .Z(n8275) );
  AND U9439 ( .A(n8276), .B(n8275), .Z(n8408) );
  XNOR U9440 ( .A(n8409), .B(n8408), .Z(n8410) );
  XOR U9441 ( .A(n8411), .B(n8410), .Z(n8291) );
  XOR U9442 ( .A(n8290), .B(n8291), .Z(n8282) );
  XOR U9443 ( .A(n8283), .B(n8282), .Z(n8284) );
  XNOR U9444 ( .A(n8285), .B(n8284), .Z(n8420) );
  XNOR U9445 ( .A(n8420), .B(sreg[289]), .Z(n8422) );
  NAND U9446 ( .A(n8277), .B(sreg[288]), .Z(n8281) );
  OR U9447 ( .A(n8279), .B(n8278), .Z(n8280) );
  AND U9448 ( .A(n8281), .B(n8280), .Z(n8421) );
  XOR U9449 ( .A(n8422), .B(n8421), .Z(c[289]) );
  NAND U9450 ( .A(n8283), .B(n8282), .Z(n8287) );
  NAND U9451 ( .A(n8285), .B(n8284), .Z(n8286) );
  NAND U9452 ( .A(n8287), .B(n8286), .Z(n8428) );
  NANDN U9453 ( .A(n8289), .B(n8288), .Z(n8293) );
  NAND U9454 ( .A(n8291), .B(n8290), .Z(n8292) );
  NAND U9455 ( .A(n8293), .B(n8292), .Z(n8425) );
  NANDN U9456 ( .A(n8295), .B(n8294), .Z(n8299) );
  NAND U9457 ( .A(n8297), .B(n8296), .Z(n8298) );
  NAND U9458 ( .A(n8299), .B(n8298), .Z(n8437) );
  XNOR U9459 ( .A(n8437), .B(n8438), .Z(n8439) );
  NANDN U9460 ( .A(n8305), .B(n8304), .Z(n8309) );
  NAND U9461 ( .A(n8307), .B(n8306), .Z(n8308) );
  NAND U9462 ( .A(n8309), .B(n8308), .Z(n8510) );
  XNOR U9463 ( .A(b[19]), .B(a[48]), .Z(n8453) );
  NANDN U9464 ( .A(n8453), .B(n37934), .Z(n8312) );
  NANDN U9465 ( .A(n8310), .B(n37935), .Z(n8311) );
  NAND U9466 ( .A(n8312), .B(n8311), .Z(n8520) );
  XOR U9467 ( .A(b[27]), .B(a[40]), .Z(n8456) );
  NAND U9468 ( .A(n38423), .B(n8456), .Z(n8315) );
  NAND U9469 ( .A(n8313), .B(n38424), .Z(n8314) );
  NAND U9470 ( .A(n8315), .B(n8314), .Z(n8517) );
  XOR U9471 ( .A(b[5]), .B(n12493), .Z(n8459) );
  NANDN U9472 ( .A(n8459), .B(n36587), .Z(n8318) );
  NANDN U9473 ( .A(n8316), .B(n36588), .Z(n8317) );
  AND U9474 ( .A(n8318), .B(n8317), .Z(n8518) );
  XNOR U9475 ( .A(n8517), .B(n8518), .Z(n8519) );
  XNOR U9476 ( .A(n8520), .B(n8519), .Z(n8508) );
  NAND U9477 ( .A(n8319), .B(n37762), .Z(n8321) );
  XNOR U9478 ( .A(b[17]), .B(a[50]), .Z(n8462) );
  NANDN U9479 ( .A(n8462), .B(n37764), .Z(n8320) );
  NAND U9480 ( .A(n8321), .B(n8320), .Z(n8480) );
  XNOR U9481 ( .A(b[31]), .B(a[36]), .Z(n8465) );
  NANDN U9482 ( .A(n8465), .B(n38552), .Z(n8324) );
  NANDN U9483 ( .A(n8322), .B(n38553), .Z(n8323) );
  NAND U9484 ( .A(n8324), .B(n8323), .Z(n8477) );
  OR U9485 ( .A(n8325), .B(n36105), .Z(n8327) );
  XNOR U9486 ( .A(b[3]), .B(a[64]), .Z(n8468) );
  NANDN U9487 ( .A(n8468), .B(n36107), .Z(n8326) );
  AND U9488 ( .A(n8327), .B(n8326), .Z(n8478) );
  XNOR U9489 ( .A(n8477), .B(n8478), .Z(n8479) );
  XOR U9490 ( .A(n8480), .B(n8479), .Z(n8507) );
  XNOR U9491 ( .A(n8508), .B(n8507), .Z(n8509) );
  XNOR U9492 ( .A(n8510), .B(n8509), .Z(n8553) );
  NANDN U9493 ( .A(n8329), .B(n8328), .Z(n8333) );
  NAND U9494 ( .A(n8331), .B(n8330), .Z(n8332) );
  NAND U9495 ( .A(n8333), .B(n8332), .Z(n8498) );
  NANDN U9496 ( .A(n8335), .B(n8334), .Z(n8339) );
  NAND U9497 ( .A(n8337), .B(n8336), .Z(n8338) );
  NAND U9498 ( .A(n8339), .B(n8338), .Z(n8496) );
  OR U9499 ( .A(n8341), .B(n8340), .Z(n8345) );
  NANDN U9500 ( .A(n8343), .B(n8342), .Z(n8344) );
  NAND U9501 ( .A(n8345), .B(n8344), .Z(n8495) );
  XNOR U9502 ( .A(n8498), .B(n8497), .Z(n8554) );
  XNOR U9503 ( .A(n8553), .B(n8554), .Z(n8555) );
  NANDN U9504 ( .A(n8347), .B(n8346), .Z(n8351) );
  NANDN U9505 ( .A(n8349), .B(n8348), .Z(n8350) );
  AND U9506 ( .A(n8351), .B(n8350), .Z(n8556) );
  XOR U9507 ( .A(n8555), .B(n8556), .Z(n8446) );
  NANDN U9508 ( .A(n8357), .B(n8356), .Z(n8361) );
  NANDN U9509 ( .A(n8359), .B(n8358), .Z(n8360) );
  NAND U9510 ( .A(n8361), .B(n8360), .Z(n8562) );
  NANDN U9511 ( .A(n8367), .B(n8366), .Z(n8371) );
  NAND U9512 ( .A(n8369), .B(n8368), .Z(n8370) );
  NAND U9513 ( .A(n8371), .B(n8370), .Z(n8501) );
  NANDN U9514 ( .A(n8373), .B(n8372), .Z(n8377) );
  NAND U9515 ( .A(n8375), .B(n8374), .Z(n8376) );
  AND U9516 ( .A(n8377), .B(n8376), .Z(n8502) );
  XNOR U9517 ( .A(n8501), .B(n8502), .Z(n8503) );
  XNOR U9518 ( .A(b[9]), .B(a[58]), .Z(n8523) );
  NANDN U9519 ( .A(n8523), .B(n36925), .Z(n8380) );
  NANDN U9520 ( .A(n8378), .B(n36926), .Z(n8379) );
  NAND U9521 ( .A(n8380), .B(n8379), .Z(n8485) );
  XNOR U9522 ( .A(b[15]), .B(a[52]), .Z(n8526) );
  OR U9523 ( .A(n8526), .B(n37665), .Z(n8383) );
  NANDN U9524 ( .A(n8381), .B(n37604), .Z(n8382) );
  AND U9525 ( .A(n8383), .B(n8382), .Z(n8483) );
  XNOR U9526 ( .A(b[21]), .B(a[46]), .Z(n8529) );
  NANDN U9527 ( .A(n8529), .B(n38101), .Z(n8386) );
  NANDN U9528 ( .A(n8384), .B(n38102), .Z(n8385) );
  AND U9529 ( .A(n8386), .B(n8385), .Z(n8484) );
  XOR U9530 ( .A(n8485), .B(n8486), .Z(n8474) );
  XNOR U9531 ( .A(b[11]), .B(a[56]), .Z(n8532) );
  OR U9532 ( .A(n8532), .B(n37311), .Z(n8389) );
  NANDN U9533 ( .A(n8387), .B(n37218), .Z(n8388) );
  NAND U9534 ( .A(n8389), .B(n8388), .Z(n8472) );
  XOR U9535 ( .A(n1053), .B(a[54]), .Z(n8535) );
  NANDN U9536 ( .A(n8535), .B(n37424), .Z(n8392) );
  NANDN U9537 ( .A(n8390), .B(n37425), .Z(n8391) );
  AND U9538 ( .A(n8392), .B(n8391), .Z(n8471) );
  XNOR U9539 ( .A(n8472), .B(n8471), .Z(n8473) );
  XOR U9540 ( .A(n8474), .B(n8473), .Z(n8491) );
  NANDN U9541 ( .A(n1049), .B(a[66]), .Z(n8393) );
  XNOR U9542 ( .A(b[1]), .B(n8393), .Z(n8395) );
  NANDN U9543 ( .A(b[0]), .B(a[65]), .Z(n8394) );
  AND U9544 ( .A(n8395), .B(n8394), .Z(n8449) );
  NAND U9545 ( .A(n38490), .B(n8396), .Z(n8398) );
  XNOR U9546 ( .A(n1058), .B(a[38]), .Z(n8541) );
  NANDN U9547 ( .A(n1048), .B(n8541), .Z(n8397) );
  NAND U9548 ( .A(n8398), .B(n8397), .Z(n8447) );
  NANDN U9549 ( .A(n1059), .B(a[34]), .Z(n8448) );
  XNOR U9550 ( .A(n8447), .B(n8448), .Z(n8450) );
  XOR U9551 ( .A(n8449), .B(n8450), .Z(n8489) );
  NANDN U9552 ( .A(n8399), .B(n38205), .Z(n8401) );
  XOR U9553 ( .A(b[23]), .B(n9873), .Z(n8544) );
  OR U9554 ( .A(n8544), .B(n38268), .Z(n8400) );
  NAND U9555 ( .A(n8401), .B(n8400), .Z(n8514) );
  XOR U9556 ( .A(b[7]), .B(a[60]), .Z(n8547) );
  NAND U9557 ( .A(n8547), .B(n36701), .Z(n8404) );
  NANDN U9558 ( .A(n8402), .B(n36702), .Z(n8403) );
  NAND U9559 ( .A(n8404), .B(n8403), .Z(n8511) );
  XOR U9560 ( .A(b[25]), .B(a[42]), .Z(n8550) );
  NAND U9561 ( .A(n8550), .B(n38325), .Z(n8407) );
  NAND U9562 ( .A(n8405), .B(n38326), .Z(n8406) );
  AND U9563 ( .A(n8407), .B(n8406), .Z(n8512) );
  XNOR U9564 ( .A(n8511), .B(n8512), .Z(n8513) );
  XNOR U9565 ( .A(n8514), .B(n8513), .Z(n8490) );
  XOR U9566 ( .A(n8489), .B(n8490), .Z(n8492) );
  XNOR U9567 ( .A(n8491), .B(n8492), .Z(n8504) );
  XNOR U9568 ( .A(n8503), .B(n8504), .Z(n8559) );
  XNOR U9569 ( .A(n8560), .B(n8559), .Z(n8561) );
  XOR U9570 ( .A(n8562), .B(n8561), .Z(n8443) );
  XNOR U9571 ( .A(n8444), .B(n8443), .Z(n8445) );
  XOR U9572 ( .A(n8446), .B(n8445), .Z(n8440) );
  XOR U9573 ( .A(n8439), .B(n8440), .Z(n8434) );
  NANDN U9574 ( .A(n8409), .B(n8408), .Z(n8413) );
  NAND U9575 ( .A(n8411), .B(n8410), .Z(n8412) );
  NAND U9576 ( .A(n8413), .B(n8412), .Z(n8431) );
  NANDN U9577 ( .A(n8415), .B(n8414), .Z(n8419) );
  OR U9578 ( .A(n8417), .B(n8416), .Z(n8418) );
  NAND U9579 ( .A(n8419), .B(n8418), .Z(n8432) );
  XNOR U9580 ( .A(n8431), .B(n8432), .Z(n8433) );
  XNOR U9581 ( .A(n8434), .B(n8433), .Z(n8426) );
  XNOR U9582 ( .A(n8425), .B(n8426), .Z(n8427) );
  XNOR U9583 ( .A(n8428), .B(n8427), .Z(n8565) );
  XNOR U9584 ( .A(n8565), .B(sreg[290]), .Z(n8567) );
  NAND U9585 ( .A(n8420), .B(sreg[289]), .Z(n8424) );
  OR U9586 ( .A(n8422), .B(n8421), .Z(n8423) );
  AND U9587 ( .A(n8424), .B(n8423), .Z(n8566) );
  XOR U9588 ( .A(n8567), .B(n8566), .Z(c[290]) );
  NANDN U9589 ( .A(n8426), .B(n8425), .Z(n8430) );
  NAND U9590 ( .A(n8428), .B(n8427), .Z(n8429) );
  NAND U9591 ( .A(n8430), .B(n8429), .Z(n8573) );
  NANDN U9592 ( .A(n8432), .B(n8431), .Z(n8436) );
  NAND U9593 ( .A(n8434), .B(n8433), .Z(n8435) );
  NAND U9594 ( .A(n8436), .B(n8435), .Z(n8571) );
  NANDN U9595 ( .A(n8438), .B(n8437), .Z(n8442) );
  NANDN U9596 ( .A(n8440), .B(n8439), .Z(n8441) );
  NAND U9597 ( .A(n8442), .B(n8441), .Z(n8577) );
  XNOR U9598 ( .A(n8577), .B(n8576), .Z(n8578) );
  NANDN U9599 ( .A(n8448), .B(n8447), .Z(n8452) );
  NAND U9600 ( .A(n8450), .B(n8449), .Z(n8451) );
  NAND U9601 ( .A(n8452), .B(n8451), .Z(n8657) );
  XNOR U9602 ( .A(b[19]), .B(a[49]), .Z(n8600) );
  NANDN U9603 ( .A(n8600), .B(n37934), .Z(n8455) );
  NANDN U9604 ( .A(n8453), .B(n37935), .Z(n8454) );
  NAND U9605 ( .A(n8455), .B(n8454), .Z(n8667) );
  XOR U9606 ( .A(b[27]), .B(a[41]), .Z(n8603) );
  NAND U9607 ( .A(n38423), .B(n8603), .Z(n8458) );
  NAND U9608 ( .A(n8456), .B(n38424), .Z(n8457) );
  NAND U9609 ( .A(n8458), .B(n8457), .Z(n8664) );
  XNOR U9610 ( .A(b[5]), .B(a[63]), .Z(n8606) );
  NANDN U9611 ( .A(n8606), .B(n36587), .Z(n8461) );
  NANDN U9612 ( .A(n8459), .B(n36588), .Z(n8460) );
  AND U9613 ( .A(n8461), .B(n8460), .Z(n8665) );
  XNOR U9614 ( .A(n8664), .B(n8665), .Z(n8666) );
  XNOR U9615 ( .A(n8667), .B(n8666), .Z(n8655) );
  NANDN U9616 ( .A(n8462), .B(n37762), .Z(n8464) );
  XOR U9617 ( .A(b[17]), .B(a[51]), .Z(n8609) );
  NAND U9618 ( .A(n8609), .B(n37764), .Z(n8463) );
  NAND U9619 ( .A(n8464), .B(n8463), .Z(n8627) );
  XOR U9620 ( .A(b[31]), .B(n8832), .Z(n8612) );
  NANDN U9621 ( .A(n8612), .B(n38552), .Z(n8467) );
  NANDN U9622 ( .A(n8465), .B(n38553), .Z(n8466) );
  NAND U9623 ( .A(n8467), .B(n8466), .Z(n8624) );
  OR U9624 ( .A(n8468), .B(n36105), .Z(n8470) );
  XNOR U9625 ( .A(b[3]), .B(a[65]), .Z(n8615) );
  NANDN U9626 ( .A(n8615), .B(n36107), .Z(n8469) );
  AND U9627 ( .A(n8470), .B(n8469), .Z(n8625) );
  XNOR U9628 ( .A(n8624), .B(n8625), .Z(n8626) );
  XOR U9629 ( .A(n8627), .B(n8626), .Z(n8654) );
  XNOR U9630 ( .A(n8655), .B(n8654), .Z(n8656) );
  XNOR U9631 ( .A(n8657), .B(n8656), .Z(n8700) );
  NANDN U9632 ( .A(n8472), .B(n8471), .Z(n8476) );
  NAND U9633 ( .A(n8474), .B(n8473), .Z(n8475) );
  NAND U9634 ( .A(n8476), .B(n8475), .Z(n8645) );
  NANDN U9635 ( .A(n8478), .B(n8477), .Z(n8482) );
  NAND U9636 ( .A(n8480), .B(n8479), .Z(n8481) );
  NAND U9637 ( .A(n8482), .B(n8481), .Z(n8643) );
  OR U9638 ( .A(n8484), .B(n8483), .Z(n8488) );
  NANDN U9639 ( .A(n8486), .B(n8485), .Z(n8487) );
  NAND U9640 ( .A(n8488), .B(n8487), .Z(n8642) );
  XNOR U9641 ( .A(n8645), .B(n8644), .Z(n8701) );
  XOR U9642 ( .A(n8700), .B(n8701), .Z(n8703) );
  NANDN U9643 ( .A(n8490), .B(n8489), .Z(n8494) );
  OR U9644 ( .A(n8492), .B(n8491), .Z(n8493) );
  NAND U9645 ( .A(n8494), .B(n8493), .Z(n8702) );
  XOR U9646 ( .A(n8703), .B(n8702), .Z(n8590) );
  OR U9647 ( .A(n8496), .B(n8495), .Z(n8500) );
  NAND U9648 ( .A(n8498), .B(n8497), .Z(n8499) );
  NAND U9649 ( .A(n8500), .B(n8499), .Z(n8589) );
  NANDN U9650 ( .A(n8502), .B(n8501), .Z(n8506) );
  NANDN U9651 ( .A(n8504), .B(n8503), .Z(n8505) );
  NAND U9652 ( .A(n8506), .B(n8505), .Z(n8708) );
  NANDN U9653 ( .A(n8512), .B(n8511), .Z(n8516) );
  NAND U9654 ( .A(n8514), .B(n8513), .Z(n8515) );
  NAND U9655 ( .A(n8516), .B(n8515), .Z(n8648) );
  NANDN U9656 ( .A(n8518), .B(n8517), .Z(n8522) );
  NAND U9657 ( .A(n8520), .B(n8519), .Z(n8521) );
  AND U9658 ( .A(n8522), .B(n8521), .Z(n8649) );
  XNOR U9659 ( .A(n8648), .B(n8649), .Z(n8650) );
  XOR U9660 ( .A(b[9]), .B(n12056), .Z(n8670) );
  NANDN U9661 ( .A(n8670), .B(n36925), .Z(n8525) );
  NANDN U9662 ( .A(n8523), .B(n36926), .Z(n8524) );
  NAND U9663 ( .A(n8525), .B(n8524), .Z(n8632) );
  XNOR U9664 ( .A(b[15]), .B(a[53]), .Z(n8673) );
  OR U9665 ( .A(n8673), .B(n37665), .Z(n8528) );
  NANDN U9666 ( .A(n8526), .B(n37604), .Z(n8527) );
  AND U9667 ( .A(n8528), .B(n8527), .Z(n8630) );
  XNOR U9668 ( .A(b[21]), .B(a[47]), .Z(n8676) );
  NANDN U9669 ( .A(n8676), .B(n38101), .Z(n8531) );
  NANDN U9670 ( .A(n8529), .B(n38102), .Z(n8530) );
  AND U9671 ( .A(n8531), .B(n8530), .Z(n8631) );
  XOR U9672 ( .A(n8632), .B(n8633), .Z(n8621) );
  XNOR U9673 ( .A(b[11]), .B(a[57]), .Z(n8679) );
  OR U9674 ( .A(n8679), .B(n37311), .Z(n8534) );
  NANDN U9675 ( .A(n8532), .B(n37218), .Z(n8533) );
  NAND U9676 ( .A(n8534), .B(n8533), .Z(n8619) );
  XOR U9677 ( .A(n1053), .B(a[55]), .Z(n8682) );
  NANDN U9678 ( .A(n8682), .B(n37424), .Z(n8537) );
  NANDN U9679 ( .A(n8535), .B(n37425), .Z(n8536) );
  AND U9680 ( .A(n8537), .B(n8536), .Z(n8618) );
  XNOR U9681 ( .A(n8619), .B(n8618), .Z(n8620) );
  XOR U9682 ( .A(n8621), .B(n8620), .Z(n8638) );
  NANDN U9683 ( .A(n1049), .B(a[67]), .Z(n8538) );
  XNOR U9684 ( .A(b[1]), .B(n8538), .Z(n8540) );
  NANDN U9685 ( .A(b[0]), .B(a[66]), .Z(n8539) );
  AND U9686 ( .A(n8540), .B(n8539), .Z(n8596) );
  NAND U9687 ( .A(n38490), .B(n8541), .Z(n8543) );
  XNOR U9688 ( .A(n1058), .B(a[39]), .Z(n8685) );
  NANDN U9689 ( .A(n1048), .B(n8685), .Z(n8542) );
  NAND U9690 ( .A(n8543), .B(n8542), .Z(n8594) );
  NANDN U9691 ( .A(n1059), .B(a[35]), .Z(n8595) );
  XNOR U9692 ( .A(n8594), .B(n8595), .Z(n8597) );
  XOR U9693 ( .A(n8596), .B(n8597), .Z(n8636) );
  NANDN U9694 ( .A(n8544), .B(n38205), .Z(n8546) );
  XNOR U9695 ( .A(b[23]), .B(a[45]), .Z(n8691) );
  OR U9696 ( .A(n8691), .B(n38268), .Z(n8545) );
  NAND U9697 ( .A(n8546), .B(n8545), .Z(n8661) );
  XOR U9698 ( .A(b[7]), .B(a[61]), .Z(n8694) );
  NAND U9699 ( .A(n8694), .B(n36701), .Z(n8549) );
  NAND U9700 ( .A(n8547), .B(n36702), .Z(n8548) );
  NAND U9701 ( .A(n8549), .B(n8548), .Z(n8658) );
  XOR U9702 ( .A(b[25]), .B(a[43]), .Z(n8697) );
  NAND U9703 ( .A(n8697), .B(n38325), .Z(n8552) );
  NAND U9704 ( .A(n8550), .B(n38326), .Z(n8551) );
  AND U9705 ( .A(n8552), .B(n8551), .Z(n8659) );
  XNOR U9706 ( .A(n8658), .B(n8659), .Z(n8660) );
  XNOR U9707 ( .A(n8661), .B(n8660), .Z(n8637) );
  XOR U9708 ( .A(n8636), .B(n8637), .Z(n8639) );
  XNOR U9709 ( .A(n8638), .B(n8639), .Z(n8651) );
  XNOR U9710 ( .A(n8650), .B(n8651), .Z(n8706) );
  XNOR U9711 ( .A(n8707), .B(n8706), .Z(n8709) );
  XNOR U9712 ( .A(n8708), .B(n8709), .Z(n8588) );
  XOR U9713 ( .A(n8589), .B(n8588), .Z(n8591) );
  NANDN U9714 ( .A(n8554), .B(n8553), .Z(n8558) );
  NAND U9715 ( .A(n8556), .B(n8555), .Z(n8557) );
  NAND U9716 ( .A(n8558), .B(n8557), .Z(n8582) );
  NAND U9717 ( .A(n8560), .B(n8559), .Z(n8564) );
  OR U9718 ( .A(n8562), .B(n8561), .Z(n8563) );
  NAND U9719 ( .A(n8564), .B(n8563), .Z(n8583) );
  XNOR U9720 ( .A(n8582), .B(n8583), .Z(n8584) );
  XOR U9721 ( .A(n8585), .B(n8584), .Z(n8579) );
  XOR U9722 ( .A(n8578), .B(n8579), .Z(n8570) );
  XOR U9723 ( .A(n8571), .B(n8570), .Z(n8572) );
  XNOR U9724 ( .A(n8573), .B(n8572), .Z(n8712) );
  XNOR U9725 ( .A(n8712), .B(sreg[291]), .Z(n8714) );
  NAND U9726 ( .A(n8565), .B(sreg[290]), .Z(n8569) );
  OR U9727 ( .A(n8567), .B(n8566), .Z(n8568) );
  AND U9728 ( .A(n8569), .B(n8568), .Z(n8713) );
  XOR U9729 ( .A(n8714), .B(n8713), .Z(c[291]) );
  NAND U9730 ( .A(n8571), .B(n8570), .Z(n8575) );
  NAND U9731 ( .A(n8573), .B(n8572), .Z(n8574) );
  NAND U9732 ( .A(n8575), .B(n8574), .Z(n8720) );
  NANDN U9733 ( .A(n8577), .B(n8576), .Z(n8581) );
  NAND U9734 ( .A(n8579), .B(n8578), .Z(n8580) );
  NAND U9735 ( .A(n8581), .B(n8580), .Z(n8718) );
  NANDN U9736 ( .A(n8583), .B(n8582), .Z(n8587) );
  NAND U9737 ( .A(n8585), .B(n8584), .Z(n8586) );
  NAND U9738 ( .A(n8587), .B(n8586), .Z(n8723) );
  NANDN U9739 ( .A(n8589), .B(n8588), .Z(n8593) );
  OR U9740 ( .A(n8591), .B(n8590), .Z(n8592) );
  NAND U9741 ( .A(n8593), .B(n8592), .Z(n8724) );
  XNOR U9742 ( .A(n8723), .B(n8724), .Z(n8725) );
  NANDN U9743 ( .A(n8595), .B(n8594), .Z(n8599) );
  NAND U9744 ( .A(n8597), .B(n8596), .Z(n8598) );
  NAND U9745 ( .A(n8599), .B(n8598), .Z(n8804) );
  XOR U9746 ( .A(b[19]), .B(n10724), .Z(n8747) );
  NANDN U9747 ( .A(n8747), .B(n37934), .Z(n8602) );
  NANDN U9748 ( .A(n8600), .B(n37935), .Z(n8601) );
  NAND U9749 ( .A(n8602), .B(n8601), .Z(n8814) );
  XOR U9750 ( .A(b[27]), .B(a[42]), .Z(n8750) );
  NAND U9751 ( .A(n38423), .B(n8750), .Z(n8605) );
  NAND U9752 ( .A(n8603), .B(n38424), .Z(n8604) );
  NAND U9753 ( .A(n8605), .B(n8604), .Z(n8811) );
  XNOR U9754 ( .A(b[5]), .B(a[64]), .Z(n8753) );
  NANDN U9755 ( .A(n8753), .B(n36587), .Z(n8608) );
  NANDN U9756 ( .A(n8606), .B(n36588), .Z(n8607) );
  AND U9757 ( .A(n8608), .B(n8607), .Z(n8812) );
  XNOR U9758 ( .A(n8811), .B(n8812), .Z(n8813) );
  XNOR U9759 ( .A(n8814), .B(n8813), .Z(n8802) );
  NAND U9760 ( .A(n8609), .B(n37762), .Z(n8611) );
  XOR U9761 ( .A(b[17]), .B(a[52]), .Z(n8756) );
  NAND U9762 ( .A(n8756), .B(n37764), .Z(n8610) );
  NAND U9763 ( .A(n8611), .B(n8610), .Z(n8774) );
  XNOR U9764 ( .A(b[31]), .B(a[38]), .Z(n8759) );
  NANDN U9765 ( .A(n8759), .B(n38552), .Z(n8614) );
  NANDN U9766 ( .A(n8612), .B(n38553), .Z(n8613) );
  NAND U9767 ( .A(n8614), .B(n8613), .Z(n8771) );
  OR U9768 ( .A(n8615), .B(n36105), .Z(n8617) );
  XNOR U9769 ( .A(b[3]), .B(a[66]), .Z(n8762) );
  NANDN U9770 ( .A(n8762), .B(n36107), .Z(n8616) );
  AND U9771 ( .A(n8617), .B(n8616), .Z(n8772) );
  XNOR U9772 ( .A(n8771), .B(n8772), .Z(n8773) );
  XOR U9773 ( .A(n8774), .B(n8773), .Z(n8801) );
  XNOR U9774 ( .A(n8802), .B(n8801), .Z(n8803) );
  XNOR U9775 ( .A(n8804), .B(n8803), .Z(n8848) );
  NANDN U9776 ( .A(n8619), .B(n8618), .Z(n8623) );
  NAND U9777 ( .A(n8621), .B(n8620), .Z(n8622) );
  NAND U9778 ( .A(n8623), .B(n8622), .Z(n8792) );
  NANDN U9779 ( .A(n8625), .B(n8624), .Z(n8629) );
  NAND U9780 ( .A(n8627), .B(n8626), .Z(n8628) );
  NAND U9781 ( .A(n8629), .B(n8628), .Z(n8790) );
  OR U9782 ( .A(n8631), .B(n8630), .Z(n8635) );
  NANDN U9783 ( .A(n8633), .B(n8632), .Z(n8634) );
  NAND U9784 ( .A(n8635), .B(n8634), .Z(n8789) );
  XNOR U9785 ( .A(n8792), .B(n8791), .Z(n8849) );
  XOR U9786 ( .A(n8848), .B(n8849), .Z(n8851) );
  NANDN U9787 ( .A(n8637), .B(n8636), .Z(n8641) );
  OR U9788 ( .A(n8639), .B(n8638), .Z(n8640) );
  NAND U9789 ( .A(n8641), .B(n8640), .Z(n8850) );
  XOR U9790 ( .A(n8851), .B(n8850), .Z(n8737) );
  OR U9791 ( .A(n8643), .B(n8642), .Z(n8647) );
  NAND U9792 ( .A(n8645), .B(n8644), .Z(n8646) );
  NAND U9793 ( .A(n8647), .B(n8646), .Z(n8736) );
  NANDN U9794 ( .A(n8649), .B(n8648), .Z(n8653) );
  NANDN U9795 ( .A(n8651), .B(n8650), .Z(n8652) );
  NAND U9796 ( .A(n8653), .B(n8652), .Z(n8856) );
  NANDN U9797 ( .A(n8659), .B(n8658), .Z(n8663) );
  NAND U9798 ( .A(n8661), .B(n8660), .Z(n8662) );
  NAND U9799 ( .A(n8663), .B(n8662), .Z(n8795) );
  NANDN U9800 ( .A(n8665), .B(n8664), .Z(n8669) );
  NAND U9801 ( .A(n8667), .B(n8666), .Z(n8668) );
  AND U9802 ( .A(n8669), .B(n8668), .Z(n8796) );
  XNOR U9803 ( .A(n8795), .B(n8796), .Z(n8797) );
  XNOR U9804 ( .A(b[9]), .B(a[60]), .Z(n8817) );
  NANDN U9805 ( .A(n8817), .B(n36925), .Z(n8672) );
  NANDN U9806 ( .A(n8670), .B(n36926), .Z(n8671) );
  NAND U9807 ( .A(n8672), .B(n8671), .Z(n8779) );
  XOR U9808 ( .A(b[15]), .B(n11319), .Z(n8820) );
  OR U9809 ( .A(n8820), .B(n37665), .Z(n8675) );
  NANDN U9810 ( .A(n8673), .B(n37604), .Z(n8674) );
  AND U9811 ( .A(n8675), .B(n8674), .Z(n8777) );
  XNOR U9812 ( .A(b[21]), .B(a[48]), .Z(n8823) );
  NANDN U9813 ( .A(n8823), .B(n38101), .Z(n8678) );
  NANDN U9814 ( .A(n8676), .B(n38102), .Z(n8677) );
  AND U9815 ( .A(n8678), .B(n8677), .Z(n8778) );
  XOR U9816 ( .A(n8779), .B(n8780), .Z(n8768) );
  XNOR U9817 ( .A(b[11]), .B(a[58]), .Z(n8826) );
  OR U9818 ( .A(n8826), .B(n37311), .Z(n8681) );
  NANDN U9819 ( .A(n8679), .B(n37218), .Z(n8680) );
  NAND U9820 ( .A(n8681), .B(n8680), .Z(n8766) );
  XOR U9821 ( .A(n1053), .B(a[56]), .Z(n8829) );
  NANDN U9822 ( .A(n8829), .B(n37424), .Z(n8684) );
  NANDN U9823 ( .A(n8682), .B(n37425), .Z(n8683) );
  AND U9824 ( .A(n8684), .B(n8683), .Z(n8765) );
  XNOR U9825 ( .A(n8766), .B(n8765), .Z(n8767) );
  XOR U9826 ( .A(n8768), .B(n8767), .Z(n8785) );
  NAND U9827 ( .A(n38490), .B(n8685), .Z(n8687) );
  XNOR U9828 ( .A(b[29]), .B(a[40]), .Z(n8833) );
  OR U9829 ( .A(n8833), .B(n1048), .Z(n8686) );
  NAND U9830 ( .A(n8687), .B(n8686), .Z(n8741) );
  NANDN U9831 ( .A(n1059), .B(a[36]), .Z(n8742) );
  XNOR U9832 ( .A(n8741), .B(n8742), .Z(n8744) );
  NANDN U9833 ( .A(n1049), .B(a[68]), .Z(n8688) );
  XNOR U9834 ( .A(b[1]), .B(n8688), .Z(n8690) );
  IV U9835 ( .A(a[67]), .Z(n13219) );
  NANDN U9836 ( .A(n13219), .B(n1049), .Z(n8689) );
  AND U9837 ( .A(n8690), .B(n8689), .Z(n8743) );
  XOR U9838 ( .A(n8744), .B(n8743), .Z(n8783) );
  NANDN U9839 ( .A(n8691), .B(n38205), .Z(n8693) );
  XNOR U9840 ( .A(b[23]), .B(a[46]), .Z(n8839) );
  OR U9841 ( .A(n8839), .B(n38268), .Z(n8692) );
  NAND U9842 ( .A(n8693), .B(n8692), .Z(n8808) );
  XNOR U9843 ( .A(b[7]), .B(a[62]), .Z(n8842) );
  NANDN U9844 ( .A(n8842), .B(n36701), .Z(n8696) );
  NAND U9845 ( .A(n8694), .B(n36702), .Z(n8695) );
  NAND U9846 ( .A(n8696), .B(n8695), .Z(n8805) );
  XNOR U9847 ( .A(b[25]), .B(a[44]), .Z(n8845) );
  NANDN U9848 ( .A(n8845), .B(n38325), .Z(n8699) );
  NAND U9849 ( .A(n8697), .B(n38326), .Z(n8698) );
  AND U9850 ( .A(n8699), .B(n8698), .Z(n8806) );
  XNOR U9851 ( .A(n8805), .B(n8806), .Z(n8807) );
  XNOR U9852 ( .A(n8808), .B(n8807), .Z(n8784) );
  XOR U9853 ( .A(n8783), .B(n8784), .Z(n8786) );
  XNOR U9854 ( .A(n8785), .B(n8786), .Z(n8798) );
  XNOR U9855 ( .A(n8797), .B(n8798), .Z(n8854) );
  XNOR U9856 ( .A(n8855), .B(n8854), .Z(n8857) );
  XNOR U9857 ( .A(n8856), .B(n8857), .Z(n8735) );
  XOR U9858 ( .A(n8736), .B(n8735), .Z(n8738) );
  NANDN U9859 ( .A(n8701), .B(n8700), .Z(n8705) );
  OR U9860 ( .A(n8703), .B(n8702), .Z(n8704) );
  NAND U9861 ( .A(n8705), .B(n8704), .Z(n8729) );
  NAND U9862 ( .A(n8707), .B(n8706), .Z(n8711) );
  NANDN U9863 ( .A(n8709), .B(n8708), .Z(n8710) );
  NAND U9864 ( .A(n8711), .B(n8710), .Z(n8730) );
  XNOR U9865 ( .A(n8729), .B(n8730), .Z(n8731) );
  XOR U9866 ( .A(n8732), .B(n8731), .Z(n8726) );
  XOR U9867 ( .A(n8725), .B(n8726), .Z(n8717) );
  XOR U9868 ( .A(n8718), .B(n8717), .Z(n8719) );
  XNOR U9869 ( .A(n8720), .B(n8719), .Z(n8860) );
  XNOR U9870 ( .A(n8860), .B(sreg[292]), .Z(n8862) );
  NAND U9871 ( .A(n8712), .B(sreg[291]), .Z(n8716) );
  OR U9872 ( .A(n8714), .B(n8713), .Z(n8715) );
  AND U9873 ( .A(n8716), .B(n8715), .Z(n8861) );
  XOR U9874 ( .A(n8862), .B(n8861), .Z(c[292]) );
  NAND U9875 ( .A(n8718), .B(n8717), .Z(n8722) );
  NAND U9876 ( .A(n8720), .B(n8719), .Z(n8721) );
  NAND U9877 ( .A(n8722), .B(n8721), .Z(n8868) );
  NANDN U9878 ( .A(n8724), .B(n8723), .Z(n8728) );
  NAND U9879 ( .A(n8726), .B(n8725), .Z(n8727) );
  NAND U9880 ( .A(n8728), .B(n8727), .Z(n8866) );
  NANDN U9881 ( .A(n8730), .B(n8729), .Z(n8734) );
  NAND U9882 ( .A(n8732), .B(n8731), .Z(n8733) );
  NAND U9883 ( .A(n8734), .B(n8733), .Z(n8871) );
  NANDN U9884 ( .A(n8736), .B(n8735), .Z(n8740) );
  OR U9885 ( .A(n8738), .B(n8737), .Z(n8739) );
  NAND U9886 ( .A(n8740), .B(n8739), .Z(n8872) );
  XNOR U9887 ( .A(n8871), .B(n8872), .Z(n8873) );
  NANDN U9888 ( .A(n8742), .B(n8741), .Z(n8746) );
  NAND U9889 ( .A(n8744), .B(n8743), .Z(n8745) );
  NAND U9890 ( .A(n8746), .B(n8745), .Z(n8952) );
  XNOR U9891 ( .A(b[19]), .B(a[51]), .Z(n8919) );
  NANDN U9892 ( .A(n8919), .B(n37934), .Z(n8749) );
  NANDN U9893 ( .A(n8747), .B(n37935), .Z(n8748) );
  NAND U9894 ( .A(n8749), .B(n8748), .Z(n8988) );
  XOR U9895 ( .A(b[27]), .B(a[43]), .Z(n8922) );
  NAND U9896 ( .A(n38423), .B(n8922), .Z(n8752) );
  NAND U9897 ( .A(n8750), .B(n38424), .Z(n8751) );
  NAND U9898 ( .A(n8752), .B(n8751), .Z(n8985) );
  XNOR U9899 ( .A(b[5]), .B(a[65]), .Z(n8925) );
  NANDN U9900 ( .A(n8925), .B(n36587), .Z(n8755) );
  NANDN U9901 ( .A(n8753), .B(n36588), .Z(n8754) );
  AND U9902 ( .A(n8755), .B(n8754), .Z(n8986) );
  XNOR U9903 ( .A(n8985), .B(n8986), .Z(n8987) );
  XNOR U9904 ( .A(n8988), .B(n8987), .Z(n8949) );
  NAND U9905 ( .A(n8756), .B(n37762), .Z(n8758) );
  XOR U9906 ( .A(b[17]), .B(a[53]), .Z(n8928) );
  NAND U9907 ( .A(n8928), .B(n37764), .Z(n8757) );
  NAND U9908 ( .A(n8758), .B(n8757), .Z(n8903) );
  XNOR U9909 ( .A(b[31]), .B(a[39]), .Z(n8931) );
  NANDN U9910 ( .A(n8931), .B(n38552), .Z(n8761) );
  NANDN U9911 ( .A(n8759), .B(n38553), .Z(n8760) );
  AND U9912 ( .A(n8761), .B(n8760), .Z(n8901) );
  OR U9913 ( .A(n8762), .B(n36105), .Z(n8764) );
  XOR U9914 ( .A(b[3]), .B(n13219), .Z(n8934) );
  NANDN U9915 ( .A(n8934), .B(n36107), .Z(n8763) );
  AND U9916 ( .A(n8764), .B(n8763), .Z(n8902) );
  XOR U9917 ( .A(n8903), .B(n8904), .Z(n8950) );
  XOR U9918 ( .A(n8949), .B(n8950), .Z(n8951) );
  XNOR U9919 ( .A(n8952), .B(n8951), .Z(n8997) );
  NANDN U9920 ( .A(n8766), .B(n8765), .Z(n8770) );
  NAND U9921 ( .A(n8768), .B(n8767), .Z(n8769) );
  NAND U9922 ( .A(n8770), .B(n8769), .Z(n8940) );
  NANDN U9923 ( .A(n8772), .B(n8771), .Z(n8776) );
  NAND U9924 ( .A(n8774), .B(n8773), .Z(n8775) );
  NAND U9925 ( .A(n8776), .B(n8775), .Z(n8938) );
  OR U9926 ( .A(n8778), .B(n8777), .Z(n8782) );
  NANDN U9927 ( .A(n8780), .B(n8779), .Z(n8781) );
  NAND U9928 ( .A(n8782), .B(n8781), .Z(n8937) );
  XNOR U9929 ( .A(n8940), .B(n8939), .Z(n8998) );
  XOR U9930 ( .A(n8997), .B(n8998), .Z(n9000) );
  NANDN U9931 ( .A(n8784), .B(n8783), .Z(n8788) );
  OR U9932 ( .A(n8786), .B(n8785), .Z(n8787) );
  NAND U9933 ( .A(n8788), .B(n8787), .Z(n8999) );
  XOR U9934 ( .A(n9000), .B(n8999), .Z(n8885) );
  OR U9935 ( .A(n8790), .B(n8789), .Z(n8794) );
  NAND U9936 ( .A(n8792), .B(n8791), .Z(n8793) );
  NAND U9937 ( .A(n8794), .B(n8793), .Z(n8884) );
  NANDN U9938 ( .A(n8796), .B(n8795), .Z(n8800) );
  NANDN U9939 ( .A(n8798), .B(n8797), .Z(n8799) );
  NAND U9940 ( .A(n8800), .B(n8799), .Z(n9005) );
  NANDN U9941 ( .A(n8806), .B(n8805), .Z(n8810) );
  NAND U9942 ( .A(n8808), .B(n8807), .Z(n8809) );
  NAND U9943 ( .A(n8810), .B(n8809), .Z(n8943) );
  NANDN U9944 ( .A(n8812), .B(n8811), .Z(n8816) );
  NAND U9945 ( .A(n8814), .B(n8813), .Z(n8815) );
  AND U9946 ( .A(n8816), .B(n8815), .Z(n8944) );
  XNOR U9947 ( .A(n8943), .B(n8944), .Z(n8945) );
  XNOR U9948 ( .A(b[9]), .B(a[61]), .Z(n8955) );
  NANDN U9949 ( .A(n8955), .B(n36925), .Z(n8819) );
  NANDN U9950 ( .A(n8817), .B(n36926), .Z(n8818) );
  NAND U9951 ( .A(n8819), .B(n8818), .Z(n8909) );
  XNOR U9952 ( .A(b[15]), .B(a[55]), .Z(n8958) );
  OR U9953 ( .A(n8958), .B(n37665), .Z(n8822) );
  NANDN U9954 ( .A(n8820), .B(n37604), .Z(n8821) );
  AND U9955 ( .A(n8822), .B(n8821), .Z(n8907) );
  XNOR U9956 ( .A(b[21]), .B(a[49]), .Z(n8961) );
  NANDN U9957 ( .A(n8961), .B(n38101), .Z(n8825) );
  NANDN U9958 ( .A(n8823), .B(n38102), .Z(n8824) );
  AND U9959 ( .A(n8825), .B(n8824), .Z(n8908) );
  XOR U9960 ( .A(n8909), .B(n8910), .Z(n8898) );
  XOR U9961 ( .A(b[11]), .B(n12056), .Z(n8964) );
  OR U9962 ( .A(n8964), .B(n37311), .Z(n8828) );
  NANDN U9963 ( .A(n8826), .B(n37218), .Z(n8827) );
  NAND U9964 ( .A(n8828), .B(n8827), .Z(n8896) );
  XOR U9965 ( .A(n1053), .B(a[57]), .Z(n8967) );
  NANDN U9966 ( .A(n8967), .B(n37424), .Z(n8831) );
  NANDN U9967 ( .A(n8829), .B(n37425), .Z(n8830) );
  NAND U9968 ( .A(n8831), .B(n8830), .Z(n8895) );
  XOR U9969 ( .A(n8898), .B(n8897), .Z(n8892) );
  ANDN U9970 ( .B(b[31]), .A(n8832), .Z(n8913) );
  NANDN U9971 ( .A(n8833), .B(n38490), .Z(n8835) );
  XNOR U9972 ( .A(n1058), .B(a[41]), .Z(n8973) );
  NANDN U9973 ( .A(n1048), .B(n8973), .Z(n8834) );
  NAND U9974 ( .A(n8835), .B(n8834), .Z(n8914) );
  XOR U9975 ( .A(n8913), .B(n8914), .Z(n8915) );
  NANDN U9976 ( .A(n1049), .B(a[69]), .Z(n8836) );
  XNOR U9977 ( .A(b[1]), .B(n8836), .Z(n8838) );
  NANDN U9978 ( .A(b[0]), .B(a[68]), .Z(n8837) );
  AND U9979 ( .A(n8838), .B(n8837), .Z(n8916) );
  XNOR U9980 ( .A(n8915), .B(n8916), .Z(n8889) );
  NANDN U9981 ( .A(n8839), .B(n38205), .Z(n8841) );
  XNOR U9982 ( .A(b[23]), .B(a[47]), .Z(n8976) );
  OR U9983 ( .A(n8976), .B(n38268), .Z(n8840) );
  NAND U9984 ( .A(n8841), .B(n8840), .Z(n8994) );
  XOR U9985 ( .A(b[7]), .B(a[63]), .Z(n8979) );
  NAND U9986 ( .A(n8979), .B(n36701), .Z(n8844) );
  NANDN U9987 ( .A(n8842), .B(n36702), .Z(n8843) );
  NAND U9988 ( .A(n8844), .B(n8843), .Z(n8991) );
  XOR U9989 ( .A(b[25]), .B(a[45]), .Z(n8982) );
  NAND U9990 ( .A(n8982), .B(n38325), .Z(n8847) );
  NANDN U9991 ( .A(n8845), .B(n38326), .Z(n8846) );
  AND U9992 ( .A(n8847), .B(n8846), .Z(n8992) );
  XNOR U9993 ( .A(n8991), .B(n8992), .Z(n8993) );
  XNOR U9994 ( .A(n8994), .B(n8993), .Z(n8890) );
  XOR U9995 ( .A(n8892), .B(n8891), .Z(n8946) );
  XNOR U9996 ( .A(n8945), .B(n8946), .Z(n9003) );
  XNOR U9997 ( .A(n9004), .B(n9003), .Z(n9006) );
  XNOR U9998 ( .A(n9005), .B(n9006), .Z(n8883) );
  XOR U9999 ( .A(n8884), .B(n8883), .Z(n8886) );
  NANDN U10000 ( .A(n8849), .B(n8848), .Z(n8853) );
  OR U10001 ( .A(n8851), .B(n8850), .Z(n8852) );
  NAND U10002 ( .A(n8853), .B(n8852), .Z(n8877) );
  NAND U10003 ( .A(n8855), .B(n8854), .Z(n8859) );
  NANDN U10004 ( .A(n8857), .B(n8856), .Z(n8858) );
  NAND U10005 ( .A(n8859), .B(n8858), .Z(n8878) );
  XNOR U10006 ( .A(n8877), .B(n8878), .Z(n8879) );
  XOR U10007 ( .A(n8880), .B(n8879), .Z(n8874) );
  XOR U10008 ( .A(n8873), .B(n8874), .Z(n8865) );
  XOR U10009 ( .A(n8866), .B(n8865), .Z(n8867) );
  XNOR U10010 ( .A(n8868), .B(n8867), .Z(n9009) );
  XNOR U10011 ( .A(n9009), .B(sreg[293]), .Z(n9011) );
  NAND U10012 ( .A(n8860), .B(sreg[292]), .Z(n8864) );
  OR U10013 ( .A(n8862), .B(n8861), .Z(n8863) );
  AND U10014 ( .A(n8864), .B(n8863), .Z(n9010) );
  XOR U10015 ( .A(n9011), .B(n9010), .Z(c[293]) );
  NAND U10016 ( .A(n8866), .B(n8865), .Z(n8870) );
  NAND U10017 ( .A(n8868), .B(n8867), .Z(n8869) );
  NAND U10018 ( .A(n8870), .B(n8869), .Z(n9017) );
  NANDN U10019 ( .A(n8872), .B(n8871), .Z(n8876) );
  NAND U10020 ( .A(n8874), .B(n8873), .Z(n8875) );
  NAND U10021 ( .A(n8876), .B(n8875), .Z(n9015) );
  NANDN U10022 ( .A(n8878), .B(n8877), .Z(n8882) );
  NAND U10023 ( .A(n8880), .B(n8879), .Z(n8881) );
  NAND U10024 ( .A(n8882), .B(n8881), .Z(n9020) );
  NANDN U10025 ( .A(n8884), .B(n8883), .Z(n8888) );
  OR U10026 ( .A(n8886), .B(n8885), .Z(n8887) );
  NAND U10027 ( .A(n8888), .B(n8887), .Z(n9021) );
  XNOR U10028 ( .A(n9020), .B(n9021), .Z(n9022) );
  OR U10029 ( .A(n8890), .B(n8889), .Z(n8894) );
  NANDN U10030 ( .A(n8892), .B(n8891), .Z(n8893) );
  NAND U10031 ( .A(n8894), .B(n8893), .Z(n9137) );
  OR U10032 ( .A(n8896), .B(n8895), .Z(n8900) );
  NAND U10033 ( .A(n8898), .B(n8897), .Z(n8899) );
  NAND U10034 ( .A(n8900), .B(n8899), .Z(n9076) );
  OR U10035 ( .A(n8902), .B(n8901), .Z(n8906) );
  NANDN U10036 ( .A(n8904), .B(n8903), .Z(n8905) );
  NAND U10037 ( .A(n8906), .B(n8905), .Z(n9075) );
  OR U10038 ( .A(n8908), .B(n8907), .Z(n8912) );
  NANDN U10039 ( .A(n8910), .B(n8909), .Z(n8911) );
  NAND U10040 ( .A(n8912), .B(n8911), .Z(n9074) );
  XOR U10041 ( .A(n9076), .B(n9077), .Z(n9135) );
  OR U10042 ( .A(n8914), .B(n8913), .Z(n8918) );
  NANDN U10043 ( .A(n8916), .B(n8915), .Z(n8917) );
  NAND U10044 ( .A(n8918), .B(n8917), .Z(n9088) );
  XNOR U10045 ( .A(b[19]), .B(a[52]), .Z(n9032) );
  NANDN U10046 ( .A(n9032), .B(n37934), .Z(n8921) );
  NANDN U10047 ( .A(n8919), .B(n37935), .Z(n8920) );
  NAND U10048 ( .A(n8921), .B(n8920), .Z(n9101) );
  XNOR U10049 ( .A(b[27]), .B(a[44]), .Z(n9035) );
  NANDN U10050 ( .A(n9035), .B(n38423), .Z(n8924) );
  NAND U10051 ( .A(n8922), .B(n38424), .Z(n8923) );
  NAND U10052 ( .A(n8924), .B(n8923), .Z(n9098) );
  XNOR U10053 ( .A(b[5]), .B(a[66]), .Z(n9038) );
  NANDN U10054 ( .A(n9038), .B(n36587), .Z(n8927) );
  NANDN U10055 ( .A(n8925), .B(n36588), .Z(n8926) );
  AND U10056 ( .A(n8927), .B(n8926), .Z(n9099) );
  XNOR U10057 ( .A(n9098), .B(n9099), .Z(n9100) );
  XNOR U10058 ( .A(n9101), .B(n9100), .Z(n9087) );
  NAND U10059 ( .A(n8928), .B(n37762), .Z(n8930) );
  XNOR U10060 ( .A(b[17]), .B(a[54]), .Z(n9041) );
  NANDN U10061 ( .A(n9041), .B(n37764), .Z(n8929) );
  NAND U10062 ( .A(n8930), .B(n8929), .Z(n9059) );
  XNOR U10063 ( .A(b[31]), .B(a[40]), .Z(n9044) );
  NANDN U10064 ( .A(n9044), .B(n38552), .Z(n8933) );
  NANDN U10065 ( .A(n8931), .B(n38553), .Z(n8932) );
  NAND U10066 ( .A(n8933), .B(n8932), .Z(n9056) );
  OR U10067 ( .A(n8934), .B(n36105), .Z(n8936) );
  XNOR U10068 ( .A(b[3]), .B(a[68]), .Z(n9047) );
  NANDN U10069 ( .A(n9047), .B(n36107), .Z(n8935) );
  AND U10070 ( .A(n8936), .B(n8935), .Z(n9057) );
  XNOR U10071 ( .A(n9056), .B(n9057), .Z(n9058) );
  XOR U10072 ( .A(n9059), .B(n9058), .Z(n9086) );
  XOR U10073 ( .A(n9087), .B(n9086), .Z(n9089) );
  XOR U10074 ( .A(n9088), .B(n9089), .Z(n9134) );
  XOR U10075 ( .A(n9135), .B(n9134), .Z(n9136) );
  XNOR U10076 ( .A(n9137), .B(n9136), .Z(n9155) );
  OR U10077 ( .A(n8938), .B(n8937), .Z(n8942) );
  NAND U10078 ( .A(n8940), .B(n8939), .Z(n8941) );
  NAND U10079 ( .A(n8942), .B(n8941), .Z(n9153) );
  NANDN U10080 ( .A(n8944), .B(n8943), .Z(n8948) );
  NANDN U10081 ( .A(n8946), .B(n8945), .Z(n8947) );
  NAND U10082 ( .A(n8948), .B(n8947), .Z(n9143) );
  OR U10083 ( .A(n8950), .B(n8949), .Z(n8954) );
  NAND U10084 ( .A(n8952), .B(n8951), .Z(n8953) );
  NAND U10085 ( .A(n8954), .B(n8953), .Z(n9140) );
  XOR U10086 ( .A(b[9]), .B(n12493), .Z(n9104) );
  NANDN U10087 ( .A(n9104), .B(n36925), .Z(n8957) );
  NANDN U10088 ( .A(n8955), .B(n36926), .Z(n8956) );
  NAND U10089 ( .A(n8957), .B(n8956), .Z(n9064) );
  XNOR U10090 ( .A(b[15]), .B(a[56]), .Z(n9107) );
  OR U10091 ( .A(n9107), .B(n37665), .Z(n8960) );
  NANDN U10092 ( .A(n8958), .B(n37604), .Z(n8959) );
  AND U10093 ( .A(n8960), .B(n8959), .Z(n9062) );
  XOR U10094 ( .A(b[21]), .B(n10724), .Z(n9110) );
  NANDN U10095 ( .A(n9110), .B(n38101), .Z(n8963) );
  NANDN U10096 ( .A(n8961), .B(n38102), .Z(n8962) );
  AND U10097 ( .A(n8963), .B(n8962), .Z(n9063) );
  XOR U10098 ( .A(n9064), .B(n9065), .Z(n9053) );
  XNOR U10099 ( .A(b[11]), .B(a[60]), .Z(n9113) );
  OR U10100 ( .A(n9113), .B(n37311), .Z(n8966) );
  NANDN U10101 ( .A(n8964), .B(n37218), .Z(n8965) );
  NAND U10102 ( .A(n8966), .B(n8965), .Z(n9051) );
  XOR U10103 ( .A(n1053), .B(a[58]), .Z(n9116) );
  NANDN U10104 ( .A(n9116), .B(n37424), .Z(n8969) );
  NANDN U10105 ( .A(n8967), .B(n37425), .Z(n8968) );
  AND U10106 ( .A(n8969), .B(n8968), .Z(n9050) );
  XNOR U10107 ( .A(n9051), .B(n9050), .Z(n9052) );
  XOR U10108 ( .A(n9053), .B(n9052), .Z(n9071) );
  NANDN U10109 ( .A(n1049), .B(a[70]), .Z(n8970) );
  XNOR U10110 ( .A(b[1]), .B(n8970), .Z(n8972) );
  NANDN U10111 ( .A(b[0]), .B(a[69]), .Z(n8971) );
  AND U10112 ( .A(n8972), .B(n8971), .Z(n9028) );
  NAND U10113 ( .A(n8973), .B(n38490), .Z(n8975) );
  XNOR U10114 ( .A(n1058), .B(a[42]), .Z(n9122) );
  NANDN U10115 ( .A(n1048), .B(n9122), .Z(n8974) );
  NAND U10116 ( .A(n8975), .B(n8974), .Z(n9026) );
  NANDN U10117 ( .A(n1059), .B(a[38]), .Z(n9027) );
  XNOR U10118 ( .A(n9026), .B(n9027), .Z(n9029) );
  XOR U10119 ( .A(n9028), .B(n9029), .Z(n9068) );
  NANDN U10120 ( .A(n8976), .B(n38205), .Z(n8978) );
  XNOR U10121 ( .A(b[23]), .B(a[48]), .Z(n9125) );
  OR U10122 ( .A(n9125), .B(n38268), .Z(n8977) );
  NAND U10123 ( .A(n8978), .B(n8977), .Z(n9095) );
  XOR U10124 ( .A(b[7]), .B(a[64]), .Z(n9128) );
  NAND U10125 ( .A(n9128), .B(n36701), .Z(n8981) );
  NAND U10126 ( .A(n8979), .B(n36702), .Z(n8980) );
  NAND U10127 ( .A(n8981), .B(n8980), .Z(n9092) );
  XOR U10128 ( .A(b[25]), .B(a[46]), .Z(n9131) );
  NAND U10129 ( .A(n9131), .B(n38325), .Z(n8984) );
  NAND U10130 ( .A(n8982), .B(n38326), .Z(n8983) );
  AND U10131 ( .A(n8984), .B(n8983), .Z(n9093) );
  XNOR U10132 ( .A(n9092), .B(n9093), .Z(n9094) );
  XNOR U10133 ( .A(n9095), .B(n9094), .Z(n9069) );
  XNOR U10134 ( .A(n9068), .B(n9069), .Z(n9070) );
  XNOR U10135 ( .A(n9071), .B(n9070), .Z(n9083) );
  NANDN U10136 ( .A(n8986), .B(n8985), .Z(n8990) );
  NAND U10137 ( .A(n8988), .B(n8987), .Z(n8989) );
  NAND U10138 ( .A(n8990), .B(n8989), .Z(n9081) );
  NANDN U10139 ( .A(n8992), .B(n8991), .Z(n8996) );
  NAND U10140 ( .A(n8994), .B(n8993), .Z(n8995) );
  AND U10141 ( .A(n8996), .B(n8995), .Z(n9080) );
  XNOR U10142 ( .A(n9081), .B(n9080), .Z(n9082) );
  XNOR U10143 ( .A(n9083), .B(n9082), .Z(n9141) );
  XNOR U10144 ( .A(n9140), .B(n9141), .Z(n9142) );
  XOR U10145 ( .A(n9143), .B(n9142), .Z(n9152) );
  XNOR U10146 ( .A(n9153), .B(n9152), .Z(n9154) );
  XOR U10147 ( .A(n9155), .B(n9154), .Z(n9149) );
  NANDN U10148 ( .A(n8998), .B(n8997), .Z(n9002) );
  OR U10149 ( .A(n9000), .B(n8999), .Z(n9001) );
  NAND U10150 ( .A(n9002), .B(n9001), .Z(n9146) );
  NAND U10151 ( .A(n9004), .B(n9003), .Z(n9008) );
  NANDN U10152 ( .A(n9006), .B(n9005), .Z(n9007) );
  NAND U10153 ( .A(n9008), .B(n9007), .Z(n9147) );
  XNOR U10154 ( .A(n9146), .B(n9147), .Z(n9148) );
  XOR U10155 ( .A(n9149), .B(n9148), .Z(n9023) );
  XOR U10156 ( .A(n9022), .B(n9023), .Z(n9014) );
  XOR U10157 ( .A(n9015), .B(n9014), .Z(n9016) );
  XNOR U10158 ( .A(n9017), .B(n9016), .Z(n9158) );
  XNOR U10159 ( .A(n9158), .B(sreg[294]), .Z(n9160) );
  NAND U10160 ( .A(n9009), .B(sreg[293]), .Z(n9013) );
  OR U10161 ( .A(n9011), .B(n9010), .Z(n9012) );
  AND U10162 ( .A(n9013), .B(n9012), .Z(n9159) );
  XOR U10163 ( .A(n9160), .B(n9159), .Z(c[294]) );
  NAND U10164 ( .A(n9015), .B(n9014), .Z(n9019) );
  NAND U10165 ( .A(n9017), .B(n9016), .Z(n9018) );
  NAND U10166 ( .A(n9019), .B(n9018), .Z(n9166) );
  NANDN U10167 ( .A(n9021), .B(n9020), .Z(n9025) );
  NAND U10168 ( .A(n9023), .B(n9022), .Z(n9024) );
  NAND U10169 ( .A(n9025), .B(n9024), .Z(n9164) );
  NANDN U10170 ( .A(n9027), .B(n9026), .Z(n9031) );
  NAND U10171 ( .A(n9029), .B(n9028), .Z(n9030) );
  NAND U10172 ( .A(n9031), .B(n9030), .Z(n9250) );
  XNOR U10173 ( .A(b[19]), .B(a[53]), .Z(n9193) );
  NANDN U10174 ( .A(n9193), .B(n37934), .Z(n9034) );
  NANDN U10175 ( .A(n9032), .B(n37935), .Z(n9033) );
  NAND U10176 ( .A(n9034), .B(n9033), .Z(n9260) );
  XOR U10177 ( .A(b[27]), .B(a[45]), .Z(n9196) );
  NAND U10178 ( .A(n38423), .B(n9196), .Z(n9037) );
  NANDN U10179 ( .A(n9035), .B(n38424), .Z(n9036) );
  NAND U10180 ( .A(n9037), .B(n9036), .Z(n9257) );
  XOR U10181 ( .A(b[5]), .B(n13219), .Z(n9199) );
  NANDN U10182 ( .A(n9199), .B(n36587), .Z(n9040) );
  NANDN U10183 ( .A(n9038), .B(n36588), .Z(n9039) );
  AND U10184 ( .A(n9040), .B(n9039), .Z(n9258) );
  XNOR U10185 ( .A(n9257), .B(n9258), .Z(n9259) );
  XNOR U10186 ( .A(n9260), .B(n9259), .Z(n9248) );
  NANDN U10187 ( .A(n9041), .B(n37762), .Z(n9043) );
  XOR U10188 ( .A(b[17]), .B(a[55]), .Z(n9202) );
  NAND U10189 ( .A(n9202), .B(n37764), .Z(n9042) );
  NAND U10190 ( .A(n9043), .B(n9042), .Z(n9220) );
  XNOR U10191 ( .A(b[31]), .B(a[41]), .Z(n9205) );
  NANDN U10192 ( .A(n9205), .B(n38552), .Z(n9046) );
  NANDN U10193 ( .A(n9044), .B(n38553), .Z(n9045) );
  NAND U10194 ( .A(n9046), .B(n9045), .Z(n9217) );
  OR U10195 ( .A(n9047), .B(n36105), .Z(n9049) );
  XNOR U10196 ( .A(b[3]), .B(a[69]), .Z(n9208) );
  NANDN U10197 ( .A(n9208), .B(n36107), .Z(n9048) );
  AND U10198 ( .A(n9049), .B(n9048), .Z(n9218) );
  XNOR U10199 ( .A(n9217), .B(n9218), .Z(n9219) );
  XOR U10200 ( .A(n9220), .B(n9219), .Z(n9247) );
  XNOR U10201 ( .A(n9248), .B(n9247), .Z(n9249) );
  XNOR U10202 ( .A(n9250), .B(n9249), .Z(n9293) );
  NANDN U10203 ( .A(n9051), .B(n9050), .Z(n9055) );
  NAND U10204 ( .A(n9053), .B(n9052), .Z(n9054) );
  NAND U10205 ( .A(n9055), .B(n9054), .Z(n9238) );
  NANDN U10206 ( .A(n9057), .B(n9056), .Z(n9061) );
  NAND U10207 ( .A(n9059), .B(n9058), .Z(n9060) );
  NAND U10208 ( .A(n9061), .B(n9060), .Z(n9236) );
  OR U10209 ( .A(n9063), .B(n9062), .Z(n9067) );
  NANDN U10210 ( .A(n9065), .B(n9064), .Z(n9066) );
  NAND U10211 ( .A(n9067), .B(n9066), .Z(n9235) );
  XNOR U10212 ( .A(n9238), .B(n9237), .Z(n9294) );
  XOR U10213 ( .A(n9293), .B(n9294), .Z(n9296) );
  NANDN U10214 ( .A(n9069), .B(n9068), .Z(n9073) );
  NANDN U10215 ( .A(n9071), .B(n9070), .Z(n9072) );
  NAND U10216 ( .A(n9073), .B(n9072), .Z(n9295) );
  XOR U10217 ( .A(n9296), .B(n9295), .Z(n9183) );
  OR U10218 ( .A(n9075), .B(n9074), .Z(n9079) );
  NANDN U10219 ( .A(n9077), .B(n9076), .Z(n9078) );
  NAND U10220 ( .A(n9079), .B(n9078), .Z(n9182) );
  NANDN U10221 ( .A(n9081), .B(n9080), .Z(n9085) );
  NANDN U10222 ( .A(n9083), .B(n9082), .Z(n9084) );
  NAND U10223 ( .A(n9085), .B(n9084), .Z(n9301) );
  NANDN U10224 ( .A(n9087), .B(n9086), .Z(n9091) );
  OR U10225 ( .A(n9089), .B(n9088), .Z(n9090) );
  NAND U10226 ( .A(n9091), .B(n9090), .Z(n9300) );
  NANDN U10227 ( .A(n9093), .B(n9092), .Z(n9097) );
  NAND U10228 ( .A(n9095), .B(n9094), .Z(n9096) );
  NAND U10229 ( .A(n9097), .B(n9096), .Z(n9241) );
  NANDN U10230 ( .A(n9099), .B(n9098), .Z(n9103) );
  NAND U10231 ( .A(n9101), .B(n9100), .Z(n9102) );
  AND U10232 ( .A(n9103), .B(n9102), .Z(n9242) );
  XNOR U10233 ( .A(n9241), .B(n9242), .Z(n9243) );
  XNOR U10234 ( .A(b[9]), .B(a[63]), .Z(n9263) );
  NANDN U10235 ( .A(n9263), .B(n36925), .Z(n9106) );
  NANDN U10236 ( .A(n9104), .B(n36926), .Z(n9105) );
  NAND U10237 ( .A(n9106), .B(n9105), .Z(n9225) );
  XNOR U10238 ( .A(b[15]), .B(a[57]), .Z(n9266) );
  OR U10239 ( .A(n9266), .B(n37665), .Z(n9109) );
  NANDN U10240 ( .A(n9107), .B(n37604), .Z(n9108) );
  AND U10241 ( .A(n9109), .B(n9108), .Z(n9223) );
  XNOR U10242 ( .A(b[21]), .B(a[51]), .Z(n9269) );
  NANDN U10243 ( .A(n9269), .B(n38101), .Z(n9112) );
  NANDN U10244 ( .A(n9110), .B(n38102), .Z(n9111) );
  AND U10245 ( .A(n9112), .B(n9111), .Z(n9224) );
  XOR U10246 ( .A(n9225), .B(n9226), .Z(n9214) );
  XNOR U10247 ( .A(b[11]), .B(a[61]), .Z(n9272) );
  OR U10248 ( .A(n9272), .B(n37311), .Z(n9115) );
  NANDN U10249 ( .A(n9113), .B(n37218), .Z(n9114) );
  NAND U10250 ( .A(n9115), .B(n9114), .Z(n9212) );
  XOR U10251 ( .A(n1053), .B(a[59]), .Z(n9275) );
  NANDN U10252 ( .A(n9275), .B(n37424), .Z(n9118) );
  NANDN U10253 ( .A(n9116), .B(n37425), .Z(n9117) );
  AND U10254 ( .A(n9118), .B(n9117), .Z(n9211) );
  XNOR U10255 ( .A(n9212), .B(n9211), .Z(n9213) );
  XOR U10256 ( .A(n9214), .B(n9213), .Z(n9231) );
  NANDN U10257 ( .A(n1049), .B(a[71]), .Z(n9119) );
  XNOR U10258 ( .A(b[1]), .B(n9119), .Z(n9121) );
  NANDN U10259 ( .A(b[0]), .B(a[70]), .Z(n9120) );
  AND U10260 ( .A(n9121), .B(n9120), .Z(n9189) );
  NAND U10261 ( .A(n38490), .B(n9122), .Z(n9124) );
  XNOR U10262 ( .A(n1058), .B(a[43]), .Z(n9281) );
  NANDN U10263 ( .A(n1048), .B(n9281), .Z(n9123) );
  NAND U10264 ( .A(n9124), .B(n9123), .Z(n9187) );
  NANDN U10265 ( .A(n1059), .B(a[39]), .Z(n9188) );
  XNOR U10266 ( .A(n9187), .B(n9188), .Z(n9190) );
  XOR U10267 ( .A(n9189), .B(n9190), .Z(n9229) );
  NANDN U10268 ( .A(n9125), .B(n38205), .Z(n9127) );
  XNOR U10269 ( .A(b[23]), .B(a[49]), .Z(n9284) );
  OR U10270 ( .A(n9284), .B(n38268), .Z(n9126) );
  NAND U10271 ( .A(n9127), .B(n9126), .Z(n9254) );
  XOR U10272 ( .A(b[7]), .B(a[65]), .Z(n9287) );
  NAND U10273 ( .A(n9287), .B(n36701), .Z(n9130) );
  NAND U10274 ( .A(n9128), .B(n36702), .Z(n9129) );
  NAND U10275 ( .A(n9130), .B(n9129), .Z(n9251) );
  XOR U10276 ( .A(b[25]), .B(a[47]), .Z(n9290) );
  NAND U10277 ( .A(n9290), .B(n38325), .Z(n9133) );
  NAND U10278 ( .A(n9131), .B(n38326), .Z(n9132) );
  AND U10279 ( .A(n9133), .B(n9132), .Z(n9252) );
  XNOR U10280 ( .A(n9251), .B(n9252), .Z(n9253) );
  XNOR U10281 ( .A(n9254), .B(n9253), .Z(n9230) );
  XOR U10282 ( .A(n9229), .B(n9230), .Z(n9232) );
  XNOR U10283 ( .A(n9231), .B(n9232), .Z(n9244) );
  XNOR U10284 ( .A(n9243), .B(n9244), .Z(n9299) );
  XNOR U10285 ( .A(n9300), .B(n9299), .Z(n9302) );
  XOR U10286 ( .A(n9301), .B(n9302), .Z(n9181) );
  XOR U10287 ( .A(n9182), .B(n9181), .Z(n9184) );
  NAND U10288 ( .A(n9135), .B(n9134), .Z(n9139) );
  NAND U10289 ( .A(n9137), .B(n9136), .Z(n9138) );
  NAND U10290 ( .A(n9139), .B(n9138), .Z(n9176) );
  NANDN U10291 ( .A(n9141), .B(n9140), .Z(n9145) );
  NAND U10292 ( .A(n9143), .B(n9142), .Z(n9144) );
  AND U10293 ( .A(n9145), .B(n9144), .Z(n9175) );
  XNOR U10294 ( .A(n9176), .B(n9175), .Z(n9177) );
  XOR U10295 ( .A(n9178), .B(n9177), .Z(n9171) );
  NANDN U10296 ( .A(n9147), .B(n9146), .Z(n9151) );
  NAND U10297 ( .A(n9149), .B(n9148), .Z(n9150) );
  NAND U10298 ( .A(n9151), .B(n9150), .Z(n9169) );
  NANDN U10299 ( .A(n9153), .B(n9152), .Z(n9157) );
  NANDN U10300 ( .A(n9155), .B(n9154), .Z(n9156) );
  NAND U10301 ( .A(n9157), .B(n9156), .Z(n9170) );
  XNOR U10302 ( .A(n9169), .B(n9170), .Z(n9172) );
  XOR U10303 ( .A(n9171), .B(n9172), .Z(n9163) );
  XOR U10304 ( .A(n9164), .B(n9163), .Z(n9165) );
  XNOR U10305 ( .A(n9166), .B(n9165), .Z(n9303) );
  XNOR U10306 ( .A(n9303), .B(sreg[295]), .Z(n9305) );
  NAND U10307 ( .A(n9158), .B(sreg[294]), .Z(n9162) );
  OR U10308 ( .A(n9160), .B(n9159), .Z(n9161) );
  AND U10309 ( .A(n9162), .B(n9161), .Z(n9304) );
  XOR U10310 ( .A(n9305), .B(n9304), .Z(c[295]) );
  NAND U10311 ( .A(n9164), .B(n9163), .Z(n9168) );
  NAND U10312 ( .A(n9166), .B(n9165), .Z(n9167) );
  NAND U10313 ( .A(n9168), .B(n9167), .Z(n9311) );
  NANDN U10314 ( .A(n9170), .B(n9169), .Z(n9174) );
  NAND U10315 ( .A(n9172), .B(n9171), .Z(n9173) );
  NAND U10316 ( .A(n9174), .B(n9173), .Z(n9309) );
  NANDN U10317 ( .A(n9176), .B(n9175), .Z(n9180) );
  NAND U10318 ( .A(n9178), .B(n9177), .Z(n9179) );
  NAND U10319 ( .A(n9180), .B(n9179), .Z(n9314) );
  NANDN U10320 ( .A(n9182), .B(n9181), .Z(n9186) );
  OR U10321 ( .A(n9184), .B(n9183), .Z(n9185) );
  NAND U10322 ( .A(n9186), .B(n9185), .Z(n9315) );
  XNOR U10323 ( .A(n9314), .B(n9315), .Z(n9316) );
  NANDN U10324 ( .A(n9188), .B(n9187), .Z(n9192) );
  NAND U10325 ( .A(n9190), .B(n9189), .Z(n9191) );
  NAND U10326 ( .A(n9192), .B(n9191), .Z(n9395) );
  XOR U10327 ( .A(b[19]), .B(n11319), .Z(n9362) );
  NANDN U10328 ( .A(n9362), .B(n37934), .Z(n9195) );
  NANDN U10329 ( .A(n9193), .B(n37935), .Z(n9194) );
  NAND U10330 ( .A(n9195), .B(n9194), .Z(n9407) );
  XOR U10331 ( .A(b[27]), .B(a[46]), .Z(n9365) );
  NAND U10332 ( .A(n38423), .B(n9365), .Z(n9198) );
  NAND U10333 ( .A(n9196), .B(n38424), .Z(n9197) );
  NAND U10334 ( .A(n9198), .B(n9197), .Z(n9404) );
  XNOR U10335 ( .A(b[5]), .B(a[68]), .Z(n9368) );
  NANDN U10336 ( .A(n9368), .B(n36587), .Z(n9201) );
  NANDN U10337 ( .A(n9199), .B(n36588), .Z(n9200) );
  AND U10338 ( .A(n9201), .B(n9200), .Z(n9405) );
  XNOR U10339 ( .A(n9404), .B(n9405), .Z(n9406) );
  XNOR U10340 ( .A(n9407), .B(n9406), .Z(n9392) );
  NAND U10341 ( .A(n9202), .B(n37762), .Z(n9204) );
  XOR U10342 ( .A(b[17]), .B(a[56]), .Z(n9371) );
  NAND U10343 ( .A(n9371), .B(n37764), .Z(n9203) );
  NAND U10344 ( .A(n9204), .B(n9203), .Z(n9346) );
  XNOR U10345 ( .A(b[31]), .B(a[42]), .Z(n9374) );
  NANDN U10346 ( .A(n9374), .B(n38552), .Z(n9207) );
  NANDN U10347 ( .A(n9205), .B(n38553), .Z(n9206) );
  AND U10348 ( .A(n9207), .B(n9206), .Z(n9344) );
  OR U10349 ( .A(n9208), .B(n36105), .Z(n9210) );
  XNOR U10350 ( .A(b[3]), .B(a[70]), .Z(n9377) );
  NANDN U10351 ( .A(n9377), .B(n36107), .Z(n9209) );
  AND U10352 ( .A(n9210), .B(n9209), .Z(n9345) );
  XOR U10353 ( .A(n9346), .B(n9347), .Z(n9393) );
  XOR U10354 ( .A(n9392), .B(n9393), .Z(n9394) );
  XNOR U10355 ( .A(n9395), .B(n9394), .Z(n9440) );
  NANDN U10356 ( .A(n9212), .B(n9211), .Z(n9216) );
  NAND U10357 ( .A(n9214), .B(n9213), .Z(n9215) );
  NAND U10358 ( .A(n9216), .B(n9215), .Z(n9383) );
  NANDN U10359 ( .A(n9218), .B(n9217), .Z(n9222) );
  NAND U10360 ( .A(n9220), .B(n9219), .Z(n9221) );
  NAND U10361 ( .A(n9222), .B(n9221), .Z(n9381) );
  OR U10362 ( .A(n9224), .B(n9223), .Z(n9228) );
  NANDN U10363 ( .A(n9226), .B(n9225), .Z(n9227) );
  NAND U10364 ( .A(n9228), .B(n9227), .Z(n9380) );
  XNOR U10365 ( .A(n9383), .B(n9382), .Z(n9441) );
  XOR U10366 ( .A(n9440), .B(n9441), .Z(n9443) );
  NANDN U10367 ( .A(n9230), .B(n9229), .Z(n9234) );
  OR U10368 ( .A(n9232), .B(n9231), .Z(n9233) );
  NAND U10369 ( .A(n9234), .B(n9233), .Z(n9442) );
  XOR U10370 ( .A(n9443), .B(n9442), .Z(n9328) );
  OR U10371 ( .A(n9236), .B(n9235), .Z(n9240) );
  NAND U10372 ( .A(n9238), .B(n9237), .Z(n9239) );
  NAND U10373 ( .A(n9240), .B(n9239), .Z(n9327) );
  NANDN U10374 ( .A(n9242), .B(n9241), .Z(n9246) );
  NANDN U10375 ( .A(n9244), .B(n9243), .Z(n9245) );
  NAND U10376 ( .A(n9246), .B(n9245), .Z(n9448) );
  NANDN U10377 ( .A(n9252), .B(n9251), .Z(n9256) );
  NAND U10378 ( .A(n9254), .B(n9253), .Z(n9255) );
  NAND U10379 ( .A(n9256), .B(n9255), .Z(n9386) );
  NANDN U10380 ( .A(n9258), .B(n9257), .Z(n9262) );
  NAND U10381 ( .A(n9260), .B(n9259), .Z(n9261) );
  AND U10382 ( .A(n9262), .B(n9261), .Z(n9387) );
  XNOR U10383 ( .A(n9386), .B(n9387), .Z(n9388) );
  XNOR U10384 ( .A(b[9]), .B(a[64]), .Z(n9410) );
  NANDN U10385 ( .A(n9410), .B(n36925), .Z(n9265) );
  NANDN U10386 ( .A(n9263), .B(n36926), .Z(n9264) );
  NAND U10387 ( .A(n9265), .B(n9264), .Z(n9352) );
  XNOR U10388 ( .A(b[15]), .B(a[58]), .Z(n9413) );
  OR U10389 ( .A(n9413), .B(n37665), .Z(n9268) );
  NANDN U10390 ( .A(n9266), .B(n37604), .Z(n9267) );
  AND U10391 ( .A(n9268), .B(n9267), .Z(n9350) );
  XNOR U10392 ( .A(b[21]), .B(a[52]), .Z(n9416) );
  NANDN U10393 ( .A(n9416), .B(n38101), .Z(n9271) );
  NANDN U10394 ( .A(n9269), .B(n38102), .Z(n9270) );
  AND U10395 ( .A(n9271), .B(n9270), .Z(n9351) );
  XOR U10396 ( .A(n9352), .B(n9353), .Z(n9341) );
  XOR U10397 ( .A(b[11]), .B(n12493), .Z(n9419) );
  OR U10398 ( .A(n9419), .B(n37311), .Z(n9274) );
  NANDN U10399 ( .A(n9272), .B(n37218), .Z(n9273) );
  NAND U10400 ( .A(n9274), .B(n9273), .Z(n9339) );
  XOR U10401 ( .A(n1053), .B(a[60]), .Z(n9422) );
  NANDN U10402 ( .A(n9422), .B(n37424), .Z(n9277) );
  NANDN U10403 ( .A(n9275), .B(n37425), .Z(n9276) );
  NAND U10404 ( .A(n9277), .B(n9276), .Z(n9338) );
  XOR U10405 ( .A(n9341), .B(n9340), .Z(n9335) );
  NANDN U10406 ( .A(n1049), .B(a[72]), .Z(n9278) );
  XNOR U10407 ( .A(b[1]), .B(n9278), .Z(n9280) );
  NANDN U10408 ( .A(b[0]), .B(a[71]), .Z(n9279) );
  AND U10409 ( .A(n9280), .B(n9279), .Z(n9358) );
  NAND U10410 ( .A(n38490), .B(n9281), .Z(n9283) );
  XOR U10411 ( .A(n1058), .B(n9873), .Z(n9428) );
  NANDN U10412 ( .A(n1048), .B(n9428), .Z(n9282) );
  NAND U10413 ( .A(n9283), .B(n9282), .Z(n9356) );
  NANDN U10414 ( .A(n1059), .B(a[40]), .Z(n9357) );
  XNOR U10415 ( .A(n9356), .B(n9357), .Z(n9359) );
  XNOR U10416 ( .A(n9358), .B(n9359), .Z(n9333) );
  NANDN U10417 ( .A(n9284), .B(n38205), .Z(n9286) );
  XOR U10418 ( .A(b[23]), .B(n10724), .Z(n9431) );
  OR U10419 ( .A(n9431), .B(n38268), .Z(n9285) );
  NAND U10420 ( .A(n9286), .B(n9285), .Z(n9401) );
  XOR U10421 ( .A(b[7]), .B(a[66]), .Z(n9434) );
  NAND U10422 ( .A(n9434), .B(n36701), .Z(n9289) );
  NAND U10423 ( .A(n9287), .B(n36702), .Z(n9288) );
  NAND U10424 ( .A(n9289), .B(n9288), .Z(n9398) );
  XOR U10425 ( .A(b[25]), .B(a[48]), .Z(n9437) );
  NAND U10426 ( .A(n9437), .B(n38325), .Z(n9292) );
  NAND U10427 ( .A(n9290), .B(n38326), .Z(n9291) );
  AND U10428 ( .A(n9292), .B(n9291), .Z(n9399) );
  XNOR U10429 ( .A(n9398), .B(n9399), .Z(n9400) );
  XOR U10430 ( .A(n9401), .B(n9400), .Z(n9332) );
  XOR U10431 ( .A(n9335), .B(n9334), .Z(n9389) );
  XNOR U10432 ( .A(n9388), .B(n9389), .Z(n9446) );
  XNOR U10433 ( .A(n9447), .B(n9446), .Z(n9449) );
  XNOR U10434 ( .A(n9448), .B(n9449), .Z(n9326) );
  XOR U10435 ( .A(n9327), .B(n9326), .Z(n9329) );
  NANDN U10436 ( .A(n9294), .B(n9293), .Z(n9298) );
  OR U10437 ( .A(n9296), .B(n9295), .Z(n9297) );
  NAND U10438 ( .A(n9298), .B(n9297), .Z(n9320) );
  XNOR U10439 ( .A(n9320), .B(n9321), .Z(n9322) );
  XOR U10440 ( .A(n9323), .B(n9322), .Z(n9317) );
  XOR U10441 ( .A(n9316), .B(n9317), .Z(n9308) );
  XOR U10442 ( .A(n9309), .B(n9308), .Z(n9310) );
  XNOR U10443 ( .A(n9311), .B(n9310), .Z(n9452) );
  XNOR U10444 ( .A(n9452), .B(sreg[296]), .Z(n9454) );
  NAND U10445 ( .A(n9303), .B(sreg[295]), .Z(n9307) );
  OR U10446 ( .A(n9305), .B(n9304), .Z(n9306) );
  AND U10447 ( .A(n9307), .B(n9306), .Z(n9453) );
  XOR U10448 ( .A(n9454), .B(n9453), .Z(c[296]) );
  NAND U10449 ( .A(n9309), .B(n9308), .Z(n9313) );
  NAND U10450 ( .A(n9311), .B(n9310), .Z(n9312) );
  NAND U10451 ( .A(n9313), .B(n9312), .Z(n9460) );
  NANDN U10452 ( .A(n9315), .B(n9314), .Z(n9319) );
  NAND U10453 ( .A(n9317), .B(n9316), .Z(n9318) );
  NAND U10454 ( .A(n9319), .B(n9318), .Z(n9458) );
  NANDN U10455 ( .A(n9321), .B(n9320), .Z(n9325) );
  NAND U10456 ( .A(n9323), .B(n9322), .Z(n9324) );
  NAND U10457 ( .A(n9325), .B(n9324), .Z(n9463) );
  NANDN U10458 ( .A(n9327), .B(n9326), .Z(n9331) );
  OR U10459 ( .A(n9329), .B(n9328), .Z(n9330) );
  NAND U10460 ( .A(n9331), .B(n9330), .Z(n9464) );
  XNOR U10461 ( .A(n9463), .B(n9464), .Z(n9465) );
  NANDN U10462 ( .A(n9333), .B(n9332), .Z(n9337) );
  NANDN U10463 ( .A(n9335), .B(n9334), .Z(n9336) );
  NAND U10464 ( .A(n9337), .B(n9336), .Z(n9580) );
  OR U10465 ( .A(n9339), .B(n9338), .Z(n9343) );
  NAND U10466 ( .A(n9341), .B(n9340), .Z(n9342) );
  NAND U10467 ( .A(n9343), .B(n9342), .Z(n9519) );
  OR U10468 ( .A(n9345), .B(n9344), .Z(n9349) );
  NANDN U10469 ( .A(n9347), .B(n9346), .Z(n9348) );
  NAND U10470 ( .A(n9349), .B(n9348), .Z(n9518) );
  OR U10471 ( .A(n9351), .B(n9350), .Z(n9355) );
  NANDN U10472 ( .A(n9353), .B(n9352), .Z(n9354) );
  NAND U10473 ( .A(n9355), .B(n9354), .Z(n9517) );
  XOR U10474 ( .A(n9519), .B(n9520), .Z(n9577) );
  NANDN U10475 ( .A(n9357), .B(n9356), .Z(n9361) );
  NAND U10476 ( .A(n9359), .B(n9358), .Z(n9360) );
  NAND U10477 ( .A(n9361), .B(n9360), .Z(n9532) );
  XNOR U10478 ( .A(b[19]), .B(a[55]), .Z(n9475) );
  NANDN U10479 ( .A(n9475), .B(n37934), .Z(n9364) );
  NANDN U10480 ( .A(n9362), .B(n37935), .Z(n9363) );
  NAND U10481 ( .A(n9364), .B(n9363), .Z(n9568) );
  XOR U10482 ( .A(b[27]), .B(a[47]), .Z(n9478) );
  NAND U10483 ( .A(n38423), .B(n9478), .Z(n9367) );
  NAND U10484 ( .A(n9365), .B(n38424), .Z(n9366) );
  NAND U10485 ( .A(n9367), .B(n9366), .Z(n9565) );
  XNOR U10486 ( .A(b[5]), .B(a[69]), .Z(n9481) );
  NANDN U10487 ( .A(n9481), .B(n36587), .Z(n9370) );
  NANDN U10488 ( .A(n9368), .B(n36588), .Z(n9369) );
  AND U10489 ( .A(n9370), .B(n9369), .Z(n9566) );
  XNOR U10490 ( .A(n9565), .B(n9566), .Z(n9567) );
  XNOR U10491 ( .A(n9568), .B(n9567), .Z(n9530) );
  NAND U10492 ( .A(n9371), .B(n37762), .Z(n9373) );
  XOR U10493 ( .A(b[17]), .B(a[57]), .Z(n9484) );
  NAND U10494 ( .A(n9484), .B(n37764), .Z(n9372) );
  NAND U10495 ( .A(n9373), .B(n9372), .Z(n9502) );
  XNOR U10496 ( .A(b[31]), .B(a[43]), .Z(n9487) );
  NANDN U10497 ( .A(n9487), .B(n38552), .Z(n9376) );
  NANDN U10498 ( .A(n9374), .B(n38553), .Z(n9375) );
  NAND U10499 ( .A(n9376), .B(n9375), .Z(n9499) );
  OR U10500 ( .A(n9377), .B(n36105), .Z(n9379) );
  XNOR U10501 ( .A(b[3]), .B(a[71]), .Z(n9490) );
  NANDN U10502 ( .A(n9490), .B(n36107), .Z(n9378) );
  AND U10503 ( .A(n9379), .B(n9378), .Z(n9500) );
  XNOR U10504 ( .A(n9499), .B(n9500), .Z(n9501) );
  XOR U10505 ( .A(n9502), .B(n9501), .Z(n9529) );
  XNOR U10506 ( .A(n9530), .B(n9529), .Z(n9531) );
  XNOR U10507 ( .A(n9532), .B(n9531), .Z(n9578) );
  XNOR U10508 ( .A(n9577), .B(n9578), .Z(n9579) );
  XNOR U10509 ( .A(n9580), .B(n9579), .Z(n9598) );
  OR U10510 ( .A(n9381), .B(n9380), .Z(n9385) );
  NAND U10511 ( .A(n9383), .B(n9382), .Z(n9384) );
  NAND U10512 ( .A(n9385), .B(n9384), .Z(n9596) );
  NANDN U10513 ( .A(n9387), .B(n9386), .Z(n9391) );
  NANDN U10514 ( .A(n9389), .B(n9388), .Z(n9390) );
  NAND U10515 ( .A(n9391), .B(n9390), .Z(n9585) );
  OR U10516 ( .A(n9393), .B(n9392), .Z(n9397) );
  NAND U10517 ( .A(n9395), .B(n9394), .Z(n9396) );
  NAND U10518 ( .A(n9397), .B(n9396), .Z(n9584) );
  NANDN U10519 ( .A(n9399), .B(n9398), .Z(n9403) );
  NAND U10520 ( .A(n9401), .B(n9400), .Z(n9402) );
  NAND U10521 ( .A(n9403), .B(n9402), .Z(n9523) );
  NANDN U10522 ( .A(n9405), .B(n9404), .Z(n9409) );
  NAND U10523 ( .A(n9407), .B(n9406), .Z(n9408) );
  AND U10524 ( .A(n9409), .B(n9408), .Z(n9524) );
  XNOR U10525 ( .A(n9523), .B(n9524), .Z(n9525) );
  XNOR U10526 ( .A(b[9]), .B(a[65]), .Z(n9535) );
  NANDN U10527 ( .A(n9535), .B(n36925), .Z(n9412) );
  NANDN U10528 ( .A(n9410), .B(n36926), .Z(n9411) );
  NAND U10529 ( .A(n9412), .B(n9411), .Z(n9513) );
  XOR U10530 ( .A(b[15]), .B(n12056), .Z(n9538) );
  OR U10531 ( .A(n9538), .B(n37665), .Z(n9415) );
  NANDN U10532 ( .A(n9413), .B(n37604), .Z(n9414) );
  AND U10533 ( .A(n9415), .B(n9414), .Z(n9511) );
  XNOR U10534 ( .A(b[21]), .B(a[53]), .Z(n9541) );
  NANDN U10535 ( .A(n9541), .B(n38101), .Z(n9418) );
  NANDN U10536 ( .A(n9416), .B(n38102), .Z(n9417) );
  AND U10537 ( .A(n9418), .B(n9417), .Z(n9512) );
  XOR U10538 ( .A(n9513), .B(n9514), .Z(n9508) );
  XNOR U10539 ( .A(b[11]), .B(a[63]), .Z(n9544) );
  OR U10540 ( .A(n9544), .B(n37311), .Z(n9421) );
  NANDN U10541 ( .A(n9419), .B(n37218), .Z(n9420) );
  NAND U10542 ( .A(n9421), .B(n9420), .Z(n9506) );
  XOR U10543 ( .A(n1053), .B(a[61]), .Z(n9547) );
  NANDN U10544 ( .A(n9547), .B(n37424), .Z(n9424) );
  NANDN U10545 ( .A(n9422), .B(n37425), .Z(n9423) );
  AND U10546 ( .A(n9424), .B(n9423), .Z(n9505) );
  XNOR U10547 ( .A(n9506), .B(n9505), .Z(n9507) );
  XOR U10548 ( .A(n9508), .B(n9507), .Z(n9495) );
  NANDN U10549 ( .A(n1049), .B(a[73]), .Z(n9425) );
  XNOR U10550 ( .A(b[1]), .B(n9425), .Z(n9427) );
  NANDN U10551 ( .A(b[0]), .B(a[72]), .Z(n9426) );
  AND U10552 ( .A(n9427), .B(n9426), .Z(n9471) );
  NAND U10553 ( .A(n38490), .B(n9428), .Z(n9430) );
  XNOR U10554 ( .A(n1058), .B(a[45]), .Z(n9553) );
  NANDN U10555 ( .A(n1048), .B(n9553), .Z(n9429) );
  NAND U10556 ( .A(n9430), .B(n9429), .Z(n9469) );
  NANDN U10557 ( .A(n1059), .B(a[41]), .Z(n9470) );
  XNOR U10558 ( .A(n9469), .B(n9470), .Z(n9472) );
  XOR U10559 ( .A(n9471), .B(n9472), .Z(n9493) );
  NANDN U10560 ( .A(n9431), .B(n38205), .Z(n9433) );
  XNOR U10561 ( .A(b[23]), .B(a[51]), .Z(n9556) );
  OR U10562 ( .A(n9556), .B(n38268), .Z(n9432) );
  NAND U10563 ( .A(n9433), .B(n9432), .Z(n9574) );
  XNOR U10564 ( .A(b[7]), .B(a[67]), .Z(n9559) );
  NANDN U10565 ( .A(n9559), .B(n36701), .Z(n9436) );
  NAND U10566 ( .A(n9434), .B(n36702), .Z(n9435) );
  NAND U10567 ( .A(n9436), .B(n9435), .Z(n9571) );
  XOR U10568 ( .A(b[25]), .B(a[49]), .Z(n9562) );
  NAND U10569 ( .A(n9562), .B(n38325), .Z(n9439) );
  NAND U10570 ( .A(n9437), .B(n38326), .Z(n9438) );
  AND U10571 ( .A(n9439), .B(n9438), .Z(n9572) );
  XNOR U10572 ( .A(n9571), .B(n9572), .Z(n9573) );
  XNOR U10573 ( .A(n9574), .B(n9573), .Z(n9494) );
  XOR U10574 ( .A(n9493), .B(n9494), .Z(n9496) );
  XNOR U10575 ( .A(n9495), .B(n9496), .Z(n9526) );
  XNOR U10576 ( .A(n9525), .B(n9526), .Z(n9583) );
  XNOR U10577 ( .A(n9584), .B(n9583), .Z(n9586) );
  XNOR U10578 ( .A(n9585), .B(n9586), .Z(n9595) );
  XNOR U10579 ( .A(n9596), .B(n9595), .Z(n9597) );
  XOR U10580 ( .A(n9598), .B(n9597), .Z(n9592) );
  NANDN U10581 ( .A(n9441), .B(n9440), .Z(n9445) );
  OR U10582 ( .A(n9443), .B(n9442), .Z(n9444) );
  NAND U10583 ( .A(n9445), .B(n9444), .Z(n9589) );
  NAND U10584 ( .A(n9447), .B(n9446), .Z(n9451) );
  NANDN U10585 ( .A(n9449), .B(n9448), .Z(n9450) );
  NAND U10586 ( .A(n9451), .B(n9450), .Z(n9590) );
  XNOR U10587 ( .A(n9589), .B(n9590), .Z(n9591) );
  XOR U10588 ( .A(n9592), .B(n9591), .Z(n9466) );
  XOR U10589 ( .A(n9465), .B(n9466), .Z(n9457) );
  XOR U10590 ( .A(n9458), .B(n9457), .Z(n9459) );
  XNOR U10591 ( .A(n9460), .B(n9459), .Z(n9601) );
  XNOR U10592 ( .A(n9601), .B(sreg[297]), .Z(n9603) );
  NAND U10593 ( .A(n9452), .B(sreg[296]), .Z(n9456) );
  OR U10594 ( .A(n9454), .B(n9453), .Z(n9455) );
  AND U10595 ( .A(n9456), .B(n9455), .Z(n9602) );
  XOR U10596 ( .A(n9603), .B(n9602), .Z(c[297]) );
  NAND U10597 ( .A(n9458), .B(n9457), .Z(n9462) );
  NAND U10598 ( .A(n9460), .B(n9459), .Z(n9461) );
  NAND U10599 ( .A(n9462), .B(n9461), .Z(n9609) );
  NANDN U10600 ( .A(n9464), .B(n9463), .Z(n9468) );
  NAND U10601 ( .A(n9466), .B(n9465), .Z(n9467) );
  NAND U10602 ( .A(n9468), .B(n9467), .Z(n9607) );
  NANDN U10603 ( .A(n9470), .B(n9469), .Z(n9474) );
  NAND U10604 ( .A(n9472), .B(n9471), .Z(n9473) );
  NAND U10605 ( .A(n9474), .B(n9473), .Z(n9691) );
  XNOR U10606 ( .A(b[19]), .B(a[56]), .Z(n9658) );
  NANDN U10607 ( .A(n9658), .B(n37934), .Z(n9477) );
  NANDN U10608 ( .A(n9475), .B(n37935), .Z(n9476) );
  NAND U10609 ( .A(n9477), .B(n9476), .Z(n9703) );
  XOR U10610 ( .A(b[27]), .B(a[48]), .Z(n9661) );
  NAND U10611 ( .A(n38423), .B(n9661), .Z(n9480) );
  NAND U10612 ( .A(n9478), .B(n38424), .Z(n9479) );
  NAND U10613 ( .A(n9480), .B(n9479), .Z(n9700) );
  XNOR U10614 ( .A(b[5]), .B(a[70]), .Z(n9664) );
  NANDN U10615 ( .A(n9664), .B(n36587), .Z(n9483) );
  NANDN U10616 ( .A(n9481), .B(n36588), .Z(n9482) );
  AND U10617 ( .A(n9483), .B(n9482), .Z(n9701) );
  XNOR U10618 ( .A(n9700), .B(n9701), .Z(n9702) );
  XNOR U10619 ( .A(n9703), .B(n9702), .Z(n9688) );
  NAND U10620 ( .A(n9484), .B(n37762), .Z(n9486) );
  XOR U10621 ( .A(b[17]), .B(a[58]), .Z(n9667) );
  NAND U10622 ( .A(n9667), .B(n37764), .Z(n9485) );
  NAND U10623 ( .A(n9486), .B(n9485), .Z(n9642) );
  XOR U10624 ( .A(b[31]), .B(n9873), .Z(n9670) );
  NANDN U10625 ( .A(n9670), .B(n38552), .Z(n9489) );
  NANDN U10626 ( .A(n9487), .B(n38553), .Z(n9488) );
  AND U10627 ( .A(n9489), .B(n9488), .Z(n9640) );
  OR U10628 ( .A(n9490), .B(n36105), .Z(n9492) );
  XNOR U10629 ( .A(b[3]), .B(a[72]), .Z(n9673) );
  NANDN U10630 ( .A(n9673), .B(n36107), .Z(n9491) );
  AND U10631 ( .A(n9492), .B(n9491), .Z(n9641) );
  XOR U10632 ( .A(n9642), .B(n9643), .Z(n9689) );
  XOR U10633 ( .A(n9688), .B(n9689), .Z(n9690) );
  XNOR U10634 ( .A(n9691), .B(n9690), .Z(n9618) );
  NANDN U10635 ( .A(n9494), .B(n9493), .Z(n9498) );
  OR U10636 ( .A(n9496), .B(n9495), .Z(n9497) );
  NAND U10637 ( .A(n9498), .B(n9497), .Z(n9619) );
  XNOR U10638 ( .A(n9618), .B(n9619), .Z(n9620) );
  NANDN U10639 ( .A(n9500), .B(n9499), .Z(n9504) );
  NAND U10640 ( .A(n9502), .B(n9501), .Z(n9503) );
  NAND U10641 ( .A(n9504), .B(n9503), .Z(n9679) );
  NANDN U10642 ( .A(n9506), .B(n9505), .Z(n9510) );
  NAND U10643 ( .A(n9508), .B(n9507), .Z(n9509) );
  NAND U10644 ( .A(n9510), .B(n9509), .Z(n9676) );
  OR U10645 ( .A(n9512), .B(n9511), .Z(n9516) );
  NANDN U10646 ( .A(n9514), .B(n9513), .Z(n9515) );
  NAND U10647 ( .A(n9516), .B(n9515), .Z(n9677) );
  XNOR U10648 ( .A(n9676), .B(n9677), .Z(n9678) );
  XOR U10649 ( .A(n9679), .B(n9678), .Z(n9621) );
  XNOR U10650 ( .A(n9620), .B(n9621), .Z(n9745) );
  OR U10651 ( .A(n9518), .B(n9517), .Z(n9522) );
  NANDN U10652 ( .A(n9520), .B(n9519), .Z(n9521) );
  NAND U10653 ( .A(n9522), .B(n9521), .Z(n9743) );
  NANDN U10654 ( .A(n9524), .B(n9523), .Z(n9528) );
  NANDN U10655 ( .A(n9526), .B(n9525), .Z(n9527) );
  NAND U10656 ( .A(n9528), .B(n9527), .Z(n9625) );
  NANDN U10657 ( .A(n9530), .B(n9529), .Z(n9534) );
  NAND U10658 ( .A(n9532), .B(n9531), .Z(n9533) );
  NAND U10659 ( .A(n9534), .B(n9533), .Z(n9622) );
  XNOR U10660 ( .A(b[9]), .B(a[66]), .Z(n9706) );
  NANDN U10661 ( .A(n9706), .B(n36925), .Z(n9537) );
  NANDN U10662 ( .A(n9535), .B(n36926), .Z(n9536) );
  NAND U10663 ( .A(n9537), .B(n9536), .Z(n9648) );
  XNOR U10664 ( .A(b[15]), .B(a[60]), .Z(n9709) );
  OR U10665 ( .A(n9709), .B(n37665), .Z(n9540) );
  NANDN U10666 ( .A(n9538), .B(n37604), .Z(n9539) );
  AND U10667 ( .A(n9540), .B(n9539), .Z(n9646) );
  XOR U10668 ( .A(b[21]), .B(n11319), .Z(n9712) );
  NANDN U10669 ( .A(n9712), .B(n38101), .Z(n9543) );
  NANDN U10670 ( .A(n9541), .B(n38102), .Z(n9542) );
  AND U10671 ( .A(n9543), .B(n9542), .Z(n9647) );
  XOR U10672 ( .A(n9648), .B(n9649), .Z(n9637) );
  XNOR U10673 ( .A(b[11]), .B(a[64]), .Z(n9715) );
  OR U10674 ( .A(n9715), .B(n37311), .Z(n9546) );
  NANDN U10675 ( .A(n9544), .B(n37218), .Z(n9545) );
  NAND U10676 ( .A(n9546), .B(n9545), .Z(n9635) );
  XOR U10677 ( .A(n1053), .B(a[62]), .Z(n9718) );
  NANDN U10678 ( .A(n9718), .B(n37424), .Z(n9549) );
  NANDN U10679 ( .A(n9547), .B(n37425), .Z(n9548) );
  NAND U10680 ( .A(n9549), .B(n9548), .Z(n9634) );
  XOR U10681 ( .A(n9637), .B(n9636), .Z(n9631) );
  NANDN U10682 ( .A(n1049), .B(a[74]), .Z(n9550) );
  XNOR U10683 ( .A(b[1]), .B(n9550), .Z(n9552) );
  NANDN U10684 ( .A(b[0]), .B(a[73]), .Z(n9551) );
  AND U10685 ( .A(n9552), .B(n9551), .Z(n9654) );
  NAND U10686 ( .A(n38490), .B(n9553), .Z(n9555) );
  XNOR U10687 ( .A(n1058), .B(a[46]), .Z(n9724) );
  NANDN U10688 ( .A(n1048), .B(n9724), .Z(n9554) );
  NAND U10689 ( .A(n9555), .B(n9554), .Z(n9652) );
  NANDN U10690 ( .A(n1059), .B(a[42]), .Z(n9653) );
  XNOR U10691 ( .A(n9652), .B(n9653), .Z(n9655) );
  XNOR U10692 ( .A(n9654), .B(n9655), .Z(n9629) );
  NANDN U10693 ( .A(n9556), .B(n38205), .Z(n9558) );
  XNOR U10694 ( .A(b[23]), .B(a[52]), .Z(n9727) );
  OR U10695 ( .A(n9727), .B(n38268), .Z(n9557) );
  NAND U10696 ( .A(n9558), .B(n9557), .Z(n9697) );
  XOR U10697 ( .A(b[7]), .B(a[68]), .Z(n9730) );
  NAND U10698 ( .A(n9730), .B(n36701), .Z(n9561) );
  NANDN U10699 ( .A(n9559), .B(n36702), .Z(n9560) );
  NAND U10700 ( .A(n9561), .B(n9560), .Z(n9694) );
  XNOR U10701 ( .A(b[25]), .B(a[50]), .Z(n9733) );
  NANDN U10702 ( .A(n9733), .B(n38325), .Z(n9564) );
  NAND U10703 ( .A(n9562), .B(n38326), .Z(n9563) );
  AND U10704 ( .A(n9564), .B(n9563), .Z(n9695) );
  XNOR U10705 ( .A(n9694), .B(n9695), .Z(n9696) );
  XOR U10706 ( .A(n9697), .B(n9696), .Z(n9628) );
  XNOR U10707 ( .A(n9631), .B(n9630), .Z(n9685) );
  NANDN U10708 ( .A(n9566), .B(n9565), .Z(n9570) );
  NAND U10709 ( .A(n9568), .B(n9567), .Z(n9569) );
  NAND U10710 ( .A(n9570), .B(n9569), .Z(n9683) );
  NANDN U10711 ( .A(n9572), .B(n9571), .Z(n9576) );
  NAND U10712 ( .A(n9574), .B(n9573), .Z(n9575) );
  AND U10713 ( .A(n9576), .B(n9575), .Z(n9682) );
  XNOR U10714 ( .A(n9683), .B(n9682), .Z(n9684) );
  XNOR U10715 ( .A(n9685), .B(n9684), .Z(n9623) );
  XNOR U10716 ( .A(n9622), .B(n9623), .Z(n9624) );
  XOR U10717 ( .A(n9625), .B(n9624), .Z(n9742) );
  XOR U10718 ( .A(n9743), .B(n9742), .Z(n9744) );
  XNOR U10719 ( .A(n9745), .B(n9744), .Z(n9739) );
  NANDN U10720 ( .A(n9578), .B(n9577), .Z(n9582) );
  NAND U10721 ( .A(n9580), .B(n9579), .Z(n9581) );
  NAND U10722 ( .A(n9582), .B(n9581), .Z(n9737) );
  NAND U10723 ( .A(n9584), .B(n9583), .Z(n9588) );
  NANDN U10724 ( .A(n9586), .B(n9585), .Z(n9587) );
  AND U10725 ( .A(n9588), .B(n9587), .Z(n9736) );
  XNOR U10726 ( .A(n9737), .B(n9736), .Z(n9738) );
  XOR U10727 ( .A(n9739), .B(n9738), .Z(n9614) );
  NANDN U10728 ( .A(n9590), .B(n9589), .Z(n9594) );
  NAND U10729 ( .A(n9592), .B(n9591), .Z(n9593) );
  NAND U10730 ( .A(n9594), .B(n9593), .Z(n9612) );
  NANDN U10731 ( .A(n9596), .B(n9595), .Z(n9600) );
  NANDN U10732 ( .A(n9598), .B(n9597), .Z(n9599) );
  NAND U10733 ( .A(n9600), .B(n9599), .Z(n9613) );
  XNOR U10734 ( .A(n9612), .B(n9613), .Z(n9615) );
  XOR U10735 ( .A(n9614), .B(n9615), .Z(n9606) );
  XOR U10736 ( .A(n9607), .B(n9606), .Z(n9608) );
  XNOR U10737 ( .A(n9609), .B(n9608), .Z(n9748) );
  XNOR U10738 ( .A(n9748), .B(sreg[298]), .Z(n9750) );
  NAND U10739 ( .A(n9601), .B(sreg[297]), .Z(n9605) );
  OR U10740 ( .A(n9603), .B(n9602), .Z(n9604) );
  AND U10741 ( .A(n9605), .B(n9604), .Z(n9749) );
  XOR U10742 ( .A(n9750), .B(n9749), .Z(c[298]) );
  NAND U10743 ( .A(n9607), .B(n9606), .Z(n9611) );
  NAND U10744 ( .A(n9609), .B(n9608), .Z(n9610) );
  NAND U10745 ( .A(n9611), .B(n9610), .Z(n9756) );
  NANDN U10746 ( .A(n9613), .B(n9612), .Z(n9617) );
  NAND U10747 ( .A(n9615), .B(n9614), .Z(n9616) );
  NAND U10748 ( .A(n9617), .B(n9616), .Z(n9754) );
  NANDN U10749 ( .A(n9623), .B(n9622), .Z(n9627) );
  NAND U10750 ( .A(n9625), .B(n9624), .Z(n9626) );
  NAND U10751 ( .A(n9627), .B(n9626), .Z(n9772) );
  XNOR U10752 ( .A(n9771), .B(n9772), .Z(n9773) );
  NANDN U10753 ( .A(n9629), .B(n9628), .Z(n9633) );
  NANDN U10754 ( .A(n9631), .B(n9630), .Z(n9632) );
  NAND U10755 ( .A(n9633), .B(n9632), .Z(n9889) );
  OR U10756 ( .A(n9635), .B(n9634), .Z(n9639) );
  NAND U10757 ( .A(n9637), .B(n9636), .Z(n9638) );
  NAND U10758 ( .A(n9639), .B(n9638), .Z(n9827) );
  OR U10759 ( .A(n9641), .B(n9640), .Z(n9645) );
  NANDN U10760 ( .A(n9643), .B(n9642), .Z(n9644) );
  NAND U10761 ( .A(n9645), .B(n9644), .Z(n9826) );
  OR U10762 ( .A(n9647), .B(n9646), .Z(n9651) );
  NANDN U10763 ( .A(n9649), .B(n9648), .Z(n9650) );
  NAND U10764 ( .A(n9651), .B(n9650), .Z(n9825) );
  XOR U10765 ( .A(n9827), .B(n9828), .Z(n9886) );
  NANDN U10766 ( .A(n9653), .B(n9652), .Z(n9657) );
  NAND U10767 ( .A(n9655), .B(n9654), .Z(n9656) );
  NAND U10768 ( .A(n9657), .B(n9656), .Z(n9840) );
  XNOR U10769 ( .A(b[19]), .B(a[57]), .Z(n9783) );
  NANDN U10770 ( .A(n9783), .B(n37934), .Z(n9660) );
  NANDN U10771 ( .A(n9658), .B(n37935), .Z(n9659) );
  NAND U10772 ( .A(n9660), .B(n9659), .Z(n9852) );
  XOR U10773 ( .A(b[27]), .B(a[49]), .Z(n9786) );
  NAND U10774 ( .A(n38423), .B(n9786), .Z(n9663) );
  NAND U10775 ( .A(n9661), .B(n38424), .Z(n9662) );
  NAND U10776 ( .A(n9663), .B(n9662), .Z(n9849) );
  XNOR U10777 ( .A(b[5]), .B(a[71]), .Z(n9789) );
  NANDN U10778 ( .A(n9789), .B(n36587), .Z(n9666) );
  NANDN U10779 ( .A(n9664), .B(n36588), .Z(n9665) );
  AND U10780 ( .A(n9666), .B(n9665), .Z(n9850) );
  XNOR U10781 ( .A(n9849), .B(n9850), .Z(n9851) );
  XNOR U10782 ( .A(n9852), .B(n9851), .Z(n9838) );
  NAND U10783 ( .A(n9667), .B(n37762), .Z(n9669) );
  XNOR U10784 ( .A(b[17]), .B(a[59]), .Z(n9792) );
  NANDN U10785 ( .A(n9792), .B(n37764), .Z(n9668) );
  NAND U10786 ( .A(n9669), .B(n9668), .Z(n9810) );
  XNOR U10787 ( .A(b[31]), .B(a[45]), .Z(n9795) );
  NANDN U10788 ( .A(n9795), .B(n38552), .Z(n9672) );
  NANDN U10789 ( .A(n9670), .B(n38553), .Z(n9671) );
  NAND U10790 ( .A(n9672), .B(n9671), .Z(n9807) );
  OR U10791 ( .A(n9673), .B(n36105), .Z(n9675) );
  XNOR U10792 ( .A(b[3]), .B(a[73]), .Z(n9798) );
  NANDN U10793 ( .A(n9798), .B(n36107), .Z(n9674) );
  AND U10794 ( .A(n9675), .B(n9674), .Z(n9808) );
  XNOR U10795 ( .A(n9807), .B(n9808), .Z(n9809) );
  XOR U10796 ( .A(n9810), .B(n9809), .Z(n9837) );
  XNOR U10797 ( .A(n9838), .B(n9837), .Z(n9839) );
  XNOR U10798 ( .A(n9840), .B(n9839), .Z(n9887) );
  XNOR U10799 ( .A(n9886), .B(n9887), .Z(n9888) );
  XNOR U10800 ( .A(n9889), .B(n9888), .Z(n9768) );
  NANDN U10801 ( .A(n9677), .B(n9676), .Z(n9681) );
  NANDN U10802 ( .A(n9679), .B(n9678), .Z(n9680) );
  NAND U10803 ( .A(n9681), .B(n9680), .Z(n9765) );
  NANDN U10804 ( .A(n9683), .B(n9682), .Z(n9687) );
  NANDN U10805 ( .A(n9685), .B(n9684), .Z(n9686) );
  NAND U10806 ( .A(n9687), .B(n9686), .Z(n9893) );
  OR U10807 ( .A(n9689), .B(n9688), .Z(n9693) );
  NAND U10808 ( .A(n9691), .B(n9690), .Z(n9692) );
  NAND U10809 ( .A(n9693), .B(n9692), .Z(n9891) );
  NANDN U10810 ( .A(n9695), .B(n9694), .Z(n9699) );
  NAND U10811 ( .A(n9697), .B(n9696), .Z(n9698) );
  NAND U10812 ( .A(n9699), .B(n9698), .Z(n9831) );
  NANDN U10813 ( .A(n9701), .B(n9700), .Z(n9705) );
  NAND U10814 ( .A(n9703), .B(n9702), .Z(n9704) );
  AND U10815 ( .A(n9705), .B(n9704), .Z(n9832) );
  XNOR U10816 ( .A(n9831), .B(n9832), .Z(n9833) );
  XOR U10817 ( .A(b[9]), .B(n13219), .Z(n9855) );
  NANDN U10818 ( .A(n9855), .B(n36925), .Z(n9708) );
  NANDN U10819 ( .A(n9706), .B(n36926), .Z(n9707) );
  NAND U10820 ( .A(n9708), .B(n9707), .Z(n9815) );
  XNOR U10821 ( .A(b[15]), .B(a[61]), .Z(n9858) );
  OR U10822 ( .A(n9858), .B(n37665), .Z(n9711) );
  NANDN U10823 ( .A(n9709), .B(n37604), .Z(n9710) );
  AND U10824 ( .A(n9711), .B(n9710), .Z(n9813) );
  XNOR U10825 ( .A(b[21]), .B(a[55]), .Z(n9861) );
  NANDN U10826 ( .A(n9861), .B(n38101), .Z(n9714) );
  NANDN U10827 ( .A(n9712), .B(n38102), .Z(n9713) );
  AND U10828 ( .A(n9714), .B(n9713), .Z(n9814) );
  XOR U10829 ( .A(n9815), .B(n9816), .Z(n9804) );
  XNOR U10830 ( .A(b[11]), .B(a[65]), .Z(n9864) );
  OR U10831 ( .A(n9864), .B(n37311), .Z(n9717) );
  NANDN U10832 ( .A(n9715), .B(n37218), .Z(n9716) );
  NAND U10833 ( .A(n9717), .B(n9716), .Z(n9802) );
  XOR U10834 ( .A(n1053), .B(a[63]), .Z(n9867) );
  NANDN U10835 ( .A(n9867), .B(n37424), .Z(n9720) );
  NANDN U10836 ( .A(n9718), .B(n37425), .Z(n9719) );
  AND U10837 ( .A(n9720), .B(n9719), .Z(n9801) );
  XNOR U10838 ( .A(n9802), .B(n9801), .Z(n9803) );
  XOR U10839 ( .A(n9804), .B(n9803), .Z(n9821) );
  NANDN U10840 ( .A(n1049), .B(a[75]), .Z(n9721) );
  XNOR U10841 ( .A(b[1]), .B(n9721), .Z(n9723) );
  NANDN U10842 ( .A(b[0]), .B(a[74]), .Z(n9722) );
  AND U10843 ( .A(n9723), .B(n9722), .Z(n9779) );
  NAND U10844 ( .A(n38490), .B(n9724), .Z(n9726) );
  XNOR U10845 ( .A(b[29]), .B(a[47]), .Z(n9874) );
  OR U10846 ( .A(n9874), .B(n1048), .Z(n9725) );
  NAND U10847 ( .A(n9726), .B(n9725), .Z(n9777) );
  NANDN U10848 ( .A(n1059), .B(a[43]), .Z(n9778) );
  XNOR U10849 ( .A(n9777), .B(n9778), .Z(n9780) );
  XOR U10850 ( .A(n9779), .B(n9780), .Z(n9819) );
  NANDN U10851 ( .A(n9727), .B(n38205), .Z(n9729) );
  XNOR U10852 ( .A(b[23]), .B(a[53]), .Z(n9877) );
  OR U10853 ( .A(n9877), .B(n38268), .Z(n9728) );
  NAND U10854 ( .A(n9729), .B(n9728), .Z(n9846) );
  XOR U10855 ( .A(b[7]), .B(a[69]), .Z(n9880) );
  NAND U10856 ( .A(n9880), .B(n36701), .Z(n9732) );
  NAND U10857 ( .A(n9730), .B(n36702), .Z(n9731) );
  NAND U10858 ( .A(n9732), .B(n9731), .Z(n9843) );
  XOR U10859 ( .A(b[25]), .B(a[51]), .Z(n9883) );
  NAND U10860 ( .A(n9883), .B(n38325), .Z(n9735) );
  NANDN U10861 ( .A(n9733), .B(n38326), .Z(n9734) );
  AND U10862 ( .A(n9735), .B(n9734), .Z(n9844) );
  XNOR U10863 ( .A(n9843), .B(n9844), .Z(n9845) );
  XNOR U10864 ( .A(n9846), .B(n9845), .Z(n9820) );
  XOR U10865 ( .A(n9819), .B(n9820), .Z(n9822) );
  XNOR U10866 ( .A(n9821), .B(n9822), .Z(n9834) );
  XNOR U10867 ( .A(n9833), .B(n9834), .Z(n9890) );
  XNOR U10868 ( .A(n9891), .B(n9890), .Z(n9892) );
  XOR U10869 ( .A(n9893), .B(n9892), .Z(n9766) );
  XNOR U10870 ( .A(n9765), .B(n9766), .Z(n9767) );
  XOR U10871 ( .A(n9768), .B(n9767), .Z(n9774) );
  XOR U10872 ( .A(n9773), .B(n9774), .Z(n9761) );
  NANDN U10873 ( .A(n9737), .B(n9736), .Z(n9741) );
  NAND U10874 ( .A(n9739), .B(n9738), .Z(n9740) );
  NAND U10875 ( .A(n9741), .B(n9740), .Z(n9759) );
  NANDN U10876 ( .A(n9743), .B(n9742), .Z(n9747) );
  OR U10877 ( .A(n9745), .B(n9744), .Z(n9746) );
  NAND U10878 ( .A(n9747), .B(n9746), .Z(n9760) );
  XNOR U10879 ( .A(n9759), .B(n9760), .Z(n9762) );
  XOR U10880 ( .A(n9761), .B(n9762), .Z(n9753) );
  XOR U10881 ( .A(n9754), .B(n9753), .Z(n9755) );
  XNOR U10882 ( .A(n9756), .B(n9755), .Z(n9896) );
  XNOR U10883 ( .A(n9896), .B(sreg[299]), .Z(n9898) );
  NAND U10884 ( .A(n9748), .B(sreg[298]), .Z(n9752) );
  OR U10885 ( .A(n9750), .B(n9749), .Z(n9751) );
  AND U10886 ( .A(n9752), .B(n9751), .Z(n9897) );
  XOR U10887 ( .A(n9898), .B(n9897), .Z(c[299]) );
  NAND U10888 ( .A(n9754), .B(n9753), .Z(n9758) );
  NAND U10889 ( .A(n9756), .B(n9755), .Z(n9757) );
  NAND U10890 ( .A(n9758), .B(n9757), .Z(n9904) );
  NANDN U10891 ( .A(n9760), .B(n9759), .Z(n9764) );
  NAND U10892 ( .A(n9762), .B(n9761), .Z(n9763) );
  NAND U10893 ( .A(n9764), .B(n9763), .Z(n9902) );
  NANDN U10894 ( .A(n9766), .B(n9765), .Z(n9770) );
  NAND U10895 ( .A(n9768), .B(n9767), .Z(n9769) );
  NAND U10896 ( .A(n9770), .B(n9769), .Z(n9907) );
  NANDN U10897 ( .A(n9772), .B(n9771), .Z(n9776) );
  NAND U10898 ( .A(n9774), .B(n9773), .Z(n9775) );
  AND U10899 ( .A(n9776), .B(n9775), .Z(n9908) );
  XNOR U10900 ( .A(n9907), .B(n9908), .Z(n9909) );
  NANDN U10901 ( .A(n9778), .B(n9777), .Z(n9782) );
  NAND U10902 ( .A(n9780), .B(n9779), .Z(n9781) );
  NAND U10903 ( .A(n9782), .B(n9781), .Z(n9988) );
  XNOR U10904 ( .A(b[19]), .B(a[58]), .Z(n9955) );
  NANDN U10905 ( .A(n9955), .B(n37934), .Z(n9785) );
  NANDN U10906 ( .A(n9783), .B(n37935), .Z(n9784) );
  NAND U10907 ( .A(n9785), .B(n9784), .Z(n10000) );
  XNOR U10908 ( .A(b[27]), .B(a[50]), .Z(n9958) );
  NANDN U10909 ( .A(n9958), .B(n38423), .Z(n9788) );
  NAND U10910 ( .A(n9786), .B(n38424), .Z(n9787) );
  NAND U10911 ( .A(n9788), .B(n9787), .Z(n9997) );
  XNOR U10912 ( .A(b[5]), .B(a[72]), .Z(n9961) );
  NANDN U10913 ( .A(n9961), .B(n36587), .Z(n9791) );
  NANDN U10914 ( .A(n9789), .B(n36588), .Z(n9790) );
  AND U10915 ( .A(n9791), .B(n9790), .Z(n9998) );
  XNOR U10916 ( .A(n9997), .B(n9998), .Z(n9999) );
  XNOR U10917 ( .A(n10000), .B(n9999), .Z(n9985) );
  NANDN U10918 ( .A(n9792), .B(n37762), .Z(n9794) );
  XOR U10919 ( .A(b[17]), .B(a[60]), .Z(n9964) );
  NAND U10920 ( .A(n9964), .B(n37764), .Z(n9793) );
  NAND U10921 ( .A(n9794), .B(n9793), .Z(n9939) );
  XNOR U10922 ( .A(b[31]), .B(a[46]), .Z(n9967) );
  NANDN U10923 ( .A(n9967), .B(n38552), .Z(n9797) );
  NANDN U10924 ( .A(n9795), .B(n38553), .Z(n9796) );
  AND U10925 ( .A(n9797), .B(n9796), .Z(n9937) );
  OR U10926 ( .A(n9798), .B(n36105), .Z(n9800) );
  XNOR U10927 ( .A(b[3]), .B(a[74]), .Z(n9970) );
  NANDN U10928 ( .A(n9970), .B(n36107), .Z(n9799) );
  AND U10929 ( .A(n9800), .B(n9799), .Z(n9938) );
  XOR U10930 ( .A(n9939), .B(n9940), .Z(n9986) );
  XOR U10931 ( .A(n9985), .B(n9986), .Z(n9987) );
  XNOR U10932 ( .A(n9988), .B(n9987), .Z(n10033) );
  NANDN U10933 ( .A(n9802), .B(n9801), .Z(n9806) );
  NAND U10934 ( .A(n9804), .B(n9803), .Z(n9805) );
  NAND U10935 ( .A(n9806), .B(n9805), .Z(n9976) );
  NANDN U10936 ( .A(n9808), .B(n9807), .Z(n9812) );
  NAND U10937 ( .A(n9810), .B(n9809), .Z(n9811) );
  NAND U10938 ( .A(n9812), .B(n9811), .Z(n9974) );
  OR U10939 ( .A(n9814), .B(n9813), .Z(n9818) );
  NANDN U10940 ( .A(n9816), .B(n9815), .Z(n9817) );
  NAND U10941 ( .A(n9818), .B(n9817), .Z(n9973) );
  XNOR U10942 ( .A(n9976), .B(n9975), .Z(n10034) );
  XOR U10943 ( .A(n10033), .B(n10034), .Z(n10036) );
  NANDN U10944 ( .A(n9820), .B(n9819), .Z(n9824) );
  OR U10945 ( .A(n9822), .B(n9821), .Z(n9823) );
  NAND U10946 ( .A(n9824), .B(n9823), .Z(n10035) );
  XOR U10947 ( .A(n10036), .B(n10035), .Z(n9921) );
  OR U10948 ( .A(n9826), .B(n9825), .Z(n9830) );
  NANDN U10949 ( .A(n9828), .B(n9827), .Z(n9829) );
  NAND U10950 ( .A(n9830), .B(n9829), .Z(n9920) );
  NANDN U10951 ( .A(n9832), .B(n9831), .Z(n9836) );
  NANDN U10952 ( .A(n9834), .B(n9833), .Z(n9835) );
  NAND U10953 ( .A(n9836), .B(n9835), .Z(n10041) );
  NANDN U10954 ( .A(n9838), .B(n9837), .Z(n9842) );
  NAND U10955 ( .A(n9840), .B(n9839), .Z(n9841) );
  NAND U10956 ( .A(n9842), .B(n9841), .Z(n10040) );
  NANDN U10957 ( .A(n9844), .B(n9843), .Z(n9848) );
  NAND U10958 ( .A(n9846), .B(n9845), .Z(n9847) );
  NAND U10959 ( .A(n9848), .B(n9847), .Z(n9979) );
  NANDN U10960 ( .A(n9850), .B(n9849), .Z(n9854) );
  NAND U10961 ( .A(n9852), .B(n9851), .Z(n9853) );
  AND U10962 ( .A(n9854), .B(n9853), .Z(n9980) );
  XNOR U10963 ( .A(n9979), .B(n9980), .Z(n9981) );
  XNOR U10964 ( .A(n1052), .B(a[68]), .Z(n10003) );
  NAND U10965 ( .A(n36925), .B(n10003), .Z(n9857) );
  NANDN U10966 ( .A(n9855), .B(n36926), .Z(n9856) );
  NAND U10967 ( .A(n9857), .B(n9856), .Z(n9945) );
  XOR U10968 ( .A(b[15]), .B(n12493), .Z(n10006) );
  OR U10969 ( .A(n10006), .B(n37665), .Z(n9860) );
  NANDN U10970 ( .A(n9858), .B(n37604), .Z(n9859) );
  AND U10971 ( .A(n9860), .B(n9859), .Z(n9943) );
  XNOR U10972 ( .A(n1056), .B(a[56]), .Z(n10009) );
  NAND U10973 ( .A(n10009), .B(n38101), .Z(n9863) );
  NANDN U10974 ( .A(n9861), .B(n38102), .Z(n9862) );
  AND U10975 ( .A(n9863), .B(n9862), .Z(n9944) );
  XOR U10976 ( .A(n9945), .B(n9946), .Z(n9934) );
  XNOR U10977 ( .A(b[11]), .B(a[66]), .Z(n10012) );
  OR U10978 ( .A(n10012), .B(n37311), .Z(n9866) );
  NANDN U10979 ( .A(n9864), .B(n37218), .Z(n9865) );
  NAND U10980 ( .A(n9866), .B(n9865), .Z(n9932) );
  XOR U10981 ( .A(n1053), .B(a[64]), .Z(n10015) );
  NANDN U10982 ( .A(n10015), .B(n37424), .Z(n9869) );
  NANDN U10983 ( .A(n9867), .B(n37425), .Z(n9868) );
  NAND U10984 ( .A(n9869), .B(n9868), .Z(n9931) );
  XOR U10985 ( .A(n9934), .B(n9933), .Z(n9928) );
  NANDN U10986 ( .A(n1049), .B(a[76]), .Z(n9870) );
  XNOR U10987 ( .A(b[1]), .B(n9870), .Z(n9872) );
  NANDN U10988 ( .A(b[0]), .B(a[75]), .Z(n9871) );
  AND U10989 ( .A(n9872), .B(n9871), .Z(n9952) );
  ANDN U10990 ( .B(b[31]), .A(n9873), .Z(n9949) );
  NANDN U10991 ( .A(n9874), .B(n38490), .Z(n9876) );
  XNOR U10992 ( .A(n1058), .B(a[48]), .Z(n10021) );
  NANDN U10993 ( .A(n1048), .B(n10021), .Z(n9875) );
  NAND U10994 ( .A(n9876), .B(n9875), .Z(n9950) );
  XOR U10995 ( .A(n9949), .B(n9950), .Z(n9951) );
  XNOR U10996 ( .A(n9952), .B(n9951), .Z(n9925) );
  NANDN U10997 ( .A(n9877), .B(n38205), .Z(n9879) );
  XOR U10998 ( .A(b[23]), .B(n11319), .Z(n10024) );
  OR U10999 ( .A(n10024), .B(n38268), .Z(n9878) );
  NAND U11000 ( .A(n9879), .B(n9878), .Z(n9994) );
  XOR U11001 ( .A(b[7]), .B(a[70]), .Z(n10027) );
  NAND U11002 ( .A(n10027), .B(n36701), .Z(n9882) );
  NAND U11003 ( .A(n9880), .B(n36702), .Z(n9881) );
  NAND U11004 ( .A(n9882), .B(n9881), .Z(n9991) );
  XOR U11005 ( .A(b[25]), .B(a[52]), .Z(n10030) );
  NAND U11006 ( .A(n10030), .B(n38325), .Z(n9885) );
  NAND U11007 ( .A(n9883), .B(n38326), .Z(n9884) );
  AND U11008 ( .A(n9885), .B(n9884), .Z(n9992) );
  XNOR U11009 ( .A(n9991), .B(n9992), .Z(n9993) );
  XNOR U11010 ( .A(n9994), .B(n9993), .Z(n9926) );
  XOR U11011 ( .A(n9928), .B(n9927), .Z(n9982) );
  XNOR U11012 ( .A(n9981), .B(n9982), .Z(n10039) );
  XNOR U11013 ( .A(n10040), .B(n10039), .Z(n10042) );
  XNOR U11014 ( .A(n10041), .B(n10042), .Z(n9919) );
  XOR U11015 ( .A(n9920), .B(n9919), .Z(n9922) );
  NAND U11016 ( .A(n9891), .B(n9890), .Z(n9895) );
  OR U11017 ( .A(n9893), .B(n9892), .Z(n9894) );
  AND U11018 ( .A(n9895), .B(n9894), .Z(n9913) );
  XNOR U11019 ( .A(n9914), .B(n9913), .Z(n9915) );
  XOR U11020 ( .A(n9916), .B(n9915), .Z(n9910) );
  XOR U11021 ( .A(n9909), .B(n9910), .Z(n9901) );
  XOR U11022 ( .A(n9902), .B(n9901), .Z(n9903) );
  XNOR U11023 ( .A(n9904), .B(n9903), .Z(n10045) );
  XNOR U11024 ( .A(n10045), .B(sreg[300]), .Z(n10047) );
  NAND U11025 ( .A(n9896), .B(sreg[299]), .Z(n9900) );
  OR U11026 ( .A(n9898), .B(n9897), .Z(n9899) );
  AND U11027 ( .A(n9900), .B(n9899), .Z(n10046) );
  XOR U11028 ( .A(n10047), .B(n10046), .Z(c[300]) );
  NAND U11029 ( .A(n9902), .B(n9901), .Z(n9906) );
  NAND U11030 ( .A(n9904), .B(n9903), .Z(n9905) );
  NAND U11031 ( .A(n9906), .B(n9905), .Z(n10053) );
  NANDN U11032 ( .A(n9908), .B(n9907), .Z(n9912) );
  NAND U11033 ( .A(n9910), .B(n9909), .Z(n9911) );
  NAND U11034 ( .A(n9912), .B(n9911), .Z(n10051) );
  NANDN U11035 ( .A(n9914), .B(n9913), .Z(n9918) );
  NAND U11036 ( .A(n9916), .B(n9915), .Z(n9917) );
  NAND U11037 ( .A(n9918), .B(n9917), .Z(n10056) );
  NANDN U11038 ( .A(n9920), .B(n9919), .Z(n9924) );
  OR U11039 ( .A(n9922), .B(n9921), .Z(n9923) );
  NAND U11040 ( .A(n9924), .B(n9923), .Z(n10057) );
  XNOR U11041 ( .A(n10056), .B(n10057), .Z(n10058) );
  OR U11042 ( .A(n9926), .B(n9925), .Z(n9930) );
  NANDN U11043 ( .A(n9928), .B(n9927), .Z(n9929) );
  NAND U11044 ( .A(n9930), .B(n9929), .Z(n10183) );
  OR U11045 ( .A(n9932), .B(n9931), .Z(n9936) );
  NAND U11046 ( .A(n9934), .B(n9933), .Z(n9935) );
  NAND U11047 ( .A(n9936), .B(n9935), .Z(n10122) );
  OR U11048 ( .A(n9938), .B(n9937), .Z(n9942) );
  NANDN U11049 ( .A(n9940), .B(n9939), .Z(n9941) );
  NAND U11050 ( .A(n9942), .B(n9941), .Z(n10121) );
  OR U11051 ( .A(n9944), .B(n9943), .Z(n9948) );
  NANDN U11052 ( .A(n9946), .B(n9945), .Z(n9947) );
  NAND U11053 ( .A(n9948), .B(n9947), .Z(n10120) );
  XOR U11054 ( .A(n10122), .B(n10123), .Z(n10181) );
  OR U11055 ( .A(n9950), .B(n9949), .Z(n9954) );
  NANDN U11056 ( .A(n9952), .B(n9951), .Z(n9953) );
  NAND U11057 ( .A(n9954), .B(n9953), .Z(n10134) );
  XOR U11058 ( .A(b[19]), .B(n12056), .Z(n10080) );
  NANDN U11059 ( .A(n10080), .B(n37934), .Z(n9957) );
  NANDN U11060 ( .A(n9955), .B(n37935), .Z(n9956) );
  NAND U11061 ( .A(n9957), .B(n9956), .Z(n10147) );
  XOR U11062 ( .A(b[27]), .B(a[51]), .Z(n10083) );
  NAND U11063 ( .A(n38423), .B(n10083), .Z(n9960) );
  NANDN U11064 ( .A(n9958), .B(n38424), .Z(n9959) );
  NAND U11065 ( .A(n9960), .B(n9959), .Z(n10144) );
  XNOR U11066 ( .A(b[5]), .B(a[73]), .Z(n10086) );
  NANDN U11067 ( .A(n10086), .B(n36587), .Z(n9963) );
  NANDN U11068 ( .A(n9961), .B(n36588), .Z(n9962) );
  AND U11069 ( .A(n9963), .B(n9962), .Z(n10145) );
  XNOR U11070 ( .A(n10144), .B(n10145), .Z(n10146) );
  XNOR U11071 ( .A(n10147), .B(n10146), .Z(n10133) );
  NAND U11072 ( .A(n9964), .B(n37762), .Z(n9966) );
  XOR U11073 ( .A(b[17]), .B(a[61]), .Z(n10089) );
  NAND U11074 ( .A(n10089), .B(n37764), .Z(n9965) );
  NAND U11075 ( .A(n9966), .B(n9965), .Z(n10107) );
  XNOR U11076 ( .A(b[31]), .B(a[47]), .Z(n10092) );
  NANDN U11077 ( .A(n10092), .B(n38552), .Z(n9969) );
  NANDN U11078 ( .A(n9967), .B(n38553), .Z(n9968) );
  NAND U11079 ( .A(n9969), .B(n9968), .Z(n10104) );
  OR U11080 ( .A(n9970), .B(n36105), .Z(n9972) );
  XNOR U11081 ( .A(b[3]), .B(a[75]), .Z(n10095) );
  NANDN U11082 ( .A(n10095), .B(n36107), .Z(n9971) );
  AND U11083 ( .A(n9972), .B(n9971), .Z(n10105) );
  XNOR U11084 ( .A(n10104), .B(n10105), .Z(n10106) );
  XOR U11085 ( .A(n10107), .B(n10106), .Z(n10132) );
  XOR U11086 ( .A(n10133), .B(n10132), .Z(n10135) );
  XOR U11087 ( .A(n10134), .B(n10135), .Z(n10180) );
  XOR U11088 ( .A(n10181), .B(n10180), .Z(n10182) );
  XNOR U11089 ( .A(n10183), .B(n10182), .Z(n10071) );
  OR U11090 ( .A(n9974), .B(n9973), .Z(n9978) );
  NAND U11091 ( .A(n9976), .B(n9975), .Z(n9977) );
  NAND U11092 ( .A(n9978), .B(n9977), .Z(n10069) );
  NANDN U11093 ( .A(n9980), .B(n9979), .Z(n9984) );
  NANDN U11094 ( .A(n9982), .B(n9981), .Z(n9983) );
  NAND U11095 ( .A(n9984), .B(n9983), .Z(n10188) );
  OR U11096 ( .A(n9986), .B(n9985), .Z(n9990) );
  NAND U11097 ( .A(n9988), .B(n9987), .Z(n9989) );
  NAND U11098 ( .A(n9990), .B(n9989), .Z(n10187) );
  NANDN U11099 ( .A(n9992), .B(n9991), .Z(n9996) );
  NAND U11100 ( .A(n9994), .B(n9993), .Z(n9995) );
  NAND U11101 ( .A(n9996), .B(n9995), .Z(n10126) );
  NANDN U11102 ( .A(n9998), .B(n9997), .Z(n10002) );
  NAND U11103 ( .A(n10000), .B(n9999), .Z(n10001) );
  AND U11104 ( .A(n10002), .B(n10001), .Z(n10127) );
  XNOR U11105 ( .A(n10126), .B(n10127), .Z(n10128) );
  XOR U11106 ( .A(n1052), .B(a[69]), .Z(n10156) );
  NANDN U11107 ( .A(n10156), .B(n36925), .Z(n10005) );
  NAND U11108 ( .A(n36926), .B(n10003), .Z(n10004) );
  NAND U11109 ( .A(n10005), .B(n10004), .Z(n10112) );
  XNOR U11110 ( .A(n1054), .B(a[63]), .Z(n10153) );
  NANDN U11111 ( .A(n37665), .B(n10153), .Z(n10008) );
  NANDN U11112 ( .A(n10006), .B(n37604), .Z(n10007) );
  NAND U11113 ( .A(n10008), .B(n10007), .Z(n10110) );
  XOR U11114 ( .A(n1056), .B(a[57]), .Z(n10150) );
  NANDN U11115 ( .A(n10150), .B(n38101), .Z(n10011) );
  NAND U11116 ( .A(n38102), .B(n10009), .Z(n10010) );
  NAND U11117 ( .A(n10011), .B(n10010), .Z(n10111) );
  XNOR U11118 ( .A(n10110), .B(n10111), .Z(n10113) );
  XOR U11119 ( .A(n10112), .B(n10113), .Z(n10101) );
  XOR U11120 ( .A(b[11]), .B(n13219), .Z(n10159) );
  OR U11121 ( .A(n10159), .B(n37311), .Z(n10014) );
  NANDN U11122 ( .A(n10012), .B(n37218), .Z(n10013) );
  NAND U11123 ( .A(n10014), .B(n10013), .Z(n10099) );
  XOR U11124 ( .A(n1053), .B(a[65]), .Z(n10162) );
  NANDN U11125 ( .A(n10162), .B(n37424), .Z(n10017) );
  NANDN U11126 ( .A(n10015), .B(n37425), .Z(n10016) );
  AND U11127 ( .A(n10017), .B(n10016), .Z(n10098) );
  XNOR U11128 ( .A(n10099), .B(n10098), .Z(n10100) );
  XNOR U11129 ( .A(n10101), .B(n10100), .Z(n10117) );
  NANDN U11130 ( .A(n1049), .B(a[77]), .Z(n10018) );
  XNOR U11131 ( .A(b[1]), .B(n10018), .Z(n10020) );
  NANDN U11132 ( .A(b[0]), .B(a[76]), .Z(n10019) );
  AND U11133 ( .A(n10020), .B(n10019), .Z(n10076) );
  NAND U11134 ( .A(n10021), .B(n38490), .Z(n10023) );
  XNOR U11135 ( .A(n1058), .B(a[49]), .Z(n10165) );
  NANDN U11136 ( .A(n1048), .B(n10165), .Z(n10022) );
  NAND U11137 ( .A(n10023), .B(n10022), .Z(n10074) );
  NANDN U11138 ( .A(n1059), .B(a[45]), .Z(n10075) );
  XNOR U11139 ( .A(n10074), .B(n10075), .Z(n10077) );
  XNOR U11140 ( .A(n10076), .B(n10077), .Z(n10115) );
  NANDN U11141 ( .A(n10024), .B(n38205), .Z(n10026) );
  XNOR U11142 ( .A(b[23]), .B(a[55]), .Z(n10171) );
  OR U11143 ( .A(n10171), .B(n38268), .Z(n10025) );
  NAND U11144 ( .A(n10026), .B(n10025), .Z(n10141) );
  XOR U11145 ( .A(b[7]), .B(a[71]), .Z(n10174) );
  NAND U11146 ( .A(n10174), .B(n36701), .Z(n10029) );
  NAND U11147 ( .A(n10027), .B(n36702), .Z(n10028) );
  NAND U11148 ( .A(n10029), .B(n10028), .Z(n10138) );
  XOR U11149 ( .A(b[25]), .B(a[53]), .Z(n10177) );
  NAND U11150 ( .A(n10177), .B(n38325), .Z(n10032) );
  NAND U11151 ( .A(n10030), .B(n38326), .Z(n10031) );
  AND U11152 ( .A(n10032), .B(n10031), .Z(n10139) );
  XNOR U11153 ( .A(n10138), .B(n10139), .Z(n10140) );
  XOR U11154 ( .A(n10141), .B(n10140), .Z(n10114) );
  XOR U11155 ( .A(n10117), .B(n10116), .Z(n10129) );
  XOR U11156 ( .A(n10128), .B(n10129), .Z(n10186) );
  XNOR U11157 ( .A(n10187), .B(n10186), .Z(n10189) );
  XNOR U11158 ( .A(n10188), .B(n10189), .Z(n10068) );
  XNOR U11159 ( .A(n10069), .B(n10068), .Z(n10070) );
  XOR U11160 ( .A(n10071), .B(n10070), .Z(n10065) );
  NANDN U11161 ( .A(n10034), .B(n10033), .Z(n10038) );
  OR U11162 ( .A(n10036), .B(n10035), .Z(n10037) );
  NAND U11163 ( .A(n10038), .B(n10037), .Z(n10062) );
  NAND U11164 ( .A(n10040), .B(n10039), .Z(n10044) );
  NANDN U11165 ( .A(n10042), .B(n10041), .Z(n10043) );
  NAND U11166 ( .A(n10044), .B(n10043), .Z(n10063) );
  XNOR U11167 ( .A(n10062), .B(n10063), .Z(n10064) );
  XOR U11168 ( .A(n10065), .B(n10064), .Z(n10059) );
  XOR U11169 ( .A(n10058), .B(n10059), .Z(n10050) );
  XOR U11170 ( .A(n10051), .B(n10050), .Z(n10052) );
  XNOR U11171 ( .A(n10053), .B(n10052), .Z(n10192) );
  XNOR U11172 ( .A(n10192), .B(sreg[301]), .Z(n10194) );
  NAND U11173 ( .A(n10045), .B(sreg[300]), .Z(n10049) );
  OR U11174 ( .A(n10047), .B(n10046), .Z(n10048) );
  AND U11175 ( .A(n10049), .B(n10048), .Z(n10193) );
  XOR U11176 ( .A(n10194), .B(n10193), .Z(c[301]) );
  NAND U11177 ( .A(n10051), .B(n10050), .Z(n10055) );
  NAND U11178 ( .A(n10053), .B(n10052), .Z(n10054) );
  NAND U11179 ( .A(n10055), .B(n10054), .Z(n10200) );
  NANDN U11180 ( .A(n10057), .B(n10056), .Z(n10061) );
  NAND U11181 ( .A(n10059), .B(n10058), .Z(n10060) );
  NAND U11182 ( .A(n10061), .B(n10060), .Z(n10198) );
  NANDN U11183 ( .A(n10063), .B(n10062), .Z(n10067) );
  NAND U11184 ( .A(n10065), .B(n10064), .Z(n10066) );
  NAND U11185 ( .A(n10067), .B(n10066), .Z(n10203) );
  NANDN U11186 ( .A(n10069), .B(n10068), .Z(n10073) );
  NANDN U11187 ( .A(n10071), .B(n10070), .Z(n10072) );
  NAND U11188 ( .A(n10073), .B(n10072), .Z(n10204) );
  XNOR U11189 ( .A(n10203), .B(n10204), .Z(n10205) );
  NANDN U11190 ( .A(n10075), .B(n10074), .Z(n10079) );
  NAND U11191 ( .A(n10077), .B(n10076), .Z(n10078) );
  NAND U11192 ( .A(n10079), .B(n10078), .Z(n10278) );
  XNOR U11193 ( .A(b[19]), .B(a[60]), .Z(n10225) );
  NANDN U11194 ( .A(n10225), .B(n37934), .Z(n10082) );
  NANDN U11195 ( .A(n10080), .B(n37935), .Z(n10081) );
  NAND U11196 ( .A(n10082), .B(n10081), .Z(n10288) );
  XOR U11197 ( .A(b[27]), .B(a[52]), .Z(n10228) );
  NAND U11198 ( .A(n38423), .B(n10228), .Z(n10085) );
  NAND U11199 ( .A(n10083), .B(n38424), .Z(n10084) );
  NAND U11200 ( .A(n10085), .B(n10084), .Z(n10285) );
  XNOR U11201 ( .A(b[5]), .B(a[74]), .Z(n10231) );
  NANDN U11202 ( .A(n10231), .B(n36587), .Z(n10088) );
  NANDN U11203 ( .A(n10086), .B(n36588), .Z(n10087) );
  AND U11204 ( .A(n10088), .B(n10087), .Z(n10286) );
  XNOR U11205 ( .A(n10285), .B(n10286), .Z(n10287) );
  XNOR U11206 ( .A(n10288), .B(n10287), .Z(n10276) );
  NAND U11207 ( .A(n10089), .B(n37762), .Z(n10091) );
  XNOR U11208 ( .A(b[17]), .B(a[62]), .Z(n10234) );
  NANDN U11209 ( .A(n10234), .B(n37764), .Z(n10090) );
  NAND U11210 ( .A(n10091), .B(n10090), .Z(n10252) );
  XNOR U11211 ( .A(b[31]), .B(a[48]), .Z(n10237) );
  NANDN U11212 ( .A(n10237), .B(n38552), .Z(n10094) );
  NANDN U11213 ( .A(n10092), .B(n38553), .Z(n10093) );
  NAND U11214 ( .A(n10094), .B(n10093), .Z(n10249) );
  OR U11215 ( .A(n10095), .B(n36105), .Z(n10097) );
  XNOR U11216 ( .A(b[3]), .B(a[76]), .Z(n10240) );
  NANDN U11217 ( .A(n10240), .B(n36107), .Z(n10096) );
  AND U11218 ( .A(n10097), .B(n10096), .Z(n10250) );
  XNOR U11219 ( .A(n10249), .B(n10250), .Z(n10251) );
  XOR U11220 ( .A(n10252), .B(n10251), .Z(n10275) );
  XNOR U11221 ( .A(n10276), .B(n10275), .Z(n10277) );
  XNOR U11222 ( .A(n10278), .B(n10277), .Z(n10216) );
  NANDN U11223 ( .A(n10099), .B(n10098), .Z(n10103) );
  NAND U11224 ( .A(n10101), .B(n10100), .Z(n10102) );
  NAND U11225 ( .A(n10103), .B(n10102), .Z(n10267) );
  NANDN U11226 ( .A(n10105), .B(n10104), .Z(n10109) );
  NAND U11227 ( .A(n10107), .B(n10106), .Z(n10108) );
  NAND U11228 ( .A(n10109), .B(n10108), .Z(n10266) );
  XNOR U11229 ( .A(n10266), .B(n10265), .Z(n10268) );
  XOR U11230 ( .A(n10267), .B(n10268), .Z(n10215) );
  XOR U11231 ( .A(n10216), .B(n10215), .Z(n10217) );
  NANDN U11232 ( .A(n10115), .B(n10114), .Z(n10119) );
  NAND U11233 ( .A(n10117), .B(n10116), .Z(n10118) );
  NAND U11234 ( .A(n10119), .B(n10118), .Z(n10218) );
  XNOR U11235 ( .A(n10217), .B(n10218), .Z(n10329) );
  OR U11236 ( .A(n10121), .B(n10120), .Z(n10125) );
  NANDN U11237 ( .A(n10123), .B(n10122), .Z(n10124) );
  NAND U11238 ( .A(n10125), .B(n10124), .Z(n10328) );
  NANDN U11239 ( .A(n10127), .B(n10126), .Z(n10131) );
  NAND U11240 ( .A(n10129), .B(n10128), .Z(n10130) );
  NAND U11241 ( .A(n10131), .B(n10130), .Z(n10211) );
  NANDN U11242 ( .A(n10133), .B(n10132), .Z(n10137) );
  OR U11243 ( .A(n10135), .B(n10134), .Z(n10136) );
  NAND U11244 ( .A(n10137), .B(n10136), .Z(n10210) );
  NANDN U11245 ( .A(n10139), .B(n10138), .Z(n10143) );
  NAND U11246 ( .A(n10141), .B(n10140), .Z(n10142) );
  NAND U11247 ( .A(n10143), .B(n10142), .Z(n10269) );
  NANDN U11248 ( .A(n10145), .B(n10144), .Z(n10149) );
  NAND U11249 ( .A(n10147), .B(n10146), .Z(n10148) );
  AND U11250 ( .A(n10149), .B(n10148), .Z(n10270) );
  XNOR U11251 ( .A(n10269), .B(n10270), .Z(n10271) );
  XNOR U11252 ( .A(b[21]), .B(a[58]), .Z(n10297) );
  NANDN U11253 ( .A(n10297), .B(n38101), .Z(n10152) );
  NANDN U11254 ( .A(n10150), .B(n38102), .Z(n10151) );
  NAND U11255 ( .A(n10152), .B(n10151), .Z(n10261) );
  XNOR U11256 ( .A(b[15]), .B(a[64]), .Z(n10294) );
  OR U11257 ( .A(n10294), .B(n37665), .Z(n10155) );
  NAND U11258 ( .A(n10153), .B(n37604), .Z(n10154) );
  AND U11259 ( .A(n10155), .B(n10154), .Z(n10262) );
  XNOR U11260 ( .A(n10261), .B(n10262), .Z(n10264) );
  XNOR U11261 ( .A(b[9]), .B(a[70]), .Z(n10291) );
  NANDN U11262 ( .A(n10291), .B(n36925), .Z(n10158) );
  NANDN U11263 ( .A(n10156), .B(n36926), .Z(n10157) );
  NAND U11264 ( .A(n10158), .B(n10157), .Z(n10263) );
  XNOR U11265 ( .A(n10264), .B(n10263), .Z(n10257) );
  XNOR U11266 ( .A(b[11]), .B(a[68]), .Z(n10300) );
  OR U11267 ( .A(n10300), .B(n37311), .Z(n10161) );
  NANDN U11268 ( .A(n10159), .B(n37218), .Z(n10160) );
  NAND U11269 ( .A(n10161), .B(n10160), .Z(n10256) );
  XOR U11270 ( .A(n1053), .B(a[66]), .Z(n10303) );
  NANDN U11271 ( .A(n10303), .B(n37424), .Z(n10164) );
  NANDN U11272 ( .A(n10162), .B(n37425), .Z(n10163) );
  NAND U11273 ( .A(n10164), .B(n10163), .Z(n10255) );
  XNOR U11274 ( .A(n10256), .B(n10255), .Z(n10258) );
  XNOR U11275 ( .A(n10257), .B(n10258), .Z(n10246) );
  NAND U11276 ( .A(n38490), .B(n10165), .Z(n10167) );
  XOR U11277 ( .A(n1058), .B(n10724), .Z(n10309) );
  NANDN U11278 ( .A(n1048), .B(n10309), .Z(n10166) );
  NAND U11279 ( .A(n10167), .B(n10166), .Z(n10219) );
  NANDN U11280 ( .A(n1059), .B(a[46]), .Z(n10220) );
  XNOR U11281 ( .A(n10219), .B(n10220), .Z(n10222) );
  NANDN U11282 ( .A(n1049), .B(a[78]), .Z(n10168) );
  XNOR U11283 ( .A(b[1]), .B(n10168), .Z(n10170) );
  NANDN U11284 ( .A(b[0]), .B(a[77]), .Z(n10169) );
  AND U11285 ( .A(n10170), .B(n10169), .Z(n10221) );
  XNOR U11286 ( .A(n10222), .B(n10221), .Z(n10244) );
  NANDN U11287 ( .A(n10171), .B(n38205), .Z(n10173) );
  XNOR U11288 ( .A(b[23]), .B(a[56]), .Z(n10312) );
  OR U11289 ( .A(n10312), .B(n38268), .Z(n10172) );
  NAND U11290 ( .A(n10173), .B(n10172), .Z(n10282) );
  XOR U11291 ( .A(b[7]), .B(a[72]), .Z(n10315) );
  NAND U11292 ( .A(n10315), .B(n36701), .Z(n10176) );
  NAND U11293 ( .A(n10174), .B(n36702), .Z(n10175) );
  NAND U11294 ( .A(n10176), .B(n10175), .Z(n10279) );
  XNOR U11295 ( .A(b[25]), .B(a[54]), .Z(n10318) );
  NANDN U11296 ( .A(n10318), .B(n38325), .Z(n10179) );
  NAND U11297 ( .A(n10177), .B(n38326), .Z(n10178) );
  AND U11298 ( .A(n10179), .B(n10178), .Z(n10280) );
  XNOR U11299 ( .A(n10279), .B(n10280), .Z(n10281) );
  XOR U11300 ( .A(n10282), .B(n10281), .Z(n10243) );
  XOR U11301 ( .A(n10246), .B(n10245), .Z(n10272) );
  XNOR U11302 ( .A(n10271), .B(n10272), .Z(n10209) );
  XNOR U11303 ( .A(n10210), .B(n10209), .Z(n10212) );
  XNOR U11304 ( .A(n10211), .B(n10212), .Z(n10327) );
  XOR U11305 ( .A(n10328), .B(n10327), .Z(n10330) );
  NAND U11306 ( .A(n10181), .B(n10180), .Z(n10185) );
  NAND U11307 ( .A(n10183), .B(n10182), .Z(n10184) );
  NAND U11308 ( .A(n10185), .B(n10184), .Z(n10322) );
  NAND U11309 ( .A(n10187), .B(n10186), .Z(n10191) );
  NANDN U11310 ( .A(n10189), .B(n10188), .Z(n10190) );
  AND U11311 ( .A(n10191), .B(n10190), .Z(n10321) );
  XNOR U11312 ( .A(n10322), .B(n10321), .Z(n10323) );
  XOR U11313 ( .A(n10324), .B(n10323), .Z(n10206) );
  XOR U11314 ( .A(n10205), .B(n10206), .Z(n10197) );
  XOR U11315 ( .A(n10198), .B(n10197), .Z(n10199) );
  XNOR U11316 ( .A(n10200), .B(n10199), .Z(n10333) );
  XNOR U11317 ( .A(n10333), .B(sreg[302]), .Z(n10335) );
  NAND U11318 ( .A(n10192), .B(sreg[301]), .Z(n10196) );
  OR U11319 ( .A(n10194), .B(n10193), .Z(n10195) );
  AND U11320 ( .A(n10196), .B(n10195), .Z(n10334) );
  XOR U11321 ( .A(n10335), .B(n10334), .Z(c[302]) );
  NAND U11322 ( .A(n10198), .B(n10197), .Z(n10202) );
  NAND U11323 ( .A(n10200), .B(n10199), .Z(n10201) );
  NAND U11324 ( .A(n10202), .B(n10201), .Z(n10341) );
  NANDN U11325 ( .A(n10204), .B(n10203), .Z(n10208) );
  NAND U11326 ( .A(n10206), .B(n10205), .Z(n10207) );
  NAND U11327 ( .A(n10208), .B(n10207), .Z(n10338) );
  NAND U11328 ( .A(n10210), .B(n10209), .Z(n10214) );
  NANDN U11329 ( .A(n10212), .B(n10211), .Z(n10213) );
  NAND U11330 ( .A(n10214), .B(n10213), .Z(n10466) );
  XNOR U11331 ( .A(n10466), .B(n10467), .Z(n10468) );
  NANDN U11332 ( .A(n10220), .B(n10219), .Z(n10224) );
  NAND U11333 ( .A(n10222), .B(n10221), .Z(n10223) );
  NAND U11334 ( .A(n10224), .B(n10223), .Z(n10411) );
  XNOR U11335 ( .A(b[19]), .B(a[61]), .Z(n10356) );
  NANDN U11336 ( .A(n10356), .B(n37934), .Z(n10227) );
  NANDN U11337 ( .A(n10225), .B(n37935), .Z(n10226) );
  NAND U11338 ( .A(n10227), .B(n10226), .Z(n10421) );
  XOR U11339 ( .A(b[27]), .B(a[53]), .Z(n10359) );
  NAND U11340 ( .A(n38423), .B(n10359), .Z(n10230) );
  NAND U11341 ( .A(n10228), .B(n38424), .Z(n10229) );
  NAND U11342 ( .A(n10230), .B(n10229), .Z(n10418) );
  XNOR U11343 ( .A(b[5]), .B(a[75]), .Z(n10362) );
  NANDN U11344 ( .A(n10362), .B(n36587), .Z(n10233) );
  NANDN U11345 ( .A(n10231), .B(n36588), .Z(n10232) );
  AND U11346 ( .A(n10233), .B(n10232), .Z(n10419) );
  XNOR U11347 ( .A(n10418), .B(n10419), .Z(n10420) );
  XNOR U11348 ( .A(n10421), .B(n10420), .Z(n10409) );
  NANDN U11349 ( .A(n10234), .B(n37762), .Z(n10236) );
  XOR U11350 ( .A(b[17]), .B(a[63]), .Z(n10365) );
  NAND U11351 ( .A(n10365), .B(n37764), .Z(n10235) );
  NAND U11352 ( .A(n10236), .B(n10235), .Z(n10383) );
  XNOR U11353 ( .A(b[31]), .B(a[49]), .Z(n10368) );
  NANDN U11354 ( .A(n10368), .B(n38552), .Z(n10239) );
  NANDN U11355 ( .A(n10237), .B(n38553), .Z(n10238) );
  NAND U11356 ( .A(n10239), .B(n10238), .Z(n10380) );
  OR U11357 ( .A(n10240), .B(n36105), .Z(n10242) );
  XNOR U11358 ( .A(b[3]), .B(a[77]), .Z(n10371) );
  NANDN U11359 ( .A(n10371), .B(n36107), .Z(n10241) );
  AND U11360 ( .A(n10242), .B(n10241), .Z(n10381) );
  XNOR U11361 ( .A(n10380), .B(n10381), .Z(n10382) );
  XOR U11362 ( .A(n10383), .B(n10382), .Z(n10408) );
  XNOR U11363 ( .A(n10409), .B(n10408), .Z(n10410) );
  XNOR U11364 ( .A(n10411), .B(n10410), .Z(n10460) );
  NANDN U11365 ( .A(n10244), .B(n10243), .Z(n10248) );
  NANDN U11366 ( .A(n10246), .B(n10245), .Z(n10247) );
  NAND U11367 ( .A(n10248), .B(n10247), .Z(n10461) );
  XNOR U11368 ( .A(n10460), .B(n10461), .Z(n10462) );
  NANDN U11369 ( .A(n10250), .B(n10249), .Z(n10254) );
  NAND U11370 ( .A(n10252), .B(n10251), .Z(n10253) );
  NAND U11371 ( .A(n10254), .B(n10253), .Z(n10401) );
  OR U11372 ( .A(n10256), .B(n10255), .Z(n10260) );
  NANDN U11373 ( .A(n10258), .B(n10257), .Z(n10259) );
  NAND U11374 ( .A(n10260), .B(n10259), .Z(n10399) );
  XNOR U11375 ( .A(n10399), .B(n10398), .Z(n10400) );
  XOR U11376 ( .A(n10401), .B(n10400), .Z(n10463) );
  XOR U11377 ( .A(n10462), .B(n10463), .Z(n10474) );
  NANDN U11378 ( .A(n10270), .B(n10269), .Z(n10274) );
  NANDN U11379 ( .A(n10272), .B(n10271), .Z(n10273) );
  NAND U11380 ( .A(n10274), .B(n10273), .Z(n10457) );
  NANDN U11381 ( .A(n10280), .B(n10279), .Z(n10284) );
  NAND U11382 ( .A(n10282), .B(n10281), .Z(n10283) );
  NAND U11383 ( .A(n10284), .B(n10283), .Z(n10402) );
  NANDN U11384 ( .A(n10286), .B(n10285), .Z(n10290) );
  NAND U11385 ( .A(n10288), .B(n10287), .Z(n10289) );
  AND U11386 ( .A(n10290), .B(n10289), .Z(n10403) );
  XNOR U11387 ( .A(n10402), .B(n10403), .Z(n10404) );
  XNOR U11388 ( .A(b[9]), .B(a[71]), .Z(n10424) );
  NANDN U11389 ( .A(n10424), .B(n36925), .Z(n10293) );
  NANDN U11390 ( .A(n10291), .B(n36926), .Z(n10292) );
  NAND U11391 ( .A(n10293), .B(n10292), .Z(n10388) );
  XNOR U11392 ( .A(b[15]), .B(a[65]), .Z(n10427) );
  OR U11393 ( .A(n10427), .B(n37665), .Z(n10296) );
  NANDN U11394 ( .A(n10294), .B(n37604), .Z(n10295) );
  AND U11395 ( .A(n10296), .B(n10295), .Z(n10386) );
  XOR U11396 ( .A(b[21]), .B(n12056), .Z(n10430) );
  NANDN U11397 ( .A(n10430), .B(n38101), .Z(n10299) );
  NANDN U11398 ( .A(n10297), .B(n38102), .Z(n10298) );
  AND U11399 ( .A(n10299), .B(n10298), .Z(n10387) );
  XOR U11400 ( .A(n10388), .B(n10389), .Z(n10377) );
  XNOR U11401 ( .A(b[11]), .B(a[69]), .Z(n10433) );
  OR U11402 ( .A(n10433), .B(n37311), .Z(n10302) );
  NANDN U11403 ( .A(n10300), .B(n37218), .Z(n10301) );
  NAND U11404 ( .A(n10302), .B(n10301), .Z(n10375) );
  XOR U11405 ( .A(n1053), .B(a[67]), .Z(n10436) );
  NANDN U11406 ( .A(n10436), .B(n37424), .Z(n10305) );
  NANDN U11407 ( .A(n10303), .B(n37425), .Z(n10304) );
  AND U11408 ( .A(n10305), .B(n10304), .Z(n10374) );
  XNOR U11409 ( .A(n10375), .B(n10374), .Z(n10376) );
  XOR U11410 ( .A(n10377), .B(n10376), .Z(n10394) );
  NANDN U11411 ( .A(n1049), .B(a[79]), .Z(n10306) );
  XNOR U11412 ( .A(b[1]), .B(n10306), .Z(n10308) );
  NANDN U11413 ( .A(b[0]), .B(a[78]), .Z(n10307) );
  AND U11414 ( .A(n10308), .B(n10307), .Z(n10352) );
  NAND U11415 ( .A(n38490), .B(n10309), .Z(n10311) );
  XNOR U11416 ( .A(n1058), .B(a[51]), .Z(n10439) );
  NANDN U11417 ( .A(n1048), .B(n10439), .Z(n10310) );
  NAND U11418 ( .A(n10311), .B(n10310), .Z(n10350) );
  NANDN U11419 ( .A(n1059), .B(a[47]), .Z(n10351) );
  XNOR U11420 ( .A(n10350), .B(n10351), .Z(n10353) );
  XOR U11421 ( .A(n10352), .B(n10353), .Z(n10392) );
  NANDN U11422 ( .A(n10312), .B(n38205), .Z(n10314) );
  XNOR U11423 ( .A(b[23]), .B(a[57]), .Z(n10445) );
  OR U11424 ( .A(n10445), .B(n38268), .Z(n10313) );
  NAND U11425 ( .A(n10314), .B(n10313), .Z(n10415) );
  XOR U11426 ( .A(b[7]), .B(a[73]), .Z(n10448) );
  NAND U11427 ( .A(n10448), .B(n36701), .Z(n10317) );
  NAND U11428 ( .A(n10315), .B(n36702), .Z(n10316) );
  NAND U11429 ( .A(n10317), .B(n10316), .Z(n10412) );
  XOR U11430 ( .A(b[25]), .B(a[55]), .Z(n10451) );
  NAND U11431 ( .A(n10451), .B(n38325), .Z(n10320) );
  NANDN U11432 ( .A(n10318), .B(n38326), .Z(n10319) );
  AND U11433 ( .A(n10320), .B(n10319), .Z(n10413) );
  XNOR U11434 ( .A(n10412), .B(n10413), .Z(n10414) );
  XNOR U11435 ( .A(n10415), .B(n10414), .Z(n10393) );
  XOR U11436 ( .A(n10392), .B(n10393), .Z(n10395) );
  XNOR U11437 ( .A(n10394), .B(n10395), .Z(n10405) );
  XOR U11438 ( .A(n10404), .B(n10405), .Z(n10455) );
  XNOR U11439 ( .A(n10454), .B(n10455), .Z(n10456) );
  XNOR U11440 ( .A(n10457), .B(n10456), .Z(n10472) );
  XNOR U11441 ( .A(n10473), .B(n10472), .Z(n10475) );
  XNOR U11442 ( .A(n10474), .B(n10475), .Z(n10469) );
  XOR U11443 ( .A(n10468), .B(n10469), .Z(n10347) );
  NANDN U11444 ( .A(n10322), .B(n10321), .Z(n10326) );
  NAND U11445 ( .A(n10324), .B(n10323), .Z(n10325) );
  NAND U11446 ( .A(n10326), .B(n10325), .Z(n10344) );
  NANDN U11447 ( .A(n10328), .B(n10327), .Z(n10332) );
  OR U11448 ( .A(n10330), .B(n10329), .Z(n10331) );
  NAND U11449 ( .A(n10332), .B(n10331), .Z(n10345) );
  XNOR U11450 ( .A(n10344), .B(n10345), .Z(n10346) );
  XNOR U11451 ( .A(n10347), .B(n10346), .Z(n10339) );
  XNOR U11452 ( .A(n10338), .B(n10339), .Z(n10340) );
  XNOR U11453 ( .A(n10341), .B(n10340), .Z(n10478) );
  XNOR U11454 ( .A(n10478), .B(sreg[303]), .Z(n10480) );
  NAND U11455 ( .A(n10333), .B(sreg[302]), .Z(n10337) );
  OR U11456 ( .A(n10335), .B(n10334), .Z(n10336) );
  AND U11457 ( .A(n10337), .B(n10336), .Z(n10479) );
  XOR U11458 ( .A(n10480), .B(n10479), .Z(c[303]) );
  NANDN U11459 ( .A(n10339), .B(n10338), .Z(n10343) );
  NAND U11460 ( .A(n10341), .B(n10340), .Z(n10342) );
  NAND U11461 ( .A(n10343), .B(n10342), .Z(n10486) );
  NANDN U11462 ( .A(n10345), .B(n10344), .Z(n10349) );
  NAND U11463 ( .A(n10347), .B(n10346), .Z(n10348) );
  NAND U11464 ( .A(n10349), .B(n10348), .Z(n10484) );
  NANDN U11465 ( .A(n10351), .B(n10350), .Z(n10355) );
  NAND U11466 ( .A(n10353), .B(n10352), .Z(n10354) );
  NAND U11467 ( .A(n10355), .B(n10354), .Z(n10556) );
  XOR U11468 ( .A(b[19]), .B(n12493), .Z(n10499) );
  NANDN U11469 ( .A(n10499), .B(n37934), .Z(n10358) );
  NANDN U11470 ( .A(n10356), .B(n37935), .Z(n10357) );
  NAND U11471 ( .A(n10358), .B(n10357), .Z(n10566) );
  XNOR U11472 ( .A(b[27]), .B(a[54]), .Z(n10502) );
  NANDN U11473 ( .A(n10502), .B(n38423), .Z(n10361) );
  NAND U11474 ( .A(n10359), .B(n38424), .Z(n10360) );
  NAND U11475 ( .A(n10361), .B(n10360), .Z(n10563) );
  XNOR U11476 ( .A(b[5]), .B(a[76]), .Z(n10505) );
  NANDN U11477 ( .A(n10505), .B(n36587), .Z(n10364) );
  NANDN U11478 ( .A(n10362), .B(n36588), .Z(n10363) );
  AND U11479 ( .A(n10364), .B(n10363), .Z(n10564) );
  XNOR U11480 ( .A(n10563), .B(n10564), .Z(n10565) );
  XNOR U11481 ( .A(n10566), .B(n10565), .Z(n10554) );
  NAND U11482 ( .A(n10365), .B(n37762), .Z(n10367) );
  XOR U11483 ( .A(b[17]), .B(a[64]), .Z(n10508) );
  NAND U11484 ( .A(n10508), .B(n37764), .Z(n10366) );
  NAND U11485 ( .A(n10367), .B(n10366), .Z(n10526) );
  XOR U11486 ( .A(b[31]), .B(n10724), .Z(n10511) );
  NANDN U11487 ( .A(n10511), .B(n38552), .Z(n10370) );
  NANDN U11488 ( .A(n10368), .B(n38553), .Z(n10369) );
  NAND U11489 ( .A(n10370), .B(n10369), .Z(n10523) );
  OR U11490 ( .A(n10371), .B(n36105), .Z(n10373) );
  XNOR U11491 ( .A(b[3]), .B(a[78]), .Z(n10514) );
  NANDN U11492 ( .A(n10514), .B(n36107), .Z(n10372) );
  AND U11493 ( .A(n10373), .B(n10372), .Z(n10524) );
  XNOR U11494 ( .A(n10523), .B(n10524), .Z(n10525) );
  XOR U11495 ( .A(n10526), .B(n10525), .Z(n10553) );
  XNOR U11496 ( .A(n10554), .B(n10553), .Z(n10555) );
  XNOR U11497 ( .A(n10556), .B(n10555), .Z(n10599) );
  NANDN U11498 ( .A(n10375), .B(n10374), .Z(n10379) );
  NAND U11499 ( .A(n10377), .B(n10376), .Z(n10378) );
  NAND U11500 ( .A(n10379), .B(n10378), .Z(n10544) );
  NANDN U11501 ( .A(n10381), .B(n10380), .Z(n10385) );
  NAND U11502 ( .A(n10383), .B(n10382), .Z(n10384) );
  NAND U11503 ( .A(n10385), .B(n10384), .Z(n10542) );
  OR U11504 ( .A(n10387), .B(n10386), .Z(n10391) );
  NANDN U11505 ( .A(n10389), .B(n10388), .Z(n10390) );
  NAND U11506 ( .A(n10391), .B(n10390), .Z(n10541) );
  XNOR U11507 ( .A(n10544), .B(n10543), .Z(n10600) );
  XNOR U11508 ( .A(n10599), .B(n10600), .Z(n10601) );
  NANDN U11509 ( .A(n10393), .B(n10392), .Z(n10397) );
  OR U11510 ( .A(n10395), .B(n10394), .Z(n10396) );
  AND U11511 ( .A(n10397), .B(n10396), .Z(n10602) );
  XNOR U11512 ( .A(n10601), .B(n10602), .Z(n10614) );
  NANDN U11513 ( .A(n10403), .B(n10402), .Z(n10407) );
  NANDN U11514 ( .A(n10405), .B(n10404), .Z(n10406) );
  NAND U11515 ( .A(n10407), .B(n10406), .Z(n10608) );
  NANDN U11516 ( .A(n10413), .B(n10412), .Z(n10417) );
  NAND U11517 ( .A(n10415), .B(n10414), .Z(n10416) );
  NAND U11518 ( .A(n10417), .B(n10416), .Z(n10547) );
  NANDN U11519 ( .A(n10419), .B(n10418), .Z(n10423) );
  NAND U11520 ( .A(n10421), .B(n10420), .Z(n10422) );
  AND U11521 ( .A(n10423), .B(n10422), .Z(n10548) );
  XNOR U11522 ( .A(n10547), .B(n10548), .Z(n10549) );
  XNOR U11523 ( .A(n1052), .B(a[72]), .Z(n10569) );
  NAND U11524 ( .A(n36925), .B(n10569), .Z(n10426) );
  NANDN U11525 ( .A(n10424), .B(n36926), .Z(n10425) );
  NAND U11526 ( .A(n10426), .B(n10425), .Z(n10537) );
  XNOR U11527 ( .A(b[15]), .B(a[66]), .Z(n10572) );
  OR U11528 ( .A(n10572), .B(n37665), .Z(n10429) );
  NANDN U11529 ( .A(n10427), .B(n37604), .Z(n10428) );
  AND U11530 ( .A(n10429), .B(n10428), .Z(n10535) );
  XNOR U11531 ( .A(n1056), .B(a[60]), .Z(n10575) );
  NAND U11532 ( .A(n10575), .B(n38101), .Z(n10432) );
  NANDN U11533 ( .A(n10430), .B(n38102), .Z(n10431) );
  AND U11534 ( .A(n10432), .B(n10431), .Z(n10536) );
  XOR U11535 ( .A(n10537), .B(n10538), .Z(n10532) );
  XNOR U11536 ( .A(b[11]), .B(a[70]), .Z(n10578) );
  OR U11537 ( .A(n10578), .B(n37311), .Z(n10435) );
  NANDN U11538 ( .A(n10433), .B(n37218), .Z(n10434) );
  NAND U11539 ( .A(n10435), .B(n10434), .Z(n10530) );
  XOR U11540 ( .A(n1053), .B(a[68]), .Z(n10581) );
  NANDN U11541 ( .A(n10581), .B(n37424), .Z(n10438) );
  NANDN U11542 ( .A(n10436), .B(n37425), .Z(n10437) );
  NAND U11543 ( .A(n10438), .B(n10437), .Z(n10529) );
  XOR U11544 ( .A(n10532), .B(n10531), .Z(n10519) );
  NAND U11545 ( .A(n38490), .B(n10439), .Z(n10441) );
  XNOR U11546 ( .A(n1058), .B(a[52]), .Z(n10587) );
  NANDN U11547 ( .A(n1048), .B(n10587), .Z(n10440) );
  NAND U11548 ( .A(n10441), .B(n10440), .Z(n10493) );
  NANDN U11549 ( .A(n1059), .B(a[48]), .Z(n10494) );
  XNOR U11550 ( .A(n10493), .B(n10494), .Z(n10496) );
  NANDN U11551 ( .A(n1049), .B(a[80]), .Z(n10442) );
  XNOR U11552 ( .A(b[1]), .B(n10442), .Z(n10444) );
  NANDN U11553 ( .A(b[0]), .B(a[79]), .Z(n10443) );
  AND U11554 ( .A(n10444), .B(n10443), .Z(n10495) );
  XOR U11555 ( .A(n10496), .B(n10495), .Z(n10517) );
  NANDN U11556 ( .A(n10445), .B(n38205), .Z(n10447) );
  XNOR U11557 ( .A(b[23]), .B(a[58]), .Z(n10590) );
  OR U11558 ( .A(n10590), .B(n38268), .Z(n10446) );
  NAND U11559 ( .A(n10447), .B(n10446), .Z(n10560) );
  XOR U11560 ( .A(b[7]), .B(a[74]), .Z(n10593) );
  NAND U11561 ( .A(n10593), .B(n36701), .Z(n10450) );
  NAND U11562 ( .A(n10448), .B(n36702), .Z(n10449) );
  NAND U11563 ( .A(n10450), .B(n10449), .Z(n10557) );
  XOR U11564 ( .A(b[25]), .B(a[56]), .Z(n10596) );
  NAND U11565 ( .A(n10596), .B(n38325), .Z(n10453) );
  NAND U11566 ( .A(n10451), .B(n38326), .Z(n10452) );
  AND U11567 ( .A(n10453), .B(n10452), .Z(n10558) );
  XNOR U11568 ( .A(n10557), .B(n10558), .Z(n10559) );
  XNOR U11569 ( .A(n10560), .B(n10559), .Z(n10518) );
  XOR U11570 ( .A(n10517), .B(n10518), .Z(n10520) );
  XNOR U11571 ( .A(n10519), .B(n10520), .Z(n10550) );
  XOR U11572 ( .A(n10549), .B(n10550), .Z(n10606) );
  XNOR U11573 ( .A(n10605), .B(n10606), .Z(n10607) );
  XOR U11574 ( .A(n10608), .B(n10607), .Z(n10612) );
  XNOR U11575 ( .A(n10611), .B(n10612), .Z(n10613) );
  XNOR U11576 ( .A(n10614), .B(n10613), .Z(n10618) );
  NANDN U11577 ( .A(n10455), .B(n10454), .Z(n10459) );
  NAND U11578 ( .A(n10457), .B(n10456), .Z(n10458) );
  NAND U11579 ( .A(n10459), .B(n10458), .Z(n10615) );
  NANDN U11580 ( .A(n10461), .B(n10460), .Z(n10465) );
  NAND U11581 ( .A(n10463), .B(n10462), .Z(n10464) );
  NAND U11582 ( .A(n10465), .B(n10464), .Z(n10616) );
  XNOR U11583 ( .A(n10615), .B(n10616), .Z(n10617) );
  XNOR U11584 ( .A(n10618), .B(n10617), .Z(n10490) );
  NANDN U11585 ( .A(n10467), .B(n10466), .Z(n10471) );
  NANDN U11586 ( .A(n10469), .B(n10468), .Z(n10470) );
  NAND U11587 ( .A(n10471), .B(n10470), .Z(n10488) );
  OR U11588 ( .A(n10473), .B(n10472), .Z(n10477) );
  OR U11589 ( .A(n10475), .B(n10474), .Z(n10476) );
  AND U11590 ( .A(n10477), .B(n10476), .Z(n10487) );
  XNOR U11591 ( .A(n10488), .B(n10487), .Z(n10489) );
  XNOR U11592 ( .A(n10490), .B(n10489), .Z(n10483) );
  XOR U11593 ( .A(n10484), .B(n10483), .Z(n10485) );
  XNOR U11594 ( .A(n10486), .B(n10485), .Z(n10621) );
  XNOR U11595 ( .A(n10621), .B(sreg[304]), .Z(n10623) );
  NAND U11596 ( .A(n10478), .B(sreg[303]), .Z(n10482) );
  OR U11597 ( .A(n10480), .B(n10479), .Z(n10481) );
  AND U11598 ( .A(n10482), .B(n10481), .Z(n10622) );
  XOR U11599 ( .A(n10623), .B(n10622), .Z(c[304]) );
  NANDN U11600 ( .A(n10488), .B(n10487), .Z(n10492) );
  NANDN U11601 ( .A(n10490), .B(n10489), .Z(n10491) );
  NAND U11602 ( .A(n10492), .B(n10491), .Z(n10627) );
  NANDN U11603 ( .A(n10494), .B(n10493), .Z(n10498) );
  NAND U11604 ( .A(n10496), .B(n10495), .Z(n10497) );
  NAND U11605 ( .A(n10498), .B(n10497), .Z(n10693) );
  XNOR U11606 ( .A(b[19]), .B(a[63]), .Z(n10644) );
  NANDN U11607 ( .A(n10644), .B(n37934), .Z(n10501) );
  NANDN U11608 ( .A(n10499), .B(n37935), .Z(n10500) );
  NAND U11609 ( .A(n10501), .B(n10500), .Z(n10703) );
  XOR U11610 ( .A(b[27]), .B(a[55]), .Z(n10647) );
  NAND U11611 ( .A(n38423), .B(n10647), .Z(n10504) );
  NANDN U11612 ( .A(n10502), .B(n38424), .Z(n10503) );
  NAND U11613 ( .A(n10504), .B(n10503), .Z(n10700) );
  XNOR U11614 ( .A(b[5]), .B(a[77]), .Z(n10650) );
  NANDN U11615 ( .A(n10650), .B(n36587), .Z(n10507) );
  NANDN U11616 ( .A(n10505), .B(n36588), .Z(n10506) );
  AND U11617 ( .A(n10507), .B(n10506), .Z(n10701) );
  XNOR U11618 ( .A(n10700), .B(n10701), .Z(n10702) );
  XNOR U11619 ( .A(n10703), .B(n10702), .Z(n10691) );
  NAND U11620 ( .A(n10508), .B(n37762), .Z(n10510) );
  XOR U11621 ( .A(b[17]), .B(a[65]), .Z(n10653) );
  NAND U11622 ( .A(n10653), .B(n37764), .Z(n10509) );
  NAND U11623 ( .A(n10510), .B(n10509), .Z(n10671) );
  XNOR U11624 ( .A(b[31]), .B(a[51]), .Z(n10656) );
  NANDN U11625 ( .A(n10656), .B(n38552), .Z(n10513) );
  NANDN U11626 ( .A(n10511), .B(n38553), .Z(n10512) );
  NAND U11627 ( .A(n10513), .B(n10512), .Z(n10668) );
  OR U11628 ( .A(n10514), .B(n36105), .Z(n10516) );
  XNOR U11629 ( .A(b[3]), .B(a[79]), .Z(n10659) );
  NANDN U11630 ( .A(n10659), .B(n36107), .Z(n10515) );
  AND U11631 ( .A(n10516), .B(n10515), .Z(n10669) );
  XNOR U11632 ( .A(n10668), .B(n10669), .Z(n10670) );
  XOR U11633 ( .A(n10671), .B(n10670), .Z(n10690) );
  XNOR U11634 ( .A(n10691), .B(n10690), .Z(n10692) );
  XNOR U11635 ( .A(n10693), .B(n10692), .Z(n10743) );
  NANDN U11636 ( .A(n10518), .B(n10517), .Z(n10522) );
  OR U11637 ( .A(n10520), .B(n10519), .Z(n10521) );
  NAND U11638 ( .A(n10522), .B(n10521), .Z(n10744) );
  XNOR U11639 ( .A(n10743), .B(n10744), .Z(n10745) );
  NANDN U11640 ( .A(n10524), .B(n10523), .Z(n10528) );
  NAND U11641 ( .A(n10526), .B(n10525), .Z(n10527) );
  NAND U11642 ( .A(n10528), .B(n10527), .Z(n10740) );
  OR U11643 ( .A(n10530), .B(n10529), .Z(n10534) );
  NAND U11644 ( .A(n10532), .B(n10531), .Z(n10533) );
  AND U11645 ( .A(n10534), .B(n10533), .Z(n10737) );
  OR U11646 ( .A(n10536), .B(n10535), .Z(n10540) );
  NANDN U11647 ( .A(n10538), .B(n10537), .Z(n10539) );
  NAND U11648 ( .A(n10540), .B(n10539), .Z(n10738) );
  XOR U11649 ( .A(n10740), .B(n10739), .Z(n10746) );
  XNOR U11650 ( .A(n10745), .B(n10746), .Z(n10762) );
  OR U11651 ( .A(n10542), .B(n10541), .Z(n10546) );
  NAND U11652 ( .A(n10544), .B(n10543), .Z(n10545) );
  NAND U11653 ( .A(n10546), .B(n10545), .Z(n10760) );
  NANDN U11654 ( .A(n10548), .B(n10547), .Z(n10552) );
  NANDN U11655 ( .A(n10550), .B(n10549), .Z(n10551) );
  NAND U11656 ( .A(n10552), .B(n10551), .Z(n10749) );
  NANDN U11657 ( .A(n10558), .B(n10557), .Z(n10562) );
  NAND U11658 ( .A(n10560), .B(n10559), .Z(n10561) );
  NAND U11659 ( .A(n10562), .B(n10561), .Z(n10684) );
  NANDN U11660 ( .A(n10564), .B(n10563), .Z(n10568) );
  NAND U11661 ( .A(n10566), .B(n10565), .Z(n10567) );
  AND U11662 ( .A(n10568), .B(n10567), .Z(n10685) );
  XNOR U11663 ( .A(n10684), .B(n10685), .Z(n10686) );
  XNOR U11664 ( .A(b[9]), .B(a[73]), .Z(n10706) );
  NANDN U11665 ( .A(n10706), .B(n36925), .Z(n10571) );
  NAND U11666 ( .A(n36926), .B(n10569), .Z(n10570) );
  NAND U11667 ( .A(n10571), .B(n10570), .Z(n10676) );
  XNOR U11668 ( .A(n1054), .B(a[67]), .Z(n10709) );
  NANDN U11669 ( .A(n37665), .B(n10709), .Z(n10574) );
  NANDN U11670 ( .A(n10572), .B(n37604), .Z(n10573) );
  NAND U11671 ( .A(n10574), .B(n10573), .Z(n10674) );
  XNOR U11672 ( .A(b[21]), .B(a[61]), .Z(n10712) );
  NANDN U11673 ( .A(n10712), .B(n38101), .Z(n10577) );
  NAND U11674 ( .A(n38102), .B(n10575), .Z(n10576) );
  NAND U11675 ( .A(n10577), .B(n10576), .Z(n10675) );
  XNOR U11676 ( .A(n10674), .B(n10675), .Z(n10677) );
  XOR U11677 ( .A(n10676), .B(n10677), .Z(n10665) );
  XNOR U11678 ( .A(b[11]), .B(a[71]), .Z(n10715) );
  OR U11679 ( .A(n10715), .B(n37311), .Z(n10580) );
  NANDN U11680 ( .A(n10578), .B(n37218), .Z(n10579) );
  NAND U11681 ( .A(n10580), .B(n10579), .Z(n10663) );
  XOR U11682 ( .A(n1053), .B(a[69]), .Z(n10718) );
  NANDN U11683 ( .A(n10718), .B(n37424), .Z(n10583) );
  NANDN U11684 ( .A(n10581), .B(n37425), .Z(n10582) );
  AND U11685 ( .A(n10583), .B(n10582), .Z(n10662) );
  XNOR U11686 ( .A(n10663), .B(n10662), .Z(n10664) );
  XNOR U11687 ( .A(n10665), .B(n10664), .Z(n10681) );
  NANDN U11688 ( .A(n1049), .B(a[81]), .Z(n10584) );
  XNOR U11689 ( .A(b[1]), .B(n10584), .Z(n10586) );
  IV U11690 ( .A(a[80]), .Z(n15068) );
  NANDN U11691 ( .A(n15068), .B(n1049), .Z(n10585) );
  AND U11692 ( .A(n10586), .B(n10585), .Z(n10640) );
  NAND U11693 ( .A(n38490), .B(n10587), .Z(n10589) );
  XNOR U11694 ( .A(b[29]), .B(a[53]), .Z(n10725) );
  OR U11695 ( .A(n10725), .B(n1048), .Z(n10588) );
  NAND U11696 ( .A(n10589), .B(n10588), .Z(n10638) );
  NANDN U11697 ( .A(n1059), .B(a[49]), .Z(n10639) );
  XNOR U11698 ( .A(n10638), .B(n10639), .Z(n10641) );
  XNOR U11699 ( .A(n10640), .B(n10641), .Z(n10679) );
  NANDN U11700 ( .A(n10590), .B(n38205), .Z(n10592) );
  XOR U11701 ( .A(b[23]), .B(n12056), .Z(n10728) );
  OR U11702 ( .A(n10728), .B(n38268), .Z(n10591) );
  NAND U11703 ( .A(n10592), .B(n10591), .Z(n10697) );
  XOR U11704 ( .A(b[7]), .B(a[75]), .Z(n10731) );
  NAND U11705 ( .A(n10731), .B(n36701), .Z(n10595) );
  NAND U11706 ( .A(n10593), .B(n36702), .Z(n10594) );
  NAND U11707 ( .A(n10595), .B(n10594), .Z(n10694) );
  XOR U11708 ( .A(b[25]), .B(a[57]), .Z(n10734) );
  NAND U11709 ( .A(n10734), .B(n38325), .Z(n10598) );
  NAND U11710 ( .A(n10596), .B(n38326), .Z(n10597) );
  AND U11711 ( .A(n10598), .B(n10597), .Z(n10695) );
  XNOR U11712 ( .A(n10694), .B(n10695), .Z(n10696) );
  XOR U11713 ( .A(n10697), .B(n10696), .Z(n10678) );
  XOR U11714 ( .A(n10681), .B(n10680), .Z(n10687) );
  XOR U11715 ( .A(n10686), .B(n10687), .Z(n10747) );
  XNOR U11716 ( .A(n10748), .B(n10747), .Z(n10750) );
  XNOR U11717 ( .A(n10749), .B(n10750), .Z(n10759) );
  XOR U11718 ( .A(n10760), .B(n10759), .Z(n10761) );
  XNOR U11719 ( .A(n10762), .B(n10761), .Z(n10756) );
  NANDN U11720 ( .A(n10600), .B(n10599), .Z(n10604) );
  NAND U11721 ( .A(n10602), .B(n10601), .Z(n10603) );
  NAND U11722 ( .A(n10604), .B(n10603), .Z(n10753) );
  NANDN U11723 ( .A(n10606), .B(n10605), .Z(n10610) );
  NAND U11724 ( .A(n10608), .B(n10607), .Z(n10609) );
  NAND U11725 ( .A(n10610), .B(n10609), .Z(n10754) );
  XNOR U11726 ( .A(n10753), .B(n10754), .Z(n10755) );
  XOR U11727 ( .A(n10756), .B(n10755), .Z(n10634) );
  NANDN U11728 ( .A(n10616), .B(n10615), .Z(n10620) );
  NANDN U11729 ( .A(n10618), .B(n10617), .Z(n10619) );
  NAND U11730 ( .A(n10620), .B(n10619), .Z(n10633) );
  XNOR U11731 ( .A(n10632), .B(n10633), .Z(n10635) );
  XOR U11732 ( .A(n10634), .B(n10635), .Z(n10626) );
  XOR U11733 ( .A(n10627), .B(n10626), .Z(n10628) );
  XNOR U11734 ( .A(n10629), .B(n10628), .Z(n10765) );
  XNOR U11735 ( .A(n10765), .B(sreg[305]), .Z(n10767) );
  NAND U11736 ( .A(n10621), .B(sreg[304]), .Z(n10625) );
  OR U11737 ( .A(n10623), .B(n10622), .Z(n10624) );
  AND U11738 ( .A(n10625), .B(n10624), .Z(n10766) );
  XOR U11739 ( .A(n10767), .B(n10766), .Z(c[305]) );
  NAND U11740 ( .A(n10627), .B(n10626), .Z(n10631) );
  NAND U11741 ( .A(n10629), .B(n10628), .Z(n10630) );
  NAND U11742 ( .A(n10631), .B(n10630), .Z(n10773) );
  NANDN U11743 ( .A(n10633), .B(n10632), .Z(n10637) );
  NAND U11744 ( .A(n10635), .B(n10634), .Z(n10636) );
  NAND U11745 ( .A(n10637), .B(n10636), .Z(n10771) );
  NANDN U11746 ( .A(n10639), .B(n10638), .Z(n10643) );
  NAND U11747 ( .A(n10641), .B(n10640), .Z(n10642) );
  NAND U11748 ( .A(n10643), .B(n10642), .Z(n10853) );
  XNOR U11749 ( .A(b[19]), .B(a[64]), .Z(n10822) );
  NANDN U11750 ( .A(n10822), .B(n37934), .Z(n10646) );
  NANDN U11751 ( .A(n10644), .B(n37935), .Z(n10645) );
  NAND U11752 ( .A(n10646), .B(n10645), .Z(n10865) );
  XOR U11753 ( .A(b[27]), .B(a[56]), .Z(n10825) );
  NAND U11754 ( .A(n38423), .B(n10825), .Z(n10649) );
  NAND U11755 ( .A(n10647), .B(n38424), .Z(n10648) );
  NAND U11756 ( .A(n10649), .B(n10648), .Z(n10862) );
  XNOR U11757 ( .A(b[5]), .B(a[78]), .Z(n10828) );
  NANDN U11758 ( .A(n10828), .B(n36587), .Z(n10652) );
  NANDN U11759 ( .A(n10650), .B(n36588), .Z(n10651) );
  AND U11760 ( .A(n10652), .B(n10651), .Z(n10863) );
  XNOR U11761 ( .A(n10862), .B(n10863), .Z(n10864) );
  XNOR U11762 ( .A(n10865), .B(n10864), .Z(n10850) );
  NAND U11763 ( .A(n10653), .B(n37762), .Z(n10655) );
  XOR U11764 ( .A(b[17]), .B(a[66]), .Z(n10831) );
  NAND U11765 ( .A(n10831), .B(n37764), .Z(n10654) );
  NAND U11766 ( .A(n10655), .B(n10654), .Z(n10806) );
  XNOR U11767 ( .A(b[31]), .B(a[52]), .Z(n10834) );
  NANDN U11768 ( .A(n10834), .B(n38552), .Z(n10658) );
  NANDN U11769 ( .A(n10656), .B(n38553), .Z(n10657) );
  AND U11770 ( .A(n10658), .B(n10657), .Z(n10804) );
  OR U11771 ( .A(n10659), .B(n36105), .Z(n10661) );
  XOR U11772 ( .A(b[3]), .B(n15068), .Z(n10837) );
  NANDN U11773 ( .A(n10837), .B(n36107), .Z(n10660) );
  AND U11774 ( .A(n10661), .B(n10660), .Z(n10805) );
  XOR U11775 ( .A(n10806), .B(n10807), .Z(n10851) );
  XOR U11776 ( .A(n10850), .B(n10851), .Z(n10852) );
  XNOR U11777 ( .A(n10853), .B(n10852), .Z(n10789) );
  NANDN U11778 ( .A(n10663), .B(n10662), .Z(n10667) );
  NAND U11779 ( .A(n10665), .B(n10664), .Z(n10666) );
  NAND U11780 ( .A(n10667), .B(n10666), .Z(n10842) );
  NANDN U11781 ( .A(n10669), .B(n10668), .Z(n10673) );
  NAND U11782 ( .A(n10671), .B(n10670), .Z(n10672) );
  NAND U11783 ( .A(n10673), .B(n10672), .Z(n10841) );
  XNOR U11784 ( .A(n10841), .B(n10840), .Z(n10843) );
  XOR U11785 ( .A(n10842), .B(n10843), .Z(n10788) );
  XOR U11786 ( .A(n10789), .B(n10788), .Z(n10790) );
  NANDN U11787 ( .A(n10679), .B(n10678), .Z(n10683) );
  NAND U11788 ( .A(n10681), .B(n10680), .Z(n10682) );
  NAND U11789 ( .A(n10683), .B(n10682), .Z(n10791) );
  XNOR U11790 ( .A(n10790), .B(n10791), .Z(n10906) );
  NANDN U11791 ( .A(n10685), .B(n10684), .Z(n10689) );
  NAND U11792 ( .A(n10687), .B(n10686), .Z(n10688) );
  NAND U11793 ( .A(n10689), .B(n10688), .Z(n10784) );
  NANDN U11794 ( .A(n10695), .B(n10694), .Z(n10699) );
  NAND U11795 ( .A(n10697), .B(n10696), .Z(n10698) );
  NAND U11796 ( .A(n10699), .B(n10698), .Z(n10844) );
  NANDN U11797 ( .A(n10701), .B(n10700), .Z(n10705) );
  NAND U11798 ( .A(n10703), .B(n10702), .Z(n10704) );
  AND U11799 ( .A(n10705), .B(n10704), .Z(n10845) );
  XNOR U11800 ( .A(n10844), .B(n10845), .Z(n10846) );
  XNOR U11801 ( .A(b[9]), .B(a[74]), .Z(n10868) );
  NANDN U11802 ( .A(n10868), .B(n36925), .Z(n10708) );
  NANDN U11803 ( .A(n10706), .B(n36926), .Z(n10707) );
  NAND U11804 ( .A(n10708), .B(n10707), .Z(n10812) );
  XNOR U11805 ( .A(b[15]), .B(a[68]), .Z(n10871) );
  OR U11806 ( .A(n10871), .B(n37665), .Z(n10711) );
  NAND U11807 ( .A(n10709), .B(n37604), .Z(n10710) );
  AND U11808 ( .A(n10711), .B(n10710), .Z(n10810) );
  XOR U11809 ( .A(b[21]), .B(n12493), .Z(n10874) );
  NANDN U11810 ( .A(n10874), .B(n38101), .Z(n10714) );
  NANDN U11811 ( .A(n10712), .B(n38102), .Z(n10713) );
  AND U11812 ( .A(n10714), .B(n10713), .Z(n10811) );
  XOR U11813 ( .A(n10812), .B(n10813), .Z(n10801) );
  XNOR U11814 ( .A(b[11]), .B(a[72]), .Z(n10877) );
  OR U11815 ( .A(n10877), .B(n37311), .Z(n10717) );
  NANDN U11816 ( .A(n10715), .B(n37218), .Z(n10716) );
  NAND U11817 ( .A(n10717), .B(n10716), .Z(n10799) );
  XOR U11818 ( .A(n1053), .B(a[70]), .Z(n10880) );
  NANDN U11819 ( .A(n10880), .B(n37424), .Z(n10720) );
  NANDN U11820 ( .A(n10718), .B(n37425), .Z(n10719) );
  NAND U11821 ( .A(n10720), .B(n10719), .Z(n10798) );
  XOR U11822 ( .A(n10801), .B(n10800), .Z(n10795) );
  NANDN U11823 ( .A(n1049), .B(a[82]), .Z(n10721) );
  XNOR U11824 ( .A(b[1]), .B(n10721), .Z(n10723) );
  NANDN U11825 ( .A(b[0]), .B(a[81]), .Z(n10722) );
  AND U11826 ( .A(n10723), .B(n10722), .Z(n10819) );
  ANDN U11827 ( .B(b[31]), .A(n10724), .Z(n10816) );
  NANDN U11828 ( .A(n10725), .B(n38490), .Z(n10727) );
  XNOR U11829 ( .A(n1058), .B(a[54]), .Z(n10883) );
  NANDN U11830 ( .A(n1048), .B(n10883), .Z(n10726) );
  NAND U11831 ( .A(n10727), .B(n10726), .Z(n10817) );
  XOR U11832 ( .A(n10816), .B(n10817), .Z(n10818) );
  XNOR U11833 ( .A(n10819), .B(n10818), .Z(n10792) );
  NANDN U11834 ( .A(n10728), .B(n38205), .Z(n10730) );
  XNOR U11835 ( .A(b[23]), .B(a[60]), .Z(n10889) );
  OR U11836 ( .A(n10889), .B(n38268), .Z(n10729) );
  NAND U11837 ( .A(n10730), .B(n10729), .Z(n10859) );
  XOR U11838 ( .A(b[7]), .B(a[76]), .Z(n10892) );
  NAND U11839 ( .A(n10892), .B(n36701), .Z(n10733) );
  NAND U11840 ( .A(n10731), .B(n36702), .Z(n10732) );
  NAND U11841 ( .A(n10733), .B(n10732), .Z(n10856) );
  XOR U11842 ( .A(b[25]), .B(a[58]), .Z(n10895) );
  NAND U11843 ( .A(n10895), .B(n38325), .Z(n10736) );
  NAND U11844 ( .A(n10734), .B(n38326), .Z(n10735) );
  AND U11845 ( .A(n10736), .B(n10735), .Z(n10857) );
  XNOR U11846 ( .A(n10856), .B(n10857), .Z(n10858) );
  XNOR U11847 ( .A(n10859), .B(n10858), .Z(n10793) );
  XOR U11848 ( .A(n10795), .B(n10794), .Z(n10847) );
  XNOR U11849 ( .A(n10846), .B(n10847), .Z(n10782) );
  XNOR U11850 ( .A(n10783), .B(n10782), .Z(n10785) );
  XNOR U11851 ( .A(n10784), .B(n10785), .Z(n10904) );
  OR U11852 ( .A(n10738), .B(n10737), .Z(n10742) );
  NANDN U11853 ( .A(n10740), .B(n10739), .Z(n10741) );
  NAND U11854 ( .A(n10742), .B(n10741), .Z(n10905) );
  XOR U11855 ( .A(n10904), .B(n10905), .Z(n10907) );
  NAND U11856 ( .A(n10748), .B(n10747), .Z(n10752) );
  NANDN U11857 ( .A(n10750), .B(n10749), .Z(n10751) );
  NAND U11858 ( .A(n10752), .B(n10751), .Z(n10899) );
  XNOR U11859 ( .A(n10898), .B(n10899), .Z(n10900) );
  XOR U11860 ( .A(n10901), .B(n10900), .Z(n10778) );
  NANDN U11861 ( .A(n10754), .B(n10753), .Z(n10758) );
  NAND U11862 ( .A(n10756), .B(n10755), .Z(n10757) );
  NAND U11863 ( .A(n10758), .B(n10757), .Z(n10776) );
  NANDN U11864 ( .A(n10760), .B(n10759), .Z(n10764) );
  OR U11865 ( .A(n10762), .B(n10761), .Z(n10763) );
  NAND U11866 ( .A(n10764), .B(n10763), .Z(n10777) );
  XNOR U11867 ( .A(n10776), .B(n10777), .Z(n10779) );
  XOR U11868 ( .A(n10778), .B(n10779), .Z(n10770) );
  XOR U11869 ( .A(n10771), .B(n10770), .Z(n10772) );
  XNOR U11870 ( .A(n10773), .B(n10772), .Z(n10910) );
  XNOR U11871 ( .A(n10910), .B(sreg[306]), .Z(n10912) );
  NAND U11872 ( .A(n10765), .B(sreg[305]), .Z(n10769) );
  OR U11873 ( .A(n10767), .B(n10766), .Z(n10768) );
  AND U11874 ( .A(n10769), .B(n10768), .Z(n10911) );
  XOR U11875 ( .A(n10912), .B(n10911), .Z(c[306]) );
  NAND U11876 ( .A(n10771), .B(n10770), .Z(n10775) );
  NAND U11877 ( .A(n10773), .B(n10772), .Z(n10774) );
  NAND U11878 ( .A(n10775), .B(n10774), .Z(n10918) );
  NANDN U11879 ( .A(n10777), .B(n10776), .Z(n10781) );
  NAND U11880 ( .A(n10779), .B(n10778), .Z(n10780) );
  NAND U11881 ( .A(n10781), .B(n10780), .Z(n10915) );
  NAND U11882 ( .A(n10783), .B(n10782), .Z(n10787) );
  NANDN U11883 ( .A(n10785), .B(n10784), .Z(n10786) );
  NAND U11884 ( .A(n10787), .B(n10786), .Z(n11047) );
  XNOR U11885 ( .A(n11047), .B(n11048), .Z(n11049) );
  OR U11886 ( .A(n10793), .B(n10792), .Z(n10797) );
  NANDN U11887 ( .A(n10795), .B(n10794), .Z(n10796) );
  NAND U11888 ( .A(n10797), .B(n10796), .Z(n11038) );
  OR U11889 ( .A(n10799), .B(n10798), .Z(n10803) );
  NAND U11890 ( .A(n10801), .B(n10800), .Z(n10802) );
  NAND U11891 ( .A(n10803), .B(n10802), .Z(n10977) );
  OR U11892 ( .A(n10805), .B(n10804), .Z(n10809) );
  NANDN U11893 ( .A(n10807), .B(n10806), .Z(n10808) );
  NAND U11894 ( .A(n10809), .B(n10808), .Z(n10976) );
  OR U11895 ( .A(n10811), .B(n10810), .Z(n10815) );
  NANDN U11896 ( .A(n10813), .B(n10812), .Z(n10814) );
  NAND U11897 ( .A(n10815), .B(n10814), .Z(n10975) );
  XOR U11898 ( .A(n10977), .B(n10978), .Z(n11036) );
  OR U11899 ( .A(n10817), .B(n10816), .Z(n10821) );
  NANDN U11900 ( .A(n10819), .B(n10818), .Z(n10820) );
  NAND U11901 ( .A(n10821), .B(n10820), .Z(n10989) );
  XNOR U11902 ( .A(b[19]), .B(a[65]), .Z(n10933) );
  NANDN U11903 ( .A(n10933), .B(n37934), .Z(n10824) );
  NANDN U11904 ( .A(n10822), .B(n37935), .Z(n10823) );
  NAND U11905 ( .A(n10824), .B(n10823), .Z(n11002) );
  XOR U11906 ( .A(b[27]), .B(a[57]), .Z(n10936) );
  NAND U11907 ( .A(n38423), .B(n10936), .Z(n10827) );
  NAND U11908 ( .A(n10825), .B(n38424), .Z(n10826) );
  NAND U11909 ( .A(n10827), .B(n10826), .Z(n10999) );
  XNOR U11910 ( .A(b[5]), .B(a[79]), .Z(n10939) );
  NANDN U11911 ( .A(n10939), .B(n36587), .Z(n10830) );
  NANDN U11912 ( .A(n10828), .B(n36588), .Z(n10829) );
  AND U11913 ( .A(n10830), .B(n10829), .Z(n11000) );
  XNOR U11914 ( .A(n10999), .B(n11000), .Z(n11001) );
  XNOR U11915 ( .A(n11002), .B(n11001), .Z(n10988) );
  NAND U11916 ( .A(n10831), .B(n37762), .Z(n10833) );
  XNOR U11917 ( .A(b[17]), .B(a[67]), .Z(n10942) );
  NANDN U11918 ( .A(n10942), .B(n37764), .Z(n10832) );
  NAND U11919 ( .A(n10833), .B(n10832), .Z(n10960) );
  XNOR U11920 ( .A(b[31]), .B(a[53]), .Z(n10945) );
  NANDN U11921 ( .A(n10945), .B(n38552), .Z(n10836) );
  NANDN U11922 ( .A(n10834), .B(n38553), .Z(n10835) );
  NAND U11923 ( .A(n10836), .B(n10835), .Z(n10957) );
  OR U11924 ( .A(n10837), .B(n36105), .Z(n10839) );
  XNOR U11925 ( .A(b[3]), .B(a[81]), .Z(n10948) );
  NANDN U11926 ( .A(n10948), .B(n36107), .Z(n10838) );
  AND U11927 ( .A(n10839), .B(n10838), .Z(n10958) );
  XNOR U11928 ( .A(n10957), .B(n10958), .Z(n10959) );
  XOR U11929 ( .A(n10960), .B(n10959), .Z(n10987) );
  XOR U11930 ( .A(n10988), .B(n10987), .Z(n10990) );
  XOR U11931 ( .A(n10989), .B(n10990), .Z(n11035) );
  XOR U11932 ( .A(n11036), .B(n11035), .Z(n11037) );
  XNOR U11933 ( .A(n11038), .B(n11037), .Z(n11056) );
  NANDN U11934 ( .A(n10845), .B(n10844), .Z(n10849) );
  NANDN U11935 ( .A(n10847), .B(n10846), .Z(n10848) );
  NAND U11936 ( .A(n10849), .B(n10848), .Z(n11043) );
  OR U11937 ( .A(n10851), .B(n10850), .Z(n10855) );
  NAND U11938 ( .A(n10853), .B(n10852), .Z(n10854) );
  NAND U11939 ( .A(n10855), .B(n10854), .Z(n11042) );
  NANDN U11940 ( .A(n10857), .B(n10856), .Z(n10861) );
  NAND U11941 ( .A(n10859), .B(n10858), .Z(n10860) );
  NAND U11942 ( .A(n10861), .B(n10860), .Z(n10981) );
  NANDN U11943 ( .A(n10863), .B(n10862), .Z(n10867) );
  NAND U11944 ( .A(n10865), .B(n10864), .Z(n10866) );
  AND U11945 ( .A(n10867), .B(n10866), .Z(n10982) );
  XNOR U11946 ( .A(n10981), .B(n10982), .Z(n10983) );
  XNOR U11947 ( .A(b[9]), .B(a[75]), .Z(n11005) );
  NANDN U11948 ( .A(n11005), .B(n36925), .Z(n10870) );
  NANDN U11949 ( .A(n10868), .B(n36926), .Z(n10869) );
  NAND U11950 ( .A(n10870), .B(n10869), .Z(n10965) );
  XNOR U11951 ( .A(b[15]), .B(a[69]), .Z(n11008) );
  OR U11952 ( .A(n11008), .B(n37665), .Z(n10873) );
  NANDN U11953 ( .A(n10871), .B(n37604), .Z(n10872) );
  AND U11954 ( .A(n10873), .B(n10872), .Z(n10963) );
  XNOR U11955 ( .A(b[21]), .B(a[63]), .Z(n11011) );
  NANDN U11956 ( .A(n11011), .B(n38101), .Z(n10876) );
  NANDN U11957 ( .A(n10874), .B(n38102), .Z(n10875) );
  AND U11958 ( .A(n10876), .B(n10875), .Z(n10964) );
  XOR U11959 ( .A(n10965), .B(n10966), .Z(n10954) );
  XNOR U11960 ( .A(b[11]), .B(a[73]), .Z(n11014) );
  OR U11961 ( .A(n11014), .B(n37311), .Z(n10879) );
  NANDN U11962 ( .A(n10877), .B(n37218), .Z(n10878) );
  NAND U11963 ( .A(n10879), .B(n10878), .Z(n10952) );
  XOR U11964 ( .A(n1053), .B(a[71]), .Z(n11017) );
  NANDN U11965 ( .A(n11017), .B(n37424), .Z(n10882) );
  NANDN U11966 ( .A(n10880), .B(n37425), .Z(n10881) );
  AND U11967 ( .A(n10882), .B(n10881), .Z(n10951) );
  XNOR U11968 ( .A(n10952), .B(n10951), .Z(n10953) );
  XOR U11969 ( .A(n10954), .B(n10953), .Z(n10971) );
  NAND U11970 ( .A(n10883), .B(n38490), .Z(n10885) );
  XNOR U11971 ( .A(n1058), .B(a[55]), .Z(n11023) );
  NANDN U11972 ( .A(n1048), .B(n11023), .Z(n10884) );
  NAND U11973 ( .A(n10885), .B(n10884), .Z(n10927) );
  NANDN U11974 ( .A(n1059), .B(a[51]), .Z(n10928) );
  XNOR U11975 ( .A(n10927), .B(n10928), .Z(n10930) );
  NANDN U11976 ( .A(n1049), .B(a[83]), .Z(n10886) );
  XNOR U11977 ( .A(b[1]), .B(n10886), .Z(n10888) );
  IV U11978 ( .A(a[82]), .Z(n15424) );
  NANDN U11979 ( .A(n15424), .B(n1049), .Z(n10887) );
  AND U11980 ( .A(n10888), .B(n10887), .Z(n10929) );
  XOR U11981 ( .A(n10930), .B(n10929), .Z(n10969) );
  NANDN U11982 ( .A(n10889), .B(n38205), .Z(n10891) );
  XNOR U11983 ( .A(b[23]), .B(a[61]), .Z(n11026) );
  OR U11984 ( .A(n11026), .B(n38268), .Z(n10890) );
  NAND U11985 ( .A(n10891), .B(n10890), .Z(n10996) );
  XOR U11986 ( .A(b[7]), .B(a[77]), .Z(n11029) );
  NAND U11987 ( .A(n11029), .B(n36701), .Z(n10894) );
  NAND U11988 ( .A(n10892), .B(n36702), .Z(n10893) );
  NAND U11989 ( .A(n10894), .B(n10893), .Z(n10993) );
  XNOR U11990 ( .A(b[25]), .B(a[59]), .Z(n11032) );
  NANDN U11991 ( .A(n11032), .B(n38325), .Z(n10897) );
  NAND U11992 ( .A(n10895), .B(n38326), .Z(n10896) );
  AND U11993 ( .A(n10897), .B(n10896), .Z(n10994) );
  XNOR U11994 ( .A(n10993), .B(n10994), .Z(n10995) );
  XNOR U11995 ( .A(n10996), .B(n10995), .Z(n10970) );
  XOR U11996 ( .A(n10969), .B(n10970), .Z(n10972) );
  XNOR U11997 ( .A(n10971), .B(n10972), .Z(n10984) );
  XNOR U11998 ( .A(n10983), .B(n10984), .Z(n11041) );
  XNOR U11999 ( .A(n11042), .B(n11041), .Z(n11044) );
  XNOR U12000 ( .A(n11043), .B(n11044), .Z(n11053) );
  XNOR U12001 ( .A(n11054), .B(n11053), .Z(n11055) );
  XOR U12002 ( .A(n11056), .B(n11055), .Z(n11050) );
  XOR U12003 ( .A(n11049), .B(n11050), .Z(n10924) );
  NANDN U12004 ( .A(n10899), .B(n10898), .Z(n10903) );
  NAND U12005 ( .A(n10901), .B(n10900), .Z(n10902) );
  NAND U12006 ( .A(n10903), .B(n10902), .Z(n10921) );
  NANDN U12007 ( .A(n10905), .B(n10904), .Z(n10909) );
  OR U12008 ( .A(n10907), .B(n10906), .Z(n10908) );
  NAND U12009 ( .A(n10909), .B(n10908), .Z(n10922) );
  XNOR U12010 ( .A(n10921), .B(n10922), .Z(n10923) );
  XNOR U12011 ( .A(n10924), .B(n10923), .Z(n10916) );
  XNOR U12012 ( .A(n10915), .B(n10916), .Z(n10917) );
  XNOR U12013 ( .A(n10918), .B(n10917), .Z(n11059) );
  XNOR U12014 ( .A(n11059), .B(sreg[307]), .Z(n11061) );
  NAND U12015 ( .A(n10910), .B(sreg[306]), .Z(n10914) );
  OR U12016 ( .A(n10912), .B(n10911), .Z(n10913) );
  AND U12017 ( .A(n10914), .B(n10913), .Z(n11060) );
  XOR U12018 ( .A(n11061), .B(n11060), .Z(c[307]) );
  NANDN U12019 ( .A(n10916), .B(n10915), .Z(n10920) );
  NAND U12020 ( .A(n10918), .B(n10917), .Z(n10919) );
  NAND U12021 ( .A(n10920), .B(n10919), .Z(n11067) );
  NANDN U12022 ( .A(n10922), .B(n10921), .Z(n10926) );
  NAND U12023 ( .A(n10924), .B(n10923), .Z(n10925) );
  NAND U12024 ( .A(n10926), .B(n10925), .Z(n11065) );
  NANDN U12025 ( .A(n10928), .B(n10927), .Z(n10932) );
  NAND U12026 ( .A(n10930), .B(n10929), .Z(n10931) );
  NAND U12027 ( .A(n10932), .B(n10931), .Z(n11151) );
  XNOR U12028 ( .A(b[19]), .B(a[66]), .Z(n11094) );
  NANDN U12029 ( .A(n11094), .B(n37934), .Z(n10935) );
  NANDN U12030 ( .A(n10933), .B(n37935), .Z(n10934) );
  NAND U12031 ( .A(n10935), .B(n10934), .Z(n11161) );
  XOR U12032 ( .A(b[27]), .B(a[58]), .Z(n11097) );
  NAND U12033 ( .A(n38423), .B(n11097), .Z(n10938) );
  NAND U12034 ( .A(n10936), .B(n38424), .Z(n10937) );
  NAND U12035 ( .A(n10938), .B(n10937), .Z(n11158) );
  XOR U12036 ( .A(b[5]), .B(n15068), .Z(n11100) );
  NANDN U12037 ( .A(n11100), .B(n36587), .Z(n10941) );
  NANDN U12038 ( .A(n10939), .B(n36588), .Z(n10940) );
  AND U12039 ( .A(n10941), .B(n10940), .Z(n11159) );
  XNOR U12040 ( .A(n11158), .B(n11159), .Z(n11160) );
  XNOR U12041 ( .A(n11161), .B(n11160), .Z(n11149) );
  NANDN U12042 ( .A(n10942), .B(n37762), .Z(n10944) );
  XOR U12043 ( .A(b[17]), .B(a[68]), .Z(n11103) );
  NAND U12044 ( .A(n11103), .B(n37764), .Z(n10943) );
  NAND U12045 ( .A(n10944), .B(n10943), .Z(n11121) );
  XOR U12046 ( .A(b[31]), .B(n11319), .Z(n11106) );
  NANDN U12047 ( .A(n11106), .B(n38552), .Z(n10947) );
  NANDN U12048 ( .A(n10945), .B(n38553), .Z(n10946) );
  NAND U12049 ( .A(n10947), .B(n10946), .Z(n11118) );
  OR U12050 ( .A(n10948), .B(n36105), .Z(n10950) );
  XOR U12051 ( .A(b[3]), .B(n15424), .Z(n11109) );
  NANDN U12052 ( .A(n11109), .B(n36107), .Z(n10949) );
  AND U12053 ( .A(n10950), .B(n10949), .Z(n11119) );
  XNOR U12054 ( .A(n11118), .B(n11119), .Z(n11120) );
  XOR U12055 ( .A(n11121), .B(n11120), .Z(n11148) );
  XNOR U12056 ( .A(n11149), .B(n11148), .Z(n11150) );
  XNOR U12057 ( .A(n11151), .B(n11150), .Z(n11194) );
  NANDN U12058 ( .A(n10952), .B(n10951), .Z(n10956) );
  NAND U12059 ( .A(n10954), .B(n10953), .Z(n10955) );
  NAND U12060 ( .A(n10956), .B(n10955), .Z(n11139) );
  NANDN U12061 ( .A(n10958), .B(n10957), .Z(n10962) );
  NAND U12062 ( .A(n10960), .B(n10959), .Z(n10961) );
  NAND U12063 ( .A(n10962), .B(n10961), .Z(n11137) );
  OR U12064 ( .A(n10964), .B(n10963), .Z(n10968) );
  NANDN U12065 ( .A(n10966), .B(n10965), .Z(n10967) );
  NAND U12066 ( .A(n10968), .B(n10967), .Z(n11136) );
  XNOR U12067 ( .A(n11139), .B(n11138), .Z(n11195) );
  XOR U12068 ( .A(n11194), .B(n11195), .Z(n11197) );
  NANDN U12069 ( .A(n10970), .B(n10969), .Z(n10974) );
  OR U12070 ( .A(n10972), .B(n10971), .Z(n10973) );
  NAND U12071 ( .A(n10974), .B(n10973), .Z(n11196) );
  XOR U12072 ( .A(n11197), .B(n11196), .Z(n11084) );
  OR U12073 ( .A(n10976), .B(n10975), .Z(n10980) );
  NANDN U12074 ( .A(n10978), .B(n10977), .Z(n10979) );
  NAND U12075 ( .A(n10980), .B(n10979), .Z(n11083) );
  NANDN U12076 ( .A(n10982), .B(n10981), .Z(n10986) );
  NANDN U12077 ( .A(n10984), .B(n10983), .Z(n10985) );
  NAND U12078 ( .A(n10986), .B(n10985), .Z(n11202) );
  NANDN U12079 ( .A(n10988), .B(n10987), .Z(n10992) );
  OR U12080 ( .A(n10990), .B(n10989), .Z(n10991) );
  NAND U12081 ( .A(n10992), .B(n10991), .Z(n11201) );
  NANDN U12082 ( .A(n10994), .B(n10993), .Z(n10998) );
  NAND U12083 ( .A(n10996), .B(n10995), .Z(n10997) );
  NAND U12084 ( .A(n10998), .B(n10997), .Z(n11142) );
  NANDN U12085 ( .A(n11000), .B(n10999), .Z(n11004) );
  NAND U12086 ( .A(n11002), .B(n11001), .Z(n11003) );
  AND U12087 ( .A(n11004), .B(n11003), .Z(n11143) );
  XNOR U12088 ( .A(n11142), .B(n11143), .Z(n11144) );
  XNOR U12089 ( .A(b[9]), .B(a[76]), .Z(n11164) );
  NANDN U12090 ( .A(n11164), .B(n36925), .Z(n11007) );
  NANDN U12091 ( .A(n11005), .B(n36926), .Z(n11006) );
  NAND U12092 ( .A(n11007), .B(n11006), .Z(n11126) );
  XNOR U12093 ( .A(b[15]), .B(a[70]), .Z(n11167) );
  OR U12094 ( .A(n11167), .B(n37665), .Z(n11010) );
  NANDN U12095 ( .A(n11008), .B(n37604), .Z(n11009) );
  AND U12096 ( .A(n11010), .B(n11009), .Z(n11124) );
  XNOR U12097 ( .A(b[21]), .B(a[64]), .Z(n11170) );
  NANDN U12098 ( .A(n11170), .B(n38101), .Z(n11013) );
  NANDN U12099 ( .A(n11011), .B(n38102), .Z(n11012) );
  AND U12100 ( .A(n11013), .B(n11012), .Z(n11125) );
  XOR U12101 ( .A(n11126), .B(n11127), .Z(n11115) );
  XNOR U12102 ( .A(b[11]), .B(a[74]), .Z(n11173) );
  OR U12103 ( .A(n11173), .B(n37311), .Z(n11016) );
  NANDN U12104 ( .A(n11014), .B(n37218), .Z(n11015) );
  NAND U12105 ( .A(n11016), .B(n11015), .Z(n11113) );
  XOR U12106 ( .A(n1053), .B(a[72]), .Z(n11176) );
  NANDN U12107 ( .A(n11176), .B(n37424), .Z(n11019) );
  NANDN U12108 ( .A(n11017), .B(n37425), .Z(n11018) );
  AND U12109 ( .A(n11019), .B(n11018), .Z(n11112) );
  XNOR U12110 ( .A(n11113), .B(n11112), .Z(n11114) );
  XOR U12111 ( .A(n11115), .B(n11114), .Z(n11132) );
  NANDN U12112 ( .A(n1049), .B(a[84]), .Z(n11020) );
  XNOR U12113 ( .A(b[1]), .B(n11020), .Z(n11022) );
  IV U12114 ( .A(a[83]), .Z(n15562) );
  NANDN U12115 ( .A(n15562), .B(n1049), .Z(n11021) );
  AND U12116 ( .A(n11022), .B(n11021), .Z(n11090) );
  NAND U12117 ( .A(n38490), .B(n11023), .Z(n11025) );
  XNOR U12118 ( .A(n1058), .B(a[56]), .Z(n11182) );
  NANDN U12119 ( .A(n1048), .B(n11182), .Z(n11024) );
  NAND U12120 ( .A(n11025), .B(n11024), .Z(n11088) );
  NANDN U12121 ( .A(n1059), .B(a[52]), .Z(n11089) );
  XNOR U12122 ( .A(n11088), .B(n11089), .Z(n11091) );
  XOR U12123 ( .A(n11090), .B(n11091), .Z(n11130) );
  NANDN U12124 ( .A(n11026), .B(n38205), .Z(n11028) );
  XOR U12125 ( .A(b[23]), .B(n12493), .Z(n11185) );
  OR U12126 ( .A(n11185), .B(n38268), .Z(n11027) );
  NAND U12127 ( .A(n11028), .B(n11027), .Z(n11155) );
  XOR U12128 ( .A(b[7]), .B(a[78]), .Z(n11188) );
  NAND U12129 ( .A(n11188), .B(n36701), .Z(n11031) );
  NAND U12130 ( .A(n11029), .B(n36702), .Z(n11030) );
  NAND U12131 ( .A(n11031), .B(n11030), .Z(n11152) );
  XOR U12132 ( .A(b[25]), .B(a[60]), .Z(n11191) );
  NAND U12133 ( .A(n11191), .B(n38325), .Z(n11034) );
  NANDN U12134 ( .A(n11032), .B(n38326), .Z(n11033) );
  AND U12135 ( .A(n11034), .B(n11033), .Z(n11153) );
  XNOR U12136 ( .A(n11152), .B(n11153), .Z(n11154) );
  XNOR U12137 ( .A(n11155), .B(n11154), .Z(n11131) );
  XOR U12138 ( .A(n11130), .B(n11131), .Z(n11133) );
  XNOR U12139 ( .A(n11132), .B(n11133), .Z(n11145) );
  XNOR U12140 ( .A(n11144), .B(n11145), .Z(n11200) );
  XNOR U12141 ( .A(n11201), .B(n11200), .Z(n11203) );
  XNOR U12142 ( .A(n11202), .B(n11203), .Z(n11082) );
  XOR U12143 ( .A(n11083), .B(n11082), .Z(n11085) );
  NAND U12144 ( .A(n11036), .B(n11035), .Z(n11040) );
  NAND U12145 ( .A(n11038), .B(n11037), .Z(n11039) );
  NAND U12146 ( .A(n11040), .B(n11039), .Z(n11077) );
  NAND U12147 ( .A(n11042), .B(n11041), .Z(n11046) );
  NANDN U12148 ( .A(n11044), .B(n11043), .Z(n11045) );
  AND U12149 ( .A(n11046), .B(n11045), .Z(n11076) );
  XNOR U12150 ( .A(n11077), .B(n11076), .Z(n11078) );
  XOR U12151 ( .A(n11079), .B(n11078), .Z(n11072) );
  NANDN U12152 ( .A(n11048), .B(n11047), .Z(n11052) );
  NANDN U12153 ( .A(n11050), .B(n11049), .Z(n11051) );
  NAND U12154 ( .A(n11052), .B(n11051), .Z(n11071) );
  NANDN U12155 ( .A(n11054), .B(n11053), .Z(n11058) );
  NANDN U12156 ( .A(n11056), .B(n11055), .Z(n11057) );
  AND U12157 ( .A(n11058), .B(n11057), .Z(n11070) );
  XNOR U12158 ( .A(n11071), .B(n11070), .Z(n11073) );
  XOR U12159 ( .A(n11072), .B(n11073), .Z(n11064) );
  XOR U12160 ( .A(n11065), .B(n11064), .Z(n11066) );
  XNOR U12161 ( .A(n11067), .B(n11066), .Z(n11206) );
  XNOR U12162 ( .A(n11206), .B(sreg[308]), .Z(n11208) );
  NAND U12163 ( .A(n11059), .B(sreg[307]), .Z(n11063) );
  OR U12164 ( .A(n11061), .B(n11060), .Z(n11062) );
  AND U12165 ( .A(n11063), .B(n11062), .Z(n11207) );
  XOR U12166 ( .A(n11208), .B(n11207), .Z(c[308]) );
  NAND U12167 ( .A(n11065), .B(n11064), .Z(n11069) );
  NAND U12168 ( .A(n11067), .B(n11066), .Z(n11068) );
  NAND U12169 ( .A(n11069), .B(n11068), .Z(n11214) );
  NANDN U12170 ( .A(n11071), .B(n11070), .Z(n11075) );
  NAND U12171 ( .A(n11073), .B(n11072), .Z(n11074) );
  NAND U12172 ( .A(n11075), .B(n11074), .Z(n11212) );
  NANDN U12173 ( .A(n11077), .B(n11076), .Z(n11081) );
  NAND U12174 ( .A(n11079), .B(n11078), .Z(n11080) );
  NAND U12175 ( .A(n11081), .B(n11080), .Z(n11217) );
  NANDN U12176 ( .A(n11083), .B(n11082), .Z(n11087) );
  OR U12177 ( .A(n11085), .B(n11084), .Z(n11086) );
  NAND U12178 ( .A(n11087), .B(n11086), .Z(n11218) );
  XNOR U12179 ( .A(n11217), .B(n11218), .Z(n11219) );
  NANDN U12180 ( .A(n11089), .B(n11088), .Z(n11093) );
  NAND U12181 ( .A(n11091), .B(n11090), .Z(n11092) );
  NAND U12182 ( .A(n11093), .B(n11092), .Z(n11286) );
  XOR U12183 ( .A(b[19]), .B(n13219), .Z(n11253) );
  NANDN U12184 ( .A(n11253), .B(n37934), .Z(n11096) );
  NANDN U12185 ( .A(n11094), .B(n37935), .Z(n11095) );
  NAND U12186 ( .A(n11096), .B(n11095), .Z(n11298) );
  XNOR U12187 ( .A(b[27]), .B(a[59]), .Z(n11256) );
  NANDN U12188 ( .A(n11256), .B(n38423), .Z(n11099) );
  NAND U12189 ( .A(n11097), .B(n38424), .Z(n11098) );
  NAND U12190 ( .A(n11099), .B(n11098), .Z(n11295) );
  XNOR U12191 ( .A(b[5]), .B(a[81]), .Z(n11259) );
  NANDN U12192 ( .A(n11259), .B(n36587), .Z(n11102) );
  NANDN U12193 ( .A(n11100), .B(n36588), .Z(n11101) );
  AND U12194 ( .A(n11102), .B(n11101), .Z(n11296) );
  XNOR U12195 ( .A(n11295), .B(n11296), .Z(n11297) );
  XNOR U12196 ( .A(n11298), .B(n11297), .Z(n11283) );
  NAND U12197 ( .A(n11103), .B(n37762), .Z(n11105) );
  XOR U12198 ( .A(b[17]), .B(a[69]), .Z(n11262) );
  NAND U12199 ( .A(n11262), .B(n37764), .Z(n11104) );
  NAND U12200 ( .A(n11105), .B(n11104), .Z(n11237) );
  XNOR U12201 ( .A(b[31]), .B(a[55]), .Z(n11265) );
  NANDN U12202 ( .A(n11265), .B(n38552), .Z(n11108) );
  NANDN U12203 ( .A(n11106), .B(n38553), .Z(n11107) );
  AND U12204 ( .A(n11108), .B(n11107), .Z(n11235) );
  OR U12205 ( .A(n11109), .B(n36105), .Z(n11111) );
  XOR U12206 ( .A(b[3]), .B(n15562), .Z(n11268) );
  NANDN U12207 ( .A(n11268), .B(n36107), .Z(n11110) );
  AND U12208 ( .A(n11111), .B(n11110), .Z(n11236) );
  XOR U12209 ( .A(n11237), .B(n11238), .Z(n11284) );
  XOR U12210 ( .A(n11283), .B(n11284), .Z(n11285) );
  XNOR U12211 ( .A(n11286), .B(n11285), .Z(n11332) );
  NANDN U12212 ( .A(n11113), .B(n11112), .Z(n11117) );
  NAND U12213 ( .A(n11115), .B(n11114), .Z(n11116) );
  NAND U12214 ( .A(n11117), .B(n11116), .Z(n11274) );
  NANDN U12215 ( .A(n11119), .B(n11118), .Z(n11123) );
  NAND U12216 ( .A(n11121), .B(n11120), .Z(n11122) );
  NAND U12217 ( .A(n11123), .B(n11122), .Z(n11272) );
  OR U12218 ( .A(n11125), .B(n11124), .Z(n11129) );
  NANDN U12219 ( .A(n11127), .B(n11126), .Z(n11128) );
  NAND U12220 ( .A(n11129), .B(n11128), .Z(n11271) );
  XNOR U12221 ( .A(n11274), .B(n11273), .Z(n11333) );
  XOR U12222 ( .A(n11332), .B(n11333), .Z(n11335) );
  NANDN U12223 ( .A(n11131), .B(n11130), .Z(n11135) );
  OR U12224 ( .A(n11133), .B(n11132), .Z(n11134) );
  NAND U12225 ( .A(n11135), .B(n11134), .Z(n11334) );
  XOR U12226 ( .A(n11335), .B(n11334), .Z(n11352) );
  OR U12227 ( .A(n11137), .B(n11136), .Z(n11141) );
  NAND U12228 ( .A(n11139), .B(n11138), .Z(n11140) );
  NAND U12229 ( .A(n11141), .B(n11140), .Z(n11351) );
  NANDN U12230 ( .A(n11143), .B(n11142), .Z(n11147) );
  NANDN U12231 ( .A(n11145), .B(n11144), .Z(n11146) );
  NAND U12232 ( .A(n11147), .B(n11146), .Z(n11340) );
  NANDN U12233 ( .A(n11153), .B(n11152), .Z(n11157) );
  NAND U12234 ( .A(n11155), .B(n11154), .Z(n11156) );
  NAND U12235 ( .A(n11157), .B(n11156), .Z(n11277) );
  NANDN U12236 ( .A(n11159), .B(n11158), .Z(n11163) );
  NAND U12237 ( .A(n11161), .B(n11160), .Z(n11162) );
  AND U12238 ( .A(n11163), .B(n11162), .Z(n11278) );
  XNOR U12239 ( .A(n11277), .B(n11278), .Z(n11279) );
  XNOR U12240 ( .A(b[9]), .B(a[77]), .Z(n11301) );
  NANDN U12241 ( .A(n11301), .B(n36925), .Z(n11166) );
  NANDN U12242 ( .A(n11164), .B(n36926), .Z(n11165) );
  NAND U12243 ( .A(n11166), .B(n11165), .Z(n11243) );
  XNOR U12244 ( .A(b[15]), .B(a[71]), .Z(n11304) );
  OR U12245 ( .A(n11304), .B(n37665), .Z(n11169) );
  NANDN U12246 ( .A(n11167), .B(n37604), .Z(n11168) );
  AND U12247 ( .A(n11169), .B(n11168), .Z(n11241) );
  XNOR U12248 ( .A(b[21]), .B(a[65]), .Z(n11307) );
  NANDN U12249 ( .A(n11307), .B(n38101), .Z(n11172) );
  NANDN U12250 ( .A(n11170), .B(n38102), .Z(n11171) );
  AND U12251 ( .A(n11172), .B(n11171), .Z(n11242) );
  XOR U12252 ( .A(n11243), .B(n11244), .Z(n11232) );
  XNOR U12253 ( .A(b[11]), .B(a[75]), .Z(n11310) );
  OR U12254 ( .A(n11310), .B(n37311), .Z(n11175) );
  NANDN U12255 ( .A(n11173), .B(n37218), .Z(n11174) );
  NAND U12256 ( .A(n11175), .B(n11174), .Z(n11230) );
  XOR U12257 ( .A(n1053), .B(a[73]), .Z(n11313) );
  NANDN U12258 ( .A(n11313), .B(n37424), .Z(n11178) );
  NANDN U12259 ( .A(n11176), .B(n37425), .Z(n11177) );
  NAND U12260 ( .A(n11178), .B(n11177), .Z(n11229) );
  XOR U12261 ( .A(n11232), .B(n11231), .Z(n11226) );
  NANDN U12262 ( .A(n1049), .B(a[85]), .Z(n11179) );
  XNOR U12263 ( .A(b[1]), .B(n11179), .Z(n11181) );
  NANDN U12264 ( .A(b[0]), .B(a[84]), .Z(n11180) );
  AND U12265 ( .A(n11181), .B(n11180), .Z(n11249) );
  NAND U12266 ( .A(n38490), .B(n11182), .Z(n11184) );
  XNOR U12267 ( .A(b[29]), .B(a[57]), .Z(n11320) );
  OR U12268 ( .A(n11320), .B(n1048), .Z(n11183) );
  NAND U12269 ( .A(n11184), .B(n11183), .Z(n11247) );
  NANDN U12270 ( .A(n1059), .B(a[53]), .Z(n11248) );
  XNOR U12271 ( .A(n11247), .B(n11248), .Z(n11250) );
  XNOR U12272 ( .A(n11249), .B(n11250), .Z(n11224) );
  NANDN U12273 ( .A(n11185), .B(n38205), .Z(n11187) );
  XNOR U12274 ( .A(b[23]), .B(a[63]), .Z(n11323) );
  OR U12275 ( .A(n11323), .B(n38268), .Z(n11186) );
  NAND U12276 ( .A(n11187), .B(n11186), .Z(n11292) );
  XOR U12277 ( .A(b[7]), .B(a[79]), .Z(n11326) );
  NAND U12278 ( .A(n11326), .B(n36701), .Z(n11190) );
  NAND U12279 ( .A(n11188), .B(n36702), .Z(n11189) );
  NAND U12280 ( .A(n11190), .B(n11189), .Z(n11289) );
  XOR U12281 ( .A(b[25]), .B(a[61]), .Z(n11329) );
  NAND U12282 ( .A(n11329), .B(n38325), .Z(n11193) );
  NAND U12283 ( .A(n11191), .B(n38326), .Z(n11192) );
  AND U12284 ( .A(n11193), .B(n11192), .Z(n11290) );
  XNOR U12285 ( .A(n11289), .B(n11290), .Z(n11291) );
  XOR U12286 ( .A(n11292), .B(n11291), .Z(n11223) );
  XOR U12287 ( .A(n11226), .B(n11225), .Z(n11280) );
  XNOR U12288 ( .A(n11279), .B(n11280), .Z(n11338) );
  XNOR U12289 ( .A(n11339), .B(n11338), .Z(n11341) );
  XNOR U12290 ( .A(n11340), .B(n11341), .Z(n11350) );
  XOR U12291 ( .A(n11351), .B(n11350), .Z(n11353) );
  NANDN U12292 ( .A(n11195), .B(n11194), .Z(n11199) );
  OR U12293 ( .A(n11197), .B(n11196), .Z(n11198) );
  NAND U12294 ( .A(n11199), .B(n11198), .Z(n11344) );
  NAND U12295 ( .A(n11201), .B(n11200), .Z(n11205) );
  NANDN U12296 ( .A(n11203), .B(n11202), .Z(n11204) );
  NAND U12297 ( .A(n11205), .B(n11204), .Z(n11345) );
  XNOR U12298 ( .A(n11344), .B(n11345), .Z(n11346) );
  XOR U12299 ( .A(n11347), .B(n11346), .Z(n11220) );
  XOR U12300 ( .A(n11219), .B(n11220), .Z(n11211) );
  XOR U12301 ( .A(n11212), .B(n11211), .Z(n11213) );
  XNOR U12302 ( .A(n11214), .B(n11213), .Z(n11356) );
  XNOR U12303 ( .A(n11356), .B(sreg[309]), .Z(n11358) );
  NAND U12304 ( .A(n11206), .B(sreg[308]), .Z(n11210) );
  OR U12305 ( .A(n11208), .B(n11207), .Z(n11209) );
  AND U12306 ( .A(n11210), .B(n11209), .Z(n11357) );
  XOR U12307 ( .A(n11358), .B(n11357), .Z(c[309]) );
  NAND U12308 ( .A(n11212), .B(n11211), .Z(n11216) );
  NAND U12309 ( .A(n11214), .B(n11213), .Z(n11215) );
  NAND U12310 ( .A(n11216), .B(n11215), .Z(n11364) );
  NANDN U12311 ( .A(n11218), .B(n11217), .Z(n11222) );
  NAND U12312 ( .A(n11220), .B(n11219), .Z(n11221) );
  NAND U12313 ( .A(n11222), .B(n11221), .Z(n11362) );
  NANDN U12314 ( .A(n11224), .B(n11223), .Z(n11228) );
  NANDN U12315 ( .A(n11226), .B(n11225), .Z(n11227) );
  NAND U12316 ( .A(n11228), .B(n11227), .Z(n11482) );
  OR U12317 ( .A(n11230), .B(n11229), .Z(n11234) );
  NAND U12318 ( .A(n11232), .B(n11231), .Z(n11233) );
  NAND U12319 ( .A(n11234), .B(n11233), .Z(n11421) );
  OR U12320 ( .A(n11236), .B(n11235), .Z(n11240) );
  NANDN U12321 ( .A(n11238), .B(n11237), .Z(n11239) );
  NAND U12322 ( .A(n11240), .B(n11239), .Z(n11420) );
  OR U12323 ( .A(n11242), .B(n11241), .Z(n11246) );
  NANDN U12324 ( .A(n11244), .B(n11243), .Z(n11245) );
  NAND U12325 ( .A(n11246), .B(n11245), .Z(n11419) );
  XOR U12326 ( .A(n11421), .B(n11422), .Z(n11479) );
  NANDN U12327 ( .A(n11248), .B(n11247), .Z(n11252) );
  NAND U12328 ( .A(n11250), .B(n11249), .Z(n11251) );
  NAND U12329 ( .A(n11252), .B(n11251), .Z(n11434) );
  XNOR U12330 ( .A(b[19]), .B(a[68]), .Z(n11401) );
  NANDN U12331 ( .A(n11401), .B(n37934), .Z(n11255) );
  NANDN U12332 ( .A(n11253), .B(n37935), .Z(n11254) );
  NAND U12333 ( .A(n11255), .B(n11254), .Z(n11446) );
  XOR U12334 ( .A(b[27]), .B(a[60]), .Z(n11404) );
  NAND U12335 ( .A(n38423), .B(n11404), .Z(n11258) );
  NANDN U12336 ( .A(n11256), .B(n38424), .Z(n11257) );
  NAND U12337 ( .A(n11258), .B(n11257), .Z(n11443) );
  XOR U12338 ( .A(b[5]), .B(n15424), .Z(n11407) );
  NANDN U12339 ( .A(n11407), .B(n36587), .Z(n11261) );
  NANDN U12340 ( .A(n11259), .B(n36588), .Z(n11260) );
  AND U12341 ( .A(n11261), .B(n11260), .Z(n11444) );
  XNOR U12342 ( .A(n11443), .B(n11444), .Z(n11445) );
  XNOR U12343 ( .A(n11446), .B(n11445), .Z(n11431) );
  NAND U12344 ( .A(n11262), .B(n37762), .Z(n11264) );
  XOR U12345 ( .A(b[17]), .B(a[70]), .Z(n11410) );
  NAND U12346 ( .A(n11410), .B(n37764), .Z(n11263) );
  NAND U12347 ( .A(n11264), .B(n11263), .Z(n11385) );
  XNOR U12348 ( .A(b[31]), .B(a[56]), .Z(n11413) );
  NANDN U12349 ( .A(n11413), .B(n38552), .Z(n11267) );
  NANDN U12350 ( .A(n11265), .B(n38553), .Z(n11266) );
  AND U12351 ( .A(n11267), .B(n11266), .Z(n11383) );
  OR U12352 ( .A(n11268), .B(n36105), .Z(n11270) );
  XNOR U12353 ( .A(b[3]), .B(a[84]), .Z(n11416) );
  NANDN U12354 ( .A(n11416), .B(n36107), .Z(n11269) );
  AND U12355 ( .A(n11270), .B(n11269), .Z(n11384) );
  XOR U12356 ( .A(n11385), .B(n11386), .Z(n11432) );
  XOR U12357 ( .A(n11431), .B(n11432), .Z(n11433) );
  XNOR U12358 ( .A(n11434), .B(n11433), .Z(n11480) );
  XNOR U12359 ( .A(n11479), .B(n11480), .Z(n11481) );
  XNOR U12360 ( .A(n11482), .B(n11481), .Z(n11500) );
  OR U12361 ( .A(n11272), .B(n11271), .Z(n11276) );
  NAND U12362 ( .A(n11274), .B(n11273), .Z(n11275) );
  NAND U12363 ( .A(n11276), .B(n11275), .Z(n11498) );
  NANDN U12364 ( .A(n11278), .B(n11277), .Z(n11282) );
  NANDN U12365 ( .A(n11280), .B(n11279), .Z(n11281) );
  NAND U12366 ( .A(n11282), .B(n11281), .Z(n11487) );
  OR U12367 ( .A(n11284), .B(n11283), .Z(n11288) );
  NAND U12368 ( .A(n11286), .B(n11285), .Z(n11287) );
  NAND U12369 ( .A(n11288), .B(n11287), .Z(n11486) );
  NANDN U12370 ( .A(n11290), .B(n11289), .Z(n11294) );
  NAND U12371 ( .A(n11292), .B(n11291), .Z(n11293) );
  NAND U12372 ( .A(n11294), .B(n11293), .Z(n11425) );
  NANDN U12373 ( .A(n11296), .B(n11295), .Z(n11300) );
  NAND U12374 ( .A(n11298), .B(n11297), .Z(n11299) );
  AND U12375 ( .A(n11300), .B(n11299), .Z(n11426) );
  XNOR U12376 ( .A(n11425), .B(n11426), .Z(n11427) );
  XNOR U12377 ( .A(n1052), .B(a[78]), .Z(n11455) );
  NAND U12378 ( .A(n36925), .B(n11455), .Z(n11303) );
  NANDN U12379 ( .A(n11301), .B(n36926), .Z(n11302) );
  NAND U12380 ( .A(n11303), .B(n11302), .Z(n11391) );
  XNOR U12381 ( .A(b[15]), .B(a[72]), .Z(n11452) );
  OR U12382 ( .A(n11452), .B(n37665), .Z(n11306) );
  NANDN U12383 ( .A(n11304), .B(n37604), .Z(n11305) );
  AND U12384 ( .A(n11306), .B(n11305), .Z(n11389) );
  XNOR U12385 ( .A(n1056), .B(a[66]), .Z(n11449) );
  NAND U12386 ( .A(n11449), .B(n38101), .Z(n11309) );
  NANDN U12387 ( .A(n11307), .B(n38102), .Z(n11308) );
  AND U12388 ( .A(n11309), .B(n11308), .Z(n11390) );
  XOR U12389 ( .A(n11391), .B(n11392), .Z(n11380) );
  XNOR U12390 ( .A(b[11]), .B(a[76]), .Z(n11458) );
  OR U12391 ( .A(n11458), .B(n37311), .Z(n11312) );
  NANDN U12392 ( .A(n11310), .B(n37218), .Z(n11311) );
  NAND U12393 ( .A(n11312), .B(n11311), .Z(n11378) );
  XOR U12394 ( .A(n1053), .B(a[74]), .Z(n11461) );
  NANDN U12395 ( .A(n11461), .B(n37424), .Z(n11315) );
  NANDN U12396 ( .A(n11313), .B(n37425), .Z(n11314) );
  NAND U12397 ( .A(n11315), .B(n11314), .Z(n11377) );
  XOR U12398 ( .A(n11380), .B(n11379), .Z(n11374) );
  NANDN U12399 ( .A(n1049), .B(a[86]), .Z(n11316) );
  XNOR U12400 ( .A(b[1]), .B(n11316), .Z(n11318) );
  NANDN U12401 ( .A(b[0]), .B(a[85]), .Z(n11317) );
  AND U12402 ( .A(n11318), .B(n11317), .Z(n11398) );
  ANDN U12403 ( .B(b[31]), .A(n11319), .Z(n11395) );
  NANDN U12404 ( .A(n11320), .B(n38490), .Z(n11322) );
  XNOR U12405 ( .A(n1058), .B(a[58]), .Z(n11464) );
  NANDN U12406 ( .A(n1048), .B(n11464), .Z(n11321) );
  NAND U12407 ( .A(n11322), .B(n11321), .Z(n11396) );
  XOR U12408 ( .A(n11395), .B(n11396), .Z(n11397) );
  XNOR U12409 ( .A(n11398), .B(n11397), .Z(n11371) );
  NANDN U12410 ( .A(n11323), .B(n38205), .Z(n11325) );
  XNOR U12411 ( .A(b[23]), .B(a[64]), .Z(n11470) );
  OR U12412 ( .A(n11470), .B(n38268), .Z(n11324) );
  NAND U12413 ( .A(n11325), .B(n11324), .Z(n11440) );
  XNOR U12414 ( .A(b[7]), .B(a[80]), .Z(n11473) );
  NANDN U12415 ( .A(n11473), .B(n36701), .Z(n11328) );
  NAND U12416 ( .A(n11326), .B(n36702), .Z(n11327) );
  NAND U12417 ( .A(n11328), .B(n11327), .Z(n11437) );
  XNOR U12418 ( .A(b[25]), .B(a[62]), .Z(n11476) );
  NANDN U12419 ( .A(n11476), .B(n38325), .Z(n11331) );
  NAND U12420 ( .A(n11329), .B(n38326), .Z(n11330) );
  AND U12421 ( .A(n11331), .B(n11330), .Z(n11438) );
  XNOR U12422 ( .A(n11437), .B(n11438), .Z(n11439) );
  XNOR U12423 ( .A(n11440), .B(n11439), .Z(n11372) );
  XOR U12424 ( .A(n11374), .B(n11373), .Z(n11428) );
  XNOR U12425 ( .A(n11427), .B(n11428), .Z(n11485) );
  XNOR U12426 ( .A(n11486), .B(n11485), .Z(n11488) );
  XNOR U12427 ( .A(n11487), .B(n11488), .Z(n11497) );
  XNOR U12428 ( .A(n11498), .B(n11497), .Z(n11499) );
  XOR U12429 ( .A(n11500), .B(n11499), .Z(n11494) );
  NANDN U12430 ( .A(n11333), .B(n11332), .Z(n11337) );
  OR U12431 ( .A(n11335), .B(n11334), .Z(n11336) );
  NAND U12432 ( .A(n11337), .B(n11336), .Z(n11491) );
  NAND U12433 ( .A(n11339), .B(n11338), .Z(n11343) );
  NANDN U12434 ( .A(n11341), .B(n11340), .Z(n11342) );
  NAND U12435 ( .A(n11343), .B(n11342), .Z(n11492) );
  XNOR U12436 ( .A(n11491), .B(n11492), .Z(n11493) );
  XNOR U12437 ( .A(n11494), .B(n11493), .Z(n11368) );
  NANDN U12438 ( .A(n11345), .B(n11344), .Z(n11349) );
  NAND U12439 ( .A(n11347), .B(n11346), .Z(n11348) );
  NAND U12440 ( .A(n11349), .B(n11348), .Z(n11365) );
  NANDN U12441 ( .A(n11351), .B(n11350), .Z(n11355) );
  OR U12442 ( .A(n11353), .B(n11352), .Z(n11354) );
  NAND U12443 ( .A(n11355), .B(n11354), .Z(n11366) );
  XNOR U12444 ( .A(n11365), .B(n11366), .Z(n11367) );
  XNOR U12445 ( .A(n11368), .B(n11367), .Z(n11361) );
  XOR U12446 ( .A(n11362), .B(n11361), .Z(n11363) );
  XNOR U12447 ( .A(n11364), .B(n11363), .Z(n11503) );
  XNOR U12448 ( .A(n11503), .B(sreg[310]), .Z(n11505) );
  NAND U12449 ( .A(n11356), .B(sreg[309]), .Z(n11360) );
  OR U12450 ( .A(n11358), .B(n11357), .Z(n11359) );
  AND U12451 ( .A(n11360), .B(n11359), .Z(n11504) );
  XOR U12452 ( .A(n11505), .B(n11504), .Z(c[310]) );
  NANDN U12453 ( .A(n11366), .B(n11365), .Z(n11370) );
  NANDN U12454 ( .A(n11368), .B(n11367), .Z(n11369) );
  NAND U12455 ( .A(n11370), .B(n11369), .Z(n11509) );
  OR U12456 ( .A(n11372), .B(n11371), .Z(n11376) );
  NANDN U12457 ( .A(n11374), .B(n11373), .Z(n11375) );
  NAND U12458 ( .A(n11376), .B(n11375), .Z(n11627) );
  OR U12459 ( .A(n11378), .B(n11377), .Z(n11382) );
  NAND U12460 ( .A(n11380), .B(n11379), .Z(n11381) );
  NAND U12461 ( .A(n11382), .B(n11381), .Z(n11566) );
  OR U12462 ( .A(n11384), .B(n11383), .Z(n11388) );
  NANDN U12463 ( .A(n11386), .B(n11385), .Z(n11387) );
  NAND U12464 ( .A(n11388), .B(n11387), .Z(n11565) );
  OR U12465 ( .A(n11390), .B(n11389), .Z(n11394) );
  NANDN U12466 ( .A(n11392), .B(n11391), .Z(n11393) );
  NAND U12467 ( .A(n11394), .B(n11393), .Z(n11564) );
  XOR U12468 ( .A(n11566), .B(n11567), .Z(n11625) );
  OR U12469 ( .A(n11396), .B(n11395), .Z(n11400) );
  NANDN U12470 ( .A(n11398), .B(n11397), .Z(n11399) );
  NAND U12471 ( .A(n11400), .B(n11399), .Z(n11578) );
  XNOR U12472 ( .A(b[19]), .B(a[69]), .Z(n11524) );
  NANDN U12473 ( .A(n11524), .B(n37934), .Z(n11403) );
  NANDN U12474 ( .A(n11401), .B(n37935), .Z(n11402) );
  NAND U12475 ( .A(n11403), .B(n11402), .Z(n11591) );
  XOR U12476 ( .A(b[27]), .B(a[61]), .Z(n11527) );
  NAND U12477 ( .A(n38423), .B(n11527), .Z(n11406) );
  NAND U12478 ( .A(n11404), .B(n38424), .Z(n11405) );
  NAND U12479 ( .A(n11406), .B(n11405), .Z(n11588) );
  XOR U12480 ( .A(b[5]), .B(n15562), .Z(n11530) );
  NANDN U12481 ( .A(n11530), .B(n36587), .Z(n11409) );
  NANDN U12482 ( .A(n11407), .B(n36588), .Z(n11408) );
  AND U12483 ( .A(n11409), .B(n11408), .Z(n11589) );
  XNOR U12484 ( .A(n11588), .B(n11589), .Z(n11590) );
  XNOR U12485 ( .A(n11591), .B(n11590), .Z(n11577) );
  NAND U12486 ( .A(n11410), .B(n37762), .Z(n11412) );
  XOR U12487 ( .A(b[17]), .B(a[71]), .Z(n11533) );
  NAND U12488 ( .A(n11533), .B(n37764), .Z(n11411) );
  NAND U12489 ( .A(n11412), .B(n11411), .Z(n11551) );
  XNOR U12490 ( .A(b[31]), .B(a[57]), .Z(n11536) );
  NANDN U12491 ( .A(n11536), .B(n38552), .Z(n11415) );
  NANDN U12492 ( .A(n11413), .B(n38553), .Z(n11414) );
  NAND U12493 ( .A(n11415), .B(n11414), .Z(n11548) );
  OR U12494 ( .A(n11416), .B(n36105), .Z(n11418) );
  XNOR U12495 ( .A(b[3]), .B(a[85]), .Z(n11539) );
  NANDN U12496 ( .A(n11539), .B(n36107), .Z(n11417) );
  AND U12497 ( .A(n11418), .B(n11417), .Z(n11549) );
  XNOR U12498 ( .A(n11548), .B(n11549), .Z(n11550) );
  XOR U12499 ( .A(n11551), .B(n11550), .Z(n11576) );
  XOR U12500 ( .A(n11577), .B(n11576), .Z(n11579) );
  XOR U12501 ( .A(n11578), .B(n11579), .Z(n11624) );
  XOR U12502 ( .A(n11625), .B(n11624), .Z(n11626) );
  XNOR U12503 ( .A(n11627), .B(n11626), .Z(n11645) );
  OR U12504 ( .A(n11420), .B(n11419), .Z(n11424) );
  NANDN U12505 ( .A(n11422), .B(n11421), .Z(n11423) );
  NAND U12506 ( .A(n11424), .B(n11423), .Z(n11643) );
  NANDN U12507 ( .A(n11426), .B(n11425), .Z(n11430) );
  NANDN U12508 ( .A(n11428), .B(n11427), .Z(n11429) );
  NAND U12509 ( .A(n11430), .B(n11429), .Z(n11632) );
  OR U12510 ( .A(n11432), .B(n11431), .Z(n11436) );
  NAND U12511 ( .A(n11434), .B(n11433), .Z(n11435) );
  NAND U12512 ( .A(n11436), .B(n11435), .Z(n11631) );
  NANDN U12513 ( .A(n11438), .B(n11437), .Z(n11442) );
  NAND U12514 ( .A(n11440), .B(n11439), .Z(n11441) );
  NAND U12515 ( .A(n11442), .B(n11441), .Z(n11570) );
  NANDN U12516 ( .A(n11444), .B(n11443), .Z(n11448) );
  NAND U12517 ( .A(n11446), .B(n11445), .Z(n11447) );
  AND U12518 ( .A(n11448), .B(n11447), .Z(n11571) );
  XNOR U12519 ( .A(n11570), .B(n11571), .Z(n11572) );
  XOR U12520 ( .A(b[21]), .B(n13219), .Z(n11600) );
  NANDN U12521 ( .A(n11600), .B(n38101), .Z(n11451) );
  NAND U12522 ( .A(n38102), .B(n11449), .Z(n11450) );
  NAND U12523 ( .A(n11451), .B(n11450), .Z(n11560) );
  XNOR U12524 ( .A(b[15]), .B(a[73]), .Z(n11597) );
  OR U12525 ( .A(n11597), .B(n37665), .Z(n11454) );
  NANDN U12526 ( .A(n11452), .B(n37604), .Z(n11453) );
  AND U12527 ( .A(n11454), .B(n11453), .Z(n11561) );
  XNOR U12528 ( .A(n11560), .B(n11561), .Z(n11563) );
  XNOR U12529 ( .A(b[9]), .B(a[79]), .Z(n11594) );
  NANDN U12530 ( .A(n11594), .B(n36925), .Z(n11457) );
  NAND U12531 ( .A(n36926), .B(n11455), .Z(n11456) );
  NAND U12532 ( .A(n11457), .B(n11456), .Z(n11562) );
  XNOR U12533 ( .A(n11563), .B(n11562), .Z(n11556) );
  XNOR U12534 ( .A(b[11]), .B(a[77]), .Z(n11603) );
  OR U12535 ( .A(n11603), .B(n37311), .Z(n11460) );
  NANDN U12536 ( .A(n11458), .B(n37218), .Z(n11459) );
  NAND U12537 ( .A(n11460), .B(n11459), .Z(n11555) );
  XOR U12538 ( .A(n1053), .B(a[75]), .Z(n11606) );
  NANDN U12539 ( .A(n11606), .B(n37424), .Z(n11463) );
  NANDN U12540 ( .A(n11461), .B(n37425), .Z(n11462) );
  NAND U12541 ( .A(n11463), .B(n11462), .Z(n11554) );
  XNOR U12542 ( .A(n11555), .B(n11554), .Z(n11557) );
  XNOR U12543 ( .A(n11556), .B(n11557), .Z(n11545) );
  NAND U12544 ( .A(n11464), .B(n38490), .Z(n11466) );
  XOR U12545 ( .A(n1058), .B(n12056), .Z(n11612) );
  NANDN U12546 ( .A(n1048), .B(n11612), .Z(n11465) );
  NAND U12547 ( .A(n11466), .B(n11465), .Z(n11518) );
  NANDN U12548 ( .A(n1059), .B(a[55]), .Z(n11519) );
  XNOR U12549 ( .A(n11518), .B(n11519), .Z(n11521) );
  NANDN U12550 ( .A(n1049), .B(a[87]), .Z(n11467) );
  XNOR U12551 ( .A(b[1]), .B(n11467), .Z(n11469) );
  NANDN U12552 ( .A(b[0]), .B(a[86]), .Z(n11468) );
  AND U12553 ( .A(n11469), .B(n11468), .Z(n11520) );
  XNOR U12554 ( .A(n11521), .B(n11520), .Z(n11543) );
  NANDN U12555 ( .A(n11470), .B(n38205), .Z(n11472) );
  XNOR U12556 ( .A(b[23]), .B(a[65]), .Z(n11615) );
  OR U12557 ( .A(n11615), .B(n38268), .Z(n11471) );
  NAND U12558 ( .A(n11472), .B(n11471), .Z(n11585) );
  XOR U12559 ( .A(b[7]), .B(a[81]), .Z(n11618) );
  NAND U12560 ( .A(n11618), .B(n36701), .Z(n11475) );
  NANDN U12561 ( .A(n11473), .B(n36702), .Z(n11474) );
  NAND U12562 ( .A(n11475), .B(n11474), .Z(n11582) );
  XOR U12563 ( .A(b[25]), .B(a[63]), .Z(n11621) );
  NAND U12564 ( .A(n11621), .B(n38325), .Z(n11478) );
  NANDN U12565 ( .A(n11476), .B(n38326), .Z(n11477) );
  AND U12566 ( .A(n11478), .B(n11477), .Z(n11583) );
  XNOR U12567 ( .A(n11582), .B(n11583), .Z(n11584) );
  XOR U12568 ( .A(n11585), .B(n11584), .Z(n11542) );
  XOR U12569 ( .A(n11545), .B(n11544), .Z(n11573) );
  XNOR U12570 ( .A(n11572), .B(n11573), .Z(n11630) );
  XNOR U12571 ( .A(n11631), .B(n11630), .Z(n11633) );
  XNOR U12572 ( .A(n11632), .B(n11633), .Z(n11642) );
  XNOR U12573 ( .A(n11643), .B(n11642), .Z(n11644) );
  XOR U12574 ( .A(n11645), .B(n11644), .Z(n11639) );
  NANDN U12575 ( .A(n11480), .B(n11479), .Z(n11484) );
  NAND U12576 ( .A(n11482), .B(n11481), .Z(n11483) );
  NAND U12577 ( .A(n11484), .B(n11483), .Z(n11637) );
  NAND U12578 ( .A(n11486), .B(n11485), .Z(n11490) );
  NANDN U12579 ( .A(n11488), .B(n11487), .Z(n11489) );
  AND U12580 ( .A(n11490), .B(n11489), .Z(n11636) );
  XNOR U12581 ( .A(n11637), .B(n11636), .Z(n11638) );
  XNOR U12582 ( .A(n11639), .B(n11638), .Z(n11515) );
  NANDN U12583 ( .A(n11492), .B(n11491), .Z(n11496) );
  NAND U12584 ( .A(n11494), .B(n11493), .Z(n11495) );
  NAND U12585 ( .A(n11496), .B(n11495), .Z(n11512) );
  NANDN U12586 ( .A(n11498), .B(n11497), .Z(n11502) );
  NANDN U12587 ( .A(n11500), .B(n11499), .Z(n11501) );
  NAND U12588 ( .A(n11502), .B(n11501), .Z(n11513) );
  XNOR U12589 ( .A(n11512), .B(n11513), .Z(n11514) );
  XNOR U12590 ( .A(n11515), .B(n11514), .Z(n11508) );
  XOR U12591 ( .A(n11509), .B(n11508), .Z(n11510) );
  XNOR U12592 ( .A(n11511), .B(n11510), .Z(n11648) );
  XNOR U12593 ( .A(n11648), .B(sreg[311]), .Z(n11650) );
  NAND U12594 ( .A(n11503), .B(sreg[310]), .Z(n11507) );
  OR U12595 ( .A(n11505), .B(n11504), .Z(n11506) );
  AND U12596 ( .A(n11507), .B(n11506), .Z(n11649) );
  XOR U12597 ( .A(n11650), .B(n11649), .Z(c[311]) );
  NANDN U12598 ( .A(n11513), .B(n11512), .Z(n11517) );
  NANDN U12599 ( .A(n11515), .B(n11514), .Z(n11516) );
  NAND U12600 ( .A(n11517), .B(n11516), .Z(n11654) );
  NANDN U12601 ( .A(n11519), .B(n11518), .Z(n11523) );
  NAND U12602 ( .A(n11521), .B(n11520), .Z(n11522) );
  NAND U12603 ( .A(n11523), .B(n11522), .Z(n11726) );
  XNOR U12604 ( .A(b[19]), .B(a[70]), .Z(n11671) );
  NANDN U12605 ( .A(n11671), .B(n37934), .Z(n11526) );
  NANDN U12606 ( .A(n11524), .B(n37935), .Z(n11525) );
  NAND U12607 ( .A(n11526), .B(n11525), .Z(n11736) );
  XNOR U12608 ( .A(b[27]), .B(a[62]), .Z(n11674) );
  NANDN U12609 ( .A(n11674), .B(n38423), .Z(n11529) );
  NAND U12610 ( .A(n11527), .B(n38424), .Z(n11528) );
  NAND U12611 ( .A(n11529), .B(n11528), .Z(n11733) );
  XNOR U12612 ( .A(b[5]), .B(a[84]), .Z(n11677) );
  NANDN U12613 ( .A(n11677), .B(n36587), .Z(n11532) );
  NANDN U12614 ( .A(n11530), .B(n36588), .Z(n11531) );
  AND U12615 ( .A(n11532), .B(n11531), .Z(n11734) );
  XNOR U12616 ( .A(n11733), .B(n11734), .Z(n11735) );
  XNOR U12617 ( .A(n11736), .B(n11735), .Z(n11724) );
  NAND U12618 ( .A(n11533), .B(n37762), .Z(n11535) );
  XOR U12619 ( .A(b[17]), .B(a[72]), .Z(n11680) );
  NAND U12620 ( .A(n11680), .B(n37764), .Z(n11534) );
  NAND U12621 ( .A(n11535), .B(n11534), .Z(n11698) );
  XNOR U12622 ( .A(b[31]), .B(a[58]), .Z(n11683) );
  NANDN U12623 ( .A(n11683), .B(n38552), .Z(n11538) );
  NANDN U12624 ( .A(n11536), .B(n38553), .Z(n11537) );
  NAND U12625 ( .A(n11538), .B(n11537), .Z(n11695) );
  OR U12626 ( .A(n11539), .B(n36105), .Z(n11541) );
  XNOR U12627 ( .A(b[3]), .B(a[86]), .Z(n11686) );
  NANDN U12628 ( .A(n11686), .B(n36107), .Z(n11540) );
  AND U12629 ( .A(n11541), .B(n11540), .Z(n11696) );
  XNOR U12630 ( .A(n11695), .B(n11696), .Z(n11697) );
  XOR U12631 ( .A(n11698), .B(n11697), .Z(n11723) );
  XNOR U12632 ( .A(n11724), .B(n11723), .Z(n11725) );
  XNOR U12633 ( .A(n11726), .B(n11725), .Z(n11775) );
  NANDN U12634 ( .A(n11543), .B(n11542), .Z(n11547) );
  NANDN U12635 ( .A(n11545), .B(n11544), .Z(n11546) );
  NAND U12636 ( .A(n11547), .B(n11546), .Z(n11776) );
  XNOR U12637 ( .A(n11775), .B(n11776), .Z(n11777) );
  NANDN U12638 ( .A(n11549), .B(n11548), .Z(n11553) );
  NAND U12639 ( .A(n11551), .B(n11550), .Z(n11552) );
  NAND U12640 ( .A(n11553), .B(n11552), .Z(n11716) );
  OR U12641 ( .A(n11555), .B(n11554), .Z(n11559) );
  NANDN U12642 ( .A(n11557), .B(n11556), .Z(n11558) );
  NAND U12643 ( .A(n11559), .B(n11558), .Z(n11714) );
  XNOR U12644 ( .A(n11714), .B(n11713), .Z(n11715) );
  XOR U12645 ( .A(n11716), .B(n11715), .Z(n11778) );
  XOR U12646 ( .A(n11777), .B(n11778), .Z(n11788) );
  OR U12647 ( .A(n11565), .B(n11564), .Z(n11569) );
  NANDN U12648 ( .A(n11567), .B(n11566), .Z(n11568) );
  NAND U12649 ( .A(n11569), .B(n11568), .Z(n11786) );
  NANDN U12650 ( .A(n11571), .B(n11570), .Z(n11575) );
  NANDN U12651 ( .A(n11573), .B(n11572), .Z(n11574) );
  NAND U12652 ( .A(n11575), .B(n11574), .Z(n11771) );
  NANDN U12653 ( .A(n11577), .B(n11576), .Z(n11581) );
  OR U12654 ( .A(n11579), .B(n11578), .Z(n11580) );
  NAND U12655 ( .A(n11581), .B(n11580), .Z(n11770) );
  NANDN U12656 ( .A(n11583), .B(n11582), .Z(n11587) );
  NAND U12657 ( .A(n11585), .B(n11584), .Z(n11586) );
  NAND U12658 ( .A(n11587), .B(n11586), .Z(n11717) );
  NANDN U12659 ( .A(n11589), .B(n11588), .Z(n11593) );
  NAND U12660 ( .A(n11591), .B(n11590), .Z(n11592) );
  AND U12661 ( .A(n11593), .B(n11592), .Z(n11718) );
  XNOR U12662 ( .A(n11717), .B(n11718), .Z(n11719) );
  XOR U12663 ( .A(b[9]), .B(n15068), .Z(n11739) );
  NANDN U12664 ( .A(n11739), .B(n36925), .Z(n11596) );
  NANDN U12665 ( .A(n11594), .B(n36926), .Z(n11595) );
  NAND U12666 ( .A(n11596), .B(n11595), .Z(n11703) );
  XNOR U12667 ( .A(b[15]), .B(a[74]), .Z(n11742) );
  OR U12668 ( .A(n11742), .B(n37665), .Z(n11599) );
  NANDN U12669 ( .A(n11597), .B(n37604), .Z(n11598) );
  AND U12670 ( .A(n11599), .B(n11598), .Z(n11701) );
  XNOR U12671 ( .A(b[21]), .B(a[68]), .Z(n11745) );
  NANDN U12672 ( .A(n11745), .B(n38101), .Z(n11602) );
  NANDN U12673 ( .A(n11600), .B(n38102), .Z(n11601) );
  AND U12674 ( .A(n11602), .B(n11601), .Z(n11702) );
  XOR U12675 ( .A(n11703), .B(n11704), .Z(n11692) );
  XNOR U12676 ( .A(b[11]), .B(a[78]), .Z(n11748) );
  OR U12677 ( .A(n11748), .B(n37311), .Z(n11605) );
  NANDN U12678 ( .A(n11603), .B(n37218), .Z(n11604) );
  NAND U12679 ( .A(n11605), .B(n11604), .Z(n11690) );
  XOR U12680 ( .A(n1053), .B(a[76]), .Z(n11751) );
  NANDN U12681 ( .A(n11751), .B(n37424), .Z(n11608) );
  NANDN U12682 ( .A(n11606), .B(n37425), .Z(n11607) );
  AND U12683 ( .A(n11608), .B(n11607), .Z(n11689) );
  XNOR U12684 ( .A(n11690), .B(n11689), .Z(n11691) );
  XOR U12685 ( .A(n11692), .B(n11691), .Z(n11709) );
  NANDN U12686 ( .A(n1049), .B(a[88]), .Z(n11609) );
  XNOR U12687 ( .A(b[1]), .B(n11609), .Z(n11611) );
  NANDN U12688 ( .A(b[0]), .B(a[87]), .Z(n11610) );
  AND U12689 ( .A(n11611), .B(n11610), .Z(n11667) );
  NAND U12690 ( .A(n38490), .B(n11612), .Z(n11614) );
  XNOR U12691 ( .A(n1058), .B(a[60]), .Z(n11757) );
  NANDN U12692 ( .A(n1048), .B(n11757), .Z(n11613) );
  NAND U12693 ( .A(n11614), .B(n11613), .Z(n11665) );
  NANDN U12694 ( .A(n1059), .B(a[56]), .Z(n11666) );
  XNOR U12695 ( .A(n11665), .B(n11666), .Z(n11668) );
  XOR U12696 ( .A(n11667), .B(n11668), .Z(n11707) );
  NANDN U12697 ( .A(n11615), .B(n38205), .Z(n11617) );
  XNOR U12698 ( .A(b[23]), .B(a[66]), .Z(n11760) );
  OR U12699 ( .A(n11760), .B(n38268), .Z(n11616) );
  NAND U12700 ( .A(n11617), .B(n11616), .Z(n11730) );
  XNOR U12701 ( .A(b[7]), .B(a[82]), .Z(n11763) );
  NANDN U12702 ( .A(n11763), .B(n36701), .Z(n11620) );
  NAND U12703 ( .A(n11618), .B(n36702), .Z(n11619) );
  NAND U12704 ( .A(n11620), .B(n11619), .Z(n11727) );
  XOR U12705 ( .A(b[25]), .B(a[64]), .Z(n11766) );
  NAND U12706 ( .A(n11766), .B(n38325), .Z(n11623) );
  NAND U12707 ( .A(n11621), .B(n38326), .Z(n11622) );
  AND U12708 ( .A(n11623), .B(n11622), .Z(n11728) );
  XNOR U12709 ( .A(n11727), .B(n11728), .Z(n11729) );
  XNOR U12710 ( .A(n11730), .B(n11729), .Z(n11708) );
  XOR U12711 ( .A(n11707), .B(n11708), .Z(n11710) );
  XNOR U12712 ( .A(n11709), .B(n11710), .Z(n11720) );
  XNOR U12713 ( .A(n11719), .B(n11720), .Z(n11769) );
  XNOR U12714 ( .A(n11770), .B(n11769), .Z(n11772) );
  XNOR U12715 ( .A(n11771), .B(n11772), .Z(n11785) );
  XOR U12716 ( .A(n11786), .B(n11785), .Z(n11787) );
  XNOR U12717 ( .A(n11788), .B(n11787), .Z(n11782) );
  NAND U12718 ( .A(n11625), .B(n11624), .Z(n11629) );
  NAND U12719 ( .A(n11627), .B(n11626), .Z(n11628) );
  NAND U12720 ( .A(n11629), .B(n11628), .Z(n11780) );
  NAND U12721 ( .A(n11631), .B(n11630), .Z(n11635) );
  NANDN U12722 ( .A(n11633), .B(n11632), .Z(n11634) );
  AND U12723 ( .A(n11635), .B(n11634), .Z(n11779) );
  XNOR U12724 ( .A(n11780), .B(n11779), .Z(n11781) );
  XOR U12725 ( .A(n11782), .B(n11781), .Z(n11661) );
  NANDN U12726 ( .A(n11637), .B(n11636), .Z(n11641) );
  NAND U12727 ( .A(n11639), .B(n11638), .Z(n11640) );
  NAND U12728 ( .A(n11641), .B(n11640), .Z(n11659) );
  NANDN U12729 ( .A(n11643), .B(n11642), .Z(n11647) );
  NANDN U12730 ( .A(n11645), .B(n11644), .Z(n11646) );
  NAND U12731 ( .A(n11647), .B(n11646), .Z(n11660) );
  XNOR U12732 ( .A(n11659), .B(n11660), .Z(n11662) );
  XOR U12733 ( .A(n11661), .B(n11662), .Z(n11653) );
  XOR U12734 ( .A(n11654), .B(n11653), .Z(n11655) );
  XNOR U12735 ( .A(n11656), .B(n11655), .Z(n11791) );
  XNOR U12736 ( .A(n11791), .B(sreg[312]), .Z(n11793) );
  NAND U12737 ( .A(n11648), .B(sreg[311]), .Z(n11652) );
  OR U12738 ( .A(n11650), .B(n11649), .Z(n11651) );
  AND U12739 ( .A(n11652), .B(n11651), .Z(n11792) );
  XOR U12740 ( .A(n11793), .B(n11792), .Z(c[312]) );
  NAND U12741 ( .A(n11654), .B(n11653), .Z(n11658) );
  NAND U12742 ( .A(n11656), .B(n11655), .Z(n11657) );
  NAND U12743 ( .A(n11658), .B(n11657), .Z(n11799) );
  NANDN U12744 ( .A(n11660), .B(n11659), .Z(n11664) );
  NAND U12745 ( .A(n11662), .B(n11661), .Z(n11663) );
  NAND U12746 ( .A(n11664), .B(n11663), .Z(n11797) );
  NANDN U12747 ( .A(n11666), .B(n11665), .Z(n11670) );
  NAND U12748 ( .A(n11668), .B(n11667), .Z(n11669) );
  NAND U12749 ( .A(n11670), .B(n11669), .Z(n11869) );
  XNOR U12750 ( .A(b[19]), .B(a[71]), .Z(n11836) );
  NANDN U12751 ( .A(n11836), .B(n37934), .Z(n11673) );
  NANDN U12752 ( .A(n11671), .B(n37935), .Z(n11672) );
  NAND U12753 ( .A(n11673), .B(n11672), .Z(n11881) );
  XOR U12754 ( .A(b[27]), .B(a[63]), .Z(n11839) );
  NAND U12755 ( .A(n38423), .B(n11839), .Z(n11676) );
  NANDN U12756 ( .A(n11674), .B(n38424), .Z(n11675) );
  NAND U12757 ( .A(n11676), .B(n11675), .Z(n11878) );
  XNOR U12758 ( .A(b[5]), .B(a[85]), .Z(n11842) );
  NANDN U12759 ( .A(n11842), .B(n36587), .Z(n11679) );
  NANDN U12760 ( .A(n11677), .B(n36588), .Z(n11678) );
  AND U12761 ( .A(n11679), .B(n11678), .Z(n11879) );
  XNOR U12762 ( .A(n11878), .B(n11879), .Z(n11880) );
  XNOR U12763 ( .A(n11881), .B(n11880), .Z(n11866) );
  NAND U12764 ( .A(n11680), .B(n37762), .Z(n11682) );
  XOR U12765 ( .A(b[17]), .B(a[73]), .Z(n11845) );
  NAND U12766 ( .A(n11845), .B(n37764), .Z(n11681) );
  NAND U12767 ( .A(n11682), .B(n11681), .Z(n11820) );
  XOR U12768 ( .A(b[31]), .B(n12056), .Z(n11848) );
  NANDN U12769 ( .A(n11848), .B(n38552), .Z(n11685) );
  NANDN U12770 ( .A(n11683), .B(n38553), .Z(n11684) );
  AND U12771 ( .A(n11685), .B(n11684), .Z(n11818) );
  OR U12772 ( .A(n11686), .B(n36105), .Z(n11688) );
  XNOR U12773 ( .A(b[3]), .B(a[87]), .Z(n11851) );
  NANDN U12774 ( .A(n11851), .B(n36107), .Z(n11687) );
  AND U12775 ( .A(n11688), .B(n11687), .Z(n11819) );
  XOR U12776 ( .A(n11820), .B(n11821), .Z(n11867) );
  XOR U12777 ( .A(n11866), .B(n11867), .Z(n11868) );
  XNOR U12778 ( .A(n11869), .B(n11868), .Z(n11914) );
  NANDN U12779 ( .A(n11690), .B(n11689), .Z(n11694) );
  NAND U12780 ( .A(n11692), .B(n11691), .Z(n11693) );
  NAND U12781 ( .A(n11694), .B(n11693), .Z(n11857) );
  NANDN U12782 ( .A(n11696), .B(n11695), .Z(n11700) );
  NAND U12783 ( .A(n11698), .B(n11697), .Z(n11699) );
  NAND U12784 ( .A(n11700), .B(n11699), .Z(n11855) );
  OR U12785 ( .A(n11702), .B(n11701), .Z(n11706) );
  NANDN U12786 ( .A(n11704), .B(n11703), .Z(n11705) );
  NAND U12787 ( .A(n11706), .B(n11705), .Z(n11854) );
  XNOR U12788 ( .A(n11857), .B(n11856), .Z(n11915) );
  XNOR U12789 ( .A(n11914), .B(n11915), .Z(n11916) );
  NANDN U12790 ( .A(n11708), .B(n11707), .Z(n11712) );
  OR U12791 ( .A(n11710), .B(n11709), .Z(n11711) );
  AND U12792 ( .A(n11712), .B(n11711), .Z(n11917) );
  XNOR U12793 ( .A(n11916), .B(n11917), .Z(n11929) );
  NANDN U12794 ( .A(n11718), .B(n11717), .Z(n11722) );
  NANDN U12795 ( .A(n11720), .B(n11719), .Z(n11721) );
  NAND U12796 ( .A(n11722), .B(n11721), .Z(n11923) );
  NANDN U12797 ( .A(n11728), .B(n11727), .Z(n11732) );
  NAND U12798 ( .A(n11730), .B(n11729), .Z(n11731) );
  NAND U12799 ( .A(n11732), .B(n11731), .Z(n11860) );
  NANDN U12800 ( .A(n11734), .B(n11733), .Z(n11738) );
  NAND U12801 ( .A(n11736), .B(n11735), .Z(n11737) );
  AND U12802 ( .A(n11738), .B(n11737), .Z(n11861) );
  XNOR U12803 ( .A(n11860), .B(n11861), .Z(n11862) );
  XNOR U12804 ( .A(b[9]), .B(a[81]), .Z(n11884) );
  NANDN U12805 ( .A(n11884), .B(n36925), .Z(n11741) );
  NANDN U12806 ( .A(n11739), .B(n36926), .Z(n11740) );
  NAND U12807 ( .A(n11741), .B(n11740), .Z(n11826) );
  XNOR U12808 ( .A(b[15]), .B(a[75]), .Z(n11887) );
  OR U12809 ( .A(n11887), .B(n37665), .Z(n11744) );
  NANDN U12810 ( .A(n11742), .B(n37604), .Z(n11743) );
  AND U12811 ( .A(n11744), .B(n11743), .Z(n11824) );
  XNOR U12812 ( .A(b[21]), .B(a[69]), .Z(n11890) );
  NANDN U12813 ( .A(n11890), .B(n38101), .Z(n11747) );
  NANDN U12814 ( .A(n11745), .B(n38102), .Z(n11746) );
  AND U12815 ( .A(n11747), .B(n11746), .Z(n11825) );
  XOR U12816 ( .A(n11826), .B(n11827), .Z(n11815) );
  XNOR U12817 ( .A(b[11]), .B(a[79]), .Z(n11893) );
  OR U12818 ( .A(n11893), .B(n37311), .Z(n11750) );
  NANDN U12819 ( .A(n11748), .B(n37218), .Z(n11749) );
  NAND U12820 ( .A(n11750), .B(n11749), .Z(n11813) );
  XOR U12821 ( .A(n1053), .B(a[77]), .Z(n11896) );
  NANDN U12822 ( .A(n11896), .B(n37424), .Z(n11753) );
  NANDN U12823 ( .A(n11751), .B(n37425), .Z(n11752) );
  NAND U12824 ( .A(n11753), .B(n11752), .Z(n11812) );
  XOR U12825 ( .A(n11815), .B(n11814), .Z(n11809) );
  NANDN U12826 ( .A(n1049), .B(a[89]), .Z(n11754) );
  XNOR U12827 ( .A(b[1]), .B(n11754), .Z(n11756) );
  NANDN U12828 ( .A(b[0]), .B(a[88]), .Z(n11755) );
  AND U12829 ( .A(n11756), .B(n11755), .Z(n11832) );
  NAND U12830 ( .A(n38490), .B(n11757), .Z(n11759) );
  XNOR U12831 ( .A(n1058), .B(a[61]), .Z(n11902) );
  NANDN U12832 ( .A(n1048), .B(n11902), .Z(n11758) );
  NAND U12833 ( .A(n11759), .B(n11758), .Z(n11830) );
  NANDN U12834 ( .A(n1059), .B(a[57]), .Z(n11831) );
  XNOR U12835 ( .A(n11830), .B(n11831), .Z(n11833) );
  XNOR U12836 ( .A(n11832), .B(n11833), .Z(n11807) );
  NANDN U12837 ( .A(n11760), .B(n38205), .Z(n11762) );
  XOR U12838 ( .A(b[23]), .B(n13219), .Z(n11905) );
  OR U12839 ( .A(n11905), .B(n38268), .Z(n11761) );
  NAND U12840 ( .A(n11762), .B(n11761), .Z(n11875) );
  XNOR U12841 ( .A(b[7]), .B(a[83]), .Z(n11908) );
  NANDN U12842 ( .A(n11908), .B(n36701), .Z(n11765) );
  NANDN U12843 ( .A(n11763), .B(n36702), .Z(n11764) );
  NAND U12844 ( .A(n11765), .B(n11764), .Z(n11872) );
  XOR U12845 ( .A(b[25]), .B(a[65]), .Z(n11911) );
  NAND U12846 ( .A(n11911), .B(n38325), .Z(n11768) );
  NAND U12847 ( .A(n11766), .B(n38326), .Z(n11767) );
  AND U12848 ( .A(n11768), .B(n11767), .Z(n11873) );
  XNOR U12849 ( .A(n11872), .B(n11873), .Z(n11874) );
  XOR U12850 ( .A(n11875), .B(n11874), .Z(n11806) );
  XOR U12851 ( .A(n11809), .B(n11808), .Z(n11863) );
  XNOR U12852 ( .A(n11862), .B(n11863), .Z(n11920) );
  XOR U12853 ( .A(n11921), .B(n11920), .Z(n11922) );
  XOR U12854 ( .A(n11923), .B(n11922), .Z(n11927) );
  XNOR U12855 ( .A(n11926), .B(n11927), .Z(n11928) );
  XNOR U12856 ( .A(n11929), .B(n11928), .Z(n11933) );
  NAND U12857 ( .A(n11770), .B(n11769), .Z(n11774) );
  NANDN U12858 ( .A(n11772), .B(n11771), .Z(n11773) );
  NAND U12859 ( .A(n11774), .B(n11773), .Z(n11930) );
  XNOR U12860 ( .A(n11930), .B(n11931), .Z(n11932) );
  XNOR U12861 ( .A(n11933), .B(n11932), .Z(n11803) );
  NANDN U12862 ( .A(n11780), .B(n11779), .Z(n11784) );
  NAND U12863 ( .A(n11782), .B(n11781), .Z(n11783) );
  NAND U12864 ( .A(n11784), .B(n11783), .Z(n11800) );
  NANDN U12865 ( .A(n11786), .B(n11785), .Z(n11790) );
  OR U12866 ( .A(n11788), .B(n11787), .Z(n11789) );
  NAND U12867 ( .A(n11790), .B(n11789), .Z(n11801) );
  XNOR U12868 ( .A(n11800), .B(n11801), .Z(n11802) );
  XNOR U12869 ( .A(n11803), .B(n11802), .Z(n11796) );
  XOR U12870 ( .A(n11797), .B(n11796), .Z(n11798) );
  XNOR U12871 ( .A(n11799), .B(n11798), .Z(n11936) );
  XNOR U12872 ( .A(n11936), .B(sreg[313]), .Z(n11938) );
  NAND U12873 ( .A(n11791), .B(sreg[312]), .Z(n11795) );
  OR U12874 ( .A(n11793), .B(n11792), .Z(n11794) );
  AND U12875 ( .A(n11795), .B(n11794), .Z(n11937) );
  XOR U12876 ( .A(n11938), .B(n11937), .Z(c[313]) );
  NANDN U12877 ( .A(n11801), .B(n11800), .Z(n11805) );
  NANDN U12878 ( .A(n11803), .B(n11802), .Z(n11804) );
  NAND U12879 ( .A(n11805), .B(n11804), .Z(n11942) );
  NANDN U12880 ( .A(n11807), .B(n11806), .Z(n11811) );
  NANDN U12881 ( .A(n11809), .B(n11808), .Z(n11810) );
  NAND U12882 ( .A(n11811), .B(n11810), .Z(n12075) );
  OR U12883 ( .A(n11813), .B(n11812), .Z(n11817) );
  NAND U12884 ( .A(n11815), .B(n11814), .Z(n11816) );
  NAND U12885 ( .A(n11817), .B(n11816), .Z(n12013) );
  OR U12886 ( .A(n11819), .B(n11818), .Z(n11823) );
  NANDN U12887 ( .A(n11821), .B(n11820), .Z(n11822) );
  NAND U12888 ( .A(n11823), .B(n11822), .Z(n12012) );
  OR U12889 ( .A(n11825), .B(n11824), .Z(n11829) );
  NANDN U12890 ( .A(n11827), .B(n11826), .Z(n11828) );
  NAND U12891 ( .A(n11829), .B(n11828), .Z(n12011) );
  XOR U12892 ( .A(n12013), .B(n12014), .Z(n12072) );
  NANDN U12893 ( .A(n11831), .B(n11830), .Z(n11835) );
  NAND U12894 ( .A(n11833), .B(n11832), .Z(n11834) );
  NAND U12895 ( .A(n11835), .B(n11834), .Z(n12026) );
  XNOR U12896 ( .A(b[19]), .B(a[72]), .Z(n11969) );
  NANDN U12897 ( .A(n11969), .B(n37934), .Z(n11838) );
  NANDN U12898 ( .A(n11836), .B(n37935), .Z(n11837) );
  NAND U12899 ( .A(n11838), .B(n11837), .Z(n12038) );
  XOR U12900 ( .A(b[27]), .B(a[64]), .Z(n11972) );
  NAND U12901 ( .A(n38423), .B(n11972), .Z(n11841) );
  NAND U12902 ( .A(n11839), .B(n38424), .Z(n11840) );
  NAND U12903 ( .A(n11841), .B(n11840), .Z(n12035) );
  XNOR U12904 ( .A(b[5]), .B(a[86]), .Z(n11975) );
  NANDN U12905 ( .A(n11975), .B(n36587), .Z(n11844) );
  NANDN U12906 ( .A(n11842), .B(n36588), .Z(n11843) );
  AND U12907 ( .A(n11844), .B(n11843), .Z(n12036) );
  XNOR U12908 ( .A(n12035), .B(n12036), .Z(n12037) );
  XNOR U12909 ( .A(n12038), .B(n12037), .Z(n12024) );
  NAND U12910 ( .A(n11845), .B(n37762), .Z(n11847) );
  XOR U12911 ( .A(b[17]), .B(a[74]), .Z(n11978) );
  NAND U12912 ( .A(n11978), .B(n37764), .Z(n11846) );
  NAND U12913 ( .A(n11847), .B(n11846), .Z(n11996) );
  XNOR U12914 ( .A(b[31]), .B(a[60]), .Z(n11981) );
  NANDN U12915 ( .A(n11981), .B(n38552), .Z(n11850) );
  NANDN U12916 ( .A(n11848), .B(n38553), .Z(n11849) );
  NAND U12917 ( .A(n11850), .B(n11849), .Z(n11993) );
  OR U12918 ( .A(n11851), .B(n36105), .Z(n11853) );
  XNOR U12919 ( .A(b[3]), .B(a[88]), .Z(n11984) );
  NANDN U12920 ( .A(n11984), .B(n36107), .Z(n11852) );
  AND U12921 ( .A(n11853), .B(n11852), .Z(n11994) );
  XNOR U12922 ( .A(n11993), .B(n11994), .Z(n11995) );
  XOR U12923 ( .A(n11996), .B(n11995), .Z(n12023) );
  XNOR U12924 ( .A(n12024), .B(n12023), .Z(n12025) );
  XNOR U12925 ( .A(n12026), .B(n12025), .Z(n12073) );
  XNOR U12926 ( .A(n12072), .B(n12073), .Z(n12074) );
  XNOR U12927 ( .A(n12075), .B(n12074), .Z(n11960) );
  OR U12928 ( .A(n11855), .B(n11854), .Z(n11859) );
  NAND U12929 ( .A(n11857), .B(n11856), .Z(n11858) );
  NAND U12930 ( .A(n11859), .B(n11858), .Z(n11958) );
  NANDN U12931 ( .A(n11861), .B(n11860), .Z(n11865) );
  NANDN U12932 ( .A(n11863), .B(n11862), .Z(n11864) );
  NAND U12933 ( .A(n11865), .B(n11864), .Z(n12080) );
  OR U12934 ( .A(n11867), .B(n11866), .Z(n11871) );
  NAND U12935 ( .A(n11869), .B(n11868), .Z(n11870) );
  NAND U12936 ( .A(n11871), .B(n11870), .Z(n12079) );
  NANDN U12937 ( .A(n11873), .B(n11872), .Z(n11877) );
  NAND U12938 ( .A(n11875), .B(n11874), .Z(n11876) );
  NAND U12939 ( .A(n11877), .B(n11876), .Z(n12017) );
  NANDN U12940 ( .A(n11879), .B(n11878), .Z(n11883) );
  NAND U12941 ( .A(n11881), .B(n11880), .Z(n11882) );
  AND U12942 ( .A(n11883), .B(n11882), .Z(n12018) );
  XNOR U12943 ( .A(n12017), .B(n12018), .Z(n12019) );
  XOR U12944 ( .A(b[9]), .B(n15424), .Z(n12041) );
  NANDN U12945 ( .A(n12041), .B(n36925), .Z(n11886) );
  NANDN U12946 ( .A(n11884), .B(n36926), .Z(n11885) );
  NAND U12947 ( .A(n11886), .B(n11885), .Z(n12001) );
  XNOR U12948 ( .A(b[15]), .B(a[76]), .Z(n12044) );
  OR U12949 ( .A(n12044), .B(n37665), .Z(n11889) );
  NANDN U12950 ( .A(n11887), .B(n37604), .Z(n11888) );
  AND U12951 ( .A(n11889), .B(n11888), .Z(n11999) );
  XNOR U12952 ( .A(b[21]), .B(a[70]), .Z(n12047) );
  NANDN U12953 ( .A(n12047), .B(n38101), .Z(n11892) );
  NANDN U12954 ( .A(n11890), .B(n38102), .Z(n11891) );
  AND U12955 ( .A(n11892), .B(n11891), .Z(n12000) );
  XOR U12956 ( .A(n12001), .B(n12002), .Z(n11990) );
  XOR U12957 ( .A(b[11]), .B(n15068), .Z(n12050) );
  OR U12958 ( .A(n12050), .B(n37311), .Z(n11895) );
  NANDN U12959 ( .A(n11893), .B(n37218), .Z(n11894) );
  NAND U12960 ( .A(n11895), .B(n11894), .Z(n11988) );
  XOR U12961 ( .A(n1053), .B(a[78]), .Z(n12053) );
  NANDN U12962 ( .A(n12053), .B(n37424), .Z(n11898) );
  NANDN U12963 ( .A(n11896), .B(n37425), .Z(n11897) );
  AND U12964 ( .A(n11898), .B(n11897), .Z(n11987) );
  XNOR U12965 ( .A(n11988), .B(n11987), .Z(n11989) );
  XOR U12966 ( .A(n11990), .B(n11989), .Z(n12007) );
  NANDN U12967 ( .A(n1049), .B(a[90]), .Z(n11899) );
  XNOR U12968 ( .A(b[1]), .B(n11899), .Z(n11901) );
  NANDN U12969 ( .A(b[0]), .B(a[89]), .Z(n11900) );
  AND U12970 ( .A(n11901), .B(n11900), .Z(n11965) );
  NAND U12971 ( .A(n38490), .B(n11902), .Z(n11904) );
  XOR U12972 ( .A(b[29]), .B(n12493), .Z(n12057) );
  OR U12973 ( .A(n12057), .B(n1048), .Z(n11903) );
  NAND U12974 ( .A(n11904), .B(n11903), .Z(n11963) );
  NANDN U12975 ( .A(n1059), .B(a[58]), .Z(n11964) );
  XNOR U12976 ( .A(n11963), .B(n11964), .Z(n11966) );
  XOR U12977 ( .A(n11965), .B(n11966), .Z(n12005) );
  NANDN U12978 ( .A(n11905), .B(n38205), .Z(n11907) );
  XNOR U12979 ( .A(b[23]), .B(a[68]), .Z(n12063) );
  OR U12980 ( .A(n12063), .B(n38268), .Z(n11906) );
  NAND U12981 ( .A(n11907), .B(n11906), .Z(n12032) );
  XOR U12982 ( .A(b[7]), .B(a[84]), .Z(n12066) );
  NAND U12983 ( .A(n12066), .B(n36701), .Z(n11910) );
  NANDN U12984 ( .A(n11908), .B(n36702), .Z(n11909) );
  NAND U12985 ( .A(n11910), .B(n11909), .Z(n12029) );
  XOR U12986 ( .A(b[25]), .B(a[66]), .Z(n12069) );
  NAND U12987 ( .A(n12069), .B(n38325), .Z(n11913) );
  NAND U12988 ( .A(n11911), .B(n38326), .Z(n11912) );
  AND U12989 ( .A(n11913), .B(n11912), .Z(n12030) );
  XNOR U12990 ( .A(n12029), .B(n12030), .Z(n12031) );
  XNOR U12991 ( .A(n12032), .B(n12031), .Z(n12006) );
  XOR U12992 ( .A(n12005), .B(n12006), .Z(n12008) );
  XNOR U12993 ( .A(n12007), .B(n12008), .Z(n12020) );
  XNOR U12994 ( .A(n12019), .B(n12020), .Z(n12078) );
  XNOR U12995 ( .A(n12079), .B(n12078), .Z(n12081) );
  XNOR U12996 ( .A(n12080), .B(n12081), .Z(n11957) );
  XNOR U12997 ( .A(n11958), .B(n11957), .Z(n11959) );
  XOR U12998 ( .A(n11960), .B(n11959), .Z(n11954) );
  NANDN U12999 ( .A(n11915), .B(n11914), .Z(n11919) );
  NAND U13000 ( .A(n11917), .B(n11916), .Z(n11918) );
  NAND U13001 ( .A(n11919), .B(n11918), .Z(n11951) );
  NAND U13002 ( .A(n11921), .B(n11920), .Z(n11925) );
  NAND U13003 ( .A(n11923), .B(n11922), .Z(n11924) );
  NAND U13004 ( .A(n11925), .B(n11924), .Z(n11952) );
  XNOR U13005 ( .A(n11951), .B(n11952), .Z(n11953) );
  XNOR U13006 ( .A(n11954), .B(n11953), .Z(n11948) );
  NANDN U13007 ( .A(n11931), .B(n11930), .Z(n11935) );
  NANDN U13008 ( .A(n11933), .B(n11932), .Z(n11934) );
  NAND U13009 ( .A(n11935), .B(n11934), .Z(n11946) );
  XNOR U13010 ( .A(n11945), .B(n11946), .Z(n11947) );
  XNOR U13011 ( .A(n11948), .B(n11947), .Z(n11941) );
  XOR U13012 ( .A(n11942), .B(n11941), .Z(n11943) );
  XNOR U13013 ( .A(n11944), .B(n11943), .Z(n12084) );
  XNOR U13014 ( .A(n12084), .B(sreg[314]), .Z(n12086) );
  NAND U13015 ( .A(n11936), .B(sreg[313]), .Z(n11940) );
  OR U13016 ( .A(n11938), .B(n11937), .Z(n11939) );
  AND U13017 ( .A(n11940), .B(n11939), .Z(n12085) );
  XOR U13018 ( .A(n12086), .B(n12085), .Z(c[314]) );
  NANDN U13019 ( .A(n11946), .B(n11945), .Z(n11950) );
  NANDN U13020 ( .A(n11948), .B(n11947), .Z(n11949) );
  NAND U13021 ( .A(n11950), .B(n11949), .Z(n12090) );
  NANDN U13022 ( .A(n11952), .B(n11951), .Z(n11956) );
  NAND U13023 ( .A(n11954), .B(n11953), .Z(n11955) );
  NAND U13024 ( .A(n11956), .B(n11955), .Z(n12095) );
  NANDN U13025 ( .A(n11958), .B(n11957), .Z(n11962) );
  NANDN U13026 ( .A(n11960), .B(n11959), .Z(n11961) );
  NAND U13027 ( .A(n11962), .B(n11961), .Z(n12096) );
  XNOR U13028 ( .A(n12095), .B(n12096), .Z(n12097) );
  NANDN U13029 ( .A(n11964), .B(n11963), .Z(n11968) );
  NAND U13030 ( .A(n11966), .B(n11965), .Z(n11967) );
  NAND U13031 ( .A(n11968), .B(n11967), .Z(n12164) );
  XNOR U13032 ( .A(b[19]), .B(a[73]), .Z(n12131) );
  NANDN U13033 ( .A(n12131), .B(n37934), .Z(n11971) );
  NANDN U13034 ( .A(n11969), .B(n37935), .Z(n11970) );
  NAND U13035 ( .A(n11971), .B(n11970), .Z(n12176) );
  XOR U13036 ( .A(b[27]), .B(a[65]), .Z(n12134) );
  NAND U13037 ( .A(n38423), .B(n12134), .Z(n11974) );
  NAND U13038 ( .A(n11972), .B(n38424), .Z(n11973) );
  NAND U13039 ( .A(n11974), .B(n11973), .Z(n12173) );
  XNOR U13040 ( .A(b[5]), .B(a[87]), .Z(n12137) );
  NANDN U13041 ( .A(n12137), .B(n36587), .Z(n11977) );
  NANDN U13042 ( .A(n11975), .B(n36588), .Z(n11976) );
  AND U13043 ( .A(n11977), .B(n11976), .Z(n12174) );
  XNOR U13044 ( .A(n12173), .B(n12174), .Z(n12175) );
  XNOR U13045 ( .A(n12176), .B(n12175), .Z(n12161) );
  NAND U13046 ( .A(n11978), .B(n37762), .Z(n11980) );
  XOR U13047 ( .A(b[17]), .B(a[75]), .Z(n12140) );
  NAND U13048 ( .A(n12140), .B(n37764), .Z(n11979) );
  NAND U13049 ( .A(n11980), .B(n11979), .Z(n12115) );
  XNOR U13050 ( .A(b[31]), .B(a[61]), .Z(n12143) );
  NANDN U13051 ( .A(n12143), .B(n38552), .Z(n11983) );
  NANDN U13052 ( .A(n11981), .B(n38553), .Z(n11982) );
  AND U13053 ( .A(n11983), .B(n11982), .Z(n12113) );
  OR U13054 ( .A(n11984), .B(n36105), .Z(n11986) );
  XNOR U13055 ( .A(b[3]), .B(a[89]), .Z(n12146) );
  NANDN U13056 ( .A(n12146), .B(n36107), .Z(n11985) );
  AND U13057 ( .A(n11986), .B(n11985), .Z(n12114) );
  XOR U13058 ( .A(n12115), .B(n12116), .Z(n12162) );
  XOR U13059 ( .A(n12161), .B(n12162), .Z(n12163) );
  XNOR U13060 ( .A(n12164), .B(n12163), .Z(n12209) );
  NANDN U13061 ( .A(n11988), .B(n11987), .Z(n11992) );
  NAND U13062 ( .A(n11990), .B(n11989), .Z(n11991) );
  NAND U13063 ( .A(n11992), .B(n11991), .Z(n12152) );
  NANDN U13064 ( .A(n11994), .B(n11993), .Z(n11998) );
  NAND U13065 ( .A(n11996), .B(n11995), .Z(n11997) );
  NAND U13066 ( .A(n11998), .B(n11997), .Z(n12150) );
  OR U13067 ( .A(n12000), .B(n11999), .Z(n12004) );
  NANDN U13068 ( .A(n12002), .B(n12001), .Z(n12003) );
  NAND U13069 ( .A(n12004), .B(n12003), .Z(n12149) );
  XNOR U13070 ( .A(n12152), .B(n12151), .Z(n12210) );
  XOR U13071 ( .A(n12209), .B(n12210), .Z(n12212) );
  NANDN U13072 ( .A(n12006), .B(n12005), .Z(n12010) );
  OR U13073 ( .A(n12008), .B(n12007), .Z(n12009) );
  NAND U13074 ( .A(n12010), .B(n12009), .Z(n12211) );
  XOR U13075 ( .A(n12212), .B(n12211), .Z(n12229) );
  OR U13076 ( .A(n12012), .B(n12011), .Z(n12016) );
  NANDN U13077 ( .A(n12014), .B(n12013), .Z(n12015) );
  NAND U13078 ( .A(n12016), .B(n12015), .Z(n12228) );
  NANDN U13079 ( .A(n12018), .B(n12017), .Z(n12022) );
  NANDN U13080 ( .A(n12020), .B(n12019), .Z(n12021) );
  NAND U13081 ( .A(n12022), .B(n12021), .Z(n12217) );
  NANDN U13082 ( .A(n12024), .B(n12023), .Z(n12028) );
  NAND U13083 ( .A(n12026), .B(n12025), .Z(n12027) );
  NAND U13084 ( .A(n12028), .B(n12027), .Z(n12216) );
  NANDN U13085 ( .A(n12030), .B(n12029), .Z(n12034) );
  NAND U13086 ( .A(n12032), .B(n12031), .Z(n12033) );
  NAND U13087 ( .A(n12034), .B(n12033), .Z(n12155) );
  NANDN U13088 ( .A(n12036), .B(n12035), .Z(n12040) );
  NAND U13089 ( .A(n12038), .B(n12037), .Z(n12039) );
  AND U13090 ( .A(n12040), .B(n12039), .Z(n12156) );
  XNOR U13091 ( .A(n12155), .B(n12156), .Z(n12157) );
  XOR U13092 ( .A(b[9]), .B(n15562), .Z(n12179) );
  NANDN U13093 ( .A(n12179), .B(n36925), .Z(n12043) );
  NANDN U13094 ( .A(n12041), .B(n36926), .Z(n12042) );
  NAND U13095 ( .A(n12043), .B(n12042), .Z(n12121) );
  XNOR U13096 ( .A(b[15]), .B(a[77]), .Z(n12182) );
  OR U13097 ( .A(n12182), .B(n37665), .Z(n12046) );
  NANDN U13098 ( .A(n12044), .B(n37604), .Z(n12045) );
  AND U13099 ( .A(n12046), .B(n12045), .Z(n12119) );
  XNOR U13100 ( .A(b[21]), .B(a[71]), .Z(n12185) );
  NANDN U13101 ( .A(n12185), .B(n38101), .Z(n12049) );
  NANDN U13102 ( .A(n12047), .B(n38102), .Z(n12048) );
  AND U13103 ( .A(n12049), .B(n12048), .Z(n12120) );
  XOR U13104 ( .A(n12121), .B(n12122), .Z(n12110) );
  XNOR U13105 ( .A(b[11]), .B(a[81]), .Z(n12188) );
  OR U13106 ( .A(n12188), .B(n37311), .Z(n12052) );
  NANDN U13107 ( .A(n12050), .B(n37218), .Z(n12051) );
  NAND U13108 ( .A(n12052), .B(n12051), .Z(n12108) );
  XOR U13109 ( .A(n1053), .B(a[79]), .Z(n12191) );
  NANDN U13110 ( .A(n12191), .B(n37424), .Z(n12055) );
  NANDN U13111 ( .A(n12053), .B(n37425), .Z(n12054) );
  NAND U13112 ( .A(n12055), .B(n12054), .Z(n12107) );
  XOR U13113 ( .A(n12110), .B(n12109), .Z(n12104) );
  ANDN U13114 ( .B(b[31]), .A(n12056), .Z(n12125) );
  NANDN U13115 ( .A(n12057), .B(n38490), .Z(n12059) );
  XNOR U13116 ( .A(n1058), .B(a[63]), .Z(n12197) );
  NANDN U13117 ( .A(n1048), .B(n12197), .Z(n12058) );
  NAND U13118 ( .A(n12059), .B(n12058), .Z(n12126) );
  XOR U13119 ( .A(n12125), .B(n12126), .Z(n12127) );
  NANDN U13120 ( .A(n1049), .B(a[91]), .Z(n12060) );
  XNOR U13121 ( .A(b[1]), .B(n12060), .Z(n12062) );
  NANDN U13122 ( .A(b[0]), .B(a[90]), .Z(n12061) );
  AND U13123 ( .A(n12062), .B(n12061), .Z(n12128) );
  XNOR U13124 ( .A(n12127), .B(n12128), .Z(n12101) );
  NANDN U13125 ( .A(n12063), .B(n38205), .Z(n12065) );
  XNOR U13126 ( .A(b[23]), .B(a[69]), .Z(n12200) );
  OR U13127 ( .A(n12200), .B(n38268), .Z(n12064) );
  NAND U13128 ( .A(n12065), .B(n12064), .Z(n12170) );
  XOR U13129 ( .A(b[7]), .B(a[85]), .Z(n12203) );
  NAND U13130 ( .A(n12203), .B(n36701), .Z(n12068) );
  NAND U13131 ( .A(n12066), .B(n36702), .Z(n12067) );
  NAND U13132 ( .A(n12068), .B(n12067), .Z(n12167) );
  XNOR U13133 ( .A(b[25]), .B(a[67]), .Z(n12206) );
  NANDN U13134 ( .A(n12206), .B(n38325), .Z(n12071) );
  NAND U13135 ( .A(n12069), .B(n38326), .Z(n12070) );
  AND U13136 ( .A(n12071), .B(n12070), .Z(n12168) );
  XNOR U13137 ( .A(n12167), .B(n12168), .Z(n12169) );
  XNOR U13138 ( .A(n12170), .B(n12169), .Z(n12102) );
  XOR U13139 ( .A(n12104), .B(n12103), .Z(n12158) );
  XNOR U13140 ( .A(n12157), .B(n12158), .Z(n12215) );
  XNOR U13141 ( .A(n12216), .B(n12215), .Z(n12218) );
  XNOR U13142 ( .A(n12217), .B(n12218), .Z(n12227) );
  XOR U13143 ( .A(n12228), .B(n12227), .Z(n12230) );
  NANDN U13144 ( .A(n12073), .B(n12072), .Z(n12077) );
  NAND U13145 ( .A(n12075), .B(n12074), .Z(n12076) );
  NAND U13146 ( .A(n12077), .B(n12076), .Z(n12222) );
  NAND U13147 ( .A(n12079), .B(n12078), .Z(n12083) );
  NANDN U13148 ( .A(n12081), .B(n12080), .Z(n12082) );
  AND U13149 ( .A(n12083), .B(n12082), .Z(n12221) );
  XNOR U13150 ( .A(n12222), .B(n12221), .Z(n12223) );
  XOR U13151 ( .A(n12224), .B(n12223), .Z(n12098) );
  XOR U13152 ( .A(n12097), .B(n12098), .Z(n12089) );
  XOR U13153 ( .A(n12090), .B(n12089), .Z(n12091) );
  XNOR U13154 ( .A(n12092), .B(n12091), .Z(n12233) );
  XNOR U13155 ( .A(n12233), .B(sreg[315]), .Z(n12235) );
  NAND U13156 ( .A(n12084), .B(sreg[314]), .Z(n12088) );
  OR U13157 ( .A(n12086), .B(n12085), .Z(n12087) );
  AND U13158 ( .A(n12088), .B(n12087), .Z(n12234) );
  XOR U13159 ( .A(n12235), .B(n12234), .Z(c[315]) );
  NAND U13160 ( .A(n12090), .B(n12089), .Z(n12094) );
  NAND U13161 ( .A(n12092), .B(n12091), .Z(n12093) );
  NAND U13162 ( .A(n12094), .B(n12093), .Z(n12241) );
  NANDN U13163 ( .A(n12096), .B(n12095), .Z(n12100) );
  NAND U13164 ( .A(n12098), .B(n12097), .Z(n12099) );
  NAND U13165 ( .A(n12100), .B(n12099), .Z(n12239) );
  OR U13166 ( .A(n12102), .B(n12101), .Z(n12106) );
  NANDN U13167 ( .A(n12104), .B(n12103), .Z(n12105) );
  NAND U13168 ( .A(n12106), .B(n12105), .Z(n12371) );
  OR U13169 ( .A(n12108), .B(n12107), .Z(n12112) );
  NAND U13170 ( .A(n12110), .B(n12109), .Z(n12111) );
  NAND U13171 ( .A(n12112), .B(n12111), .Z(n12310) );
  OR U13172 ( .A(n12114), .B(n12113), .Z(n12118) );
  NANDN U13173 ( .A(n12116), .B(n12115), .Z(n12117) );
  NAND U13174 ( .A(n12118), .B(n12117), .Z(n12309) );
  OR U13175 ( .A(n12120), .B(n12119), .Z(n12124) );
  NANDN U13176 ( .A(n12122), .B(n12121), .Z(n12123) );
  NAND U13177 ( .A(n12124), .B(n12123), .Z(n12308) );
  XOR U13178 ( .A(n12310), .B(n12311), .Z(n12369) );
  OR U13179 ( .A(n12126), .B(n12125), .Z(n12130) );
  NANDN U13180 ( .A(n12128), .B(n12127), .Z(n12129) );
  NAND U13181 ( .A(n12130), .B(n12129), .Z(n12322) );
  XNOR U13182 ( .A(b[19]), .B(a[74]), .Z(n12266) );
  NANDN U13183 ( .A(n12266), .B(n37934), .Z(n12133) );
  NANDN U13184 ( .A(n12131), .B(n37935), .Z(n12132) );
  NAND U13185 ( .A(n12133), .B(n12132), .Z(n12335) );
  XOR U13186 ( .A(b[27]), .B(a[66]), .Z(n12269) );
  NAND U13187 ( .A(n38423), .B(n12269), .Z(n12136) );
  NAND U13188 ( .A(n12134), .B(n38424), .Z(n12135) );
  NAND U13189 ( .A(n12136), .B(n12135), .Z(n12332) );
  XNOR U13190 ( .A(b[5]), .B(a[88]), .Z(n12272) );
  NANDN U13191 ( .A(n12272), .B(n36587), .Z(n12139) );
  NANDN U13192 ( .A(n12137), .B(n36588), .Z(n12138) );
  AND U13193 ( .A(n12139), .B(n12138), .Z(n12333) );
  XNOR U13194 ( .A(n12332), .B(n12333), .Z(n12334) );
  XNOR U13195 ( .A(n12335), .B(n12334), .Z(n12321) );
  NAND U13196 ( .A(n12140), .B(n37762), .Z(n12142) );
  XOR U13197 ( .A(b[17]), .B(a[76]), .Z(n12275) );
  NAND U13198 ( .A(n12275), .B(n37764), .Z(n12141) );
  NAND U13199 ( .A(n12142), .B(n12141), .Z(n12293) );
  XOR U13200 ( .A(b[31]), .B(n12493), .Z(n12278) );
  NANDN U13201 ( .A(n12278), .B(n38552), .Z(n12145) );
  NANDN U13202 ( .A(n12143), .B(n38553), .Z(n12144) );
  NAND U13203 ( .A(n12145), .B(n12144), .Z(n12290) );
  OR U13204 ( .A(n12146), .B(n36105), .Z(n12148) );
  XNOR U13205 ( .A(b[3]), .B(a[90]), .Z(n12281) );
  NANDN U13206 ( .A(n12281), .B(n36107), .Z(n12147) );
  AND U13207 ( .A(n12148), .B(n12147), .Z(n12291) );
  XNOR U13208 ( .A(n12290), .B(n12291), .Z(n12292) );
  XOR U13209 ( .A(n12293), .B(n12292), .Z(n12320) );
  XOR U13210 ( .A(n12321), .B(n12320), .Z(n12323) );
  XOR U13211 ( .A(n12322), .B(n12323), .Z(n12368) );
  XOR U13212 ( .A(n12369), .B(n12368), .Z(n12370) );
  XNOR U13213 ( .A(n12371), .B(n12370), .Z(n12257) );
  OR U13214 ( .A(n12150), .B(n12149), .Z(n12154) );
  NAND U13215 ( .A(n12152), .B(n12151), .Z(n12153) );
  NAND U13216 ( .A(n12154), .B(n12153), .Z(n12255) );
  NANDN U13217 ( .A(n12156), .B(n12155), .Z(n12160) );
  NANDN U13218 ( .A(n12158), .B(n12157), .Z(n12159) );
  NAND U13219 ( .A(n12160), .B(n12159), .Z(n12376) );
  OR U13220 ( .A(n12162), .B(n12161), .Z(n12166) );
  NAND U13221 ( .A(n12164), .B(n12163), .Z(n12165) );
  NAND U13222 ( .A(n12166), .B(n12165), .Z(n12375) );
  NANDN U13223 ( .A(n12168), .B(n12167), .Z(n12172) );
  NAND U13224 ( .A(n12170), .B(n12169), .Z(n12171) );
  NAND U13225 ( .A(n12172), .B(n12171), .Z(n12314) );
  NANDN U13226 ( .A(n12174), .B(n12173), .Z(n12178) );
  NAND U13227 ( .A(n12176), .B(n12175), .Z(n12177) );
  AND U13228 ( .A(n12178), .B(n12177), .Z(n12315) );
  XNOR U13229 ( .A(n12314), .B(n12315), .Z(n12316) );
  XNOR U13230 ( .A(b[9]), .B(a[84]), .Z(n12338) );
  NANDN U13231 ( .A(n12338), .B(n36925), .Z(n12181) );
  NANDN U13232 ( .A(n12179), .B(n36926), .Z(n12180) );
  NAND U13233 ( .A(n12181), .B(n12180), .Z(n12298) );
  XNOR U13234 ( .A(b[15]), .B(a[78]), .Z(n12341) );
  OR U13235 ( .A(n12341), .B(n37665), .Z(n12184) );
  NANDN U13236 ( .A(n12182), .B(n37604), .Z(n12183) );
  AND U13237 ( .A(n12184), .B(n12183), .Z(n12296) );
  XNOR U13238 ( .A(b[21]), .B(a[72]), .Z(n12344) );
  NANDN U13239 ( .A(n12344), .B(n38101), .Z(n12187) );
  NANDN U13240 ( .A(n12185), .B(n38102), .Z(n12186) );
  AND U13241 ( .A(n12187), .B(n12186), .Z(n12297) );
  XOR U13242 ( .A(n12298), .B(n12299), .Z(n12287) );
  XOR U13243 ( .A(b[11]), .B(n15424), .Z(n12347) );
  OR U13244 ( .A(n12347), .B(n37311), .Z(n12190) );
  NANDN U13245 ( .A(n12188), .B(n37218), .Z(n12189) );
  NAND U13246 ( .A(n12190), .B(n12189), .Z(n12285) );
  XOR U13247 ( .A(n1053), .B(a[80]), .Z(n12350) );
  NANDN U13248 ( .A(n12350), .B(n37424), .Z(n12193) );
  NANDN U13249 ( .A(n12191), .B(n37425), .Z(n12192) );
  AND U13250 ( .A(n12193), .B(n12192), .Z(n12284) );
  XNOR U13251 ( .A(n12285), .B(n12284), .Z(n12286) );
  XOR U13252 ( .A(n12287), .B(n12286), .Z(n12304) );
  NANDN U13253 ( .A(n1049), .B(a[92]), .Z(n12194) );
  XNOR U13254 ( .A(b[1]), .B(n12194), .Z(n12196) );
  NANDN U13255 ( .A(b[0]), .B(a[91]), .Z(n12195) );
  AND U13256 ( .A(n12196), .B(n12195), .Z(n12262) );
  NAND U13257 ( .A(n12197), .B(n38490), .Z(n12199) );
  XNOR U13258 ( .A(n1058), .B(a[64]), .Z(n12353) );
  NANDN U13259 ( .A(n1048), .B(n12353), .Z(n12198) );
  NAND U13260 ( .A(n12199), .B(n12198), .Z(n12260) );
  NANDN U13261 ( .A(n1059), .B(a[60]), .Z(n12261) );
  XNOR U13262 ( .A(n12260), .B(n12261), .Z(n12263) );
  XOR U13263 ( .A(n12262), .B(n12263), .Z(n12302) );
  NANDN U13264 ( .A(n12200), .B(n38205), .Z(n12202) );
  XNOR U13265 ( .A(b[23]), .B(a[70]), .Z(n12359) );
  OR U13266 ( .A(n12359), .B(n38268), .Z(n12201) );
  NAND U13267 ( .A(n12202), .B(n12201), .Z(n12329) );
  XOR U13268 ( .A(b[7]), .B(a[86]), .Z(n12362) );
  NAND U13269 ( .A(n12362), .B(n36701), .Z(n12205) );
  NAND U13270 ( .A(n12203), .B(n36702), .Z(n12204) );
  NAND U13271 ( .A(n12205), .B(n12204), .Z(n12326) );
  XOR U13272 ( .A(b[25]), .B(a[68]), .Z(n12365) );
  NAND U13273 ( .A(n12365), .B(n38325), .Z(n12208) );
  NANDN U13274 ( .A(n12206), .B(n38326), .Z(n12207) );
  AND U13275 ( .A(n12208), .B(n12207), .Z(n12327) );
  XNOR U13276 ( .A(n12326), .B(n12327), .Z(n12328) );
  XNOR U13277 ( .A(n12329), .B(n12328), .Z(n12303) );
  XOR U13278 ( .A(n12302), .B(n12303), .Z(n12305) );
  XNOR U13279 ( .A(n12304), .B(n12305), .Z(n12317) );
  XNOR U13280 ( .A(n12316), .B(n12317), .Z(n12374) );
  XNOR U13281 ( .A(n12375), .B(n12374), .Z(n12377) );
  XNOR U13282 ( .A(n12376), .B(n12377), .Z(n12254) );
  XNOR U13283 ( .A(n12255), .B(n12254), .Z(n12256) );
  XOR U13284 ( .A(n12257), .B(n12256), .Z(n12251) );
  NANDN U13285 ( .A(n12210), .B(n12209), .Z(n12214) );
  OR U13286 ( .A(n12212), .B(n12211), .Z(n12213) );
  NAND U13287 ( .A(n12214), .B(n12213), .Z(n12248) );
  NAND U13288 ( .A(n12216), .B(n12215), .Z(n12220) );
  NANDN U13289 ( .A(n12218), .B(n12217), .Z(n12219) );
  NAND U13290 ( .A(n12220), .B(n12219), .Z(n12249) );
  XNOR U13291 ( .A(n12248), .B(n12249), .Z(n12250) );
  XNOR U13292 ( .A(n12251), .B(n12250), .Z(n12245) );
  NANDN U13293 ( .A(n12222), .B(n12221), .Z(n12226) );
  NAND U13294 ( .A(n12224), .B(n12223), .Z(n12225) );
  NAND U13295 ( .A(n12226), .B(n12225), .Z(n12242) );
  NANDN U13296 ( .A(n12228), .B(n12227), .Z(n12232) );
  OR U13297 ( .A(n12230), .B(n12229), .Z(n12231) );
  NAND U13298 ( .A(n12232), .B(n12231), .Z(n12243) );
  XNOR U13299 ( .A(n12242), .B(n12243), .Z(n12244) );
  XNOR U13300 ( .A(n12245), .B(n12244), .Z(n12238) );
  XOR U13301 ( .A(n12239), .B(n12238), .Z(n12240) );
  XNOR U13302 ( .A(n12241), .B(n12240), .Z(n12380) );
  XNOR U13303 ( .A(n12380), .B(sreg[316]), .Z(n12382) );
  NAND U13304 ( .A(n12233), .B(sreg[315]), .Z(n12237) );
  OR U13305 ( .A(n12235), .B(n12234), .Z(n12236) );
  AND U13306 ( .A(n12237), .B(n12236), .Z(n12381) );
  XOR U13307 ( .A(n12382), .B(n12381), .Z(c[316]) );
  NANDN U13308 ( .A(n12243), .B(n12242), .Z(n12247) );
  NANDN U13309 ( .A(n12245), .B(n12244), .Z(n12246) );
  NAND U13310 ( .A(n12247), .B(n12246), .Z(n12386) );
  NANDN U13311 ( .A(n12249), .B(n12248), .Z(n12253) );
  NAND U13312 ( .A(n12251), .B(n12250), .Z(n12252) );
  NAND U13313 ( .A(n12253), .B(n12252), .Z(n12391) );
  NANDN U13314 ( .A(n12255), .B(n12254), .Z(n12259) );
  NANDN U13315 ( .A(n12257), .B(n12256), .Z(n12258) );
  NAND U13316 ( .A(n12259), .B(n12258), .Z(n12392) );
  XNOR U13317 ( .A(n12391), .B(n12392), .Z(n12393) );
  NANDN U13318 ( .A(n12261), .B(n12260), .Z(n12265) );
  NAND U13319 ( .A(n12263), .B(n12262), .Z(n12264) );
  NAND U13320 ( .A(n12265), .B(n12264), .Z(n12460) );
  XNOR U13321 ( .A(b[19]), .B(a[75]), .Z(n12427) );
  NANDN U13322 ( .A(n12427), .B(n37934), .Z(n12268) );
  NANDN U13323 ( .A(n12266), .B(n37935), .Z(n12267) );
  NAND U13324 ( .A(n12268), .B(n12267), .Z(n12472) );
  XNOR U13325 ( .A(b[27]), .B(a[67]), .Z(n12430) );
  NANDN U13326 ( .A(n12430), .B(n38423), .Z(n12271) );
  NAND U13327 ( .A(n12269), .B(n38424), .Z(n12270) );
  NAND U13328 ( .A(n12271), .B(n12270), .Z(n12469) );
  XNOR U13329 ( .A(b[5]), .B(a[89]), .Z(n12433) );
  NANDN U13330 ( .A(n12433), .B(n36587), .Z(n12274) );
  NANDN U13331 ( .A(n12272), .B(n36588), .Z(n12273) );
  AND U13332 ( .A(n12274), .B(n12273), .Z(n12470) );
  XNOR U13333 ( .A(n12469), .B(n12470), .Z(n12471) );
  XNOR U13334 ( .A(n12472), .B(n12471), .Z(n12457) );
  NAND U13335 ( .A(n12275), .B(n37762), .Z(n12277) );
  XOR U13336 ( .A(b[17]), .B(a[77]), .Z(n12436) );
  NAND U13337 ( .A(n12436), .B(n37764), .Z(n12276) );
  NAND U13338 ( .A(n12277), .B(n12276), .Z(n12411) );
  XNOR U13339 ( .A(b[31]), .B(a[63]), .Z(n12439) );
  NANDN U13340 ( .A(n12439), .B(n38552), .Z(n12280) );
  NANDN U13341 ( .A(n12278), .B(n38553), .Z(n12279) );
  AND U13342 ( .A(n12280), .B(n12279), .Z(n12409) );
  OR U13343 ( .A(n12281), .B(n36105), .Z(n12283) );
  XNOR U13344 ( .A(b[3]), .B(a[91]), .Z(n12442) );
  NANDN U13345 ( .A(n12442), .B(n36107), .Z(n12282) );
  AND U13346 ( .A(n12283), .B(n12282), .Z(n12410) );
  XOR U13347 ( .A(n12411), .B(n12412), .Z(n12458) );
  XOR U13348 ( .A(n12457), .B(n12458), .Z(n12459) );
  XNOR U13349 ( .A(n12460), .B(n12459), .Z(n12506) );
  NANDN U13350 ( .A(n12285), .B(n12284), .Z(n12289) );
  NAND U13351 ( .A(n12287), .B(n12286), .Z(n12288) );
  NAND U13352 ( .A(n12289), .B(n12288), .Z(n12448) );
  NANDN U13353 ( .A(n12291), .B(n12290), .Z(n12295) );
  NAND U13354 ( .A(n12293), .B(n12292), .Z(n12294) );
  NAND U13355 ( .A(n12295), .B(n12294), .Z(n12446) );
  OR U13356 ( .A(n12297), .B(n12296), .Z(n12301) );
  NANDN U13357 ( .A(n12299), .B(n12298), .Z(n12300) );
  NAND U13358 ( .A(n12301), .B(n12300), .Z(n12445) );
  XNOR U13359 ( .A(n12448), .B(n12447), .Z(n12507) );
  XOR U13360 ( .A(n12506), .B(n12507), .Z(n12509) );
  NANDN U13361 ( .A(n12303), .B(n12302), .Z(n12307) );
  OR U13362 ( .A(n12305), .B(n12304), .Z(n12306) );
  NAND U13363 ( .A(n12307), .B(n12306), .Z(n12508) );
  XOR U13364 ( .A(n12509), .B(n12508), .Z(n12526) );
  OR U13365 ( .A(n12309), .B(n12308), .Z(n12313) );
  NANDN U13366 ( .A(n12311), .B(n12310), .Z(n12312) );
  NAND U13367 ( .A(n12313), .B(n12312), .Z(n12525) );
  NANDN U13368 ( .A(n12315), .B(n12314), .Z(n12319) );
  NANDN U13369 ( .A(n12317), .B(n12316), .Z(n12318) );
  NAND U13370 ( .A(n12319), .B(n12318), .Z(n12514) );
  NANDN U13371 ( .A(n12321), .B(n12320), .Z(n12325) );
  OR U13372 ( .A(n12323), .B(n12322), .Z(n12324) );
  NAND U13373 ( .A(n12325), .B(n12324), .Z(n12513) );
  NANDN U13374 ( .A(n12327), .B(n12326), .Z(n12331) );
  NAND U13375 ( .A(n12329), .B(n12328), .Z(n12330) );
  NAND U13376 ( .A(n12331), .B(n12330), .Z(n12451) );
  NANDN U13377 ( .A(n12333), .B(n12332), .Z(n12337) );
  NAND U13378 ( .A(n12335), .B(n12334), .Z(n12336) );
  AND U13379 ( .A(n12337), .B(n12336), .Z(n12452) );
  XNOR U13380 ( .A(n12451), .B(n12452), .Z(n12453) );
  XNOR U13381 ( .A(n1052), .B(a[85]), .Z(n12481) );
  NAND U13382 ( .A(n36925), .B(n12481), .Z(n12340) );
  NANDN U13383 ( .A(n12338), .B(n36926), .Z(n12339) );
  NAND U13384 ( .A(n12340), .B(n12339), .Z(n12417) );
  XNOR U13385 ( .A(b[15]), .B(a[79]), .Z(n12478) );
  OR U13386 ( .A(n12478), .B(n37665), .Z(n12343) );
  NANDN U13387 ( .A(n12341), .B(n37604), .Z(n12342) );
  AND U13388 ( .A(n12343), .B(n12342), .Z(n12415) );
  XNOR U13389 ( .A(n1056), .B(a[73]), .Z(n12475) );
  NAND U13390 ( .A(n12475), .B(n38101), .Z(n12346) );
  NANDN U13391 ( .A(n12344), .B(n38102), .Z(n12345) );
  AND U13392 ( .A(n12346), .B(n12345), .Z(n12416) );
  XOR U13393 ( .A(n12417), .B(n12418), .Z(n12406) );
  XOR U13394 ( .A(b[11]), .B(n15562), .Z(n12484) );
  OR U13395 ( .A(n12484), .B(n37311), .Z(n12349) );
  NANDN U13396 ( .A(n12347), .B(n37218), .Z(n12348) );
  NAND U13397 ( .A(n12349), .B(n12348), .Z(n12404) );
  XOR U13398 ( .A(n1053), .B(a[81]), .Z(n12487) );
  NANDN U13399 ( .A(n12487), .B(n37424), .Z(n12352) );
  NANDN U13400 ( .A(n12350), .B(n37425), .Z(n12351) );
  NAND U13401 ( .A(n12352), .B(n12351), .Z(n12403) );
  XOR U13402 ( .A(n12406), .B(n12405), .Z(n12400) );
  NAND U13403 ( .A(n38490), .B(n12353), .Z(n12355) );
  XNOR U13404 ( .A(b[29]), .B(a[65]), .Z(n12494) );
  OR U13405 ( .A(n12494), .B(n1048), .Z(n12354) );
  NAND U13406 ( .A(n12355), .B(n12354), .Z(n12421) );
  NANDN U13407 ( .A(n1059), .B(a[61]), .Z(n12422) );
  XNOR U13408 ( .A(n12421), .B(n12422), .Z(n12424) );
  NANDN U13409 ( .A(n1049), .B(a[93]), .Z(n12356) );
  XNOR U13410 ( .A(b[1]), .B(n12356), .Z(n12358) );
  NANDN U13411 ( .A(b[0]), .B(a[92]), .Z(n12357) );
  AND U13412 ( .A(n12358), .B(n12357), .Z(n12423) );
  XNOR U13413 ( .A(n12424), .B(n12423), .Z(n12398) );
  NANDN U13414 ( .A(n12359), .B(n38205), .Z(n12361) );
  XNOR U13415 ( .A(b[23]), .B(a[71]), .Z(n12497) );
  OR U13416 ( .A(n12497), .B(n38268), .Z(n12360) );
  NAND U13417 ( .A(n12361), .B(n12360), .Z(n12466) );
  XOR U13418 ( .A(b[7]), .B(a[87]), .Z(n12500) );
  NAND U13419 ( .A(n12500), .B(n36701), .Z(n12364) );
  NAND U13420 ( .A(n12362), .B(n36702), .Z(n12363) );
  NAND U13421 ( .A(n12364), .B(n12363), .Z(n12463) );
  XOR U13422 ( .A(b[25]), .B(a[69]), .Z(n12503) );
  NAND U13423 ( .A(n12503), .B(n38325), .Z(n12367) );
  NAND U13424 ( .A(n12365), .B(n38326), .Z(n12366) );
  AND U13425 ( .A(n12367), .B(n12366), .Z(n12464) );
  XNOR U13426 ( .A(n12463), .B(n12464), .Z(n12465) );
  XOR U13427 ( .A(n12466), .B(n12465), .Z(n12397) );
  XOR U13428 ( .A(n12400), .B(n12399), .Z(n12454) );
  XNOR U13429 ( .A(n12453), .B(n12454), .Z(n12512) );
  XNOR U13430 ( .A(n12513), .B(n12512), .Z(n12515) );
  XNOR U13431 ( .A(n12514), .B(n12515), .Z(n12524) );
  XOR U13432 ( .A(n12525), .B(n12524), .Z(n12527) );
  NAND U13433 ( .A(n12369), .B(n12368), .Z(n12373) );
  NAND U13434 ( .A(n12371), .B(n12370), .Z(n12372) );
  NAND U13435 ( .A(n12373), .B(n12372), .Z(n12519) );
  NAND U13436 ( .A(n12375), .B(n12374), .Z(n12379) );
  NANDN U13437 ( .A(n12377), .B(n12376), .Z(n12378) );
  AND U13438 ( .A(n12379), .B(n12378), .Z(n12518) );
  XNOR U13439 ( .A(n12519), .B(n12518), .Z(n12520) );
  XOR U13440 ( .A(n12521), .B(n12520), .Z(n12394) );
  XOR U13441 ( .A(n12393), .B(n12394), .Z(n12385) );
  XOR U13442 ( .A(n12386), .B(n12385), .Z(n12387) );
  XNOR U13443 ( .A(n12388), .B(n12387), .Z(n12530) );
  XNOR U13444 ( .A(n12530), .B(sreg[317]), .Z(n12532) );
  NAND U13445 ( .A(n12380), .B(sreg[316]), .Z(n12384) );
  OR U13446 ( .A(n12382), .B(n12381), .Z(n12383) );
  AND U13447 ( .A(n12384), .B(n12383), .Z(n12531) );
  XOR U13448 ( .A(n12532), .B(n12531), .Z(c[317]) );
  NAND U13449 ( .A(n12386), .B(n12385), .Z(n12390) );
  NAND U13450 ( .A(n12388), .B(n12387), .Z(n12389) );
  NAND U13451 ( .A(n12390), .B(n12389), .Z(n12538) );
  NANDN U13452 ( .A(n12392), .B(n12391), .Z(n12396) );
  NAND U13453 ( .A(n12394), .B(n12393), .Z(n12395) );
  NAND U13454 ( .A(n12396), .B(n12395), .Z(n12536) );
  NANDN U13455 ( .A(n12398), .B(n12397), .Z(n12402) );
  NANDN U13456 ( .A(n12400), .B(n12399), .Z(n12401) );
  NAND U13457 ( .A(n12402), .B(n12401), .Z(n12654) );
  OR U13458 ( .A(n12404), .B(n12403), .Z(n12408) );
  NAND U13459 ( .A(n12406), .B(n12405), .Z(n12407) );
  NAND U13460 ( .A(n12408), .B(n12407), .Z(n12593) );
  OR U13461 ( .A(n12410), .B(n12409), .Z(n12414) );
  NANDN U13462 ( .A(n12412), .B(n12411), .Z(n12413) );
  NAND U13463 ( .A(n12414), .B(n12413), .Z(n12592) );
  OR U13464 ( .A(n12416), .B(n12415), .Z(n12420) );
  NANDN U13465 ( .A(n12418), .B(n12417), .Z(n12419) );
  NAND U13466 ( .A(n12420), .B(n12419), .Z(n12591) );
  XOR U13467 ( .A(n12593), .B(n12594), .Z(n12651) );
  NANDN U13468 ( .A(n12422), .B(n12421), .Z(n12426) );
  NAND U13469 ( .A(n12424), .B(n12423), .Z(n12425) );
  NAND U13470 ( .A(n12426), .B(n12425), .Z(n12606) );
  XNOR U13471 ( .A(b[19]), .B(a[76]), .Z(n12551) );
  NANDN U13472 ( .A(n12551), .B(n37934), .Z(n12429) );
  NANDN U13473 ( .A(n12427), .B(n37935), .Z(n12428) );
  NAND U13474 ( .A(n12429), .B(n12428), .Z(n12642) );
  XOR U13475 ( .A(b[27]), .B(a[68]), .Z(n12554) );
  NAND U13476 ( .A(n38423), .B(n12554), .Z(n12432) );
  NANDN U13477 ( .A(n12430), .B(n38424), .Z(n12431) );
  NAND U13478 ( .A(n12432), .B(n12431), .Z(n12639) );
  XNOR U13479 ( .A(b[5]), .B(a[90]), .Z(n12557) );
  NANDN U13480 ( .A(n12557), .B(n36587), .Z(n12435) );
  NANDN U13481 ( .A(n12433), .B(n36588), .Z(n12434) );
  AND U13482 ( .A(n12435), .B(n12434), .Z(n12640) );
  XNOR U13483 ( .A(n12639), .B(n12640), .Z(n12641) );
  XNOR U13484 ( .A(n12642), .B(n12641), .Z(n12604) );
  NAND U13485 ( .A(n12436), .B(n37762), .Z(n12438) );
  XOR U13486 ( .A(b[17]), .B(a[78]), .Z(n12560) );
  NAND U13487 ( .A(n12560), .B(n37764), .Z(n12437) );
  NAND U13488 ( .A(n12438), .B(n12437), .Z(n12578) );
  XNOR U13489 ( .A(b[31]), .B(a[64]), .Z(n12563) );
  NANDN U13490 ( .A(n12563), .B(n38552), .Z(n12441) );
  NANDN U13491 ( .A(n12439), .B(n38553), .Z(n12440) );
  NAND U13492 ( .A(n12441), .B(n12440), .Z(n12575) );
  OR U13493 ( .A(n12442), .B(n36105), .Z(n12444) );
  XNOR U13494 ( .A(b[3]), .B(a[92]), .Z(n12566) );
  NANDN U13495 ( .A(n12566), .B(n36107), .Z(n12443) );
  AND U13496 ( .A(n12444), .B(n12443), .Z(n12576) );
  XNOR U13497 ( .A(n12575), .B(n12576), .Z(n12577) );
  XOR U13498 ( .A(n12578), .B(n12577), .Z(n12603) );
  XNOR U13499 ( .A(n12604), .B(n12603), .Z(n12605) );
  XNOR U13500 ( .A(n12606), .B(n12605), .Z(n12652) );
  XNOR U13501 ( .A(n12651), .B(n12652), .Z(n12653) );
  XNOR U13502 ( .A(n12654), .B(n12653), .Z(n12672) );
  OR U13503 ( .A(n12446), .B(n12445), .Z(n12450) );
  NAND U13504 ( .A(n12448), .B(n12447), .Z(n12449) );
  NAND U13505 ( .A(n12450), .B(n12449), .Z(n12670) );
  NANDN U13506 ( .A(n12452), .B(n12451), .Z(n12456) );
  NANDN U13507 ( .A(n12454), .B(n12453), .Z(n12455) );
  NAND U13508 ( .A(n12456), .B(n12455), .Z(n12659) );
  OR U13509 ( .A(n12458), .B(n12457), .Z(n12462) );
  NAND U13510 ( .A(n12460), .B(n12459), .Z(n12461) );
  NAND U13511 ( .A(n12462), .B(n12461), .Z(n12658) );
  NANDN U13512 ( .A(n12464), .B(n12463), .Z(n12468) );
  NAND U13513 ( .A(n12466), .B(n12465), .Z(n12467) );
  NAND U13514 ( .A(n12468), .B(n12467), .Z(n12597) );
  NANDN U13515 ( .A(n12470), .B(n12469), .Z(n12474) );
  NAND U13516 ( .A(n12472), .B(n12471), .Z(n12473) );
  AND U13517 ( .A(n12474), .B(n12473), .Z(n12598) );
  XNOR U13518 ( .A(n12597), .B(n12598), .Z(n12599) );
  XOR U13519 ( .A(n1056), .B(a[74]), .Z(n12615) );
  NANDN U13520 ( .A(n12615), .B(n38101), .Z(n12477) );
  NAND U13521 ( .A(n38102), .B(n12475), .Z(n12476) );
  NAND U13522 ( .A(n12477), .B(n12476), .Z(n12587) );
  XOR U13523 ( .A(b[15]), .B(n15068), .Z(n12612) );
  OR U13524 ( .A(n12612), .B(n37665), .Z(n12480) );
  NANDN U13525 ( .A(n12478), .B(n37604), .Z(n12479) );
  AND U13526 ( .A(n12480), .B(n12479), .Z(n12588) );
  XNOR U13527 ( .A(n12587), .B(n12588), .Z(n12590) );
  XOR U13528 ( .A(n1052), .B(a[86]), .Z(n12609) );
  NANDN U13529 ( .A(n12609), .B(n36925), .Z(n12483) );
  NAND U13530 ( .A(n36926), .B(n12481), .Z(n12482) );
  NAND U13531 ( .A(n12483), .B(n12482), .Z(n12589) );
  XNOR U13532 ( .A(n12590), .B(n12589), .Z(n12583) );
  XNOR U13533 ( .A(b[11]), .B(a[84]), .Z(n12618) );
  OR U13534 ( .A(n12618), .B(n37311), .Z(n12486) );
  NANDN U13535 ( .A(n12484), .B(n37218), .Z(n12485) );
  NAND U13536 ( .A(n12486), .B(n12485), .Z(n12582) );
  XOR U13537 ( .A(n1053), .B(a[82]), .Z(n12621) );
  NANDN U13538 ( .A(n12621), .B(n37424), .Z(n12489) );
  NANDN U13539 ( .A(n12487), .B(n37425), .Z(n12488) );
  NAND U13540 ( .A(n12489), .B(n12488), .Z(n12581) );
  XNOR U13541 ( .A(n12582), .B(n12581), .Z(n12584) );
  XNOR U13542 ( .A(n12583), .B(n12584), .Z(n12572) );
  NANDN U13543 ( .A(n1049), .B(a[94]), .Z(n12490) );
  XNOR U13544 ( .A(b[1]), .B(n12490), .Z(n12492) );
  IV U13545 ( .A(a[93]), .Z(n17031) );
  NANDN U13546 ( .A(n17031), .B(n1049), .Z(n12491) );
  AND U13547 ( .A(n12492), .B(n12491), .Z(n12548) );
  ANDN U13548 ( .B(b[31]), .A(n12493), .Z(n12545) );
  NANDN U13549 ( .A(n12494), .B(n38490), .Z(n12496) );
  XNOR U13550 ( .A(n1058), .B(a[66]), .Z(n12624) );
  NANDN U13551 ( .A(n1048), .B(n12624), .Z(n12495) );
  NAND U13552 ( .A(n12496), .B(n12495), .Z(n12546) );
  XOR U13553 ( .A(n12545), .B(n12546), .Z(n12547) );
  XNOR U13554 ( .A(n12548), .B(n12547), .Z(n12569) );
  NANDN U13555 ( .A(n12497), .B(n38205), .Z(n12499) );
  XNOR U13556 ( .A(b[23]), .B(a[72]), .Z(n12630) );
  OR U13557 ( .A(n12630), .B(n38268), .Z(n12498) );
  NAND U13558 ( .A(n12499), .B(n12498), .Z(n12648) );
  XOR U13559 ( .A(b[7]), .B(a[88]), .Z(n12633) );
  NAND U13560 ( .A(n12633), .B(n36701), .Z(n12502) );
  NAND U13561 ( .A(n12500), .B(n36702), .Z(n12501) );
  NAND U13562 ( .A(n12502), .B(n12501), .Z(n12645) );
  XOR U13563 ( .A(b[25]), .B(a[70]), .Z(n12636) );
  NAND U13564 ( .A(n12636), .B(n38325), .Z(n12505) );
  NAND U13565 ( .A(n12503), .B(n38326), .Z(n12504) );
  AND U13566 ( .A(n12505), .B(n12504), .Z(n12646) );
  XNOR U13567 ( .A(n12645), .B(n12646), .Z(n12647) );
  XNOR U13568 ( .A(n12648), .B(n12647), .Z(n12570) );
  XOR U13569 ( .A(n12572), .B(n12571), .Z(n12600) );
  XNOR U13570 ( .A(n12599), .B(n12600), .Z(n12657) );
  XNOR U13571 ( .A(n12658), .B(n12657), .Z(n12660) );
  XNOR U13572 ( .A(n12659), .B(n12660), .Z(n12669) );
  XNOR U13573 ( .A(n12670), .B(n12669), .Z(n12671) );
  XOR U13574 ( .A(n12672), .B(n12671), .Z(n12666) );
  NANDN U13575 ( .A(n12507), .B(n12506), .Z(n12511) );
  OR U13576 ( .A(n12509), .B(n12508), .Z(n12510) );
  NAND U13577 ( .A(n12511), .B(n12510), .Z(n12663) );
  NAND U13578 ( .A(n12513), .B(n12512), .Z(n12517) );
  NANDN U13579 ( .A(n12515), .B(n12514), .Z(n12516) );
  NAND U13580 ( .A(n12517), .B(n12516), .Z(n12664) );
  XNOR U13581 ( .A(n12663), .B(n12664), .Z(n12665) );
  XNOR U13582 ( .A(n12666), .B(n12665), .Z(n12542) );
  NANDN U13583 ( .A(n12519), .B(n12518), .Z(n12523) );
  NAND U13584 ( .A(n12521), .B(n12520), .Z(n12522) );
  NAND U13585 ( .A(n12523), .B(n12522), .Z(n12539) );
  NANDN U13586 ( .A(n12525), .B(n12524), .Z(n12529) );
  OR U13587 ( .A(n12527), .B(n12526), .Z(n12528) );
  NAND U13588 ( .A(n12529), .B(n12528), .Z(n12540) );
  XNOR U13589 ( .A(n12539), .B(n12540), .Z(n12541) );
  XNOR U13590 ( .A(n12542), .B(n12541), .Z(n12535) );
  XOR U13591 ( .A(n12536), .B(n12535), .Z(n12537) );
  XNOR U13592 ( .A(n12538), .B(n12537), .Z(n12675) );
  XNOR U13593 ( .A(n12675), .B(sreg[318]), .Z(n12677) );
  NAND U13594 ( .A(n12530), .B(sreg[317]), .Z(n12534) );
  OR U13595 ( .A(n12532), .B(n12531), .Z(n12533) );
  AND U13596 ( .A(n12534), .B(n12533), .Z(n12676) );
  XOR U13597 ( .A(n12677), .B(n12676), .Z(c[318]) );
  NANDN U13598 ( .A(n12540), .B(n12539), .Z(n12544) );
  NANDN U13599 ( .A(n12542), .B(n12541), .Z(n12543) );
  NAND U13600 ( .A(n12544), .B(n12543), .Z(n12681) );
  OR U13601 ( .A(n12546), .B(n12545), .Z(n12550) );
  NANDN U13602 ( .A(n12548), .B(n12547), .Z(n12549) );
  NAND U13603 ( .A(n12550), .B(n12549), .Z(n12750) );
  XNOR U13604 ( .A(b[19]), .B(a[77]), .Z(n12698) );
  NANDN U13605 ( .A(n12698), .B(n37934), .Z(n12553) );
  NANDN U13606 ( .A(n12551), .B(n37935), .Z(n12552) );
  NAND U13607 ( .A(n12553), .B(n12552), .Z(n12763) );
  XOR U13608 ( .A(b[27]), .B(a[69]), .Z(n12701) );
  NAND U13609 ( .A(n38423), .B(n12701), .Z(n12556) );
  NAND U13610 ( .A(n12554), .B(n38424), .Z(n12555) );
  NAND U13611 ( .A(n12556), .B(n12555), .Z(n12760) );
  XNOR U13612 ( .A(b[5]), .B(a[91]), .Z(n12704) );
  NANDN U13613 ( .A(n12704), .B(n36587), .Z(n12559) );
  NANDN U13614 ( .A(n12557), .B(n36588), .Z(n12558) );
  AND U13615 ( .A(n12559), .B(n12558), .Z(n12761) );
  XNOR U13616 ( .A(n12760), .B(n12761), .Z(n12762) );
  XNOR U13617 ( .A(n12763), .B(n12762), .Z(n12749) );
  NAND U13618 ( .A(n12560), .B(n37762), .Z(n12562) );
  XOR U13619 ( .A(b[17]), .B(a[79]), .Z(n12707) );
  NAND U13620 ( .A(n12707), .B(n37764), .Z(n12561) );
  NAND U13621 ( .A(n12562), .B(n12561), .Z(n12725) );
  XNOR U13622 ( .A(b[31]), .B(a[65]), .Z(n12710) );
  NANDN U13623 ( .A(n12710), .B(n38552), .Z(n12565) );
  NANDN U13624 ( .A(n12563), .B(n38553), .Z(n12564) );
  NAND U13625 ( .A(n12565), .B(n12564), .Z(n12722) );
  OR U13626 ( .A(n12566), .B(n36105), .Z(n12568) );
  XOR U13627 ( .A(b[3]), .B(n17031), .Z(n12713) );
  NANDN U13628 ( .A(n12713), .B(n36107), .Z(n12567) );
  AND U13629 ( .A(n12568), .B(n12567), .Z(n12723) );
  XNOR U13630 ( .A(n12722), .B(n12723), .Z(n12724) );
  XOR U13631 ( .A(n12725), .B(n12724), .Z(n12748) );
  XOR U13632 ( .A(n12749), .B(n12748), .Z(n12751) );
  XNOR U13633 ( .A(n12750), .B(n12751), .Z(n12802) );
  OR U13634 ( .A(n12570), .B(n12569), .Z(n12574) );
  NANDN U13635 ( .A(n12572), .B(n12571), .Z(n12573) );
  NAND U13636 ( .A(n12574), .B(n12573), .Z(n12803) );
  XNOR U13637 ( .A(n12802), .B(n12803), .Z(n12804) );
  NANDN U13638 ( .A(n12576), .B(n12575), .Z(n12580) );
  NAND U13639 ( .A(n12578), .B(n12577), .Z(n12579) );
  NAND U13640 ( .A(n12580), .B(n12579), .Z(n12741) );
  OR U13641 ( .A(n12582), .B(n12581), .Z(n12586) );
  NANDN U13642 ( .A(n12584), .B(n12583), .Z(n12585) );
  NAND U13643 ( .A(n12586), .B(n12585), .Z(n12739) );
  XNOR U13644 ( .A(n12739), .B(n12738), .Z(n12740) );
  XOR U13645 ( .A(n12741), .B(n12740), .Z(n12805) );
  XOR U13646 ( .A(n12804), .B(n12805), .Z(n12817) );
  OR U13647 ( .A(n12592), .B(n12591), .Z(n12596) );
  NANDN U13648 ( .A(n12594), .B(n12593), .Z(n12595) );
  NAND U13649 ( .A(n12596), .B(n12595), .Z(n12815) );
  NANDN U13650 ( .A(n12598), .B(n12597), .Z(n12602) );
  NANDN U13651 ( .A(n12600), .B(n12599), .Z(n12601) );
  NAND U13652 ( .A(n12602), .B(n12601), .Z(n12799) );
  NANDN U13653 ( .A(n12604), .B(n12603), .Z(n12608) );
  NAND U13654 ( .A(n12606), .B(n12605), .Z(n12607) );
  NAND U13655 ( .A(n12608), .B(n12607), .Z(n12796) );
  XNOR U13656 ( .A(b[9]), .B(a[87]), .Z(n12766) );
  NANDN U13657 ( .A(n12766), .B(n36925), .Z(n12611) );
  NANDN U13658 ( .A(n12609), .B(n36926), .Z(n12610) );
  NAND U13659 ( .A(n12611), .B(n12610), .Z(n12730) );
  XNOR U13660 ( .A(n1054), .B(a[81]), .Z(n12769) );
  NANDN U13661 ( .A(n37665), .B(n12769), .Z(n12614) );
  NANDN U13662 ( .A(n12612), .B(n37604), .Z(n12613) );
  NAND U13663 ( .A(n12614), .B(n12613), .Z(n12728) );
  XNOR U13664 ( .A(b[21]), .B(a[75]), .Z(n12772) );
  NANDN U13665 ( .A(n12772), .B(n38101), .Z(n12617) );
  NANDN U13666 ( .A(n12615), .B(n38102), .Z(n12616) );
  NAND U13667 ( .A(n12617), .B(n12616), .Z(n12729) );
  XNOR U13668 ( .A(n12728), .B(n12729), .Z(n12731) );
  XOR U13669 ( .A(n12730), .B(n12731), .Z(n12719) );
  XNOR U13670 ( .A(b[11]), .B(a[85]), .Z(n12775) );
  OR U13671 ( .A(n12775), .B(n37311), .Z(n12620) );
  NANDN U13672 ( .A(n12618), .B(n37218), .Z(n12619) );
  NAND U13673 ( .A(n12620), .B(n12619), .Z(n12717) );
  XOR U13674 ( .A(n1053), .B(a[83]), .Z(n12778) );
  NANDN U13675 ( .A(n12778), .B(n37424), .Z(n12623) );
  NANDN U13676 ( .A(n12621), .B(n37425), .Z(n12622) );
  AND U13677 ( .A(n12623), .B(n12622), .Z(n12716) );
  XNOR U13678 ( .A(n12717), .B(n12716), .Z(n12718) );
  XNOR U13679 ( .A(n12719), .B(n12718), .Z(n12735) );
  NAND U13680 ( .A(n12624), .B(n38490), .Z(n12626) );
  XOR U13681 ( .A(n1058), .B(n13219), .Z(n12784) );
  NANDN U13682 ( .A(n1048), .B(n12784), .Z(n12625) );
  NAND U13683 ( .A(n12626), .B(n12625), .Z(n12692) );
  NANDN U13684 ( .A(n1059), .B(a[63]), .Z(n12693) );
  XNOR U13685 ( .A(n12692), .B(n12693), .Z(n12695) );
  NANDN U13686 ( .A(n1049), .B(a[95]), .Z(n12627) );
  XNOR U13687 ( .A(b[1]), .B(n12627), .Z(n12629) );
  NANDN U13688 ( .A(b[0]), .B(a[94]), .Z(n12628) );
  AND U13689 ( .A(n12629), .B(n12628), .Z(n12694) );
  XNOR U13690 ( .A(n12695), .B(n12694), .Z(n12733) );
  NANDN U13691 ( .A(n12630), .B(n38205), .Z(n12632) );
  XNOR U13692 ( .A(b[23]), .B(a[73]), .Z(n12787) );
  OR U13693 ( .A(n12787), .B(n38268), .Z(n12631) );
  NAND U13694 ( .A(n12632), .B(n12631), .Z(n12757) );
  XOR U13695 ( .A(b[7]), .B(a[89]), .Z(n12790) );
  NAND U13696 ( .A(n12790), .B(n36701), .Z(n12635) );
  NAND U13697 ( .A(n12633), .B(n36702), .Z(n12634) );
  NAND U13698 ( .A(n12635), .B(n12634), .Z(n12754) );
  XOR U13699 ( .A(b[25]), .B(a[71]), .Z(n12793) );
  NAND U13700 ( .A(n12793), .B(n38325), .Z(n12638) );
  NAND U13701 ( .A(n12636), .B(n38326), .Z(n12637) );
  AND U13702 ( .A(n12638), .B(n12637), .Z(n12755) );
  XNOR U13703 ( .A(n12754), .B(n12755), .Z(n12756) );
  XOR U13704 ( .A(n12757), .B(n12756), .Z(n12732) );
  XOR U13705 ( .A(n12735), .B(n12734), .Z(n12745) );
  NANDN U13706 ( .A(n12640), .B(n12639), .Z(n12644) );
  NAND U13707 ( .A(n12642), .B(n12641), .Z(n12643) );
  NAND U13708 ( .A(n12644), .B(n12643), .Z(n12743) );
  NANDN U13709 ( .A(n12646), .B(n12645), .Z(n12650) );
  NAND U13710 ( .A(n12648), .B(n12647), .Z(n12649) );
  AND U13711 ( .A(n12650), .B(n12649), .Z(n12742) );
  XNOR U13712 ( .A(n12743), .B(n12742), .Z(n12744) );
  XNOR U13713 ( .A(n12745), .B(n12744), .Z(n12797) );
  XNOR U13714 ( .A(n12796), .B(n12797), .Z(n12798) );
  XOR U13715 ( .A(n12799), .B(n12798), .Z(n12814) );
  XOR U13716 ( .A(n12815), .B(n12814), .Z(n12816) );
  XNOR U13717 ( .A(n12817), .B(n12816), .Z(n12811) );
  NANDN U13718 ( .A(n12652), .B(n12651), .Z(n12656) );
  NAND U13719 ( .A(n12654), .B(n12653), .Z(n12655) );
  NAND U13720 ( .A(n12656), .B(n12655), .Z(n12809) );
  NAND U13721 ( .A(n12658), .B(n12657), .Z(n12662) );
  NANDN U13722 ( .A(n12660), .B(n12659), .Z(n12661) );
  AND U13723 ( .A(n12662), .B(n12661), .Z(n12808) );
  XNOR U13724 ( .A(n12809), .B(n12808), .Z(n12810) );
  XOR U13725 ( .A(n12811), .B(n12810), .Z(n12688) );
  NANDN U13726 ( .A(n12664), .B(n12663), .Z(n12668) );
  NAND U13727 ( .A(n12666), .B(n12665), .Z(n12667) );
  NAND U13728 ( .A(n12668), .B(n12667), .Z(n12686) );
  NANDN U13729 ( .A(n12670), .B(n12669), .Z(n12674) );
  NANDN U13730 ( .A(n12672), .B(n12671), .Z(n12673) );
  NAND U13731 ( .A(n12674), .B(n12673), .Z(n12687) );
  XNOR U13732 ( .A(n12686), .B(n12687), .Z(n12689) );
  XOR U13733 ( .A(n12688), .B(n12689), .Z(n12680) );
  XOR U13734 ( .A(n12681), .B(n12680), .Z(n12682) );
  XNOR U13735 ( .A(n12683), .B(n12682), .Z(n12820) );
  XNOR U13736 ( .A(n12820), .B(sreg[319]), .Z(n12822) );
  NAND U13737 ( .A(n12675), .B(sreg[318]), .Z(n12679) );
  OR U13738 ( .A(n12677), .B(n12676), .Z(n12678) );
  AND U13739 ( .A(n12679), .B(n12678), .Z(n12821) );
  XOR U13740 ( .A(n12822), .B(n12821), .Z(c[319]) );
  NAND U13741 ( .A(n12681), .B(n12680), .Z(n12685) );
  NAND U13742 ( .A(n12683), .B(n12682), .Z(n12684) );
  NAND U13743 ( .A(n12685), .B(n12684), .Z(n12828) );
  NANDN U13744 ( .A(n12687), .B(n12686), .Z(n12691) );
  NAND U13745 ( .A(n12689), .B(n12688), .Z(n12690) );
  NAND U13746 ( .A(n12691), .B(n12690), .Z(n12826) );
  NANDN U13747 ( .A(n12693), .B(n12692), .Z(n12697) );
  NAND U13748 ( .A(n12695), .B(n12694), .Z(n12696) );
  NAND U13749 ( .A(n12697), .B(n12696), .Z(n12906) );
  XNOR U13750 ( .A(b[19]), .B(a[78]), .Z(n12851) );
  NANDN U13751 ( .A(n12851), .B(n37934), .Z(n12700) );
  NANDN U13752 ( .A(n12698), .B(n37935), .Z(n12699) );
  NAND U13753 ( .A(n12700), .B(n12699), .Z(n12916) );
  XOR U13754 ( .A(b[27]), .B(a[70]), .Z(n12854) );
  NAND U13755 ( .A(n38423), .B(n12854), .Z(n12703) );
  NAND U13756 ( .A(n12701), .B(n38424), .Z(n12702) );
  NAND U13757 ( .A(n12703), .B(n12702), .Z(n12913) );
  XNOR U13758 ( .A(b[5]), .B(a[92]), .Z(n12857) );
  NANDN U13759 ( .A(n12857), .B(n36587), .Z(n12706) );
  NANDN U13760 ( .A(n12704), .B(n36588), .Z(n12705) );
  AND U13761 ( .A(n12706), .B(n12705), .Z(n12914) );
  XNOR U13762 ( .A(n12913), .B(n12914), .Z(n12915) );
  XNOR U13763 ( .A(n12916), .B(n12915), .Z(n12904) );
  NAND U13764 ( .A(n12707), .B(n37762), .Z(n12709) );
  XNOR U13765 ( .A(b[17]), .B(a[80]), .Z(n12860) );
  NANDN U13766 ( .A(n12860), .B(n37764), .Z(n12708) );
  NAND U13767 ( .A(n12709), .B(n12708), .Z(n12878) );
  XNOR U13768 ( .A(b[31]), .B(a[66]), .Z(n12863) );
  NANDN U13769 ( .A(n12863), .B(n38552), .Z(n12712) );
  NANDN U13770 ( .A(n12710), .B(n38553), .Z(n12711) );
  NAND U13771 ( .A(n12712), .B(n12711), .Z(n12875) );
  OR U13772 ( .A(n12713), .B(n36105), .Z(n12715) );
  XNOR U13773 ( .A(b[3]), .B(a[94]), .Z(n12866) );
  NANDN U13774 ( .A(n12866), .B(n36107), .Z(n12714) );
  AND U13775 ( .A(n12715), .B(n12714), .Z(n12876) );
  XNOR U13776 ( .A(n12875), .B(n12876), .Z(n12877) );
  XOR U13777 ( .A(n12878), .B(n12877), .Z(n12903) );
  XNOR U13778 ( .A(n12904), .B(n12903), .Z(n12905) );
  XNOR U13779 ( .A(n12906), .B(n12905), .Z(n12842) );
  NANDN U13780 ( .A(n12717), .B(n12716), .Z(n12721) );
  NAND U13781 ( .A(n12719), .B(n12718), .Z(n12720) );
  NAND U13782 ( .A(n12721), .B(n12720), .Z(n12895) );
  NANDN U13783 ( .A(n12723), .B(n12722), .Z(n12727) );
  NAND U13784 ( .A(n12725), .B(n12724), .Z(n12726) );
  NAND U13785 ( .A(n12727), .B(n12726), .Z(n12894) );
  XNOR U13786 ( .A(n12894), .B(n12893), .Z(n12896) );
  XOR U13787 ( .A(n12895), .B(n12896), .Z(n12841) );
  XOR U13788 ( .A(n12842), .B(n12841), .Z(n12843) );
  NANDN U13789 ( .A(n12733), .B(n12732), .Z(n12737) );
  NAND U13790 ( .A(n12735), .B(n12734), .Z(n12736) );
  AND U13791 ( .A(n12737), .B(n12736), .Z(n12844) );
  XNOR U13792 ( .A(n12843), .B(n12844), .Z(n12952) );
  NANDN U13793 ( .A(n12743), .B(n12742), .Z(n12747) );
  NANDN U13794 ( .A(n12745), .B(n12744), .Z(n12746) );
  NAND U13795 ( .A(n12747), .B(n12746), .Z(n12838) );
  NANDN U13796 ( .A(n12749), .B(n12748), .Z(n12753) );
  OR U13797 ( .A(n12751), .B(n12750), .Z(n12752) );
  NAND U13798 ( .A(n12753), .B(n12752), .Z(n12836) );
  NANDN U13799 ( .A(n12755), .B(n12754), .Z(n12759) );
  NAND U13800 ( .A(n12757), .B(n12756), .Z(n12758) );
  NAND U13801 ( .A(n12759), .B(n12758), .Z(n12897) );
  NANDN U13802 ( .A(n12761), .B(n12760), .Z(n12765) );
  NAND U13803 ( .A(n12763), .B(n12762), .Z(n12764) );
  AND U13804 ( .A(n12765), .B(n12764), .Z(n12898) );
  XNOR U13805 ( .A(n12897), .B(n12898), .Z(n12899) );
  XNOR U13806 ( .A(b[9]), .B(a[88]), .Z(n12919) );
  NANDN U13807 ( .A(n12919), .B(n36925), .Z(n12768) );
  NANDN U13808 ( .A(n12766), .B(n36926), .Z(n12767) );
  NAND U13809 ( .A(n12768), .B(n12767), .Z(n12883) );
  XOR U13810 ( .A(b[15]), .B(n15424), .Z(n12922) );
  OR U13811 ( .A(n12922), .B(n37665), .Z(n12771) );
  NAND U13812 ( .A(n12769), .B(n37604), .Z(n12770) );
  AND U13813 ( .A(n12771), .B(n12770), .Z(n12881) );
  XNOR U13814 ( .A(b[21]), .B(a[76]), .Z(n12925) );
  NANDN U13815 ( .A(n12925), .B(n38101), .Z(n12774) );
  NANDN U13816 ( .A(n12772), .B(n38102), .Z(n12773) );
  AND U13817 ( .A(n12774), .B(n12773), .Z(n12882) );
  XOR U13818 ( .A(n12883), .B(n12884), .Z(n12872) );
  XNOR U13819 ( .A(b[11]), .B(a[86]), .Z(n12928) );
  OR U13820 ( .A(n12928), .B(n37311), .Z(n12777) );
  NANDN U13821 ( .A(n12775), .B(n37218), .Z(n12776) );
  NAND U13822 ( .A(n12777), .B(n12776), .Z(n12870) );
  XOR U13823 ( .A(n1053), .B(a[84]), .Z(n12931) );
  NANDN U13824 ( .A(n12931), .B(n37424), .Z(n12780) );
  NANDN U13825 ( .A(n12778), .B(n37425), .Z(n12779) );
  AND U13826 ( .A(n12780), .B(n12779), .Z(n12869) );
  XNOR U13827 ( .A(n12870), .B(n12869), .Z(n12871) );
  XOR U13828 ( .A(n12872), .B(n12871), .Z(n12889) );
  NANDN U13829 ( .A(n1049), .B(a[96]), .Z(n12781) );
  XNOR U13830 ( .A(b[1]), .B(n12781), .Z(n12783) );
  NANDN U13831 ( .A(b[0]), .B(a[95]), .Z(n12782) );
  AND U13832 ( .A(n12783), .B(n12782), .Z(n12847) );
  NAND U13833 ( .A(n38490), .B(n12784), .Z(n12786) );
  XNOR U13834 ( .A(n1058), .B(a[68]), .Z(n12937) );
  NANDN U13835 ( .A(n1048), .B(n12937), .Z(n12785) );
  NAND U13836 ( .A(n12786), .B(n12785), .Z(n12845) );
  NANDN U13837 ( .A(n1059), .B(a[64]), .Z(n12846) );
  XNOR U13838 ( .A(n12845), .B(n12846), .Z(n12848) );
  XOR U13839 ( .A(n12847), .B(n12848), .Z(n12887) );
  NANDN U13840 ( .A(n12787), .B(n38205), .Z(n12789) );
  XNOR U13841 ( .A(b[23]), .B(a[74]), .Z(n12940) );
  OR U13842 ( .A(n12940), .B(n38268), .Z(n12788) );
  NAND U13843 ( .A(n12789), .B(n12788), .Z(n12910) );
  XOR U13844 ( .A(b[7]), .B(a[90]), .Z(n12943) );
  NAND U13845 ( .A(n12943), .B(n36701), .Z(n12792) );
  NAND U13846 ( .A(n12790), .B(n36702), .Z(n12791) );
  NAND U13847 ( .A(n12792), .B(n12791), .Z(n12907) );
  XOR U13848 ( .A(b[25]), .B(a[72]), .Z(n12946) );
  NAND U13849 ( .A(n12946), .B(n38325), .Z(n12795) );
  NAND U13850 ( .A(n12793), .B(n38326), .Z(n12794) );
  AND U13851 ( .A(n12795), .B(n12794), .Z(n12908) );
  XNOR U13852 ( .A(n12907), .B(n12908), .Z(n12909) );
  XNOR U13853 ( .A(n12910), .B(n12909), .Z(n12888) );
  XOR U13854 ( .A(n12887), .B(n12888), .Z(n12890) );
  XNOR U13855 ( .A(n12889), .B(n12890), .Z(n12900) );
  XNOR U13856 ( .A(n12899), .B(n12900), .Z(n12835) );
  XNOR U13857 ( .A(n12836), .B(n12835), .Z(n12837) );
  XOR U13858 ( .A(n12838), .B(n12837), .Z(n12950) );
  XNOR U13859 ( .A(n12949), .B(n12950), .Z(n12951) );
  XNOR U13860 ( .A(n12952), .B(n12951), .Z(n12956) );
  NANDN U13861 ( .A(n12797), .B(n12796), .Z(n12801) );
  NAND U13862 ( .A(n12799), .B(n12798), .Z(n12800) );
  NAND U13863 ( .A(n12801), .B(n12800), .Z(n12953) );
  NANDN U13864 ( .A(n12803), .B(n12802), .Z(n12807) );
  NAND U13865 ( .A(n12805), .B(n12804), .Z(n12806) );
  NAND U13866 ( .A(n12807), .B(n12806), .Z(n12954) );
  XNOR U13867 ( .A(n12953), .B(n12954), .Z(n12955) );
  XNOR U13868 ( .A(n12956), .B(n12955), .Z(n12832) );
  NANDN U13869 ( .A(n12809), .B(n12808), .Z(n12813) );
  NAND U13870 ( .A(n12811), .B(n12810), .Z(n12812) );
  NAND U13871 ( .A(n12813), .B(n12812), .Z(n12829) );
  NANDN U13872 ( .A(n12815), .B(n12814), .Z(n12819) );
  OR U13873 ( .A(n12817), .B(n12816), .Z(n12818) );
  NAND U13874 ( .A(n12819), .B(n12818), .Z(n12830) );
  XNOR U13875 ( .A(n12829), .B(n12830), .Z(n12831) );
  XNOR U13876 ( .A(n12832), .B(n12831), .Z(n12825) );
  XOR U13877 ( .A(n12826), .B(n12825), .Z(n12827) );
  XNOR U13878 ( .A(n12828), .B(n12827), .Z(n12959) );
  XNOR U13879 ( .A(n12959), .B(sreg[320]), .Z(n12961) );
  NAND U13880 ( .A(n12820), .B(sreg[319]), .Z(n12824) );
  OR U13881 ( .A(n12822), .B(n12821), .Z(n12823) );
  AND U13882 ( .A(n12824), .B(n12823), .Z(n12960) );
  XOR U13883 ( .A(n12961), .B(n12960), .Z(c[320]) );
  NANDN U13884 ( .A(n12830), .B(n12829), .Z(n12834) );
  NANDN U13885 ( .A(n12832), .B(n12831), .Z(n12833) );
  NAND U13886 ( .A(n12834), .B(n12833), .Z(n12964) );
  NAND U13887 ( .A(n12836), .B(n12835), .Z(n12840) );
  OR U13888 ( .A(n12838), .B(n12837), .Z(n12839) );
  NAND U13889 ( .A(n12840), .B(n12839), .Z(n13096) );
  XNOR U13890 ( .A(n13096), .B(n13097), .Z(n13098) );
  NANDN U13891 ( .A(n12846), .B(n12845), .Z(n12850) );
  NAND U13892 ( .A(n12848), .B(n12847), .Z(n12849) );
  NAND U13893 ( .A(n12850), .B(n12849), .Z(n13039) );
  XNOR U13894 ( .A(b[19]), .B(a[79]), .Z(n13006) );
  NANDN U13895 ( .A(n13006), .B(n37934), .Z(n12853) );
  NANDN U13896 ( .A(n12851), .B(n37935), .Z(n12852) );
  NAND U13897 ( .A(n12853), .B(n12852), .Z(n13051) );
  XOR U13898 ( .A(b[27]), .B(a[71]), .Z(n13009) );
  NAND U13899 ( .A(n38423), .B(n13009), .Z(n12856) );
  NAND U13900 ( .A(n12854), .B(n38424), .Z(n12855) );
  NAND U13901 ( .A(n12856), .B(n12855), .Z(n13048) );
  XOR U13902 ( .A(b[5]), .B(n17031), .Z(n13012) );
  NANDN U13903 ( .A(n13012), .B(n36587), .Z(n12859) );
  NANDN U13904 ( .A(n12857), .B(n36588), .Z(n12858) );
  AND U13905 ( .A(n12859), .B(n12858), .Z(n13049) );
  XNOR U13906 ( .A(n13048), .B(n13049), .Z(n13050) );
  XNOR U13907 ( .A(n13051), .B(n13050), .Z(n13036) );
  NANDN U13908 ( .A(n12860), .B(n37762), .Z(n12862) );
  XOR U13909 ( .A(b[17]), .B(a[81]), .Z(n13015) );
  NAND U13910 ( .A(n13015), .B(n37764), .Z(n12861) );
  NAND U13911 ( .A(n12862), .B(n12861), .Z(n12990) );
  XOR U13912 ( .A(b[31]), .B(n13219), .Z(n13018) );
  NANDN U13913 ( .A(n13018), .B(n38552), .Z(n12865) );
  NANDN U13914 ( .A(n12863), .B(n38553), .Z(n12864) );
  AND U13915 ( .A(n12865), .B(n12864), .Z(n12988) );
  OR U13916 ( .A(n12866), .B(n36105), .Z(n12868) );
  XNOR U13917 ( .A(b[3]), .B(a[95]), .Z(n13021) );
  NANDN U13918 ( .A(n13021), .B(n36107), .Z(n12867) );
  AND U13919 ( .A(n12868), .B(n12867), .Z(n12989) );
  XOR U13920 ( .A(n12990), .B(n12991), .Z(n13037) );
  XOR U13921 ( .A(n13036), .B(n13037), .Z(n13038) );
  XNOR U13922 ( .A(n13039), .B(n13038), .Z(n13084) );
  NANDN U13923 ( .A(n12870), .B(n12869), .Z(n12874) );
  NAND U13924 ( .A(n12872), .B(n12871), .Z(n12873) );
  NAND U13925 ( .A(n12874), .B(n12873), .Z(n13027) );
  NANDN U13926 ( .A(n12876), .B(n12875), .Z(n12880) );
  NAND U13927 ( .A(n12878), .B(n12877), .Z(n12879) );
  NAND U13928 ( .A(n12880), .B(n12879), .Z(n13025) );
  OR U13929 ( .A(n12882), .B(n12881), .Z(n12886) );
  NANDN U13930 ( .A(n12884), .B(n12883), .Z(n12885) );
  NAND U13931 ( .A(n12886), .B(n12885), .Z(n13024) );
  XNOR U13932 ( .A(n13027), .B(n13026), .Z(n13085) );
  XNOR U13933 ( .A(n13084), .B(n13085), .Z(n13086) );
  NANDN U13934 ( .A(n12888), .B(n12887), .Z(n12892) );
  OR U13935 ( .A(n12890), .B(n12889), .Z(n12891) );
  AND U13936 ( .A(n12892), .B(n12891), .Z(n13087) );
  XOR U13937 ( .A(n13086), .B(n13087), .Z(n13104) );
  NANDN U13938 ( .A(n12898), .B(n12897), .Z(n12902) );
  NANDN U13939 ( .A(n12900), .B(n12899), .Z(n12901) );
  NAND U13940 ( .A(n12902), .B(n12901), .Z(n13093) );
  NANDN U13941 ( .A(n12908), .B(n12907), .Z(n12912) );
  NAND U13942 ( .A(n12910), .B(n12909), .Z(n12911) );
  NAND U13943 ( .A(n12912), .B(n12911), .Z(n13030) );
  NANDN U13944 ( .A(n12914), .B(n12913), .Z(n12918) );
  NAND U13945 ( .A(n12916), .B(n12915), .Z(n12917) );
  AND U13946 ( .A(n12918), .B(n12917), .Z(n13031) );
  XNOR U13947 ( .A(n13030), .B(n13031), .Z(n13032) );
  XNOR U13948 ( .A(b[9]), .B(a[89]), .Z(n13054) );
  NANDN U13949 ( .A(n13054), .B(n36925), .Z(n12921) );
  NANDN U13950 ( .A(n12919), .B(n36926), .Z(n12920) );
  NAND U13951 ( .A(n12921), .B(n12920), .Z(n12996) );
  XOR U13952 ( .A(b[15]), .B(n15562), .Z(n13057) );
  OR U13953 ( .A(n13057), .B(n37665), .Z(n12924) );
  NANDN U13954 ( .A(n12922), .B(n37604), .Z(n12923) );
  AND U13955 ( .A(n12924), .B(n12923), .Z(n12994) );
  XNOR U13956 ( .A(b[21]), .B(a[77]), .Z(n13060) );
  NANDN U13957 ( .A(n13060), .B(n38101), .Z(n12927) );
  NANDN U13958 ( .A(n12925), .B(n38102), .Z(n12926) );
  AND U13959 ( .A(n12927), .B(n12926), .Z(n12995) );
  XOR U13960 ( .A(n12996), .B(n12997), .Z(n12985) );
  XNOR U13961 ( .A(b[11]), .B(a[87]), .Z(n13063) );
  OR U13962 ( .A(n13063), .B(n37311), .Z(n12930) );
  NANDN U13963 ( .A(n12928), .B(n37218), .Z(n12929) );
  NAND U13964 ( .A(n12930), .B(n12929), .Z(n12983) );
  XOR U13965 ( .A(n1053), .B(a[85]), .Z(n13066) );
  NANDN U13966 ( .A(n13066), .B(n37424), .Z(n12933) );
  NANDN U13967 ( .A(n12931), .B(n37425), .Z(n12932) );
  NAND U13968 ( .A(n12933), .B(n12932), .Z(n12982) );
  XOR U13969 ( .A(n12985), .B(n12984), .Z(n12979) );
  NANDN U13970 ( .A(n1049), .B(a[97]), .Z(n12934) );
  XNOR U13971 ( .A(b[1]), .B(n12934), .Z(n12936) );
  NANDN U13972 ( .A(b[0]), .B(a[96]), .Z(n12935) );
  AND U13973 ( .A(n12936), .B(n12935), .Z(n13002) );
  NAND U13974 ( .A(n38490), .B(n12937), .Z(n12939) );
  XNOR U13975 ( .A(n1058), .B(a[69]), .Z(n13072) );
  NANDN U13976 ( .A(n1048), .B(n13072), .Z(n12938) );
  NAND U13977 ( .A(n12939), .B(n12938), .Z(n13000) );
  NANDN U13978 ( .A(n1059), .B(a[65]), .Z(n13001) );
  XNOR U13979 ( .A(n13000), .B(n13001), .Z(n13003) );
  XNOR U13980 ( .A(n13002), .B(n13003), .Z(n12977) );
  NANDN U13981 ( .A(n12940), .B(n38205), .Z(n12942) );
  XNOR U13982 ( .A(b[23]), .B(a[75]), .Z(n13075) );
  OR U13983 ( .A(n13075), .B(n38268), .Z(n12941) );
  NAND U13984 ( .A(n12942), .B(n12941), .Z(n13045) );
  XOR U13985 ( .A(b[7]), .B(a[91]), .Z(n13078) );
  NAND U13986 ( .A(n13078), .B(n36701), .Z(n12945) );
  NAND U13987 ( .A(n12943), .B(n36702), .Z(n12944) );
  NAND U13988 ( .A(n12945), .B(n12944), .Z(n13042) );
  XOR U13989 ( .A(b[25]), .B(a[73]), .Z(n13081) );
  NAND U13990 ( .A(n13081), .B(n38325), .Z(n12948) );
  NAND U13991 ( .A(n12946), .B(n38326), .Z(n12947) );
  AND U13992 ( .A(n12948), .B(n12947), .Z(n13043) );
  XNOR U13993 ( .A(n13042), .B(n13043), .Z(n13044) );
  XOR U13994 ( .A(n13045), .B(n13044), .Z(n12976) );
  XOR U13995 ( .A(n12979), .B(n12978), .Z(n13033) );
  XNOR U13996 ( .A(n13032), .B(n13033), .Z(n13090) );
  XOR U13997 ( .A(n13091), .B(n13090), .Z(n13092) );
  XNOR U13998 ( .A(n13093), .B(n13092), .Z(n13102) );
  XNOR U13999 ( .A(n13103), .B(n13102), .Z(n13105) );
  XNOR U14000 ( .A(n13104), .B(n13105), .Z(n13099) );
  XOR U14001 ( .A(n13098), .B(n13099), .Z(n12973) );
  NANDN U14002 ( .A(n12954), .B(n12953), .Z(n12958) );
  NANDN U14003 ( .A(n12956), .B(n12955), .Z(n12957) );
  NAND U14004 ( .A(n12958), .B(n12957), .Z(n12971) );
  XNOR U14005 ( .A(n12970), .B(n12971), .Z(n12972) );
  XNOR U14006 ( .A(n12973), .B(n12972), .Z(n12965) );
  XNOR U14007 ( .A(n12964), .B(n12965), .Z(n12966) );
  XNOR U14008 ( .A(n12967), .B(n12966), .Z(n13108) );
  XNOR U14009 ( .A(n13108), .B(sreg[321]), .Z(n13110) );
  NAND U14010 ( .A(n12959), .B(sreg[320]), .Z(n12963) );
  OR U14011 ( .A(n12961), .B(n12960), .Z(n12962) );
  AND U14012 ( .A(n12963), .B(n12962), .Z(n13109) );
  XOR U14013 ( .A(n13110), .B(n13109), .Z(c[321]) );
  NANDN U14014 ( .A(n12965), .B(n12964), .Z(n12969) );
  NAND U14015 ( .A(n12967), .B(n12966), .Z(n12968) );
  NAND U14016 ( .A(n12969), .B(n12968), .Z(n13116) );
  NANDN U14017 ( .A(n12971), .B(n12970), .Z(n12975) );
  NAND U14018 ( .A(n12973), .B(n12972), .Z(n12974) );
  NAND U14019 ( .A(n12975), .B(n12974), .Z(n13114) );
  NANDN U14020 ( .A(n12977), .B(n12976), .Z(n12981) );
  NANDN U14021 ( .A(n12979), .B(n12978), .Z(n12980) );
  NAND U14022 ( .A(n12981), .B(n12980), .Z(n13235) );
  OR U14023 ( .A(n12983), .B(n12982), .Z(n12987) );
  NAND U14024 ( .A(n12985), .B(n12984), .Z(n12986) );
  NAND U14025 ( .A(n12987), .B(n12986), .Z(n13173) );
  OR U14026 ( .A(n12989), .B(n12988), .Z(n12993) );
  NANDN U14027 ( .A(n12991), .B(n12990), .Z(n12992) );
  NAND U14028 ( .A(n12993), .B(n12992), .Z(n13172) );
  OR U14029 ( .A(n12995), .B(n12994), .Z(n12999) );
  NANDN U14030 ( .A(n12997), .B(n12996), .Z(n12998) );
  NAND U14031 ( .A(n12999), .B(n12998), .Z(n13171) );
  XOR U14032 ( .A(n13173), .B(n13174), .Z(n13232) );
  NANDN U14033 ( .A(n13001), .B(n13000), .Z(n13005) );
  NAND U14034 ( .A(n13003), .B(n13002), .Z(n13004) );
  NAND U14035 ( .A(n13005), .B(n13004), .Z(n13186) );
  XOR U14036 ( .A(b[19]), .B(n15068), .Z(n13129) );
  NANDN U14037 ( .A(n13129), .B(n37934), .Z(n13008) );
  NANDN U14038 ( .A(n13006), .B(n37935), .Z(n13007) );
  NAND U14039 ( .A(n13008), .B(n13007), .Z(n13198) );
  XOR U14040 ( .A(b[27]), .B(a[72]), .Z(n13132) );
  NAND U14041 ( .A(n38423), .B(n13132), .Z(n13011) );
  NAND U14042 ( .A(n13009), .B(n38424), .Z(n13010) );
  NAND U14043 ( .A(n13011), .B(n13010), .Z(n13195) );
  XNOR U14044 ( .A(b[5]), .B(a[94]), .Z(n13135) );
  NANDN U14045 ( .A(n13135), .B(n36587), .Z(n13014) );
  NANDN U14046 ( .A(n13012), .B(n36588), .Z(n13013) );
  AND U14047 ( .A(n13014), .B(n13013), .Z(n13196) );
  XNOR U14048 ( .A(n13195), .B(n13196), .Z(n13197) );
  XNOR U14049 ( .A(n13198), .B(n13197), .Z(n13184) );
  NAND U14050 ( .A(n13015), .B(n37762), .Z(n13017) );
  XNOR U14051 ( .A(b[17]), .B(a[82]), .Z(n13138) );
  NANDN U14052 ( .A(n13138), .B(n37764), .Z(n13016) );
  NAND U14053 ( .A(n13017), .B(n13016), .Z(n13156) );
  XNOR U14054 ( .A(b[31]), .B(a[68]), .Z(n13141) );
  NANDN U14055 ( .A(n13141), .B(n38552), .Z(n13020) );
  NANDN U14056 ( .A(n13018), .B(n38553), .Z(n13019) );
  NAND U14057 ( .A(n13020), .B(n13019), .Z(n13153) );
  OR U14058 ( .A(n13021), .B(n36105), .Z(n13023) );
  XNOR U14059 ( .A(b[3]), .B(a[96]), .Z(n13144) );
  NANDN U14060 ( .A(n13144), .B(n36107), .Z(n13022) );
  AND U14061 ( .A(n13023), .B(n13022), .Z(n13154) );
  XNOR U14062 ( .A(n13153), .B(n13154), .Z(n13155) );
  XOR U14063 ( .A(n13156), .B(n13155), .Z(n13183) );
  XNOR U14064 ( .A(n13184), .B(n13183), .Z(n13185) );
  XNOR U14065 ( .A(n13186), .B(n13185), .Z(n13233) );
  XNOR U14066 ( .A(n13232), .B(n13233), .Z(n13234) );
  XNOR U14067 ( .A(n13235), .B(n13234), .Z(n13253) );
  OR U14068 ( .A(n13025), .B(n13024), .Z(n13029) );
  NAND U14069 ( .A(n13027), .B(n13026), .Z(n13028) );
  NAND U14070 ( .A(n13029), .B(n13028), .Z(n13251) );
  NANDN U14071 ( .A(n13031), .B(n13030), .Z(n13035) );
  NANDN U14072 ( .A(n13033), .B(n13032), .Z(n13034) );
  NAND U14073 ( .A(n13035), .B(n13034), .Z(n13240) );
  OR U14074 ( .A(n13037), .B(n13036), .Z(n13041) );
  NAND U14075 ( .A(n13039), .B(n13038), .Z(n13040) );
  NAND U14076 ( .A(n13041), .B(n13040), .Z(n13239) );
  NANDN U14077 ( .A(n13043), .B(n13042), .Z(n13047) );
  NAND U14078 ( .A(n13045), .B(n13044), .Z(n13046) );
  NAND U14079 ( .A(n13047), .B(n13046), .Z(n13177) );
  NANDN U14080 ( .A(n13049), .B(n13048), .Z(n13053) );
  NAND U14081 ( .A(n13051), .B(n13050), .Z(n13052) );
  AND U14082 ( .A(n13053), .B(n13052), .Z(n13178) );
  XNOR U14083 ( .A(n13177), .B(n13178), .Z(n13179) );
  XNOR U14084 ( .A(b[9]), .B(a[90]), .Z(n13201) );
  NANDN U14085 ( .A(n13201), .B(n36925), .Z(n13056) );
  NANDN U14086 ( .A(n13054), .B(n36926), .Z(n13055) );
  NAND U14087 ( .A(n13056), .B(n13055), .Z(n13161) );
  XNOR U14088 ( .A(b[15]), .B(a[84]), .Z(n13204) );
  OR U14089 ( .A(n13204), .B(n37665), .Z(n13059) );
  NANDN U14090 ( .A(n13057), .B(n37604), .Z(n13058) );
  AND U14091 ( .A(n13059), .B(n13058), .Z(n13159) );
  XNOR U14092 ( .A(b[21]), .B(a[78]), .Z(n13207) );
  NANDN U14093 ( .A(n13207), .B(n38101), .Z(n13062) );
  NANDN U14094 ( .A(n13060), .B(n38102), .Z(n13061) );
  AND U14095 ( .A(n13062), .B(n13061), .Z(n13160) );
  XOR U14096 ( .A(n13161), .B(n13162), .Z(n13150) );
  XNOR U14097 ( .A(b[11]), .B(a[88]), .Z(n13210) );
  OR U14098 ( .A(n13210), .B(n37311), .Z(n13065) );
  NANDN U14099 ( .A(n13063), .B(n37218), .Z(n13064) );
  NAND U14100 ( .A(n13065), .B(n13064), .Z(n13148) );
  XOR U14101 ( .A(n1053), .B(a[86]), .Z(n13213) );
  NANDN U14102 ( .A(n13213), .B(n37424), .Z(n13068) );
  NANDN U14103 ( .A(n13066), .B(n37425), .Z(n13067) );
  AND U14104 ( .A(n13068), .B(n13067), .Z(n13147) );
  XNOR U14105 ( .A(n13148), .B(n13147), .Z(n13149) );
  XOR U14106 ( .A(n13150), .B(n13149), .Z(n13167) );
  NANDN U14107 ( .A(n1049), .B(a[98]), .Z(n13069) );
  XNOR U14108 ( .A(b[1]), .B(n13069), .Z(n13071) );
  NANDN U14109 ( .A(b[0]), .B(a[97]), .Z(n13070) );
  AND U14110 ( .A(n13071), .B(n13070), .Z(n13125) );
  NAND U14111 ( .A(n38490), .B(n13072), .Z(n13074) );
  XNOR U14112 ( .A(b[29]), .B(a[70]), .Z(n13220) );
  OR U14113 ( .A(n13220), .B(n1048), .Z(n13073) );
  NAND U14114 ( .A(n13074), .B(n13073), .Z(n13123) );
  NANDN U14115 ( .A(n1059), .B(a[66]), .Z(n13124) );
  XNOR U14116 ( .A(n13123), .B(n13124), .Z(n13126) );
  XOR U14117 ( .A(n13125), .B(n13126), .Z(n13165) );
  NANDN U14118 ( .A(n13075), .B(n38205), .Z(n13077) );
  XNOR U14119 ( .A(b[23]), .B(a[76]), .Z(n13223) );
  OR U14120 ( .A(n13223), .B(n38268), .Z(n13076) );
  NAND U14121 ( .A(n13077), .B(n13076), .Z(n13192) );
  XOR U14122 ( .A(b[7]), .B(a[92]), .Z(n13226) );
  NAND U14123 ( .A(n13226), .B(n36701), .Z(n13080) );
  NAND U14124 ( .A(n13078), .B(n36702), .Z(n13079) );
  NAND U14125 ( .A(n13080), .B(n13079), .Z(n13189) );
  XOR U14126 ( .A(b[25]), .B(a[74]), .Z(n13229) );
  NAND U14127 ( .A(n13229), .B(n38325), .Z(n13083) );
  NAND U14128 ( .A(n13081), .B(n38326), .Z(n13082) );
  AND U14129 ( .A(n13083), .B(n13082), .Z(n13190) );
  XNOR U14130 ( .A(n13189), .B(n13190), .Z(n13191) );
  XNOR U14131 ( .A(n13192), .B(n13191), .Z(n13166) );
  XOR U14132 ( .A(n13165), .B(n13166), .Z(n13168) );
  XNOR U14133 ( .A(n13167), .B(n13168), .Z(n13180) );
  XNOR U14134 ( .A(n13179), .B(n13180), .Z(n13238) );
  XNOR U14135 ( .A(n13239), .B(n13238), .Z(n13241) );
  XNOR U14136 ( .A(n13240), .B(n13241), .Z(n13250) );
  XNOR U14137 ( .A(n13251), .B(n13250), .Z(n13252) );
  XOR U14138 ( .A(n13253), .B(n13252), .Z(n13247) );
  NANDN U14139 ( .A(n13085), .B(n13084), .Z(n13089) );
  NAND U14140 ( .A(n13087), .B(n13086), .Z(n13088) );
  NAND U14141 ( .A(n13089), .B(n13088), .Z(n13244) );
  NAND U14142 ( .A(n13091), .B(n13090), .Z(n13095) );
  NAND U14143 ( .A(n13093), .B(n13092), .Z(n13094) );
  NAND U14144 ( .A(n13095), .B(n13094), .Z(n13245) );
  XNOR U14145 ( .A(n13244), .B(n13245), .Z(n13246) );
  XNOR U14146 ( .A(n13247), .B(n13246), .Z(n13120) );
  NANDN U14147 ( .A(n13097), .B(n13096), .Z(n13101) );
  NANDN U14148 ( .A(n13099), .B(n13098), .Z(n13100) );
  NAND U14149 ( .A(n13101), .B(n13100), .Z(n13118) );
  OR U14150 ( .A(n13103), .B(n13102), .Z(n13107) );
  OR U14151 ( .A(n13105), .B(n13104), .Z(n13106) );
  AND U14152 ( .A(n13107), .B(n13106), .Z(n13117) );
  XNOR U14153 ( .A(n13118), .B(n13117), .Z(n13119) );
  XNOR U14154 ( .A(n13120), .B(n13119), .Z(n13113) );
  XOR U14155 ( .A(n13114), .B(n13113), .Z(n13115) );
  XNOR U14156 ( .A(n13116), .B(n13115), .Z(n13256) );
  XNOR U14157 ( .A(n13256), .B(sreg[322]), .Z(n13258) );
  NAND U14158 ( .A(n13108), .B(sreg[321]), .Z(n13112) );
  OR U14159 ( .A(n13110), .B(n13109), .Z(n13111) );
  AND U14160 ( .A(n13112), .B(n13111), .Z(n13257) );
  XOR U14161 ( .A(n13258), .B(n13257), .Z(c[322]) );
  NANDN U14162 ( .A(n13118), .B(n13117), .Z(n13122) );
  NANDN U14163 ( .A(n13120), .B(n13119), .Z(n13121) );
  NAND U14164 ( .A(n13122), .B(n13121), .Z(n13262) );
  NANDN U14165 ( .A(n13124), .B(n13123), .Z(n13128) );
  NAND U14166 ( .A(n13126), .B(n13125), .Z(n13127) );
  NAND U14167 ( .A(n13128), .B(n13127), .Z(n13336) );
  XNOR U14168 ( .A(b[19]), .B(a[81]), .Z(n13303) );
  NANDN U14169 ( .A(n13303), .B(n37934), .Z(n13131) );
  NANDN U14170 ( .A(n13129), .B(n37935), .Z(n13130) );
  NAND U14171 ( .A(n13131), .B(n13130), .Z(n13348) );
  XOR U14172 ( .A(b[27]), .B(a[73]), .Z(n13306) );
  NAND U14173 ( .A(n38423), .B(n13306), .Z(n13134) );
  NAND U14174 ( .A(n13132), .B(n38424), .Z(n13133) );
  NAND U14175 ( .A(n13134), .B(n13133), .Z(n13345) );
  XNOR U14176 ( .A(b[5]), .B(a[95]), .Z(n13309) );
  NANDN U14177 ( .A(n13309), .B(n36587), .Z(n13137) );
  NANDN U14178 ( .A(n13135), .B(n36588), .Z(n13136) );
  AND U14179 ( .A(n13137), .B(n13136), .Z(n13346) );
  XNOR U14180 ( .A(n13345), .B(n13346), .Z(n13347) );
  XNOR U14181 ( .A(n13348), .B(n13347), .Z(n13333) );
  NANDN U14182 ( .A(n13138), .B(n37762), .Z(n13140) );
  XNOR U14183 ( .A(b[17]), .B(a[83]), .Z(n13312) );
  NANDN U14184 ( .A(n13312), .B(n37764), .Z(n13139) );
  NAND U14185 ( .A(n13140), .B(n13139), .Z(n13287) );
  XNOR U14186 ( .A(b[31]), .B(a[69]), .Z(n13315) );
  NANDN U14187 ( .A(n13315), .B(n38552), .Z(n13143) );
  NANDN U14188 ( .A(n13141), .B(n38553), .Z(n13142) );
  AND U14189 ( .A(n13143), .B(n13142), .Z(n13285) );
  OR U14190 ( .A(n13144), .B(n36105), .Z(n13146) );
  XNOR U14191 ( .A(b[3]), .B(a[97]), .Z(n13318) );
  NANDN U14192 ( .A(n13318), .B(n36107), .Z(n13145) );
  AND U14193 ( .A(n13146), .B(n13145), .Z(n13286) );
  XOR U14194 ( .A(n13287), .B(n13288), .Z(n13334) );
  XOR U14195 ( .A(n13333), .B(n13334), .Z(n13335) );
  XNOR U14196 ( .A(n13336), .B(n13335), .Z(n13381) );
  NANDN U14197 ( .A(n13148), .B(n13147), .Z(n13152) );
  NAND U14198 ( .A(n13150), .B(n13149), .Z(n13151) );
  NAND U14199 ( .A(n13152), .B(n13151), .Z(n13324) );
  NANDN U14200 ( .A(n13154), .B(n13153), .Z(n13158) );
  NAND U14201 ( .A(n13156), .B(n13155), .Z(n13157) );
  NAND U14202 ( .A(n13158), .B(n13157), .Z(n13322) );
  OR U14203 ( .A(n13160), .B(n13159), .Z(n13164) );
  NANDN U14204 ( .A(n13162), .B(n13161), .Z(n13163) );
  NAND U14205 ( .A(n13164), .B(n13163), .Z(n13321) );
  XNOR U14206 ( .A(n13324), .B(n13323), .Z(n13382) );
  XOR U14207 ( .A(n13381), .B(n13382), .Z(n13384) );
  NANDN U14208 ( .A(n13166), .B(n13165), .Z(n13170) );
  OR U14209 ( .A(n13168), .B(n13167), .Z(n13169) );
  NAND U14210 ( .A(n13170), .B(n13169), .Z(n13383) );
  XOR U14211 ( .A(n13384), .B(n13383), .Z(n13401) );
  OR U14212 ( .A(n13172), .B(n13171), .Z(n13176) );
  NANDN U14213 ( .A(n13174), .B(n13173), .Z(n13175) );
  NAND U14214 ( .A(n13176), .B(n13175), .Z(n13400) );
  NANDN U14215 ( .A(n13178), .B(n13177), .Z(n13182) );
  NANDN U14216 ( .A(n13180), .B(n13179), .Z(n13181) );
  NAND U14217 ( .A(n13182), .B(n13181), .Z(n13389) );
  NANDN U14218 ( .A(n13184), .B(n13183), .Z(n13188) );
  NAND U14219 ( .A(n13186), .B(n13185), .Z(n13187) );
  NAND U14220 ( .A(n13188), .B(n13187), .Z(n13388) );
  NANDN U14221 ( .A(n13190), .B(n13189), .Z(n13194) );
  NAND U14222 ( .A(n13192), .B(n13191), .Z(n13193) );
  NAND U14223 ( .A(n13194), .B(n13193), .Z(n13327) );
  NANDN U14224 ( .A(n13196), .B(n13195), .Z(n13200) );
  NAND U14225 ( .A(n13198), .B(n13197), .Z(n13199) );
  AND U14226 ( .A(n13200), .B(n13199), .Z(n13328) );
  XNOR U14227 ( .A(n13327), .B(n13328), .Z(n13329) );
  XNOR U14228 ( .A(b[9]), .B(a[91]), .Z(n13351) );
  NANDN U14229 ( .A(n13351), .B(n36925), .Z(n13203) );
  NANDN U14230 ( .A(n13201), .B(n36926), .Z(n13202) );
  NAND U14231 ( .A(n13203), .B(n13202), .Z(n13293) );
  XNOR U14232 ( .A(b[15]), .B(a[85]), .Z(n13354) );
  OR U14233 ( .A(n13354), .B(n37665), .Z(n13206) );
  NANDN U14234 ( .A(n13204), .B(n37604), .Z(n13205) );
  AND U14235 ( .A(n13206), .B(n13205), .Z(n13291) );
  XNOR U14236 ( .A(b[21]), .B(a[79]), .Z(n13357) );
  NANDN U14237 ( .A(n13357), .B(n38101), .Z(n13209) );
  NANDN U14238 ( .A(n13207), .B(n38102), .Z(n13208) );
  AND U14239 ( .A(n13209), .B(n13208), .Z(n13292) );
  XOR U14240 ( .A(n13293), .B(n13294), .Z(n13282) );
  XNOR U14241 ( .A(b[11]), .B(a[89]), .Z(n13360) );
  OR U14242 ( .A(n13360), .B(n37311), .Z(n13212) );
  NANDN U14243 ( .A(n13210), .B(n37218), .Z(n13211) );
  NAND U14244 ( .A(n13212), .B(n13211), .Z(n13280) );
  XOR U14245 ( .A(n1053), .B(a[87]), .Z(n13363) );
  NANDN U14246 ( .A(n13363), .B(n37424), .Z(n13215) );
  NANDN U14247 ( .A(n13213), .B(n37425), .Z(n13214) );
  NAND U14248 ( .A(n13215), .B(n13214), .Z(n13279) );
  XOR U14249 ( .A(n13282), .B(n13281), .Z(n13276) );
  NANDN U14250 ( .A(n1049), .B(a[99]), .Z(n13216) );
  XNOR U14251 ( .A(b[1]), .B(n13216), .Z(n13218) );
  NANDN U14252 ( .A(b[0]), .B(a[98]), .Z(n13217) );
  AND U14253 ( .A(n13218), .B(n13217), .Z(n13300) );
  ANDN U14254 ( .B(b[31]), .A(n13219), .Z(n13297) );
  NANDN U14255 ( .A(n13220), .B(n38490), .Z(n13222) );
  XNOR U14256 ( .A(n1058), .B(a[71]), .Z(n13366) );
  NANDN U14257 ( .A(n1048), .B(n13366), .Z(n13221) );
  NAND U14258 ( .A(n13222), .B(n13221), .Z(n13298) );
  XOR U14259 ( .A(n13297), .B(n13298), .Z(n13299) );
  XNOR U14260 ( .A(n13300), .B(n13299), .Z(n13273) );
  NANDN U14261 ( .A(n13223), .B(n38205), .Z(n13225) );
  XNOR U14262 ( .A(b[23]), .B(a[77]), .Z(n13372) );
  OR U14263 ( .A(n13372), .B(n38268), .Z(n13224) );
  NAND U14264 ( .A(n13225), .B(n13224), .Z(n13342) );
  XNOR U14265 ( .A(b[7]), .B(a[93]), .Z(n13375) );
  NANDN U14266 ( .A(n13375), .B(n36701), .Z(n13228) );
  NAND U14267 ( .A(n13226), .B(n36702), .Z(n13227) );
  NAND U14268 ( .A(n13228), .B(n13227), .Z(n13339) );
  XOR U14269 ( .A(b[25]), .B(a[75]), .Z(n13378) );
  NAND U14270 ( .A(n13378), .B(n38325), .Z(n13231) );
  NAND U14271 ( .A(n13229), .B(n38326), .Z(n13230) );
  AND U14272 ( .A(n13231), .B(n13230), .Z(n13340) );
  XNOR U14273 ( .A(n13339), .B(n13340), .Z(n13341) );
  XNOR U14274 ( .A(n13342), .B(n13341), .Z(n13274) );
  XOR U14275 ( .A(n13276), .B(n13275), .Z(n13330) );
  XNOR U14276 ( .A(n13329), .B(n13330), .Z(n13387) );
  XNOR U14277 ( .A(n13388), .B(n13387), .Z(n13390) );
  XNOR U14278 ( .A(n13389), .B(n13390), .Z(n13399) );
  XOR U14279 ( .A(n13400), .B(n13399), .Z(n13402) );
  NANDN U14280 ( .A(n13233), .B(n13232), .Z(n13237) );
  NAND U14281 ( .A(n13235), .B(n13234), .Z(n13236) );
  NAND U14282 ( .A(n13237), .B(n13236), .Z(n13394) );
  NAND U14283 ( .A(n13239), .B(n13238), .Z(n13243) );
  NANDN U14284 ( .A(n13241), .B(n13240), .Z(n13242) );
  AND U14285 ( .A(n13243), .B(n13242), .Z(n13393) );
  XNOR U14286 ( .A(n13394), .B(n13393), .Z(n13395) );
  XOR U14287 ( .A(n13396), .B(n13395), .Z(n13269) );
  NANDN U14288 ( .A(n13245), .B(n13244), .Z(n13249) );
  NAND U14289 ( .A(n13247), .B(n13246), .Z(n13248) );
  NAND U14290 ( .A(n13249), .B(n13248), .Z(n13267) );
  NANDN U14291 ( .A(n13251), .B(n13250), .Z(n13255) );
  NANDN U14292 ( .A(n13253), .B(n13252), .Z(n13254) );
  NAND U14293 ( .A(n13255), .B(n13254), .Z(n13268) );
  XNOR U14294 ( .A(n13267), .B(n13268), .Z(n13270) );
  XOR U14295 ( .A(n13269), .B(n13270), .Z(n13261) );
  XOR U14296 ( .A(n13262), .B(n13261), .Z(n13263) );
  XNOR U14297 ( .A(n13264), .B(n13263), .Z(n13405) );
  XNOR U14298 ( .A(n13405), .B(sreg[323]), .Z(n13407) );
  NAND U14299 ( .A(n13256), .B(sreg[322]), .Z(n13260) );
  OR U14300 ( .A(n13258), .B(n13257), .Z(n13259) );
  AND U14301 ( .A(n13260), .B(n13259), .Z(n13406) );
  XOR U14302 ( .A(n13407), .B(n13406), .Z(c[323]) );
  NAND U14303 ( .A(n13262), .B(n13261), .Z(n13266) );
  NAND U14304 ( .A(n13264), .B(n13263), .Z(n13265) );
  NAND U14305 ( .A(n13266), .B(n13265), .Z(n13413) );
  NANDN U14306 ( .A(n13268), .B(n13267), .Z(n13272) );
  NAND U14307 ( .A(n13270), .B(n13269), .Z(n13271) );
  NAND U14308 ( .A(n13272), .B(n13271), .Z(n13411) );
  OR U14309 ( .A(n13274), .B(n13273), .Z(n13278) );
  NANDN U14310 ( .A(n13276), .B(n13275), .Z(n13277) );
  NAND U14311 ( .A(n13278), .B(n13277), .Z(n13543) );
  OR U14312 ( .A(n13280), .B(n13279), .Z(n13284) );
  NAND U14313 ( .A(n13282), .B(n13281), .Z(n13283) );
  NAND U14314 ( .A(n13284), .B(n13283), .Z(n13482) );
  OR U14315 ( .A(n13286), .B(n13285), .Z(n13290) );
  NANDN U14316 ( .A(n13288), .B(n13287), .Z(n13289) );
  NAND U14317 ( .A(n13290), .B(n13289), .Z(n13481) );
  OR U14318 ( .A(n13292), .B(n13291), .Z(n13296) );
  NANDN U14319 ( .A(n13294), .B(n13293), .Z(n13295) );
  NAND U14320 ( .A(n13296), .B(n13295), .Z(n13480) );
  XOR U14321 ( .A(n13482), .B(n13483), .Z(n13541) );
  OR U14322 ( .A(n13298), .B(n13297), .Z(n13302) );
  NANDN U14323 ( .A(n13300), .B(n13299), .Z(n13301) );
  NAND U14324 ( .A(n13302), .B(n13301), .Z(n13494) );
  XOR U14325 ( .A(b[19]), .B(n15424), .Z(n13438) );
  NANDN U14326 ( .A(n13438), .B(n37934), .Z(n13305) );
  NANDN U14327 ( .A(n13303), .B(n37935), .Z(n13304) );
  NAND U14328 ( .A(n13305), .B(n13304), .Z(n13507) );
  XOR U14329 ( .A(b[27]), .B(a[74]), .Z(n13441) );
  NAND U14330 ( .A(n38423), .B(n13441), .Z(n13308) );
  NAND U14331 ( .A(n13306), .B(n38424), .Z(n13307) );
  NAND U14332 ( .A(n13308), .B(n13307), .Z(n13504) );
  XNOR U14333 ( .A(b[5]), .B(a[96]), .Z(n13444) );
  NANDN U14334 ( .A(n13444), .B(n36587), .Z(n13311) );
  NANDN U14335 ( .A(n13309), .B(n36588), .Z(n13310) );
  AND U14336 ( .A(n13311), .B(n13310), .Z(n13505) );
  XNOR U14337 ( .A(n13504), .B(n13505), .Z(n13506) );
  XNOR U14338 ( .A(n13507), .B(n13506), .Z(n13493) );
  NANDN U14339 ( .A(n13312), .B(n37762), .Z(n13314) );
  XOR U14340 ( .A(b[17]), .B(a[84]), .Z(n13447) );
  NAND U14341 ( .A(n13447), .B(n37764), .Z(n13313) );
  NAND U14342 ( .A(n13314), .B(n13313), .Z(n13465) );
  XNOR U14343 ( .A(b[31]), .B(a[70]), .Z(n13450) );
  NANDN U14344 ( .A(n13450), .B(n38552), .Z(n13317) );
  NANDN U14345 ( .A(n13315), .B(n38553), .Z(n13316) );
  NAND U14346 ( .A(n13317), .B(n13316), .Z(n13462) );
  OR U14347 ( .A(n13318), .B(n36105), .Z(n13320) );
  XNOR U14348 ( .A(b[3]), .B(a[98]), .Z(n13453) );
  NANDN U14349 ( .A(n13453), .B(n36107), .Z(n13319) );
  AND U14350 ( .A(n13320), .B(n13319), .Z(n13463) );
  XNOR U14351 ( .A(n13462), .B(n13463), .Z(n13464) );
  XOR U14352 ( .A(n13465), .B(n13464), .Z(n13492) );
  XOR U14353 ( .A(n13493), .B(n13492), .Z(n13495) );
  XOR U14354 ( .A(n13494), .B(n13495), .Z(n13540) );
  XOR U14355 ( .A(n13541), .B(n13540), .Z(n13542) );
  XNOR U14356 ( .A(n13543), .B(n13542), .Z(n13429) );
  OR U14357 ( .A(n13322), .B(n13321), .Z(n13326) );
  NAND U14358 ( .A(n13324), .B(n13323), .Z(n13325) );
  NAND U14359 ( .A(n13326), .B(n13325), .Z(n13427) );
  NANDN U14360 ( .A(n13328), .B(n13327), .Z(n13332) );
  NANDN U14361 ( .A(n13330), .B(n13329), .Z(n13331) );
  NAND U14362 ( .A(n13332), .B(n13331), .Z(n13548) );
  OR U14363 ( .A(n13334), .B(n13333), .Z(n13338) );
  NAND U14364 ( .A(n13336), .B(n13335), .Z(n13337) );
  NAND U14365 ( .A(n13338), .B(n13337), .Z(n13547) );
  NANDN U14366 ( .A(n13340), .B(n13339), .Z(n13344) );
  NAND U14367 ( .A(n13342), .B(n13341), .Z(n13343) );
  NAND U14368 ( .A(n13344), .B(n13343), .Z(n13486) );
  NANDN U14369 ( .A(n13346), .B(n13345), .Z(n13350) );
  NAND U14370 ( .A(n13348), .B(n13347), .Z(n13349) );
  AND U14371 ( .A(n13350), .B(n13349), .Z(n13487) );
  XNOR U14372 ( .A(n13486), .B(n13487), .Z(n13488) );
  XNOR U14373 ( .A(b[9]), .B(a[92]), .Z(n13510) );
  NANDN U14374 ( .A(n13510), .B(n36925), .Z(n13353) );
  NANDN U14375 ( .A(n13351), .B(n36926), .Z(n13352) );
  NAND U14376 ( .A(n13353), .B(n13352), .Z(n13470) );
  XNOR U14377 ( .A(b[15]), .B(a[86]), .Z(n13513) );
  OR U14378 ( .A(n13513), .B(n37665), .Z(n13356) );
  NANDN U14379 ( .A(n13354), .B(n37604), .Z(n13355) );
  AND U14380 ( .A(n13356), .B(n13355), .Z(n13468) );
  XOR U14381 ( .A(b[21]), .B(n15068), .Z(n13516) );
  NANDN U14382 ( .A(n13516), .B(n38101), .Z(n13359) );
  NANDN U14383 ( .A(n13357), .B(n38102), .Z(n13358) );
  AND U14384 ( .A(n13359), .B(n13358), .Z(n13469) );
  XOR U14385 ( .A(n13470), .B(n13471), .Z(n13459) );
  XNOR U14386 ( .A(b[11]), .B(a[90]), .Z(n13519) );
  OR U14387 ( .A(n13519), .B(n37311), .Z(n13362) );
  NANDN U14388 ( .A(n13360), .B(n37218), .Z(n13361) );
  NAND U14389 ( .A(n13362), .B(n13361), .Z(n13457) );
  XOR U14390 ( .A(n1053), .B(a[88]), .Z(n13522) );
  NANDN U14391 ( .A(n13522), .B(n37424), .Z(n13365) );
  NANDN U14392 ( .A(n13363), .B(n37425), .Z(n13364) );
  AND U14393 ( .A(n13365), .B(n13364), .Z(n13456) );
  XNOR U14394 ( .A(n13457), .B(n13456), .Z(n13458) );
  XOR U14395 ( .A(n13459), .B(n13458), .Z(n13476) );
  NAND U14396 ( .A(n13366), .B(n38490), .Z(n13368) );
  XNOR U14397 ( .A(n1058), .B(a[72]), .Z(n13528) );
  NANDN U14398 ( .A(n1048), .B(n13528), .Z(n13367) );
  NAND U14399 ( .A(n13368), .B(n13367), .Z(n13432) );
  NANDN U14400 ( .A(n1059), .B(a[68]), .Z(n13433) );
  XNOR U14401 ( .A(n13432), .B(n13433), .Z(n13435) );
  NANDN U14402 ( .A(n1049), .B(a[100]), .Z(n13369) );
  XNOR U14403 ( .A(b[1]), .B(n13369), .Z(n13371) );
  IV U14404 ( .A(a[99]), .Z(n17884) );
  NANDN U14405 ( .A(n17884), .B(n1049), .Z(n13370) );
  AND U14406 ( .A(n13371), .B(n13370), .Z(n13434) );
  XOR U14407 ( .A(n13435), .B(n13434), .Z(n13474) );
  NANDN U14408 ( .A(n13372), .B(n38205), .Z(n13374) );
  XNOR U14409 ( .A(b[23]), .B(a[78]), .Z(n13531) );
  OR U14410 ( .A(n13531), .B(n38268), .Z(n13373) );
  NAND U14411 ( .A(n13374), .B(n13373), .Z(n13501) );
  XOR U14412 ( .A(b[7]), .B(a[94]), .Z(n13534) );
  NAND U14413 ( .A(n13534), .B(n36701), .Z(n13377) );
  NANDN U14414 ( .A(n13375), .B(n36702), .Z(n13376) );
  NAND U14415 ( .A(n13377), .B(n13376), .Z(n13498) );
  XOR U14416 ( .A(b[25]), .B(a[76]), .Z(n13537) );
  NAND U14417 ( .A(n13537), .B(n38325), .Z(n13380) );
  NAND U14418 ( .A(n13378), .B(n38326), .Z(n13379) );
  AND U14419 ( .A(n13380), .B(n13379), .Z(n13499) );
  XNOR U14420 ( .A(n13498), .B(n13499), .Z(n13500) );
  XNOR U14421 ( .A(n13501), .B(n13500), .Z(n13475) );
  XOR U14422 ( .A(n13474), .B(n13475), .Z(n13477) );
  XNOR U14423 ( .A(n13476), .B(n13477), .Z(n13489) );
  XNOR U14424 ( .A(n13488), .B(n13489), .Z(n13546) );
  XNOR U14425 ( .A(n13547), .B(n13546), .Z(n13549) );
  XNOR U14426 ( .A(n13548), .B(n13549), .Z(n13426) );
  XNOR U14427 ( .A(n13427), .B(n13426), .Z(n13428) );
  XOR U14428 ( .A(n13429), .B(n13428), .Z(n13423) );
  NANDN U14429 ( .A(n13382), .B(n13381), .Z(n13386) );
  OR U14430 ( .A(n13384), .B(n13383), .Z(n13385) );
  NAND U14431 ( .A(n13386), .B(n13385), .Z(n13420) );
  NAND U14432 ( .A(n13388), .B(n13387), .Z(n13392) );
  NANDN U14433 ( .A(n13390), .B(n13389), .Z(n13391) );
  NAND U14434 ( .A(n13392), .B(n13391), .Z(n13421) );
  XNOR U14435 ( .A(n13420), .B(n13421), .Z(n13422) );
  XNOR U14436 ( .A(n13423), .B(n13422), .Z(n13417) );
  NANDN U14437 ( .A(n13394), .B(n13393), .Z(n13398) );
  NAND U14438 ( .A(n13396), .B(n13395), .Z(n13397) );
  NAND U14439 ( .A(n13398), .B(n13397), .Z(n13414) );
  NANDN U14440 ( .A(n13400), .B(n13399), .Z(n13404) );
  OR U14441 ( .A(n13402), .B(n13401), .Z(n13403) );
  NAND U14442 ( .A(n13404), .B(n13403), .Z(n13415) );
  XNOR U14443 ( .A(n13414), .B(n13415), .Z(n13416) );
  XNOR U14444 ( .A(n13417), .B(n13416), .Z(n13410) );
  XOR U14445 ( .A(n13411), .B(n13410), .Z(n13412) );
  XNOR U14446 ( .A(n13413), .B(n13412), .Z(n13552) );
  XNOR U14447 ( .A(n13552), .B(sreg[324]), .Z(n13554) );
  NAND U14448 ( .A(n13405), .B(sreg[323]), .Z(n13409) );
  OR U14449 ( .A(n13407), .B(n13406), .Z(n13408) );
  AND U14450 ( .A(n13409), .B(n13408), .Z(n13553) );
  XOR U14451 ( .A(n13554), .B(n13553), .Z(c[324]) );
  NANDN U14452 ( .A(n13415), .B(n13414), .Z(n13419) );
  NANDN U14453 ( .A(n13417), .B(n13416), .Z(n13418) );
  NAND U14454 ( .A(n13419), .B(n13418), .Z(n13558) );
  NANDN U14455 ( .A(n13421), .B(n13420), .Z(n13425) );
  NAND U14456 ( .A(n13423), .B(n13422), .Z(n13424) );
  NAND U14457 ( .A(n13425), .B(n13424), .Z(n13563) );
  NANDN U14458 ( .A(n13427), .B(n13426), .Z(n13431) );
  NANDN U14459 ( .A(n13429), .B(n13428), .Z(n13430) );
  NAND U14460 ( .A(n13431), .B(n13430), .Z(n13564) );
  XNOR U14461 ( .A(n13563), .B(n13564), .Z(n13565) );
  NANDN U14462 ( .A(n13433), .B(n13432), .Z(n13437) );
  NAND U14463 ( .A(n13435), .B(n13434), .Z(n13436) );
  NAND U14464 ( .A(n13437), .B(n13436), .Z(n13632) );
  XOR U14465 ( .A(b[19]), .B(n15562), .Z(n13575) );
  NANDN U14466 ( .A(n13575), .B(n37934), .Z(n13440) );
  NANDN U14467 ( .A(n13438), .B(n37935), .Z(n13439) );
  NAND U14468 ( .A(n13440), .B(n13439), .Z(n13642) );
  XOR U14469 ( .A(b[27]), .B(a[75]), .Z(n13578) );
  NAND U14470 ( .A(n38423), .B(n13578), .Z(n13443) );
  NAND U14471 ( .A(n13441), .B(n38424), .Z(n13442) );
  NAND U14472 ( .A(n13443), .B(n13442), .Z(n13639) );
  XNOR U14473 ( .A(b[5]), .B(a[97]), .Z(n13581) );
  NANDN U14474 ( .A(n13581), .B(n36587), .Z(n13446) );
  NANDN U14475 ( .A(n13444), .B(n36588), .Z(n13445) );
  AND U14476 ( .A(n13446), .B(n13445), .Z(n13640) );
  XNOR U14477 ( .A(n13639), .B(n13640), .Z(n13641) );
  XNOR U14478 ( .A(n13642), .B(n13641), .Z(n13630) );
  NAND U14479 ( .A(n13447), .B(n37762), .Z(n13449) );
  XOR U14480 ( .A(b[17]), .B(a[85]), .Z(n13584) );
  NAND U14481 ( .A(n13584), .B(n37764), .Z(n13448) );
  NAND U14482 ( .A(n13449), .B(n13448), .Z(n13602) );
  XNOR U14483 ( .A(b[31]), .B(a[71]), .Z(n13587) );
  NANDN U14484 ( .A(n13587), .B(n38552), .Z(n13452) );
  NANDN U14485 ( .A(n13450), .B(n38553), .Z(n13451) );
  NAND U14486 ( .A(n13452), .B(n13451), .Z(n13599) );
  OR U14487 ( .A(n13453), .B(n36105), .Z(n13455) );
  XOR U14488 ( .A(b[3]), .B(n17884), .Z(n13590) );
  NANDN U14489 ( .A(n13590), .B(n36107), .Z(n13454) );
  AND U14490 ( .A(n13455), .B(n13454), .Z(n13600) );
  XNOR U14491 ( .A(n13599), .B(n13600), .Z(n13601) );
  XOR U14492 ( .A(n13602), .B(n13601), .Z(n13629) );
  XNOR U14493 ( .A(n13630), .B(n13629), .Z(n13631) );
  XNOR U14494 ( .A(n13632), .B(n13631), .Z(n13675) );
  NANDN U14495 ( .A(n13457), .B(n13456), .Z(n13461) );
  NAND U14496 ( .A(n13459), .B(n13458), .Z(n13460) );
  NAND U14497 ( .A(n13461), .B(n13460), .Z(n13620) );
  NANDN U14498 ( .A(n13463), .B(n13462), .Z(n13467) );
  NAND U14499 ( .A(n13465), .B(n13464), .Z(n13466) );
  NAND U14500 ( .A(n13467), .B(n13466), .Z(n13618) );
  OR U14501 ( .A(n13469), .B(n13468), .Z(n13473) );
  NANDN U14502 ( .A(n13471), .B(n13470), .Z(n13472) );
  NAND U14503 ( .A(n13473), .B(n13472), .Z(n13617) );
  XNOR U14504 ( .A(n13620), .B(n13619), .Z(n13676) );
  XOR U14505 ( .A(n13675), .B(n13676), .Z(n13678) );
  NANDN U14506 ( .A(n13475), .B(n13474), .Z(n13479) );
  OR U14507 ( .A(n13477), .B(n13476), .Z(n13478) );
  NAND U14508 ( .A(n13479), .B(n13478), .Z(n13677) );
  XOR U14509 ( .A(n13678), .B(n13677), .Z(n13695) );
  OR U14510 ( .A(n13481), .B(n13480), .Z(n13485) );
  NANDN U14511 ( .A(n13483), .B(n13482), .Z(n13484) );
  NAND U14512 ( .A(n13485), .B(n13484), .Z(n13694) );
  NANDN U14513 ( .A(n13487), .B(n13486), .Z(n13491) );
  NANDN U14514 ( .A(n13489), .B(n13488), .Z(n13490) );
  NAND U14515 ( .A(n13491), .B(n13490), .Z(n13683) );
  NANDN U14516 ( .A(n13493), .B(n13492), .Z(n13497) );
  OR U14517 ( .A(n13495), .B(n13494), .Z(n13496) );
  NAND U14518 ( .A(n13497), .B(n13496), .Z(n13682) );
  NANDN U14519 ( .A(n13499), .B(n13498), .Z(n13503) );
  NAND U14520 ( .A(n13501), .B(n13500), .Z(n13502) );
  NAND U14521 ( .A(n13503), .B(n13502), .Z(n13623) );
  NANDN U14522 ( .A(n13505), .B(n13504), .Z(n13509) );
  NAND U14523 ( .A(n13507), .B(n13506), .Z(n13508) );
  AND U14524 ( .A(n13509), .B(n13508), .Z(n13624) );
  XNOR U14525 ( .A(n13623), .B(n13624), .Z(n13625) );
  XOR U14526 ( .A(b[9]), .B(n17031), .Z(n13645) );
  NANDN U14527 ( .A(n13645), .B(n36925), .Z(n13512) );
  NANDN U14528 ( .A(n13510), .B(n36926), .Z(n13511) );
  NAND U14529 ( .A(n13512), .B(n13511), .Z(n13607) );
  XNOR U14530 ( .A(b[15]), .B(a[87]), .Z(n13648) );
  OR U14531 ( .A(n13648), .B(n37665), .Z(n13515) );
  NANDN U14532 ( .A(n13513), .B(n37604), .Z(n13514) );
  AND U14533 ( .A(n13515), .B(n13514), .Z(n13605) );
  XNOR U14534 ( .A(b[21]), .B(a[81]), .Z(n13651) );
  NANDN U14535 ( .A(n13651), .B(n38101), .Z(n13518) );
  NANDN U14536 ( .A(n13516), .B(n38102), .Z(n13517) );
  AND U14537 ( .A(n13518), .B(n13517), .Z(n13606) );
  XOR U14538 ( .A(n13607), .B(n13608), .Z(n13596) );
  XNOR U14539 ( .A(b[11]), .B(a[91]), .Z(n13654) );
  OR U14540 ( .A(n13654), .B(n37311), .Z(n13521) );
  NANDN U14541 ( .A(n13519), .B(n37218), .Z(n13520) );
  NAND U14542 ( .A(n13521), .B(n13520), .Z(n13594) );
  XOR U14543 ( .A(n1053), .B(a[89]), .Z(n13657) );
  NANDN U14544 ( .A(n13657), .B(n37424), .Z(n13524) );
  NANDN U14545 ( .A(n13522), .B(n37425), .Z(n13523) );
  AND U14546 ( .A(n13524), .B(n13523), .Z(n13593) );
  XNOR U14547 ( .A(n13594), .B(n13593), .Z(n13595) );
  XOR U14548 ( .A(n13596), .B(n13595), .Z(n13613) );
  ANDN U14549 ( .B(a[101]), .A(n1049), .Z(n13525) );
  XOR U14550 ( .A(b[1]), .B(n13525), .Z(n13527) );
  NANDN U14551 ( .A(b[0]), .B(a[100]), .Z(n13526) );
  NAND U14552 ( .A(n13527), .B(n13526), .Z(n13572) );
  NAND U14553 ( .A(n38490), .B(n13528), .Z(n13530) );
  XNOR U14554 ( .A(n1058), .B(a[73]), .Z(n13663) );
  NANDN U14555 ( .A(n1048), .B(n13663), .Z(n13529) );
  NAND U14556 ( .A(n13530), .B(n13529), .Z(n13569) );
  NANDN U14557 ( .A(n1059), .B(a[69]), .Z(n13570) );
  XNOR U14558 ( .A(n13569), .B(n13570), .Z(n13571) );
  XNOR U14559 ( .A(n13572), .B(n13571), .Z(n13611) );
  NANDN U14560 ( .A(n13531), .B(n38205), .Z(n13533) );
  XNOR U14561 ( .A(b[23]), .B(a[79]), .Z(n13666) );
  OR U14562 ( .A(n13666), .B(n38268), .Z(n13532) );
  NAND U14563 ( .A(n13533), .B(n13532), .Z(n13636) );
  XOR U14564 ( .A(b[7]), .B(a[95]), .Z(n13669) );
  NAND U14565 ( .A(n13669), .B(n36701), .Z(n13536) );
  NAND U14566 ( .A(n13534), .B(n36702), .Z(n13535) );
  NAND U14567 ( .A(n13536), .B(n13535), .Z(n13633) );
  XOR U14568 ( .A(b[25]), .B(a[77]), .Z(n13672) );
  NAND U14569 ( .A(n13672), .B(n38325), .Z(n13539) );
  NAND U14570 ( .A(n13537), .B(n38326), .Z(n13538) );
  AND U14571 ( .A(n13539), .B(n13538), .Z(n13634) );
  XNOR U14572 ( .A(n13633), .B(n13634), .Z(n13635) );
  XNOR U14573 ( .A(n13636), .B(n13635), .Z(n13612) );
  XOR U14574 ( .A(n13611), .B(n13612), .Z(n13614) );
  XNOR U14575 ( .A(n13613), .B(n13614), .Z(n13626) );
  XNOR U14576 ( .A(n13625), .B(n13626), .Z(n13681) );
  XNOR U14577 ( .A(n13682), .B(n13681), .Z(n13684) );
  XNOR U14578 ( .A(n13683), .B(n13684), .Z(n13693) );
  XOR U14579 ( .A(n13694), .B(n13693), .Z(n13696) );
  NAND U14580 ( .A(n13541), .B(n13540), .Z(n13545) );
  NAND U14581 ( .A(n13543), .B(n13542), .Z(n13544) );
  NAND U14582 ( .A(n13545), .B(n13544), .Z(n13688) );
  NAND U14583 ( .A(n13547), .B(n13546), .Z(n13551) );
  NANDN U14584 ( .A(n13549), .B(n13548), .Z(n13550) );
  AND U14585 ( .A(n13551), .B(n13550), .Z(n13687) );
  XNOR U14586 ( .A(n13688), .B(n13687), .Z(n13689) );
  XOR U14587 ( .A(n13690), .B(n13689), .Z(n13566) );
  XOR U14588 ( .A(n13565), .B(n13566), .Z(n13557) );
  XOR U14589 ( .A(n13558), .B(n13557), .Z(n13559) );
  XNOR U14590 ( .A(n13560), .B(n13559), .Z(n13699) );
  XNOR U14591 ( .A(n13699), .B(sreg[325]), .Z(n13701) );
  NAND U14592 ( .A(n13552), .B(sreg[324]), .Z(n13556) );
  OR U14593 ( .A(n13554), .B(n13553), .Z(n13555) );
  AND U14594 ( .A(n13556), .B(n13555), .Z(n13700) );
  XOR U14595 ( .A(n13701), .B(n13700), .Z(c[325]) );
  NAND U14596 ( .A(n13558), .B(n13557), .Z(n13562) );
  NAND U14597 ( .A(n13560), .B(n13559), .Z(n13561) );
  NAND U14598 ( .A(n13562), .B(n13561), .Z(n13707) );
  NANDN U14599 ( .A(n13564), .B(n13563), .Z(n13568) );
  NAND U14600 ( .A(n13566), .B(n13565), .Z(n13567) );
  NAND U14601 ( .A(n13568), .B(n13567), .Z(n13705) );
  NANDN U14602 ( .A(n13570), .B(n13569), .Z(n13574) );
  NANDN U14603 ( .A(n13572), .B(n13571), .Z(n13573) );
  NAND U14604 ( .A(n13574), .B(n13573), .Z(n13779) );
  XNOR U14605 ( .A(b[19]), .B(a[84]), .Z(n13746) );
  NANDN U14606 ( .A(n13746), .B(n37934), .Z(n13577) );
  NANDN U14607 ( .A(n13575), .B(n37935), .Z(n13576) );
  NAND U14608 ( .A(n13577), .B(n13576), .Z(n13815) );
  XOR U14609 ( .A(b[27]), .B(a[76]), .Z(n13749) );
  NAND U14610 ( .A(n38423), .B(n13749), .Z(n13580) );
  NAND U14611 ( .A(n13578), .B(n38424), .Z(n13579) );
  NAND U14612 ( .A(n13580), .B(n13579), .Z(n13812) );
  XNOR U14613 ( .A(b[5]), .B(a[98]), .Z(n13752) );
  NANDN U14614 ( .A(n13752), .B(n36587), .Z(n13583) );
  NANDN U14615 ( .A(n13581), .B(n36588), .Z(n13582) );
  AND U14616 ( .A(n13583), .B(n13582), .Z(n13813) );
  XNOR U14617 ( .A(n13812), .B(n13813), .Z(n13814) );
  XNOR U14618 ( .A(n13815), .B(n13814), .Z(n13776) );
  NAND U14619 ( .A(n13584), .B(n37762), .Z(n13586) );
  XOR U14620 ( .A(b[17]), .B(a[86]), .Z(n13755) );
  NAND U14621 ( .A(n13755), .B(n37764), .Z(n13585) );
  NAND U14622 ( .A(n13586), .B(n13585), .Z(n13730) );
  XNOR U14623 ( .A(b[31]), .B(a[72]), .Z(n13758) );
  NANDN U14624 ( .A(n13758), .B(n38552), .Z(n13589) );
  NANDN U14625 ( .A(n13587), .B(n38553), .Z(n13588) );
  AND U14626 ( .A(n13589), .B(n13588), .Z(n13728) );
  OR U14627 ( .A(n13590), .B(n36105), .Z(n13592) );
  XNOR U14628 ( .A(b[3]), .B(a[100]), .Z(n13761) );
  NANDN U14629 ( .A(n13761), .B(n36107), .Z(n13591) );
  AND U14630 ( .A(n13592), .B(n13591), .Z(n13729) );
  XOR U14631 ( .A(n13730), .B(n13731), .Z(n13777) );
  XOR U14632 ( .A(n13776), .B(n13777), .Z(n13778) );
  XNOR U14633 ( .A(n13779), .B(n13778), .Z(n13824) );
  NANDN U14634 ( .A(n13594), .B(n13593), .Z(n13598) );
  NAND U14635 ( .A(n13596), .B(n13595), .Z(n13597) );
  NAND U14636 ( .A(n13598), .B(n13597), .Z(n13767) );
  NANDN U14637 ( .A(n13600), .B(n13599), .Z(n13604) );
  NAND U14638 ( .A(n13602), .B(n13601), .Z(n13603) );
  NAND U14639 ( .A(n13604), .B(n13603), .Z(n13765) );
  OR U14640 ( .A(n13606), .B(n13605), .Z(n13610) );
  NANDN U14641 ( .A(n13608), .B(n13607), .Z(n13609) );
  NAND U14642 ( .A(n13610), .B(n13609), .Z(n13764) );
  XNOR U14643 ( .A(n13767), .B(n13766), .Z(n13825) );
  XOR U14644 ( .A(n13824), .B(n13825), .Z(n13827) );
  NANDN U14645 ( .A(n13612), .B(n13611), .Z(n13616) );
  OR U14646 ( .A(n13614), .B(n13613), .Z(n13615) );
  NAND U14647 ( .A(n13616), .B(n13615), .Z(n13826) );
  XOR U14648 ( .A(n13827), .B(n13826), .Z(n13844) );
  OR U14649 ( .A(n13618), .B(n13617), .Z(n13622) );
  NAND U14650 ( .A(n13620), .B(n13619), .Z(n13621) );
  NAND U14651 ( .A(n13622), .B(n13621), .Z(n13843) );
  NANDN U14652 ( .A(n13624), .B(n13623), .Z(n13628) );
  NANDN U14653 ( .A(n13626), .B(n13625), .Z(n13627) );
  NAND U14654 ( .A(n13628), .B(n13627), .Z(n13832) );
  NANDN U14655 ( .A(n13634), .B(n13633), .Z(n13638) );
  NAND U14656 ( .A(n13636), .B(n13635), .Z(n13637) );
  NAND U14657 ( .A(n13638), .B(n13637), .Z(n13770) );
  NANDN U14658 ( .A(n13640), .B(n13639), .Z(n13644) );
  NAND U14659 ( .A(n13642), .B(n13641), .Z(n13643) );
  AND U14660 ( .A(n13644), .B(n13643), .Z(n13771) );
  XNOR U14661 ( .A(n13770), .B(n13771), .Z(n13772) );
  XNOR U14662 ( .A(b[9]), .B(a[94]), .Z(n13782) );
  NANDN U14663 ( .A(n13782), .B(n36925), .Z(n13647) );
  NANDN U14664 ( .A(n13645), .B(n36926), .Z(n13646) );
  NAND U14665 ( .A(n13647), .B(n13646), .Z(n13736) );
  XNOR U14666 ( .A(b[15]), .B(a[88]), .Z(n13785) );
  OR U14667 ( .A(n13785), .B(n37665), .Z(n13650) );
  NANDN U14668 ( .A(n13648), .B(n37604), .Z(n13649) );
  AND U14669 ( .A(n13650), .B(n13649), .Z(n13734) );
  XOR U14670 ( .A(b[21]), .B(n15424), .Z(n13788) );
  NANDN U14671 ( .A(n13788), .B(n38101), .Z(n13653) );
  NANDN U14672 ( .A(n13651), .B(n38102), .Z(n13652) );
  AND U14673 ( .A(n13653), .B(n13652), .Z(n13735) );
  XOR U14674 ( .A(n13736), .B(n13737), .Z(n13725) );
  XNOR U14675 ( .A(b[11]), .B(a[92]), .Z(n13791) );
  OR U14676 ( .A(n13791), .B(n37311), .Z(n13656) );
  NANDN U14677 ( .A(n13654), .B(n37218), .Z(n13655) );
  NAND U14678 ( .A(n13656), .B(n13655), .Z(n13723) );
  XOR U14679 ( .A(n1053), .B(a[90]), .Z(n13794) );
  NANDN U14680 ( .A(n13794), .B(n37424), .Z(n13659) );
  NANDN U14681 ( .A(n13657), .B(n37425), .Z(n13658) );
  NAND U14682 ( .A(n13659), .B(n13658), .Z(n13722) );
  XOR U14683 ( .A(n13725), .B(n13724), .Z(n13719) );
  NANDN U14684 ( .A(n1049), .B(a[102]), .Z(n13660) );
  XNOR U14685 ( .A(b[1]), .B(n13660), .Z(n13662) );
  IV U14686 ( .A(a[101]), .Z(n17812) );
  NANDN U14687 ( .A(n17812), .B(n1049), .Z(n13661) );
  AND U14688 ( .A(n13662), .B(n13661), .Z(n13742) );
  NAND U14689 ( .A(n38490), .B(n13663), .Z(n13665) );
  XNOR U14690 ( .A(n1058), .B(a[74]), .Z(n13800) );
  NANDN U14691 ( .A(n1048), .B(n13800), .Z(n13664) );
  NAND U14692 ( .A(n13665), .B(n13664), .Z(n13740) );
  NANDN U14693 ( .A(n1059), .B(a[70]), .Z(n13741) );
  XNOR U14694 ( .A(n13740), .B(n13741), .Z(n13743) );
  XNOR U14695 ( .A(n13742), .B(n13743), .Z(n13717) );
  NANDN U14696 ( .A(n13666), .B(n38205), .Z(n13668) );
  XOR U14697 ( .A(b[23]), .B(n15068), .Z(n13803) );
  OR U14698 ( .A(n13803), .B(n38268), .Z(n13667) );
  NAND U14699 ( .A(n13668), .B(n13667), .Z(n13821) );
  XOR U14700 ( .A(b[7]), .B(a[96]), .Z(n13806) );
  NAND U14701 ( .A(n13806), .B(n36701), .Z(n13671) );
  NAND U14702 ( .A(n13669), .B(n36702), .Z(n13670) );
  NAND U14703 ( .A(n13671), .B(n13670), .Z(n13818) );
  XOR U14704 ( .A(b[25]), .B(a[78]), .Z(n13809) );
  NAND U14705 ( .A(n13809), .B(n38325), .Z(n13674) );
  NAND U14706 ( .A(n13672), .B(n38326), .Z(n13673) );
  AND U14707 ( .A(n13674), .B(n13673), .Z(n13819) );
  XNOR U14708 ( .A(n13818), .B(n13819), .Z(n13820) );
  XOR U14709 ( .A(n13821), .B(n13820), .Z(n13716) );
  XOR U14710 ( .A(n13719), .B(n13718), .Z(n13773) );
  XNOR U14711 ( .A(n13772), .B(n13773), .Z(n13830) );
  XNOR U14712 ( .A(n13831), .B(n13830), .Z(n13833) );
  XNOR U14713 ( .A(n13832), .B(n13833), .Z(n13842) );
  XOR U14714 ( .A(n13843), .B(n13842), .Z(n13845) );
  NANDN U14715 ( .A(n13676), .B(n13675), .Z(n13680) );
  OR U14716 ( .A(n13678), .B(n13677), .Z(n13679) );
  NAND U14717 ( .A(n13680), .B(n13679), .Z(n13836) );
  NAND U14718 ( .A(n13682), .B(n13681), .Z(n13686) );
  NANDN U14719 ( .A(n13684), .B(n13683), .Z(n13685) );
  NAND U14720 ( .A(n13686), .B(n13685), .Z(n13837) );
  XNOR U14721 ( .A(n13836), .B(n13837), .Z(n13838) );
  XOR U14722 ( .A(n13839), .B(n13838), .Z(n13712) );
  NANDN U14723 ( .A(n13688), .B(n13687), .Z(n13692) );
  NAND U14724 ( .A(n13690), .B(n13689), .Z(n13691) );
  NAND U14725 ( .A(n13692), .B(n13691), .Z(n13710) );
  NANDN U14726 ( .A(n13694), .B(n13693), .Z(n13698) );
  OR U14727 ( .A(n13696), .B(n13695), .Z(n13697) );
  NAND U14728 ( .A(n13698), .B(n13697), .Z(n13711) );
  XNOR U14729 ( .A(n13710), .B(n13711), .Z(n13713) );
  XOR U14730 ( .A(n13712), .B(n13713), .Z(n13704) );
  XOR U14731 ( .A(n13705), .B(n13704), .Z(n13706) );
  XNOR U14732 ( .A(n13707), .B(n13706), .Z(n13848) );
  XNOR U14733 ( .A(n13848), .B(sreg[326]), .Z(n13850) );
  NAND U14734 ( .A(n13699), .B(sreg[325]), .Z(n13703) );
  OR U14735 ( .A(n13701), .B(n13700), .Z(n13702) );
  AND U14736 ( .A(n13703), .B(n13702), .Z(n13849) );
  XOR U14737 ( .A(n13850), .B(n13849), .Z(c[326]) );
  NAND U14738 ( .A(n13705), .B(n13704), .Z(n13709) );
  NAND U14739 ( .A(n13707), .B(n13706), .Z(n13708) );
  NAND U14740 ( .A(n13709), .B(n13708), .Z(n13856) );
  NANDN U14741 ( .A(n13711), .B(n13710), .Z(n13715) );
  NAND U14742 ( .A(n13713), .B(n13712), .Z(n13714) );
  NAND U14743 ( .A(n13715), .B(n13714), .Z(n13854) );
  NANDN U14744 ( .A(n13717), .B(n13716), .Z(n13721) );
  NANDN U14745 ( .A(n13719), .B(n13718), .Z(n13720) );
  NAND U14746 ( .A(n13721), .B(n13720), .Z(n13974) );
  OR U14747 ( .A(n13723), .B(n13722), .Z(n13727) );
  NAND U14748 ( .A(n13725), .B(n13724), .Z(n13726) );
  NAND U14749 ( .A(n13727), .B(n13726), .Z(n13913) );
  OR U14750 ( .A(n13729), .B(n13728), .Z(n13733) );
  NANDN U14751 ( .A(n13731), .B(n13730), .Z(n13732) );
  NAND U14752 ( .A(n13733), .B(n13732), .Z(n13912) );
  OR U14753 ( .A(n13735), .B(n13734), .Z(n13739) );
  NANDN U14754 ( .A(n13737), .B(n13736), .Z(n13738) );
  NAND U14755 ( .A(n13739), .B(n13738), .Z(n13911) );
  XOR U14756 ( .A(n13913), .B(n13914), .Z(n13971) );
  NANDN U14757 ( .A(n13741), .B(n13740), .Z(n13745) );
  NAND U14758 ( .A(n13743), .B(n13742), .Z(n13744) );
  NAND U14759 ( .A(n13745), .B(n13744), .Z(n13926) );
  XNOR U14760 ( .A(b[19]), .B(a[85]), .Z(n13869) );
  NANDN U14761 ( .A(n13869), .B(n37934), .Z(n13748) );
  NANDN U14762 ( .A(n13746), .B(n37935), .Z(n13747) );
  NAND U14763 ( .A(n13748), .B(n13747), .Z(n13938) );
  XOR U14764 ( .A(b[27]), .B(a[77]), .Z(n13872) );
  NAND U14765 ( .A(n38423), .B(n13872), .Z(n13751) );
  NAND U14766 ( .A(n13749), .B(n38424), .Z(n13750) );
  NAND U14767 ( .A(n13751), .B(n13750), .Z(n13935) );
  XOR U14768 ( .A(b[5]), .B(n17884), .Z(n13875) );
  NANDN U14769 ( .A(n13875), .B(n36587), .Z(n13754) );
  NANDN U14770 ( .A(n13752), .B(n36588), .Z(n13753) );
  AND U14771 ( .A(n13754), .B(n13753), .Z(n13936) );
  XNOR U14772 ( .A(n13935), .B(n13936), .Z(n13937) );
  XNOR U14773 ( .A(n13938), .B(n13937), .Z(n13924) );
  NAND U14774 ( .A(n13755), .B(n37762), .Z(n13757) );
  XOR U14775 ( .A(b[17]), .B(a[87]), .Z(n13878) );
  NAND U14776 ( .A(n13878), .B(n37764), .Z(n13756) );
  NAND U14777 ( .A(n13757), .B(n13756), .Z(n13896) );
  XNOR U14778 ( .A(b[31]), .B(a[73]), .Z(n13881) );
  NANDN U14779 ( .A(n13881), .B(n38552), .Z(n13760) );
  NANDN U14780 ( .A(n13758), .B(n38553), .Z(n13759) );
  NAND U14781 ( .A(n13760), .B(n13759), .Z(n13893) );
  OR U14782 ( .A(n13761), .B(n36105), .Z(n13763) );
  XOR U14783 ( .A(b[3]), .B(n17812), .Z(n13884) );
  NANDN U14784 ( .A(n13884), .B(n36107), .Z(n13762) );
  AND U14785 ( .A(n13763), .B(n13762), .Z(n13894) );
  XNOR U14786 ( .A(n13893), .B(n13894), .Z(n13895) );
  XOR U14787 ( .A(n13896), .B(n13895), .Z(n13923) );
  XNOR U14788 ( .A(n13924), .B(n13923), .Z(n13925) );
  XNOR U14789 ( .A(n13926), .B(n13925), .Z(n13972) );
  XNOR U14790 ( .A(n13971), .B(n13972), .Z(n13973) );
  XNOR U14791 ( .A(n13974), .B(n13973), .Z(n13992) );
  OR U14792 ( .A(n13765), .B(n13764), .Z(n13769) );
  NAND U14793 ( .A(n13767), .B(n13766), .Z(n13768) );
  NAND U14794 ( .A(n13769), .B(n13768), .Z(n13990) );
  NANDN U14795 ( .A(n13771), .B(n13770), .Z(n13775) );
  NANDN U14796 ( .A(n13773), .B(n13772), .Z(n13774) );
  NAND U14797 ( .A(n13775), .B(n13774), .Z(n13980) );
  OR U14798 ( .A(n13777), .B(n13776), .Z(n13781) );
  NAND U14799 ( .A(n13779), .B(n13778), .Z(n13780) );
  NAND U14800 ( .A(n13781), .B(n13780), .Z(n13977) );
  XNOR U14801 ( .A(b[9]), .B(a[95]), .Z(n13941) );
  NANDN U14802 ( .A(n13941), .B(n36925), .Z(n13784) );
  NANDN U14803 ( .A(n13782), .B(n36926), .Z(n13783) );
  NAND U14804 ( .A(n13784), .B(n13783), .Z(n13901) );
  XNOR U14805 ( .A(b[15]), .B(a[89]), .Z(n13944) );
  OR U14806 ( .A(n13944), .B(n37665), .Z(n13787) );
  NANDN U14807 ( .A(n13785), .B(n37604), .Z(n13786) );
  AND U14808 ( .A(n13787), .B(n13786), .Z(n13899) );
  XOR U14809 ( .A(b[21]), .B(n15562), .Z(n13947) );
  NANDN U14810 ( .A(n13947), .B(n38101), .Z(n13790) );
  NANDN U14811 ( .A(n13788), .B(n38102), .Z(n13789) );
  AND U14812 ( .A(n13790), .B(n13789), .Z(n13900) );
  XOR U14813 ( .A(n13901), .B(n13902), .Z(n13890) );
  XOR U14814 ( .A(b[11]), .B(n17031), .Z(n13950) );
  OR U14815 ( .A(n13950), .B(n37311), .Z(n13793) );
  NANDN U14816 ( .A(n13791), .B(n37218), .Z(n13792) );
  NAND U14817 ( .A(n13793), .B(n13792), .Z(n13888) );
  XOR U14818 ( .A(n1053), .B(a[91]), .Z(n13953) );
  NANDN U14819 ( .A(n13953), .B(n37424), .Z(n13796) );
  NANDN U14820 ( .A(n13794), .B(n37425), .Z(n13795) );
  AND U14821 ( .A(n13796), .B(n13795), .Z(n13887) );
  XNOR U14822 ( .A(n13888), .B(n13887), .Z(n13889) );
  XOR U14823 ( .A(n13890), .B(n13889), .Z(n13908) );
  NANDN U14824 ( .A(n1049), .B(a[103]), .Z(n13797) );
  XNOR U14825 ( .A(b[1]), .B(n13797), .Z(n13799) );
  NANDN U14826 ( .A(b[0]), .B(a[102]), .Z(n13798) );
  AND U14827 ( .A(n13799), .B(n13798), .Z(n13865) );
  NAND U14828 ( .A(n38490), .B(n13800), .Z(n13802) );
  XNOR U14829 ( .A(n1058), .B(a[75]), .Z(n13959) );
  NANDN U14830 ( .A(n1048), .B(n13959), .Z(n13801) );
  NAND U14831 ( .A(n13802), .B(n13801), .Z(n13863) );
  NANDN U14832 ( .A(n1059), .B(a[71]), .Z(n13864) );
  XNOR U14833 ( .A(n13863), .B(n13864), .Z(n13866) );
  XOR U14834 ( .A(n13865), .B(n13866), .Z(n13905) );
  NANDN U14835 ( .A(n13803), .B(n38205), .Z(n13805) );
  XNOR U14836 ( .A(b[23]), .B(a[81]), .Z(n13962) );
  OR U14837 ( .A(n13962), .B(n38268), .Z(n13804) );
  NAND U14838 ( .A(n13805), .B(n13804), .Z(n13932) );
  XOR U14839 ( .A(b[7]), .B(a[97]), .Z(n13965) );
  NAND U14840 ( .A(n13965), .B(n36701), .Z(n13808) );
  NAND U14841 ( .A(n13806), .B(n36702), .Z(n13807) );
  NAND U14842 ( .A(n13808), .B(n13807), .Z(n13929) );
  XOR U14843 ( .A(b[25]), .B(a[79]), .Z(n13968) );
  NAND U14844 ( .A(n13968), .B(n38325), .Z(n13811) );
  NAND U14845 ( .A(n13809), .B(n38326), .Z(n13810) );
  AND U14846 ( .A(n13811), .B(n13810), .Z(n13930) );
  XNOR U14847 ( .A(n13929), .B(n13930), .Z(n13931) );
  XNOR U14848 ( .A(n13932), .B(n13931), .Z(n13906) );
  XNOR U14849 ( .A(n13905), .B(n13906), .Z(n13907) );
  XNOR U14850 ( .A(n13908), .B(n13907), .Z(n13920) );
  NANDN U14851 ( .A(n13813), .B(n13812), .Z(n13817) );
  NAND U14852 ( .A(n13815), .B(n13814), .Z(n13816) );
  NAND U14853 ( .A(n13817), .B(n13816), .Z(n13918) );
  NANDN U14854 ( .A(n13819), .B(n13818), .Z(n13823) );
  NAND U14855 ( .A(n13821), .B(n13820), .Z(n13822) );
  AND U14856 ( .A(n13823), .B(n13822), .Z(n13917) );
  XNOR U14857 ( .A(n13918), .B(n13917), .Z(n13919) );
  XNOR U14858 ( .A(n13920), .B(n13919), .Z(n13978) );
  XNOR U14859 ( .A(n13977), .B(n13978), .Z(n13979) );
  XOR U14860 ( .A(n13980), .B(n13979), .Z(n13989) );
  XNOR U14861 ( .A(n13990), .B(n13989), .Z(n13991) );
  XOR U14862 ( .A(n13992), .B(n13991), .Z(n13986) );
  NANDN U14863 ( .A(n13825), .B(n13824), .Z(n13829) );
  OR U14864 ( .A(n13827), .B(n13826), .Z(n13828) );
  NAND U14865 ( .A(n13829), .B(n13828), .Z(n13983) );
  NAND U14866 ( .A(n13831), .B(n13830), .Z(n13835) );
  NANDN U14867 ( .A(n13833), .B(n13832), .Z(n13834) );
  NAND U14868 ( .A(n13835), .B(n13834), .Z(n13984) );
  XNOR U14869 ( .A(n13983), .B(n13984), .Z(n13985) );
  XNOR U14870 ( .A(n13986), .B(n13985), .Z(n13860) );
  NANDN U14871 ( .A(n13837), .B(n13836), .Z(n13841) );
  NAND U14872 ( .A(n13839), .B(n13838), .Z(n13840) );
  NAND U14873 ( .A(n13841), .B(n13840), .Z(n13857) );
  NANDN U14874 ( .A(n13843), .B(n13842), .Z(n13847) );
  OR U14875 ( .A(n13845), .B(n13844), .Z(n13846) );
  NAND U14876 ( .A(n13847), .B(n13846), .Z(n13858) );
  XNOR U14877 ( .A(n13857), .B(n13858), .Z(n13859) );
  XNOR U14878 ( .A(n13860), .B(n13859), .Z(n13853) );
  XOR U14879 ( .A(n13854), .B(n13853), .Z(n13855) );
  XNOR U14880 ( .A(n13856), .B(n13855), .Z(n13995) );
  XNOR U14881 ( .A(n13995), .B(sreg[327]), .Z(n13997) );
  NAND U14882 ( .A(n13848), .B(sreg[326]), .Z(n13852) );
  OR U14883 ( .A(n13850), .B(n13849), .Z(n13851) );
  AND U14884 ( .A(n13852), .B(n13851), .Z(n13996) );
  XOR U14885 ( .A(n13997), .B(n13996), .Z(c[327]) );
  NANDN U14886 ( .A(n13858), .B(n13857), .Z(n13862) );
  NANDN U14887 ( .A(n13860), .B(n13859), .Z(n13861) );
  NAND U14888 ( .A(n13862), .B(n13861), .Z(n14001) );
  NANDN U14889 ( .A(n13864), .B(n13863), .Z(n13868) );
  NAND U14890 ( .A(n13866), .B(n13865), .Z(n13867) );
  NAND U14891 ( .A(n13868), .B(n13867), .Z(n14075) );
  XNOR U14892 ( .A(b[19]), .B(a[86]), .Z(n14018) );
  NANDN U14893 ( .A(n14018), .B(n37934), .Z(n13871) );
  NANDN U14894 ( .A(n13869), .B(n37935), .Z(n13870) );
  NAND U14895 ( .A(n13871), .B(n13870), .Z(n14085) );
  XOR U14896 ( .A(b[27]), .B(a[78]), .Z(n14021) );
  NAND U14897 ( .A(n38423), .B(n14021), .Z(n13874) );
  NAND U14898 ( .A(n13872), .B(n38424), .Z(n13873) );
  NAND U14899 ( .A(n13874), .B(n13873), .Z(n14082) );
  XNOR U14900 ( .A(b[5]), .B(a[100]), .Z(n14024) );
  NANDN U14901 ( .A(n14024), .B(n36587), .Z(n13877) );
  NANDN U14902 ( .A(n13875), .B(n36588), .Z(n13876) );
  AND U14903 ( .A(n13877), .B(n13876), .Z(n14083) );
  XNOR U14904 ( .A(n14082), .B(n14083), .Z(n14084) );
  XNOR U14905 ( .A(n14085), .B(n14084), .Z(n14073) );
  NAND U14906 ( .A(n13878), .B(n37762), .Z(n13880) );
  XOR U14907 ( .A(b[17]), .B(a[88]), .Z(n14027) );
  NAND U14908 ( .A(n14027), .B(n37764), .Z(n13879) );
  NAND U14909 ( .A(n13880), .B(n13879), .Z(n14045) );
  XNOR U14910 ( .A(b[31]), .B(a[74]), .Z(n14030) );
  NANDN U14911 ( .A(n14030), .B(n38552), .Z(n13883) );
  NANDN U14912 ( .A(n13881), .B(n38553), .Z(n13882) );
  NAND U14913 ( .A(n13883), .B(n13882), .Z(n14042) );
  OR U14914 ( .A(n13884), .B(n36105), .Z(n13886) );
  XNOR U14915 ( .A(b[3]), .B(a[102]), .Z(n14033) );
  NANDN U14916 ( .A(n14033), .B(n36107), .Z(n13885) );
  AND U14917 ( .A(n13886), .B(n13885), .Z(n14043) );
  XNOR U14918 ( .A(n14042), .B(n14043), .Z(n14044) );
  XOR U14919 ( .A(n14045), .B(n14044), .Z(n14072) );
  XNOR U14920 ( .A(n14073), .B(n14072), .Z(n14074) );
  XNOR U14921 ( .A(n14075), .B(n14074), .Z(n14118) );
  NANDN U14922 ( .A(n13888), .B(n13887), .Z(n13892) );
  NAND U14923 ( .A(n13890), .B(n13889), .Z(n13891) );
  NAND U14924 ( .A(n13892), .B(n13891), .Z(n14063) );
  NANDN U14925 ( .A(n13894), .B(n13893), .Z(n13898) );
  NAND U14926 ( .A(n13896), .B(n13895), .Z(n13897) );
  NAND U14927 ( .A(n13898), .B(n13897), .Z(n14061) );
  OR U14928 ( .A(n13900), .B(n13899), .Z(n13904) );
  NANDN U14929 ( .A(n13902), .B(n13901), .Z(n13903) );
  NAND U14930 ( .A(n13904), .B(n13903), .Z(n14060) );
  XNOR U14931 ( .A(n14063), .B(n14062), .Z(n14119) );
  XOR U14932 ( .A(n14118), .B(n14119), .Z(n14121) );
  NANDN U14933 ( .A(n13906), .B(n13905), .Z(n13910) );
  NANDN U14934 ( .A(n13908), .B(n13907), .Z(n13909) );
  NAND U14935 ( .A(n13910), .B(n13909), .Z(n14120) );
  XOR U14936 ( .A(n14121), .B(n14120), .Z(n14136) );
  OR U14937 ( .A(n13912), .B(n13911), .Z(n13916) );
  NANDN U14938 ( .A(n13914), .B(n13913), .Z(n13915) );
  NAND U14939 ( .A(n13916), .B(n13915), .Z(n14135) );
  NANDN U14940 ( .A(n13918), .B(n13917), .Z(n13922) );
  NANDN U14941 ( .A(n13920), .B(n13919), .Z(n13921) );
  NAND U14942 ( .A(n13922), .B(n13921), .Z(n14126) );
  NANDN U14943 ( .A(n13924), .B(n13923), .Z(n13928) );
  NAND U14944 ( .A(n13926), .B(n13925), .Z(n13927) );
  NAND U14945 ( .A(n13928), .B(n13927), .Z(n14125) );
  NANDN U14946 ( .A(n13930), .B(n13929), .Z(n13934) );
  NAND U14947 ( .A(n13932), .B(n13931), .Z(n13933) );
  NAND U14948 ( .A(n13934), .B(n13933), .Z(n14066) );
  NANDN U14949 ( .A(n13936), .B(n13935), .Z(n13940) );
  NAND U14950 ( .A(n13938), .B(n13937), .Z(n13939) );
  AND U14951 ( .A(n13940), .B(n13939), .Z(n14067) );
  XNOR U14952 ( .A(n14066), .B(n14067), .Z(n14068) );
  XNOR U14953 ( .A(n1052), .B(a[96]), .Z(n14088) );
  NAND U14954 ( .A(n36925), .B(n14088), .Z(n13943) );
  NANDN U14955 ( .A(n13941), .B(n36926), .Z(n13942) );
  NAND U14956 ( .A(n13943), .B(n13942), .Z(n14050) );
  XNOR U14957 ( .A(b[15]), .B(a[90]), .Z(n14091) );
  OR U14958 ( .A(n14091), .B(n37665), .Z(n13946) );
  NANDN U14959 ( .A(n13944), .B(n37604), .Z(n13945) );
  AND U14960 ( .A(n13946), .B(n13945), .Z(n14048) );
  XNOR U14961 ( .A(n1056), .B(a[84]), .Z(n14094) );
  NAND U14962 ( .A(n14094), .B(n38101), .Z(n13949) );
  NANDN U14963 ( .A(n13947), .B(n38102), .Z(n13948) );
  AND U14964 ( .A(n13949), .B(n13948), .Z(n14049) );
  XOR U14965 ( .A(n14050), .B(n14051), .Z(n14039) );
  XNOR U14966 ( .A(b[11]), .B(a[94]), .Z(n14097) );
  OR U14967 ( .A(n14097), .B(n37311), .Z(n13952) );
  NANDN U14968 ( .A(n13950), .B(n37218), .Z(n13951) );
  NAND U14969 ( .A(n13952), .B(n13951), .Z(n14037) );
  XOR U14970 ( .A(n1053), .B(a[92]), .Z(n14100) );
  NANDN U14971 ( .A(n14100), .B(n37424), .Z(n13955) );
  NANDN U14972 ( .A(n13953), .B(n37425), .Z(n13954) );
  AND U14973 ( .A(n13955), .B(n13954), .Z(n14036) );
  XNOR U14974 ( .A(n14037), .B(n14036), .Z(n14038) );
  XOR U14975 ( .A(n14039), .B(n14038), .Z(n14056) );
  NANDN U14976 ( .A(n1049), .B(a[104]), .Z(n13956) );
  XNOR U14977 ( .A(b[1]), .B(n13956), .Z(n13958) );
  NANDN U14978 ( .A(b[0]), .B(a[103]), .Z(n13957) );
  AND U14979 ( .A(n13958), .B(n13957), .Z(n14014) );
  NAND U14980 ( .A(n38490), .B(n13959), .Z(n13961) );
  XNOR U14981 ( .A(n1058), .B(a[76]), .Z(n14103) );
  NANDN U14982 ( .A(n1048), .B(n14103), .Z(n13960) );
  NAND U14983 ( .A(n13961), .B(n13960), .Z(n14012) );
  NANDN U14984 ( .A(n1059), .B(a[72]), .Z(n14013) );
  XNOR U14985 ( .A(n14012), .B(n14013), .Z(n14015) );
  XOR U14986 ( .A(n14014), .B(n14015), .Z(n14054) );
  NANDN U14987 ( .A(n13962), .B(n38205), .Z(n13964) );
  XOR U14988 ( .A(b[23]), .B(n15424), .Z(n14109) );
  OR U14989 ( .A(n14109), .B(n38268), .Z(n13963) );
  NAND U14990 ( .A(n13964), .B(n13963), .Z(n14079) );
  XOR U14991 ( .A(b[7]), .B(a[98]), .Z(n14112) );
  NAND U14992 ( .A(n14112), .B(n36701), .Z(n13967) );
  NAND U14993 ( .A(n13965), .B(n36702), .Z(n13966) );
  NAND U14994 ( .A(n13967), .B(n13966), .Z(n14076) );
  XNOR U14995 ( .A(b[25]), .B(a[80]), .Z(n14115) );
  NANDN U14996 ( .A(n14115), .B(n38325), .Z(n13970) );
  NAND U14997 ( .A(n13968), .B(n38326), .Z(n13969) );
  AND U14998 ( .A(n13970), .B(n13969), .Z(n14077) );
  XNOR U14999 ( .A(n14076), .B(n14077), .Z(n14078) );
  XNOR U15000 ( .A(n14079), .B(n14078), .Z(n14055) );
  XOR U15001 ( .A(n14054), .B(n14055), .Z(n14057) );
  XNOR U15002 ( .A(n14056), .B(n14057), .Z(n14069) );
  XNOR U15003 ( .A(n14068), .B(n14069), .Z(n14124) );
  XNOR U15004 ( .A(n14125), .B(n14124), .Z(n14127) );
  XOR U15005 ( .A(n14126), .B(n14127), .Z(n14134) );
  XOR U15006 ( .A(n14135), .B(n14134), .Z(n14137) );
  NANDN U15007 ( .A(n13972), .B(n13971), .Z(n13976) );
  NAND U15008 ( .A(n13974), .B(n13973), .Z(n13975) );
  NAND U15009 ( .A(n13976), .B(n13975), .Z(n14129) );
  NANDN U15010 ( .A(n13978), .B(n13977), .Z(n13982) );
  NAND U15011 ( .A(n13980), .B(n13979), .Z(n13981) );
  AND U15012 ( .A(n13982), .B(n13981), .Z(n14128) );
  XNOR U15013 ( .A(n14129), .B(n14128), .Z(n14130) );
  XOR U15014 ( .A(n14131), .B(n14130), .Z(n14008) );
  NANDN U15015 ( .A(n13984), .B(n13983), .Z(n13988) );
  NAND U15016 ( .A(n13986), .B(n13985), .Z(n13987) );
  NAND U15017 ( .A(n13988), .B(n13987), .Z(n14006) );
  NANDN U15018 ( .A(n13990), .B(n13989), .Z(n13994) );
  NANDN U15019 ( .A(n13992), .B(n13991), .Z(n13993) );
  NAND U15020 ( .A(n13994), .B(n13993), .Z(n14007) );
  XNOR U15021 ( .A(n14006), .B(n14007), .Z(n14009) );
  XOR U15022 ( .A(n14008), .B(n14009), .Z(n14000) );
  XOR U15023 ( .A(n14001), .B(n14000), .Z(n14002) );
  XNOR U15024 ( .A(n14003), .B(n14002), .Z(n14140) );
  XNOR U15025 ( .A(n14140), .B(sreg[328]), .Z(n14142) );
  NAND U15026 ( .A(n13995), .B(sreg[327]), .Z(n13999) );
  OR U15027 ( .A(n13997), .B(n13996), .Z(n13998) );
  AND U15028 ( .A(n13999), .B(n13998), .Z(n14141) );
  XOR U15029 ( .A(n14142), .B(n14141), .Z(c[328]) );
  NAND U15030 ( .A(n14001), .B(n14000), .Z(n14005) );
  NAND U15031 ( .A(n14003), .B(n14002), .Z(n14004) );
  NAND U15032 ( .A(n14005), .B(n14004), .Z(n14148) );
  NANDN U15033 ( .A(n14007), .B(n14006), .Z(n14011) );
  NAND U15034 ( .A(n14009), .B(n14008), .Z(n14010) );
  NAND U15035 ( .A(n14011), .B(n14010), .Z(n14146) );
  NANDN U15036 ( .A(n14013), .B(n14012), .Z(n14017) );
  NAND U15037 ( .A(n14015), .B(n14014), .Z(n14016) );
  NAND U15038 ( .A(n14017), .B(n14016), .Z(n14218) );
  XNOR U15039 ( .A(b[19]), .B(a[87]), .Z(n14163) );
  NANDN U15040 ( .A(n14163), .B(n37934), .Z(n14020) );
  NANDN U15041 ( .A(n14018), .B(n37935), .Z(n14019) );
  NAND U15042 ( .A(n14020), .B(n14019), .Z(n14228) );
  XOR U15043 ( .A(b[27]), .B(a[79]), .Z(n14166) );
  NAND U15044 ( .A(n38423), .B(n14166), .Z(n14023) );
  NAND U15045 ( .A(n14021), .B(n38424), .Z(n14022) );
  NAND U15046 ( .A(n14023), .B(n14022), .Z(n14225) );
  XOR U15047 ( .A(b[5]), .B(n17812), .Z(n14169) );
  NANDN U15048 ( .A(n14169), .B(n36587), .Z(n14026) );
  NANDN U15049 ( .A(n14024), .B(n36588), .Z(n14025) );
  AND U15050 ( .A(n14026), .B(n14025), .Z(n14226) );
  XNOR U15051 ( .A(n14225), .B(n14226), .Z(n14227) );
  XNOR U15052 ( .A(n14228), .B(n14227), .Z(n14216) );
  NAND U15053 ( .A(n14027), .B(n37762), .Z(n14029) );
  XOR U15054 ( .A(b[17]), .B(a[89]), .Z(n14172) );
  NAND U15055 ( .A(n14172), .B(n37764), .Z(n14028) );
  NAND U15056 ( .A(n14029), .B(n14028), .Z(n14190) );
  XNOR U15057 ( .A(b[31]), .B(a[75]), .Z(n14175) );
  NANDN U15058 ( .A(n14175), .B(n38552), .Z(n14032) );
  NANDN U15059 ( .A(n14030), .B(n38553), .Z(n14031) );
  NAND U15060 ( .A(n14032), .B(n14031), .Z(n14187) );
  OR U15061 ( .A(n14033), .B(n36105), .Z(n14035) );
  XNOR U15062 ( .A(b[3]), .B(a[103]), .Z(n14178) );
  NANDN U15063 ( .A(n14178), .B(n36107), .Z(n14034) );
  AND U15064 ( .A(n14035), .B(n14034), .Z(n14188) );
  XNOR U15065 ( .A(n14187), .B(n14188), .Z(n14189) );
  XOR U15066 ( .A(n14190), .B(n14189), .Z(n14215) );
  XNOR U15067 ( .A(n14216), .B(n14215), .Z(n14217) );
  XNOR U15068 ( .A(n14218), .B(n14217), .Z(n14261) );
  NANDN U15069 ( .A(n14037), .B(n14036), .Z(n14041) );
  NAND U15070 ( .A(n14039), .B(n14038), .Z(n14040) );
  NAND U15071 ( .A(n14041), .B(n14040), .Z(n14206) );
  NANDN U15072 ( .A(n14043), .B(n14042), .Z(n14047) );
  NAND U15073 ( .A(n14045), .B(n14044), .Z(n14046) );
  NAND U15074 ( .A(n14047), .B(n14046), .Z(n14204) );
  OR U15075 ( .A(n14049), .B(n14048), .Z(n14053) );
  NANDN U15076 ( .A(n14051), .B(n14050), .Z(n14052) );
  NAND U15077 ( .A(n14053), .B(n14052), .Z(n14203) );
  XNOR U15078 ( .A(n14206), .B(n14205), .Z(n14262) );
  XOR U15079 ( .A(n14261), .B(n14262), .Z(n14264) );
  NANDN U15080 ( .A(n14055), .B(n14054), .Z(n14059) );
  OR U15081 ( .A(n14057), .B(n14056), .Z(n14058) );
  NAND U15082 ( .A(n14059), .B(n14058), .Z(n14263) );
  XOR U15083 ( .A(n14264), .B(n14263), .Z(n14281) );
  OR U15084 ( .A(n14061), .B(n14060), .Z(n14065) );
  NAND U15085 ( .A(n14063), .B(n14062), .Z(n14064) );
  NAND U15086 ( .A(n14065), .B(n14064), .Z(n14280) );
  NANDN U15087 ( .A(n14067), .B(n14066), .Z(n14071) );
  NANDN U15088 ( .A(n14069), .B(n14068), .Z(n14070) );
  NAND U15089 ( .A(n14071), .B(n14070), .Z(n14269) );
  NANDN U15090 ( .A(n14077), .B(n14076), .Z(n14081) );
  NAND U15091 ( .A(n14079), .B(n14078), .Z(n14080) );
  NAND U15092 ( .A(n14081), .B(n14080), .Z(n14209) );
  NANDN U15093 ( .A(n14083), .B(n14082), .Z(n14087) );
  NAND U15094 ( .A(n14085), .B(n14084), .Z(n14086) );
  AND U15095 ( .A(n14087), .B(n14086), .Z(n14210) );
  XNOR U15096 ( .A(n14209), .B(n14210), .Z(n14211) );
  XNOR U15097 ( .A(b[9]), .B(a[97]), .Z(n14231) );
  NANDN U15098 ( .A(n14231), .B(n36925), .Z(n14090) );
  NAND U15099 ( .A(n36926), .B(n14088), .Z(n14089) );
  NAND U15100 ( .A(n14090), .B(n14089), .Z(n14195) );
  XNOR U15101 ( .A(n1054), .B(a[91]), .Z(n14234) );
  NANDN U15102 ( .A(n37665), .B(n14234), .Z(n14093) );
  NANDN U15103 ( .A(n14091), .B(n37604), .Z(n14092) );
  NAND U15104 ( .A(n14093), .B(n14092), .Z(n14193) );
  XNOR U15105 ( .A(b[21]), .B(a[85]), .Z(n14237) );
  NANDN U15106 ( .A(n14237), .B(n38101), .Z(n14096) );
  NAND U15107 ( .A(n38102), .B(n14094), .Z(n14095) );
  NAND U15108 ( .A(n14096), .B(n14095), .Z(n14194) );
  XNOR U15109 ( .A(n14193), .B(n14194), .Z(n14196) );
  XOR U15110 ( .A(n14195), .B(n14196), .Z(n14184) );
  XNOR U15111 ( .A(b[11]), .B(a[95]), .Z(n14240) );
  OR U15112 ( .A(n14240), .B(n37311), .Z(n14099) );
  NANDN U15113 ( .A(n14097), .B(n37218), .Z(n14098) );
  NAND U15114 ( .A(n14099), .B(n14098), .Z(n14182) );
  XOR U15115 ( .A(n1053), .B(a[93]), .Z(n14243) );
  NANDN U15116 ( .A(n14243), .B(n37424), .Z(n14102) );
  NANDN U15117 ( .A(n14100), .B(n37425), .Z(n14101) );
  AND U15118 ( .A(n14102), .B(n14101), .Z(n14181) );
  XNOR U15119 ( .A(n14182), .B(n14181), .Z(n14183) );
  XNOR U15120 ( .A(n14184), .B(n14183), .Z(n14200) );
  NAND U15121 ( .A(n38490), .B(n14103), .Z(n14105) );
  XNOR U15122 ( .A(n1058), .B(a[77]), .Z(n14249) );
  NANDN U15123 ( .A(n1048), .B(n14249), .Z(n14104) );
  NAND U15124 ( .A(n14105), .B(n14104), .Z(n14157) );
  NANDN U15125 ( .A(n1059), .B(a[73]), .Z(n14158) );
  XNOR U15126 ( .A(n14157), .B(n14158), .Z(n14160) );
  NANDN U15127 ( .A(n1049), .B(a[105]), .Z(n14106) );
  XNOR U15128 ( .A(b[1]), .B(n14106), .Z(n14108) );
  NANDN U15129 ( .A(b[0]), .B(a[104]), .Z(n14107) );
  AND U15130 ( .A(n14108), .B(n14107), .Z(n14159) );
  XNOR U15131 ( .A(n14160), .B(n14159), .Z(n14198) );
  NANDN U15132 ( .A(n14109), .B(n38205), .Z(n14111) );
  XOR U15133 ( .A(b[23]), .B(n15562), .Z(n14252) );
  OR U15134 ( .A(n14252), .B(n38268), .Z(n14110) );
  NAND U15135 ( .A(n14111), .B(n14110), .Z(n14222) );
  XNOR U15136 ( .A(b[7]), .B(a[99]), .Z(n14255) );
  NANDN U15137 ( .A(n14255), .B(n36701), .Z(n14114) );
  NAND U15138 ( .A(n14112), .B(n36702), .Z(n14113) );
  NAND U15139 ( .A(n14114), .B(n14113), .Z(n14219) );
  XOR U15140 ( .A(b[25]), .B(a[81]), .Z(n14258) );
  NAND U15141 ( .A(n14258), .B(n38325), .Z(n14117) );
  NANDN U15142 ( .A(n14115), .B(n38326), .Z(n14116) );
  AND U15143 ( .A(n14117), .B(n14116), .Z(n14220) );
  XNOR U15144 ( .A(n14219), .B(n14220), .Z(n14221) );
  XOR U15145 ( .A(n14222), .B(n14221), .Z(n14197) );
  XOR U15146 ( .A(n14200), .B(n14199), .Z(n14212) );
  XOR U15147 ( .A(n14211), .B(n14212), .Z(n14267) );
  XNOR U15148 ( .A(n14268), .B(n14267), .Z(n14270) );
  XNOR U15149 ( .A(n14269), .B(n14270), .Z(n14279) );
  XOR U15150 ( .A(n14280), .B(n14279), .Z(n14282) );
  NANDN U15151 ( .A(n14119), .B(n14118), .Z(n14123) );
  OR U15152 ( .A(n14121), .B(n14120), .Z(n14122) );
  NAND U15153 ( .A(n14123), .B(n14122), .Z(n14273) );
  XNOR U15154 ( .A(n14273), .B(n14274), .Z(n14275) );
  XOR U15155 ( .A(n14276), .B(n14275), .Z(n14153) );
  NANDN U15156 ( .A(n14129), .B(n14128), .Z(n14133) );
  NAND U15157 ( .A(n14131), .B(n14130), .Z(n14132) );
  NAND U15158 ( .A(n14133), .B(n14132), .Z(n14151) );
  NANDN U15159 ( .A(n14135), .B(n14134), .Z(n14139) );
  OR U15160 ( .A(n14137), .B(n14136), .Z(n14138) );
  NAND U15161 ( .A(n14139), .B(n14138), .Z(n14152) );
  XNOR U15162 ( .A(n14151), .B(n14152), .Z(n14154) );
  XOR U15163 ( .A(n14153), .B(n14154), .Z(n14145) );
  XOR U15164 ( .A(n14146), .B(n14145), .Z(n14147) );
  XNOR U15165 ( .A(n14148), .B(n14147), .Z(n14285) );
  XNOR U15166 ( .A(n14285), .B(sreg[329]), .Z(n14287) );
  NAND U15167 ( .A(n14140), .B(sreg[328]), .Z(n14144) );
  OR U15168 ( .A(n14142), .B(n14141), .Z(n14143) );
  AND U15169 ( .A(n14144), .B(n14143), .Z(n14286) );
  XOR U15170 ( .A(n14287), .B(n14286), .Z(c[329]) );
  NAND U15171 ( .A(n14146), .B(n14145), .Z(n14150) );
  NAND U15172 ( .A(n14148), .B(n14147), .Z(n14149) );
  NAND U15173 ( .A(n14150), .B(n14149), .Z(n14293) );
  NANDN U15174 ( .A(n14152), .B(n14151), .Z(n14156) );
  NAND U15175 ( .A(n14154), .B(n14153), .Z(n14155) );
  NAND U15176 ( .A(n14156), .B(n14155), .Z(n14291) );
  NANDN U15177 ( .A(n14158), .B(n14157), .Z(n14162) );
  NAND U15178 ( .A(n14160), .B(n14159), .Z(n14161) );
  NAND U15179 ( .A(n14162), .B(n14161), .Z(n14373) );
  XNOR U15180 ( .A(b[19]), .B(a[88]), .Z(n14318) );
  NANDN U15181 ( .A(n14318), .B(n37934), .Z(n14165) );
  NANDN U15182 ( .A(n14163), .B(n37935), .Z(n14164) );
  NAND U15183 ( .A(n14165), .B(n14164), .Z(n14383) );
  XNOR U15184 ( .A(b[27]), .B(a[80]), .Z(n14321) );
  NANDN U15185 ( .A(n14321), .B(n38423), .Z(n14168) );
  NAND U15186 ( .A(n14166), .B(n38424), .Z(n14167) );
  NAND U15187 ( .A(n14168), .B(n14167), .Z(n14380) );
  XNOR U15188 ( .A(b[5]), .B(a[102]), .Z(n14324) );
  NANDN U15189 ( .A(n14324), .B(n36587), .Z(n14171) );
  NANDN U15190 ( .A(n14169), .B(n36588), .Z(n14170) );
  AND U15191 ( .A(n14171), .B(n14170), .Z(n14381) );
  XNOR U15192 ( .A(n14380), .B(n14381), .Z(n14382) );
  XNOR U15193 ( .A(n14383), .B(n14382), .Z(n14371) );
  NAND U15194 ( .A(n14172), .B(n37762), .Z(n14174) );
  XOR U15195 ( .A(b[17]), .B(a[90]), .Z(n14327) );
  NAND U15196 ( .A(n14327), .B(n37764), .Z(n14173) );
  NAND U15197 ( .A(n14174), .B(n14173), .Z(n14345) );
  XNOR U15198 ( .A(b[31]), .B(a[76]), .Z(n14330) );
  NANDN U15199 ( .A(n14330), .B(n38552), .Z(n14177) );
  NANDN U15200 ( .A(n14175), .B(n38553), .Z(n14176) );
  NAND U15201 ( .A(n14177), .B(n14176), .Z(n14342) );
  OR U15202 ( .A(n14178), .B(n36105), .Z(n14180) );
  XNOR U15203 ( .A(b[3]), .B(a[104]), .Z(n14333) );
  NANDN U15204 ( .A(n14333), .B(n36107), .Z(n14179) );
  AND U15205 ( .A(n14180), .B(n14179), .Z(n14343) );
  XNOR U15206 ( .A(n14342), .B(n14343), .Z(n14344) );
  XOR U15207 ( .A(n14345), .B(n14344), .Z(n14370) );
  XNOR U15208 ( .A(n14371), .B(n14370), .Z(n14372) );
  XNOR U15209 ( .A(n14373), .B(n14372), .Z(n14309) );
  NANDN U15210 ( .A(n14182), .B(n14181), .Z(n14186) );
  NAND U15211 ( .A(n14184), .B(n14183), .Z(n14185) );
  NAND U15212 ( .A(n14186), .B(n14185), .Z(n14362) );
  NANDN U15213 ( .A(n14188), .B(n14187), .Z(n14192) );
  NAND U15214 ( .A(n14190), .B(n14189), .Z(n14191) );
  NAND U15215 ( .A(n14192), .B(n14191), .Z(n14361) );
  XNOR U15216 ( .A(n14361), .B(n14360), .Z(n14363) );
  XOR U15217 ( .A(n14362), .B(n14363), .Z(n14308) );
  XOR U15218 ( .A(n14309), .B(n14308), .Z(n14310) );
  NANDN U15219 ( .A(n14198), .B(n14197), .Z(n14202) );
  NAND U15220 ( .A(n14200), .B(n14199), .Z(n14201) );
  NAND U15221 ( .A(n14202), .B(n14201), .Z(n14311) );
  XNOR U15222 ( .A(n14310), .B(n14311), .Z(n14424) );
  OR U15223 ( .A(n14204), .B(n14203), .Z(n14208) );
  NAND U15224 ( .A(n14206), .B(n14205), .Z(n14207) );
  NAND U15225 ( .A(n14208), .B(n14207), .Z(n14423) );
  NANDN U15226 ( .A(n14210), .B(n14209), .Z(n14214) );
  NAND U15227 ( .A(n14212), .B(n14211), .Z(n14213) );
  NAND U15228 ( .A(n14214), .B(n14213), .Z(n14304) );
  NANDN U15229 ( .A(n14220), .B(n14219), .Z(n14224) );
  NAND U15230 ( .A(n14222), .B(n14221), .Z(n14223) );
  NAND U15231 ( .A(n14224), .B(n14223), .Z(n14364) );
  NANDN U15232 ( .A(n14226), .B(n14225), .Z(n14230) );
  NAND U15233 ( .A(n14228), .B(n14227), .Z(n14229) );
  AND U15234 ( .A(n14230), .B(n14229), .Z(n14365) );
  XNOR U15235 ( .A(n14364), .B(n14365), .Z(n14366) );
  XNOR U15236 ( .A(b[9]), .B(a[98]), .Z(n14386) );
  NANDN U15237 ( .A(n14386), .B(n36925), .Z(n14233) );
  NANDN U15238 ( .A(n14231), .B(n36926), .Z(n14232) );
  NAND U15239 ( .A(n14233), .B(n14232), .Z(n14356) );
  XNOR U15240 ( .A(b[15]), .B(a[92]), .Z(n14389) );
  OR U15241 ( .A(n14389), .B(n37665), .Z(n14236) );
  NAND U15242 ( .A(n14234), .B(n37604), .Z(n14235) );
  AND U15243 ( .A(n14236), .B(n14235), .Z(n14354) );
  XNOR U15244 ( .A(b[21]), .B(a[86]), .Z(n14392) );
  NANDN U15245 ( .A(n14392), .B(n38101), .Z(n14239) );
  NANDN U15246 ( .A(n14237), .B(n38102), .Z(n14238) );
  AND U15247 ( .A(n14239), .B(n14238), .Z(n14355) );
  XOR U15248 ( .A(n14356), .B(n14357), .Z(n14351) );
  XNOR U15249 ( .A(b[11]), .B(a[96]), .Z(n14395) );
  OR U15250 ( .A(n14395), .B(n37311), .Z(n14242) );
  NANDN U15251 ( .A(n14240), .B(n37218), .Z(n14241) );
  NAND U15252 ( .A(n14242), .B(n14241), .Z(n14349) );
  XOR U15253 ( .A(n1053), .B(a[94]), .Z(n14398) );
  NANDN U15254 ( .A(n14398), .B(n37424), .Z(n14245) );
  NANDN U15255 ( .A(n14243), .B(n37425), .Z(n14244) );
  AND U15256 ( .A(n14245), .B(n14244), .Z(n14348) );
  XNOR U15257 ( .A(n14349), .B(n14348), .Z(n14350) );
  XOR U15258 ( .A(n14351), .B(n14350), .Z(n14338) );
  NANDN U15259 ( .A(n1049), .B(a[106]), .Z(n14246) );
  XNOR U15260 ( .A(b[1]), .B(n14246), .Z(n14248) );
  NANDN U15261 ( .A(b[0]), .B(a[105]), .Z(n14247) );
  AND U15262 ( .A(n14248), .B(n14247), .Z(n14314) );
  NAND U15263 ( .A(n38490), .B(n14249), .Z(n14251) );
  XNOR U15264 ( .A(n1058), .B(a[78]), .Z(n14404) );
  NANDN U15265 ( .A(n1048), .B(n14404), .Z(n14250) );
  NAND U15266 ( .A(n14251), .B(n14250), .Z(n14312) );
  NANDN U15267 ( .A(n1059), .B(a[74]), .Z(n14313) );
  XNOR U15268 ( .A(n14312), .B(n14313), .Z(n14315) );
  XOR U15269 ( .A(n14314), .B(n14315), .Z(n14336) );
  NANDN U15270 ( .A(n14252), .B(n38205), .Z(n14254) );
  XNOR U15271 ( .A(b[23]), .B(a[84]), .Z(n14407) );
  OR U15272 ( .A(n14407), .B(n38268), .Z(n14253) );
  NAND U15273 ( .A(n14254), .B(n14253), .Z(n14377) );
  XOR U15274 ( .A(b[7]), .B(a[100]), .Z(n14410) );
  NAND U15275 ( .A(n14410), .B(n36701), .Z(n14257) );
  NANDN U15276 ( .A(n14255), .B(n36702), .Z(n14256) );
  NAND U15277 ( .A(n14257), .B(n14256), .Z(n14374) );
  XNOR U15278 ( .A(b[25]), .B(a[82]), .Z(n14413) );
  NANDN U15279 ( .A(n14413), .B(n38325), .Z(n14260) );
  NAND U15280 ( .A(n14258), .B(n38326), .Z(n14259) );
  AND U15281 ( .A(n14260), .B(n14259), .Z(n14375) );
  XNOR U15282 ( .A(n14374), .B(n14375), .Z(n14376) );
  XNOR U15283 ( .A(n14377), .B(n14376), .Z(n14337) );
  XOR U15284 ( .A(n14336), .B(n14337), .Z(n14339) );
  XNOR U15285 ( .A(n14338), .B(n14339), .Z(n14367) );
  XNOR U15286 ( .A(n14366), .B(n14367), .Z(n14302) );
  XNOR U15287 ( .A(n14303), .B(n14302), .Z(n14305) );
  XNOR U15288 ( .A(n14304), .B(n14305), .Z(n14422) );
  XOR U15289 ( .A(n14423), .B(n14422), .Z(n14425) );
  NANDN U15290 ( .A(n14262), .B(n14261), .Z(n14266) );
  OR U15291 ( .A(n14264), .B(n14263), .Z(n14265) );
  NAND U15292 ( .A(n14266), .B(n14265), .Z(n14416) );
  NAND U15293 ( .A(n14268), .B(n14267), .Z(n14272) );
  NANDN U15294 ( .A(n14270), .B(n14269), .Z(n14271) );
  NAND U15295 ( .A(n14272), .B(n14271), .Z(n14417) );
  XNOR U15296 ( .A(n14416), .B(n14417), .Z(n14418) );
  XOR U15297 ( .A(n14419), .B(n14418), .Z(n14298) );
  NANDN U15298 ( .A(n14274), .B(n14273), .Z(n14278) );
  NAND U15299 ( .A(n14276), .B(n14275), .Z(n14277) );
  NAND U15300 ( .A(n14278), .B(n14277), .Z(n14296) );
  NANDN U15301 ( .A(n14280), .B(n14279), .Z(n14284) );
  OR U15302 ( .A(n14282), .B(n14281), .Z(n14283) );
  NAND U15303 ( .A(n14284), .B(n14283), .Z(n14297) );
  XNOR U15304 ( .A(n14296), .B(n14297), .Z(n14299) );
  XOR U15305 ( .A(n14298), .B(n14299), .Z(n14290) );
  XOR U15306 ( .A(n14291), .B(n14290), .Z(n14292) );
  XNOR U15307 ( .A(n14293), .B(n14292), .Z(n14428) );
  XNOR U15308 ( .A(n14428), .B(sreg[330]), .Z(n14430) );
  NAND U15309 ( .A(n14285), .B(sreg[329]), .Z(n14289) );
  OR U15310 ( .A(n14287), .B(n14286), .Z(n14288) );
  AND U15311 ( .A(n14289), .B(n14288), .Z(n14429) );
  XOR U15312 ( .A(n14430), .B(n14429), .Z(c[330]) );
  NAND U15313 ( .A(n14291), .B(n14290), .Z(n14295) );
  NAND U15314 ( .A(n14293), .B(n14292), .Z(n14294) );
  NAND U15315 ( .A(n14295), .B(n14294), .Z(n14436) );
  NANDN U15316 ( .A(n14297), .B(n14296), .Z(n14301) );
  NAND U15317 ( .A(n14299), .B(n14298), .Z(n14300) );
  NAND U15318 ( .A(n14301), .B(n14300), .Z(n14433) );
  NAND U15319 ( .A(n14303), .B(n14302), .Z(n14307) );
  NANDN U15320 ( .A(n14305), .B(n14304), .Z(n14306) );
  NAND U15321 ( .A(n14307), .B(n14306), .Z(n14565) );
  XNOR U15322 ( .A(n14565), .B(n14566), .Z(n14567) );
  NANDN U15323 ( .A(n14313), .B(n14312), .Z(n14317) );
  NAND U15324 ( .A(n14315), .B(n14314), .Z(n14316) );
  NAND U15325 ( .A(n14317), .B(n14316), .Z(n14520) );
  XNOR U15326 ( .A(b[19]), .B(a[89]), .Z(n14487) );
  NANDN U15327 ( .A(n14487), .B(n37934), .Z(n14320) );
  NANDN U15328 ( .A(n14318), .B(n37935), .Z(n14319) );
  NAND U15329 ( .A(n14320), .B(n14319), .Z(n14532) );
  XOR U15330 ( .A(b[27]), .B(a[81]), .Z(n14490) );
  NAND U15331 ( .A(n38423), .B(n14490), .Z(n14323) );
  NANDN U15332 ( .A(n14321), .B(n38424), .Z(n14322) );
  NAND U15333 ( .A(n14323), .B(n14322), .Z(n14529) );
  XNOR U15334 ( .A(b[5]), .B(a[103]), .Z(n14493) );
  NANDN U15335 ( .A(n14493), .B(n36587), .Z(n14326) );
  NANDN U15336 ( .A(n14324), .B(n36588), .Z(n14325) );
  AND U15337 ( .A(n14326), .B(n14325), .Z(n14530) );
  XNOR U15338 ( .A(n14529), .B(n14530), .Z(n14531) );
  XNOR U15339 ( .A(n14532), .B(n14531), .Z(n14517) );
  NAND U15340 ( .A(n14327), .B(n37762), .Z(n14329) );
  XOR U15341 ( .A(b[17]), .B(a[91]), .Z(n14496) );
  NAND U15342 ( .A(n14496), .B(n37764), .Z(n14328) );
  NAND U15343 ( .A(n14329), .B(n14328), .Z(n14471) );
  XNOR U15344 ( .A(b[31]), .B(a[77]), .Z(n14499) );
  NANDN U15345 ( .A(n14499), .B(n38552), .Z(n14332) );
  NANDN U15346 ( .A(n14330), .B(n38553), .Z(n14331) );
  AND U15347 ( .A(n14332), .B(n14331), .Z(n14469) );
  OR U15348 ( .A(n14333), .B(n36105), .Z(n14335) );
  XNOR U15349 ( .A(b[3]), .B(a[105]), .Z(n14502) );
  NANDN U15350 ( .A(n14502), .B(n36107), .Z(n14334) );
  AND U15351 ( .A(n14335), .B(n14334), .Z(n14470) );
  XOR U15352 ( .A(n14471), .B(n14472), .Z(n14518) );
  XOR U15353 ( .A(n14517), .B(n14518), .Z(n14519) );
  XNOR U15354 ( .A(n14520), .B(n14519), .Z(n14445) );
  NANDN U15355 ( .A(n14337), .B(n14336), .Z(n14341) );
  OR U15356 ( .A(n14339), .B(n14338), .Z(n14340) );
  NAND U15357 ( .A(n14341), .B(n14340), .Z(n14446) );
  XNOR U15358 ( .A(n14445), .B(n14446), .Z(n14447) );
  NANDN U15359 ( .A(n14343), .B(n14342), .Z(n14347) );
  NAND U15360 ( .A(n14345), .B(n14344), .Z(n14346) );
  NAND U15361 ( .A(n14347), .B(n14346), .Z(n14508) );
  NANDN U15362 ( .A(n14349), .B(n14348), .Z(n14353) );
  NAND U15363 ( .A(n14351), .B(n14350), .Z(n14352) );
  NAND U15364 ( .A(n14353), .B(n14352), .Z(n14505) );
  OR U15365 ( .A(n14355), .B(n14354), .Z(n14359) );
  NANDN U15366 ( .A(n14357), .B(n14356), .Z(n14358) );
  NAND U15367 ( .A(n14359), .B(n14358), .Z(n14506) );
  XNOR U15368 ( .A(n14505), .B(n14506), .Z(n14507) );
  XOR U15369 ( .A(n14508), .B(n14507), .Z(n14448) );
  XNOR U15370 ( .A(n14447), .B(n14448), .Z(n14573) );
  NANDN U15371 ( .A(n14365), .B(n14364), .Z(n14369) );
  NANDN U15372 ( .A(n14367), .B(n14366), .Z(n14368) );
  NAND U15373 ( .A(n14369), .B(n14368), .Z(n14454) );
  NANDN U15374 ( .A(n14375), .B(n14374), .Z(n14379) );
  NAND U15375 ( .A(n14377), .B(n14376), .Z(n14378) );
  NAND U15376 ( .A(n14379), .B(n14378), .Z(n14511) );
  NANDN U15377 ( .A(n14381), .B(n14380), .Z(n14385) );
  NAND U15378 ( .A(n14383), .B(n14382), .Z(n14384) );
  AND U15379 ( .A(n14385), .B(n14384), .Z(n14512) );
  XNOR U15380 ( .A(n14511), .B(n14512), .Z(n14513) );
  XOR U15381 ( .A(b[9]), .B(n17884), .Z(n14535) );
  NANDN U15382 ( .A(n14535), .B(n36925), .Z(n14388) );
  NANDN U15383 ( .A(n14386), .B(n36926), .Z(n14387) );
  NAND U15384 ( .A(n14388), .B(n14387), .Z(n14477) );
  XOR U15385 ( .A(b[15]), .B(n17031), .Z(n14538) );
  OR U15386 ( .A(n14538), .B(n37665), .Z(n14391) );
  NANDN U15387 ( .A(n14389), .B(n37604), .Z(n14390) );
  AND U15388 ( .A(n14391), .B(n14390), .Z(n14475) );
  XNOR U15389 ( .A(b[21]), .B(a[87]), .Z(n14541) );
  NANDN U15390 ( .A(n14541), .B(n38101), .Z(n14394) );
  NANDN U15391 ( .A(n14392), .B(n38102), .Z(n14393) );
  AND U15392 ( .A(n14394), .B(n14393), .Z(n14476) );
  XOR U15393 ( .A(n14477), .B(n14478), .Z(n14466) );
  XNOR U15394 ( .A(b[11]), .B(a[97]), .Z(n14544) );
  OR U15395 ( .A(n14544), .B(n37311), .Z(n14397) );
  NANDN U15396 ( .A(n14395), .B(n37218), .Z(n14396) );
  NAND U15397 ( .A(n14397), .B(n14396), .Z(n14464) );
  XOR U15398 ( .A(n1053), .B(a[95]), .Z(n14547) );
  NANDN U15399 ( .A(n14547), .B(n37424), .Z(n14400) );
  NANDN U15400 ( .A(n14398), .B(n37425), .Z(n14399) );
  NAND U15401 ( .A(n14400), .B(n14399), .Z(n14463) );
  XOR U15402 ( .A(n14466), .B(n14465), .Z(n14460) );
  NANDN U15403 ( .A(n1049), .B(a[107]), .Z(n14401) );
  XNOR U15404 ( .A(b[1]), .B(n14401), .Z(n14403) );
  NANDN U15405 ( .A(b[0]), .B(a[106]), .Z(n14402) );
  AND U15406 ( .A(n14403), .B(n14402), .Z(n14483) );
  NAND U15407 ( .A(n38490), .B(n14404), .Z(n14406) );
  XNOR U15408 ( .A(n1058), .B(a[79]), .Z(n14553) );
  NANDN U15409 ( .A(n1048), .B(n14553), .Z(n14405) );
  NAND U15410 ( .A(n14406), .B(n14405), .Z(n14481) );
  NANDN U15411 ( .A(n1059), .B(a[75]), .Z(n14482) );
  XNOR U15412 ( .A(n14481), .B(n14482), .Z(n14484) );
  XNOR U15413 ( .A(n14483), .B(n14484), .Z(n14458) );
  NANDN U15414 ( .A(n14407), .B(n38205), .Z(n14409) );
  XNOR U15415 ( .A(b[23]), .B(a[85]), .Z(n14556) );
  OR U15416 ( .A(n14556), .B(n38268), .Z(n14408) );
  NAND U15417 ( .A(n14409), .B(n14408), .Z(n14526) );
  XNOR U15418 ( .A(b[7]), .B(a[101]), .Z(n14559) );
  NANDN U15419 ( .A(n14559), .B(n36701), .Z(n14412) );
  NAND U15420 ( .A(n14410), .B(n36702), .Z(n14411) );
  NAND U15421 ( .A(n14412), .B(n14411), .Z(n14523) );
  XNOR U15422 ( .A(b[25]), .B(a[83]), .Z(n14562) );
  NANDN U15423 ( .A(n14562), .B(n38325), .Z(n14415) );
  NANDN U15424 ( .A(n14413), .B(n38326), .Z(n14414) );
  AND U15425 ( .A(n14415), .B(n14414), .Z(n14524) );
  XNOR U15426 ( .A(n14523), .B(n14524), .Z(n14525) );
  XOR U15427 ( .A(n14526), .B(n14525), .Z(n14457) );
  XOR U15428 ( .A(n14460), .B(n14459), .Z(n14514) );
  XNOR U15429 ( .A(n14513), .B(n14514), .Z(n14451) );
  XOR U15430 ( .A(n14452), .B(n14451), .Z(n14453) );
  XNOR U15431 ( .A(n14454), .B(n14453), .Z(n14571) );
  XNOR U15432 ( .A(n14572), .B(n14571), .Z(n14574) );
  XNOR U15433 ( .A(n14573), .B(n14574), .Z(n14568) );
  XOR U15434 ( .A(n14567), .B(n14568), .Z(n14442) );
  NANDN U15435 ( .A(n14417), .B(n14416), .Z(n14421) );
  NAND U15436 ( .A(n14419), .B(n14418), .Z(n14420) );
  NAND U15437 ( .A(n14421), .B(n14420), .Z(n14439) );
  NANDN U15438 ( .A(n14423), .B(n14422), .Z(n14427) );
  OR U15439 ( .A(n14425), .B(n14424), .Z(n14426) );
  NAND U15440 ( .A(n14427), .B(n14426), .Z(n14440) );
  XNOR U15441 ( .A(n14439), .B(n14440), .Z(n14441) );
  XNOR U15442 ( .A(n14442), .B(n14441), .Z(n14434) );
  XNOR U15443 ( .A(n14433), .B(n14434), .Z(n14435) );
  XNOR U15444 ( .A(n14436), .B(n14435), .Z(n14577) );
  XNOR U15445 ( .A(n14577), .B(sreg[331]), .Z(n14579) );
  NAND U15446 ( .A(n14428), .B(sreg[330]), .Z(n14432) );
  OR U15447 ( .A(n14430), .B(n14429), .Z(n14431) );
  AND U15448 ( .A(n14432), .B(n14431), .Z(n14578) );
  XOR U15449 ( .A(n14579), .B(n14578), .Z(c[331]) );
  NANDN U15450 ( .A(n14434), .B(n14433), .Z(n14438) );
  NAND U15451 ( .A(n14436), .B(n14435), .Z(n14437) );
  NAND U15452 ( .A(n14438), .B(n14437), .Z(n14585) );
  NANDN U15453 ( .A(n14440), .B(n14439), .Z(n14444) );
  NAND U15454 ( .A(n14442), .B(n14441), .Z(n14443) );
  NAND U15455 ( .A(n14444), .B(n14443), .Z(n14583) );
  NANDN U15456 ( .A(n14446), .B(n14445), .Z(n14450) );
  NANDN U15457 ( .A(n14448), .B(n14447), .Z(n14449) );
  NAND U15458 ( .A(n14450), .B(n14449), .Z(n14718) );
  NAND U15459 ( .A(n14452), .B(n14451), .Z(n14456) );
  NAND U15460 ( .A(n14454), .B(n14453), .Z(n14455) );
  NAND U15461 ( .A(n14456), .B(n14455), .Z(n14719) );
  XNOR U15462 ( .A(n14718), .B(n14719), .Z(n14720) );
  NANDN U15463 ( .A(n14458), .B(n14457), .Z(n14462) );
  NANDN U15464 ( .A(n14460), .B(n14459), .Z(n14461) );
  NAND U15465 ( .A(n14462), .B(n14461), .Z(n14705) );
  OR U15466 ( .A(n14464), .B(n14463), .Z(n14468) );
  NAND U15467 ( .A(n14466), .B(n14465), .Z(n14467) );
  NAND U15468 ( .A(n14468), .B(n14467), .Z(n14644) );
  OR U15469 ( .A(n14470), .B(n14469), .Z(n14474) );
  NANDN U15470 ( .A(n14472), .B(n14471), .Z(n14473) );
  NAND U15471 ( .A(n14474), .B(n14473), .Z(n14643) );
  OR U15472 ( .A(n14476), .B(n14475), .Z(n14480) );
  NANDN U15473 ( .A(n14478), .B(n14477), .Z(n14479) );
  NAND U15474 ( .A(n14480), .B(n14479), .Z(n14642) );
  XOR U15475 ( .A(n14644), .B(n14645), .Z(n14702) );
  NANDN U15476 ( .A(n14482), .B(n14481), .Z(n14486) );
  NAND U15477 ( .A(n14484), .B(n14483), .Z(n14485) );
  NAND U15478 ( .A(n14486), .B(n14485), .Z(n14657) );
  XNOR U15479 ( .A(b[19]), .B(a[90]), .Z(n14600) );
  NANDN U15480 ( .A(n14600), .B(n37934), .Z(n14489) );
  NANDN U15481 ( .A(n14487), .B(n37935), .Z(n14488) );
  NAND U15482 ( .A(n14489), .B(n14488), .Z(n14669) );
  XNOR U15483 ( .A(b[27]), .B(a[82]), .Z(n14603) );
  NANDN U15484 ( .A(n14603), .B(n38423), .Z(n14492) );
  NAND U15485 ( .A(n14490), .B(n38424), .Z(n14491) );
  NAND U15486 ( .A(n14492), .B(n14491), .Z(n14666) );
  XNOR U15487 ( .A(b[5]), .B(a[104]), .Z(n14606) );
  NANDN U15488 ( .A(n14606), .B(n36587), .Z(n14495) );
  NANDN U15489 ( .A(n14493), .B(n36588), .Z(n14494) );
  AND U15490 ( .A(n14495), .B(n14494), .Z(n14667) );
  XNOR U15491 ( .A(n14666), .B(n14667), .Z(n14668) );
  XNOR U15492 ( .A(n14669), .B(n14668), .Z(n14655) );
  NAND U15493 ( .A(n14496), .B(n37762), .Z(n14498) );
  XOR U15494 ( .A(b[17]), .B(a[92]), .Z(n14609) );
  NAND U15495 ( .A(n14609), .B(n37764), .Z(n14497) );
  NAND U15496 ( .A(n14498), .B(n14497), .Z(n14627) );
  XNOR U15497 ( .A(b[31]), .B(a[78]), .Z(n14612) );
  NANDN U15498 ( .A(n14612), .B(n38552), .Z(n14501) );
  NANDN U15499 ( .A(n14499), .B(n38553), .Z(n14500) );
  NAND U15500 ( .A(n14501), .B(n14500), .Z(n14624) );
  OR U15501 ( .A(n14502), .B(n36105), .Z(n14504) );
  XNOR U15502 ( .A(b[3]), .B(a[106]), .Z(n14615) );
  NANDN U15503 ( .A(n14615), .B(n36107), .Z(n14503) );
  AND U15504 ( .A(n14504), .B(n14503), .Z(n14625) );
  XNOR U15505 ( .A(n14624), .B(n14625), .Z(n14626) );
  XOR U15506 ( .A(n14627), .B(n14626), .Z(n14654) );
  XNOR U15507 ( .A(n14655), .B(n14654), .Z(n14656) );
  XNOR U15508 ( .A(n14657), .B(n14656), .Z(n14703) );
  XNOR U15509 ( .A(n14702), .B(n14703), .Z(n14704) );
  XNOR U15510 ( .A(n14705), .B(n14704), .Z(n14715) );
  NANDN U15511 ( .A(n14506), .B(n14505), .Z(n14510) );
  NANDN U15512 ( .A(n14508), .B(n14507), .Z(n14509) );
  NAND U15513 ( .A(n14510), .B(n14509), .Z(n14712) );
  NANDN U15514 ( .A(n14512), .B(n14511), .Z(n14516) );
  NANDN U15515 ( .A(n14514), .B(n14513), .Z(n14515) );
  NAND U15516 ( .A(n14516), .B(n14515), .Z(n14709) );
  OR U15517 ( .A(n14518), .B(n14517), .Z(n14522) );
  NAND U15518 ( .A(n14520), .B(n14519), .Z(n14521) );
  NAND U15519 ( .A(n14522), .B(n14521), .Z(n14706) );
  NANDN U15520 ( .A(n14524), .B(n14523), .Z(n14528) );
  NAND U15521 ( .A(n14526), .B(n14525), .Z(n14527) );
  NAND U15522 ( .A(n14528), .B(n14527), .Z(n14648) );
  NANDN U15523 ( .A(n14530), .B(n14529), .Z(n14534) );
  NAND U15524 ( .A(n14532), .B(n14531), .Z(n14533) );
  AND U15525 ( .A(n14534), .B(n14533), .Z(n14649) );
  XNOR U15526 ( .A(n14648), .B(n14649), .Z(n14650) );
  XNOR U15527 ( .A(n1052), .B(a[100]), .Z(n14672) );
  NAND U15528 ( .A(n36925), .B(n14672), .Z(n14537) );
  NANDN U15529 ( .A(n14535), .B(n36926), .Z(n14536) );
  NAND U15530 ( .A(n14537), .B(n14536), .Z(n14632) );
  XNOR U15531 ( .A(b[15]), .B(a[94]), .Z(n14675) );
  OR U15532 ( .A(n14675), .B(n37665), .Z(n14540) );
  NANDN U15533 ( .A(n14538), .B(n37604), .Z(n14539) );
  AND U15534 ( .A(n14540), .B(n14539), .Z(n14630) );
  XNOR U15535 ( .A(n1056), .B(a[88]), .Z(n14678) );
  NAND U15536 ( .A(n14678), .B(n38101), .Z(n14543) );
  NANDN U15537 ( .A(n14541), .B(n38102), .Z(n14542) );
  AND U15538 ( .A(n14543), .B(n14542), .Z(n14631) );
  XOR U15539 ( .A(n14632), .B(n14633), .Z(n14621) );
  XNOR U15540 ( .A(b[11]), .B(a[98]), .Z(n14681) );
  OR U15541 ( .A(n14681), .B(n37311), .Z(n14546) );
  NANDN U15542 ( .A(n14544), .B(n37218), .Z(n14545) );
  NAND U15543 ( .A(n14546), .B(n14545), .Z(n14619) );
  XOR U15544 ( .A(n1053), .B(a[96]), .Z(n14684) );
  NANDN U15545 ( .A(n14684), .B(n37424), .Z(n14549) );
  NANDN U15546 ( .A(n14547), .B(n37425), .Z(n14548) );
  AND U15547 ( .A(n14549), .B(n14548), .Z(n14618) );
  XNOR U15548 ( .A(n14619), .B(n14618), .Z(n14620) );
  XOR U15549 ( .A(n14621), .B(n14620), .Z(n14638) );
  NANDN U15550 ( .A(n1049), .B(a[108]), .Z(n14550) );
  XNOR U15551 ( .A(b[1]), .B(n14550), .Z(n14552) );
  IV U15552 ( .A(a[107]), .Z(n18980) );
  NANDN U15553 ( .A(n18980), .B(n1049), .Z(n14551) );
  AND U15554 ( .A(n14552), .B(n14551), .Z(n14596) );
  NAND U15555 ( .A(n38490), .B(n14553), .Z(n14555) );
  XOR U15556 ( .A(n1058), .B(n15068), .Z(n14687) );
  NANDN U15557 ( .A(n1048), .B(n14687), .Z(n14554) );
  NAND U15558 ( .A(n14555), .B(n14554), .Z(n14594) );
  NANDN U15559 ( .A(n1059), .B(a[76]), .Z(n14595) );
  XNOR U15560 ( .A(n14594), .B(n14595), .Z(n14597) );
  XOR U15561 ( .A(n14596), .B(n14597), .Z(n14636) );
  NANDN U15562 ( .A(n14556), .B(n38205), .Z(n14558) );
  XNOR U15563 ( .A(b[23]), .B(a[86]), .Z(n14693) );
  OR U15564 ( .A(n14693), .B(n38268), .Z(n14557) );
  NAND U15565 ( .A(n14558), .B(n14557), .Z(n14663) );
  XOR U15566 ( .A(b[7]), .B(a[102]), .Z(n14696) );
  NAND U15567 ( .A(n14696), .B(n36701), .Z(n14561) );
  NANDN U15568 ( .A(n14559), .B(n36702), .Z(n14560) );
  NAND U15569 ( .A(n14561), .B(n14560), .Z(n14660) );
  XOR U15570 ( .A(b[25]), .B(a[84]), .Z(n14699) );
  NAND U15571 ( .A(n14699), .B(n38325), .Z(n14564) );
  NANDN U15572 ( .A(n14562), .B(n38326), .Z(n14563) );
  AND U15573 ( .A(n14564), .B(n14563), .Z(n14661) );
  XNOR U15574 ( .A(n14660), .B(n14661), .Z(n14662) );
  XNOR U15575 ( .A(n14663), .B(n14662), .Z(n14637) );
  XOR U15576 ( .A(n14636), .B(n14637), .Z(n14639) );
  XNOR U15577 ( .A(n14638), .B(n14639), .Z(n14651) );
  XOR U15578 ( .A(n14650), .B(n14651), .Z(n14707) );
  XNOR U15579 ( .A(n14706), .B(n14707), .Z(n14708) );
  XOR U15580 ( .A(n14709), .B(n14708), .Z(n14713) );
  XNOR U15581 ( .A(n14712), .B(n14713), .Z(n14714) );
  XOR U15582 ( .A(n14715), .B(n14714), .Z(n14721) );
  XOR U15583 ( .A(n14720), .B(n14721), .Z(n14590) );
  NANDN U15584 ( .A(n14566), .B(n14565), .Z(n14570) );
  NANDN U15585 ( .A(n14568), .B(n14567), .Z(n14569) );
  NAND U15586 ( .A(n14570), .B(n14569), .Z(n14589) );
  OR U15587 ( .A(n14572), .B(n14571), .Z(n14576) );
  OR U15588 ( .A(n14574), .B(n14573), .Z(n14575) );
  AND U15589 ( .A(n14576), .B(n14575), .Z(n14588) );
  XNOR U15590 ( .A(n14589), .B(n14588), .Z(n14591) );
  XOR U15591 ( .A(n14590), .B(n14591), .Z(n14582) );
  XOR U15592 ( .A(n14583), .B(n14582), .Z(n14584) );
  XNOR U15593 ( .A(n14585), .B(n14584), .Z(n14724) );
  XNOR U15594 ( .A(n14724), .B(sreg[332]), .Z(n14726) );
  NAND U15595 ( .A(n14577), .B(sreg[331]), .Z(n14581) );
  OR U15596 ( .A(n14579), .B(n14578), .Z(n14580) );
  AND U15597 ( .A(n14581), .B(n14580), .Z(n14725) );
  XOR U15598 ( .A(n14726), .B(n14725), .Z(c[332]) );
  NAND U15599 ( .A(n14583), .B(n14582), .Z(n14587) );
  NAND U15600 ( .A(n14585), .B(n14584), .Z(n14586) );
  NAND U15601 ( .A(n14587), .B(n14586), .Z(n14732) );
  NANDN U15602 ( .A(n14589), .B(n14588), .Z(n14593) );
  NAND U15603 ( .A(n14591), .B(n14590), .Z(n14592) );
  NAND U15604 ( .A(n14593), .B(n14592), .Z(n14730) );
  NANDN U15605 ( .A(n14595), .B(n14594), .Z(n14599) );
  NAND U15606 ( .A(n14597), .B(n14596), .Z(n14598) );
  NAND U15607 ( .A(n14599), .B(n14598), .Z(n14814) );
  XNOR U15608 ( .A(b[19]), .B(a[91]), .Z(n14759) );
  NANDN U15609 ( .A(n14759), .B(n37934), .Z(n14602) );
  NANDN U15610 ( .A(n14600), .B(n37935), .Z(n14601) );
  NAND U15611 ( .A(n14602), .B(n14601), .Z(n14824) );
  XNOR U15612 ( .A(b[27]), .B(a[83]), .Z(n14762) );
  NANDN U15613 ( .A(n14762), .B(n38423), .Z(n14605) );
  NANDN U15614 ( .A(n14603), .B(n38424), .Z(n14604) );
  NAND U15615 ( .A(n14605), .B(n14604), .Z(n14821) );
  XNOR U15616 ( .A(b[5]), .B(a[105]), .Z(n14765) );
  NANDN U15617 ( .A(n14765), .B(n36587), .Z(n14608) );
  NANDN U15618 ( .A(n14606), .B(n36588), .Z(n14607) );
  AND U15619 ( .A(n14608), .B(n14607), .Z(n14822) );
  XNOR U15620 ( .A(n14821), .B(n14822), .Z(n14823) );
  XNOR U15621 ( .A(n14824), .B(n14823), .Z(n14812) );
  NAND U15622 ( .A(n14609), .B(n37762), .Z(n14611) );
  XNOR U15623 ( .A(b[17]), .B(a[93]), .Z(n14768) );
  NANDN U15624 ( .A(n14768), .B(n37764), .Z(n14610) );
  NAND U15625 ( .A(n14611), .B(n14610), .Z(n14786) );
  XNOR U15626 ( .A(b[31]), .B(a[79]), .Z(n14771) );
  NANDN U15627 ( .A(n14771), .B(n38552), .Z(n14614) );
  NANDN U15628 ( .A(n14612), .B(n38553), .Z(n14613) );
  NAND U15629 ( .A(n14614), .B(n14613), .Z(n14783) );
  OR U15630 ( .A(n14615), .B(n36105), .Z(n14617) );
  XOR U15631 ( .A(b[3]), .B(n18980), .Z(n14774) );
  NANDN U15632 ( .A(n14774), .B(n36107), .Z(n14616) );
  AND U15633 ( .A(n14617), .B(n14616), .Z(n14784) );
  XNOR U15634 ( .A(n14783), .B(n14784), .Z(n14785) );
  XOR U15635 ( .A(n14786), .B(n14785), .Z(n14811) );
  XNOR U15636 ( .A(n14812), .B(n14811), .Z(n14813) );
  XNOR U15637 ( .A(n14814), .B(n14813), .Z(n14857) );
  NANDN U15638 ( .A(n14619), .B(n14618), .Z(n14623) );
  NAND U15639 ( .A(n14621), .B(n14620), .Z(n14622) );
  NAND U15640 ( .A(n14623), .B(n14622), .Z(n14802) );
  NANDN U15641 ( .A(n14625), .B(n14624), .Z(n14629) );
  NAND U15642 ( .A(n14627), .B(n14626), .Z(n14628) );
  NAND U15643 ( .A(n14629), .B(n14628), .Z(n14800) );
  OR U15644 ( .A(n14631), .B(n14630), .Z(n14635) );
  NANDN U15645 ( .A(n14633), .B(n14632), .Z(n14634) );
  NAND U15646 ( .A(n14635), .B(n14634), .Z(n14799) );
  XNOR U15647 ( .A(n14802), .B(n14801), .Z(n14858) );
  XOR U15648 ( .A(n14857), .B(n14858), .Z(n14860) );
  NANDN U15649 ( .A(n14637), .B(n14636), .Z(n14641) );
  OR U15650 ( .A(n14639), .B(n14638), .Z(n14640) );
  NAND U15651 ( .A(n14641), .B(n14640), .Z(n14859) );
  XOR U15652 ( .A(n14860), .B(n14859), .Z(n14749) );
  OR U15653 ( .A(n14643), .B(n14642), .Z(n14647) );
  NANDN U15654 ( .A(n14645), .B(n14644), .Z(n14646) );
  NAND U15655 ( .A(n14647), .B(n14646), .Z(n14748) );
  NANDN U15656 ( .A(n14649), .B(n14648), .Z(n14653) );
  NANDN U15657 ( .A(n14651), .B(n14650), .Z(n14652) );
  NAND U15658 ( .A(n14653), .B(n14652), .Z(n14865) );
  NANDN U15659 ( .A(n14655), .B(n14654), .Z(n14659) );
  NAND U15660 ( .A(n14657), .B(n14656), .Z(n14658) );
  NAND U15661 ( .A(n14659), .B(n14658), .Z(n14864) );
  NANDN U15662 ( .A(n14661), .B(n14660), .Z(n14665) );
  NAND U15663 ( .A(n14663), .B(n14662), .Z(n14664) );
  NAND U15664 ( .A(n14665), .B(n14664), .Z(n14805) );
  NANDN U15665 ( .A(n14667), .B(n14666), .Z(n14671) );
  NAND U15666 ( .A(n14669), .B(n14668), .Z(n14670) );
  AND U15667 ( .A(n14671), .B(n14670), .Z(n14806) );
  XNOR U15668 ( .A(n14805), .B(n14806), .Z(n14807) );
  XOR U15669 ( .A(n1052), .B(a[101]), .Z(n14833) );
  NANDN U15670 ( .A(n14833), .B(n36925), .Z(n14674) );
  NAND U15671 ( .A(n36926), .B(n14672), .Z(n14673) );
  NAND U15672 ( .A(n14674), .B(n14673), .Z(n14791) );
  XNOR U15673 ( .A(n1054), .B(a[95]), .Z(n14830) );
  NANDN U15674 ( .A(n37665), .B(n14830), .Z(n14677) );
  NANDN U15675 ( .A(n14675), .B(n37604), .Z(n14676) );
  NAND U15676 ( .A(n14677), .B(n14676), .Z(n14789) );
  XOR U15677 ( .A(n1056), .B(a[89]), .Z(n14827) );
  NANDN U15678 ( .A(n14827), .B(n38101), .Z(n14680) );
  NAND U15679 ( .A(n38102), .B(n14678), .Z(n14679) );
  NAND U15680 ( .A(n14680), .B(n14679), .Z(n14790) );
  XNOR U15681 ( .A(n14789), .B(n14790), .Z(n14792) );
  XOR U15682 ( .A(n14791), .B(n14792), .Z(n14780) );
  XOR U15683 ( .A(b[11]), .B(n17884), .Z(n14836) );
  OR U15684 ( .A(n14836), .B(n37311), .Z(n14683) );
  NANDN U15685 ( .A(n14681), .B(n37218), .Z(n14682) );
  NAND U15686 ( .A(n14683), .B(n14682), .Z(n14778) );
  XOR U15687 ( .A(n1053), .B(a[97]), .Z(n14839) );
  NANDN U15688 ( .A(n14839), .B(n37424), .Z(n14686) );
  NANDN U15689 ( .A(n14684), .B(n37425), .Z(n14685) );
  AND U15690 ( .A(n14686), .B(n14685), .Z(n14777) );
  XNOR U15691 ( .A(n14778), .B(n14777), .Z(n14779) );
  XNOR U15692 ( .A(n14780), .B(n14779), .Z(n14796) );
  NAND U15693 ( .A(n38490), .B(n14687), .Z(n14689) );
  XNOR U15694 ( .A(n1058), .B(a[81]), .Z(n14845) );
  NANDN U15695 ( .A(n1048), .B(n14845), .Z(n14688) );
  NAND U15696 ( .A(n14689), .B(n14688), .Z(n14753) );
  NANDN U15697 ( .A(n1059), .B(a[77]), .Z(n14754) );
  XNOR U15698 ( .A(n14753), .B(n14754), .Z(n14756) );
  NANDN U15699 ( .A(n1049), .B(a[109]), .Z(n14690) );
  XNOR U15700 ( .A(b[1]), .B(n14690), .Z(n14692) );
  NANDN U15701 ( .A(b[0]), .B(a[108]), .Z(n14691) );
  AND U15702 ( .A(n14692), .B(n14691), .Z(n14755) );
  XNOR U15703 ( .A(n14756), .B(n14755), .Z(n14794) );
  NANDN U15704 ( .A(n14693), .B(n38205), .Z(n14695) );
  XNOR U15705 ( .A(b[23]), .B(a[87]), .Z(n14848) );
  OR U15706 ( .A(n14848), .B(n38268), .Z(n14694) );
  NAND U15707 ( .A(n14695), .B(n14694), .Z(n14818) );
  XOR U15708 ( .A(b[7]), .B(a[103]), .Z(n14851) );
  NAND U15709 ( .A(n14851), .B(n36701), .Z(n14698) );
  NAND U15710 ( .A(n14696), .B(n36702), .Z(n14697) );
  NAND U15711 ( .A(n14698), .B(n14697), .Z(n14815) );
  XOR U15712 ( .A(b[25]), .B(a[85]), .Z(n14854) );
  NAND U15713 ( .A(n14854), .B(n38325), .Z(n14701) );
  NAND U15714 ( .A(n14699), .B(n38326), .Z(n14700) );
  AND U15715 ( .A(n14701), .B(n14700), .Z(n14816) );
  XNOR U15716 ( .A(n14815), .B(n14816), .Z(n14817) );
  XOR U15717 ( .A(n14818), .B(n14817), .Z(n14793) );
  XOR U15718 ( .A(n14796), .B(n14795), .Z(n14808) );
  XOR U15719 ( .A(n14807), .B(n14808), .Z(n14863) );
  XNOR U15720 ( .A(n14864), .B(n14863), .Z(n14866) );
  XNOR U15721 ( .A(n14865), .B(n14866), .Z(n14747) );
  XOR U15722 ( .A(n14748), .B(n14747), .Z(n14750) );
  NANDN U15723 ( .A(n14707), .B(n14706), .Z(n14711) );
  NAND U15724 ( .A(n14709), .B(n14708), .Z(n14710) );
  AND U15725 ( .A(n14711), .B(n14710), .Z(n14741) );
  XNOR U15726 ( .A(n14742), .B(n14741), .Z(n14743) );
  XOR U15727 ( .A(n14744), .B(n14743), .Z(n14737) );
  NANDN U15728 ( .A(n14713), .B(n14712), .Z(n14717) );
  NAND U15729 ( .A(n14715), .B(n14714), .Z(n14716) );
  NAND U15730 ( .A(n14717), .B(n14716), .Z(n14735) );
  NANDN U15731 ( .A(n14719), .B(n14718), .Z(n14723) );
  NAND U15732 ( .A(n14721), .B(n14720), .Z(n14722) );
  AND U15733 ( .A(n14723), .B(n14722), .Z(n14736) );
  XNOR U15734 ( .A(n14735), .B(n14736), .Z(n14738) );
  XOR U15735 ( .A(n14737), .B(n14738), .Z(n14729) );
  XOR U15736 ( .A(n14730), .B(n14729), .Z(n14731) );
  XNOR U15737 ( .A(n14732), .B(n14731), .Z(n14869) );
  XNOR U15738 ( .A(n14869), .B(sreg[333]), .Z(n14871) );
  NAND U15739 ( .A(n14724), .B(sreg[332]), .Z(n14728) );
  OR U15740 ( .A(n14726), .B(n14725), .Z(n14727) );
  AND U15741 ( .A(n14728), .B(n14727), .Z(n14870) );
  XOR U15742 ( .A(n14871), .B(n14870), .Z(c[333]) );
  NAND U15743 ( .A(n14730), .B(n14729), .Z(n14734) );
  NAND U15744 ( .A(n14732), .B(n14731), .Z(n14733) );
  NAND U15745 ( .A(n14734), .B(n14733), .Z(n14877) );
  NANDN U15746 ( .A(n14736), .B(n14735), .Z(n14740) );
  NAND U15747 ( .A(n14738), .B(n14737), .Z(n14739) );
  NAND U15748 ( .A(n14740), .B(n14739), .Z(n14875) );
  NANDN U15749 ( .A(n14742), .B(n14741), .Z(n14746) );
  NAND U15750 ( .A(n14744), .B(n14743), .Z(n14745) );
  NAND U15751 ( .A(n14746), .B(n14745), .Z(n14880) );
  NANDN U15752 ( .A(n14748), .B(n14747), .Z(n14752) );
  OR U15753 ( .A(n14750), .B(n14749), .Z(n14751) );
  NAND U15754 ( .A(n14752), .B(n14751), .Z(n14881) );
  XNOR U15755 ( .A(n14880), .B(n14881), .Z(n14882) );
  NANDN U15756 ( .A(n14754), .B(n14753), .Z(n14758) );
  NAND U15757 ( .A(n14756), .B(n14755), .Z(n14757) );
  NAND U15758 ( .A(n14758), .B(n14757), .Z(n14955) );
  XNOR U15759 ( .A(b[19]), .B(a[92]), .Z(n14902) );
  NANDN U15760 ( .A(n14902), .B(n37934), .Z(n14761) );
  NANDN U15761 ( .A(n14759), .B(n37935), .Z(n14760) );
  NAND U15762 ( .A(n14761), .B(n14760), .Z(n14965) );
  XOR U15763 ( .A(b[27]), .B(a[84]), .Z(n14905) );
  NAND U15764 ( .A(n38423), .B(n14905), .Z(n14764) );
  NANDN U15765 ( .A(n14762), .B(n38424), .Z(n14763) );
  NAND U15766 ( .A(n14764), .B(n14763), .Z(n14962) );
  XNOR U15767 ( .A(b[5]), .B(a[106]), .Z(n14908) );
  NANDN U15768 ( .A(n14908), .B(n36587), .Z(n14767) );
  NANDN U15769 ( .A(n14765), .B(n36588), .Z(n14766) );
  AND U15770 ( .A(n14767), .B(n14766), .Z(n14963) );
  XNOR U15771 ( .A(n14962), .B(n14963), .Z(n14964) );
  XNOR U15772 ( .A(n14965), .B(n14964), .Z(n14953) );
  NANDN U15773 ( .A(n14768), .B(n37762), .Z(n14770) );
  XOR U15774 ( .A(b[17]), .B(a[94]), .Z(n14911) );
  NAND U15775 ( .A(n14911), .B(n37764), .Z(n14769) );
  NAND U15776 ( .A(n14770), .B(n14769), .Z(n14929) );
  XOR U15777 ( .A(b[31]), .B(n15068), .Z(n14914) );
  NANDN U15778 ( .A(n14914), .B(n38552), .Z(n14773) );
  NANDN U15779 ( .A(n14771), .B(n38553), .Z(n14772) );
  NAND U15780 ( .A(n14773), .B(n14772), .Z(n14926) );
  OR U15781 ( .A(n14774), .B(n36105), .Z(n14776) );
  XNOR U15782 ( .A(b[3]), .B(a[108]), .Z(n14917) );
  NANDN U15783 ( .A(n14917), .B(n36107), .Z(n14775) );
  AND U15784 ( .A(n14776), .B(n14775), .Z(n14927) );
  XNOR U15785 ( .A(n14926), .B(n14927), .Z(n14928) );
  XOR U15786 ( .A(n14929), .B(n14928), .Z(n14952) );
  XNOR U15787 ( .A(n14953), .B(n14952), .Z(n14954) );
  XNOR U15788 ( .A(n14955), .B(n14954), .Z(n14893) );
  NANDN U15789 ( .A(n14778), .B(n14777), .Z(n14782) );
  NAND U15790 ( .A(n14780), .B(n14779), .Z(n14781) );
  NAND U15791 ( .A(n14782), .B(n14781), .Z(n14944) );
  NANDN U15792 ( .A(n14784), .B(n14783), .Z(n14788) );
  NAND U15793 ( .A(n14786), .B(n14785), .Z(n14787) );
  NAND U15794 ( .A(n14788), .B(n14787), .Z(n14943) );
  XNOR U15795 ( .A(n14943), .B(n14942), .Z(n14945) );
  XOR U15796 ( .A(n14944), .B(n14945), .Z(n14892) );
  XOR U15797 ( .A(n14893), .B(n14892), .Z(n14894) );
  NANDN U15798 ( .A(n14794), .B(n14793), .Z(n14798) );
  NAND U15799 ( .A(n14796), .B(n14795), .Z(n14797) );
  NAND U15800 ( .A(n14798), .B(n14797), .Z(n14895) );
  XNOR U15801 ( .A(n14894), .B(n14895), .Z(n15006) );
  OR U15802 ( .A(n14800), .B(n14799), .Z(n14804) );
  NAND U15803 ( .A(n14802), .B(n14801), .Z(n14803) );
  NAND U15804 ( .A(n14804), .B(n14803), .Z(n15005) );
  NANDN U15805 ( .A(n14806), .B(n14805), .Z(n14810) );
  NAND U15806 ( .A(n14808), .B(n14807), .Z(n14809) );
  NAND U15807 ( .A(n14810), .B(n14809), .Z(n14888) );
  NANDN U15808 ( .A(n14816), .B(n14815), .Z(n14820) );
  NAND U15809 ( .A(n14818), .B(n14817), .Z(n14819) );
  NAND U15810 ( .A(n14820), .B(n14819), .Z(n14946) );
  NANDN U15811 ( .A(n14822), .B(n14821), .Z(n14826) );
  NAND U15812 ( .A(n14824), .B(n14823), .Z(n14825) );
  AND U15813 ( .A(n14826), .B(n14825), .Z(n14947) );
  XNOR U15814 ( .A(n14946), .B(n14947), .Z(n14948) );
  XNOR U15815 ( .A(b[21]), .B(a[90]), .Z(n14974) );
  NANDN U15816 ( .A(n14974), .B(n38101), .Z(n14829) );
  NANDN U15817 ( .A(n14827), .B(n38102), .Z(n14828) );
  NAND U15818 ( .A(n14829), .B(n14828), .Z(n14938) );
  XNOR U15819 ( .A(b[15]), .B(a[96]), .Z(n14971) );
  OR U15820 ( .A(n14971), .B(n37665), .Z(n14832) );
  NAND U15821 ( .A(n14830), .B(n37604), .Z(n14831) );
  AND U15822 ( .A(n14832), .B(n14831), .Z(n14939) );
  XNOR U15823 ( .A(n14938), .B(n14939), .Z(n14941) );
  XNOR U15824 ( .A(b[9]), .B(a[102]), .Z(n14968) );
  NANDN U15825 ( .A(n14968), .B(n36925), .Z(n14835) );
  NANDN U15826 ( .A(n14833), .B(n36926), .Z(n14834) );
  NAND U15827 ( .A(n14835), .B(n14834), .Z(n14940) );
  XNOR U15828 ( .A(n14941), .B(n14940), .Z(n14934) );
  XNOR U15829 ( .A(b[11]), .B(a[100]), .Z(n14977) );
  OR U15830 ( .A(n14977), .B(n37311), .Z(n14838) );
  NANDN U15831 ( .A(n14836), .B(n37218), .Z(n14837) );
  NAND U15832 ( .A(n14838), .B(n14837), .Z(n14933) );
  XOR U15833 ( .A(n1053), .B(a[98]), .Z(n14980) );
  NANDN U15834 ( .A(n14980), .B(n37424), .Z(n14841) );
  NANDN U15835 ( .A(n14839), .B(n37425), .Z(n14840) );
  NAND U15836 ( .A(n14841), .B(n14840), .Z(n14932) );
  XNOR U15837 ( .A(n14933), .B(n14932), .Z(n14935) );
  XNOR U15838 ( .A(n14934), .B(n14935), .Z(n14923) );
  NANDN U15839 ( .A(n1049), .B(a[110]), .Z(n14842) );
  XNOR U15840 ( .A(b[1]), .B(n14842), .Z(n14844) );
  NANDN U15841 ( .A(b[0]), .B(a[109]), .Z(n14843) );
  AND U15842 ( .A(n14844), .B(n14843), .Z(n14898) );
  NAND U15843 ( .A(n38490), .B(n14845), .Z(n14847) );
  XOR U15844 ( .A(n1058), .B(n15424), .Z(n14986) );
  NANDN U15845 ( .A(n1048), .B(n14986), .Z(n14846) );
  NAND U15846 ( .A(n14847), .B(n14846), .Z(n14896) );
  NANDN U15847 ( .A(n1059), .B(a[78]), .Z(n14897) );
  XNOR U15848 ( .A(n14896), .B(n14897), .Z(n14899) );
  XNOR U15849 ( .A(n14898), .B(n14899), .Z(n14921) );
  NANDN U15850 ( .A(n14848), .B(n38205), .Z(n14850) );
  XNOR U15851 ( .A(b[23]), .B(a[88]), .Z(n14989) );
  OR U15852 ( .A(n14989), .B(n38268), .Z(n14849) );
  NAND U15853 ( .A(n14850), .B(n14849), .Z(n14959) );
  XOR U15854 ( .A(b[7]), .B(a[104]), .Z(n14992) );
  NAND U15855 ( .A(n14992), .B(n36701), .Z(n14853) );
  NAND U15856 ( .A(n14851), .B(n36702), .Z(n14852) );
  NAND U15857 ( .A(n14853), .B(n14852), .Z(n14956) );
  XOR U15858 ( .A(b[25]), .B(a[86]), .Z(n14995) );
  NAND U15859 ( .A(n14995), .B(n38325), .Z(n14856) );
  NAND U15860 ( .A(n14854), .B(n38326), .Z(n14855) );
  AND U15861 ( .A(n14856), .B(n14855), .Z(n14957) );
  XNOR U15862 ( .A(n14956), .B(n14957), .Z(n14958) );
  XOR U15863 ( .A(n14959), .B(n14958), .Z(n14920) );
  XOR U15864 ( .A(n14923), .B(n14922), .Z(n14949) );
  XNOR U15865 ( .A(n14948), .B(n14949), .Z(n14886) );
  XNOR U15866 ( .A(n14887), .B(n14886), .Z(n14889) );
  XNOR U15867 ( .A(n14888), .B(n14889), .Z(n15004) );
  XOR U15868 ( .A(n15005), .B(n15004), .Z(n15007) );
  NANDN U15869 ( .A(n14858), .B(n14857), .Z(n14862) );
  OR U15870 ( .A(n14860), .B(n14859), .Z(n14861) );
  NAND U15871 ( .A(n14862), .B(n14861), .Z(n14998) );
  NAND U15872 ( .A(n14864), .B(n14863), .Z(n14868) );
  NANDN U15873 ( .A(n14866), .B(n14865), .Z(n14867) );
  NAND U15874 ( .A(n14868), .B(n14867), .Z(n14999) );
  XNOR U15875 ( .A(n14998), .B(n14999), .Z(n15000) );
  XOR U15876 ( .A(n15001), .B(n15000), .Z(n14883) );
  XOR U15877 ( .A(n14882), .B(n14883), .Z(n14874) );
  XOR U15878 ( .A(n14875), .B(n14874), .Z(n14876) );
  XNOR U15879 ( .A(n14877), .B(n14876), .Z(n15010) );
  XNOR U15880 ( .A(n15010), .B(sreg[334]), .Z(n15012) );
  NAND U15881 ( .A(n14869), .B(sreg[333]), .Z(n14873) );
  OR U15882 ( .A(n14871), .B(n14870), .Z(n14872) );
  AND U15883 ( .A(n14873), .B(n14872), .Z(n15011) );
  XOR U15884 ( .A(n15012), .B(n15011), .Z(c[334]) );
  NAND U15885 ( .A(n14875), .B(n14874), .Z(n14879) );
  NAND U15886 ( .A(n14877), .B(n14876), .Z(n14878) );
  NAND U15887 ( .A(n14879), .B(n14878), .Z(n15018) );
  NANDN U15888 ( .A(n14881), .B(n14880), .Z(n14885) );
  NAND U15889 ( .A(n14883), .B(n14882), .Z(n14884) );
  NAND U15890 ( .A(n14885), .B(n14884), .Z(n15015) );
  NAND U15891 ( .A(n14887), .B(n14886), .Z(n14891) );
  NANDN U15892 ( .A(n14889), .B(n14888), .Z(n14890) );
  NAND U15893 ( .A(n14891), .B(n14890), .Z(n15144) );
  XNOR U15894 ( .A(n15144), .B(n15145), .Z(n15146) );
  NANDN U15895 ( .A(n14897), .B(n14896), .Z(n14901) );
  NAND U15896 ( .A(n14899), .B(n14898), .Z(n14900) );
  NAND U15897 ( .A(n14901), .B(n14900), .Z(n15040) );
  XOR U15898 ( .A(b[19]), .B(n17031), .Z(n15090) );
  NANDN U15899 ( .A(n15090), .B(n37934), .Z(n14904) );
  NANDN U15900 ( .A(n14902), .B(n37935), .Z(n14903) );
  NAND U15901 ( .A(n14904), .B(n14903), .Z(n15050) );
  XOR U15902 ( .A(b[27]), .B(a[85]), .Z(n15093) );
  NAND U15903 ( .A(n38423), .B(n15093), .Z(n14907) );
  NAND U15904 ( .A(n14905), .B(n38424), .Z(n14906) );
  NAND U15905 ( .A(n14907), .B(n14906), .Z(n15047) );
  XOR U15906 ( .A(b[5]), .B(n18980), .Z(n15096) );
  NANDN U15907 ( .A(n15096), .B(n36587), .Z(n14910) );
  NANDN U15908 ( .A(n14908), .B(n36588), .Z(n14909) );
  AND U15909 ( .A(n14910), .B(n14909), .Z(n15048) );
  XNOR U15910 ( .A(n15047), .B(n15048), .Z(n15049) );
  XNOR U15911 ( .A(n15050), .B(n15049), .Z(n15038) );
  NAND U15912 ( .A(n14911), .B(n37762), .Z(n14913) );
  XOR U15913 ( .A(b[17]), .B(a[95]), .Z(n15099) );
  NAND U15914 ( .A(n15099), .B(n37764), .Z(n14912) );
  NAND U15915 ( .A(n14913), .B(n14912), .Z(n15117) );
  XNOR U15916 ( .A(b[31]), .B(a[81]), .Z(n15102) );
  NANDN U15917 ( .A(n15102), .B(n38552), .Z(n14916) );
  NANDN U15918 ( .A(n14914), .B(n38553), .Z(n14915) );
  NAND U15919 ( .A(n14916), .B(n14915), .Z(n15114) );
  OR U15920 ( .A(n14917), .B(n36105), .Z(n14919) );
  XNOR U15921 ( .A(b[3]), .B(a[109]), .Z(n15105) );
  NANDN U15922 ( .A(n15105), .B(n36107), .Z(n14918) );
  AND U15923 ( .A(n14919), .B(n14918), .Z(n15115) );
  XNOR U15924 ( .A(n15114), .B(n15115), .Z(n15116) );
  XOR U15925 ( .A(n15117), .B(n15116), .Z(n15037) );
  XNOR U15926 ( .A(n15038), .B(n15037), .Z(n15039) );
  XNOR U15927 ( .A(n15040), .B(n15039), .Z(n15138) );
  NANDN U15928 ( .A(n14921), .B(n14920), .Z(n14925) );
  NANDN U15929 ( .A(n14923), .B(n14922), .Z(n14924) );
  NAND U15930 ( .A(n14925), .B(n14924), .Z(n15139) );
  XNOR U15931 ( .A(n15138), .B(n15139), .Z(n15140) );
  NANDN U15932 ( .A(n14927), .B(n14926), .Z(n14931) );
  NAND U15933 ( .A(n14929), .B(n14928), .Z(n14930) );
  NAND U15934 ( .A(n14931), .B(n14930), .Z(n15030) );
  OR U15935 ( .A(n14933), .B(n14932), .Z(n14937) );
  NANDN U15936 ( .A(n14935), .B(n14934), .Z(n14936) );
  NAND U15937 ( .A(n14937), .B(n14936), .Z(n15028) );
  XNOR U15938 ( .A(n15028), .B(n15027), .Z(n15029) );
  XOR U15939 ( .A(n15030), .B(n15029), .Z(n15141) );
  XOR U15940 ( .A(n15140), .B(n15141), .Z(n15152) );
  NANDN U15941 ( .A(n14947), .B(n14946), .Z(n14951) );
  NANDN U15942 ( .A(n14949), .B(n14948), .Z(n14950) );
  NAND U15943 ( .A(n14951), .B(n14950), .Z(n15135) );
  NANDN U15944 ( .A(n14957), .B(n14956), .Z(n14961) );
  NAND U15945 ( .A(n14959), .B(n14958), .Z(n14960) );
  NAND U15946 ( .A(n14961), .B(n14960), .Z(n15031) );
  NANDN U15947 ( .A(n14963), .B(n14962), .Z(n14967) );
  NAND U15948 ( .A(n14965), .B(n14964), .Z(n14966) );
  AND U15949 ( .A(n14967), .B(n14966), .Z(n15032) );
  XNOR U15950 ( .A(n15031), .B(n15032), .Z(n15033) );
  XNOR U15951 ( .A(b[9]), .B(a[103]), .Z(n15053) );
  NANDN U15952 ( .A(n15053), .B(n36925), .Z(n14970) );
  NANDN U15953 ( .A(n14968), .B(n36926), .Z(n14969) );
  NAND U15954 ( .A(n14970), .B(n14969), .Z(n15128) );
  XNOR U15955 ( .A(b[15]), .B(a[97]), .Z(n15056) );
  OR U15956 ( .A(n15056), .B(n37665), .Z(n14973) );
  NANDN U15957 ( .A(n14971), .B(n37604), .Z(n14972) );
  AND U15958 ( .A(n14973), .B(n14972), .Z(n15126) );
  XNOR U15959 ( .A(b[21]), .B(a[91]), .Z(n15059) );
  NANDN U15960 ( .A(n15059), .B(n38101), .Z(n14976) );
  NANDN U15961 ( .A(n14974), .B(n38102), .Z(n14975) );
  AND U15962 ( .A(n14976), .B(n14975), .Z(n15127) );
  XOR U15963 ( .A(n15128), .B(n15129), .Z(n15123) );
  XOR U15964 ( .A(b[11]), .B(n17812), .Z(n15062) );
  OR U15965 ( .A(n15062), .B(n37311), .Z(n14979) );
  NANDN U15966 ( .A(n14977), .B(n37218), .Z(n14978) );
  NAND U15967 ( .A(n14979), .B(n14978), .Z(n15121) );
  XOR U15968 ( .A(n1053), .B(a[99]), .Z(n15065) );
  NANDN U15969 ( .A(n15065), .B(n37424), .Z(n14982) );
  NANDN U15970 ( .A(n14980), .B(n37425), .Z(n14981) );
  AND U15971 ( .A(n14982), .B(n14981), .Z(n15120) );
  XNOR U15972 ( .A(n15121), .B(n15120), .Z(n15122) );
  XOR U15973 ( .A(n15123), .B(n15122), .Z(n15110) );
  NANDN U15974 ( .A(n1049), .B(a[111]), .Z(n14983) );
  XNOR U15975 ( .A(b[1]), .B(n14983), .Z(n14985) );
  NANDN U15976 ( .A(b[0]), .B(a[110]), .Z(n14984) );
  AND U15977 ( .A(n14985), .B(n14984), .Z(n15086) );
  NAND U15978 ( .A(n38490), .B(n14986), .Z(n14988) );
  XOR U15979 ( .A(b[29]), .B(n15562), .Z(n15069) );
  OR U15980 ( .A(n15069), .B(n1048), .Z(n14987) );
  NAND U15981 ( .A(n14988), .B(n14987), .Z(n15084) );
  NANDN U15982 ( .A(n1059), .B(a[79]), .Z(n15085) );
  XNOR U15983 ( .A(n15084), .B(n15085), .Z(n15087) );
  XOR U15984 ( .A(n15086), .B(n15087), .Z(n15108) );
  NANDN U15985 ( .A(n14989), .B(n38205), .Z(n14991) );
  XNOR U15986 ( .A(b[23]), .B(a[89]), .Z(n15075) );
  OR U15987 ( .A(n15075), .B(n38268), .Z(n14990) );
  NAND U15988 ( .A(n14991), .B(n14990), .Z(n15044) );
  XOR U15989 ( .A(b[7]), .B(a[105]), .Z(n15078) );
  NAND U15990 ( .A(n15078), .B(n36701), .Z(n14994) );
  NAND U15991 ( .A(n14992), .B(n36702), .Z(n14993) );
  NAND U15992 ( .A(n14994), .B(n14993), .Z(n15041) );
  XOR U15993 ( .A(b[25]), .B(a[87]), .Z(n15081) );
  NAND U15994 ( .A(n15081), .B(n38325), .Z(n14997) );
  NAND U15995 ( .A(n14995), .B(n38326), .Z(n14996) );
  AND U15996 ( .A(n14997), .B(n14996), .Z(n15042) );
  XNOR U15997 ( .A(n15041), .B(n15042), .Z(n15043) );
  XNOR U15998 ( .A(n15044), .B(n15043), .Z(n15109) );
  XOR U15999 ( .A(n15108), .B(n15109), .Z(n15111) );
  XNOR U16000 ( .A(n15110), .B(n15111), .Z(n15034) );
  XOR U16001 ( .A(n15033), .B(n15034), .Z(n15133) );
  XNOR U16002 ( .A(n15132), .B(n15133), .Z(n15134) );
  XNOR U16003 ( .A(n15135), .B(n15134), .Z(n15150) );
  XNOR U16004 ( .A(n15151), .B(n15150), .Z(n15153) );
  XNOR U16005 ( .A(n15152), .B(n15153), .Z(n15147) );
  XOR U16006 ( .A(n15146), .B(n15147), .Z(n15024) );
  NANDN U16007 ( .A(n14999), .B(n14998), .Z(n15003) );
  NAND U16008 ( .A(n15001), .B(n15000), .Z(n15002) );
  NAND U16009 ( .A(n15003), .B(n15002), .Z(n15021) );
  NANDN U16010 ( .A(n15005), .B(n15004), .Z(n15009) );
  OR U16011 ( .A(n15007), .B(n15006), .Z(n15008) );
  NAND U16012 ( .A(n15009), .B(n15008), .Z(n15022) );
  XNOR U16013 ( .A(n15021), .B(n15022), .Z(n15023) );
  XNOR U16014 ( .A(n15024), .B(n15023), .Z(n15016) );
  XNOR U16015 ( .A(n15015), .B(n15016), .Z(n15017) );
  XNOR U16016 ( .A(n15018), .B(n15017), .Z(n15156) );
  XNOR U16017 ( .A(n15156), .B(sreg[335]), .Z(n15158) );
  NAND U16018 ( .A(n15010), .B(sreg[334]), .Z(n15014) );
  OR U16019 ( .A(n15012), .B(n15011), .Z(n15013) );
  AND U16020 ( .A(n15014), .B(n15013), .Z(n15157) );
  XOR U16021 ( .A(n15158), .B(n15157), .Z(c[335]) );
  NANDN U16022 ( .A(n15016), .B(n15015), .Z(n15020) );
  NAND U16023 ( .A(n15018), .B(n15017), .Z(n15019) );
  NAND U16024 ( .A(n15020), .B(n15019), .Z(n15164) );
  NANDN U16025 ( .A(n15022), .B(n15021), .Z(n15026) );
  NAND U16026 ( .A(n15024), .B(n15023), .Z(n15025) );
  NAND U16027 ( .A(n15026), .B(n15025), .Z(n15162) );
  NANDN U16028 ( .A(n15032), .B(n15031), .Z(n15036) );
  NANDN U16029 ( .A(n15034), .B(n15033), .Z(n15035) );
  NAND U16030 ( .A(n15036), .B(n15035), .Z(n15178) );
  NANDN U16031 ( .A(n15042), .B(n15041), .Z(n15046) );
  NAND U16032 ( .A(n15044), .B(n15043), .Z(n15045) );
  NAND U16033 ( .A(n15046), .B(n15045), .Z(n15235) );
  NANDN U16034 ( .A(n15048), .B(n15047), .Z(n15052) );
  NAND U16035 ( .A(n15050), .B(n15049), .Z(n15051) );
  AND U16036 ( .A(n15052), .B(n15051), .Z(n15236) );
  XNOR U16037 ( .A(n15235), .B(n15236), .Z(n15237) );
  XNOR U16038 ( .A(b[9]), .B(a[104]), .Z(n15259) );
  NANDN U16039 ( .A(n15259), .B(n36925), .Z(n15055) );
  NANDN U16040 ( .A(n15053), .B(n36926), .Z(n15054) );
  NAND U16041 ( .A(n15055), .B(n15054), .Z(n15201) );
  XNOR U16042 ( .A(b[15]), .B(a[98]), .Z(n15262) );
  OR U16043 ( .A(n15262), .B(n37665), .Z(n15058) );
  NANDN U16044 ( .A(n15056), .B(n37604), .Z(n15057) );
  AND U16045 ( .A(n15058), .B(n15057), .Z(n15199) );
  XNOR U16046 ( .A(b[21]), .B(a[92]), .Z(n15265) );
  NANDN U16047 ( .A(n15265), .B(n38101), .Z(n15061) );
  NANDN U16048 ( .A(n15059), .B(n38102), .Z(n15060) );
  AND U16049 ( .A(n15061), .B(n15060), .Z(n15200) );
  XOR U16050 ( .A(n15201), .B(n15202), .Z(n15190) );
  XNOR U16051 ( .A(b[11]), .B(a[102]), .Z(n15268) );
  OR U16052 ( .A(n15268), .B(n37311), .Z(n15064) );
  NANDN U16053 ( .A(n15062), .B(n37218), .Z(n15063) );
  NAND U16054 ( .A(n15064), .B(n15063), .Z(n15188) );
  XOR U16055 ( .A(n1053), .B(a[100]), .Z(n15271) );
  NANDN U16056 ( .A(n15271), .B(n37424), .Z(n15067) );
  NANDN U16057 ( .A(n15065), .B(n37425), .Z(n15066) );
  NAND U16058 ( .A(n15067), .B(n15066), .Z(n15187) );
  XOR U16059 ( .A(n15190), .B(n15189), .Z(n15184) );
  ANDN U16060 ( .B(b[31]), .A(n15068), .Z(n15205) );
  NANDN U16061 ( .A(n15069), .B(n38490), .Z(n15071) );
  XNOR U16062 ( .A(n1058), .B(a[84]), .Z(n15277) );
  NANDN U16063 ( .A(n1048), .B(n15277), .Z(n15070) );
  NAND U16064 ( .A(n15071), .B(n15070), .Z(n15206) );
  XOR U16065 ( .A(n15205), .B(n15206), .Z(n15207) );
  NANDN U16066 ( .A(n1049), .B(a[112]), .Z(n15072) );
  XNOR U16067 ( .A(b[1]), .B(n15072), .Z(n15074) );
  NANDN U16068 ( .A(b[0]), .B(a[111]), .Z(n15073) );
  AND U16069 ( .A(n15074), .B(n15073), .Z(n15208) );
  XNOR U16070 ( .A(n15207), .B(n15208), .Z(n15181) );
  NANDN U16071 ( .A(n15075), .B(n38205), .Z(n15077) );
  XNOR U16072 ( .A(b[23]), .B(a[90]), .Z(n15280) );
  OR U16073 ( .A(n15280), .B(n38268), .Z(n15076) );
  NAND U16074 ( .A(n15077), .B(n15076), .Z(n15250) );
  XOR U16075 ( .A(b[7]), .B(a[106]), .Z(n15283) );
  NAND U16076 ( .A(n15283), .B(n36701), .Z(n15080) );
  NAND U16077 ( .A(n15078), .B(n36702), .Z(n15079) );
  NAND U16078 ( .A(n15080), .B(n15079), .Z(n15247) );
  XOR U16079 ( .A(b[25]), .B(a[88]), .Z(n15286) );
  NAND U16080 ( .A(n15286), .B(n38325), .Z(n15083) );
  NAND U16081 ( .A(n15081), .B(n38326), .Z(n15082) );
  AND U16082 ( .A(n15083), .B(n15082), .Z(n15248) );
  XNOR U16083 ( .A(n15247), .B(n15248), .Z(n15249) );
  XNOR U16084 ( .A(n15250), .B(n15249), .Z(n15182) );
  XOR U16085 ( .A(n15184), .B(n15183), .Z(n15238) );
  XNOR U16086 ( .A(n15237), .B(n15238), .Z(n15175) );
  XOR U16087 ( .A(n15176), .B(n15175), .Z(n15177) );
  XOR U16088 ( .A(n15178), .B(n15177), .Z(n15290) );
  XNOR U16089 ( .A(n15289), .B(n15290), .Z(n15292) );
  NANDN U16090 ( .A(n15085), .B(n15084), .Z(n15089) );
  NAND U16091 ( .A(n15087), .B(n15086), .Z(n15088) );
  NAND U16092 ( .A(n15089), .B(n15088), .Z(n15244) );
  XNOR U16093 ( .A(b[19]), .B(a[94]), .Z(n15211) );
  NANDN U16094 ( .A(n15211), .B(n37934), .Z(n15092) );
  NANDN U16095 ( .A(n15090), .B(n37935), .Z(n15091) );
  NAND U16096 ( .A(n15092), .B(n15091), .Z(n15256) );
  XOR U16097 ( .A(b[27]), .B(a[86]), .Z(n15214) );
  NAND U16098 ( .A(n38423), .B(n15214), .Z(n15095) );
  NAND U16099 ( .A(n15093), .B(n38424), .Z(n15094) );
  NAND U16100 ( .A(n15095), .B(n15094), .Z(n15253) );
  XNOR U16101 ( .A(b[5]), .B(a[108]), .Z(n15217) );
  NANDN U16102 ( .A(n15217), .B(n36587), .Z(n15098) );
  NANDN U16103 ( .A(n15096), .B(n36588), .Z(n15097) );
  AND U16104 ( .A(n15098), .B(n15097), .Z(n15254) );
  XNOR U16105 ( .A(n15253), .B(n15254), .Z(n15255) );
  XNOR U16106 ( .A(n15256), .B(n15255), .Z(n15241) );
  NAND U16107 ( .A(n15099), .B(n37762), .Z(n15101) );
  XOR U16108 ( .A(b[17]), .B(a[96]), .Z(n15220) );
  NAND U16109 ( .A(n15220), .B(n37764), .Z(n15100) );
  NAND U16110 ( .A(n15101), .B(n15100), .Z(n15195) );
  XOR U16111 ( .A(b[31]), .B(n15424), .Z(n15223) );
  NANDN U16112 ( .A(n15223), .B(n38552), .Z(n15104) );
  NANDN U16113 ( .A(n15102), .B(n38553), .Z(n15103) );
  AND U16114 ( .A(n15104), .B(n15103), .Z(n15193) );
  OR U16115 ( .A(n15105), .B(n36105), .Z(n15107) );
  XNOR U16116 ( .A(b[3]), .B(a[110]), .Z(n15226) );
  NANDN U16117 ( .A(n15226), .B(n36107), .Z(n15106) );
  AND U16118 ( .A(n15107), .B(n15106), .Z(n15194) );
  XOR U16119 ( .A(n15195), .B(n15196), .Z(n15242) );
  XOR U16120 ( .A(n15241), .B(n15242), .Z(n15243) );
  XNOR U16121 ( .A(n15244), .B(n15243), .Z(n15171) );
  NANDN U16122 ( .A(n15109), .B(n15108), .Z(n15113) );
  OR U16123 ( .A(n15111), .B(n15110), .Z(n15112) );
  NAND U16124 ( .A(n15113), .B(n15112), .Z(n15172) );
  XNOR U16125 ( .A(n15171), .B(n15172), .Z(n15173) );
  NANDN U16126 ( .A(n15115), .B(n15114), .Z(n15119) );
  NAND U16127 ( .A(n15117), .B(n15116), .Z(n15118) );
  NAND U16128 ( .A(n15119), .B(n15118), .Z(n15232) );
  NANDN U16129 ( .A(n15121), .B(n15120), .Z(n15125) );
  NAND U16130 ( .A(n15123), .B(n15122), .Z(n15124) );
  NAND U16131 ( .A(n15125), .B(n15124), .Z(n15229) );
  OR U16132 ( .A(n15127), .B(n15126), .Z(n15131) );
  NANDN U16133 ( .A(n15129), .B(n15128), .Z(n15130) );
  NAND U16134 ( .A(n15131), .B(n15130), .Z(n15230) );
  XNOR U16135 ( .A(n15229), .B(n15230), .Z(n15231) );
  XOR U16136 ( .A(n15232), .B(n15231), .Z(n15174) );
  XNOR U16137 ( .A(n15173), .B(n15174), .Z(n15291) );
  XOR U16138 ( .A(n15292), .B(n15291), .Z(n15296) );
  NANDN U16139 ( .A(n15133), .B(n15132), .Z(n15137) );
  NAND U16140 ( .A(n15135), .B(n15134), .Z(n15136) );
  NAND U16141 ( .A(n15137), .B(n15136), .Z(n15293) );
  NANDN U16142 ( .A(n15139), .B(n15138), .Z(n15143) );
  NAND U16143 ( .A(n15141), .B(n15140), .Z(n15142) );
  NAND U16144 ( .A(n15143), .B(n15142), .Z(n15294) );
  XNOR U16145 ( .A(n15293), .B(n15294), .Z(n15295) );
  XNOR U16146 ( .A(n15296), .B(n15295), .Z(n15168) );
  NANDN U16147 ( .A(n15145), .B(n15144), .Z(n15149) );
  NANDN U16148 ( .A(n15147), .B(n15146), .Z(n15148) );
  NAND U16149 ( .A(n15149), .B(n15148), .Z(n15166) );
  OR U16150 ( .A(n15151), .B(n15150), .Z(n15155) );
  OR U16151 ( .A(n15153), .B(n15152), .Z(n15154) );
  AND U16152 ( .A(n15155), .B(n15154), .Z(n15165) );
  XNOR U16153 ( .A(n15166), .B(n15165), .Z(n15167) );
  XNOR U16154 ( .A(n15168), .B(n15167), .Z(n15161) );
  XOR U16155 ( .A(n15162), .B(n15161), .Z(n15163) );
  XNOR U16156 ( .A(n15164), .B(n15163), .Z(n15299) );
  XNOR U16157 ( .A(n15299), .B(sreg[336]), .Z(n15301) );
  NAND U16158 ( .A(n15156), .B(sreg[335]), .Z(n15160) );
  OR U16159 ( .A(n15158), .B(n15157), .Z(n15159) );
  AND U16160 ( .A(n15160), .B(n15159), .Z(n15300) );
  XOR U16161 ( .A(n15301), .B(n15300), .Z(c[336]) );
  NANDN U16162 ( .A(n15166), .B(n15165), .Z(n15170) );
  NANDN U16163 ( .A(n15168), .B(n15167), .Z(n15169) );
  NAND U16164 ( .A(n15170), .B(n15169), .Z(n15305) );
  NAND U16165 ( .A(n15176), .B(n15175), .Z(n15180) );
  NAND U16166 ( .A(n15178), .B(n15177), .Z(n15179) );
  NAND U16167 ( .A(n15180), .B(n15179), .Z(n15323) );
  XNOR U16168 ( .A(n15322), .B(n15323), .Z(n15324) );
  OR U16169 ( .A(n15182), .B(n15181), .Z(n15186) );
  NANDN U16170 ( .A(n15184), .B(n15183), .Z(n15185) );
  NAND U16171 ( .A(n15186), .B(n15185), .Z(n15440) );
  OR U16172 ( .A(n15188), .B(n15187), .Z(n15192) );
  NAND U16173 ( .A(n15190), .B(n15189), .Z(n15191) );
  NAND U16174 ( .A(n15192), .B(n15191), .Z(n15378) );
  OR U16175 ( .A(n15194), .B(n15193), .Z(n15198) );
  NANDN U16176 ( .A(n15196), .B(n15195), .Z(n15197) );
  NAND U16177 ( .A(n15198), .B(n15197), .Z(n15377) );
  OR U16178 ( .A(n15200), .B(n15199), .Z(n15204) );
  NANDN U16179 ( .A(n15202), .B(n15201), .Z(n15203) );
  NAND U16180 ( .A(n15204), .B(n15203), .Z(n15376) );
  XOR U16181 ( .A(n15378), .B(n15379), .Z(n15438) );
  OR U16182 ( .A(n15206), .B(n15205), .Z(n15210) );
  NANDN U16183 ( .A(n15208), .B(n15207), .Z(n15209) );
  NAND U16184 ( .A(n15210), .B(n15209), .Z(n15390) );
  XNOR U16185 ( .A(b[19]), .B(a[95]), .Z(n15334) );
  NANDN U16186 ( .A(n15334), .B(n37934), .Z(n15213) );
  NANDN U16187 ( .A(n15211), .B(n37935), .Z(n15212) );
  NAND U16188 ( .A(n15213), .B(n15212), .Z(n15403) );
  XOR U16189 ( .A(b[27]), .B(a[87]), .Z(n15337) );
  NAND U16190 ( .A(n38423), .B(n15337), .Z(n15216) );
  NAND U16191 ( .A(n15214), .B(n38424), .Z(n15215) );
  NAND U16192 ( .A(n15216), .B(n15215), .Z(n15400) );
  XNOR U16193 ( .A(b[5]), .B(a[109]), .Z(n15340) );
  NANDN U16194 ( .A(n15340), .B(n36587), .Z(n15219) );
  NANDN U16195 ( .A(n15217), .B(n36588), .Z(n15218) );
  AND U16196 ( .A(n15219), .B(n15218), .Z(n15401) );
  XNOR U16197 ( .A(n15400), .B(n15401), .Z(n15402) );
  XNOR U16198 ( .A(n15403), .B(n15402), .Z(n15389) );
  NAND U16199 ( .A(n15220), .B(n37762), .Z(n15222) );
  XOR U16200 ( .A(b[17]), .B(a[97]), .Z(n15343) );
  NAND U16201 ( .A(n15343), .B(n37764), .Z(n15221) );
  NAND U16202 ( .A(n15222), .B(n15221), .Z(n15361) );
  XOR U16203 ( .A(b[31]), .B(n15562), .Z(n15346) );
  NANDN U16204 ( .A(n15346), .B(n38552), .Z(n15225) );
  NANDN U16205 ( .A(n15223), .B(n38553), .Z(n15224) );
  NAND U16206 ( .A(n15225), .B(n15224), .Z(n15358) );
  OR U16207 ( .A(n15226), .B(n36105), .Z(n15228) );
  XNOR U16208 ( .A(b[3]), .B(a[111]), .Z(n15349) );
  NANDN U16209 ( .A(n15349), .B(n36107), .Z(n15227) );
  AND U16210 ( .A(n15228), .B(n15227), .Z(n15359) );
  XNOR U16211 ( .A(n15358), .B(n15359), .Z(n15360) );
  XOR U16212 ( .A(n15361), .B(n15360), .Z(n15388) );
  XOR U16213 ( .A(n15389), .B(n15388), .Z(n15391) );
  XOR U16214 ( .A(n15390), .B(n15391), .Z(n15437) );
  XOR U16215 ( .A(n15438), .B(n15437), .Z(n15439) );
  XNOR U16216 ( .A(n15440), .B(n15439), .Z(n15319) );
  NANDN U16217 ( .A(n15230), .B(n15229), .Z(n15234) );
  NANDN U16218 ( .A(n15232), .B(n15231), .Z(n15233) );
  NAND U16219 ( .A(n15234), .B(n15233), .Z(n15316) );
  NANDN U16220 ( .A(n15236), .B(n15235), .Z(n15240) );
  NANDN U16221 ( .A(n15238), .B(n15237), .Z(n15239) );
  NAND U16222 ( .A(n15240), .B(n15239), .Z(n15446) );
  OR U16223 ( .A(n15242), .B(n15241), .Z(n15246) );
  NAND U16224 ( .A(n15244), .B(n15243), .Z(n15245) );
  NAND U16225 ( .A(n15246), .B(n15245), .Z(n15443) );
  NANDN U16226 ( .A(n15248), .B(n15247), .Z(n15252) );
  NAND U16227 ( .A(n15250), .B(n15249), .Z(n15251) );
  NAND U16228 ( .A(n15252), .B(n15251), .Z(n15382) );
  NANDN U16229 ( .A(n15254), .B(n15253), .Z(n15258) );
  NAND U16230 ( .A(n15256), .B(n15255), .Z(n15257) );
  AND U16231 ( .A(n15258), .B(n15257), .Z(n15383) );
  XNOR U16232 ( .A(n15382), .B(n15383), .Z(n15384) );
  XNOR U16233 ( .A(b[9]), .B(a[105]), .Z(n15406) );
  NANDN U16234 ( .A(n15406), .B(n36925), .Z(n15261) );
  NANDN U16235 ( .A(n15259), .B(n36926), .Z(n15260) );
  NAND U16236 ( .A(n15261), .B(n15260), .Z(n15366) );
  XOR U16237 ( .A(b[15]), .B(n17884), .Z(n15409) );
  OR U16238 ( .A(n15409), .B(n37665), .Z(n15264) );
  NANDN U16239 ( .A(n15262), .B(n37604), .Z(n15263) );
  AND U16240 ( .A(n15264), .B(n15263), .Z(n15364) );
  XOR U16241 ( .A(b[21]), .B(n17031), .Z(n15412) );
  NANDN U16242 ( .A(n15412), .B(n38101), .Z(n15267) );
  NANDN U16243 ( .A(n15265), .B(n38102), .Z(n15266) );
  AND U16244 ( .A(n15267), .B(n15266), .Z(n15365) );
  XOR U16245 ( .A(n15366), .B(n15367), .Z(n15355) );
  XNOR U16246 ( .A(b[11]), .B(a[103]), .Z(n15415) );
  OR U16247 ( .A(n15415), .B(n37311), .Z(n15270) );
  NANDN U16248 ( .A(n15268), .B(n37218), .Z(n15269) );
  NAND U16249 ( .A(n15270), .B(n15269), .Z(n15353) );
  XOR U16250 ( .A(n1053), .B(a[101]), .Z(n15418) );
  NANDN U16251 ( .A(n15418), .B(n37424), .Z(n15273) );
  NANDN U16252 ( .A(n15271), .B(n37425), .Z(n15272) );
  AND U16253 ( .A(n15273), .B(n15272), .Z(n15352) );
  XNOR U16254 ( .A(n15353), .B(n15352), .Z(n15354) );
  XOR U16255 ( .A(n15355), .B(n15354), .Z(n15372) );
  NANDN U16256 ( .A(n1049), .B(a[113]), .Z(n15274) );
  XNOR U16257 ( .A(b[1]), .B(n15274), .Z(n15276) );
  NANDN U16258 ( .A(b[0]), .B(a[112]), .Z(n15275) );
  AND U16259 ( .A(n15276), .B(n15275), .Z(n15330) );
  NAND U16260 ( .A(n15277), .B(n38490), .Z(n15279) );
  XNOR U16261 ( .A(b[29]), .B(a[85]), .Z(n15425) );
  OR U16262 ( .A(n15425), .B(n1048), .Z(n15278) );
  NAND U16263 ( .A(n15279), .B(n15278), .Z(n15328) );
  NANDN U16264 ( .A(n1059), .B(a[81]), .Z(n15329) );
  XNOR U16265 ( .A(n15328), .B(n15329), .Z(n15331) );
  XOR U16266 ( .A(n15330), .B(n15331), .Z(n15370) );
  NANDN U16267 ( .A(n15280), .B(n38205), .Z(n15282) );
  XNOR U16268 ( .A(b[23]), .B(a[91]), .Z(n15428) );
  OR U16269 ( .A(n15428), .B(n38268), .Z(n15281) );
  NAND U16270 ( .A(n15282), .B(n15281), .Z(n15397) );
  XNOR U16271 ( .A(b[7]), .B(a[107]), .Z(n15431) );
  NANDN U16272 ( .A(n15431), .B(n36701), .Z(n15285) );
  NAND U16273 ( .A(n15283), .B(n36702), .Z(n15284) );
  NAND U16274 ( .A(n15285), .B(n15284), .Z(n15394) );
  XOR U16275 ( .A(b[25]), .B(a[89]), .Z(n15434) );
  NAND U16276 ( .A(n15434), .B(n38325), .Z(n15288) );
  NAND U16277 ( .A(n15286), .B(n38326), .Z(n15287) );
  AND U16278 ( .A(n15288), .B(n15287), .Z(n15395) );
  XNOR U16279 ( .A(n15394), .B(n15395), .Z(n15396) );
  XNOR U16280 ( .A(n15397), .B(n15396), .Z(n15371) );
  XOR U16281 ( .A(n15370), .B(n15371), .Z(n15373) );
  XNOR U16282 ( .A(n15372), .B(n15373), .Z(n15385) );
  XOR U16283 ( .A(n15384), .B(n15385), .Z(n15444) );
  XNOR U16284 ( .A(n15443), .B(n15444), .Z(n15445) );
  XOR U16285 ( .A(n15446), .B(n15445), .Z(n15317) );
  XNOR U16286 ( .A(n15316), .B(n15317), .Z(n15318) );
  XOR U16287 ( .A(n15319), .B(n15318), .Z(n15325) );
  XOR U16288 ( .A(n15324), .B(n15325), .Z(n15312) );
  NANDN U16289 ( .A(n15294), .B(n15293), .Z(n15298) );
  NANDN U16290 ( .A(n15296), .B(n15295), .Z(n15297) );
  NAND U16291 ( .A(n15298), .B(n15297), .Z(n15311) );
  XNOR U16292 ( .A(n15310), .B(n15311), .Z(n15313) );
  XOR U16293 ( .A(n15312), .B(n15313), .Z(n15304) );
  XOR U16294 ( .A(n15305), .B(n15304), .Z(n15306) );
  XNOR U16295 ( .A(n15307), .B(n15306), .Z(n15449) );
  XNOR U16296 ( .A(n15449), .B(sreg[337]), .Z(n15451) );
  NAND U16297 ( .A(n15299), .B(sreg[336]), .Z(n15303) );
  OR U16298 ( .A(n15301), .B(n15300), .Z(n15302) );
  AND U16299 ( .A(n15303), .B(n15302), .Z(n15450) );
  XOR U16300 ( .A(n15451), .B(n15450), .Z(c[337]) );
  NAND U16301 ( .A(n15305), .B(n15304), .Z(n15309) );
  NAND U16302 ( .A(n15307), .B(n15306), .Z(n15308) );
  NAND U16303 ( .A(n15309), .B(n15308), .Z(n15457) );
  NANDN U16304 ( .A(n15311), .B(n15310), .Z(n15315) );
  NAND U16305 ( .A(n15313), .B(n15312), .Z(n15314) );
  NAND U16306 ( .A(n15315), .B(n15314), .Z(n15455) );
  NANDN U16307 ( .A(n15317), .B(n15316), .Z(n15321) );
  NAND U16308 ( .A(n15319), .B(n15318), .Z(n15320) );
  NAND U16309 ( .A(n15321), .B(n15320), .Z(n15460) );
  NANDN U16310 ( .A(n15323), .B(n15322), .Z(n15327) );
  NAND U16311 ( .A(n15325), .B(n15324), .Z(n15326) );
  AND U16312 ( .A(n15327), .B(n15326), .Z(n15461) );
  XNOR U16313 ( .A(n15460), .B(n15461), .Z(n15462) );
  NANDN U16314 ( .A(n15329), .B(n15328), .Z(n15333) );
  NAND U16315 ( .A(n15331), .B(n15330), .Z(n15332) );
  NAND U16316 ( .A(n15333), .B(n15332), .Z(n15529) );
  XNOR U16317 ( .A(b[19]), .B(a[96]), .Z(n15496) );
  NANDN U16318 ( .A(n15496), .B(n37934), .Z(n15336) );
  NANDN U16319 ( .A(n15334), .B(n37935), .Z(n15335) );
  NAND U16320 ( .A(n15336), .B(n15335), .Z(n15541) );
  XOR U16321 ( .A(b[27]), .B(a[88]), .Z(n15499) );
  NAND U16322 ( .A(n38423), .B(n15499), .Z(n15339) );
  NAND U16323 ( .A(n15337), .B(n38424), .Z(n15338) );
  NAND U16324 ( .A(n15339), .B(n15338), .Z(n15538) );
  XNOR U16325 ( .A(b[5]), .B(a[110]), .Z(n15502) );
  NANDN U16326 ( .A(n15502), .B(n36587), .Z(n15342) );
  NANDN U16327 ( .A(n15340), .B(n36588), .Z(n15341) );
  AND U16328 ( .A(n15342), .B(n15341), .Z(n15539) );
  XNOR U16329 ( .A(n15538), .B(n15539), .Z(n15540) );
  XNOR U16330 ( .A(n15541), .B(n15540), .Z(n15526) );
  NAND U16331 ( .A(n15343), .B(n37762), .Z(n15345) );
  XOR U16332 ( .A(b[17]), .B(a[98]), .Z(n15505) );
  NAND U16333 ( .A(n15505), .B(n37764), .Z(n15344) );
  NAND U16334 ( .A(n15345), .B(n15344), .Z(n15480) );
  XNOR U16335 ( .A(b[31]), .B(a[84]), .Z(n15508) );
  NANDN U16336 ( .A(n15508), .B(n38552), .Z(n15348) );
  NANDN U16337 ( .A(n15346), .B(n38553), .Z(n15347) );
  AND U16338 ( .A(n15348), .B(n15347), .Z(n15478) );
  OR U16339 ( .A(n15349), .B(n36105), .Z(n15351) );
  XNOR U16340 ( .A(b[3]), .B(a[112]), .Z(n15511) );
  NANDN U16341 ( .A(n15511), .B(n36107), .Z(n15350) );
  AND U16342 ( .A(n15351), .B(n15350), .Z(n15479) );
  XOR U16343 ( .A(n15480), .B(n15481), .Z(n15527) );
  XOR U16344 ( .A(n15526), .B(n15527), .Z(n15528) );
  XNOR U16345 ( .A(n15529), .B(n15528), .Z(n15575) );
  NANDN U16346 ( .A(n15353), .B(n15352), .Z(n15357) );
  NAND U16347 ( .A(n15355), .B(n15354), .Z(n15356) );
  NAND U16348 ( .A(n15357), .B(n15356), .Z(n15517) );
  NANDN U16349 ( .A(n15359), .B(n15358), .Z(n15363) );
  NAND U16350 ( .A(n15361), .B(n15360), .Z(n15362) );
  NAND U16351 ( .A(n15363), .B(n15362), .Z(n15515) );
  OR U16352 ( .A(n15365), .B(n15364), .Z(n15369) );
  NANDN U16353 ( .A(n15367), .B(n15366), .Z(n15368) );
  NAND U16354 ( .A(n15369), .B(n15368), .Z(n15514) );
  XNOR U16355 ( .A(n15517), .B(n15516), .Z(n15576) );
  XOR U16356 ( .A(n15575), .B(n15576), .Z(n15578) );
  NANDN U16357 ( .A(n15371), .B(n15370), .Z(n15375) );
  OR U16358 ( .A(n15373), .B(n15372), .Z(n15374) );
  NAND U16359 ( .A(n15375), .B(n15374), .Z(n15577) );
  XOR U16360 ( .A(n15578), .B(n15577), .Z(n15595) );
  OR U16361 ( .A(n15377), .B(n15376), .Z(n15381) );
  NANDN U16362 ( .A(n15379), .B(n15378), .Z(n15380) );
  NAND U16363 ( .A(n15381), .B(n15380), .Z(n15594) );
  NANDN U16364 ( .A(n15383), .B(n15382), .Z(n15387) );
  NANDN U16365 ( .A(n15385), .B(n15384), .Z(n15386) );
  NAND U16366 ( .A(n15387), .B(n15386), .Z(n15583) );
  NANDN U16367 ( .A(n15389), .B(n15388), .Z(n15393) );
  OR U16368 ( .A(n15391), .B(n15390), .Z(n15392) );
  NAND U16369 ( .A(n15393), .B(n15392), .Z(n15582) );
  NANDN U16370 ( .A(n15395), .B(n15394), .Z(n15399) );
  NAND U16371 ( .A(n15397), .B(n15396), .Z(n15398) );
  NAND U16372 ( .A(n15399), .B(n15398), .Z(n15520) );
  NANDN U16373 ( .A(n15401), .B(n15400), .Z(n15405) );
  NAND U16374 ( .A(n15403), .B(n15402), .Z(n15404) );
  AND U16375 ( .A(n15405), .B(n15404), .Z(n15521) );
  XNOR U16376 ( .A(n15520), .B(n15521), .Z(n15522) );
  XNOR U16377 ( .A(b[9]), .B(a[106]), .Z(n15544) );
  NANDN U16378 ( .A(n15544), .B(n36925), .Z(n15408) );
  NANDN U16379 ( .A(n15406), .B(n36926), .Z(n15407) );
  NAND U16380 ( .A(n15408), .B(n15407), .Z(n15486) );
  XNOR U16381 ( .A(b[15]), .B(a[100]), .Z(n15547) );
  OR U16382 ( .A(n15547), .B(n37665), .Z(n15411) );
  NANDN U16383 ( .A(n15409), .B(n37604), .Z(n15410) );
  AND U16384 ( .A(n15411), .B(n15410), .Z(n15484) );
  XNOR U16385 ( .A(b[21]), .B(a[94]), .Z(n15550) );
  NANDN U16386 ( .A(n15550), .B(n38101), .Z(n15414) );
  NANDN U16387 ( .A(n15412), .B(n38102), .Z(n15413) );
  AND U16388 ( .A(n15414), .B(n15413), .Z(n15485) );
  XOR U16389 ( .A(n15486), .B(n15487), .Z(n15475) );
  XNOR U16390 ( .A(b[11]), .B(a[104]), .Z(n15553) );
  OR U16391 ( .A(n15553), .B(n37311), .Z(n15417) );
  NANDN U16392 ( .A(n15415), .B(n37218), .Z(n15416) );
  NAND U16393 ( .A(n15417), .B(n15416), .Z(n15473) );
  XOR U16394 ( .A(n1053), .B(a[102]), .Z(n15556) );
  NANDN U16395 ( .A(n15556), .B(n37424), .Z(n15420) );
  NANDN U16396 ( .A(n15418), .B(n37425), .Z(n15419) );
  NAND U16397 ( .A(n15420), .B(n15419), .Z(n15472) );
  XOR U16398 ( .A(n15475), .B(n15474), .Z(n15469) );
  NANDN U16399 ( .A(n1049), .B(a[114]), .Z(n15421) );
  XNOR U16400 ( .A(b[1]), .B(n15421), .Z(n15423) );
  IV U16401 ( .A(a[113]), .Z(n19909) );
  NANDN U16402 ( .A(n19909), .B(n1049), .Z(n15422) );
  AND U16403 ( .A(n15423), .B(n15422), .Z(n15493) );
  ANDN U16404 ( .B(b[31]), .A(n15424), .Z(n15490) );
  NANDN U16405 ( .A(n15425), .B(n38490), .Z(n15427) );
  XNOR U16406 ( .A(b[29]), .B(a[86]), .Z(n15563) );
  OR U16407 ( .A(n15563), .B(n1048), .Z(n15426) );
  NAND U16408 ( .A(n15427), .B(n15426), .Z(n15491) );
  XOR U16409 ( .A(n15490), .B(n15491), .Z(n15492) );
  XNOR U16410 ( .A(n15493), .B(n15492), .Z(n15466) );
  NANDN U16411 ( .A(n15428), .B(n38205), .Z(n15430) );
  XNOR U16412 ( .A(b[23]), .B(a[92]), .Z(n15566) );
  OR U16413 ( .A(n15566), .B(n38268), .Z(n15429) );
  NAND U16414 ( .A(n15430), .B(n15429), .Z(n15535) );
  XOR U16415 ( .A(b[7]), .B(a[108]), .Z(n15569) );
  NAND U16416 ( .A(n15569), .B(n36701), .Z(n15433) );
  NANDN U16417 ( .A(n15431), .B(n36702), .Z(n15432) );
  NAND U16418 ( .A(n15433), .B(n15432), .Z(n15532) );
  XOR U16419 ( .A(b[25]), .B(a[90]), .Z(n15572) );
  NAND U16420 ( .A(n15572), .B(n38325), .Z(n15436) );
  NAND U16421 ( .A(n15434), .B(n38326), .Z(n15435) );
  AND U16422 ( .A(n15436), .B(n15435), .Z(n15533) );
  XNOR U16423 ( .A(n15532), .B(n15533), .Z(n15534) );
  XNOR U16424 ( .A(n15535), .B(n15534), .Z(n15467) );
  XOR U16425 ( .A(n15469), .B(n15468), .Z(n15523) );
  XNOR U16426 ( .A(n15522), .B(n15523), .Z(n15581) );
  XNOR U16427 ( .A(n15582), .B(n15581), .Z(n15584) );
  XNOR U16428 ( .A(n15583), .B(n15584), .Z(n15593) );
  XOR U16429 ( .A(n15594), .B(n15593), .Z(n15596) );
  NAND U16430 ( .A(n15438), .B(n15437), .Z(n15442) );
  NAND U16431 ( .A(n15440), .B(n15439), .Z(n15441) );
  NAND U16432 ( .A(n15442), .B(n15441), .Z(n15588) );
  NANDN U16433 ( .A(n15444), .B(n15443), .Z(n15448) );
  NAND U16434 ( .A(n15446), .B(n15445), .Z(n15447) );
  AND U16435 ( .A(n15448), .B(n15447), .Z(n15587) );
  XNOR U16436 ( .A(n15588), .B(n15587), .Z(n15589) );
  XOR U16437 ( .A(n15590), .B(n15589), .Z(n15463) );
  XOR U16438 ( .A(n15462), .B(n15463), .Z(n15454) );
  XOR U16439 ( .A(n15455), .B(n15454), .Z(n15456) );
  XNOR U16440 ( .A(n15457), .B(n15456), .Z(n15599) );
  XNOR U16441 ( .A(n15599), .B(sreg[338]), .Z(n15601) );
  NAND U16442 ( .A(n15449), .B(sreg[337]), .Z(n15453) );
  OR U16443 ( .A(n15451), .B(n15450), .Z(n15452) );
  AND U16444 ( .A(n15453), .B(n15452), .Z(n15600) );
  XOR U16445 ( .A(n15601), .B(n15600), .Z(c[338]) );
  NAND U16446 ( .A(n15455), .B(n15454), .Z(n15459) );
  NAND U16447 ( .A(n15457), .B(n15456), .Z(n15458) );
  NAND U16448 ( .A(n15459), .B(n15458), .Z(n15607) );
  NANDN U16449 ( .A(n15461), .B(n15460), .Z(n15465) );
  NAND U16450 ( .A(n15463), .B(n15462), .Z(n15464) );
  NAND U16451 ( .A(n15465), .B(n15464), .Z(n15605) );
  OR U16452 ( .A(n15467), .B(n15466), .Z(n15471) );
  NANDN U16453 ( .A(n15469), .B(n15468), .Z(n15470) );
  NAND U16454 ( .A(n15471), .B(n15470), .Z(n15725) );
  OR U16455 ( .A(n15473), .B(n15472), .Z(n15477) );
  NAND U16456 ( .A(n15475), .B(n15474), .Z(n15476) );
  NAND U16457 ( .A(n15477), .B(n15476), .Z(n15664) );
  OR U16458 ( .A(n15479), .B(n15478), .Z(n15483) );
  NANDN U16459 ( .A(n15481), .B(n15480), .Z(n15482) );
  NAND U16460 ( .A(n15483), .B(n15482), .Z(n15663) );
  OR U16461 ( .A(n15485), .B(n15484), .Z(n15489) );
  NANDN U16462 ( .A(n15487), .B(n15486), .Z(n15488) );
  NAND U16463 ( .A(n15489), .B(n15488), .Z(n15662) );
  XOR U16464 ( .A(n15664), .B(n15665), .Z(n15723) );
  OR U16465 ( .A(n15491), .B(n15490), .Z(n15495) );
  NANDN U16466 ( .A(n15493), .B(n15492), .Z(n15494) );
  NAND U16467 ( .A(n15495), .B(n15494), .Z(n15677) );
  XNOR U16468 ( .A(b[19]), .B(a[97]), .Z(n15644) );
  NANDN U16469 ( .A(n15644), .B(n37934), .Z(n15498) );
  NANDN U16470 ( .A(n15496), .B(n37935), .Z(n15497) );
  NAND U16471 ( .A(n15498), .B(n15497), .Z(n15689) );
  XOR U16472 ( .A(b[27]), .B(a[89]), .Z(n15647) );
  NAND U16473 ( .A(n38423), .B(n15647), .Z(n15501) );
  NAND U16474 ( .A(n15499), .B(n38424), .Z(n15500) );
  NAND U16475 ( .A(n15501), .B(n15500), .Z(n15686) );
  XNOR U16476 ( .A(b[5]), .B(a[111]), .Z(n15650) );
  NANDN U16477 ( .A(n15650), .B(n36587), .Z(n15504) );
  NANDN U16478 ( .A(n15502), .B(n36588), .Z(n15503) );
  AND U16479 ( .A(n15504), .B(n15503), .Z(n15687) );
  XNOR U16480 ( .A(n15686), .B(n15687), .Z(n15688) );
  XNOR U16481 ( .A(n15689), .B(n15688), .Z(n15674) );
  NAND U16482 ( .A(n15505), .B(n37762), .Z(n15507) );
  XNOR U16483 ( .A(b[17]), .B(a[99]), .Z(n15653) );
  NANDN U16484 ( .A(n15653), .B(n37764), .Z(n15506) );
  NAND U16485 ( .A(n15507), .B(n15506), .Z(n15628) );
  XNOR U16486 ( .A(b[31]), .B(a[85]), .Z(n15656) );
  NANDN U16487 ( .A(n15656), .B(n38552), .Z(n15510) );
  NANDN U16488 ( .A(n15508), .B(n38553), .Z(n15509) );
  AND U16489 ( .A(n15510), .B(n15509), .Z(n15626) );
  OR U16490 ( .A(n15511), .B(n36105), .Z(n15513) );
  XOR U16491 ( .A(b[3]), .B(n19909), .Z(n15659) );
  NANDN U16492 ( .A(n15659), .B(n36107), .Z(n15512) );
  AND U16493 ( .A(n15513), .B(n15512), .Z(n15627) );
  XOR U16494 ( .A(n15628), .B(n15629), .Z(n15675) );
  XOR U16495 ( .A(n15674), .B(n15675), .Z(n15676) );
  XNOR U16496 ( .A(n15677), .B(n15676), .Z(n15722) );
  XOR U16497 ( .A(n15723), .B(n15722), .Z(n15724) );
  XNOR U16498 ( .A(n15725), .B(n15724), .Z(n15741) );
  OR U16499 ( .A(n15515), .B(n15514), .Z(n15519) );
  NAND U16500 ( .A(n15517), .B(n15516), .Z(n15518) );
  NAND U16501 ( .A(n15519), .B(n15518), .Z(n15739) );
  NANDN U16502 ( .A(n15521), .B(n15520), .Z(n15525) );
  NANDN U16503 ( .A(n15523), .B(n15522), .Z(n15524) );
  NAND U16504 ( .A(n15525), .B(n15524), .Z(n15728) );
  OR U16505 ( .A(n15527), .B(n15526), .Z(n15531) );
  NAND U16506 ( .A(n15529), .B(n15528), .Z(n15530) );
  NAND U16507 ( .A(n15531), .B(n15530), .Z(n15727) );
  NANDN U16508 ( .A(n15533), .B(n15532), .Z(n15537) );
  NAND U16509 ( .A(n15535), .B(n15534), .Z(n15536) );
  NAND U16510 ( .A(n15537), .B(n15536), .Z(n15668) );
  NANDN U16511 ( .A(n15539), .B(n15538), .Z(n15543) );
  NAND U16512 ( .A(n15541), .B(n15540), .Z(n15542) );
  AND U16513 ( .A(n15543), .B(n15542), .Z(n15669) );
  XNOR U16514 ( .A(n15668), .B(n15669), .Z(n15670) );
  XOR U16515 ( .A(b[9]), .B(n18980), .Z(n15692) );
  NANDN U16516 ( .A(n15692), .B(n36925), .Z(n15546) );
  NANDN U16517 ( .A(n15544), .B(n36926), .Z(n15545) );
  NAND U16518 ( .A(n15546), .B(n15545), .Z(n15634) );
  XOR U16519 ( .A(b[15]), .B(n17812), .Z(n15695) );
  OR U16520 ( .A(n15695), .B(n37665), .Z(n15549) );
  NANDN U16521 ( .A(n15547), .B(n37604), .Z(n15548) );
  AND U16522 ( .A(n15549), .B(n15548), .Z(n15632) );
  XNOR U16523 ( .A(b[21]), .B(a[95]), .Z(n15698) );
  NANDN U16524 ( .A(n15698), .B(n38101), .Z(n15552) );
  NANDN U16525 ( .A(n15550), .B(n38102), .Z(n15551) );
  AND U16526 ( .A(n15552), .B(n15551), .Z(n15633) );
  XOR U16527 ( .A(n15634), .B(n15635), .Z(n15623) );
  XNOR U16528 ( .A(b[11]), .B(a[105]), .Z(n15701) );
  OR U16529 ( .A(n15701), .B(n37311), .Z(n15555) );
  NANDN U16530 ( .A(n15553), .B(n37218), .Z(n15554) );
  NAND U16531 ( .A(n15555), .B(n15554), .Z(n15621) );
  XOR U16532 ( .A(n1053), .B(a[103]), .Z(n15704) );
  NANDN U16533 ( .A(n15704), .B(n37424), .Z(n15558) );
  NANDN U16534 ( .A(n15556), .B(n37425), .Z(n15557) );
  NAND U16535 ( .A(n15558), .B(n15557), .Z(n15620) );
  XOR U16536 ( .A(n15623), .B(n15622), .Z(n15617) );
  NANDN U16537 ( .A(n1049), .B(a[115]), .Z(n15559) );
  XNOR U16538 ( .A(b[1]), .B(n15559), .Z(n15561) );
  NANDN U16539 ( .A(b[0]), .B(a[114]), .Z(n15560) );
  AND U16540 ( .A(n15561), .B(n15560), .Z(n15641) );
  ANDN U16541 ( .B(b[31]), .A(n15562), .Z(n15638) );
  NANDN U16542 ( .A(n15563), .B(n38490), .Z(n15565) );
  XNOR U16543 ( .A(n1058), .B(a[87]), .Z(n15710) );
  NANDN U16544 ( .A(n1048), .B(n15710), .Z(n15564) );
  NAND U16545 ( .A(n15565), .B(n15564), .Z(n15639) );
  XOR U16546 ( .A(n15638), .B(n15639), .Z(n15640) );
  XNOR U16547 ( .A(n15641), .B(n15640), .Z(n15614) );
  NANDN U16548 ( .A(n15566), .B(n38205), .Z(n15568) );
  XOR U16549 ( .A(b[23]), .B(n17031), .Z(n15713) );
  OR U16550 ( .A(n15713), .B(n38268), .Z(n15567) );
  NAND U16551 ( .A(n15568), .B(n15567), .Z(n15683) );
  XOR U16552 ( .A(b[7]), .B(a[109]), .Z(n15716) );
  NAND U16553 ( .A(n15716), .B(n36701), .Z(n15571) );
  NAND U16554 ( .A(n15569), .B(n36702), .Z(n15570) );
  NAND U16555 ( .A(n15571), .B(n15570), .Z(n15680) );
  XOR U16556 ( .A(b[25]), .B(a[91]), .Z(n15719) );
  NAND U16557 ( .A(n15719), .B(n38325), .Z(n15574) );
  NAND U16558 ( .A(n15572), .B(n38326), .Z(n15573) );
  AND U16559 ( .A(n15574), .B(n15573), .Z(n15681) );
  XNOR U16560 ( .A(n15680), .B(n15681), .Z(n15682) );
  XNOR U16561 ( .A(n15683), .B(n15682), .Z(n15615) );
  XOR U16562 ( .A(n15617), .B(n15616), .Z(n15671) );
  XNOR U16563 ( .A(n15670), .B(n15671), .Z(n15726) );
  XNOR U16564 ( .A(n15727), .B(n15726), .Z(n15729) );
  XNOR U16565 ( .A(n15728), .B(n15729), .Z(n15738) );
  XNOR U16566 ( .A(n15739), .B(n15738), .Z(n15740) );
  XOR U16567 ( .A(n15741), .B(n15740), .Z(n15735) );
  NANDN U16568 ( .A(n15576), .B(n15575), .Z(n15580) );
  OR U16569 ( .A(n15578), .B(n15577), .Z(n15579) );
  NAND U16570 ( .A(n15580), .B(n15579), .Z(n15732) );
  NAND U16571 ( .A(n15582), .B(n15581), .Z(n15586) );
  NANDN U16572 ( .A(n15584), .B(n15583), .Z(n15585) );
  NAND U16573 ( .A(n15586), .B(n15585), .Z(n15733) );
  XNOR U16574 ( .A(n15732), .B(n15733), .Z(n15734) );
  XNOR U16575 ( .A(n15735), .B(n15734), .Z(n15611) );
  NANDN U16576 ( .A(n15588), .B(n15587), .Z(n15592) );
  NAND U16577 ( .A(n15590), .B(n15589), .Z(n15591) );
  NAND U16578 ( .A(n15592), .B(n15591), .Z(n15608) );
  NANDN U16579 ( .A(n15594), .B(n15593), .Z(n15598) );
  OR U16580 ( .A(n15596), .B(n15595), .Z(n15597) );
  NAND U16581 ( .A(n15598), .B(n15597), .Z(n15609) );
  XNOR U16582 ( .A(n15608), .B(n15609), .Z(n15610) );
  XNOR U16583 ( .A(n15611), .B(n15610), .Z(n15604) );
  XOR U16584 ( .A(n15605), .B(n15604), .Z(n15606) );
  XNOR U16585 ( .A(n15607), .B(n15606), .Z(n15744) );
  XNOR U16586 ( .A(n15744), .B(sreg[339]), .Z(n15746) );
  NAND U16587 ( .A(n15599), .B(sreg[338]), .Z(n15603) );
  OR U16588 ( .A(n15601), .B(n15600), .Z(n15602) );
  AND U16589 ( .A(n15603), .B(n15602), .Z(n15745) );
  XOR U16590 ( .A(n15746), .B(n15745), .Z(c[339]) );
  NANDN U16591 ( .A(n15609), .B(n15608), .Z(n15613) );
  NANDN U16592 ( .A(n15611), .B(n15610), .Z(n15612) );
  NAND U16593 ( .A(n15613), .B(n15612), .Z(n15750) );
  OR U16594 ( .A(n15615), .B(n15614), .Z(n15619) );
  NANDN U16595 ( .A(n15617), .B(n15616), .Z(n15618) );
  NAND U16596 ( .A(n15619), .B(n15618), .Z(n15882) );
  OR U16597 ( .A(n15621), .B(n15620), .Z(n15625) );
  NAND U16598 ( .A(n15623), .B(n15622), .Z(n15624) );
  NAND U16599 ( .A(n15625), .B(n15624), .Z(n15821) );
  OR U16600 ( .A(n15627), .B(n15626), .Z(n15631) );
  NANDN U16601 ( .A(n15629), .B(n15628), .Z(n15630) );
  NAND U16602 ( .A(n15631), .B(n15630), .Z(n15820) );
  OR U16603 ( .A(n15633), .B(n15632), .Z(n15637) );
  NANDN U16604 ( .A(n15635), .B(n15634), .Z(n15636) );
  NAND U16605 ( .A(n15637), .B(n15636), .Z(n15819) );
  XOR U16606 ( .A(n15821), .B(n15822), .Z(n15880) );
  OR U16607 ( .A(n15639), .B(n15638), .Z(n15643) );
  NANDN U16608 ( .A(n15641), .B(n15640), .Z(n15642) );
  NAND U16609 ( .A(n15643), .B(n15642), .Z(n15833) );
  XNOR U16610 ( .A(b[19]), .B(a[98]), .Z(n15777) );
  NANDN U16611 ( .A(n15777), .B(n37934), .Z(n15646) );
  NANDN U16612 ( .A(n15644), .B(n37935), .Z(n15645) );
  NAND U16613 ( .A(n15646), .B(n15645), .Z(n15846) );
  XOR U16614 ( .A(b[27]), .B(a[90]), .Z(n15780) );
  NAND U16615 ( .A(n38423), .B(n15780), .Z(n15649) );
  NAND U16616 ( .A(n15647), .B(n38424), .Z(n15648) );
  NAND U16617 ( .A(n15649), .B(n15648), .Z(n15843) );
  XNOR U16618 ( .A(b[5]), .B(a[112]), .Z(n15783) );
  NANDN U16619 ( .A(n15783), .B(n36587), .Z(n15652) );
  NANDN U16620 ( .A(n15650), .B(n36588), .Z(n15651) );
  AND U16621 ( .A(n15652), .B(n15651), .Z(n15844) );
  XNOR U16622 ( .A(n15843), .B(n15844), .Z(n15845) );
  XNOR U16623 ( .A(n15846), .B(n15845), .Z(n15832) );
  NANDN U16624 ( .A(n15653), .B(n37762), .Z(n15655) );
  XOR U16625 ( .A(b[17]), .B(a[100]), .Z(n15786) );
  NAND U16626 ( .A(n15786), .B(n37764), .Z(n15654) );
  NAND U16627 ( .A(n15655), .B(n15654), .Z(n15804) );
  XNOR U16628 ( .A(b[31]), .B(a[86]), .Z(n15789) );
  NANDN U16629 ( .A(n15789), .B(n38552), .Z(n15658) );
  NANDN U16630 ( .A(n15656), .B(n38553), .Z(n15657) );
  NAND U16631 ( .A(n15658), .B(n15657), .Z(n15801) );
  OR U16632 ( .A(n15659), .B(n36105), .Z(n15661) );
  XNOR U16633 ( .A(b[3]), .B(a[114]), .Z(n15792) );
  NANDN U16634 ( .A(n15792), .B(n36107), .Z(n15660) );
  AND U16635 ( .A(n15661), .B(n15660), .Z(n15802) );
  XNOR U16636 ( .A(n15801), .B(n15802), .Z(n15803) );
  XOR U16637 ( .A(n15804), .B(n15803), .Z(n15831) );
  XOR U16638 ( .A(n15832), .B(n15831), .Z(n15834) );
  XOR U16639 ( .A(n15833), .B(n15834), .Z(n15879) );
  XOR U16640 ( .A(n15880), .B(n15879), .Z(n15881) );
  XNOR U16641 ( .A(n15882), .B(n15881), .Z(n15768) );
  OR U16642 ( .A(n15663), .B(n15662), .Z(n15667) );
  NANDN U16643 ( .A(n15665), .B(n15664), .Z(n15666) );
  NAND U16644 ( .A(n15667), .B(n15666), .Z(n15766) );
  NANDN U16645 ( .A(n15669), .B(n15668), .Z(n15673) );
  NANDN U16646 ( .A(n15671), .B(n15670), .Z(n15672) );
  NAND U16647 ( .A(n15673), .B(n15672), .Z(n15887) );
  OR U16648 ( .A(n15675), .B(n15674), .Z(n15679) );
  NANDN U16649 ( .A(n15677), .B(n15676), .Z(n15678) );
  NAND U16650 ( .A(n15679), .B(n15678), .Z(n15886) );
  NANDN U16651 ( .A(n15681), .B(n15680), .Z(n15685) );
  NAND U16652 ( .A(n15683), .B(n15682), .Z(n15684) );
  NAND U16653 ( .A(n15685), .B(n15684), .Z(n15825) );
  NANDN U16654 ( .A(n15687), .B(n15686), .Z(n15691) );
  NAND U16655 ( .A(n15689), .B(n15688), .Z(n15690) );
  AND U16656 ( .A(n15691), .B(n15690), .Z(n15826) );
  XNOR U16657 ( .A(n15825), .B(n15826), .Z(n15827) );
  XNOR U16658 ( .A(b[9]), .B(a[108]), .Z(n15849) );
  NANDN U16659 ( .A(n15849), .B(n36925), .Z(n15694) );
  NANDN U16660 ( .A(n15692), .B(n36926), .Z(n15693) );
  NAND U16661 ( .A(n15694), .B(n15693), .Z(n15809) );
  XNOR U16662 ( .A(b[15]), .B(a[102]), .Z(n15852) );
  OR U16663 ( .A(n15852), .B(n37665), .Z(n15697) );
  NANDN U16664 ( .A(n15695), .B(n37604), .Z(n15696) );
  AND U16665 ( .A(n15697), .B(n15696), .Z(n15807) );
  XNOR U16666 ( .A(b[21]), .B(a[96]), .Z(n15855) );
  NANDN U16667 ( .A(n15855), .B(n38101), .Z(n15700) );
  NANDN U16668 ( .A(n15698), .B(n38102), .Z(n15699) );
  AND U16669 ( .A(n15700), .B(n15699), .Z(n15808) );
  XOR U16670 ( .A(n15809), .B(n15810), .Z(n15798) );
  XNOR U16671 ( .A(b[11]), .B(a[106]), .Z(n15858) );
  OR U16672 ( .A(n15858), .B(n37311), .Z(n15703) );
  NANDN U16673 ( .A(n15701), .B(n37218), .Z(n15702) );
  NAND U16674 ( .A(n15703), .B(n15702), .Z(n15796) );
  XOR U16675 ( .A(n1053), .B(a[104]), .Z(n15861) );
  NANDN U16676 ( .A(n15861), .B(n37424), .Z(n15706) );
  NANDN U16677 ( .A(n15704), .B(n37425), .Z(n15705) );
  AND U16678 ( .A(n15706), .B(n15705), .Z(n15795) );
  XNOR U16679 ( .A(n15796), .B(n15795), .Z(n15797) );
  XOR U16680 ( .A(n15798), .B(n15797), .Z(n15815) );
  NANDN U16681 ( .A(n1049), .B(a[116]), .Z(n15707) );
  XNOR U16682 ( .A(b[1]), .B(n15707), .Z(n15709) );
  NANDN U16683 ( .A(b[0]), .B(a[115]), .Z(n15708) );
  AND U16684 ( .A(n15709), .B(n15708), .Z(n15773) );
  NAND U16685 ( .A(n15710), .B(n38490), .Z(n15712) );
  XNOR U16686 ( .A(n1058), .B(a[88]), .Z(n15864) );
  NANDN U16687 ( .A(n1048), .B(n15864), .Z(n15711) );
  NAND U16688 ( .A(n15712), .B(n15711), .Z(n15771) );
  NANDN U16689 ( .A(n1059), .B(a[84]), .Z(n15772) );
  XNOR U16690 ( .A(n15771), .B(n15772), .Z(n15774) );
  XOR U16691 ( .A(n15773), .B(n15774), .Z(n15813) );
  NANDN U16692 ( .A(n15713), .B(n38205), .Z(n15715) );
  XNOR U16693 ( .A(b[23]), .B(a[94]), .Z(n15870) );
  OR U16694 ( .A(n15870), .B(n38268), .Z(n15714) );
  NAND U16695 ( .A(n15715), .B(n15714), .Z(n15840) );
  XOR U16696 ( .A(b[7]), .B(a[110]), .Z(n15873) );
  NAND U16697 ( .A(n15873), .B(n36701), .Z(n15718) );
  NAND U16698 ( .A(n15716), .B(n36702), .Z(n15717) );
  NAND U16699 ( .A(n15718), .B(n15717), .Z(n15837) );
  XOR U16700 ( .A(b[25]), .B(a[92]), .Z(n15876) );
  NAND U16701 ( .A(n15876), .B(n38325), .Z(n15721) );
  NAND U16702 ( .A(n15719), .B(n38326), .Z(n15720) );
  AND U16703 ( .A(n15721), .B(n15720), .Z(n15838) );
  XNOR U16704 ( .A(n15837), .B(n15838), .Z(n15839) );
  XNOR U16705 ( .A(n15840), .B(n15839), .Z(n15814) );
  XOR U16706 ( .A(n15813), .B(n15814), .Z(n15816) );
  XNOR U16707 ( .A(n15815), .B(n15816), .Z(n15828) );
  XNOR U16708 ( .A(n15827), .B(n15828), .Z(n15885) );
  XNOR U16709 ( .A(n15886), .B(n15885), .Z(n15888) );
  XNOR U16710 ( .A(n15887), .B(n15888), .Z(n15765) );
  XNOR U16711 ( .A(n15766), .B(n15765), .Z(n15767) );
  XOR U16712 ( .A(n15768), .B(n15767), .Z(n15762) );
  NAND U16713 ( .A(n15727), .B(n15726), .Z(n15731) );
  NANDN U16714 ( .A(n15729), .B(n15728), .Z(n15730) );
  AND U16715 ( .A(n15731), .B(n15730), .Z(n15759) );
  XNOR U16716 ( .A(n15760), .B(n15759), .Z(n15761) );
  XNOR U16717 ( .A(n15762), .B(n15761), .Z(n15756) );
  NANDN U16718 ( .A(n15733), .B(n15732), .Z(n15737) );
  NAND U16719 ( .A(n15735), .B(n15734), .Z(n15736) );
  NAND U16720 ( .A(n15737), .B(n15736), .Z(n15753) );
  NANDN U16721 ( .A(n15739), .B(n15738), .Z(n15743) );
  NANDN U16722 ( .A(n15741), .B(n15740), .Z(n15742) );
  NAND U16723 ( .A(n15743), .B(n15742), .Z(n15754) );
  XNOR U16724 ( .A(n15753), .B(n15754), .Z(n15755) );
  XNOR U16725 ( .A(n15756), .B(n15755), .Z(n15749) );
  XOR U16726 ( .A(n15750), .B(n15749), .Z(n15751) );
  XNOR U16727 ( .A(n15752), .B(n15751), .Z(n15891) );
  XNOR U16728 ( .A(n15891), .B(sreg[340]), .Z(n15893) );
  NAND U16729 ( .A(n15744), .B(sreg[339]), .Z(n15748) );
  OR U16730 ( .A(n15746), .B(n15745), .Z(n15747) );
  AND U16731 ( .A(n15748), .B(n15747), .Z(n15892) );
  XOR U16732 ( .A(n15893), .B(n15892), .Z(c[340]) );
  NANDN U16733 ( .A(n15754), .B(n15753), .Z(n15758) );
  NANDN U16734 ( .A(n15756), .B(n15755), .Z(n15757) );
  NAND U16735 ( .A(n15758), .B(n15757), .Z(n15897) );
  NANDN U16736 ( .A(n15760), .B(n15759), .Z(n15764) );
  NAND U16737 ( .A(n15762), .B(n15761), .Z(n15763) );
  NAND U16738 ( .A(n15764), .B(n15763), .Z(n15902) );
  NANDN U16739 ( .A(n15766), .B(n15765), .Z(n15770) );
  NANDN U16740 ( .A(n15768), .B(n15767), .Z(n15769) );
  NAND U16741 ( .A(n15770), .B(n15769), .Z(n15903) );
  XNOR U16742 ( .A(n15902), .B(n15903), .Z(n15904) );
  NANDN U16743 ( .A(n15772), .B(n15771), .Z(n15776) );
  NAND U16744 ( .A(n15774), .B(n15773), .Z(n15775) );
  NAND U16745 ( .A(n15776), .B(n15775), .Z(n15983) );
  XOR U16746 ( .A(b[19]), .B(n17884), .Z(n15950) );
  NANDN U16747 ( .A(n15950), .B(n37934), .Z(n15779) );
  NANDN U16748 ( .A(n15777), .B(n37935), .Z(n15778) );
  NAND U16749 ( .A(n15779), .B(n15778), .Z(n16019) );
  XOR U16750 ( .A(b[27]), .B(a[91]), .Z(n15953) );
  NAND U16751 ( .A(n38423), .B(n15953), .Z(n15782) );
  NAND U16752 ( .A(n15780), .B(n38424), .Z(n15781) );
  NAND U16753 ( .A(n15782), .B(n15781), .Z(n16016) );
  XOR U16754 ( .A(b[5]), .B(n19909), .Z(n15956) );
  NANDN U16755 ( .A(n15956), .B(n36587), .Z(n15785) );
  NANDN U16756 ( .A(n15783), .B(n36588), .Z(n15784) );
  AND U16757 ( .A(n15785), .B(n15784), .Z(n16017) );
  XNOR U16758 ( .A(n16016), .B(n16017), .Z(n16018) );
  XNOR U16759 ( .A(n16019), .B(n16018), .Z(n15980) );
  NAND U16760 ( .A(n15786), .B(n37762), .Z(n15788) );
  XNOR U16761 ( .A(b[17]), .B(a[101]), .Z(n15959) );
  NANDN U16762 ( .A(n15959), .B(n37764), .Z(n15787) );
  NAND U16763 ( .A(n15788), .B(n15787), .Z(n15934) );
  XNOR U16764 ( .A(b[31]), .B(a[87]), .Z(n15962) );
  NANDN U16765 ( .A(n15962), .B(n38552), .Z(n15791) );
  NANDN U16766 ( .A(n15789), .B(n38553), .Z(n15790) );
  AND U16767 ( .A(n15791), .B(n15790), .Z(n15932) );
  OR U16768 ( .A(n15792), .B(n36105), .Z(n15794) );
  XNOR U16769 ( .A(b[3]), .B(a[115]), .Z(n15965) );
  NANDN U16770 ( .A(n15965), .B(n36107), .Z(n15793) );
  AND U16771 ( .A(n15794), .B(n15793), .Z(n15933) );
  XOR U16772 ( .A(n15934), .B(n15935), .Z(n15981) );
  XOR U16773 ( .A(n15980), .B(n15981), .Z(n15982) );
  XNOR U16774 ( .A(n15983), .B(n15982), .Z(n16028) );
  NANDN U16775 ( .A(n15796), .B(n15795), .Z(n15800) );
  NAND U16776 ( .A(n15798), .B(n15797), .Z(n15799) );
  NAND U16777 ( .A(n15800), .B(n15799), .Z(n15971) );
  NANDN U16778 ( .A(n15802), .B(n15801), .Z(n15806) );
  NAND U16779 ( .A(n15804), .B(n15803), .Z(n15805) );
  NAND U16780 ( .A(n15806), .B(n15805), .Z(n15969) );
  OR U16781 ( .A(n15808), .B(n15807), .Z(n15812) );
  NANDN U16782 ( .A(n15810), .B(n15809), .Z(n15811) );
  NAND U16783 ( .A(n15812), .B(n15811), .Z(n15968) );
  XNOR U16784 ( .A(n15971), .B(n15970), .Z(n16029) );
  XOR U16785 ( .A(n16028), .B(n16029), .Z(n16031) );
  NANDN U16786 ( .A(n15814), .B(n15813), .Z(n15818) );
  OR U16787 ( .A(n15816), .B(n15815), .Z(n15817) );
  NAND U16788 ( .A(n15818), .B(n15817), .Z(n16030) );
  XOR U16789 ( .A(n16031), .B(n16030), .Z(n15916) );
  OR U16790 ( .A(n15820), .B(n15819), .Z(n15824) );
  NANDN U16791 ( .A(n15822), .B(n15821), .Z(n15823) );
  NAND U16792 ( .A(n15824), .B(n15823), .Z(n15915) );
  NANDN U16793 ( .A(n15826), .B(n15825), .Z(n15830) );
  NANDN U16794 ( .A(n15828), .B(n15827), .Z(n15829) );
  NAND U16795 ( .A(n15830), .B(n15829), .Z(n16036) );
  NANDN U16796 ( .A(n15832), .B(n15831), .Z(n15836) );
  OR U16797 ( .A(n15834), .B(n15833), .Z(n15835) );
  NAND U16798 ( .A(n15836), .B(n15835), .Z(n16035) );
  NANDN U16799 ( .A(n15838), .B(n15837), .Z(n15842) );
  NAND U16800 ( .A(n15840), .B(n15839), .Z(n15841) );
  NAND U16801 ( .A(n15842), .B(n15841), .Z(n15974) );
  NANDN U16802 ( .A(n15844), .B(n15843), .Z(n15848) );
  NAND U16803 ( .A(n15846), .B(n15845), .Z(n15847) );
  AND U16804 ( .A(n15848), .B(n15847), .Z(n15975) );
  XNOR U16805 ( .A(n15974), .B(n15975), .Z(n15976) );
  XNOR U16806 ( .A(n1052), .B(a[109]), .Z(n15986) );
  NAND U16807 ( .A(n36925), .B(n15986), .Z(n15851) );
  NANDN U16808 ( .A(n15849), .B(n36926), .Z(n15850) );
  NAND U16809 ( .A(n15851), .B(n15850), .Z(n15940) );
  XNOR U16810 ( .A(b[15]), .B(a[103]), .Z(n15989) );
  OR U16811 ( .A(n15989), .B(n37665), .Z(n15854) );
  NANDN U16812 ( .A(n15852), .B(n37604), .Z(n15853) );
  AND U16813 ( .A(n15854), .B(n15853), .Z(n15938) );
  XNOR U16814 ( .A(n1056), .B(a[97]), .Z(n15992) );
  NAND U16815 ( .A(n15992), .B(n38101), .Z(n15857) );
  NANDN U16816 ( .A(n15855), .B(n38102), .Z(n15856) );
  AND U16817 ( .A(n15857), .B(n15856), .Z(n15939) );
  XOR U16818 ( .A(n15940), .B(n15941), .Z(n15929) );
  XOR U16819 ( .A(b[11]), .B(n18980), .Z(n15995) );
  OR U16820 ( .A(n15995), .B(n37311), .Z(n15860) );
  NANDN U16821 ( .A(n15858), .B(n37218), .Z(n15859) );
  NAND U16822 ( .A(n15860), .B(n15859), .Z(n15927) );
  XOR U16823 ( .A(n1053), .B(a[105]), .Z(n15998) );
  NANDN U16824 ( .A(n15998), .B(n37424), .Z(n15863) );
  NANDN U16825 ( .A(n15861), .B(n37425), .Z(n15862) );
  NAND U16826 ( .A(n15863), .B(n15862), .Z(n15926) );
  XOR U16827 ( .A(n15929), .B(n15928), .Z(n15923) );
  NAND U16828 ( .A(n38490), .B(n15864), .Z(n15866) );
  XNOR U16829 ( .A(n1058), .B(a[89]), .Z(n16004) );
  NANDN U16830 ( .A(n1048), .B(n16004), .Z(n15865) );
  NAND U16831 ( .A(n15866), .B(n15865), .Z(n15944) );
  NANDN U16832 ( .A(n1059), .B(a[85]), .Z(n15945) );
  XNOR U16833 ( .A(n15944), .B(n15945), .Z(n15947) );
  NANDN U16834 ( .A(n1049), .B(a[117]), .Z(n15867) );
  XNOR U16835 ( .A(b[1]), .B(n15867), .Z(n15869) );
  NANDN U16836 ( .A(b[0]), .B(a[116]), .Z(n15868) );
  AND U16837 ( .A(n15869), .B(n15868), .Z(n15946) );
  XNOR U16838 ( .A(n15947), .B(n15946), .Z(n15921) );
  NANDN U16839 ( .A(n15870), .B(n38205), .Z(n15872) );
  XNOR U16840 ( .A(b[23]), .B(a[95]), .Z(n16007) );
  OR U16841 ( .A(n16007), .B(n38268), .Z(n15871) );
  NAND U16842 ( .A(n15872), .B(n15871), .Z(n16025) );
  XOR U16843 ( .A(b[7]), .B(a[111]), .Z(n16010) );
  NAND U16844 ( .A(n16010), .B(n36701), .Z(n15875) );
  NAND U16845 ( .A(n15873), .B(n36702), .Z(n15874) );
  NAND U16846 ( .A(n15875), .B(n15874), .Z(n16022) );
  XNOR U16847 ( .A(b[25]), .B(a[93]), .Z(n16013) );
  NANDN U16848 ( .A(n16013), .B(n38325), .Z(n15878) );
  NAND U16849 ( .A(n15876), .B(n38326), .Z(n15877) );
  AND U16850 ( .A(n15878), .B(n15877), .Z(n16023) );
  XNOR U16851 ( .A(n16022), .B(n16023), .Z(n16024) );
  XOR U16852 ( .A(n16025), .B(n16024), .Z(n15920) );
  XOR U16853 ( .A(n15923), .B(n15922), .Z(n15977) );
  XNOR U16854 ( .A(n15976), .B(n15977), .Z(n16034) );
  XNOR U16855 ( .A(n16035), .B(n16034), .Z(n16037) );
  XNOR U16856 ( .A(n16036), .B(n16037), .Z(n15914) );
  XOR U16857 ( .A(n15915), .B(n15914), .Z(n15917) );
  NAND U16858 ( .A(n15880), .B(n15879), .Z(n15884) );
  NAND U16859 ( .A(n15882), .B(n15881), .Z(n15883) );
  NAND U16860 ( .A(n15884), .B(n15883), .Z(n15909) );
  NAND U16861 ( .A(n15886), .B(n15885), .Z(n15890) );
  NANDN U16862 ( .A(n15888), .B(n15887), .Z(n15889) );
  AND U16863 ( .A(n15890), .B(n15889), .Z(n15908) );
  XNOR U16864 ( .A(n15909), .B(n15908), .Z(n15910) );
  XOR U16865 ( .A(n15911), .B(n15910), .Z(n15905) );
  XOR U16866 ( .A(n15904), .B(n15905), .Z(n15896) );
  XOR U16867 ( .A(n15897), .B(n15896), .Z(n15898) );
  XNOR U16868 ( .A(n15899), .B(n15898), .Z(n16040) );
  XNOR U16869 ( .A(n16040), .B(sreg[341]), .Z(n16042) );
  NAND U16870 ( .A(n15891), .B(sreg[340]), .Z(n15895) );
  OR U16871 ( .A(n15893), .B(n15892), .Z(n15894) );
  AND U16872 ( .A(n15895), .B(n15894), .Z(n16041) );
  XOR U16873 ( .A(n16042), .B(n16041), .Z(c[341]) );
  NAND U16874 ( .A(n15897), .B(n15896), .Z(n15901) );
  NAND U16875 ( .A(n15899), .B(n15898), .Z(n15900) );
  NAND U16876 ( .A(n15901), .B(n15900), .Z(n16048) );
  NANDN U16877 ( .A(n15903), .B(n15902), .Z(n15907) );
  NAND U16878 ( .A(n15905), .B(n15904), .Z(n15906) );
  NAND U16879 ( .A(n15907), .B(n15906), .Z(n16046) );
  NANDN U16880 ( .A(n15909), .B(n15908), .Z(n15913) );
  NAND U16881 ( .A(n15911), .B(n15910), .Z(n15912) );
  NAND U16882 ( .A(n15913), .B(n15912), .Z(n16051) );
  NANDN U16883 ( .A(n15915), .B(n15914), .Z(n15919) );
  OR U16884 ( .A(n15917), .B(n15916), .Z(n15918) );
  NAND U16885 ( .A(n15919), .B(n15918), .Z(n16052) );
  XNOR U16886 ( .A(n16051), .B(n16052), .Z(n16053) );
  NANDN U16887 ( .A(n15921), .B(n15920), .Z(n15925) );
  NANDN U16888 ( .A(n15923), .B(n15922), .Z(n15924) );
  NAND U16889 ( .A(n15925), .B(n15924), .Z(n16166) );
  OR U16890 ( .A(n15927), .B(n15926), .Z(n15931) );
  NAND U16891 ( .A(n15929), .B(n15928), .Z(n15930) );
  NAND U16892 ( .A(n15931), .B(n15930), .Z(n16105) );
  OR U16893 ( .A(n15933), .B(n15932), .Z(n15937) );
  NANDN U16894 ( .A(n15935), .B(n15934), .Z(n15936) );
  NAND U16895 ( .A(n15937), .B(n15936), .Z(n16104) );
  OR U16896 ( .A(n15939), .B(n15938), .Z(n15943) );
  NANDN U16897 ( .A(n15941), .B(n15940), .Z(n15942) );
  NAND U16898 ( .A(n15943), .B(n15942), .Z(n16103) );
  XOR U16899 ( .A(n16105), .B(n16106), .Z(n16163) );
  NANDN U16900 ( .A(n15945), .B(n15944), .Z(n15949) );
  NAND U16901 ( .A(n15947), .B(n15946), .Z(n15948) );
  NAND U16902 ( .A(n15949), .B(n15948), .Z(n16118) );
  XNOR U16903 ( .A(b[19]), .B(a[100]), .Z(n16063) );
  NANDN U16904 ( .A(n16063), .B(n37934), .Z(n15952) );
  NANDN U16905 ( .A(n15950), .B(n37935), .Z(n15951) );
  NAND U16906 ( .A(n15952), .B(n15951), .Z(n16130) );
  XOR U16907 ( .A(b[27]), .B(a[92]), .Z(n16066) );
  NAND U16908 ( .A(n38423), .B(n16066), .Z(n15955) );
  NAND U16909 ( .A(n15953), .B(n38424), .Z(n15954) );
  NAND U16910 ( .A(n15955), .B(n15954), .Z(n16127) );
  XNOR U16911 ( .A(b[5]), .B(a[114]), .Z(n16069) );
  NANDN U16912 ( .A(n16069), .B(n36587), .Z(n15958) );
  NANDN U16913 ( .A(n15956), .B(n36588), .Z(n15957) );
  AND U16914 ( .A(n15958), .B(n15957), .Z(n16128) );
  XNOR U16915 ( .A(n16127), .B(n16128), .Z(n16129) );
  XNOR U16916 ( .A(n16130), .B(n16129), .Z(n16116) );
  NANDN U16917 ( .A(n15959), .B(n37762), .Z(n15961) );
  XOR U16918 ( .A(b[17]), .B(a[102]), .Z(n16072) );
  NAND U16919 ( .A(n16072), .B(n37764), .Z(n15960) );
  NAND U16920 ( .A(n15961), .B(n15960), .Z(n16090) );
  XNOR U16921 ( .A(b[31]), .B(a[88]), .Z(n16075) );
  NANDN U16922 ( .A(n16075), .B(n38552), .Z(n15964) );
  NANDN U16923 ( .A(n15962), .B(n38553), .Z(n15963) );
  NAND U16924 ( .A(n15964), .B(n15963), .Z(n16087) );
  OR U16925 ( .A(n15965), .B(n36105), .Z(n15967) );
  XNOR U16926 ( .A(b[3]), .B(a[116]), .Z(n16078) );
  NANDN U16927 ( .A(n16078), .B(n36107), .Z(n15966) );
  AND U16928 ( .A(n15967), .B(n15966), .Z(n16088) );
  XNOR U16929 ( .A(n16087), .B(n16088), .Z(n16089) );
  XOR U16930 ( .A(n16090), .B(n16089), .Z(n16115) );
  XNOR U16931 ( .A(n16116), .B(n16115), .Z(n16117) );
  XNOR U16932 ( .A(n16118), .B(n16117), .Z(n16164) );
  XNOR U16933 ( .A(n16163), .B(n16164), .Z(n16165) );
  XNOR U16934 ( .A(n16166), .B(n16165), .Z(n16184) );
  OR U16935 ( .A(n15969), .B(n15968), .Z(n15973) );
  NAND U16936 ( .A(n15971), .B(n15970), .Z(n15972) );
  NAND U16937 ( .A(n15973), .B(n15972), .Z(n16182) );
  NANDN U16938 ( .A(n15975), .B(n15974), .Z(n15979) );
  NANDN U16939 ( .A(n15977), .B(n15976), .Z(n15978) );
  NAND U16940 ( .A(n15979), .B(n15978), .Z(n16172) );
  OR U16941 ( .A(n15981), .B(n15980), .Z(n15985) );
  NAND U16942 ( .A(n15983), .B(n15982), .Z(n15984) );
  NAND U16943 ( .A(n15985), .B(n15984), .Z(n16169) );
  XNOR U16944 ( .A(b[9]), .B(a[110]), .Z(n16133) );
  NANDN U16945 ( .A(n16133), .B(n36925), .Z(n15988) );
  NAND U16946 ( .A(n36926), .B(n15986), .Z(n15987) );
  NAND U16947 ( .A(n15988), .B(n15987), .Z(n16095) );
  XNOR U16948 ( .A(n1054), .B(a[104]), .Z(n16136) );
  NANDN U16949 ( .A(n37665), .B(n16136), .Z(n15991) );
  NANDN U16950 ( .A(n15989), .B(n37604), .Z(n15990) );
  NAND U16951 ( .A(n15991), .B(n15990), .Z(n16093) );
  XNOR U16952 ( .A(b[21]), .B(a[98]), .Z(n16139) );
  NANDN U16953 ( .A(n16139), .B(n38101), .Z(n15994) );
  NAND U16954 ( .A(n38102), .B(n15992), .Z(n15993) );
  NAND U16955 ( .A(n15994), .B(n15993), .Z(n16094) );
  XNOR U16956 ( .A(n16093), .B(n16094), .Z(n16096) );
  XOR U16957 ( .A(n16095), .B(n16096), .Z(n16084) );
  XNOR U16958 ( .A(b[11]), .B(a[108]), .Z(n16142) );
  OR U16959 ( .A(n16142), .B(n37311), .Z(n15997) );
  NANDN U16960 ( .A(n15995), .B(n37218), .Z(n15996) );
  NAND U16961 ( .A(n15997), .B(n15996), .Z(n16082) );
  XOR U16962 ( .A(n1053), .B(a[106]), .Z(n16145) );
  NANDN U16963 ( .A(n16145), .B(n37424), .Z(n16000) );
  NANDN U16964 ( .A(n15998), .B(n37425), .Z(n15999) );
  AND U16965 ( .A(n16000), .B(n15999), .Z(n16081) );
  XNOR U16966 ( .A(n16082), .B(n16081), .Z(n16083) );
  XNOR U16967 ( .A(n16084), .B(n16083), .Z(n16100) );
  ANDN U16968 ( .B(a[118]), .A(n1049), .Z(n16001) );
  XOR U16969 ( .A(b[1]), .B(n16001), .Z(n16003) );
  NANDN U16970 ( .A(b[0]), .B(a[117]), .Z(n16002) );
  NAND U16971 ( .A(n16003), .B(n16002), .Z(n16060) );
  NAND U16972 ( .A(n38490), .B(n16004), .Z(n16006) );
  XNOR U16973 ( .A(n1058), .B(a[90]), .Z(n16151) );
  NANDN U16974 ( .A(n1048), .B(n16151), .Z(n16005) );
  NAND U16975 ( .A(n16006), .B(n16005), .Z(n16057) );
  NANDN U16976 ( .A(n1059), .B(a[86]), .Z(n16058) );
  XNOR U16977 ( .A(n16057), .B(n16058), .Z(n16059) );
  XOR U16978 ( .A(n16060), .B(n16059), .Z(n16098) );
  NANDN U16979 ( .A(n16007), .B(n38205), .Z(n16009) );
  XNOR U16980 ( .A(b[23]), .B(a[96]), .Z(n16154) );
  OR U16981 ( .A(n16154), .B(n38268), .Z(n16008) );
  NAND U16982 ( .A(n16009), .B(n16008), .Z(n16124) );
  XOR U16983 ( .A(b[7]), .B(a[112]), .Z(n16157) );
  NAND U16984 ( .A(n16157), .B(n36701), .Z(n16012) );
  NAND U16985 ( .A(n16010), .B(n36702), .Z(n16011) );
  NAND U16986 ( .A(n16012), .B(n16011), .Z(n16121) );
  XOR U16987 ( .A(b[25]), .B(a[94]), .Z(n16160) );
  NAND U16988 ( .A(n16160), .B(n38325), .Z(n16015) );
  NANDN U16989 ( .A(n16013), .B(n38326), .Z(n16014) );
  AND U16990 ( .A(n16015), .B(n16014), .Z(n16122) );
  XNOR U16991 ( .A(n16121), .B(n16122), .Z(n16123) );
  XOR U16992 ( .A(n16124), .B(n16123), .Z(n16097) );
  XNOR U16993 ( .A(n16098), .B(n16097), .Z(n16099) );
  XOR U16994 ( .A(n16100), .B(n16099), .Z(n16112) );
  NANDN U16995 ( .A(n16017), .B(n16016), .Z(n16021) );
  NAND U16996 ( .A(n16019), .B(n16018), .Z(n16020) );
  NAND U16997 ( .A(n16021), .B(n16020), .Z(n16110) );
  NANDN U16998 ( .A(n16023), .B(n16022), .Z(n16027) );
  NAND U16999 ( .A(n16025), .B(n16024), .Z(n16026) );
  AND U17000 ( .A(n16027), .B(n16026), .Z(n16109) );
  XNOR U17001 ( .A(n16110), .B(n16109), .Z(n16111) );
  XNOR U17002 ( .A(n16112), .B(n16111), .Z(n16170) );
  XNOR U17003 ( .A(n16169), .B(n16170), .Z(n16171) );
  XOR U17004 ( .A(n16172), .B(n16171), .Z(n16181) );
  XNOR U17005 ( .A(n16182), .B(n16181), .Z(n16183) );
  XOR U17006 ( .A(n16184), .B(n16183), .Z(n16178) );
  NANDN U17007 ( .A(n16029), .B(n16028), .Z(n16033) );
  OR U17008 ( .A(n16031), .B(n16030), .Z(n16032) );
  NAND U17009 ( .A(n16033), .B(n16032), .Z(n16175) );
  NAND U17010 ( .A(n16035), .B(n16034), .Z(n16039) );
  NANDN U17011 ( .A(n16037), .B(n16036), .Z(n16038) );
  NAND U17012 ( .A(n16039), .B(n16038), .Z(n16176) );
  XNOR U17013 ( .A(n16175), .B(n16176), .Z(n16177) );
  XOR U17014 ( .A(n16178), .B(n16177), .Z(n16054) );
  XOR U17015 ( .A(n16053), .B(n16054), .Z(n16045) );
  XOR U17016 ( .A(n16046), .B(n16045), .Z(n16047) );
  XNOR U17017 ( .A(n16048), .B(n16047), .Z(n16187) );
  XNOR U17018 ( .A(n16187), .B(sreg[342]), .Z(n16189) );
  NAND U17019 ( .A(n16040), .B(sreg[341]), .Z(n16044) );
  OR U17020 ( .A(n16042), .B(n16041), .Z(n16043) );
  AND U17021 ( .A(n16044), .B(n16043), .Z(n16188) );
  XOR U17022 ( .A(n16189), .B(n16188), .Z(c[342]) );
  NAND U17023 ( .A(n16046), .B(n16045), .Z(n16050) );
  NAND U17024 ( .A(n16048), .B(n16047), .Z(n16049) );
  NAND U17025 ( .A(n16050), .B(n16049), .Z(n16195) );
  NANDN U17026 ( .A(n16052), .B(n16051), .Z(n16056) );
  NAND U17027 ( .A(n16054), .B(n16053), .Z(n16055) );
  NAND U17028 ( .A(n16056), .B(n16055), .Z(n16193) );
  NANDN U17029 ( .A(n16058), .B(n16057), .Z(n16062) );
  NANDN U17030 ( .A(n16060), .B(n16059), .Z(n16061) );
  NAND U17031 ( .A(n16062), .B(n16061), .Z(n16275) );
  XOR U17032 ( .A(b[19]), .B(n17812), .Z(n16244) );
  NANDN U17033 ( .A(n16244), .B(n37934), .Z(n16065) );
  NANDN U17034 ( .A(n16063), .B(n37935), .Z(n16064) );
  NAND U17035 ( .A(n16065), .B(n16064), .Z(n16287) );
  XNOR U17036 ( .A(b[27]), .B(a[93]), .Z(n16247) );
  NANDN U17037 ( .A(n16247), .B(n38423), .Z(n16068) );
  NAND U17038 ( .A(n16066), .B(n38424), .Z(n16067) );
  NAND U17039 ( .A(n16068), .B(n16067), .Z(n16284) );
  XNOR U17040 ( .A(b[5]), .B(a[115]), .Z(n16250) );
  NANDN U17041 ( .A(n16250), .B(n36587), .Z(n16071) );
  NANDN U17042 ( .A(n16069), .B(n36588), .Z(n16070) );
  AND U17043 ( .A(n16071), .B(n16070), .Z(n16285) );
  XNOR U17044 ( .A(n16284), .B(n16285), .Z(n16286) );
  XNOR U17045 ( .A(n16287), .B(n16286), .Z(n16272) );
  NAND U17046 ( .A(n16072), .B(n37762), .Z(n16074) );
  XOR U17047 ( .A(b[17]), .B(a[103]), .Z(n16253) );
  NAND U17048 ( .A(n16253), .B(n37764), .Z(n16073) );
  NAND U17049 ( .A(n16074), .B(n16073), .Z(n16228) );
  XNOR U17050 ( .A(b[31]), .B(a[89]), .Z(n16256) );
  NANDN U17051 ( .A(n16256), .B(n38552), .Z(n16077) );
  NANDN U17052 ( .A(n16075), .B(n38553), .Z(n16076) );
  AND U17053 ( .A(n16077), .B(n16076), .Z(n16226) );
  OR U17054 ( .A(n16078), .B(n36105), .Z(n16080) );
  XNOR U17055 ( .A(b[3]), .B(a[117]), .Z(n16259) );
  NANDN U17056 ( .A(n16259), .B(n36107), .Z(n16079) );
  AND U17057 ( .A(n16080), .B(n16079), .Z(n16227) );
  XOR U17058 ( .A(n16228), .B(n16229), .Z(n16273) );
  XOR U17059 ( .A(n16272), .B(n16273), .Z(n16274) );
  XNOR U17060 ( .A(n16275), .B(n16274), .Z(n16211) );
  NANDN U17061 ( .A(n16082), .B(n16081), .Z(n16086) );
  NAND U17062 ( .A(n16084), .B(n16083), .Z(n16085) );
  NAND U17063 ( .A(n16086), .B(n16085), .Z(n16264) );
  NANDN U17064 ( .A(n16088), .B(n16087), .Z(n16092) );
  NAND U17065 ( .A(n16090), .B(n16089), .Z(n16091) );
  NAND U17066 ( .A(n16092), .B(n16091), .Z(n16263) );
  XNOR U17067 ( .A(n16263), .B(n16262), .Z(n16265) );
  XOR U17068 ( .A(n16264), .B(n16265), .Z(n16210) );
  XOR U17069 ( .A(n16211), .B(n16210), .Z(n16212) );
  NANDN U17070 ( .A(n16098), .B(n16097), .Z(n16102) );
  NAND U17071 ( .A(n16100), .B(n16099), .Z(n16101) );
  NAND U17072 ( .A(n16102), .B(n16101), .Z(n16213) );
  XNOR U17073 ( .A(n16212), .B(n16213), .Z(n16328) );
  OR U17074 ( .A(n16104), .B(n16103), .Z(n16108) );
  NANDN U17075 ( .A(n16106), .B(n16105), .Z(n16107) );
  NAND U17076 ( .A(n16108), .B(n16107), .Z(n16327) );
  NANDN U17077 ( .A(n16110), .B(n16109), .Z(n16114) );
  NANDN U17078 ( .A(n16112), .B(n16111), .Z(n16113) );
  NAND U17079 ( .A(n16114), .B(n16113), .Z(n16207) );
  NANDN U17080 ( .A(n16116), .B(n16115), .Z(n16120) );
  NAND U17081 ( .A(n16118), .B(n16117), .Z(n16119) );
  NAND U17082 ( .A(n16120), .B(n16119), .Z(n16205) );
  NANDN U17083 ( .A(n16122), .B(n16121), .Z(n16126) );
  NAND U17084 ( .A(n16124), .B(n16123), .Z(n16125) );
  NAND U17085 ( .A(n16126), .B(n16125), .Z(n16266) );
  NANDN U17086 ( .A(n16128), .B(n16127), .Z(n16132) );
  NAND U17087 ( .A(n16130), .B(n16129), .Z(n16131) );
  AND U17088 ( .A(n16132), .B(n16131), .Z(n16267) );
  XNOR U17089 ( .A(n16266), .B(n16267), .Z(n16268) );
  XNOR U17090 ( .A(b[9]), .B(a[111]), .Z(n16290) );
  NANDN U17091 ( .A(n16290), .B(n36925), .Z(n16135) );
  NANDN U17092 ( .A(n16133), .B(n36926), .Z(n16134) );
  NAND U17093 ( .A(n16135), .B(n16134), .Z(n16234) );
  XNOR U17094 ( .A(b[15]), .B(a[105]), .Z(n16293) );
  OR U17095 ( .A(n16293), .B(n37665), .Z(n16138) );
  NAND U17096 ( .A(n16136), .B(n37604), .Z(n16137) );
  AND U17097 ( .A(n16138), .B(n16137), .Z(n16232) );
  XOR U17098 ( .A(b[21]), .B(n17884), .Z(n16296) );
  NANDN U17099 ( .A(n16296), .B(n38101), .Z(n16141) );
  NANDN U17100 ( .A(n16139), .B(n38102), .Z(n16140) );
  AND U17101 ( .A(n16141), .B(n16140), .Z(n16233) );
  XOR U17102 ( .A(n16234), .B(n16235), .Z(n16223) );
  XNOR U17103 ( .A(b[11]), .B(a[109]), .Z(n16299) );
  OR U17104 ( .A(n16299), .B(n37311), .Z(n16144) );
  NANDN U17105 ( .A(n16142), .B(n37218), .Z(n16143) );
  NAND U17106 ( .A(n16144), .B(n16143), .Z(n16221) );
  XOR U17107 ( .A(n1053), .B(a[107]), .Z(n16302) );
  NANDN U17108 ( .A(n16302), .B(n37424), .Z(n16147) );
  NANDN U17109 ( .A(n16145), .B(n37425), .Z(n16146) );
  NAND U17110 ( .A(n16147), .B(n16146), .Z(n16220) );
  XOR U17111 ( .A(n16223), .B(n16222), .Z(n16217) );
  NANDN U17112 ( .A(n1049), .B(a[119]), .Z(n16148) );
  XNOR U17113 ( .A(b[1]), .B(n16148), .Z(n16150) );
  IV U17114 ( .A(a[118]), .Z(n20271) );
  NANDN U17115 ( .A(n20271), .B(n1049), .Z(n16149) );
  AND U17116 ( .A(n16150), .B(n16149), .Z(n16240) );
  NAND U17117 ( .A(n38490), .B(n16151), .Z(n16153) );
  XNOR U17118 ( .A(n1058), .B(a[91]), .Z(n16308) );
  NANDN U17119 ( .A(n1048), .B(n16308), .Z(n16152) );
  NAND U17120 ( .A(n16153), .B(n16152), .Z(n16238) );
  NANDN U17121 ( .A(n1059), .B(a[87]), .Z(n16239) );
  XNOR U17122 ( .A(n16238), .B(n16239), .Z(n16241) );
  XNOR U17123 ( .A(n16240), .B(n16241), .Z(n16215) );
  NANDN U17124 ( .A(n16154), .B(n38205), .Z(n16156) );
  XNOR U17125 ( .A(b[23]), .B(a[97]), .Z(n16311) );
  OR U17126 ( .A(n16311), .B(n38268), .Z(n16155) );
  NAND U17127 ( .A(n16156), .B(n16155), .Z(n16281) );
  XNOR U17128 ( .A(b[7]), .B(a[113]), .Z(n16314) );
  NANDN U17129 ( .A(n16314), .B(n36701), .Z(n16159) );
  NAND U17130 ( .A(n16157), .B(n36702), .Z(n16158) );
  NAND U17131 ( .A(n16159), .B(n16158), .Z(n16278) );
  XOR U17132 ( .A(b[25]), .B(a[95]), .Z(n16317) );
  NAND U17133 ( .A(n16317), .B(n38325), .Z(n16162) );
  NAND U17134 ( .A(n16160), .B(n38326), .Z(n16161) );
  AND U17135 ( .A(n16162), .B(n16161), .Z(n16279) );
  XNOR U17136 ( .A(n16278), .B(n16279), .Z(n16280) );
  XOR U17137 ( .A(n16281), .B(n16280), .Z(n16214) );
  XOR U17138 ( .A(n16217), .B(n16216), .Z(n16269) );
  XNOR U17139 ( .A(n16268), .B(n16269), .Z(n16204) );
  XOR U17140 ( .A(n16205), .B(n16204), .Z(n16206) );
  XNOR U17141 ( .A(n16207), .B(n16206), .Z(n16326) );
  XOR U17142 ( .A(n16327), .B(n16326), .Z(n16329) );
  NANDN U17143 ( .A(n16164), .B(n16163), .Z(n16168) );
  NAND U17144 ( .A(n16166), .B(n16165), .Z(n16167) );
  NAND U17145 ( .A(n16168), .B(n16167), .Z(n16321) );
  NANDN U17146 ( .A(n16170), .B(n16169), .Z(n16174) );
  NAND U17147 ( .A(n16172), .B(n16171), .Z(n16173) );
  AND U17148 ( .A(n16174), .B(n16173), .Z(n16320) );
  XNOR U17149 ( .A(n16321), .B(n16320), .Z(n16322) );
  XOR U17150 ( .A(n16323), .B(n16322), .Z(n16200) );
  NANDN U17151 ( .A(n16176), .B(n16175), .Z(n16180) );
  NAND U17152 ( .A(n16178), .B(n16177), .Z(n16179) );
  NAND U17153 ( .A(n16180), .B(n16179), .Z(n16198) );
  NANDN U17154 ( .A(n16182), .B(n16181), .Z(n16186) );
  NANDN U17155 ( .A(n16184), .B(n16183), .Z(n16185) );
  NAND U17156 ( .A(n16186), .B(n16185), .Z(n16199) );
  XNOR U17157 ( .A(n16198), .B(n16199), .Z(n16201) );
  XOR U17158 ( .A(n16200), .B(n16201), .Z(n16192) );
  XOR U17159 ( .A(n16193), .B(n16192), .Z(n16194) );
  XNOR U17160 ( .A(n16195), .B(n16194), .Z(n16332) );
  XNOR U17161 ( .A(n16332), .B(sreg[343]), .Z(n16334) );
  NAND U17162 ( .A(n16187), .B(sreg[342]), .Z(n16191) );
  OR U17163 ( .A(n16189), .B(n16188), .Z(n16190) );
  AND U17164 ( .A(n16191), .B(n16190), .Z(n16333) );
  XOR U17165 ( .A(n16334), .B(n16333), .Z(c[343]) );
  NAND U17166 ( .A(n16193), .B(n16192), .Z(n16197) );
  NAND U17167 ( .A(n16195), .B(n16194), .Z(n16196) );
  NAND U17168 ( .A(n16197), .B(n16196), .Z(n16340) );
  NANDN U17169 ( .A(n16199), .B(n16198), .Z(n16203) );
  NAND U17170 ( .A(n16201), .B(n16200), .Z(n16202) );
  NAND U17171 ( .A(n16203), .B(n16202), .Z(n16337) );
  NAND U17172 ( .A(n16205), .B(n16204), .Z(n16209) );
  NANDN U17173 ( .A(n16207), .B(n16206), .Z(n16208) );
  NAND U17174 ( .A(n16209), .B(n16208), .Z(n16349) );
  XNOR U17175 ( .A(n16349), .B(n16350), .Z(n16351) );
  NANDN U17176 ( .A(n16215), .B(n16214), .Z(n16219) );
  NANDN U17177 ( .A(n16217), .B(n16216), .Z(n16218) );
  NAND U17178 ( .A(n16219), .B(n16218), .Z(n16472) );
  OR U17179 ( .A(n16221), .B(n16220), .Z(n16225) );
  NAND U17180 ( .A(n16223), .B(n16222), .Z(n16224) );
  NAND U17181 ( .A(n16225), .B(n16224), .Z(n16411) );
  OR U17182 ( .A(n16227), .B(n16226), .Z(n16231) );
  NANDN U17183 ( .A(n16229), .B(n16228), .Z(n16230) );
  NAND U17184 ( .A(n16231), .B(n16230), .Z(n16410) );
  OR U17185 ( .A(n16233), .B(n16232), .Z(n16237) );
  NANDN U17186 ( .A(n16235), .B(n16234), .Z(n16236) );
  NAND U17187 ( .A(n16237), .B(n16236), .Z(n16409) );
  XOR U17188 ( .A(n16411), .B(n16412), .Z(n16469) );
  NANDN U17189 ( .A(n16239), .B(n16238), .Z(n16243) );
  NAND U17190 ( .A(n16241), .B(n16240), .Z(n16242) );
  NAND U17191 ( .A(n16243), .B(n16242), .Z(n16424) );
  XNOR U17192 ( .A(b[19]), .B(a[102]), .Z(n16367) );
  NANDN U17193 ( .A(n16367), .B(n37934), .Z(n16246) );
  NANDN U17194 ( .A(n16244), .B(n37935), .Z(n16245) );
  NAND U17195 ( .A(n16246), .B(n16245), .Z(n16436) );
  XOR U17196 ( .A(b[27]), .B(a[94]), .Z(n16370) );
  NAND U17197 ( .A(n38423), .B(n16370), .Z(n16249) );
  NANDN U17198 ( .A(n16247), .B(n38424), .Z(n16248) );
  NAND U17199 ( .A(n16249), .B(n16248), .Z(n16433) );
  XNOR U17200 ( .A(b[5]), .B(a[116]), .Z(n16373) );
  NANDN U17201 ( .A(n16373), .B(n36587), .Z(n16252) );
  NANDN U17202 ( .A(n16250), .B(n36588), .Z(n16251) );
  AND U17203 ( .A(n16252), .B(n16251), .Z(n16434) );
  XNOR U17204 ( .A(n16433), .B(n16434), .Z(n16435) );
  XNOR U17205 ( .A(n16436), .B(n16435), .Z(n16422) );
  NAND U17206 ( .A(n16253), .B(n37762), .Z(n16255) );
  XOR U17207 ( .A(b[17]), .B(a[104]), .Z(n16376) );
  NAND U17208 ( .A(n16376), .B(n37764), .Z(n16254) );
  NAND U17209 ( .A(n16255), .B(n16254), .Z(n16394) );
  XNOR U17210 ( .A(b[31]), .B(a[90]), .Z(n16379) );
  NANDN U17211 ( .A(n16379), .B(n38552), .Z(n16258) );
  NANDN U17212 ( .A(n16256), .B(n38553), .Z(n16257) );
  NAND U17213 ( .A(n16258), .B(n16257), .Z(n16391) );
  OR U17214 ( .A(n16259), .B(n36105), .Z(n16261) );
  XOR U17215 ( .A(b[3]), .B(n20271), .Z(n16382) );
  NANDN U17216 ( .A(n16382), .B(n36107), .Z(n16260) );
  AND U17217 ( .A(n16261), .B(n16260), .Z(n16392) );
  XNOR U17218 ( .A(n16391), .B(n16392), .Z(n16393) );
  XOR U17219 ( .A(n16394), .B(n16393), .Z(n16421) );
  XNOR U17220 ( .A(n16422), .B(n16421), .Z(n16423) );
  XNOR U17221 ( .A(n16424), .B(n16423), .Z(n16470) );
  XNOR U17222 ( .A(n16469), .B(n16470), .Z(n16471) );
  XNOR U17223 ( .A(n16472), .B(n16471), .Z(n16358) );
  NANDN U17224 ( .A(n16267), .B(n16266), .Z(n16271) );
  NANDN U17225 ( .A(n16269), .B(n16268), .Z(n16270) );
  NAND U17226 ( .A(n16271), .B(n16270), .Z(n16477) );
  OR U17227 ( .A(n16273), .B(n16272), .Z(n16277) );
  NAND U17228 ( .A(n16275), .B(n16274), .Z(n16276) );
  NAND U17229 ( .A(n16277), .B(n16276), .Z(n16476) );
  NANDN U17230 ( .A(n16279), .B(n16278), .Z(n16283) );
  NAND U17231 ( .A(n16281), .B(n16280), .Z(n16282) );
  NAND U17232 ( .A(n16283), .B(n16282), .Z(n16415) );
  NANDN U17233 ( .A(n16285), .B(n16284), .Z(n16289) );
  NAND U17234 ( .A(n16287), .B(n16286), .Z(n16288) );
  AND U17235 ( .A(n16289), .B(n16288), .Z(n16416) );
  XNOR U17236 ( .A(n16415), .B(n16416), .Z(n16417) );
  XNOR U17237 ( .A(n1052), .B(a[112]), .Z(n16439) );
  NAND U17238 ( .A(n36925), .B(n16439), .Z(n16292) );
  NANDN U17239 ( .A(n16290), .B(n36926), .Z(n16291) );
  NAND U17240 ( .A(n16292), .B(n16291), .Z(n16399) );
  XNOR U17241 ( .A(b[15]), .B(a[106]), .Z(n16442) );
  OR U17242 ( .A(n16442), .B(n37665), .Z(n16295) );
  NANDN U17243 ( .A(n16293), .B(n37604), .Z(n16294) );
  AND U17244 ( .A(n16295), .B(n16294), .Z(n16397) );
  XNOR U17245 ( .A(n1056), .B(a[100]), .Z(n16445) );
  NAND U17246 ( .A(n16445), .B(n38101), .Z(n16298) );
  NANDN U17247 ( .A(n16296), .B(n38102), .Z(n16297) );
  AND U17248 ( .A(n16298), .B(n16297), .Z(n16398) );
  XOR U17249 ( .A(n16399), .B(n16400), .Z(n16388) );
  XNOR U17250 ( .A(b[11]), .B(a[110]), .Z(n16448) );
  OR U17251 ( .A(n16448), .B(n37311), .Z(n16301) );
  NANDN U17252 ( .A(n16299), .B(n37218), .Z(n16300) );
  NAND U17253 ( .A(n16301), .B(n16300), .Z(n16386) );
  XOR U17254 ( .A(n1053), .B(a[108]), .Z(n16451) );
  NANDN U17255 ( .A(n16451), .B(n37424), .Z(n16304) );
  NANDN U17256 ( .A(n16302), .B(n37425), .Z(n16303) );
  AND U17257 ( .A(n16304), .B(n16303), .Z(n16385) );
  XNOR U17258 ( .A(n16386), .B(n16385), .Z(n16387) );
  XOR U17259 ( .A(n16388), .B(n16387), .Z(n16405) );
  NANDN U17260 ( .A(n1049), .B(a[120]), .Z(n16305) );
  XNOR U17261 ( .A(b[1]), .B(n16305), .Z(n16307) );
  NANDN U17262 ( .A(b[0]), .B(a[119]), .Z(n16306) );
  AND U17263 ( .A(n16307), .B(n16306), .Z(n16363) );
  NAND U17264 ( .A(n38490), .B(n16308), .Z(n16310) );
  XNOR U17265 ( .A(n1058), .B(a[92]), .Z(n16457) );
  NANDN U17266 ( .A(n1048), .B(n16457), .Z(n16309) );
  NAND U17267 ( .A(n16310), .B(n16309), .Z(n16361) );
  NANDN U17268 ( .A(n1059), .B(a[88]), .Z(n16362) );
  XNOR U17269 ( .A(n16361), .B(n16362), .Z(n16364) );
  XOR U17270 ( .A(n16363), .B(n16364), .Z(n16403) );
  NANDN U17271 ( .A(n16311), .B(n38205), .Z(n16313) );
  XNOR U17272 ( .A(b[23]), .B(a[98]), .Z(n16460) );
  OR U17273 ( .A(n16460), .B(n38268), .Z(n16312) );
  NAND U17274 ( .A(n16313), .B(n16312), .Z(n16430) );
  XOR U17275 ( .A(b[7]), .B(a[114]), .Z(n16463) );
  NAND U17276 ( .A(n16463), .B(n36701), .Z(n16316) );
  NANDN U17277 ( .A(n16314), .B(n36702), .Z(n16315) );
  NAND U17278 ( .A(n16316), .B(n16315), .Z(n16427) );
  XOR U17279 ( .A(b[25]), .B(a[96]), .Z(n16466) );
  NAND U17280 ( .A(n16466), .B(n38325), .Z(n16319) );
  NAND U17281 ( .A(n16317), .B(n38326), .Z(n16318) );
  AND U17282 ( .A(n16319), .B(n16318), .Z(n16428) );
  XNOR U17283 ( .A(n16427), .B(n16428), .Z(n16429) );
  XNOR U17284 ( .A(n16430), .B(n16429), .Z(n16404) );
  XOR U17285 ( .A(n16403), .B(n16404), .Z(n16406) );
  XNOR U17286 ( .A(n16405), .B(n16406), .Z(n16418) );
  XNOR U17287 ( .A(n16417), .B(n16418), .Z(n16475) );
  XNOR U17288 ( .A(n16476), .B(n16475), .Z(n16478) );
  XNOR U17289 ( .A(n16477), .B(n16478), .Z(n16355) );
  XNOR U17290 ( .A(n16356), .B(n16355), .Z(n16357) );
  XOR U17291 ( .A(n16358), .B(n16357), .Z(n16352) );
  XOR U17292 ( .A(n16351), .B(n16352), .Z(n16346) );
  NANDN U17293 ( .A(n16321), .B(n16320), .Z(n16325) );
  NAND U17294 ( .A(n16323), .B(n16322), .Z(n16324) );
  NAND U17295 ( .A(n16325), .B(n16324), .Z(n16343) );
  NANDN U17296 ( .A(n16327), .B(n16326), .Z(n16331) );
  OR U17297 ( .A(n16329), .B(n16328), .Z(n16330) );
  NAND U17298 ( .A(n16331), .B(n16330), .Z(n16344) );
  XNOR U17299 ( .A(n16343), .B(n16344), .Z(n16345) );
  XNOR U17300 ( .A(n16346), .B(n16345), .Z(n16338) );
  XNOR U17301 ( .A(n16337), .B(n16338), .Z(n16339) );
  XNOR U17302 ( .A(n16340), .B(n16339), .Z(n16481) );
  XNOR U17303 ( .A(n16481), .B(sreg[344]), .Z(n16483) );
  NAND U17304 ( .A(n16332), .B(sreg[343]), .Z(n16336) );
  OR U17305 ( .A(n16334), .B(n16333), .Z(n16335) );
  AND U17306 ( .A(n16336), .B(n16335), .Z(n16482) );
  XOR U17307 ( .A(n16483), .B(n16482), .Z(c[344]) );
  NANDN U17308 ( .A(n16338), .B(n16337), .Z(n16342) );
  NAND U17309 ( .A(n16340), .B(n16339), .Z(n16341) );
  NAND U17310 ( .A(n16342), .B(n16341), .Z(n16489) );
  NANDN U17311 ( .A(n16344), .B(n16343), .Z(n16348) );
  NAND U17312 ( .A(n16346), .B(n16345), .Z(n16347) );
  NAND U17313 ( .A(n16348), .B(n16347), .Z(n16487) );
  NANDN U17314 ( .A(n16350), .B(n16349), .Z(n16354) );
  NANDN U17315 ( .A(n16352), .B(n16351), .Z(n16353) );
  NAND U17316 ( .A(n16354), .B(n16353), .Z(n16493) );
  NANDN U17317 ( .A(n16356), .B(n16355), .Z(n16360) );
  NANDN U17318 ( .A(n16358), .B(n16357), .Z(n16359) );
  AND U17319 ( .A(n16360), .B(n16359), .Z(n16492) );
  XNOR U17320 ( .A(n16493), .B(n16492), .Z(n16494) );
  NANDN U17321 ( .A(n16362), .B(n16361), .Z(n16366) );
  NAND U17322 ( .A(n16364), .B(n16363), .Z(n16365) );
  NAND U17323 ( .A(n16366), .B(n16365), .Z(n16571) );
  XNOR U17324 ( .A(b[19]), .B(a[103]), .Z(n16516) );
  NANDN U17325 ( .A(n16516), .B(n37934), .Z(n16369) );
  NANDN U17326 ( .A(n16367), .B(n37935), .Z(n16368) );
  NAND U17327 ( .A(n16369), .B(n16368), .Z(n16581) );
  XOR U17328 ( .A(b[27]), .B(a[95]), .Z(n16519) );
  NAND U17329 ( .A(n38423), .B(n16519), .Z(n16372) );
  NAND U17330 ( .A(n16370), .B(n38424), .Z(n16371) );
  NAND U17331 ( .A(n16372), .B(n16371), .Z(n16578) );
  XNOR U17332 ( .A(b[5]), .B(a[117]), .Z(n16522) );
  NANDN U17333 ( .A(n16522), .B(n36587), .Z(n16375) );
  NANDN U17334 ( .A(n16373), .B(n36588), .Z(n16374) );
  AND U17335 ( .A(n16375), .B(n16374), .Z(n16579) );
  XNOR U17336 ( .A(n16578), .B(n16579), .Z(n16580) );
  XNOR U17337 ( .A(n16581), .B(n16580), .Z(n16569) );
  NAND U17338 ( .A(n16376), .B(n37762), .Z(n16378) );
  XOR U17339 ( .A(b[17]), .B(a[105]), .Z(n16525) );
  NAND U17340 ( .A(n16525), .B(n37764), .Z(n16377) );
  NAND U17341 ( .A(n16378), .B(n16377), .Z(n16543) );
  XNOR U17342 ( .A(b[31]), .B(a[91]), .Z(n16528) );
  NANDN U17343 ( .A(n16528), .B(n38552), .Z(n16381) );
  NANDN U17344 ( .A(n16379), .B(n38553), .Z(n16380) );
  NAND U17345 ( .A(n16381), .B(n16380), .Z(n16540) );
  OR U17346 ( .A(n16382), .B(n36105), .Z(n16384) );
  XNOR U17347 ( .A(b[3]), .B(a[119]), .Z(n16531) );
  NANDN U17348 ( .A(n16531), .B(n36107), .Z(n16383) );
  AND U17349 ( .A(n16384), .B(n16383), .Z(n16541) );
  XNOR U17350 ( .A(n16540), .B(n16541), .Z(n16542) );
  XOR U17351 ( .A(n16543), .B(n16542), .Z(n16568) );
  XNOR U17352 ( .A(n16569), .B(n16568), .Z(n16570) );
  XNOR U17353 ( .A(n16571), .B(n16570), .Z(n16614) );
  NANDN U17354 ( .A(n16386), .B(n16385), .Z(n16390) );
  NAND U17355 ( .A(n16388), .B(n16387), .Z(n16389) );
  NAND U17356 ( .A(n16390), .B(n16389), .Z(n16559) );
  NANDN U17357 ( .A(n16392), .B(n16391), .Z(n16396) );
  NAND U17358 ( .A(n16394), .B(n16393), .Z(n16395) );
  NAND U17359 ( .A(n16396), .B(n16395), .Z(n16557) );
  OR U17360 ( .A(n16398), .B(n16397), .Z(n16402) );
  NANDN U17361 ( .A(n16400), .B(n16399), .Z(n16401) );
  NAND U17362 ( .A(n16402), .B(n16401), .Z(n16556) );
  XNOR U17363 ( .A(n16559), .B(n16558), .Z(n16615) );
  XOR U17364 ( .A(n16614), .B(n16615), .Z(n16617) );
  NANDN U17365 ( .A(n16404), .B(n16403), .Z(n16408) );
  OR U17366 ( .A(n16406), .B(n16405), .Z(n16407) );
  NAND U17367 ( .A(n16408), .B(n16407), .Z(n16616) );
  XOR U17368 ( .A(n16617), .B(n16616), .Z(n16506) );
  OR U17369 ( .A(n16410), .B(n16409), .Z(n16414) );
  NANDN U17370 ( .A(n16412), .B(n16411), .Z(n16413) );
  NAND U17371 ( .A(n16414), .B(n16413), .Z(n16505) );
  NANDN U17372 ( .A(n16416), .B(n16415), .Z(n16420) );
  NANDN U17373 ( .A(n16418), .B(n16417), .Z(n16419) );
  NAND U17374 ( .A(n16420), .B(n16419), .Z(n16622) );
  NANDN U17375 ( .A(n16422), .B(n16421), .Z(n16426) );
  NAND U17376 ( .A(n16424), .B(n16423), .Z(n16425) );
  NAND U17377 ( .A(n16426), .B(n16425), .Z(n16621) );
  NANDN U17378 ( .A(n16428), .B(n16427), .Z(n16432) );
  NAND U17379 ( .A(n16430), .B(n16429), .Z(n16431) );
  NAND U17380 ( .A(n16432), .B(n16431), .Z(n16562) );
  NANDN U17381 ( .A(n16434), .B(n16433), .Z(n16438) );
  NAND U17382 ( .A(n16436), .B(n16435), .Z(n16437) );
  AND U17383 ( .A(n16438), .B(n16437), .Z(n16563) );
  XNOR U17384 ( .A(n16562), .B(n16563), .Z(n16564) );
  XOR U17385 ( .A(n1052), .B(a[113]), .Z(n16590) );
  NANDN U17386 ( .A(n16590), .B(n36925), .Z(n16441) );
  NAND U17387 ( .A(n36926), .B(n16439), .Z(n16440) );
  NAND U17388 ( .A(n16441), .B(n16440), .Z(n16548) );
  XNOR U17389 ( .A(n1054), .B(a[107]), .Z(n16587) );
  NANDN U17390 ( .A(n37665), .B(n16587), .Z(n16444) );
  NANDN U17391 ( .A(n16442), .B(n37604), .Z(n16443) );
  NAND U17392 ( .A(n16444), .B(n16443), .Z(n16546) );
  XOR U17393 ( .A(n1056), .B(a[101]), .Z(n16584) );
  NANDN U17394 ( .A(n16584), .B(n38101), .Z(n16447) );
  NAND U17395 ( .A(n38102), .B(n16445), .Z(n16446) );
  NAND U17396 ( .A(n16447), .B(n16446), .Z(n16547) );
  XNOR U17397 ( .A(n16546), .B(n16547), .Z(n16549) );
  XOR U17398 ( .A(n16548), .B(n16549), .Z(n16537) );
  XNOR U17399 ( .A(b[11]), .B(a[111]), .Z(n16593) );
  OR U17400 ( .A(n16593), .B(n37311), .Z(n16450) );
  NANDN U17401 ( .A(n16448), .B(n37218), .Z(n16449) );
  NAND U17402 ( .A(n16450), .B(n16449), .Z(n16535) );
  XOR U17403 ( .A(n1053), .B(a[109]), .Z(n16596) );
  NANDN U17404 ( .A(n16596), .B(n37424), .Z(n16453) );
  NANDN U17405 ( .A(n16451), .B(n37425), .Z(n16452) );
  AND U17406 ( .A(n16453), .B(n16452), .Z(n16534) );
  XNOR U17407 ( .A(n16535), .B(n16534), .Z(n16536) );
  XNOR U17408 ( .A(n16537), .B(n16536), .Z(n16553) );
  NANDN U17409 ( .A(n1049), .B(a[121]), .Z(n16454) );
  XNOR U17410 ( .A(b[1]), .B(n16454), .Z(n16456) );
  NANDN U17411 ( .A(b[0]), .B(a[120]), .Z(n16455) );
  AND U17412 ( .A(n16456), .B(n16455), .Z(n16512) );
  NAND U17413 ( .A(n38490), .B(n16457), .Z(n16459) );
  XOR U17414 ( .A(n1058), .B(n17031), .Z(n16602) );
  NANDN U17415 ( .A(n1048), .B(n16602), .Z(n16458) );
  NAND U17416 ( .A(n16459), .B(n16458), .Z(n16510) );
  NANDN U17417 ( .A(n1059), .B(a[89]), .Z(n16511) );
  XNOR U17418 ( .A(n16510), .B(n16511), .Z(n16513) );
  XNOR U17419 ( .A(n16512), .B(n16513), .Z(n16551) );
  NANDN U17420 ( .A(n16460), .B(n38205), .Z(n16462) );
  XOR U17421 ( .A(b[23]), .B(n17884), .Z(n16605) );
  OR U17422 ( .A(n16605), .B(n38268), .Z(n16461) );
  NAND U17423 ( .A(n16462), .B(n16461), .Z(n16575) );
  XOR U17424 ( .A(b[7]), .B(a[115]), .Z(n16608) );
  NAND U17425 ( .A(n16608), .B(n36701), .Z(n16465) );
  NAND U17426 ( .A(n16463), .B(n36702), .Z(n16464) );
  NAND U17427 ( .A(n16465), .B(n16464), .Z(n16572) );
  XOR U17428 ( .A(b[25]), .B(a[97]), .Z(n16611) );
  NAND U17429 ( .A(n16611), .B(n38325), .Z(n16468) );
  NAND U17430 ( .A(n16466), .B(n38326), .Z(n16467) );
  AND U17431 ( .A(n16468), .B(n16467), .Z(n16573) );
  XNOR U17432 ( .A(n16572), .B(n16573), .Z(n16574) );
  XOR U17433 ( .A(n16575), .B(n16574), .Z(n16550) );
  XOR U17434 ( .A(n16553), .B(n16552), .Z(n16565) );
  XOR U17435 ( .A(n16564), .B(n16565), .Z(n16620) );
  XNOR U17436 ( .A(n16621), .B(n16620), .Z(n16623) );
  XNOR U17437 ( .A(n16622), .B(n16623), .Z(n16504) );
  XOR U17438 ( .A(n16505), .B(n16504), .Z(n16507) );
  NANDN U17439 ( .A(n16470), .B(n16469), .Z(n16474) );
  NAND U17440 ( .A(n16472), .B(n16471), .Z(n16473) );
  NAND U17441 ( .A(n16474), .B(n16473), .Z(n16499) );
  NAND U17442 ( .A(n16476), .B(n16475), .Z(n16480) );
  NANDN U17443 ( .A(n16478), .B(n16477), .Z(n16479) );
  AND U17444 ( .A(n16480), .B(n16479), .Z(n16498) );
  XNOR U17445 ( .A(n16499), .B(n16498), .Z(n16500) );
  XOR U17446 ( .A(n16501), .B(n16500), .Z(n16495) );
  XOR U17447 ( .A(n16494), .B(n16495), .Z(n16486) );
  XOR U17448 ( .A(n16487), .B(n16486), .Z(n16488) );
  XNOR U17449 ( .A(n16489), .B(n16488), .Z(n16626) );
  XNOR U17450 ( .A(n16626), .B(sreg[345]), .Z(n16628) );
  NAND U17451 ( .A(n16481), .B(sreg[344]), .Z(n16485) );
  OR U17452 ( .A(n16483), .B(n16482), .Z(n16484) );
  AND U17453 ( .A(n16485), .B(n16484), .Z(n16627) );
  XOR U17454 ( .A(n16628), .B(n16627), .Z(c[345]) );
  NAND U17455 ( .A(n16487), .B(n16486), .Z(n16491) );
  NAND U17456 ( .A(n16489), .B(n16488), .Z(n16490) );
  NAND U17457 ( .A(n16491), .B(n16490), .Z(n16634) );
  NANDN U17458 ( .A(n16493), .B(n16492), .Z(n16497) );
  NAND U17459 ( .A(n16495), .B(n16494), .Z(n16496) );
  NAND U17460 ( .A(n16497), .B(n16496), .Z(n16632) );
  NANDN U17461 ( .A(n16499), .B(n16498), .Z(n16503) );
  NAND U17462 ( .A(n16501), .B(n16500), .Z(n16502) );
  NAND U17463 ( .A(n16503), .B(n16502), .Z(n16637) );
  NANDN U17464 ( .A(n16505), .B(n16504), .Z(n16509) );
  OR U17465 ( .A(n16507), .B(n16506), .Z(n16508) );
  NAND U17466 ( .A(n16509), .B(n16508), .Z(n16638) );
  XNOR U17467 ( .A(n16637), .B(n16638), .Z(n16639) );
  NANDN U17468 ( .A(n16511), .B(n16510), .Z(n16515) );
  NAND U17469 ( .A(n16513), .B(n16512), .Z(n16514) );
  NAND U17470 ( .A(n16515), .B(n16514), .Z(n16712) );
  XNOR U17471 ( .A(b[19]), .B(a[104]), .Z(n16659) );
  NANDN U17472 ( .A(n16659), .B(n37934), .Z(n16518) );
  NANDN U17473 ( .A(n16516), .B(n37935), .Z(n16517) );
  NAND U17474 ( .A(n16518), .B(n16517), .Z(n16722) );
  XOR U17475 ( .A(b[27]), .B(a[96]), .Z(n16662) );
  NAND U17476 ( .A(n38423), .B(n16662), .Z(n16521) );
  NAND U17477 ( .A(n16519), .B(n38424), .Z(n16520) );
  NAND U17478 ( .A(n16521), .B(n16520), .Z(n16719) );
  XOR U17479 ( .A(b[5]), .B(n20271), .Z(n16665) );
  NANDN U17480 ( .A(n16665), .B(n36587), .Z(n16524) );
  NANDN U17481 ( .A(n16522), .B(n36588), .Z(n16523) );
  AND U17482 ( .A(n16524), .B(n16523), .Z(n16720) );
  XNOR U17483 ( .A(n16719), .B(n16720), .Z(n16721) );
  XNOR U17484 ( .A(n16722), .B(n16721), .Z(n16710) );
  NAND U17485 ( .A(n16525), .B(n37762), .Z(n16527) );
  XOR U17486 ( .A(b[17]), .B(a[106]), .Z(n16668) );
  NAND U17487 ( .A(n16668), .B(n37764), .Z(n16526) );
  NAND U17488 ( .A(n16527), .B(n16526), .Z(n16686) );
  XNOR U17489 ( .A(b[31]), .B(a[92]), .Z(n16671) );
  NANDN U17490 ( .A(n16671), .B(n38552), .Z(n16530) );
  NANDN U17491 ( .A(n16528), .B(n38553), .Z(n16529) );
  NAND U17492 ( .A(n16530), .B(n16529), .Z(n16683) );
  OR U17493 ( .A(n16531), .B(n36105), .Z(n16533) );
  XNOR U17494 ( .A(b[3]), .B(a[120]), .Z(n16674) );
  NANDN U17495 ( .A(n16674), .B(n36107), .Z(n16532) );
  AND U17496 ( .A(n16533), .B(n16532), .Z(n16684) );
  XNOR U17497 ( .A(n16683), .B(n16684), .Z(n16685) );
  XOR U17498 ( .A(n16686), .B(n16685), .Z(n16709) );
  XNOR U17499 ( .A(n16710), .B(n16709), .Z(n16711) );
  XNOR U17500 ( .A(n16712), .B(n16711), .Z(n16650) );
  NANDN U17501 ( .A(n16535), .B(n16534), .Z(n16539) );
  NAND U17502 ( .A(n16537), .B(n16536), .Z(n16538) );
  NAND U17503 ( .A(n16539), .B(n16538), .Z(n16701) );
  NANDN U17504 ( .A(n16541), .B(n16540), .Z(n16545) );
  NAND U17505 ( .A(n16543), .B(n16542), .Z(n16544) );
  NAND U17506 ( .A(n16545), .B(n16544), .Z(n16700) );
  XNOR U17507 ( .A(n16700), .B(n16699), .Z(n16702) );
  XOR U17508 ( .A(n16701), .B(n16702), .Z(n16649) );
  XOR U17509 ( .A(n16650), .B(n16649), .Z(n16651) );
  NANDN U17510 ( .A(n16551), .B(n16550), .Z(n16555) );
  NAND U17511 ( .A(n16553), .B(n16552), .Z(n16554) );
  NAND U17512 ( .A(n16555), .B(n16554), .Z(n16652) );
  XNOR U17513 ( .A(n16651), .B(n16652), .Z(n16763) );
  OR U17514 ( .A(n16557), .B(n16556), .Z(n16561) );
  NAND U17515 ( .A(n16559), .B(n16558), .Z(n16560) );
  NAND U17516 ( .A(n16561), .B(n16560), .Z(n16762) );
  NANDN U17517 ( .A(n16563), .B(n16562), .Z(n16567) );
  NAND U17518 ( .A(n16565), .B(n16564), .Z(n16566) );
  NAND U17519 ( .A(n16567), .B(n16566), .Z(n16645) );
  NANDN U17520 ( .A(n16573), .B(n16572), .Z(n16577) );
  NAND U17521 ( .A(n16575), .B(n16574), .Z(n16576) );
  NAND U17522 ( .A(n16577), .B(n16576), .Z(n16703) );
  NANDN U17523 ( .A(n16579), .B(n16578), .Z(n16583) );
  NAND U17524 ( .A(n16581), .B(n16580), .Z(n16582) );
  AND U17525 ( .A(n16583), .B(n16582), .Z(n16704) );
  XNOR U17526 ( .A(n16703), .B(n16704), .Z(n16705) );
  XNOR U17527 ( .A(b[21]), .B(a[102]), .Z(n16731) );
  NANDN U17528 ( .A(n16731), .B(n38101), .Z(n16586) );
  NANDN U17529 ( .A(n16584), .B(n38102), .Z(n16585) );
  NAND U17530 ( .A(n16586), .B(n16585), .Z(n16695) );
  XNOR U17531 ( .A(b[15]), .B(a[108]), .Z(n16728) );
  OR U17532 ( .A(n16728), .B(n37665), .Z(n16589) );
  NAND U17533 ( .A(n16587), .B(n37604), .Z(n16588) );
  AND U17534 ( .A(n16589), .B(n16588), .Z(n16696) );
  XNOR U17535 ( .A(n16695), .B(n16696), .Z(n16698) );
  XNOR U17536 ( .A(b[9]), .B(a[114]), .Z(n16725) );
  NANDN U17537 ( .A(n16725), .B(n36925), .Z(n16592) );
  NANDN U17538 ( .A(n16590), .B(n36926), .Z(n16591) );
  NAND U17539 ( .A(n16592), .B(n16591), .Z(n16697) );
  XNOR U17540 ( .A(n16698), .B(n16697), .Z(n16691) );
  XNOR U17541 ( .A(b[11]), .B(a[112]), .Z(n16734) );
  OR U17542 ( .A(n16734), .B(n37311), .Z(n16595) );
  NANDN U17543 ( .A(n16593), .B(n37218), .Z(n16594) );
  NAND U17544 ( .A(n16595), .B(n16594), .Z(n16690) );
  XOR U17545 ( .A(n1053), .B(a[110]), .Z(n16737) );
  NANDN U17546 ( .A(n16737), .B(n37424), .Z(n16598) );
  NANDN U17547 ( .A(n16596), .B(n37425), .Z(n16597) );
  NAND U17548 ( .A(n16598), .B(n16597), .Z(n16689) );
  XNOR U17549 ( .A(n16690), .B(n16689), .Z(n16692) );
  XNOR U17550 ( .A(n16691), .B(n16692), .Z(n16680) );
  NANDN U17551 ( .A(n1049), .B(a[122]), .Z(n16599) );
  XNOR U17552 ( .A(b[1]), .B(n16599), .Z(n16601) );
  NANDN U17553 ( .A(b[0]), .B(a[121]), .Z(n16600) );
  AND U17554 ( .A(n16601), .B(n16600), .Z(n16655) );
  NAND U17555 ( .A(n38490), .B(n16602), .Z(n16604) );
  XNOR U17556 ( .A(n1058), .B(a[94]), .Z(n16740) );
  NANDN U17557 ( .A(n1048), .B(n16740), .Z(n16603) );
  NAND U17558 ( .A(n16604), .B(n16603), .Z(n16653) );
  NANDN U17559 ( .A(n1059), .B(a[90]), .Z(n16654) );
  XNOR U17560 ( .A(n16653), .B(n16654), .Z(n16656) );
  XNOR U17561 ( .A(n16655), .B(n16656), .Z(n16678) );
  NANDN U17562 ( .A(n16605), .B(n38205), .Z(n16607) );
  XNOR U17563 ( .A(b[23]), .B(a[100]), .Z(n16746) );
  OR U17564 ( .A(n16746), .B(n38268), .Z(n16606) );
  NAND U17565 ( .A(n16607), .B(n16606), .Z(n16716) );
  XOR U17566 ( .A(b[7]), .B(a[116]), .Z(n16749) );
  NAND U17567 ( .A(n16749), .B(n36701), .Z(n16610) );
  NAND U17568 ( .A(n16608), .B(n36702), .Z(n16609) );
  NAND U17569 ( .A(n16610), .B(n16609), .Z(n16713) );
  XOR U17570 ( .A(b[25]), .B(a[98]), .Z(n16752) );
  NAND U17571 ( .A(n16752), .B(n38325), .Z(n16613) );
  NAND U17572 ( .A(n16611), .B(n38326), .Z(n16612) );
  AND U17573 ( .A(n16613), .B(n16612), .Z(n16714) );
  XNOR U17574 ( .A(n16713), .B(n16714), .Z(n16715) );
  XOR U17575 ( .A(n16716), .B(n16715), .Z(n16677) );
  XOR U17576 ( .A(n16680), .B(n16679), .Z(n16706) );
  XNOR U17577 ( .A(n16705), .B(n16706), .Z(n16643) );
  XNOR U17578 ( .A(n16644), .B(n16643), .Z(n16646) );
  XNOR U17579 ( .A(n16645), .B(n16646), .Z(n16761) );
  XOR U17580 ( .A(n16762), .B(n16761), .Z(n16764) );
  NANDN U17581 ( .A(n16615), .B(n16614), .Z(n16619) );
  OR U17582 ( .A(n16617), .B(n16616), .Z(n16618) );
  NAND U17583 ( .A(n16619), .B(n16618), .Z(n16755) );
  NAND U17584 ( .A(n16621), .B(n16620), .Z(n16625) );
  NANDN U17585 ( .A(n16623), .B(n16622), .Z(n16624) );
  NAND U17586 ( .A(n16625), .B(n16624), .Z(n16756) );
  XNOR U17587 ( .A(n16755), .B(n16756), .Z(n16757) );
  XOR U17588 ( .A(n16758), .B(n16757), .Z(n16640) );
  XOR U17589 ( .A(n16639), .B(n16640), .Z(n16631) );
  XOR U17590 ( .A(n16632), .B(n16631), .Z(n16633) );
  XNOR U17591 ( .A(n16634), .B(n16633), .Z(n16767) );
  XNOR U17592 ( .A(n16767), .B(sreg[346]), .Z(n16769) );
  NAND U17593 ( .A(n16626), .B(sreg[345]), .Z(n16630) );
  OR U17594 ( .A(n16628), .B(n16627), .Z(n16629) );
  AND U17595 ( .A(n16630), .B(n16629), .Z(n16768) );
  XOR U17596 ( .A(n16769), .B(n16768), .Z(c[346]) );
  NAND U17597 ( .A(n16632), .B(n16631), .Z(n16636) );
  NAND U17598 ( .A(n16634), .B(n16633), .Z(n16635) );
  NAND U17599 ( .A(n16636), .B(n16635), .Z(n16775) );
  NANDN U17600 ( .A(n16638), .B(n16637), .Z(n16642) );
  NAND U17601 ( .A(n16640), .B(n16639), .Z(n16641) );
  NAND U17602 ( .A(n16642), .B(n16641), .Z(n16772) );
  NAND U17603 ( .A(n16644), .B(n16643), .Z(n16648) );
  NANDN U17604 ( .A(n16646), .B(n16645), .Z(n16647) );
  NAND U17605 ( .A(n16648), .B(n16647), .Z(n16900) );
  XNOR U17606 ( .A(n16900), .B(n16901), .Z(n16902) );
  NANDN U17607 ( .A(n16654), .B(n16653), .Z(n16658) );
  NAND U17608 ( .A(n16656), .B(n16655), .Z(n16657) );
  NAND U17609 ( .A(n16658), .B(n16657), .Z(n16845) );
  XNOR U17610 ( .A(b[19]), .B(a[105]), .Z(n16790) );
  NANDN U17611 ( .A(n16790), .B(n37934), .Z(n16661) );
  NANDN U17612 ( .A(n16659), .B(n37935), .Z(n16660) );
  NAND U17613 ( .A(n16661), .B(n16660), .Z(n16855) );
  XOR U17614 ( .A(b[27]), .B(a[97]), .Z(n16793) );
  NAND U17615 ( .A(n38423), .B(n16793), .Z(n16664) );
  NAND U17616 ( .A(n16662), .B(n38424), .Z(n16663) );
  NAND U17617 ( .A(n16664), .B(n16663), .Z(n16852) );
  XNOR U17618 ( .A(b[5]), .B(a[119]), .Z(n16796) );
  NANDN U17619 ( .A(n16796), .B(n36587), .Z(n16667) );
  NANDN U17620 ( .A(n16665), .B(n36588), .Z(n16666) );
  AND U17621 ( .A(n16667), .B(n16666), .Z(n16853) );
  XNOR U17622 ( .A(n16852), .B(n16853), .Z(n16854) );
  XNOR U17623 ( .A(n16855), .B(n16854), .Z(n16843) );
  NAND U17624 ( .A(n16668), .B(n37762), .Z(n16670) );
  XNOR U17625 ( .A(b[17]), .B(a[107]), .Z(n16799) );
  NANDN U17626 ( .A(n16799), .B(n37764), .Z(n16669) );
  NAND U17627 ( .A(n16670), .B(n16669), .Z(n16817) );
  XOR U17628 ( .A(b[31]), .B(n17031), .Z(n16802) );
  NANDN U17629 ( .A(n16802), .B(n38552), .Z(n16673) );
  NANDN U17630 ( .A(n16671), .B(n38553), .Z(n16672) );
  NAND U17631 ( .A(n16673), .B(n16672), .Z(n16814) );
  OR U17632 ( .A(n16674), .B(n36105), .Z(n16676) );
  XNOR U17633 ( .A(b[3]), .B(a[121]), .Z(n16805) );
  NANDN U17634 ( .A(n16805), .B(n36107), .Z(n16675) );
  AND U17635 ( .A(n16676), .B(n16675), .Z(n16815) );
  XNOR U17636 ( .A(n16814), .B(n16815), .Z(n16816) );
  XOR U17637 ( .A(n16817), .B(n16816), .Z(n16842) );
  XNOR U17638 ( .A(n16843), .B(n16842), .Z(n16844) );
  XNOR U17639 ( .A(n16845), .B(n16844), .Z(n16894) );
  NANDN U17640 ( .A(n16678), .B(n16677), .Z(n16682) );
  NANDN U17641 ( .A(n16680), .B(n16679), .Z(n16681) );
  NAND U17642 ( .A(n16682), .B(n16681), .Z(n16895) );
  XNOR U17643 ( .A(n16894), .B(n16895), .Z(n16896) );
  NANDN U17644 ( .A(n16684), .B(n16683), .Z(n16688) );
  NAND U17645 ( .A(n16686), .B(n16685), .Z(n16687) );
  NAND U17646 ( .A(n16688), .B(n16687), .Z(n16835) );
  OR U17647 ( .A(n16690), .B(n16689), .Z(n16694) );
  NANDN U17648 ( .A(n16692), .B(n16691), .Z(n16693) );
  NAND U17649 ( .A(n16694), .B(n16693), .Z(n16833) );
  XNOR U17650 ( .A(n16833), .B(n16832), .Z(n16834) );
  XOR U17651 ( .A(n16835), .B(n16834), .Z(n16897) );
  XOR U17652 ( .A(n16896), .B(n16897), .Z(n16908) );
  NANDN U17653 ( .A(n16704), .B(n16703), .Z(n16708) );
  NANDN U17654 ( .A(n16706), .B(n16705), .Z(n16707) );
  NAND U17655 ( .A(n16708), .B(n16707), .Z(n16891) );
  NANDN U17656 ( .A(n16714), .B(n16713), .Z(n16718) );
  NAND U17657 ( .A(n16716), .B(n16715), .Z(n16717) );
  NAND U17658 ( .A(n16718), .B(n16717), .Z(n16836) );
  NANDN U17659 ( .A(n16720), .B(n16719), .Z(n16724) );
  NAND U17660 ( .A(n16722), .B(n16721), .Z(n16723) );
  AND U17661 ( .A(n16724), .B(n16723), .Z(n16837) );
  XNOR U17662 ( .A(n16836), .B(n16837), .Z(n16838) );
  XNOR U17663 ( .A(b[9]), .B(a[115]), .Z(n16858) );
  NANDN U17664 ( .A(n16858), .B(n36925), .Z(n16727) );
  NANDN U17665 ( .A(n16725), .B(n36926), .Z(n16726) );
  NAND U17666 ( .A(n16727), .B(n16726), .Z(n16822) );
  XNOR U17667 ( .A(b[15]), .B(a[109]), .Z(n16861) );
  OR U17668 ( .A(n16861), .B(n37665), .Z(n16730) );
  NANDN U17669 ( .A(n16728), .B(n37604), .Z(n16729) );
  AND U17670 ( .A(n16730), .B(n16729), .Z(n16820) );
  XNOR U17671 ( .A(b[21]), .B(a[103]), .Z(n16864) );
  NANDN U17672 ( .A(n16864), .B(n38101), .Z(n16733) );
  NANDN U17673 ( .A(n16731), .B(n38102), .Z(n16732) );
  AND U17674 ( .A(n16733), .B(n16732), .Z(n16821) );
  XOR U17675 ( .A(n16822), .B(n16823), .Z(n16811) );
  XOR U17676 ( .A(b[11]), .B(n19909), .Z(n16867) );
  OR U17677 ( .A(n16867), .B(n37311), .Z(n16736) );
  NANDN U17678 ( .A(n16734), .B(n37218), .Z(n16735) );
  NAND U17679 ( .A(n16736), .B(n16735), .Z(n16809) );
  XOR U17680 ( .A(n1053), .B(a[111]), .Z(n16870) );
  NANDN U17681 ( .A(n16870), .B(n37424), .Z(n16739) );
  NANDN U17682 ( .A(n16737), .B(n37425), .Z(n16738) );
  AND U17683 ( .A(n16739), .B(n16738), .Z(n16808) );
  XNOR U17684 ( .A(n16809), .B(n16808), .Z(n16810) );
  XOR U17685 ( .A(n16811), .B(n16810), .Z(n16828) );
  NAND U17686 ( .A(n38490), .B(n16740), .Z(n16742) );
  XNOR U17687 ( .A(n1058), .B(a[95]), .Z(n16876) );
  NANDN U17688 ( .A(n1048), .B(n16876), .Z(n16741) );
  NAND U17689 ( .A(n16742), .B(n16741), .Z(n16784) );
  NANDN U17690 ( .A(n1059), .B(a[91]), .Z(n16785) );
  XNOR U17691 ( .A(n16784), .B(n16785), .Z(n16787) );
  NANDN U17692 ( .A(n1049), .B(a[123]), .Z(n16743) );
  XNOR U17693 ( .A(b[1]), .B(n16743), .Z(n16745) );
  NANDN U17694 ( .A(b[0]), .B(a[122]), .Z(n16744) );
  AND U17695 ( .A(n16745), .B(n16744), .Z(n16786) );
  XOR U17696 ( .A(n16787), .B(n16786), .Z(n16826) );
  NANDN U17697 ( .A(n16746), .B(n38205), .Z(n16748) );
  XOR U17698 ( .A(b[23]), .B(n17812), .Z(n16879) );
  OR U17699 ( .A(n16879), .B(n38268), .Z(n16747) );
  NAND U17700 ( .A(n16748), .B(n16747), .Z(n16849) );
  XOR U17701 ( .A(b[7]), .B(a[117]), .Z(n16882) );
  NAND U17702 ( .A(n16882), .B(n36701), .Z(n16751) );
  NAND U17703 ( .A(n16749), .B(n36702), .Z(n16750) );
  NAND U17704 ( .A(n16751), .B(n16750), .Z(n16846) );
  XNOR U17705 ( .A(b[25]), .B(a[99]), .Z(n16885) );
  NANDN U17706 ( .A(n16885), .B(n38325), .Z(n16754) );
  NAND U17707 ( .A(n16752), .B(n38326), .Z(n16753) );
  AND U17708 ( .A(n16754), .B(n16753), .Z(n16847) );
  XNOR U17709 ( .A(n16846), .B(n16847), .Z(n16848) );
  XNOR U17710 ( .A(n16849), .B(n16848), .Z(n16827) );
  XOR U17711 ( .A(n16826), .B(n16827), .Z(n16829) );
  XNOR U17712 ( .A(n16828), .B(n16829), .Z(n16839) );
  XOR U17713 ( .A(n16838), .B(n16839), .Z(n16889) );
  XNOR U17714 ( .A(n16888), .B(n16889), .Z(n16890) );
  XNOR U17715 ( .A(n16891), .B(n16890), .Z(n16906) );
  XNOR U17716 ( .A(n16907), .B(n16906), .Z(n16909) );
  XNOR U17717 ( .A(n16908), .B(n16909), .Z(n16903) );
  XOR U17718 ( .A(n16902), .B(n16903), .Z(n16781) );
  NANDN U17719 ( .A(n16756), .B(n16755), .Z(n16760) );
  NAND U17720 ( .A(n16758), .B(n16757), .Z(n16759) );
  NAND U17721 ( .A(n16760), .B(n16759), .Z(n16778) );
  NANDN U17722 ( .A(n16762), .B(n16761), .Z(n16766) );
  OR U17723 ( .A(n16764), .B(n16763), .Z(n16765) );
  NAND U17724 ( .A(n16766), .B(n16765), .Z(n16779) );
  XNOR U17725 ( .A(n16778), .B(n16779), .Z(n16780) );
  XNOR U17726 ( .A(n16781), .B(n16780), .Z(n16773) );
  XNOR U17727 ( .A(n16772), .B(n16773), .Z(n16774) );
  XNOR U17728 ( .A(n16775), .B(n16774), .Z(n16912) );
  XNOR U17729 ( .A(n16912), .B(sreg[347]), .Z(n16914) );
  NAND U17730 ( .A(n16767), .B(sreg[346]), .Z(n16771) );
  OR U17731 ( .A(n16769), .B(n16768), .Z(n16770) );
  AND U17732 ( .A(n16771), .B(n16770), .Z(n16913) );
  XOR U17733 ( .A(n16914), .B(n16913), .Z(c[347]) );
  NANDN U17734 ( .A(n16773), .B(n16772), .Z(n16777) );
  NAND U17735 ( .A(n16775), .B(n16774), .Z(n16776) );
  NAND U17736 ( .A(n16777), .B(n16776), .Z(n16920) );
  NANDN U17737 ( .A(n16779), .B(n16778), .Z(n16783) );
  NAND U17738 ( .A(n16781), .B(n16780), .Z(n16782) );
  NAND U17739 ( .A(n16783), .B(n16782), .Z(n16918) );
  NANDN U17740 ( .A(n16785), .B(n16784), .Z(n16789) );
  NAND U17741 ( .A(n16787), .B(n16786), .Z(n16788) );
  NAND U17742 ( .A(n16789), .B(n16788), .Z(n17000) );
  XNOR U17743 ( .A(b[19]), .B(a[106]), .Z(n16943) );
  NANDN U17744 ( .A(n16943), .B(n37934), .Z(n16792) );
  NANDN U17745 ( .A(n16790), .B(n37935), .Z(n16791) );
  NAND U17746 ( .A(n16792), .B(n16791), .Z(n17010) );
  XOR U17747 ( .A(b[27]), .B(a[98]), .Z(n16946) );
  NAND U17748 ( .A(n38423), .B(n16946), .Z(n16795) );
  NAND U17749 ( .A(n16793), .B(n38424), .Z(n16794) );
  NAND U17750 ( .A(n16795), .B(n16794), .Z(n17007) );
  XNOR U17751 ( .A(b[5]), .B(a[120]), .Z(n16949) );
  NANDN U17752 ( .A(n16949), .B(n36587), .Z(n16798) );
  NANDN U17753 ( .A(n16796), .B(n36588), .Z(n16797) );
  AND U17754 ( .A(n16798), .B(n16797), .Z(n17008) );
  XNOR U17755 ( .A(n17007), .B(n17008), .Z(n17009) );
  XNOR U17756 ( .A(n17010), .B(n17009), .Z(n16998) );
  NANDN U17757 ( .A(n16799), .B(n37762), .Z(n16801) );
  XOR U17758 ( .A(b[17]), .B(a[108]), .Z(n16952) );
  NAND U17759 ( .A(n16952), .B(n37764), .Z(n16800) );
  NAND U17760 ( .A(n16801), .B(n16800), .Z(n16970) );
  XNOR U17761 ( .A(n1059), .B(a[94]), .Z(n16955) );
  NAND U17762 ( .A(n16955), .B(n38552), .Z(n16804) );
  NANDN U17763 ( .A(n16802), .B(n38553), .Z(n16803) );
  NAND U17764 ( .A(n16804), .B(n16803), .Z(n16967) );
  OR U17765 ( .A(n16805), .B(n36105), .Z(n16807) );
  XNOR U17766 ( .A(b[3]), .B(a[122]), .Z(n16958) );
  NANDN U17767 ( .A(n16958), .B(n36107), .Z(n16806) );
  AND U17768 ( .A(n16807), .B(n16806), .Z(n16968) );
  XNOR U17769 ( .A(n16967), .B(n16968), .Z(n16969) );
  XOR U17770 ( .A(n16970), .B(n16969), .Z(n16997) );
  XNOR U17771 ( .A(n16998), .B(n16997), .Z(n16999) );
  XNOR U17772 ( .A(n17000), .B(n16999), .Z(n17044) );
  NANDN U17773 ( .A(n16809), .B(n16808), .Z(n16813) );
  NAND U17774 ( .A(n16811), .B(n16810), .Z(n16812) );
  NAND U17775 ( .A(n16813), .B(n16812), .Z(n16988) );
  NANDN U17776 ( .A(n16815), .B(n16814), .Z(n16819) );
  NAND U17777 ( .A(n16817), .B(n16816), .Z(n16818) );
  NAND U17778 ( .A(n16819), .B(n16818), .Z(n16986) );
  OR U17779 ( .A(n16821), .B(n16820), .Z(n16825) );
  NANDN U17780 ( .A(n16823), .B(n16822), .Z(n16824) );
  NAND U17781 ( .A(n16825), .B(n16824), .Z(n16985) );
  XNOR U17782 ( .A(n16988), .B(n16987), .Z(n17045) );
  XNOR U17783 ( .A(n17044), .B(n17045), .Z(n17046) );
  NANDN U17784 ( .A(n16827), .B(n16826), .Z(n16831) );
  OR U17785 ( .A(n16829), .B(n16828), .Z(n16830) );
  AND U17786 ( .A(n16831), .B(n16830), .Z(n17047) );
  XNOR U17787 ( .A(n17046), .B(n17047), .Z(n16930) );
  NANDN U17788 ( .A(n16837), .B(n16836), .Z(n16841) );
  NANDN U17789 ( .A(n16839), .B(n16838), .Z(n16840) );
  NAND U17790 ( .A(n16841), .B(n16840), .Z(n17053) );
  NANDN U17791 ( .A(n16847), .B(n16846), .Z(n16851) );
  NAND U17792 ( .A(n16849), .B(n16848), .Z(n16850) );
  NAND U17793 ( .A(n16851), .B(n16850), .Z(n16991) );
  NANDN U17794 ( .A(n16853), .B(n16852), .Z(n16857) );
  NAND U17795 ( .A(n16855), .B(n16854), .Z(n16856) );
  AND U17796 ( .A(n16857), .B(n16856), .Z(n16992) );
  XNOR U17797 ( .A(n16991), .B(n16992), .Z(n16993) );
  XNOR U17798 ( .A(n1052), .B(a[116]), .Z(n17013) );
  NAND U17799 ( .A(n36925), .B(n17013), .Z(n16860) );
  NANDN U17800 ( .A(n16858), .B(n36926), .Z(n16859) );
  NAND U17801 ( .A(n16860), .B(n16859), .Z(n16975) );
  XNOR U17802 ( .A(b[15]), .B(a[110]), .Z(n17016) );
  OR U17803 ( .A(n17016), .B(n37665), .Z(n16863) );
  NANDN U17804 ( .A(n16861), .B(n37604), .Z(n16862) );
  AND U17805 ( .A(n16863), .B(n16862), .Z(n16973) );
  XNOR U17806 ( .A(b[21]), .B(a[104]), .Z(n17019) );
  NANDN U17807 ( .A(n17019), .B(n38101), .Z(n16866) );
  NANDN U17808 ( .A(n16864), .B(n38102), .Z(n16865) );
  AND U17809 ( .A(n16866), .B(n16865), .Z(n16974) );
  XOR U17810 ( .A(n16975), .B(n16976), .Z(n16964) );
  XNOR U17811 ( .A(b[11]), .B(a[114]), .Z(n17022) );
  OR U17812 ( .A(n17022), .B(n37311), .Z(n16869) );
  NANDN U17813 ( .A(n16867), .B(n37218), .Z(n16868) );
  NAND U17814 ( .A(n16869), .B(n16868), .Z(n16962) );
  XNOR U17815 ( .A(b[13]), .B(a[112]), .Z(n17025) );
  NANDN U17816 ( .A(n17025), .B(n37424), .Z(n16872) );
  NANDN U17817 ( .A(n16870), .B(n37425), .Z(n16871) );
  AND U17818 ( .A(n16872), .B(n16871), .Z(n16961) );
  XNOR U17819 ( .A(n16962), .B(n16961), .Z(n16963) );
  XOR U17820 ( .A(n16964), .B(n16963), .Z(n16981) );
  NANDN U17821 ( .A(n1049), .B(a[124]), .Z(n16873) );
  XNOR U17822 ( .A(b[1]), .B(n16873), .Z(n16875) );
  NANDN U17823 ( .A(b[0]), .B(a[123]), .Z(n16874) );
  AND U17824 ( .A(n16875), .B(n16874), .Z(n16939) );
  NAND U17825 ( .A(n38490), .B(n16876), .Z(n16878) );
  XNOR U17826 ( .A(b[29]), .B(a[96]), .Z(n17032) );
  OR U17827 ( .A(n17032), .B(n1048), .Z(n16877) );
  NAND U17828 ( .A(n16878), .B(n16877), .Z(n16937) );
  NANDN U17829 ( .A(n1059), .B(a[92]), .Z(n16938) );
  XNOR U17830 ( .A(n16937), .B(n16938), .Z(n16940) );
  XOR U17831 ( .A(n16939), .B(n16940), .Z(n16979) );
  NANDN U17832 ( .A(n16879), .B(n38205), .Z(n16881) );
  XNOR U17833 ( .A(b[23]), .B(a[102]), .Z(n17035) );
  OR U17834 ( .A(n17035), .B(n38268), .Z(n16880) );
  NAND U17835 ( .A(n16881), .B(n16880), .Z(n17004) );
  XNOR U17836 ( .A(b[7]), .B(a[118]), .Z(n17038) );
  NANDN U17837 ( .A(n17038), .B(n36701), .Z(n16884) );
  NAND U17838 ( .A(n16882), .B(n36702), .Z(n16883) );
  NAND U17839 ( .A(n16884), .B(n16883), .Z(n17001) );
  XOR U17840 ( .A(b[25]), .B(a[100]), .Z(n17041) );
  NAND U17841 ( .A(n17041), .B(n38325), .Z(n16887) );
  NANDN U17842 ( .A(n16885), .B(n38326), .Z(n16886) );
  AND U17843 ( .A(n16887), .B(n16886), .Z(n17002) );
  XNOR U17844 ( .A(n17001), .B(n17002), .Z(n17003) );
  XNOR U17845 ( .A(n17004), .B(n17003), .Z(n16980) );
  XOR U17846 ( .A(n16979), .B(n16980), .Z(n16982) );
  XNOR U17847 ( .A(n16981), .B(n16982), .Z(n16994) );
  XOR U17848 ( .A(n16993), .B(n16994), .Z(n17051) );
  XNOR U17849 ( .A(n17050), .B(n17051), .Z(n17052) );
  XOR U17850 ( .A(n17053), .B(n17052), .Z(n16928) );
  XNOR U17851 ( .A(n16927), .B(n16928), .Z(n16929) );
  XNOR U17852 ( .A(n16930), .B(n16929), .Z(n16934) );
  NANDN U17853 ( .A(n16889), .B(n16888), .Z(n16893) );
  NAND U17854 ( .A(n16891), .B(n16890), .Z(n16892) );
  NAND U17855 ( .A(n16893), .B(n16892), .Z(n16931) );
  NANDN U17856 ( .A(n16895), .B(n16894), .Z(n16899) );
  NAND U17857 ( .A(n16897), .B(n16896), .Z(n16898) );
  NAND U17858 ( .A(n16899), .B(n16898), .Z(n16932) );
  XNOR U17859 ( .A(n16931), .B(n16932), .Z(n16933) );
  XNOR U17860 ( .A(n16934), .B(n16933), .Z(n16924) );
  NANDN U17861 ( .A(n16901), .B(n16900), .Z(n16905) );
  NANDN U17862 ( .A(n16903), .B(n16902), .Z(n16904) );
  NAND U17863 ( .A(n16905), .B(n16904), .Z(n16922) );
  OR U17864 ( .A(n16907), .B(n16906), .Z(n16911) );
  OR U17865 ( .A(n16909), .B(n16908), .Z(n16910) );
  AND U17866 ( .A(n16911), .B(n16910), .Z(n16921) );
  XNOR U17867 ( .A(n16922), .B(n16921), .Z(n16923) );
  XNOR U17868 ( .A(n16924), .B(n16923), .Z(n16917) );
  XOR U17869 ( .A(n16918), .B(n16917), .Z(n16919) );
  XNOR U17870 ( .A(n16920), .B(n16919), .Z(n17056) );
  XNOR U17871 ( .A(n17056), .B(sreg[348]), .Z(n17058) );
  NAND U17872 ( .A(n16912), .B(sreg[347]), .Z(n16916) );
  OR U17873 ( .A(n16914), .B(n16913), .Z(n16915) );
  AND U17874 ( .A(n16916), .B(n16915), .Z(n17057) );
  XOR U17875 ( .A(n17058), .B(n17057), .Z(c[348]) );
  NANDN U17876 ( .A(n16922), .B(n16921), .Z(n16926) );
  NANDN U17877 ( .A(n16924), .B(n16923), .Z(n16925) );
  NAND U17878 ( .A(n16926), .B(n16925), .Z(n17062) );
  NANDN U17879 ( .A(n16932), .B(n16931), .Z(n16936) );
  NANDN U17880 ( .A(n16934), .B(n16933), .Z(n16935) );
  NAND U17881 ( .A(n16936), .B(n16935), .Z(n17068) );
  XNOR U17882 ( .A(n17067), .B(n17068), .Z(n17069) );
  NANDN U17883 ( .A(n16938), .B(n16937), .Z(n16942) );
  NAND U17884 ( .A(n16940), .B(n16939), .Z(n16941) );
  NAND U17885 ( .A(n16942), .B(n16941), .Z(n17130) );
  XOR U17886 ( .A(b[19]), .B(n18980), .Z(n17097) );
  NANDN U17887 ( .A(n17097), .B(n37934), .Z(n16945) );
  NANDN U17888 ( .A(n16943), .B(n37935), .Z(n16944) );
  NAND U17889 ( .A(n16945), .B(n16944), .Z(n17142) );
  XNOR U17890 ( .A(b[27]), .B(a[99]), .Z(n17100) );
  NANDN U17891 ( .A(n17100), .B(n38423), .Z(n16948) );
  NAND U17892 ( .A(n16946), .B(n38424), .Z(n16947) );
  NAND U17893 ( .A(n16948), .B(n16947), .Z(n17139) );
  XNOR U17894 ( .A(b[5]), .B(a[121]), .Z(n17103) );
  NANDN U17895 ( .A(n17103), .B(n36587), .Z(n16951) );
  NANDN U17896 ( .A(n16949), .B(n36588), .Z(n16950) );
  AND U17897 ( .A(n16951), .B(n16950), .Z(n17140) );
  XNOR U17898 ( .A(n17139), .B(n17140), .Z(n17141) );
  XNOR U17899 ( .A(n17142), .B(n17141), .Z(n17127) );
  XNOR U17900 ( .A(b[17]), .B(a[109]), .Z(n17106) );
  NANDN U17901 ( .A(n17106), .B(n37764), .Z(n16954) );
  NAND U17902 ( .A(n16952), .B(n37762), .Z(n16953) );
  NAND U17903 ( .A(n16954), .B(n16953), .Z(n17085) );
  XNOR U17904 ( .A(b[31]), .B(a[95]), .Z(n17109) );
  NANDN U17905 ( .A(n17109), .B(n38552), .Z(n16957) );
  NAND U17906 ( .A(n38553), .B(n16955), .Z(n16956) );
  NAND U17907 ( .A(n16957), .B(n16956), .Z(n17083) );
  OR U17908 ( .A(n16958), .B(n36105), .Z(n16960) );
  XNOR U17909 ( .A(b[3]), .B(a[123]), .Z(n17112) );
  NANDN U17910 ( .A(n17112), .B(n36107), .Z(n16959) );
  AND U17911 ( .A(n16960), .B(n16959), .Z(n17084) );
  XNOR U17912 ( .A(n17083), .B(n17084), .Z(n17086) );
  XNOR U17913 ( .A(n17085), .B(n17086), .Z(n17128) );
  XOR U17914 ( .A(n17127), .B(n17128), .Z(n17129) );
  XNOR U17915 ( .A(n17130), .B(n17129), .Z(n17175) );
  NANDN U17916 ( .A(n16962), .B(n16961), .Z(n16966) );
  NAND U17917 ( .A(n16964), .B(n16963), .Z(n16965) );
  NAND U17918 ( .A(n16966), .B(n16965), .Z(n17118) );
  NANDN U17919 ( .A(n16968), .B(n16967), .Z(n16972) );
  NAND U17920 ( .A(n16970), .B(n16969), .Z(n16971) );
  NAND U17921 ( .A(n16972), .B(n16971), .Z(n17116) );
  OR U17922 ( .A(n16974), .B(n16973), .Z(n16978) );
  NANDN U17923 ( .A(n16976), .B(n16975), .Z(n16977) );
  NAND U17924 ( .A(n16978), .B(n16977), .Z(n17115) );
  XNOR U17925 ( .A(n17118), .B(n17117), .Z(n17176) );
  XOR U17926 ( .A(n17175), .B(n17176), .Z(n17178) );
  NANDN U17927 ( .A(n16980), .B(n16979), .Z(n16984) );
  OR U17928 ( .A(n16982), .B(n16981), .Z(n16983) );
  NAND U17929 ( .A(n16984), .B(n16983), .Z(n17177) );
  XOR U17930 ( .A(n17178), .B(n17177), .Z(n17195) );
  OR U17931 ( .A(n16986), .B(n16985), .Z(n16990) );
  NAND U17932 ( .A(n16988), .B(n16987), .Z(n16989) );
  NAND U17933 ( .A(n16990), .B(n16989), .Z(n17194) );
  NANDN U17934 ( .A(n16992), .B(n16991), .Z(n16996) );
  NANDN U17935 ( .A(n16994), .B(n16993), .Z(n16995) );
  NAND U17936 ( .A(n16996), .B(n16995), .Z(n17183) );
  NANDN U17937 ( .A(n17002), .B(n17001), .Z(n17006) );
  NAND U17938 ( .A(n17004), .B(n17003), .Z(n17005) );
  NAND U17939 ( .A(n17006), .B(n17005), .Z(n17121) );
  NANDN U17940 ( .A(n17008), .B(n17007), .Z(n17012) );
  NAND U17941 ( .A(n17010), .B(n17009), .Z(n17011) );
  AND U17942 ( .A(n17012), .B(n17011), .Z(n17122) );
  XNOR U17943 ( .A(n17121), .B(n17122), .Z(n17123) );
  XNOR U17944 ( .A(b[9]), .B(a[117]), .Z(n17145) );
  NANDN U17945 ( .A(n17145), .B(n36925), .Z(n17015) );
  NAND U17946 ( .A(n36926), .B(n17013), .Z(n17014) );
  NAND U17947 ( .A(n17015), .B(n17014), .Z(n17089) );
  XNOR U17948 ( .A(n1054), .B(a[111]), .Z(n17148) );
  NANDN U17949 ( .A(n37665), .B(n17148), .Z(n17018) );
  NANDN U17950 ( .A(n17016), .B(n37604), .Z(n17017) );
  NAND U17951 ( .A(n17018), .B(n17017), .Z(n17087) );
  XNOR U17952 ( .A(b[21]), .B(a[105]), .Z(n17151) );
  NANDN U17953 ( .A(n17151), .B(n38101), .Z(n17021) );
  NANDN U17954 ( .A(n17019), .B(n38102), .Z(n17020) );
  AND U17955 ( .A(n17021), .B(n17020), .Z(n17088) );
  XNOR U17956 ( .A(n17087), .B(n17088), .Z(n17090) );
  XOR U17957 ( .A(n17089), .B(n17090), .Z(n17082) );
  XNOR U17958 ( .A(b[11]), .B(a[115]), .Z(n17154) );
  OR U17959 ( .A(n17154), .B(n37311), .Z(n17024) );
  NANDN U17960 ( .A(n17022), .B(n37218), .Z(n17023) );
  NAND U17961 ( .A(n17024), .B(n17023), .Z(n17080) );
  XOR U17962 ( .A(n1053), .B(n19909), .Z(n17157) );
  NAND U17963 ( .A(n17157), .B(n37424), .Z(n17027) );
  NANDN U17964 ( .A(n17025), .B(n37425), .Z(n17026) );
  AND U17965 ( .A(n17027), .B(n17026), .Z(n17079) );
  XNOR U17966 ( .A(n17080), .B(n17079), .Z(n17081) );
  XNOR U17967 ( .A(n17082), .B(n17081), .Z(n17075) );
  NANDN U17968 ( .A(n1049), .B(a[125]), .Z(n17028) );
  XNOR U17969 ( .A(b[1]), .B(n17028), .Z(n17030) );
  NANDN U17970 ( .A(b[0]), .B(a[124]), .Z(n17029) );
  AND U17971 ( .A(n17030), .B(n17029), .Z(n17094) );
  ANDN U17972 ( .B(b[31]), .A(n17031), .Z(n17091) );
  NANDN U17973 ( .A(n17032), .B(n38490), .Z(n17034) );
  XNOR U17974 ( .A(n1058), .B(a[97]), .Z(n17160) );
  NANDN U17975 ( .A(n1048), .B(n17160), .Z(n17033) );
  NAND U17976 ( .A(n17034), .B(n17033), .Z(n17092) );
  XOR U17977 ( .A(n17091), .B(n17092), .Z(n17093) );
  XNOR U17978 ( .A(n17094), .B(n17093), .Z(n17073) );
  NANDN U17979 ( .A(n17035), .B(n38205), .Z(n17037) );
  XNOR U17980 ( .A(b[23]), .B(a[103]), .Z(n17166) );
  OR U17981 ( .A(n17166), .B(n38268), .Z(n17036) );
  NAND U17982 ( .A(n17037), .B(n17036), .Z(n17136) );
  XOR U17983 ( .A(b[7]), .B(a[119]), .Z(n17169) );
  NAND U17984 ( .A(n17169), .B(n36701), .Z(n17040) );
  NANDN U17985 ( .A(n17038), .B(n36702), .Z(n17039) );
  NAND U17986 ( .A(n17040), .B(n17039), .Z(n17133) );
  XNOR U17987 ( .A(b[25]), .B(a[101]), .Z(n17172) );
  NANDN U17988 ( .A(n17172), .B(n38325), .Z(n17043) );
  NAND U17989 ( .A(n17041), .B(n38326), .Z(n17042) );
  AND U17990 ( .A(n17043), .B(n17042), .Z(n17134) );
  XNOR U17991 ( .A(n17133), .B(n17134), .Z(n17135) );
  XNOR U17992 ( .A(n17136), .B(n17135), .Z(n17074) );
  XNOR U17993 ( .A(n17073), .B(n17074), .Z(n17076) );
  XOR U17994 ( .A(n17123), .B(n17124), .Z(n17181) );
  XNOR U17995 ( .A(n17182), .B(n17181), .Z(n17184) );
  XNOR U17996 ( .A(n17183), .B(n17184), .Z(n17193) );
  XOR U17997 ( .A(n17194), .B(n17193), .Z(n17196) );
  NANDN U17998 ( .A(n17045), .B(n17044), .Z(n17049) );
  NAND U17999 ( .A(n17047), .B(n17046), .Z(n17048) );
  NAND U18000 ( .A(n17049), .B(n17048), .Z(n17187) );
  NANDN U18001 ( .A(n17051), .B(n17050), .Z(n17055) );
  NAND U18002 ( .A(n17053), .B(n17052), .Z(n17054) );
  NAND U18003 ( .A(n17055), .B(n17054), .Z(n17188) );
  XNOR U18004 ( .A(n17187), .B(n17188), .Z(n17189) );
  XOR U18005 ( .A(n17190), .B(n17189), .Z(n17070) );
  XOR U18006 ( .A(n17069), .B(n17070), .Z(n17061) );
  XOR U18007 ( .A(n17062), .B(n17061), .Z(n17063) );
  XNOR U18008 ( .A(n17064), .B(n17063), .Z(n17199) );
  XNOR U18009 ( .A(n17199), .B(sreg[349]), .Z(n17201) );
  NAND U18010 ( .A(n17056), .B(sreg[348]), .Z(n17060) );
  OR U18011 ( .A(n17058), .B(n17057), .Z(n17059) );
  AND U18012 ( .A(n17060), .B(n17059), .Z(n17200) );
  XOR U18013 ( .A(n17201), .B(n17200), .Z(c[349]) );
  NAND U18014 ( .A(n17062), .B(n17061), .Z(n17066) );
  NAND U18015 ( .A(n17064), .B(n17063), .Z(n17065) );
  NAND U18016 ( .A(n17066), .B(n17065), .Z(n17207) );
  NANDN U18017 ( .A(n17068), .B(n17067), .Z(n17072) );
  NAND U18018 ( .A(n17070), .B(n17069), .Z(n17071) );
  NAND U18019 ( .A(n17072), .B(n17071), .Z(n17205) );
  OR U18020 ( .A(n17074), .B(n17073), .Z(n17078) );
  OR U18021 ( .A(n17076), .B(n17075), .Z(n17077) );
  NAND U18022 ( .A(n17078), .B(n17077), .Z(n17223) );
  XNOR U18023 ( .A(n17275), .B(n17274), .Z(n17277) );
  XNOR U18024 ( .A(n17276), .B(n17277), .Z(n17221) );
  OR U18025 ( .A(n17092), .B(n17091), .Z(n17096) );
  NANDN U18026 ( .A(n17094), .B(n17093), .Z(n17095) );
  NAND U18027 ( .A(n17096), .B(n17095), .Z(n17286) );
  XNOR U18028 ( .A(b[19]), .B(a[108]), .Z(n17232) );
  NANDN U18029 ( .A(n17232), .B(n37934), .Z(n17099) );
  NANDN U18030 ( .A(n17097), .B(n37935), .Z(n17098) );
  NAND U18031 ( .A(n17099), .B(n17098), .Z(n17299) );
  XOR U18032 ( .A(b[27]), .B(a[100]), .Z(n17235) );
  NAND U18033 ( .A(n38423), .B(n17235), .Z(n17102) );
  NANDN U18034 ( .A(n17100), .B(n38424), .Z(n17101) );
  NAND U18035 ( .A(n17102), .B(n17101), .Z(n17296) );
  XNOR U18036 ( .A(b[5]), .B(a[122]), .Z(n17238) );
  NANDN U18037 ( .A(n17238), .B(n36587), .Z(n17105) );
  NANDN U18038 ( .A(n17103), .B(n36588), .Z(n17104) );
  AND U18039 ( .A(n17105), .B(n17104), .Z(n17297) );
  XNOR U18040 ( .A(n17296), .B(n17297), .Z(n17298) );
  XNOR U18041 ( .A(n17299), .B(n17298), .Z(n17285) );
  NANDN U18042 ( .A(n17106), .B(n37762), .Z(n17108) );
  XOR U18043 ( .A(b[17]), .B(a[110]), .Z(n17241) );
  NAND U18044 ( .A(n17241), .B(n37764), .Z(n17107) );
  NAND U18045 ( .A(n17108), .B(n17107), .Z(n17259) );
  XNOR U18046 ( .A(b[31]), .B(a[96]), .Z(n17244) );
  NANDN U18047 ( .A(n17244), .B(n38552), .Z(n17111) );
  NANDN U18048 ( .A(n17109), .B(n38553), .Z(n17110) );
  NAND U18049 ( .A(n17111), .B(n17110), .Z(n17256) );
  OR U18050 ( .A(n17112), .B(n36105), .Z(n17114) );
  XNOR U18051 ( .A(b[3]), .B(a[124]), .Z(n17247) );
  NANDN U18052 ( .A(n17247), .B(n36107), .Z(n17113) );
  AND U18053 ( .A(n17114), .B(n17113), .Z(n17257) );
  XNOR U18054 ( .A(n17256), .B(n17257), .Z(n17258) );
  XOR U18055 ( .A(n17259), .B(n17258), .Z(n17284) );
  XOR U18056 ( .A(n17285), .B(n17284), .Z(n17287) );
  XOR U18057 ( .A(n17286), .B(n17287), .Z(n17220) );
  XNOR U18058 ( .A(n17221), .B(n17220), .Z(n17222) );
  XNOR U18059 ( .A(n17223), .B(n17222), .Z(n17341) );
  OR U18060 ( .A(n17116), .B(n17115), .Z(n17120) );
  NAND U18061 ( .A(n17118), .B(n17117), .Z(n17119) );
  NAND U18062 ( .A(n17120), .B(n17119), .Z(n17339) );
  NANDN U18063 ( .A(n17122), .B(n17121), .Z(n17126) );
  NAND U18064 ( .A(n17124), .B(n17123), .Z(n17125) );
  NAND U18065 ( .A(n17126), .B(n17125), .Z(n17216) );
  OR U18066 ( .A(n17128), .B(n17127), .Z(n17132) );
  NAND U18067 ( .A(n17130), .B(n17129), .Z(n17131) );
  NAND U18068 ( .A(n17132), .B(n17131), .Z(n17215) );
  NANDN U18069 ( .A(n17134), .B(n17133), .Z(n17138) );
  NAND U18070 ( .A(n17136), .B(n17135), .Z(n17137) );
  NAND U18071 ( .A(n17138), .B(n17137), .Z(n17278) );
  NANDN U18072 ( .A(n17140), .B(n17139), .Z(n17144) );
  NAND U18073 ( .A(n17142), .B(n17141), .Z(n17143) );
  AND U18074 ( .A(n17144), .B(n17143), .Z(n17279) );
  XNOR U18075 ( .A(n17278), .B(n17279), .Z(n17280) );
  XOR U18076 ( .A(b[9]), .B(n20271), .Z(n17302) );
  NANDN U18077 ( .A(n17302), .B(n36925), .Z(n17147) );
  NANDN U18078 ( .A(n17145), .B(n36926), .Z(n17146) );
  NAND U18079 ( .A(n17147), .B(n17146), .Z(n17270) );
  XNOR U18080 ( .A(b[15]), .B(a[112]), .Z(n17305) );
  OR U18081 ( .A(n17305), .B(n37665), .Z(n17150) );
  NAND U18082 ( .A(n17148), .B(n37604), .Z(n17149) );
  AND U18083 ( .A(n17150), .B(n17149), .Z(n17268) );
  XNOR U18084 ( .A(b[21]), .B(a[106]), .Z(n17308) );
  NANDN U18085 ( .A(n17308), .B(n38101), .Z(n17153) );
  NANDN U18086 ( .A(n17151), .B(n38102), .Z(n17152) );
  AND U18087 ( .A(n17153), .B(n17152), .Z(n17269) );
  XOR U18088 ( .A(n17270), .B(n17271), .Z(n17265) );
  XNOR U18089 ( .A(b[11]), .B(a[116]), .Z(n17311) );
  OR U18090 ( .A(n17311), .B(n37311), .Z(n17156) );
  NANDN U18091 ( .A(n17154), .B(n37218), .Z(n17155) );
  NAND U18092 ( .A(n17156), .B(n17155), .Z(n17263) );
  XOR U18093 ( .A(n1053), .B(a[114]), .Z(n17314) );
  NANDN U18094 ( .A(n17314), .B(n37424), .Z(n17159) );
  NAND U18095 ( .A(n37425), .B(n17157), .Z(n17158) );
  AND U18096 ( .A(n17159), .B(n17158), .Z(n17262) );
  XNOR U18097 ( .A(n17263), .B(n17262), .Z(n17264) );
  XOR U18098 ( .A(n17265), .B(n17264), .Z(n17252) );
  NAND U18099 ( .A(n17160), .B(n38490), .Z(n17162) );
  XNOR U18100 ( .A(n1058), .B(a[98]), .Z(n17320) );
  NANDN U18101 ( .A(n1048), .B(n17320), .Z(n17161) );
  NAND U18102 ( .A(n17162), .B(n17161), .Z(n17226) );
  NANDN U18103 ( .A(n1059), .B(a[94]), .Z(n17227) );
  XNOR U18104 ( .A(n17226), .B(n17227), .Z(n17229) );
  NANDN U18105 ( .A(n1049), .B(a[126]), .Z(n17163) );
  XNOR U18106 ( .A(b[1]), .B(n17163), .Z(n17165) );
  NANDN U18107 ( .A(b[0]), .B(a[125]), .Z(n17164) );
  AND U18108 ( .A(n17165), .B(n17164), .Z(n17228) );
  XOR U18109 ( .A(n17229), .B(n17228), .Z(n17250) );
  NANDN U18110 ( .A(n17166), .B(n38205), .Z(n17168) );
  XNOR U18111 ( .A(b[23]), .B(a[104]), .Z(n17323) );
  OR U18112 ( .A(n17323), .B(n38268), .Z(n17167) );
  NAND U18113 ( .A(n17168), .B(n17167), .Z(n17293) );
  XOR U18114 ( .A(b[7]), .B(a[120]), .Z(n17326) );
  NAND U18115 ( .A(n17326), .B(n36701), .Z(n17171) );
  NAND U18116 ( .A(n17169), .B(n36702), .Z(n17170) );
  NAND U18117 ( .A(n17171), .B(n17170), .Z(n17290) );
  XOR U18118 ( .A(b[25]), .B(a[102]), .Z(n17329) );
  NAND U18119 ( .A(n17329), .B(n38325), .Z(n17174) );
  NANDN U18120 ( .A(n17172), .B(n38326), .Z(n17173) );
  AND U18121 ( .A(n17174), .B(n17173), .Z(n17291) );
  XNOR U18122 ( .A(n17290), .B(n17291), .Z(n17292) );
  XNOR U18123 ( .A(n17293), .B(n17292), .Z(n17251) );
  XOR U18124 ( .A(n17250), .B(n17251), .Z(n17253) );
  XNOR U18125 ( .A(n17252), .B(n17253), .Z(n17281) );
  XNOR U18126 ( .A(n17280), .B(n17281), .Z(n17214) );
  XNOR U18127 ( .A(n17215), .B(n17214), .Z(n17217) );
  XNOR U18128 ( .A(n17216), .B(n17217), .Z(n17338) );
  XNOR U18129 ( .A(n17339), .B(n17338), .Z(n17340) );
  XOR U18130 ( .A(n17341), .B(n17340), .Z(n17335) );
  NANDN U18131 ( .A(n17176), .B(n17175), .Z(n17180) );
  OR U18132 ( .A(n17178), .B(n17177), .Z(n17179) );
  NAND U18133 ( .A(n17180), .B(n17179), .Z(n17332) );
  NAND U18134 ( .A(n17182), .B(n17181), .Z(n17186) );
  NANDN U18135 ( .A(n17184), .B(n17183), .Z(n17185) );
  NAND U18136 ( .A(n17186), .B(n17185), .Z(n17333) );
  XNOR U18137 ( .A(n17332), .B(n17333), .Z(n17334) );
  XNOR U18138 ( .A(n17335), .B(n17334), .Z(n17211) );
  NANDN U18139 ( .A(n17188), .B(n17187), .Z(n17192) );
  NAND U18140 ( .A(n17190), .B(n17189), .Z(n17191) );
  NAND U18141 ( .A(n17192), .B(n17191), .Z(n17208) );
  NANDN U18142 ( .A(n17194), .B(n17193), .Z(n17198) );
  OR U18143 ( .A(n17196), .B(n17195), .Z(n17197) );
  NAND U18144 ( .A(n17198), .B(n17197), .Z(n17209) );
  XNOR U18145 ( .A(n17208), .B(n17209), .Z(n17210) );
  XNOR U18146 ( .A(n17211), .B(n17210), .Z(n17204) );
  XOR U18147 ( .A(n17205), .B(n17204), .Z(n17206) );
  XNOR U18148 ( .A(n17207), .B(n17206), .Z(n17344) );
  XNOR U18149 ( .A(n17344), .B(sreg[350]), .Z(n17346) );
  NAND U18150 ( .A(n17199), .B(sreg[349]), .Z(n17203) );
  OR U18151 ( .A(n17201), .B(n17200), .Z(n17202) );
  AND U18152 ( .A(n17203), .B(n17202), .Z(n17345) );
  XOR U18153 ( .A(n17346), .B(n17345), .Z(c[350]) );
  NANDN U18154 ( .A(n17209), .B(n17208), .Z(n17213) );
  NANDN U18155 ( .A(n17211), .B(n17210), .Z(n17212) );
  NAND U18156 ( .A(n17213), .B(n17212), .Z(n17349) );
  NAND U18157 ( .A(n17215), .B(n17214), .Z(n17219) );
  NANDN U18158 ( .A(n17217), .B(n17216), .Z(n17218) );
  NAND U18159 ( .A(n17219), .B(n17218), .Z(n17481) );
  NANDN U18160 ( .A(n17221), .B(n17220), .Z(n17225) );
  NAND U18161 ( .A(n17223), .B(n17222), .Z(n17224) );
  AND U18162 ( .A(n17225), .B(n17224), .Z(n17482) );
  XNOR U18163 ( .A(n17481), .B(n17482), .Z(n17483) );
  NANDN U18164 ( .A(n17227), .B(n17226), .Z(n17231) );
  NAND U18165 ( .A(n17229), .B(n17228), .Z(n17230) );
  NAND U18166 ( .A(n17231), .B(n17230), .Z(n17436) );
  XNOR U18167 ( .A(b[19]), .B(a[109]), .Z(n17403) );
  NANDN U18168 ( .A(n17403), .B(n37934), .Z(n17234) );
  NANDN U18169 ( .A(n17232), .B(n37935), .Z(n17233) );
  NAND U18170 ( .A(n17234), .B(n17233), .Z(n17448) );
  XNOR U18171 ( .A(b[27]), .B(a[101]), .Z(n17406) );
  NANDN U18172 ( .A(n17406), .B(n38423), .Z(n17237) );
  NAND U18173 ( .A(n17235), .B(n38424), .Z(n17236) );
  NAND U18174 ( .A(n17237), .B(n17236), .Z(n17445) );
  XNOR U18175 ( .A(b[5]), .B(a[123]), .Z(n17409) );
  NANDN U18176 ( .A(n17409), .B(n36587), .Z(n17240) );
  NANDN U18177 ( .A(n17238), .B(n36588), .Z(n17239) );
  AND U18178 ( .A(n17240), .B(n17239), .Z(n17446) );
  XNOR U18179 ( .A(n17445), .B(n17446), .Z(n17447) );
  XNOR U18180 ( .A(n17448), .B(n17447), .Z(n17433) );
  NAND U18181 ( .A(n17241), .B(n37762), .Z(n17243) );
  XOR U18182 ( .A(b[17]), .B(a[111]), .Z(n17412) );
  NAND U18183 ( .A(n17412), .B(n37764), .Z(n17242) );
  NAND U18184 ( .A(n17243), .B(n17242), .Z(n17387) );
  XNOR U18185 ( .A(b[31]), .B(a[97]), .Z(n17415) );
  NANDN U18186 ( .A(n17415), .B(n38552), .Z(n17246) );
  NANDN U18187 ( .A(n17244), .B(n38553), .Z(n17245) );
  AND U18188 ( .A(n17246), .B(n17245), .Z(n17385) );
  OR U18189 ( .A(n17247), .B(n36105), .Z(n17249) );
  XNOR U18190 ( .A(b[3]), .B(a[125]), .Z(n17418) );
  NANDN U18191 ( .A(n17418), .B(n36107), .Z(n17248) );
  AND U18192 ( .A(n17249), .B(n17248), .Z(n17386) );
  XOR U18193 ( .A(n17387), .B(n17388), .Z(n17434) );
  XOR U18194 ( .A(n17433), .B(n17434), .Z(n17435) );
  XNOR U18195 ( .A(n17436), .B(n17435), .Z(n17361) );
  NANDN U18196 ( .A(n17251), .B(n17250), .Z(n17255) );
  OR U18197 ( .A(n17253), .B(n17252), .Z(n17254) );
  NAND U18198 ( .A(n17255), .B(n17254), .Z(n17362) );
  XNOR U18199 ( .A(n17361), .B(n17362), .Z(n17363) );
  NANDN U18200 ( .A(n17257), .B(n17256), .Z(n17261) );
  NAND U18201 ( .A(n17259), .B(n17258), .Z(n17260) );
  NAND U18202 ( .A(n17261), .B(n17260), .Z(n17424) );
  NANDN U18203 ( .A(n17263), .B(n17262), .Z(n17267) );
  NAND U18204 ( .A(n17265), .B(n17264), .Z(n17266) );
  NAND U18205 ( .A(n17267), .B(n17266), .Z(n17421) );
  OR U18206 ( .A(n17269), .B(n17268), .Z(n17273) );
  NANDN U18207 ( .A(n17271), .B(n17270), .Z(n17272) );
  NAND U18208 ( .A(n17273), .B(n17272), .Z(n17422) );
  XNOR U18209 ( .A(n17421), .B(n17422), .Z(n17423) );
  XOR U18210 ( .A(n17424), .B(n17423), .Z(n17364) );
  XNOR U18211 ( .A(n17363), .B(n17364), .Z(n17489) );
  NANDN U18212 ( .A(n17279), .B(n17278), .Z(n17283) );
  NANDN U18213 ( .A(n17281), .B(n17280), .Z(n17282) );
  NAND U18214 ( .A(n17283), .B(n17282), .Z(n17370) );
  NANDN U18215 ( .A(n17285), .B(n17284), .Z(n17289) );
  OR U18216 ( .A(n17287), .B(n17286), .Z(n17288) );
  NAND U18217 ( .A(n17289), .B(n17288), .Z(n17368) );
  NANDN U18218 ( .A(n17291), .B(n17290), .Z(n17295) );
  NAND U18219 ( .A(n17293), .B(n17292), .Z(n17294) );
  NAND U18220 ( .A(n17295), .B(n17294), .Z(n17427) );
  NANDN U18221 ( .A(n17297), .B(n17296), .Z(n17301) );
  NAND U18222 ( .A(n17299), .B(n17298), .Z(n17300) );
  AND U18223 ( .A(n17301), .B(n17300), .Z(n17428) );
  XNOR U18224 ( .A(n17427), .B(n17428), .Z(n17429) );
  XNOR U18225 ( .A(n1052), .B(a[119]), .Z(n17457) );
  NAND U18226 ( .A(n36925), .B(n17457), .Z(n17304) );
  NANDN U18227 ( .A(n17302), .B(n36926), .Z(n17303) );
  NAND U18228 ( .A(n17304), .B(n17303), .Z(n17393) );
  XOR U18229 ( .A(b[15]), .B(n19909), .Z(n17454) );
  OR U18230 ( .A(n17454), .B(n37665), .Z(n17307) );
  NANDN U18231 ( .A(n17305), .B(n37604), .Z(n17306) );
  AND U18232 ( .A(n17307), .B(n17306), .Z(n17391) );
  XOR U18233 ( .A(n1056), .B(n18980), .Z(n17451) );
  NAND U18234 ( .A(n17451), .B(n38101), .Z(n17310) );
  NANDN U18235 ( .A(n17308), .B(n38102), .Z(n17309) );
  AND U18236 ( .A(n17310), .B(n17309), .Z(n17392) );
  XOR U18237 ( .A(n17393), .B(n17394), .Z(n17382) );
  XNOR U18238 ( .A(b[11]), .B(a[117]), .Z(n17460) );
  OR U18239 ( .A(n17460), .B(n37311), .Z(n17313) );
  NANDN U18240 ( .A(n17311), .B(n37218), .Z(n17312) );
  NAND U18241 ( .A(n17313), .B(n17312), .Z(n17380) );
  XOR U18242 ( .A(n1053), .B(a[115]), .Z(n17463) );
  NANDN U18243 ( .A(n17463), .B(n37424), .Z(n17316) );
  NANDN U18244 ( .A(n17314), .B(n37425), .Z(n17315) );
  NAND U18245 ( .A(n17316), .B(n17315), .Z(n17379) );
  XOR U18246 ( .A(n17382), .B(n17381), .Z(n17376) );
  NANDN U18247 ( .A(n1049), .B(a[127]), .Z(n17317) );
  XNOR U18248 ( .A(b[1]), .B(n17317), .Z(n17319) );
  NANDN U18249 ( .A(b[0]), .B(a[126]), .Z(n17318) );
  AND U18250 ( .A(n17319), .B(n17318), .Z(n17399) );
  NAND U18251 ( .A(n38490), .B(n17320), .Z(n17322) );
  XOR U18252 ( .A(n1058), .B(n17884), .Z(n17469) );
  NANDN U18253 ( .A(n1048), .B(n17469), .Z(n17321) );
  NAND U18254 ( .A(n17322), .B(n17321), .Z(n17397) );
  NANDN U18255 ( .A(n1059), .B(a[95]), .Z(n17398) );
  XNOR U18256 ( .A(n17397), .B(n17398), .Z(n17400) );
  XNOR U18257 ( .A(n17399), .B(n17400), .Z(n17374) );
  NANDN U18258 ( .A(n17323), .B(n38205), .Z(n17325) );
  XNOR U18259 ( .A(b[23]), .B(a[105]), .Z(n17472) );
  OR U18260 ( .A(n17472), .B(n38268), .Z(n17324) );
  NAND U18261 ( .A(n17325), .B(n17324), .Z(n17442) );
  XOR U18262 ( .A(b[7]), .B(a[121]), .Z(n17475) );
  NAND U18263 ( .A(n17475), .B(n36701), .Z(n17328) );
  NAND U18264 ( .A(n17326), .B(n36702), .Z(n17327) );
  NAND U18265 ( .A(n17328), .B(n17327), .Z(n17439) );
  XOR U18266 ( .A(b[25]), .B(a[103]), .Z(n17478) );
  NAND U18267 ( .A(n17478), .B(n38325), .Z(n17331) );
  NAND U18268 ( .A(n17329), .B(n38326), .Z(n17330) );
  AND U18269 ( .A(n17331), .B(n17330), .Z(n17440) );
  XNOR U18270 ( .A(n17439), .B(n17440), .Z(n17441) );
  XOR U18271 ( .A(n17442), .B(n17441), .Z(n17373) );
  XOR U18272 ( .A(n17376), .B(n17375), .Z(n17430) );
  XNOR U18273 ( .A(n17429), .B(n17430), .Z(n17367) );
  XOR U18274 ( .A(n17368), .B(n17367), .Z(n17369) );
  XNOR U18275 ( .A(n17370), .B(n17369), .Z(n17487) );
  XNOR U18276 ( .A(n17488), .B(n17487), .Z(n17490) );
  XNOR U18277 ( .A(n17489), .B(n17490), .Z(n17484) );
  XOR U18278 ( .A(n17483), .B(n17484), .Z(n17358) );
  NANDN U18279 ( .A(n17333), .B(n17332), .Z(n17337) );
  NAND U18280 ( .A(n17335), .B(n17334), .Z(n17336) );
  NAND U18281 ( .A(n17337), .B(n17336), .Z(n17355) );
  NANDN U18282 ( .A(n17339), .B(n17338), .Z(n17343) );
  NANDN U18283 ( .A(n17341), .B(n17340), .Z(n17342) );
  NAND U18284 ( .A(n17343), .B(n17342), .Z(n17356) );
  XNOR U18285 ( .A(n17355), .B(n17356), .Z(n17357) );
  XNOR U18286 ( .A(n17358), .B(n17357), .Z(n17350) );
  XNOR U18287 ( .A(n17349), .B(n17350), .Z(n17351) );
  XNOR U18288 ( .A(n17352), .B(n17351), .Z(n17493) );
  XNOR U18289 ( .A(n17493), .B(sreg[351]), .Z(n17495) );
  NAND U18290 ( .A(n17344), .B(sreg[350]), .Z(n17348) );
  OR U18291 ( .A(n17346), .B(n17345), .Z(n17347) );
  AND U18292 ( .A(n17348), .B(n17347), .Z(n17494) );
  XOR U18293 ( .A(n17495), .B(n17494), .Z(c[351]) );
  NANDN U18294 ( .A(n17350), .B(n17349), .Z(n17354) );
  NAND U18295 ( .A(n17352), .B(n17351), .Z(n17353) );
  NAND U18296 ( .A(n17354), .B(n17353), .Z(n17501) );
  NANDN U18297 ( .A(n17356), .B(n17355), .Z(n17360) );
  NAND U18298 ( .A(n17358), .B(n17357), .Z(n17359) );
  NAND U18299 ( .A(n17360), .B(n17359), .Z(n17499) );
  NANDN U18300 ( .A(n17362), .B(n17361), .Z(n17366) );
  NANDN U18301 ( .A(n17364), .B(n17363), .Z(n17365) );
  NAND U18302 ( .A(n17366), .B(n17365), .Z(n17632) );
  NAND U18303 ( .A(n17368), .B(n17367), .Z(n17372) );
  NAND U18304 ( .A(n17370), .B(n17369), .Z(n17371) );
  NAND U18305 ( .A(n17372), .B(n17371), .Z(n17633) );
  XNOR U18306 ( .A(n17632), .B(n17633), .Z(n17634) );
  NANDN U18307 ( .A(n17374), .B(n17373), .Z(n17378) );
  NANDN U18308 ( .A(n17376), .B(n17375), .Z(n17377) );
  NAND U18309 ( .A(n17378), .B(n17377), .Z(n17619) );
  OR U18310 ( .A(n17380), .B(n17379), .Z(n17384) );
  NAND U18311 ( .A(n17382), .B(n17381), .Z(n17383) );
  NAND U18312 ( .A(n17384), .B(n17383), .Z(n17558) );
  OR U18313 ( .A(n17386), .B(n17385), .Z(n17390) );
  NANDN U18314 ( .A(n17388), .B(n17387), .Z(n17389) );
  NAND U18315 ( .A(n17390), .B(n17389), .Z(n17557) );
  OR U18316 ( .A(n17392), .B(n17391), .Z(n17396) );
  NANDN U18317 ( .A(n17394), .B(n17393), .Z(n17395) );
  NAND U18318 ( .A(n17396), .B(n17395), .Z(n17556) );
  XOR U18319 ( .A(n17558), .B(n17559), .Z(n17616) );
  NANDN U18320 ( .A(n17398), .B(n17397), .Z(n17402) );
  NAND U18321 ( .A(n17400), .B(n17399), .Z(n17401) );
  NAND U18322 ( .A(n17402), .B(n17401), .Z(n17571) );
  XNOR U18323 ( .A(b[19]), .B(a[110]), .Z(n17516) );
  NANDN U18324 ( .A(n17516), .B(n37934), .Z(n17405) );
  NANDN U18325 ( .A(n17403), .B(n37935), .Z(n17404) );
  NAND U18326 ( .A(n17405), .B(n17404), .Z(n17583) );
  XOR U18327 ( .A(b[27]), .B(a[102]), .Z(n17519) );
  NAND U18328 ( .A(n38423), .B(n17519), .Z(n17408) );
  NANDN U18329 ( .A(n17406), .B(n38424), .Z(n17407) );
  NAND U18330 ( .A(n17408), .B(n17407), .Z(n17580) );
  XNOR U18331 ( .A(b[5]), .B(a[124]), .Z(n17522) );
  NANDN U18332 ( .A(n17522), .B(n36587), .Z(n17411) );
  NANDN U18333 ( .A(n17409), .B(n36588), .Z(n17410) );
  AND U18334 ( .A(n17411), .B(n17410), .Z(n17581) );
  XNOR U18335 ( .A(n17580), .B(n17581), .Z(n17582) );
  XNOR U18336 ( .A(n17583), .B(n17582), .Z(n17569) );
  NAND U18337 ( .A(n17412), .B(n37762), .Z(n17414) );
  XOR U18338 ( .A(b[17]), .B(a[112]), .Z(n17525) );
  NAND U18339 ( .A(n17525), .B(n37764), .Z(n17413) );
  NAND U18340 ( .A(n17414), .B(n17413), .Z(n17543) );
  XNOR U18341 ( .A(b[31]), .B(a[98]), .Z(n17528) );
  NANDN U18342 ( .A(n17528), .B(n38552), .Z(n17417) );
  NANDN U18343 ( .A(n17415), .B(n38553), .Z(n17416) );
  NAND U18344 ( .A(n17417), .B(n17416), .Z(n17540) );
  OR U18345 ( .A(n17418), .B(n36105), .Z(n17420) );
  XNOR U18346 ( .A(b[3]), .B(a[126]), .Z(n17531) );
  NANDN U18347 ( .A(n17531), .B(n36107), .Z(n17419) );
  AND U18348 ( .A(n17420), .B(n17419), .Z(n17541) );
  XNOR U18349 ( .A(n17540), .B(n17541), .Z(n17542) );
  XOR U18350 ( .A(n17543), .B(n17542), .Z(n17568) );
  XNOR U18351 ( .A(n17569), .B(n17568), .Z(n17570) );
  XNOR U18352 ( .A(n17571), .B(n17570), .Z(n17617) );
  XNOR U18353 ( .A(n17616), .B(n17617), .Z(n17618) );
  XNOR U18354 ( .A(n17619), .B(n17618), .Z(n17629) );
  NANDN U18355 ( .A(n17422), .B(n17421), .Z(n17426) );
  NANDN U18356 ( .A(n17424), .B(n17423), .Z(n17425) );
  NAND U18357 ( .A(n17426), .B(n17425), .Z(n17626) );
  NANDN U18358 ( .A(n17428), .B(n17427), .Z(n17432) );
  NANDN U18359 ( .A(n17430), .B(n17429), .Z(n17431) );
  NAND U18360 ( .A(n17432), .B(n17431), .Z(n17623) );
  OR U18361 ( .A(n17434), .B(n17433), .Z(n17438) );
  NAND U18362 ( .A(n17436), .B(n17435), .Z(n17437) );
  NAND U18363 ( .A(n17438), .B(n17437), .Z(n17621) );
  NANDN U18364 ( .A(n17440), .B(n17439), .Z(n17444) );
  NAND U18365 ( .A(n17442), .B(n17441), .Z(n17443) );
  NAND U18366 ( .A(n17444), .B(n17443), .Z(n17562) );
  NANDN U18367 ( .A(n17446), .B(n17445), .Z(n17450) );
  NAND U18368 ( .A(n17448), .B(n17447), .Z(n17449) );
  AND U18369 ( .A(n17450), .B(n17449), .Z(n17563) );
  XNOR U18370 ( .A(n17562), .B(n17563), .Z(n17564) );
  XOR U18371 ( .A(n1056), .B(a[108]), .Z(n17586) );
  NANDN U18372 ( .A(n17586), .B(n38101), .Z(n17453) );
  NAND U18373 ( .A(n38102), .B(n17451), .Z(n17452) );
  NAND U18374 ( .A(n17453), .B(n17452), .Z(n17552) );
  XNOR U18375 ( .A(b[15]), .B(a[114]), .Z(n17589) );
  OR U18376 ( .A(n17589), .B(n37665), .Z(n17456) );
  NANDN U18377 ( .A(n17454), .B(n37604), .Z(n17455) );
  AND U18378 ( .A(n17456), .B(n17455), .Z(n17553) );
  XNOR U18379 ( .A(n17552), .B(n17553), .Z(n17555) );
  XOR U18380 ( .A(n1052), .B(a[120]), .Z(n17592) );
  NANDN U18381 ( .A(n17592), .B(n36925), .Z(n17459) );
  NAND U18382 ( .A(n36926), .B(n17457), .Z(n17458) );
  NAND U18383 ( .A(n17459), .B(n17458), .Z(n17554) );
  XNOR U18384 ( .A(n17555), .B(n17554), .Z(n17548) );
  XOR U18385 ( .A(b[11]), .B(n20271), .Z(n17595) );
  OR U18386 ( .A(n17595), .B(n37311), .Z(n17462) );
  NANDN U18387 ( .A(n17460), .B(n37218), .Z(n17461) );
  NAND U18388 ( .A(n17462), .B(n17461), .Z(n17547) );
  XOR U18389 ( .A(n1053), .B(a[116]), .Z(n17598) );
  NANDN U18390 ( .A(n17598), .B(n37424), .Z(n17465) );
  NANDN U18391 ( .A(n17463), .B(n37425), .Z(n17464) );
  NAND U18392 ( .A(n17465), .B(n17464), .Z(n17546) );
  XNOR U18393 ( .A(n17547), .B(n17546), .Z(n17549) );
  XNOR U18394 ( .A(n17548), .B(n17549), .Z(n17537) );
  NANDN U18395 ( .A(n1049), .B(a[128]), .Z(n17466) );
  XNOR U18396 ( .A(b[1]), .B(n17466), .Z(n17468) );
  NANDN U18397 ( .A(b[0]), .B(a[127]), .Z(n17467) );
  AND U18398 ( .A(n17468), .B(n17467), .Z(n17512) );
  NAND U18399 ( .A(n38490), .B(n17469), .Z(n17471) );
  XNOR U18400 ( .A(n1058), .B(a[100]), .Z(n17604) );
  NANDN U18401 ( .A(n1048), .B(n17604), .Z(n17470) );
  NAND U18402 ( .A(n17471), .B(n17470), .Z(n17510) );
  NANDN U18403 ( .A(n1059), .B(a[96]), .Z(n17511) );
  XNOR U18404 ( .A(n17510), .B(n17511), .Z(n17513) );
  XNOR U18405 ( .A(n17512), .B(n17513), .Z(n17535) );
  NANDN U18406 ( .A(n17472), .B(n38205), .Z(n17474) );
  XNOR U18407 ( .A(b[23]), .B(a[106]), .Z(n17607) );
  OR U18408 ( .A(n17607), .B(n38268), .Z(n17473) );
  NAND U18409 ( .A(n17474), .B(n17473), .Z(n17577) );
  XOR U18410 ( .A(b[7]), .B(a[122]), .Z(n17610) );
  NAND U18411 ( .A(n17610), .B(n36701), .Z(n17477) );
  NAND U18412 ( .A(n17475), .B(n36702), .Z(n17476) );
  NAND U18413 ( .A(n17477), .B(n17476), .Z(n17574) );
  XOR U18414 ( .A(b[25]), .B(a[104]), .Z(n17613) );
  NAND U18415 ( .A(n17613), .B(n38325), .Z(n17480) );
  NAND U18416 ( .A(n17478), .B(n38326), .Z(n17479) );
  AND U18417 ( .A(n17480), .B(n17479), .Z(n17575) );
  XNOR U18418 ( .A(n17574), .B(n17575), .Z(n17576) );
  XOR U18419 ( .A(n17577), .B(n17576), .Z(n17534) );
  XOR U18420 ( .A(n17537), .B(n17536), .Z(n17565) );
  XNOR U18421 ( .A(n17564), .B(n17565), .Z(n17620) );
  XOR U18422 ( .A(n17621), .B(n17620), .Z(n17622) );
  XOR U18423 ( .A(n17623), .B(n17622), .Z(n17627) );
  XNOR U18424 ( .A(n17626), .B(n17627), .Z(n17628) );
  XOR U18425 ( .A(n17629), .B(n17628), .Z(n17635) );
  XOR U18426 ( .A(n17634), .B(n17635), .Z(n17506) );
  NANDN U18427 ( .A(n17482), .B(n17481), .Z(n17486) );
  NANDN U18428 ( .A(n17484), .B(n17483), .Z(n17485) );
  NAND U18429 ( .A(n17486), .B(n17485), .Z(n17505) );
  OR U18430 ( .A(n17488), .B(n17487), .Z(n17492) );
  OR U18431 ( .A(n17490), .B(n17489), .Z(n17491) );
  AND U18432 ( .A(n17492), .B(n17491), .Z(n17504) );
  XNOR U18433 ( .A(n17505), .B(n17504), .Z(n17507) );
  XOR U18434 ( .A(n17506), .B(n17507), .Z(n17498) );
  XOR U18435 ( .A(n17499), .B(n17498), .Z(n17500) );
  XNOR U18436 ( .A(n17501), .B(n17500), .Z(n17638) );
  XNOR U18437 ( .A(n17638), .B(sreg[352]), .Z(n17640) );
  NAND U18438 ( .A(n17493), .B(sreg[351]), .Z(n17497) );
  OR U18439 ( .A(n17495), .B(n17494), .Z(n17496) );
  AND U18440 ( .A(n17497), .B(n17496), .Z(n17639) );
  XOR U18441 ( .A(n17640), .B(n17639), .Z(c[352]) );
  NAND U18442 ( .A(n17499), .B(n17498), .Z(n17503) );
  NAND U18443 ( .A(n17501), .B(n17500), .Z(n17502) );
  NAND U18444 ( .A(n17503), .B(n17502), .Z(n17646) );
  NANDN U18445 ( .A(n17505), .B(n17504), .Z(n17509) );
  NAND U18446 ( .A(n17507), .B(n17506), .Z(n17508) );
  NAND U18447 ( .A(n17509), .B(n17508), .Z(n17644) );
  NANDN U18448 ( .A(n17511), .B(n17510), .Z(n17515) );
  NAND U18449 ( .A(n17513), .B(n17512), .Z(n17514) );
  NAND U18450 ( .A(n17515), .B(n17514), .Z(n17668) );
  XNOR U18451 ( .A(b[19]), .B(a[111]), .Z(n17717) );
  NANDN U18452 ( .A(n17717), .B(n37934), .Z(n17518) );
  NANDN U18453 ( .A(n17516), .B(n37935), .Z(n17517) );
  NAND U18454 ( .A(n17518), .B(n17517), .Z(n17678) );
  XOR U18455 ( .A(b[27]), .B(a[103]), .Z(n17720) );
  NAND U18456 ( .A(n38423), .B(n17720), .Z(n17521) );
  NAND U18457 ( .A(n17519), .B(n38424), .Z(n17520) );
  NAND U18458 ( .A(n17521), .B(n17520), .Z(n17675) );
  XNOR U18459 ( .A(b[5]), .B(a[125]), .Z(n17723) );
  NANDN U18460 ( .A(n17723), .B(n36587), .Z(n17524) );
  NANDN U18461 ( .A(n17522), .B(n36588), .Z(n17523) );
  AND U18462 ( .A(n17524), .B(n17523), .Z(n17676) );
  XNOR U18463 ( .A(n17675), .B(n17676), .Z(n17677) );
  XNOR U18464 ( .A(n17678), .B(n17677), .Z(n17666) );
  NAND U18465 ( .A(n17525), .B(n37762), .Z(n17527) );
  XNOR U18466 ( .A(b[17]), .B(a[113]), .Z(n17726) );
  NANDN U18467 ( .A(n17726), .B(n37764), .Z(n17526) );
  NAND U18468 ( .A(n17527), .B(n17526), .Z(n17744) );
  XOR U18469 ( .A(b[31]), .B(n17884), .Z(n17729) );
  NANDN U18470 ( .A(n17729), .B(n38552), .Z(n17530) );
  NANDN U18471 ( .A(n17528), .B(n38553), .Z(n17529) );
  NAND U18472 ( .A(n17530), .B(n17529), .Z(n17741) );
  OR U18473 ( .A(n17531), .B(n36105), .Z(n17533) );
  XNOR U18474 ( .A(b[3]), .B(a[127]), .Z(n17732) );
  NANDN U18475 ( .A(n17732), .B(n36107), .Z(n17532) );
  AND U18476 ( .A(n17533), .B(n17532), .Z(n17742) );
  XNOR U18477 ( .A(n17741), .B(n17742), .Z(n17743) );
  XOR U18478 ( .A(n17744), .B(n17743), .Z(n17665) );
  XNOR U18479 ( .A(n17666), .B(n17665), .Z(n17667) );
  XNOR U18480 ( .A(n17668), .B(n17667), .Z(n17763) );
  NANDN U18481 ( .A(n17535), .B(n17534), .Z(n17539) );
  NANDN U18482 ( .A(n17537), .B(n17536), .Z(n17538) );
  NAND U18483 ( .A(n17539), .B(n17538), .Z(n17764) );
  XNOR U18484 ( .A(n17763), .B(n17764), .Z(n17765) );
  NANDN U18485 ( .A(n17541), .B(n17540), .Z(n17545) );
  NAND U18486 ( .A(n17543), .B(n17542), .Z(n17544) );
  NAND U18487 ( .A(n17545), .B(n17544), .Z(n17658) );
  OR U18488 ( .A(n17547), .B(n17546), .Z(n17551) );
  NANDN U18489 ( .A(n17549), .B(n17548), .Z(n17550) );
  NAND U18490 ( .A(n17551), .B(n17550), .Z(n17656) );
  XNOR U18491 ( .A(n17656), .B(n17655), .Z(n17657) );
  XOR U18492 ( .A(n17658), .B(n17657), .Z(n17766) );
  XOR U18493 ( .A(n17765), .B(n17766), .Z(n17776) );
  OR U18494 ( .A(n17557), .B(n17556), .Z(n17561) );
  NANDN U18495 ( .A(n17559), .B(n17558), .Z(n17560) );
  NAND U18496 ( .A(n17561), .B(n17560), .Z(n17774) );
  NANDN U18497 ( .A(n17563), .B(n17562), .Z(n17567) );
  NANDN U18498 ( .A(n17565), .B(n17564), .Z(n17566) );
  NAND U18499 ( .A(n17567), .B(n17566), .Z(n17759) );
  NANDN U18500 ( .A(n17569), .B(n17568), .Z(n17573) );
  NAND U18501 ( .A(n17571), .B(n17570), .Z(n17572) );
  NAND U18502 ( .A(n17573), .B(n17572), .Z(n17758) );
  NANDN U18503 ( .A(n17575), .B(n17574), .Z(n17579) );
  NAND U18504 ( .A(n17577), .B(n17576), .Z(n17578) );
  NAND U18505 ( .A(n17579), .B(n17578), .Z(n17659) );
  NANDN U18506 ( .A(n17581), .B(n17580), .Z(n17585) );
  NAND U18507 ( .A(n17583), .B(n17582), .Z(n17584) );
  AND U18508 ( .A(n17585), .B(n17584), .Z(n17660) );
  XNOR U18509 ( .A(n17659), .B(n17660), .Z(n17661) );
  XNOR U18510 ( .A(b[21]), .B(a[109]), .Z(n17687) );
  NANDN U18511 ( .A(n17687), .B(n38101), .Z(n17588) );
  NANDN U18512 ( .A(n17586), .B(n38102), .Z(n17587) );
  NAND U18513 ( .A(n17588), .B(n17587), .Z(n17753) );
  XNOR U18514 ( .A(b[15]), .B(a[115]), .Z(n17684) );
  OR U18515 ( .A(n17684), .B(n37665), .Z(n17591) );
  NANDN U18516 ( .A(n17589), .B(n37604), .Z(n17590) );
  AND U18517 ( .A(n17591), .B(n17590), .Z(n17754) );
  XNOR U18518 ( .A(n17753), .B(n17754), .Z(n17756) );
  XNOR U18519 ( .A(b[9]), .B(a[121]), .Z(n17681) );
  NANDN U18520 ( .A(n17681), .B(n36925), .Z(n17594) );
  NANDN U18521 ( .A(n17592), .B(n36926), .Z(n17593) );
  NAND U18522 ( .A(n17594), .B(n17593), .Z(n17755) );
  XNOR U18523 ( .A(n17756), .B(n17755), .Z(n17749) );
  XNOR U18524 ( .A(b[11]), .B(a[119]), .Z(n17690) );
  OR U18525 ( .A(n17690), .B(n37311), .Z(n17597) );
  NANDN U18526 ( .A(n17595), .B(n37218), .Z(n17596) );
  NAND U18527 ( .A(n17597), .B(n17596), .Z(n17748) );
  XOR U18528 ( .A(n1053), .B(a[117]), .Z(n17693) );
  NANDN U18529 ( .A(n17693), .B(n37424), .Z(n17600) );
  NANDN U18530 ( .A(n17598), .B(n37425), .Z(n17599) );
  NAND U18531 ( .A(n17600), .B(n17599), .Z(n17747) );
  XNOR U18532 ( .A(n17748), .B(n17747), .Z(n17750) );
  XNOR U18533 ( .A(n17749), .B(n17750), .Z(n17738) );
  NANDN U18534 ( .A(n1049), .B(a[129]), .Z(n17601) );
  XNOR U18535 ( .A(b[1]), .B(n17601), .Z(n17603) );
  NANDN U18536 ( .A(b[0]), .B(a[128]), .Z(n17602) );
  AND U18537 ( .A(n17603), .B(n17602), .Z(n17713) );
  NAND U18538 ( .A(n38490), .B(n17604), .Z(n17606) );
  XOR U18539 ( .A(n1058), .B(n17812), .Z(n17699) );
  NANDN U18540 ( .A(n1048), .B(n17699), .Z(n17605) );
  NAND U18541 ( .A(n17606), .B(n17605), .Z(n17711) );
  NANDN U18542 ( .A(n1059), .B(a[97]), .Z(n17712) );
  XNOR U18543 ( .A(n17711), .B(n17712), .Z(n17714) );
  XNOR U18544 ( .A(n17713), .B(n17714), .Z(n17736) );
  NANDN U18545 ( .A(n17607), .B(n38205), .Z(n17609) );
  XOR U18546 ( .A(b[23]), .B(n18980), .Z(n17702) );
  OR U18547 ( .A(n17702), .B(n38268), .Z(n17608) );
  NAND U18548 ( .A(n17609), .B(n17608), .Z(n17672) );
  XOR U18549 ( .A(b[7]), .B(a[123]), .Z(n17705) );
  NAND U18550 ( .A(n17705), .B(n36701), .Z(n17612) );
  NAND U18551 ( .A(n17610), .B(n36702), .Z(n17611) );
  NAND U18552 ( .A(n17612), .B(n17611), .Z(n17669) );
  XOR U18553 ( .A(b[25]), .B(a[105]), .Z(n17708) );
  NAND U18554 ( .A(n17708), .B(n38325), .Z(n17615) );
  NAND U18555 ( .A(n17613), .B(n38326), .Z(n17614) );
  AND U18556 ( .A(n17615), .B(n17614), .Z(n17670) );
  XNOR U18557 ( .A(n17669), .B(n17670), .Z(n17671) );
  XOR U18558 ( .A(n17672), .B(n17671), .Z(n17735) );
  XOR U18559 ( .A(n17738), .B(n17737), .Z(n17662) );
  XNOR U18560 ( .A(n17661), .B(n17662), .Z(n17757) );
  XNOR U18561 ( .A(n17758), .B(n17757), .Z(n17760) );
  XNOR U18562 ( .A(n17759), .B(n17760), .Z(n17773) );
  XOR U18563 ( .A(n17774), .B(n17773), .Z(n17775) );
  XNOR U18564 ( .A(n17776), .B(n17775), .Z(n17770) );
  NAND U18565 ( .A(n17621), .B(n17620), .Z(n17625) );
  NAND U18566 ( .A(n17623), .B(n17622), .Z(n17624) );
  AND U18567 ( .A(n17625), .B(n17624), .Z(n17767) );
  XNOR U18568 ( .A(n17768), .B(n17767), .Z(n17769) );
  XOR U18569 ( .A(n17770), .B(n17769), .Z(n17651) );
  NANDN U18570 ( .A(n17627), .B(n17626), .Z(n17631) );
  NAND U18571 ( .A(n17629), .B(n17628), .Z(n17630) );
  NAND U18572 ( .A(n17631), .B(n17630), .Z(n17649) );
  NANDN U18573 ( .A(n17633), .B(n17632), .Z(n17637) );
  NAND U18574 ( .A(n17635), .B(n17634), .Z(n17636) );
  AND U18575 ( .A(n17637), .B(n17636), .Z(n17650) );
  XNOR U18576 ( .A(n17649), .B(n17650), .Z(n17652) );
  XOR U18577 ( .A(n17651), .B(n17652), .Z(n17643) );
  XOR U18578 ( .A(n17644), .B(n17643), .Z(n17645) );
  XNOR U18579 ( .A(n17646), .B(n17645), .Z(n17779) );
  XNOR U18580 ( .A(n17779), .B(sreg[353]), .Z(n17781) );
  NAND U18581 ( .A(n17638), .B(sreg[352]), .Z(n17642) );
  OR U18582 ( .A(n17640), .B(n17639), .Z(n17641) );
  AND U18583 ( .A(n17642), .B(n17641), .Z(n17780) );
  XOR U18584 ( .A(n17781), .B(n17780), .Z(c[353]) );
  NAND U18585 ( .A(n17644), .B(n17643), .Z(n17648) );
  NAND U18586 ( .A(n17646), .B(n17645), .Z(n17647) );
  NAND U18587 ( .A(n17648), .B(n17647), .Z(n17787) );
  NANDN U18588 ( .A(n17650), .B(n17649), .Z(n17654) );
  NAND U18589 ( .A(n17652), .B(n17651), .Z(n17653) );
  NAND U18590 ( .A(n17654), .B(n17653), .Z(n17785) );
  NANDN U18591 ( .A(n17660), .B(n17659), .Z(n17664) );
  NANDN U18592 ( .A(n17662), .B(n17661), .Z(n17663) );
  NAND U18593 ( .A(n17664), .B(n17663), .Z(n17903) );
  NANDN U18594 ( .A(n17670), .B(n17669), .Z(n17674) );
  NAND U18595 ( .A(n17672), .B(n17671), .Z(n17673) );
  NAND U18596 ( .A(n17674), .B(n17673), .Z(n17847) );
  NANDN U18597 ( .A(n17676), .B(n17675), .Z(n17680) );
  NAND U18598 ( .A(n17678), .B(n17677), .Z(n17679) );
  AND U18599 ( .A(n17680), .B(n17679), .Z(n17848) );
  XNOR U18600 ( .A(n17847), .B(n17848), .Z(n17849) );
  XNOR U18601 ( .A(b[9]), .B(a[122]), .Z(n17869) );
  NANDN U18602 ( .A(n17869), .B(n36925), .Z(n17683) );
  NANDN U18603 ( .A(n17681), .B(n36926), .Z(n17682) );
  NAND U18604 ( .A(n17683), .B(n17682), .Z(n17833) );
  XNOR U18605 ( .A(b[15]), .B(a[116]), .Z(n17872) );
  OR U18606 ( .A(n17872), .B(n37665), .Z(n17686) );
  NANDN U18607 ( .A(n17684), .B(n37604), .Z(n17685) );
  AND U18608 ( .A(n17686), .B(n17685), .Z(n17831) );
  XNOR U18609 ( .A(b[21]), .B(a[110]), .Z(n17875) );
  NANDN U18610 ( .A(n17875), .B(n38101), .Z(n17689) );
  NANDN U18611 ( .A(n17687), .B(n38102), .Z(n17688) );
  AND U18612 ( .A(n17689), .B(n17688), .Z(n17832) );
  XOR U18613 ( .A(n17833), .B(n17834), .Z(n17822) );
  XNOR U18614 ( .A(b[11]), .B(a[120]), .Z(n17878) );
  OR U18615 ( .A(n17878), .B(n37311), .Z(n17692) );
  NANDN U18616 ( .A(n17690), .B(n37218), .Z(n17691) );
  NAND U18617 ( .A(n17692), .B(n17691), .Z(n17820) );
  XOR U18618 ( .A(n1053), .B(a[118]), .Z(n17881) );
  NANDN U18619 ( .A(n17881), .B(n37424), .Z(n17695) );
  NANDN U18620 ( .A(n17693), .B(n37425), .Z(n17694) );
  AND U18621 ( .A(n17695), .B(n17694), .Z(n17819) );
  XNOR U18622 ( .A(n17820), .B(n17819), .Z(n17821) );
  XOR U18623 ( .A(n17822), .B(n17821), .Z(n17839) );
  NANDN U18624 ( .A(n1049), .B(a[130]), .Z(n17696) );
  XNOR U18625 ( .A(b[1]), .B(n17696), .Z(n17698) );
  IV U18626 ( .A(a[129]), .Z(n22221) );
  NANDN U18627 ( .A(n22221), .B(n1049), .Z(n17697) );
  AND U18628 ( .A(n17698), .B(n17697), .Z(n17796) );
  NAND U18629 ( .A(n38490), .B(n17699), .Z(n17701) );
  XNOR U18630 ( .A(b[29]), .B(a[102]), .Z(n17885) );
  OR U18631 ( .A(n17885), .B(n1048), .Z(n17700) );
  NAND U18632 ( .A(n17701), .B(n17700), .Z(n17794) );
  NANDN U18633 ( .A(n1059), .B(a[98]), .Z(n17795) );
  XNOR U18634 ( .A(n17794), .B(n17795), .Z(n17797) );
  XOR U18635 ( .A(n17796), .B(n17797), .Z(n17837) );
  NANDN U18636 ( .A(n17702), .B(n38205), .Z(n17704) );
  XNOR U18637 ( .A(b[23]), .B(a[108]), .Z(n17891) );
  OR U18638 ( .A(n17891), .B(n38268), .Z(n17703) );
  NAND U18639 ( .A(n17704), .B(n17703), .Z(n17860) );
  XOR U18640 ( .A(b[7]), .B(a[124]), .Z(n17894) );
  NAND U18641 ( .A(n17894), .B(n36701), .Z(n17707) );
  NAND U18642 ( .A(n17705), .B(n36702), .Z(n17706) );
  NAND U18643 ( .A(n17707), .B(n17706), .Z(n17857) );
  XOR U18644 ( .A(b[25]), .B(a[106]), .Z(n17897) );
  NAND U18645 ( .A(n17897), .B(n38325), .Z(n17710) );
  NAND U18646 ( .A(n17708), .B(n38326), .Z(n17709) );
  AND U18647 ( .A(n17710), .B(n17709), .Z(n17858) );
  XNOR U18648 ( .A(n17857), .B(n17858), .Z(n17859) );
  XNOR U18649 ( .A(n17860), .B(n17859), .Z(n17838) );
  XOR U18650 ( .A(n17837), .B(n17838), .Z(n17840) );
  XNOR U18651 ( .A(n17839), .B(n17840), .Z(n17850) );
  XOR U18652 ( .A(n17849), .B(n17850), .Z(n17901) );
  XNOR U18653 ( .A(n17900), .B(n17901), .Z(n17902) );
  XOR U18654 ( .A(n17903), .B(n17902), .Z(n17911) );
  XNOR U18655 ( .A(n17910), .B(n17911), .Z(n17913) );
  NANDN U18656 ( .A(n17712), .B(n17711), .Z(n17716) );
  NAND U18657 ( .A(n17714), .B(n17713), .Z(n17715) );
  NAND U18658 ( .A(n17716), .B(n17715), .Z(n17856) );
  XNOR U18659 ( .A(b[19]), .B(a[112]), .Z(n17800) );
  NANDN U18660 ( .A(n17800), .B(n37934), .Z(n17719) );
  NANDN U18661 ( .A(n17717), .B(n37935), .Z(n17718) );
  NAND U18662 ( .A(n17719), .B(n17718), .Z(n17866) );
  XOR U18663 ( .A(b[27]), .B(a[104]), .Z(n17803) );
  NAND U18664 ( .A(n38423), .B(n17803), .Z(n17722) );
  NAND U18665 ( .A(n17720), .B(n38424), .Z(n17721) );
  NAND U18666 ( .A(n17722), .B(n17721), .Z(n17863) );
  XNOR U18667 ( .A(b[5]), .B(a[126]), .Z(n17806) );
  NANDN U18668 ( .A(n17806), .B(n36587), .Z(n17725) );
  NANDN U18669 ( .A(n17723), .B(n36588), .Z(n17724) );
  AND U18670 ( .A(n17725), .B(n17724), .Z(n17864) );
  XNOR U18671 ( .A(n17863), .B(n17864), .Z(n17865) );
  XNOR U18672 ( .A(n17866), .B(n17865), .Z(n17854) );
  NANDN U18673 ( .A(n17726), .B(n37762), .Z(n17728) );
  XOR U18674 ( .A(b[17]), .B(a[114]), .Z(n17809) );
  NAND U18675 ( .A(n17809), .B(n37764), .Z(n17727) );
  NAND U18676 ( .A(n17728), .B(n17727), .Z(n17828) );
  XNOR U18677 ( .A(b[31]), .B(a[100]), .Z(n17813) );
  NANDN U18678 ( .A(n17813), .B(n38552), .Z(n17731) );
  NANDN U18679 ( .A(n17729), .B(n38553), .Z(n17730) );
  NAND U18680 ( .A(n17731), .B(n17730), .Z(n17825) );
  OR U18681 ( .A(n17732), .B(n36105), .Z(n17734) );
  XNOR U18682 ( .A(b[3]), .B(a[128]), .Z(n17816) );
  NANDN U18683 ( .A(n17816), .B(n36107), .Z(n17733) );
  AND U18684 ( .A(n17734), .B(n17733), .Z(n17826) );
  XNOR U18685 ( .A(n17825), .B(n17826), .Z(n17827) );
  XOR U18686 ( .A(n17828), .B(n17827), .Z(n17853) );
  XNOR U18687 ( .A(n17854), .B(n17853), .Z(n17855) );
  XNOR U18688 ( .A(n17856), .B(n17855), .Z(n17906) );
  NANDN U18689 ( .A(n17736), .B(n17735), .Z(n17740) );
  NANDN U18690 ( .A(n17738), .B(n17737), .Z(n17739) );
  NAND U18691 ( .A(n17740), .B(n17739), .Z(n17907) );
  XNOR U18692 ( .A(n17906), .B(n17907), .Z(n17908) );
  NANDN U18693 ( .A(n17742), .B(n17741), .Z(n17746) );
  NAND U18694 ( .A(n17744), .B(n17743), .Z(n17745) );
  NAND U18695 ( .A(n17746), .B(n17745), .Z(n17846) );
  OR U18696 ( .A(n17748), .B(n17747), .Z(n17752) );
  NANDN U18697 ( .A(n17750), .B(n17749), .Z(n17751) );
  NAND U18698 ( .A(n17752), .B(n17751), .Z(n17844) );
  XNOR U18699 ( .A(n17844), .B(n17843), .Z(n17845) );
  XOR U18700 ( .A(n17846), .B(n17845), .Z(n17909) );
  XOR U18701 ( .A(n17908), .B(n17909), .Z(n17912) );
  XOR U18702 ( .A(n17913), .B(n17912), .Z(n17917) );
  NAND U18703 ( .A(n17758), .B(n17757), .Z(n17762) );
  NANDN U18704 ( .A(n17760), .B(n17759), .Z(n17761) );
  NAND U18705 ( .A(n17762), .B(n17761), .Z(n17914) );
  XNOR U18706 ( .A(n17914), .B(n17915), .Z(n17916) );
  XNOR U18707 ( .A(n17917), .B(n17916), .Z(n17791) );
  NANDN U18708 ( .A(n17768), .B(n17767), .Z(n17772) );
  NAND U18709 ( .A(n17770), .B(n17769), .Z(n17771) );
  NAND U18710 ( .A(n17772), .B(n17771), .Z(n17788) );
  NANDN U18711 ( .A(n17774), .B(n17773), .Z(n17778) );
  OR U18712 ( .A(n17776), .B(n17775), .Z(n17777) );
  NAND U18713 ( .A(n17778), .B(n17777), .Z(n17789) );
  XNOR U18714 ( .A(n17788), .B(n17789), .Z(n17790) );
  XNOR U18715 ( .A(n17791), .B(n17790), .Z(n17784) );
  XOR U18716 ( .A(n17785), .B(n17784), .Z(n17786) );
  XNOR U18717 ( .A(n17787), .B(n17786), .Z(n17920) );
  XNOR U18718 ( .A(n17920), .B(sreg[354]), .Z(n17922) );
  NAND U18719 ( .A(n17779), .B(sreg[353]), .Z(n17783) );
  OR U18720 ( .A(n17781), .B(n17780), .Z(n17782) );
  AND U18721 ( .A(n17783), .B(n17782), .Z(n17921) );
  XOR U18722 ( .A(n17922), .B(n17921), .Z(c[354]) );
  NANDN U18723 ( .A(n17789), .B(n17788), .Z(n17793) );
  NANDN U18724 ( .A(n17791), .B(n17790), .Z(n17792) );
  NAND U18725 ( .A(n17793), .B(n17792), .Z(n17926) );
  NANDN U18726 ( .A(n17795), .B(n17794), .Z(n17799) );
  NAND U18727 ( .A(n17797), .B(n17796), .Z(n17798) );
  NAND U18728 ( .A(n17799), .B(n17798), .Z(n17998) );
  XOR U18729 ( .A(b[19]), .B(n19909), .Z(n17965) );
  NANDN U18730 ( .A(n17965), .B(n37934), .Z(n17802) );
  NANDN U18731 ( .A(n17800), .B(n37935), .Z(n17801) );
  NAND U18732 ( .A(n17802), .B(n17801), .Z(n18010) );
  XOR U18733 ( .A(b[27]), .B(a[105]), .Z(n17968) );
  NAND U18734 ( .A(n38423), .B(n17968), .Z(n17805) );
  NAND U18735 ( .A(n17803), .B(n38424), .Z(n17804) );
  NAND U18736 ( .A(n17805), .B(n17804), .Z(n18007) );
  XNOR U18737 ( .A(b[5]), .B(a[127]), .Z(n17971) );
  NANDN U18738 ( .A(n17971), .B(n36587), .Z(n17808) );
  NANDN U18739 ( .A(n17806), .B(n36588), .Z(n17807) );
  AND U18740 ( .A(n17808), .B(n17807), .Z(n18008) );
  XNOR U18741 ( .A(n18007), .B(n18008), .Z(n18009) );
  XNOR U18742 ( .A(n18010), .B(n18009), .Z(n17995) );
  NAND U18743 ( .A(n17809), .B(n37762), .Z(n17811) );
  XOR U18744 ( .A(b[17]), .B(a[115]), .Z(n17974) );
  NAND U18745 ( .A(n17974), .B(n37764), .Z(n17810) );
  NAND U18746 ( .A(n17811), .B(n17810), .Z(n17949) );
  XOR U18747 ( .A(b[31]), .B(n17812), .Z(n17977) );
  NANDN U18748 ( .A(n17977), .B(n38552), .Z(n17815) );
  NANDN U18749 ( .A(n17813), .B(n38553), .Z(n17814) );
  AND U18750 ( .A(n17815), .B(n17814), .Z(n17947) );
  OR U18751 ( .A(n17816), .B(n36105), .Z(n17818) );
  XOR U18752 ( .A(b[3]), .B(n22221), .Z(n17980) );
  NANDN U18753 ( .A(n17980), .B(n36107), .Z(n17817) );
  AND U18754 ( .A(n17818), .B(n17817), .Z(n17948) );
  XOR U18755 ( .A(n17949), .B(n17950), .Z(n17996) );
  XOR U18756 ( .A(n17995), .B(n17996), .Z(n17997) );
  XNOR U18757 ( .A(n17998), .B(n17997), .Z(n18043) );
  NANDN U18758 ( .A(n17820), .B(n17819), .Z(n17824) );
  NAND U18759 ( .A(n17822), .B(n17821), .Z(n17823) );
  NAND U18760 ( .A(n17824), .B(n17823), .Z(n17986) );
  NANDN U18761 ( .A(n17826), .B(n17825), .Z(n17830) );
  NAND U18762 ( .A(n17828), .B(n17827), .Z(n17829) );
  NAND U18763 ( .A(n17830), .B(n17829), .Z(n17984) );
  OR U18764 ( .A(n17832), .B(n17831), .Z(n17836) );
  NANDN U18765 ( .A(n17834), .B(n17833), .Z(n17835) );
  NAND U18766 ( .A(n17836), .B(n17835), .Z(n17983) );
  XNOR U18767 ( .A(n17986), .B(n17985), .Z(n18044) );
  XNOR U18768 ( .A(n18043), .B(n18044), .Z(n18045) );
  NANDN U18769 ( .A(n17838), .B(n17837), .Z(n17842) );
  OR U18770 ( .A(n17840), .B(n17839), .Z(n17841) );
  AND U18771 ( .A(n17842), .B(n17841), .Z(n18046) );
  XNOR U18772 ( .A(n18045), .B(n18046), .Z(n18058) );
  NANDN U18773 ( .A(n17848), .B(n17847), .Z(n17852) );
  NANDN U18774 ( .A(n17850), .B(n17849), .Z(n17851) );
  NAND U18775 ( .A(n17852), .B(n17851), .Z(n18052) );
  NANDN U18776 ( .A(n17858), .B(n17857), .Z(n17862) );
  NAND U18777 ( .A(n17860), .B(n17859), .Z(n17861) );
  NAND U18778 ( .A(n17862), .B(n17861), .Z(n17989) );
  NANDN U18779 ( .A(n17864), .B(n17863), .Z(n17868) );
  NAND U18780 ( .A(n17866), .B(n17865), .Z(n17867) );
  AND U18781 ( .A(n17868), .B(n17867), .Z(n17990) );
  XNOR U18782 ( .A(n17989), .B(n17990), .Z(n17991) );
  XNOR U18783 ( .A(b[9]), .B(a[123]), .Z(n18013) );
  NANDN U18784 ( .A(n18013), .B(n36925), .Z(n17871) );
  NANDN U18785 ( .A(n17869), .B(n36926), .Z(n17870) );
  NAND U18786 ( .A(n17871), .B(n17870), .Z(n17955) );
  XNOR U18787 ( .A(b[15]), .B(a[117]), .Z(n18016) );
  OR U18788 ( .A(n18016), .B(n37665), .Z(n17874) );
  NANDN U18789 ( .A(n17872), .B(n37604), .Z(n17873) );
  AND U18790 ( .A(n17874), .B(n17873), .Z(n17953) );
  XNOR U18791 ( .A(b[21]), .B(a[111]), .Z(n18019) );
  NANDN U18792 ( .A(n18019), .B(n38101), .Z(n17877) );
  NANDN U18793 ( .A(n17875), .B(n38102), .Z(n17876) );
  AND U18794 ( .A(n17877), .B(n17876), .Z(n17954) );
  XOR U18795 ( .A(n17955), .B(n17956), .Z(n17944) );
  XNOR U18796 ( .A(b[11]), .B(a[121]), .Z(n18022) );
  OR U18797 ( .A(n18022), .B(n37311), .Z(n17880) );
  NANDN U18798 ( .A(n17878), .B(n37218), .Z(n17879) );
  NAND U18799 ( .A(n17880), .B(n17879), .Z(n17942) );
  XOR U18800 ( .A(n1053), .B(a[119]), .Z(n18025) );
  NANDN U18801 ( .A(n18025), .B(n37424), .Z(n17883) );
  NANDN U18802 ( .A(n17881), .B(n37425), .Z(n17882) );
  NAND U18803 ( .A(n17883), .B(n17882), .Z(n17941) );
  XOR U18804 ( .A(n17944), .B(n17943), .Z(n17938) );
  ANDN U18805 ( .B(b[31]), .A(n17884), .Z(n17959) );
  NANDN U18806 ( .A(n17885), .B(n38490), .Z(n17887) );
  XNOR U18807 ( .A(n1058), .B(a[103]), .Z(n18031) );
  NANDN U18808 ( .A(n1048), .B(n18031), .Z(n17886) );
  NAND U18809 ( .A(n17887), .B(n17886), .Z(n17960) );
  XOR U18810 ( .A(n17959), .B(n17960), .Z(n17961) );
  NANDN U18811 ( .A(n1049), .B(a[131]), .Z(n17888) );
  XNOR U18812 ( .A(b[1]), .B(n17888), .Z(n17890) );
  NANDN U18813 ( .A(b[0]), .B(a[130]), .Z(n17889) );
  AND U18814 ( .A(n17890), .B(n17889), .Z(n17962) );
  XNOR U18815 ( .A(n17961), .B(n17962), .Z(n17935) );
  NANDN U18816 ( .A(n17891), .B(n38205), .Z(n17893) );
  XNOR U18817 ( .A(b[23]), .B(a[109]), .Z(n18034) );
  OR U18818 ( .A(n18034), .B(n38268), .Z(n17892) );
  NAND U18819 ( .A(n17893), .B(n17892), .Z(n18004) );
  XOR U18820 ( .A(b[7]), .B(a[125]), .Z(n18037) );
  NAND U18821 ( .A(n18037), .B(n36701), .Z(n17896) );
  NAND U18822 ( .A(n17894), .B(n36702), .Z(n17895) );
  NAND U18823 ( .A(n17896), .B(n17895), .Z(n18001) );
  XNOR U18824 ( .A(b[25]), .B(a[107]), .Z(n18040) );
  NANDN U18825 ( .A(n18040), .B(n38325), .Z(n17899) );
  NAND U18826 ( .A(n17897), .B(n38326), .Z(n17898) );
  AND U18827 ( .A(n17899), .B(n17898), .Z(n18002) );
  XNOR U18828 ( .A(n18001), .B(n18002), .Z(n18003) );
  XNOR U18829 ( .A(n18004), .B(n18003), .Z(n17936) );
  XOR U18830 ( .A(n17938), .B(n17937), .Z(n17992) );
  XNOR U18831 ( .A(n17991), .B(n17992), .Z(n18049) );
  XOR U18832 ( .A(n18050), .B(n18049), .Z(n18051) );
  XOR U18833 ( .A(n18052), .B(n18051), .Z(n18056) );
  XNOR U18834 ( .A(n18055), .B(n18056), .Z(n18057) );
  XNOR U18835 ( .A(n18058), .B(n18057), .Z(n18062) );
  NANDN U18836 ( .A(n17901), .B(n17900), .Z(n17905) );
  NAND U18837 ( .A(n17903), .B(n17902), .Z(n17904) );
  NAND U18838 ( .A(n17905), .B(n17904), .Z(n18059) );
  XNOR U18839 ( .A(n18059), .B(n18060), .Z(n18061) );
  XNOR U18840 ( .A(n18062), .B(n18061), .Z(n17932) );
  NANDN U18841 ( .A(n17915), .B(n17914), .Z(n17919) );
  NANDN U18842 ( .A(n17917), .B(n17916), .Z(n17918) );
  NAND U18843 ( .A(n17919), .B(n17918), .Z(n17930) );
  XNOR U18844 ( .A(n17929), .B(n17930), .Z(n17931) );
  XNOR U18845 ( .A(n17932), .B(n17931), .Z(n17925) );
  XOR U18846 ( .A(n17926), .B(n17925), .Z(n17927) );
  XNOR U18847 ( .A(n17928), .B(n17927), .Z(n18065) );
  XNOR U18848 ( .A(n18065), .B(sreg[355]), .Z(n18067) );
  NAND U18849 ( .A(n17920), .B(sreg[354]), .Z(n17924) );
  OR U18850 ( .A(n17922), .B(n17921), .Z(n17923) );
  AND U18851 ( .A(n17924), .B(n17923), .Z(n18066) );
  XOR U18852 ( .A(n18067), .B(n18066), .Z(c[355]) );
  NANDN U18853 ( .A(n17930), .B(n17929), .Z(n17934) );
  NANDN U18854 ( .A(n17932), .B(n17931), .Z(n17933) );
  NAND U18855 ( .A(n17934), .B(n17933), .Z(n18071) );
  OR U18856 ( .A(n17936), .B(n17935), .Z(n17940) );
  NANDN U18857 ( .A(n17938), .B(n17937), .Z(n17939) );
  NAND U18858 ( .A(n17940), .B(n17939), .Z(n18203) );
  OR U18859 ( .A(n17942), .B(n17941), .Z(n17946) );
  NAND U18860 ( .A(n17944), .B(n17943), .Z(n17945) );
  NAND U18861 ( .A(n17946), .B(n17945), .Z(n18142) );
  OR U18862 ( .A(n17948), .B(n17947), .Z(n17952) );
  NANDN U18863 ( .A(n17950), .B(n17949), .Z(n17951) );
  NAND U18864 ( .A(n17952), .B(n17951), .Z(n18141) );
  OR U18865 ( .A(n17954), .B(n17953), .Z(n17958) );
  NANDN U18866 ( .A(n17956), .B(n17955), .Z(n17957) );
  NAND U18867 ( .A(n17958), .B(n17957), .Z(n18140) );
  XOR U18868 ( .A(n18142), .B(n18143), .Z(n18201) );
  OR U18869 ( .A(n17960), .B(n17959), .Z(n17964) );
  NANDN U18870 ( .A(n17962), .B(n17961), .Z(n17963) );
  NAND U18871 ( .A(n17964), .B(n17963), .Z(n18155) );
  XNOR U18872 ( .A(b[19]), .B(a[114]), .Z(n18122) );
  NANDN U18873 ( .A(n18122), .B(n37934), .Z(n17967) );
  NANDN U18874 ( .A(n17965), .B(n37935), .Z(n17966) );
  NAND U18875 ( .A(n17967), .B(n17966), .Z(n18167) );
  XOR U18876 ( .A(b[27]), .B(a[106]), .Z(n18125) );
  NAND U18877 ( .A(n38423), .B(n18125), .Z(n17970) );
  NAND U18878 ( .A(n17968), .B(n38424), .Z(n17969) );
  NAND U18879 ( .A(n17970), .B(n17969), .Z(n18164) );
  XNOR U18880 ( .A(b[5]), .B(a[128]), .Z(n18128) );
  NANDN U18881 ( .A(n18128), .B(n36587), .Z(n17973) );
  NANDN U18882 ( .A(n17971), .B(n36588), .Z(n17972) );
  AND U18883 ( .A(n17973), .B(n17972), .Z(n18165) );
  XNOR U18884 ( .A(n18164), .B(n18165), .Z(n18166) );
  XNOR U18885 ( .A(n18167), .B(n18166), .Z(n18152) );
  NAND U18886 ( .A(n17974), .B(n37762), .Z(n17976) );
  XOR U18887 ( .A(b[17]), .B(a[116]), .Z(n18131) );
  NAND U18888 ( .A(n18131), .B(n37764), .Z(n17975) );
  NAND U18889 ( .A(n17976), .B(n17975), .Z(n18106) );
  XNOR U18890 ( .A(b[31]), .B(a[102]), .Z(n18134) );
  NANDN U18891 ( .A(n18134), .B(n38552), .Z(n17979) );
  NANDN U18892 ( .A(n17977), .B(n38553), .Z(n17978) );
  AND U18893 ( .A(n17979), .B(n17978), .Z(n18104) );
  OR U18894 ( .A(n17980), .B(n36105), .Z(n17982) );
  XNOR U18895 ( .A(b[3]), .B(a[130]), .Z(n18137) );
  NANDN U18896 ( .A(n18137), .B(n36107), .Z(n17981) );
  AND U18897 ( .A(n17982), .B(n17981), .Z(n18105) );
  XOR U18898 ( .A(n18106), .B(n18107), .Z(n18153) );
  XOR U18899 ( .A(n18152), .B(n18153), .Z(n18154) );
  XNOR U18900 ( .A(n18155), .B(n18154), .Z(n18200) );
  XOR U18901 ( .A(n18201), .B(n18200), .Z(n18202) );
  XNOR U18902 ( .A(n18203), .B(n18202), .Z(n18089) );
  OR U18903 ( .A(n17984), .B(n17983), .Z(n17988) );
  NAND U18904 ( .A(n17986), .B(n17985), .Z(n17987) );
  NAND U18905 ( .A(n17988), .B(n17987), .Z(n18087) );
  NANDN U18906 ( .A(n17990), .B(n17989), .Z(n17994) );
  NANDN U18907 ( .A(n17992), .B(n17991), .Z(n17993) );
  NAND U18908 ( .A(n17994), .B(n17993), .Z(n18206) );
  OR U18909 ( .A(n17996), .B(n17995), .Z(n18000) );
  NAND U18910 ( .A(n17998), .B(n17997), .Z(n17999) );
  NAND U18911 ( .A(n18000), .B(n17999), .Z(n18205) );
  NANDN U18912 ( .A(n18002), .B(n18001), .Z(n18006) );
  NAND U18913 ( .A(n18004), .B(n18003), .Z(n18005) );
  NAND U18914 ( .A(n18006), .B(n18005), .Z(n18146) );
  NANDN U18915 ( .A(n18008), .B(n18007), .Z(n18012) );
  NAND U18916 ( .A(n18010), .B(n18009), .Z(n18011) );
  AND U18917 ( .A(n18012), .B(n18011), .Z(n18147) );
  XNOR U18918 ( .A(n18146), .B(n18147), .Z(n18148) );
  XNOR U18919 ( .A(n1052), .B(a[124]), .Z(n18170) );
  NAND U18920 ( .A(n36925), .B(n18170), .Z(n18015) );
  NANDN U18921 ( .A(n18013), .B(n36926), .Z(n18014) );
  NAND U18922 ( .A(n18015), .B(n18014), .Z(n18112) );
  XOR U18923 ( .A(b[15]), .B(n20271), .Z(n18173) );
  OR U18924 ( .A(n18173), .B(n37665), .Z(n18018) );
  NANDN U18925 ( .A(n18016), .B(n37604), .Z(n18017) );
  AND U18926 ( .A(n18018), .B(n18017), .Z(n18110) );
  XNOR U18927 ( .A(n1056), .B(a[112]), .Z(n18176) );
  NAND U18928 ( .A(n18176), .B(n38101), .Z(n18021) );
  NANDN U18929 ( .A(n18019), .B(n38102), .Z(n18020) );
  AND U18930 ( .A(n18021), .B(n18020), .Z(n18111) );
  XOR U18931 ( .A(n18112), .B(n18113), .Z(n18101) );
  XNOR U18932 ( .A(b[11]), .B(a[122]), .Z(n18179) );
  OR U18933 ( .A(n18179), .B(n37311), .Z(n18024) );
  NANDN U18934 ( .A(n18022), .B(n37218), .Z(n18023) );
  NAND U18935 ( .A(n18024), .B(n18023), .Z(n18099) );
  XOR U18936 ( .A(n1053), .B(a[120]), .Z(n18182) );
  NANDN U18937 ( .A(n18182), .B(n37424), .Z(n18027) );
  NANDN U18938 ( .A(n18025), .B(n37425), .Z(n18026) );
  NAND U18939 ( .A(n18027), .B(n18026), .Z(n18098) );
  XOR U18940 ( .A(n18101), .B(n18100), .Z(n18095) );
  NANDN U18941 ( .A(n1049), .B(a[132]), .Z(n18028) );
  XNOR U18942 ( .A(b[1]), .B(n18028), .Z(n18030) );
  IV U18943 ( .A(a[131]), .Z(n22518) );
  NANDN U18944 ( .A(n22518), .B(n1049), .Z(n18029) );
  AND U18945 ( .A(n18030), .B(n18029), .Z(n18118) );
  NAND U18946 ( .A(n18031), .B(n38490), .Z(n18033) );
  XNOR U18947 ( .A(n1058), .B(a[104]), .Z(n18188) );
  NANDN U18948 ( .A(n1048), .B(n18188), .Z(n18032) );
  NAND U18949 ( .A(n18033), .B(n18032), .Z(n18116) );
  NANDN U18950 ( .A(n1059), .B(a[100]), .Z(n18117) );
  XNOR U18951 ( .A(n18116), .B(n18117), .Z(n18119) );
  XNOR U18952 ( .A(n18118), .B(n18119), .Z(n18093) );
  NANDN U18953 ( .A(n18034), .B(n38205), .Z(n18036) );
  XNOR U18954 ( .A(b[23]), .B(a[110]), .Z(n18191) );
  OR U18955 ( .A(n18191), .B(n38268), .Z(n18035) );
  NAND U18956 ( .A(n18036), .B(n18035), .Z(n18161) );
  XOR U18957 ( .A(b[7]), .B(a[126]), .Z(n18194) );
  NAND U18958 ( .A(n18194), .B(n36701), .Z(n18039) );
  NAND U18959 ( .A(n18037), .B(n36702), .Z(n18038) );
  NAND U18960 ( .A(n18039), .B(n18038), .Z(n18158) );
  XOR U18961 ( .A(b[25]), .B(a[108]), .Z(n18197) );
  NAND U18962 ( .A(n18197), .B(n38325), .Z(n18042) );
  NANDN U18963 ( .A(n18040), .B(n38326), .Z(n18041) );
  AND U18964 ( .A(n18042), .B(n18041), .Z(n18159) );
  XNOR U18965 ( .A(n18158), .B(n18159), .Z(n18160) );
  XOR U18966 ( .A(n18161), .B(n18160), .Z(n18092) );
  XOR U18967 ( .A(n18095), .B(n18094), .Z(n18149) );
  XNOR U18968 ( .A(n18148), .B(n18149), .Z(n18204) );
  XNOR U18969 ( .A(n18205), .B(n18204), .Z(n18207) );
  XNOR U18970 ( .A(n18206), .B(n18207), .Z(n18086) );
  XNOR U18971 ( .A(n18087), .B(n18086), .Z(n18088) );
  XOR U18972 ( .A(n18089), .B(n18088), .Z(n18083) );
  NANDN U18973 ( .A(n18044), .B(n18043), .Z(n18048) );
  NAND U18974 ( .A(n18046), .B(n18045), .Z(n18047) );
  NAND U18975 ( .A(n18048), .B(n18047), .Z(n18080) );
  NAND U18976 ( .A(n18050), .B(n18049), .Z(n18054) );
  NAND U18977 ( .A(n18052), .B(n18051), .Z(n18053) );
  NAND U18978 ( .A(n18054), .B(n18053), .Z(n18081) );
  XNOR U18979 ( .A(n18080), .B(n18081), .Z(n18082) );
  XNOR U18980 ( .A(n18083), .B(n18082), .Z(n18077) );
  NANDN U18981 ( .A(n18060), .B(n18059), .Z(n18064) );
  NANDN U18982 ( .A(n18062), .B(n18061), .Z(n18063) );
  NAND U18983 ( .A(n18064), .B(n18063), .Z(n18075) );
  XNOR U18984 ( .A(n18074), .B(n18075), .Z(n18076) );
  XNOR U18985 ( .A(n18077), .B(n18076), .Z(n18070) );
  XOR U18986 ( .A(n18071), .B(n18070), .Z(n18072) );
  XNOR U18987 ( .A(n18073), .B(n18072), .Z(n18210) );
  XNOR U18988 ( .A(n18210), .B(sreg[356]), .Z(n18212) );
  NAND U18989 ( .A(n18065), .B(sreg[355]), .Z(n18069) );
  OR U18990 ( .A(n18067), .B(n18066), .Z(n18068) );
  AND U18991 ( .A(n18069), .B(n18068), .Z(n18211) );
  XOR U18992 ( .A(n18212), .B(n18211), .Z(c[356]) );
  NANDN U18993 ( .A(n18075), .B(n18074), .Z(n18079) );
  NANDN U18994 ( .A(n18077), .B(n18076), .Z(n18078) );
  NAND U18995 ( .A(n18079), .B(n18078), .Z(n18216) );
  NANDN U18996 ( .A(n18081), .B(n18080), .Z(n18085) );
  NAND U18997 ( .A(n18083), .B(n18082), .Z(n18084) );
  NAND U18998 ( .A(n18085), .B(n18084), .Z(n18221) );
  NANDN U18999 ( .A(n18087), .B(n18086), .Z(n18091) );
  NANDN U19000 ( .A(n18089), .B(n18088), .Z(n18090) );
  NAND U19001 ( .A(n18091), .B(n18090), .Z(n18222) );
  XNOR U19002 ( .A(n18221), .B(n18222), .Z(n18223) );
  NANDN U19003 ( .A(n18093), .B(n18092), .Z(n18097) );
  NANDN U19004 ( .A(n18095), .B(n18094), .Z(n18096) );
  NAND U19005 ( .A(n18097), .B(n18096), .Z(n18336) );
  OR U19006 ( .A(n18099), .B(n18098), .Z(n18103) );
  NAND U19007 ( .A(n18101), .B(n18100), .Z(n18102) );
  NAND U19008 ( .A(n18103), .B(n18102), .Z(n18275) );
  OR U19009 ( .A(n18105), .B(n18104), .Z(n18109) );
  NANDN U19010 ( .A(n18107), .B(n18106), .Z(n18108) );
  NAND U19011 ( .A(n18109), .B(n18108), .Z(n18274) );
  OR U19012 ( .A(n18111), .B(n18110), .Z(n18115) );
  NANDN U19013 ( .A(n18113), .B(n18112), .Z(n18114) );
  NAND U19014 ( .A(n18115), .B(n18114), .Z(n18273) );
  XOR U19015 ( .A(n18275), .B(n18276), .Z(n18333) );
  NANDN U19016 ( .A(n18117), .B(n18116), .Z(n18121) );
  NAND U19017 ( .A(n18119), .B(n18118), .Z(n18120) );
  NAND U19018 ( .A(n18121), .B(n18120), .Z(n18288) );
  XNOR U19019 ( .A(b[19]), .B(a[115]), .Z(n18233) );
  NANDN U19020 ( .A(n18233), .B(n37934), .Z(n18124) );
  NANDN U19021 ( .A(n18122), .B(n37935), .Z(n18123) );
  NAND U19022 ( .A(n18124), .B(n18123), .Z(n18300) );
  XNOR U19023 ( .A(b[27]), .B(a[107]), .Z(n18236) );
  NANDN U19024 ( .A(n18236), .B(n38423), .Z(n18127) );
  NAND U19025 ( .A(n18125), .B(n38424), .Z(n18126) );
  NAND U19026 ( .A(n18127), .B(n18126), .Z(n18297) );
  XOR U19027 ( .A(b[5]), .B(n22221), .Z(n18239) );
  NANDN U19028 ( .A(n18239), .B(n36587), .Z(n18130) );
  NANDN U19029 ( .A(n18128), .B(n36588), .Z(n18129) );
  AND U19030 ( .A(n18130), .B(n18129), .Z(n18298) );
  XNOR U19031 ( .A(n18297), .B(n18298), .Z(n18299) );
  XNOR U19032 ( .A(n18300), .B(n18299), .Z(n18286) );
  NAND U19033 ( .A(n18131), .B(n37762), .Z(n18133) );
  XOR U19034 ( .A(b[17]), .B(a[117]), .Z(n18242) );
  NAND U19035 ( .A(n18242), .B(n37764), .Z(n18132) );
  NAND U19036 ( .A(n18133), .B(n18132), .Z(n18260) );
  XNOR U19037 ( .A(b[31]), .B(a[103]), .Z(n18245) );
  NANDN U19038 ( .A(n18245), .B(n38552), .Z(n18136) );
  NANDN U19039 ( .A(n18134), .B(n38553), .Z(n18135) );
  NAND U19040 ( .A(n18136), .B(n18135), .Z(n18257) );
  OR U19041 ( .A(n18137), .B(n36105), .Z(n18139) );
  XOR U19042 ( .A(b[3]), .B(n22518), .Z(n18248) );
  NANDN U19043 ( .A(n18248), .B(n36107), .Z(n18138) );
  AND U19044 ( .A(n18139), .B(n18138), .Z(n18258) );
  XNOR U19045 ( .A(n18257), .B(n18258), .Z(n18259) );
  XOR U19046 ( .A(n18260), .B(n18259), .Z(n18285) );
  XNOR U19047 ( .A(n18286), .B(n18285), .Z(n18287) );
  XNOR U19048 ( .A(n18288), .B(n18287), .Z(n18334) );
  XNOR U19049 ( .A(n18333), .B(n18334), .Z(n18335) );
  XNOR U19050 ( .A(n18336), .B(n18335), .Z(n18354) );
  OR U19051 ( .A(n18141), .B(n18140), .Z(n18145) );
  NANDN U19052 ( .A(n18143), .B(n18142), .Z(n18144) );
  NAND U19053 ( .A(n18145), .B(n18144), .Z(n18352) );
  NANDN U19054 ( .A(n18147), .B(n18146), .Z(n18151) );
  NANDN U19055 ( .A(n18149), .B(n18148), .Z(n18150) );
  NAND U19056 ( .A(n18151), .B(n18150), .Z(n18341) );
  OR U19057 ( .A(n18153), .B(n18152), .Z(n18157) );
  NANDN U19058 ( .A(n18155), .B(n18154), .Z(n18156) );
  NAND U19059 ( .A(n18157), .B(n18156), .Z(n18340) );
  NANDN U19060 ( .A(n18159), .B(n18158), .Z(n18163) );
  NAND U19061 ( .A(n18161), .B(n18160), .Z(n18162) );
  NAND U19062 ( .A(n18163), .B(n18162), .Z(n18279) );
  NANDN U19063 ( .A(n18165), .B(n18164), .Z(n18169) );
  NAND U19064 ( .A(n18167), .B(n18166), .Z(n18168) );
  AND U19065 ( .A(n18169), .B(n18168), .Z(n18280) );
  XNOR U19066 ( .A(n18279), .B(n18280), .Z(n18281) );
  XOR U19067 ( .A(n1052), .B(a[125]), .Z(n18309) );
  NANDN U19068 ( .A(n18309), .B(n36925), .Z(n18172) );
  NAND U19069 ( .A(n36926), .B(n18170), .Z(n18171) );
  NAND U19070 ( .A(n18172), .B(n18171), .Z(n18265) );
  XNOR U19071 ( .A(n1054), .B(a[119]), .Z(n18306) );
  NANDN U19072 ( .A(n37665), .B(n18306), .Z(n18175) );
  NANDN U19073 ( .A(n18173), .B(n37604), .Z(n18174) );
  NAND U19074 ( .A(n18175), .B(n18174), .Z(n18263) );
  XOR U19075 ( .A(n1056), .B(a[113]), .Z(n18303) );
  NANDN U19076 ( .A(n18303), .B(n38101), .Z(n18178) );
  NAND U19077 ( .A(n38102), .B(n18176), .Z(n18177) );
  NAND U19078 ( .A(n18178), .B(n18177), .Z(n18264) );
  XNOR U19079 ( .A(n18263), .B(n18264), .Z(n18266) );
  XOR U19080 ( .A(n18265), .B(n18266), .Z(n18254) );
  XNOR U19081 ( .A(b[11]), .B(a[123]), .Z(n18312) );
  OR U19082 ( .A(n18312), .B(n37311), .Z(n18181) );
  NANDN U19083 ( .A(n18179), .B(n37218), .Z(n18180) );
  NAND U19084 ( .A(n18181), .B(n18180), .Z(n18252) );
  XOR U19085 ( .A(n1053), .B(a[121]), .Z(n18315) );
  NANDN U19086 ( .A(n18315), .B(n37424), .Z(n18184) );
  NANDN U19087 ( .A(n18182), .B(n37425), .Z(n18183) );
  AND U19088 ( .A(n18184), .B(n18183), .Z(n18251) );
  XNOR U19089 ( .A(n18252), .B(n18251), .Z(n18253) );
  XNOR U19090 ( .A(n18254), .B(n18253), .Z(n18270) );
  NANDN U19091 ( .A(n1049), .B(a[133]), .Z(n18185) );
  XNOR U19092 ( .A(b[1]), .B(n18185), .Z(n18187) );
  NANDN U19093 ( .A(b[0]), .B(a[132]), .Z(n18186) );
  AND U19094 ( .A(n18187), .B(n18186), .Z(n18229) );
  NAND U19095 ( .A(n38490), .B(n18188), .Z(n18190) );
  XNOR U19096 ( .A(n1058), .B(a[105]), .Z(n18321) );
  NANDN U19097 ( .A(n1048), .B(n18321), .Z(n18189) );
  NAND U19098 ( .A(n18190), .B(n18189), .Z(n18227) );
  NANDN U19099 ( .A(n1059), .B(a[101]), .Z(n18228) );
  XNOR U19100 ( .A(n18227), .B(n18228), .Z(n18230) );
  XNOR U19101 ( .A(n18229), .B(n18230), .Z(n18268) );
  NANDN U19102 ( .A(n18191), .B(n38205), .Z(n18193) );
  XNOR U19103 ( .A(b[23]), .B(a[111]), .Z(n18324) );
  OR U19104 ( .A(n18324), .B(n38268), .Z(n18192) );
  NAND U19105 ( .A(n18193), .B(n18192), .Z(n18294) );
  XOR U19106 ( .A(b[7]), .B(a[127]), .Z(n18327) );
  NAND U19107 ( .A(n18327), .B(n36701), .Z(n18196) );
  NAND U19108 ( .A(n18194), .B(n36702), .Z(n18195) );
  NAND U19109 ( .A(n18196), .B(n18195), .Z(n18291) );
  XOR U19110 ( .A(b[25]), .B(a[109]), .Z(n18330) );
  NAND U19111 ( .A(n18330), .B(n38325), .Z(n18199) );
  NAND U19112 ( .A(n18197), .B(n38326), .Z(n18198) );
  AND U19113 ( .A(n18199), .B(n18198), .Z(n18292) );
  XNOR U19114 ( .A(n18291), .B(n18292), .Z(n18293) );
  XOR U19115 ( .A(n18294), .B(n18293), .Z(n18267) );
  XOR U19116 ( .A(n18270), .B(n18269), .Z(n18282) );
  XOR U19117 ( .A(n18281), .B(n18282), .Z(n18339) );
  XNOR U19118 ( .A(n18340), .B(n18339), .Z(n18342) );
  XNOR U19119 ( .A(n18341), .B(n18342), .Z(n18351) );
  XNOR U19120 ( .A(n18352), .B(n18351), .Z(n18353) );
  XOR U19121 ( .A(n18354), .B(n18353), .Z(n18348) );
  NAND U19122 ( .A(n18205), .B(n18204), .Z(n18209) );
  NANDN U19123 ( .A(n18207), .B(n18206), .Z(n18208) );
  AND U19124 ( .A(n18209), .B(n18208), .Z(n18345) );
  XNOR U19125 ( .A(n18346), .B(n18345), .Z(n18347) );
  XOR U19126 ( .A(n18348), .B(n18347), .Z(n18224) );
  XOR U19127 ( .A(n18223), .B(n18224), .Z(n18215) );
  XOR U19128 ( .A(n18216), .B(n18215), .Z(n18217) );
  XNOR U19129 ( .A(n18218), .B(n18217), .Z(n18357) );
  XNOR U19130 ( .A(n18357), .B(sreg[357]), .Z(n18359) );
  NAND U19131 ( .A(n18210), .B(sreg[356]), .Z(n18214) );
  OR U19132 ( .A(n18212), .B(n18211), .Z(n18213) );
  AND U19133 ( .A(n18214), .B(n18213), .Z(n18358) );
  XOR U19134 ( .A(n18359), .B(n18358), .Z(c[357]) );
  NAND U19135 ( .A(n18216), .B(n18215), .Z(n18220) );
  NAND U19136 ( .A(n18218), .B(n18217), .Z(n18219) );
  NAND U19137 ( .A(n18220), .B(n18219), .Z(n18365) );
  NANDN U19138 ( .A(n18222), .B(n18221), .Z(n18226) );
  NAND U19139 ( .A(n18224), .B(n18223), .Z(n18225) );
  NAND U19140 ( .A(n18226), .B(n18225), .Z(n18363) );
  NANDN U19141 ( .A(n18228), .B(n18227), .Z(n18232) );
  NAND U19142 ( .A(n18230), .B(n18229), .Z(n18231) );
  NAND U19143 ( .A(n18232), .B(n18231), .Z(n18443) );
  XNOR U19144 ( .A(b[19]), .B(a[116]), .Z(n18390) );
  NANDN U19145 ( .A(n18390), .B(n37934), .Z(n18235) );
  NANDN U19146 ( .A(n18233), .B(n37935), .Z(n18234) );
  NAND U19147 ( .A(n18235), .B(n18234), .Z(n18453) );
  XOR U19148 ( .A(b[27]), .B(a[108]), .Z(n18393) );
  NAND U19149 ( .A(n38423), .B(n18393), .Z(n18238) );
  NANDN U19150 ( .A(n18236), .B(n38424), .Z(n18237) );
  NAND U19151 ( .A(n18238), .B(n18237), .Z(n18450) );
  XNOR U19152 ( .A(b[5]), .B(a[130]), .Z(n18396) );
  NANDN U19153 ( .A(n18396), .B(n36587), .Z(n18241) );
  NANDN U19154 ( .A(n18239), .B(n36588), .Z(n18240) );
  AND U19155 ( .A(n18241), .B(n18240), .Z(n18451) );
  XNOR U19156 ( .A(n18450), .B(n18451), .Z(n18452) );
  XNOR U19157 ( .A(n18453), .B(n18452), .Z(n18441) );
  NAND U19158 ( .A(n18242), .B(n37762), .Z(n18244) );
  XNOR U19159 ( .A(b[17]), .B(a[118]), .Z(n18399) );
  NANDN U19160 ( .A(n18399), .B(n37764), .Z(n18243) );
  NAND U19161 ( .A(n18244), .B(n18243), .Z(n18417) );
  XNOR U19162 ( .A(b[31]), .B(a[104]), .Z(n18402) );
  NANDN U19163 ( .A(n18402), .B(n38552), .Z(n18247) );
  NANDN U19164 ( .A(n18245), .B(n38553), .Z(n18246) );
  NAND U19165 ( .A(n18247), .B(n18246), .Z(n18414) );
  OR U19166 ( .A(n18248), .B(n36105), .Z(n18250) );
  XNOR U19167 ( .A(b[3]), .B(a[132]), .Z(n18405) );
  NANDN U19168 ( .A(n18405), .B(n36107), .Z(n18249) );
  AND U19169 ( .A(n18250), .B(n18249), .Z(n18415) );
  XNOR U19170 ( .A(n18414), .B(n18415), .Z(n18416) );
  XOR U19171 ( .A(n18417), .B(n18416), .Z(n18440) );
  XNOR U19172 ( .A(n18441), .B(n18440), .Z(n18442) );
  XNOR U19173 ( .A(n18443), .B(n18442), .Z(n18381) );
  NANDN U19174 ( .A(n18252), .B(n18251), .Z(n18256) );
  NAND U19175 ( .A(n18254), .B(n18253), .Z(n18255) );
  NAND U19176 ( .A(n18256), .B(n18255), .Z(n18432) );
  NANDN U19177 ( .A(n18258), .B(n18257), .Z(n18262) );
  NAND U19178 ( .A(n18260), .B(n18259), .Z(n18261) );
  NAND U19179 ( .A(n18262), .B(n18261), .Z(n18431) );
  XNOR U19180 ( .A(n18431), .B(n18430), .Z(n18433) );
  XOR U19181 ( .A(n18432), .B(n18433), .Z(n18380) );
  XOR U19182 ( .A(n18381), .B(n18380), .Z(n18382) );
  NANDN U19183 ( .A(n18268), .B(n18267), .Z(n18272) );
  NAND U19184 ( .A(n18270), .B(n18269), .Z(n18271) );
  NAND U19185 ( .A(n18272), .B(n18271), .Z(n18383) );
  XNOR U19186 ( .A(n18382), .B(n18383), .Z(n18494) );
  OR U19187 ( .A(n18274), .B(n18273), .Z(n18278) );
  NANDN U19188 ( .A(n18276), .B(n18275), .Z(n18277) );
  NAND U19189 ( .A(n18278), .B(n18277), .Z(n18493) );
  NANDN U19190 ( .A(n18280), .B(n18279), .Z(n18284) );
  NAND U19191 ( .A(n18282), .B(n18281), .Z(n18283) );
  NAND U19192 ( .A(n18284), .B(n18283), .Z(n18376) );
  NANDN U19193 ( .A(n18286), .B(n18285), .Z(n18290) );
  NAND U19194 ( .A(n18288), .B(n18287), .Z(n18289) );
  NAND U19195 ( .A(n18290), .B(n18289), .Z(n18375) );
  NANDN U19196 ( .A(n18292), .B(n18291), .Z(n18296) );
  NAND U19197 ( .A(n18294), .B(n18293), .Z(n18295) );
  NAND U19198 ( .A(n18296), .B(n18295), .Z(n18434) );
  NANDN U19199 ( .A(n18298), .B(n18297), .Z(n18302) );
  NAND U19200 ( .A(n18300), .B(n18299), .Z(n18301) );
  AND U19201 ( .A(n18302), .B(n18301), .Z(n18435) );
  XNOR U19202 ( .A(n18434), .B(n18435), .Z(n18436) );
  XOR U19203 ( .A(n1056), .B(a[114]), .Z(n18462) );
  NANDN U19204 ( .A(n18462), .B(n38101), .Z(n18305) );
  NANDN U19205 ( .A(n18303), .B(n38102), .Z(n18304) );
  NAND U19206 ( .A(n18305), .B(n18304), .Z(n18426) );
  XNOR U19207 ( .A(b[15]), .B(a[120]), .Z(n18459) );
  OR U19208 ( .A(n18459), .B(n37665), .Z(n18308) );
  NAND U19209 ( .A(n18306), .B(n37604), .Z(n18307) );
  AND U19210 ( .A(n18308), .B(n18307), .Z(n18427) );
  XNOR U19211 ( .A(n18426), .B(n18427), .Z(n18429) );
  XOR U19212 ( .A(n1052), .B(a[126]), .Z(n18456) );
  NANDN U19213 ( .A(n18456), .B(n36925), .Z(n18311) );
  NANDN U19214 ( .A(n18309), .B(n36926), .Z(n18310) );
  NAND U19215 ( .A(n18311), .B(n18310), .Z(n18428) );
  XNOR U19216 ( .A(n18429), .B(n18428), .Z(n18422) );
  XNOR U19217 ( .A(b[11]), .B(a[124]), .Z(n18465) );
  OR U19218 ( .A(n18465), .B(n37311), .Z(n18314) );
  NANDN U19219 ( .A(n18312), .B(n37218), .Z(n18313) );
  NAND U19220 ( .A(n18314), .B(n18313), .Z(n18421) );
  XOR U19221 ( .A(n1053), .B(a[122]), .Z(n18468) );
  NANDN U19222 ( .A(n18468), .B(n37424), .Z(n18317) );
  NANDN U19223 ( .A(n18315), .B(n37425), .Z(n18316) );
  NAND U19224 ( .A(n18317), .B(n18316), .Z(n18420) );
  XNOR U19225 ( .A(n18421), .B(n18420), .Z(n18423) );
  XNOR U19226 ( .A(n18422), .B(n18423), .Z(n18411) );
  NANDN U19227 ( .A(n1049), .B(a[134]), .Z(n18318) );
  XNOR U19228 ( .A(b[1]), .B(n18318), .Z(n18320) );
  NANDN U19229 ( .A(b[0]), .B(a[133]), .Z(n18319) );
  AND U19230 ( .A(n18320), .B(n18319), .Z(n18386) );
  NAND U19231 ( .A(n38490), .B(n18321), .Z(n18323) );
  XNOR U19232 ( .A(n1058), .B(a[106]), .Z(n18471) );
  NANDN U19233 ( .A(n1048), .B(n18471), .Z(n18322) );
  NAND U19234 ( .A(n18323), .B(n18322), .Z(n18384) );
  NANDN U19235 ( .A(n1059), .B(a[102]), .Z(n18385) );
  XNOR U19236 ( .A(n18384), .B(n18385), .Z(n18387) );
  XNOR U19237 ( .A(n18386), .B(n18387), .Z(n18409) );
  NANDN U19238 ( .A(n18324), .B(n38205), .Z(n18326) );
  XNOR U19239 ( .A(b[23]), .B(a[112]), .Z(n18477) );
  OR U19240 ( .A(n18477), .B(n38268), .Z(n18325) );
  NAND U19241 ( .A(n18326), .B(n18325), .Z(n18447) );
  XOR U19242 ( .A(b[7]), .B(a[128]), .Z(n18480) );
  NAND U19243 ( .A(n18480), .B(n36701), .Z(n18329) );
  NAND U19244 ( .A(n18327), .B(n36702), .Z(n18328) );
  NAND U19245 ( .A(n18329), .B(n18328), .Z(n18444) );
  XOR U19246 ( .A(b[25]), .B(a[110]), .Z(n18483) );
  NAND U19247 ( .A(n18483), .B(n38325), .Z(n18332) );
  NAND U19248 ( .A(n18330), .B(n38326), .Z(n18331) );
  AND U19249 ( .A(n18332), .B(n18331), .Z(n18445) );
  XNOR U19250 ( .A(n18444), .B(n18445), .Z(n18446) );
  XOR U19251 ( .A(n18447), .B(n18446), .Z(n18408) );
  XOR U19252 ( .A(n18411), .B(n18410), .Z(n18437) );
  XNOR U19253 ( .A(n18436), .B(n18437), .Z(n18374) );
  XNOR U19254 ( .A(n18375), .B(n18374), .Z(n18377) );
  XNOR U19255 ( .A(n18376), .B(n18377), .Z(n18492) );
  XOR U19256 ( .A(n18493), .B(n18492), .Z(n18495) );
  NANDN U19257 ( .A(n18334), .B(n18333), .Z(n18338) );
  NAND U19258 ( .A(n18336), .B(n18335), .Z(n18337) );
  NAND U19259 ( .A(n18338), .B(n18337), .Z(n18487) );
  NAND U19260 ( .A(n18340), .B(n18339), .Z(n18344) );
  NANDN U19261 ( .A(n18342), .B(n18341), .Z(n18343) );
  AND U19262 ( .A(n18344), .B(n18343), .Z(n18486) );
  XNOR U19263 ( .A(n18487), .B(n18486), .Z(n18488) );
  XOR U19264 ( .A(n18489), .B(n18488), .Z(n18370) );
  NANDN U19265 ( .A(n18346), .B(n18345), .Z(n18350) );
  NAND U19266 ( .A(n18348), .B(n18347), .Z(n18349) );
  NAND U19267 ( .A(n18350), .B(n18349), .Z(n18368) );
  NANDN U19268 ( .A(n18352), .B(n18351), .Z(n18356) );
  NANDN U19269 ( .A(n18354), .B(n18353), .Z(n18355) );
  NAND U19270 ( .A(n18356), .B(n18355), .Z(n18369) );
  XNOR U19271 ( .A(n18368), .B(n18369), .Z(n18371) );
  XOR U19272 ( .A(n18370), .B(n18371), .Z(n18362) );
  XOR U19273 ( .A(n18363), .B(n18362), .Z(n18364) );
  XNOR U19274 ( .A(n18365), .B(n18364), .Z(n18498) );
  XNOR U19275 ( .A(n18498), .B(sreg[358]), .Z(n18500) );
  NAND U19276 ( .A(n18357), .B(sreg[357]), .Z(n18361) );
  OR U19277 ( .A(n18359), .B(n18358), .Z(n18360) );
  AND U19278 ( .A(n18361), .B(n18360), .Z(n18499) );
  XOR U19279 ( .A(n18500), .B(n18499), .Z(c[358]) );
  NAND U19280 ( .A(n18363), .B(n18362), .Z(n18367) );
  NAND U19281 ( .A(n18365), .B(n18364), .Z(n18366) );
  NAND U19282 ( .A(n18367), .B(n18366), .Z(n18506) );
  NANDN U19283 ( .A(n18369), .B(n18368), .Z(n18373) );
  NAND U19284 ( .A(n18371), .B(n18370), .Z(n18372) );
  NAND U19285 ( .A(n18373), .B(n18372), .Z(n18503) );
  NAND U19286 ( .A(n18375), .B(n18374), .Z(n18379) );
  NANDN U19287 ( .A(n18377), .B(n18376), .Z(n18378) );
  NAND U19288 ( .A(n18379), .B(n18378), .Z(n18629) );
  XNOR U19289 ( .A(n18629), .B(n18630), .Z(n18631) );
  NANDN U19290 ( .A(n18385), .B(n18384), .Z(n18389) );
  NAND U19291 ( .A(n18387), .B(n18386), .Z(n18388) );
  NAND U19292 ( .A(n18389), .B(n18388), .Z(n18574) );
  XNOR U19293 ( .A(b[19]), .B(a[117]), .Z(n18521) );
  NANDN U19294 ( .A(n18521), .B(n37934), .Z(n18392) );
  NANDN U19295 ( .A(n18390), .B(n37935), .Z(n18391) );
  NAND U19296 ( .A(n18392), .B(n18391), .Z(n18584) );
  XOR U19297 ( .A(b[27]), .B(a[109]), .Z(n18524) );
  NAND U19298 ( .A(n38423), .B(n18524), .Z(n18395) );
  NAND U19299 ( .A(n18393), .B(n38424), .Z(n18394) );
  NAND U19300 ( .A(n18395), .B(n18394), .Z(n18581) );
  XOR U19301 ( .A(b[5]), .B(n22518), .Z(n18527) );
  NANDN U19302 ( .A(n18527), .B(n36587), .Z(n18398) );
  NANDN U19303 ( .A(n18396), .B(n36588), .Z(n18397) );
  AND U19304 ( .A(n18398), .B(n18397), .Z(n18582) );
  XNOR U19305 ( .A(n18581), .B(n18582), .Z(n18583) );
  XNOR U19306 ( .A(n18584), .B(n18583), .Z(n18572) );
  NANDN U19307 ( .A(n18399), .B(n37762), .Z(n18401) );
  XOR U19308 ( .A(b[17]), .B(a[119]), .Z(n18530) );
  NAND U19309 ( .A(n18530), .B(n37764), .Z(n18400) );
  NAND U19310 ( .A(n18401), .B(n18400), .Z(n18548) );
  XNOR U19311 ( .A(b[31]), .B(a[105]), .Z(n18533) );
  NANDN U19312 ( .A(n18533), .B(n38552), .Z(n18404) );
  NANDN U19313 ( .A(n18402), .B(n38553), .Z(n18403) );
  NAND U19314 ( .A(n18404), .B(n18403), .Z(n18545) );
  OR U19315 ( .A(n18405), .B(n36105), .Z(n18407) );
  XNOR U19316 ( .A(b[3]), .B(a[133]), .Z(n18536) );
  NANDN U19317 ( .A(n18536), .B(n36107), .Z(n18406) );
  AND U19318 ( .A(n18407), .B(n18406), .Z(n18546) );
  XNOR U19319 ( .A(n18545), .B(n18546), .Z(n18547) );
  XOR U19320 ( .A(n18548), .B(n18547), .Z(n18571) );
  XNOR U19321 ( .A(n18572), .B(n18571), .Z(n18573) );
  XNOR U19322 ( .A(n18574), .B(n18573), .Z(n18623) );
  NANDN U19323 ( .A(n18409), .B(n18408), .Z(n18413) );
  NANDN U19324 ( .A(n18411), .B(n18410), .Z(n18412) );
  NAND U19325 ( .A(n18413), .B(n18412), .Z(n18624) );
  XNOR U19326 ( .A(n18623), .B(n18624), .Z(n18625) );
  NANDN U19327 ( .A(n18415), .B(n18414), .Z(n18419) );
  NAND U19328 ( .A(n18417), .B(n18416), .Z(n18418) );
  NAND U19329 ( .A(n18419), .B(n18418), .Z(n18564) );
  OR U19330 ( .A(n18421), .B(n18420), .Z(n18425) );
  NANDN U19331 ( .A(n18423), .B(n18422), .Z(n18424) );
  NAND U19332 ( .A(n18425), .B(n18424), .Z(n18562) );
  XNOR U19333 ( .A(n18562), .B(n18561), .Z(n18563) );
  XOR U19334 ( .A(n18564), .B(n18563), .Z(n18626) );
  XOR U19335 ( .A(n18625), .B(n18626), .Z(n18637) );
  NANDN U19336 ( .A(n18435), .B(n18434), .Z(n18439) );
  NANDN U19337 ( .A(n18437), .B(n18436), .Z(n18438) );
  NAND U19338 ( .A(n18439), .B(n18438), .Z(n18620) );
  NANDN U19339 ( .A(n18445), .B(n18444), .Z(n18449) );
  NAND U19340 ( .A(n18447), .B(n18446), .Z(n18448) );
  NAND U19341 ( .A(n18449), .B(n18448), .Z(n18565) );
  NANDN U19342 ( .A(n18451), .B(n18450), .Z(n18455) );
  NAND U19343 ( .A(n18453), .B(n18452), .Z(n18454) );
  AND U19344 ( .A(n18455), .B(n18454), .Z(n18566) );
  XNOR U19345 ( .A(n18565), .B(n18566), .Z(n18567) );
  XOR U19346 ( .A(n1052), .B(a[127]), .Z(n18587) );
  NANDN U19347 ( .A(n18587), .B(n36925), .Z(n18458) );
  NANDN U19348 ( .A(n18456), .B(n36926), .Z(n18457) );
  NAND U19349 ( .A(n18458), .B(n18457), .Z(n18553) );
  XNOR U19350 ( .A(b[15]), .B(a[121]), .Z(n18590) );
  OR U19351 ( .A(n18590), .B(n37665), .Z(n18461) );
  NANDN U19352 ( .A(n18459), .B(n37604), .Z(n18460) );
  NAND U19353 ( .A(n18461), .B(n18460), .Z(n18551) );
  XOR U19354 ( .A(n1056), .B(a[115]), .Z(n18593) );
  NANDN U19355 ( .A(n18593), .B(n38101), .Z(n18464) );
  NANDN U19356 ( .A(n18462), .B(n38102), .Z(n18463) );
  NAND U19357 ( .A(n18464), .B(n18463), .Z(n18552) );
  XNOR U19358 ( .A(n18551), .B(n18552), .Z(n18554) );
  XOR U19359 ( .A(n18553), .B(n18554), .Z(n18542) );
  XNOR U19360 ( .A(b[11]), .B(a[125]), .Z(n18596) );
  OR U19361 ( .A(n18596), .B(n37311), .Z(n18467) );
  NANDN U19362 ( .A(n18465), .B(n37218), .Z(n18466) );
  NAND U19363 ( .A(n18467), .B(n18466), .Z(n18540) );
  XOR U19364 ( .A(n1053), .B(a[123]), .Z(n18599) );
  NANDN U19365 ( .A(n18599), .B(n37424), .Z(n18470) );
  NANDN U19366 ( .A(n18468), .B(n37425), .Z(n18469) );
  AND U19367 ( .A(n18470), .B(n18469), .Z(n18539) );
  XNOR U19368 ( .A(n18540), .B(n18539), .Z(n18541) );
  XNOR U19369 ( .A(n18542), .B(n18541), .Z(n18558) );
  NAND U19370 ( .A(n38490), .B(n18471), .Z(n18473) );
  XOR U19371 ( .A(n1058), .B(n18980), .Z(n18605) );
  NANDN U19372 ( .A(n1048), .B(n18605), .Z(n18472) );
  NAND U19373 ( .A(n18473), .B(n18472), .Z(n18515) );
  NANDN U19374 ( .A(n1059), .B(a[103]), .Z(n18516) );
  XNOR U19375 ( .A(n18515), .B(n18516), .Z(n18518) );
  NANDN U19376 ( .A(n1049), .B(a[135]), .Z(n18474) );
  XNOR U19377 ( .A(b[1]), .B(n18474), .Z(n18476) );
  NANDN U19378 ( .A(b[0]), .B(a[134]), .Z(n18475) );
  AND U19379 ( .A(n18476), .B(n18475), .Z(n18517) );
  XNOR U19380 ( .A(n18518), .B(n18517), .Z(n18556) );
  NANDN U19381 ( .A(n18477), .B(n38205), .Z(n18479) );
  XOR U19382 ( .A(b[23]), .B(n19909), .Z(n18608) );
  OR U19383 ( .A(n18608), .B(n38268), .Z(n18478) );
  NAND U19384 ( .A(n18479), .B(n18478), .Z(n18578) );
  XNOR U19385 ( .A(b[7]), .B(a[129]), .Z(n18611) );
  NANDN U19386 ( .A(n18611), .B(n36701), .Z(n18482) );
  NAND U19387 ( .A(n18480), .B(n36702), .Z(n18481) );
  NAND U19388 ( .A(n18482), .B(n18481), .Z(n18575) );
  XOR U19389 ( .A(b[25]), .B(a[111]), .Z(n18614) );
  NAND U19390 ( .A(n18614), .B(n38325), .Z(n18485) );
  NAND U19391 ( .A(n18483), .B(n38326), .Z(n18484) );
  AND U19392 ( .A(n18485), .B(n18484), .Z(n18576) );
  XNOR U19393 ( .A(n18575), .B(n18576), .Z(n18577) );
  XOR U19394 ( .A(n18578), .B(n18577), .Z(n18555) );
  XOR U19395 ( .A(n18558), .B(n18557), .Z(n18568) );
  XOR U19396 ( .A(n18567), .B(n18568), .Z(n18617) );
  XOR U19397 ( .A(n18618), .B(n18617), .Z(n18619) );
  XNOR U19398 ( .A(n18620), .B(n18619), .Z(n18635) );
  XNOR U19399 ( .A(n18636), .B(n18635), .Z(n18638) );
  XNOR U19400 ( .A(n18637), .B(n18638), .Z(n18632) );
  XOR U19401 ( .A(n18631), .B(n18632), .Z(n18512) );
  NANDN U19402 ( .A(n18487), .B(n18486), .Z(n18491) );
  NAND U19403 ( .A(n18489), .B(n18488), .Z(n18490) );
  NAND U19404 ( .A(n18491), .B(n18490), .Z(n18509) );
  NANDN U19405 ( .A(n18493), .B(n18492), .Z(n18497) );
  OR U19406 ( .A(n18495), .B(n18494), .Z(n18496) );
  NAND U19407 ( .A(n18497), .B(n18496), .Z(n18510) );
  XNOR U19408 ( .A(n18509), .B(n18510), .Z(n18511) );
  XNOR U19409 ( .A(n18512), .B(n18511), .Z(n18504) );
  XNOR U19410 ( .A(n18503), .B(n18504), .Z(n18505) );
  XNOR U19411 ( .A(n18506), .B(n18505), .Z(n18641) );
  XNOR U19412 ( .A(n18641), .B(sreg[359]), .Z(n18643) );
  NAND U19413 ( .A(n18498), .B(sreg[358]), .Z(n18502) );
  OR U19414 ( .A(n18500), .B(n18499), .Z(n18501) );
  AND U19415 ( .A(n18502), .B(n18501), .Z(n18642) );
  XOR U19416 ( .A(n18643), .B(n18642), .Z(c[359]) );
  NANDN U19417 ( .A(n18504), .B(n18503), .Z(n18508) );
  NAND U19418 ( .A(n18506), .B(n18505), .Z(n18507) );
  NAND U19419 ( .A(n18508), .B(n18507), .Z(n18649) );
  NANDN U19420 ( .A(n18510), .B(n18509), .Z(n18514) );
  NAND U19421 ( .A(n18512), .B(n18511), .Z(n18513) );
  NAND U19422 ( .A(n18514), .B(n18513), .Z(n18647) );
  NANDN U19423 ( .A(n18516), .B(n18515), .Z(n18520) );
  NAND U19424 ( .A(n18518), .B(n18517), .Z(n18519) );
  NAND U19425 ( .A(n18520), .B(n18519), .Z(n18725) );
  XOR U19426 ( .A(b[19]), .B(n20271), .Z(n18672) );
  NANDN U19427 ( .A(n18672), .B(n37934), .Z(n18523) );
  NANDN U19428 ( .A(n18521), .B(n37935), .Z(n18522) );
  NAND U19429 ( .A(n18523), .B(n18522), .Z(n18735) );
  XOR U19430 ( .A(b[27]), .B(a[110]), .Z(n18675) );
  NAND U19431 ( .A(n38423), .B(n18675), .Z(n18526) );
  NAND U19432 ( .A(n18524), .B(n38424), .Z(n18525) );
  NAND U19433 ( .A(n18526), .B(n18525), .Z(n18732) );
  XNOR U19434 ( .A(b[5]), .B(a[132]), .Z(n18678) );
  NANDN U19435 ( .A(n18678), .B(n36587), .Z(n18529) );
  NANDN U19436 ( .A(n18527), .B(n36588), .Z(n18528) );
  AND U19437 ( .A(n18529), .B(n18528), .Z(n18733) );
  XNOR U19438 ( .A(n18732), .B(n18733), .Z(n18734) );
  XNOR U19439 ( .A(n18735), .B(n18734), .Z(n18723) );
  NAND U19440 ( .A(n18530), .B(n37762), .Z(n18532) );
  XOR U19441 ( .A(b[17]), .B(a[120]), .Z(n18681) );
  NAND U19442 ( .A(n18681), .B(n37764), .Z(n18531) );
  NAND U19443 ( .A(n18532), .B(n18531), .Z(n18699) );
  XNOR U19444 ( .A(b[31]), .B(a[106]), .Z(n18684) );
  NANDN U19445 ( .A(n18684), .B(n38552), .Z(n18535) );
  NANDN U19446 ( .A(n18533), .B(n38553), .Z(n18534) );
  NAND U19447 ( .A(n18535), .B(n18534), .Z(n18696) );
  OR U19448 ( .A(n18536), .B(n36105), .Z(n18538) );
  XNOR U19449 ( .A(b[3]), .B(a[134]), .Z(n18687) );
  NANDN U19450 ( .A(n18687), .B(n36107), .Z(n18537) );
  AND U19451 ( .A(n18538), .B(n18537), .Z(n18697) );
  XNOR U19452 ( .A(n18696), .B(n18697), .Z(n18698) );
  XOR U19453 ( .A(n18699), .B(n18698), .Z(n18722) );
  XNOR U19454 ( .A(n18723), .B(n18722), .Z(n18724) );
  XNOR U19455 ( .A(n18725), .B(n18724), .Z(n18663) );
  NANDN U19456 ( .A(n18540), .B(n18539), .Z(n18544) );
  NAND U19457 ( .A(n18542), .B(n18541), .Z(n18543) );
  NAND U19458 ( .A(n18544), .B(n18543), .Z(n18714) );
  NANDN U19459 ( .A(n18546), .B(n18545), .Z(n18550) );
  NAND U19460 ( .A(n18548), .B(n18547), .Z(n18549) );
  NAND U19461 ( .A(n18550), .B(n18549), .Z(n18713) );
  XNOR U19462 ( .A(n18713), .B(n18712), .Z(n18715) );
  XOR U19463 ( .A(n18714), .B(n18715), .Z(n18662) );
  XOR U19464 ( .A(n18663), .B(n18662), .Z(n18664) );
  NANDN U19465 ( .A(n18556), .B(n18555), .Z(n18560) );
  NAND U19466 ( .A(n18558), .B(n18557), .Z(n18559) );
  AND U19467 ( .A(n18560), .B(n18559), .Z(n18665) );
  XNOR U19468 ( .A(n18664), .B(n18665), .Z(n18771) );
  NANDN U19469 ( .A(n18566), .B(n18565), .Z(n18570) );
  NAND U19470 ( .A(n18568), .B(n18567), .Z(n18569) );
  NAND U19471 ( .A(n18570), .B(n18569), .Z(n18659) );
  NANDN U19472 ( .A(n18576), .B(n18575), .Z(n18580) );
  NAND U19473 ( .A(n18578), .B(n18577), .Z(n18579) );
  NAND U19474 ( .A(n18580), .B(n18579), .Z(n18716) );
  NANDN U19475 ( .A(n18582), .B(n18581), .Z(n18586) );
  NAND U19476 ( .A(n18584), .B(n18583), .Z(n18585) );
  AND U19477 ( .A(n18586), .B(n18585), .Z(n18717) );
  XNOR U19478 ( .A(n18716), .B(n18717), .Z(n18718) );
  XOR U19479 ( .A(n1052), .B(a[128]), .Z(n18744) );
  NANDN U19480 ( .A(n18744), .B(n36925), .Z(n18589) );
  NANDN U19481 ( .A(n18587), .B(n36926), .Z(n18588) );
  NAND U19482 ( .A(n18589), .B(n18588), .Z(n18704) );
  XNOR U19483 ( .A(n1054), .B(a[122]), .Z(n18741) );
  NANDN U19484 ( .A(n37665), .B(n18741), .Z(n18592) );
  NANDN U19485 ( .A(n18590), .B(n37604), .Z(n18591) );
  NAND U19486 ( .A(n18592), .B(n18591), .Z(n18702) );
  XOR U19487 ( .A(n1056), .B(a[116]), .Z(n18738) );
  NANDN U19488 ( .A(n18738), .B(n38101), .Z(n18595) );
  NANDN U19489 ( .A(n18593), .B(n38102), .Z(n18594) );
  NAND U19490 ( .A(n18595), .B(n18594), .Z(n18703) );
  XNOR U19491 ( .A(n18702), .B(n18703), .Z(n18705) );
  XOR U19492 ( .A(n18704), .B(n18705), .Z(n18693) );
  XNOR U19493 ( .A(b[11]), .B(a[126]), .Z(n18747) );
  OR U19494 ( .A(n18747), .B(n37311), .Z(n18598) );
  NANDN U19495 ( .A(n18596), .B(n37218), .Z(n18597) );
  NAND U19496 ( .A(n18598), .B(n18597), .Z(n18691) );
  XOR U19497 ( .A(n1053), .B(a[124]), .Z(n18750) );
  NANDN U19498 ( .A(n18750), .B(n37424), .Z(n18601) );
  NANDN U19499 ( .A(n18599), .B(n37425), .Z(n18600) );
  AND U19500 ( .A(n18601), .B(n18600), .Z(n18690) );
  XNOR U19501 ( .A(n18691), .B(n18690), .Z(n18692) );
  XNOR U19502 ( .A(n18693), .B(n18692), .Z(n18709) );
  NANDN U19503 ( .A(n1049), .B(a[136]), .Z(n18602) );
  XNOR U19504 ( .A(b[1]), .B(n18602), .Z(n18604) );
  NANDN U19505 ( .A(b[0]), .B(a[135]), .Z(n18603) );
  AND U19506 ( .A(n18604), .B(n18603), .Z(n18668) );
  NAND U19507 ( .A(n38490), .B(n18605), .Z(n18607) );
  XNOR U19508 ( .A(n1058), .B(a[108]), .Z(n18756) );
  NANDN U19509 ( .A(n1048), .B(n18756), .Z(n18606) );
  NAND U19510 ( .A(n18607), .B(n18606), .Z(n18666) );
  NANDN U19511 ( .A(n1059), .B(a[104]), .Z(n18667) );
  XNOR U19512 ( .A(n18666), .B(n18667), .Z(n18669) );
  XNOR U19513 ( .A(n18668), .B(n18669), .Z(n18707) );
  NANDN U19514 ( .A(n18608), .B(n38205), .Z(n18610) );
  XNOR U19515 ( .A(b[23]), .B(a[114]), .Z(n18759) );
  OR U19516 ( .A(n18759), .B(n38268), .Z(n18609) );
  NAND U19517 ( .A(n18610), .B(n18609), .Z(n18729) );
  XOR U19518 ( .A(b[7]), .B(a[130]), .Z(n18762) );
  NAND U19519 ( .A(n18762), .B(n36701), .Z(n18613) );
  NANDN U19520 ( .A(n18611), .B(n36702), .Z(n18612) );
  NAND U19521 ( .A(n18613), .B(n18612), .Z(n18726) );
  XOR U19522 ( .A(b[25]), .B(a[112]), .Z(n18765) );
  NAND U19523 ( .A(n18765), .B(n38325), .Z(n18616) );
  NAND U19524 ( .A(n18614), .B(n38326), .Z(n18615) );
  AND U19525 ( .A(n18616), .B(n18615), .Z(n18727) );
  XNOR U19526 ( .A(n18726), .B(n18727), .Z(n18728) );
  XOR U19527 ( .A(n18729), .B(n18728), .Z(n18706) );
  XOR U19528 ( .A(n18709), .B(n18708), .Z(n18719) );
  XOR U19529 ( .A(n18718), .B(n18719), .Z(n18656) );
  XOR U19530 ( .A(n18657), .B(n18656), .Z(n18658) );
  XOR U19531 ( .A(n18659), .B(n18658), .Z(n18769) );
  XNOR U19532 ( .A(n18768), .B(n18769), .Z(n18770) );
  XNOR U19533 ( .A(n18771), .B(n18770), .Z(n18775) );
  NAND U19534 ( .A(n18618), .B(n18617), .Z(n18622) );
  NAND U19535 ( .A(n18620), .B(n18619), .Z(n18621) );
  NAND U19536 ( .A(n18622), .B(n18621), .Z(n18772) );
  NANDN U19537 ( .A(n18624), .B(n18623), .Z(n18628) );
  NAND U19538 ( .A(n18626), .B(n18625), .Z(n18627) );
  NAND U19539 ( .A(n18628), .B(n18627), .Z(n18773) );
  XNOR U19540 ( .A(n18772), .B(n18773), .Z(n18774) );
  XNOR U19541 ( .A(n18775), .B(n18774), .Z(n18653) );
  NANDN U19542 ( .A(n18630), .B(n18629), .Z(n18634) );
  NANDN U19543 ( .A(n18632), .B(n18631), .Z(n18633) );
  NAND U19544 ( .A(n18634), .B(n18633), .Z(n18651) );
  OR U19545 ( .A(n18636), .B(n18635), .Z(n18640) );
  OR U19546 ( .A(n18638), .B(n18637), .Z(n18639) );
  AND U19547 ( .A(n18640), .B(n18639), .Z(n18650) );
  XNOR U19548 ( .A(n18651), .B(n18650), .Z(n18652) );
  XNOR U19549 ( .A(n18653), .B(n18652), .Z(n18646) );
  XOR U19550 ( .A(n18647), .B(n18646), .Z(n18648) );
  XNOR U19551 ( .A(n18649), .B(n18648), .Z(n18778) );
  XNOR U19552 ( .A(n18778), .B(sreg[360]), .Z(n18780) );
  NAND U19553 ( .A(n18641), .B(sreg[359]), .Z(n18645) );
  OR U19554 ( .A(n18643), .B(n18642), .Z(n18644) );
  AND U19555 ( .A(n18645), .B(n18644), .Z(n18779) );
  XOR U19556 ( .A(n18780), .B(n18779), .Z(c[360]) );
  NANDN U19557 ( .A(n18651), .B(n18650), .Z(n18655) );
  NANDN U19558 ( .A(n18653), .B(n18652), .Z(n18654) );
  NAND U19559 ( .A(n18655), .B(n18654), .Z(n18783) );
  NAND U19560 ( .A(n18657), .B(n18656), .Z(n18661) );
  NAND U19561 ( .A(n18659), .B(n18658), .Z(n18660) );
  NAND U19562 ( .A(n18661), .B(n18660), .Z(n18907) );
  XNOR U19563 ( .A(n18907), .B(n18908), .Z(n18909) );
  NANDN U19564 ( .A(n18667), .B(n18666), .Z(n18671) );
  NAND U19565 ( .A(n18669), .B(n18668), .Z(n18670) );
  NAND U19566 ( .A(n18671), .B(n18670), .Z(n18864) );
  XNOR U19567 ( .A(b[19]), .B(a[119]), .Z(n18811) );
  NANDN U19568 ( .A(n18811), .B(n37934), .Z(n18674) );
  NANDN U19569 ( .A(n18672), .B(n37935), .Z(n18673) );
  NAND U19570 ( .A(n18674), .B(n18673), .Z(n18874) );
  XOR U19571 ( .A(b[27]), .B(a[111]), .Z(n18814) );
  NAND U19572 ( .A(n38423), .B(n18814), .Z(n18677) );
  NAND U19573 ( .A(n18675), .B(n38424), .Z(n18676) );
  NAND U19574 ( .A(n18677), .B(n18676), .Z(n18871) );
  XNOR U19575 ( .A(b[5]), .B(a[133]), .Z(n18817) );
  NANDN U19576 ( .A(n18817), .B(n36587), .Z(n18680) );
  NANDN U19577 ( .A(n18678), .B(n36588), .Z(n18679) );
  AND U19578 ( .A(n18680), .B(n18679), .Z(n18872) );
  XNOR U19579 ( .A(n18871), .B(n18872), .Z(n18873) );
  XNOR U19580 ( .A(n18874), .B(n18873), .Z(n18862) );
  NAND U19581 ( .A(n18681), .B(n37762), .Z(n18683) );
  XOR U19582 ( .A(b[17]), .B(a[121]), .Z(n18820) );
  NAND U19583 ( .A(n18820), .B(n37764), .Z(n18682) );
  NAND U19584 ( .A(n18683), .B(n18682), .Z(n18838) );
  XOR U19585 ( .A(b[31]), .B(n18980), .Z(n18823) );
  NANDN U19586 ( .A(n18823), .B(n38552), .Z(n18686) );
  NANDN U19587 ( .A(n18684), .B(n38553), .Z(n18685) );
  NAND U19588 ( .A(n18686), .B(n18685), .Z(n18835) );
  OR U19589 ( .A(n18687), .B(n36105), .Z(n18689) );
  XNOR U19590 ( .A(b[3]), .B(a[135]), .Z(n18826) );
  NANDN U19591 ( .A(n18826), .B(n36107), .Z(n18688) );
  AND U19592 ( .A(n18689), .B(n18688), .Z(n18836) );
  XNOR U19593 ( .A(n18835), .B(n18836), .Z(n18837) );
  XOR U19594 ( .A(n18838), .B(n18837), .Z(n18861) );
  XNOR U19595 ( .A(n18862), .B(n18861), .Z(n18863) );
  XNOR U19596 ( .A(n18864), .B(n18863), .Z(n18802) );
  NANDN U19597 ( .A(n18691), .B(n18690), .Z(n18695) );
  NAND U19598 ( .A(n18693), .B(n18692), .Z(n18694) );
  NAND U19599 ( .A(n18695), .B(n18694), .Z(n18853) );
  NANDN U19600 ( .A(n18697), .B(n18696), .Z(n18701) );
  NAND U19601 ( .A(n18699), .B(n18698), .Z(n18700) );
  NAND U19602 ( .A(n18701), .B(n18700), .Z(n18852) );
  XNOR U19603 ( .A(n18852), .B(n18851), .Z(n18854) );
  XOR U19604 ( .A(n18853), .B(n18854), .Z(n18801) );
  XOR U19605 ( .A(n18802), .B(n18801), .Z(n18803) );
  NANDN U19606 ( .A(n18707), .B(n18706), .Z(n18711) );
  NAND U19607 ( .A(n18709), .B(n18708), .Z(n18710) );
  AND U19608 ( .A(n18711), .B(n18710), .Z(n18804) );
  XOR U19609 ( .A(n18803), .B(n18804), .Z(n18915) );
  NANDN U19610 ( .A(n18717), .B(n18716), .Z(n18721) );
  NAND U19611 ( .A(n18719), .B(n18718), .Z(n18720) );
  NAND U19612 ( .A(n18721), .B(n18720), .Z(n18798) );
  NANDN U19613 ( .A(n18727), .B(n18726), .Z(n18731) );
  NAND U19614 ( .A(n18729), .B(n18728), .Z(n18730) );
  NAND U19615 ( .A(n18731), .B(n18730), .Z(n18855) );
  NANDN U19616 ( .A(n18733), .B(n18732), .Z(n18737) );
  NAND U19617 ( .A(n18735), .B(n18734), .Z(n18736) );
  AND U19618 ( .A(n18737), .B(n18736), .Z(n18856) );
  XNOR U19619 ( .A(n18855), .B(n18856), .Z(n18857) );
  XNOR U19620 ( .A(b[21]), .B(a[117]), .Z(n18883) );
  NANDN U19621 ( .A(n18883), .B(n38101), .Z(n18740) );
  NANDN U19622 ( .A(n18738), .B(n38102), .Z(n18739) );
  NAND U19623 ( .A(n18740), .B(n18739), .Z(n18847) );
  XNOR U19624 ( .A(b[15]), .B(a[123]), .Z(n18880) );
  OR U19625 ( .A(n18880), .B(n37665), .Z(n18743) );
  NAND U19626 ( .A(n18741), .B(n37604), .Z(n18742) );
  AND U19627 ( .A(n18743), .B(n18742), .Z(n18848) );
  XNOR U19628 ( .A(n18847), .B(n18848), .Z(n18850) );
  XOR U19629 ( .A(b[9]), .B(n22221), .Z(n18877) );
  NANDN U19630 ( .A(n18877), .B(n36925), .Z(n18746) );
  NANDN U19631 ( .A(n18744), .B(n36926), .Z(n18745) );
  NAND U19632 ( .A(n18746), .B(n18745), .Z(n18849) );
  XNOR U19633 ( .A(n18850), .B(n18849), .Z(n18843) );
  XNOR U19634 ( .A(b[11]), .B(a[127]), .Z(n18886) );
  OR U19635 ( .A(n18886), .B(n37311), .Z(n18749) );
  NANDN U19636 ( .A(n18747), .B(n37218), .Z(n18748) );
  NAND U19637 ( .A(n18749), .B(n18748), .Z(n18842) );
  XOR U19638 ( .A(n1053), .B(a[125]), .Z(n18889) );
  NANDN U19639 ( .A(n18889), .B(n37424), .Z(n18752) );
  NANDN U19640 ( .A(n18750), .B(n37425), .Z(n18751) );
  NAND U19641 ( .A(n18752), .B(n18751), .Z(n18841) );
  XNOR U19642 ( .A(n18842), .B(n18841), .Z(n18844) );
  XNOR U19643 ( .A(n18843), .B(n18844), .Z(n18832) );
  NANDN U19644 ( .A(n1049), .B(a[137]), .Z(n18753) );
  XNOR U19645 ( .A(b[1]), .B(n18753), .Z(n18755) );
  NANDN U19646 ( .A(b[0]), .B(a[136]), .Z(n18754) );
  AND U19647 ( .A(n18755), .B(n18754), .Z(n18807) );
  NAND U19648 ( .A(n38490), .B(n18756), .Z(n18758) );
  XNOR U19649 ( .A(n1058), .B(a[109]), .Z(n18892) );
  NANDN U19650 ( .A(n1048), .B(n18892), .Z(n18757) );
  NAND U19651 ( .A(n18758), .B(n18757), .Z(n18805) );
  NANDN U19652 ( .A(n1059), .B(a[105]), .Z(n18806) );
  XNOR U19653 ( .A(n18805), .B(n18806), .Z(n18808) );
  XNOR U19654 ( .A(n18807), .B(n18808), .Z(n18830) );
  NANDN U19655 ( .A(n18759), .B(n38205), .Z(n18761) );
  XNOR U19656 ( .A(b[23]), .B(a[115]), .Z(n18898) );
  OR U19657 ( .A(n18898), .B(n38268), .Z(n18760) );
  NAND U19658 ( .A(n18761), .B(n18760), .Z(n18868) );
  XNOR U19659 ( .A(b[7]), .B(a[131]), .Z(n18901) );
  NANDN U19660 ( .A(n18901), .B(n36701), .Z(n18764) );
  NAND U19661 ( .A(n18762), .B(n36702), .Z(n18763) );
  NAND U19662 ( .A(n18764), .B(n18763), .Z(n18865) );
  XNOR U19663 ( .A(b[25]), .B(a[113]), .Z(n18904) );
  NANDN U19664 ( .A(n18904), .B(n38325), .Z(n18767) );
  NAND U19665 ( .A(n18765), .B(n38326), .Z(n18766) );
  AND U19666 ( .A(n18767), .B(n18766), .Z(n18866) );
  XNOR U19667 ( .A(n18865), .B(n18866), .Z(n18867) );
  XOR U19668 ( .A(n18868), .B(n18867), .Z(n18829) );
  XOR U19669 ( .A(n18832), .B(n18831), .Z(n18858) );
  XNOR U19670 ( .A(n18857), .B(n18858), .Z(n18795) );
  XOR U19671 ( .A(n18796), .B(n18795), .Z(n18797) );
  XNOR U19672 ( .A(n18798), .B(n18797), .Z(n18913) );
  XNOR U19673 ( .A(n18914), .B(n18913), .Z(n18916) );
  XNOR U19674 ( .A(n18915), .B(n18916), .Z(n18910) );
  XOR U19675 ( .A(n18909), .B(n18910), .Z(n18792) );
  NANDN U19676 ( .A(n18773), .B(n18772), .Z(n18777) );
  NANDN U19677 ( .A(n18775), .B(n18774), .Z(n18776) );
  NAND U19678 ( .A(n18777), .B(n18776), .Z(n18790) );
  XNOR U19679 ( .A(n18789), .B(n18790), .Z(n18791) );
  XNOR U19680 ( .A(n18792), .B(n18791), .Z(n18784) );
  XNOR U19681 ( .A(n18783), .B(n18784), .Z(n18785) );
  XNOR U19682 ( .A(n18786), .B(n18785), .Z(n18919) );
  XNOR U19683 ( .A(n18919), .B(sreg[361]), .Z(n18921) );
  NAND U19684 ( .A(n18778), .B(sreg[360]), .Z(n18782) );
  OR U19685 ( .A(n18780), .B(n18779), .Z(n18781) );
  AND U19686 ( .A(n18782), .B(n18781), .Z(n18920) );
  XOR U19687 ( .A(n18921), .B(n18920), .Z(c[361]) );
  NANDN U19688 ( .A(n18784), .B(n18783), .Z(n18788) );
  NAND U19689 ( .A(n18786), .B(n18785), .Z(n18787) );
  NAND U19690 ( .A(n18788), .B(n18787), .Z(n18927) );
  NANDN U19691 ( .A(n18790), .B(n18789), .Z(n18794) );
  NAND U19692 ( .A(n18792), .B(n18791), .Z(n18793) );
  NAND U19693 ( .A(n18794), .B(n18793), .Z(n18924) );
  NAND U19694 ( .A(n18796), .B(n18795), .Z(n18800) );
  NAND U19695 ( .A(n18798), .B(n18797), .Z(n18799) );
  NAND U19696 ( .A(n18800), .B(n18799), .Z(n19053) );
  XNOR U19697 ( .A(n19053), .B(n19054), .Z(n19055) );
  NANDN U19698 ( .A(n18806), .B(n18805), .Z(n18810) );
  NAND U19699 ( .A(n18808), .B(n18807), .Z(n18809) );
  NAND U19700 ( .A(n18810), .B(n18809), .Z(n18949) );
  XNOR U19701 ( .A(b[19]), .B(a[120]), .Z(n18999) );
  NANDN U19702 ( .A(n18999), .B(n37934), .Z(n18813) );
  NANDN U19703 ( .A(n18811), .B(n37935), .Z(n18812) );
  NAND U19704 ( .A(n18813), .B(n18812), .Z(n18959) );
  XOR U19705 ( .A(b[27]), .B(a[112]), .Z(n19002) );
  NAND U19706 ( .A(n38423), .B(n19002), .Z(n18816) );
  NAND U19707 ( .A(n18814), .B(n38424), .Z(n18815) );
  NAND U19708 ( .A(n18816), .B(n18815), .Z(n18956) );
  XNOR U19709 ( .A(b[5]), .B(a[134]), .Z(n19005) );
  NANDN U19710 ( .A(n19005), .B(n36587), .Z(n18819) );
  NANDN U19711 ( .A(n18817), .B(n36588), .Z(n18818) );
  AND U19712 ( .A(n18819), .B(n18818), .Z(n18957) );
  XNOR U19713 ( .A(n18956), .B(n18957), .Z(n18958) );
  XNOR U19714 ( .A(n18959), .B(n18958), .Z(n18947) );
  NAND U19715 ( .A(n18820), .B(n37762), .Z(n18822) );
  XOR U19716 ( .A(b[17]), .B(a[122]), .Z(n19008) );
  NAND U19717 ( .A(n19008), .B(n37764), .Z(n18821) );
  NAND U19718 ( .A(n18822), .B(n18821), .Z(n19026) );
  XNOR U19719 ( .A(b[31]), .B(a[108]), .Z(n19011) );
  NANDN U19720 ( .A(n19011), .B(n38552), .Z(n18825) );
  NANDN U19721 ( .A(n18823), .B(n38553), .Z(n18824) );
  NAND U19722 ( .A(n18825), .B(n18824), .Z(n19023) );
  OR U19723 ( .A(n18826), .B(n36105), .Z(n18828) );
  XNOR U19724 ( .A(b[3]), .B(a[136]), .Z(n19014) );
  NANDN U19725 ( .A(n19014), .B(n36107), .Z(n18827) );
  AND U19726 ( .A(n18828), .B(n18827), .Z(n19024) );
  XNOR U19727 ( .A(n19023), .B(n19024), .Z(n19025) );
  XOR U19728 ( .A(n19026), .B(n19025), .Z(n18946) );
  XNOR U19729 ( .A(n18947), .B(n18946), .Z(n18948) );
  XNOR U19730 ( .A(n18949), .B(n18948), .Z(n19047) );
  NANDN U19731 ( .A(n18830), .B(n18829), .Z(n18834) );
  NANDN U19732 ( .A(n18832), .B(n18831), .Z(n18833) );
  NAND U19733 ( .A(n18834), .B(n18833), .Z(n19048) );
  XNOR U19734 ( .A(n19047), .B(n19048), .Z(n19049) );
  NANDN U19735 ( .A(n18836), .B(n18835), .Z(n18840) );
  NAND U19736 ( .A(n18838), .B(n18837), .Z(n18839) );
  NAND U19737 ( .A(n18840), .B(n18839), .Z(n18939) );
  OR U19738 ( .A(n18842), .B(n18841), .Z(n18846) );
  NANDN U19739 ( .A(n18844), .B(n18843), .Z(n18845) );
  NAND U19740 ( .A(n18846), .B(n18845), .Z(n18937) );
  XNOR U19741 ( .A(n18937), .B(n18936), .Z(n18938) );
  XOR U19742 ( .A(n18939), .B(n18938), .Z(n19050) );
  XOR U19743 ( .A(n19049), .B(n19050), .Z(n19061) );
  NANDN U19744 ( .A(n18856), .B(n18855), .Z(n18860) );
  NANDN U19745 ( .A(n18858), .B(n18857), .Z(n18859) );
  NAND U19746 ( .A(n18860), .B(n18859), .Z(n19044) );
  NANDN U19747 ( .A(n18866), .B(n18865), .Z(n18870) );
  NAND U19748 ( .A(n18868), .B(n18867), .Z(n18869) );
  NAND U19749 ( .A(n18870), .B(n18869), .Z(n18940) );
  NANDN U19750 ( .A(n18872), .B(n18871), .Z(n18876) );
  NAND U19751 ( .A(n18874), .B(n18873), .Z(n18875) );
  AND U19752 ( .A(n18876), .B(n18875), .Z(n18941) );
  XNOR U19753 ( .A(n18940), .B(n18941), .Z(n18942) );
  XNOR U19754 ( .A(b[9]), .B(a[130]), .Z(n18962) );
  NANDN U19755 ( .A(n18962), .B(n36925), .Z(n18879) );
  NANDN U19756 ( .A(n18877), .B(n36926), .Z(n18878) );
  NAND U19757 ( .A(n18879), .B(n18878), .Z(n19037) );
  XNOR U19758 ( .A(b[15]), .B(a[124]), .Z(n18965) );
  OR U19759 ( .A(n18965), .B(n37665), .Z(n18882) );
  NANDN U19760 ( .A(n18880), .B(n37604), .Z(n18881) );
  AND U19761 ( .A(n18882), .B(n18881), .Z(n19035) );
  XOR U19762 ( .A(b[21]), .B(n20271), .Z(n18968) );
  NANDN U19763 ( .A(n18968), .B(n38101), .Z(n18885) );
  NANDN U19764 ( .A(n18883), .B(n38102), .Z(n18884) );
  AND U19765 ( .A(n18885), .B(n18884), .Z(n19036) );
  XOR U19766 ( .A(n19037), .B(n19038), .Z(n19032) );
  XNOR U19767 ( .A(b[11]), .B(a[128]), .Z(n18971) );
  OR U19768 ( .A(n18971), .B(n37311), .Z(n18888) );
  NANDN U19769 ( .A(n18886), .B(n37218), .Z(n18887) );
  NAND U19770 ( .A(n18888), .B(n18887), .Z(n19030) );
  XOR U19771 ( .A(n1053), .B(a[126]), .Z(n18974) );
  NANDN U19772 ( .A(n18974), .B(n37424), .Z(n18891) );
  NANDN U19773 ( .A(n18889), .B(n37425), .Z(n18890) );
  AND U19774 ( .A(n18891), .B(n18890), .Z(n19029) );
  XNOR U19775 ( .A(n19030), .B(n19029), .Z(n19031) );
  XOR U19776 ( .A(n19032), .B(n19031), .Z(n19019) );
  NAND U19777 ( .A(n38490), .B(n18892), .Z(n18894) );
  XNOR U19778 ( .A(b[29]), .B(a[110]), .Z(n18981) );
  OR U19779 ( .A(n18981), .B(n1048), .Z(n18893) );
  NAND U19780 ( .A(n18894), .B(n18893), .Z(n18993) );
  NANDN U19781 ( .A(n1059), .B(a[106]), .Z(n18994) );
  XNOR U19782 ( .A(n18993), .B(n18994), .Z(n18996) );
  NANDN U19783 ( .A(n1049), .B(a[138]), .Z(n18895) );
  XNOR U19784 ( .A(b[1]), .B(n18895), .Z(n18897) );
  IV U19785 ( .A(a[137]), .Z(n23393) );
  NANDN U19786 ( .A(n23393), .B(n1049), .Z(n18896) );
  AND U19787 ( .A(n18897), .B(n18896), .Z(n18995) );
  XOR U19788 ( .A(n18996), .B(n18995), .Z(n19017) );
  NANDN U19789 ( .A(n18898), .B(n38205), .Z(n18900) );
  XNOR U19790 ( .A(b[23]), .B(a[116]), .Z(n18984) );
  OR U19791 ( .A(n18984), .B(n38268), .Z(n18899) );
  NAND U19792 ( .A(n18900), .B(n18899), .Z(n18953) );
  XOR U19793 ( .A(b[7]), .B(a[132]), .Z(n18987) );
  NAND U19794 ( .A(n18987), .B(n36701), .Z(n18903) );
  NANDN U19795 ( .A(n18901), .B(n36702), .Z(n18902) );
  NAND U19796 ( .A(n18903), .B(n18902), .Z(n18950) );
  XOR U19797 ( .A(b[25]), .B(a[114]), .Z(n18990) );
  NAND U19798 ( .A(n18990), .B(n38325), .Z(n18906) );
  NANDN U19799 ( .A(n18904), .B(n38326), .Z(n18905) );
  AND U19800 ( .A(n18906), .B(n18905), .Z(n18951) );
  XNOR U19801 ( .A(n18950), .B(n18951), .Z(n18952) );
  XNOR U19802 ( .A(n18953), .B(n18952), .Z(n19018) );
  XOR U19803 ( .A(n19017), .B(n19018), .Z(n19020) );
  XNOR U19804 ( .A(n19019), .B(n19020), .Z(n18943) );
  XOR U19805 ( .A(n18942), .B(n18943), .Z(n19042) );
  XNOR U19806 ( .A(n19041), .B(n19042), .Z(n19043) );
  XNOR U19807 ( .A(n19044), .B(n19043), .Z(n19059) );
  XNOR U19808 ( .A(n19060), .B(n19059), .Z(n19062) );
  XNOR U19809 ( .A(n19061), .B(n19062), .Z(n19056) );
  XOR U19810 ( .A(n19055), .B(n19056), .Z(n18933) );
  NANDN U19811 ( .A(n18908), .B(n18907), .Z(n18912) );
  NANDN U19812 ( .A(n18910), .B(n18909), .Z(n18911) );
  NAND U19813 ( .A(n18912), .B(n18911), .Z(n18931) );
  OR U19814 ( .A(n18914), .B(n18913), .Z(n18918) );
  OR U19815 ( .A(n18916), .B(n18915), .Z(n18917) );
  AND U19816 ( .A(n18918), .B(n18917), .Z(n18930) );
  XNOR U19817 ( .A(n18931), .B(n18930), .Z(n18932) );
  XNOR U19818 ( .A(n18933), .B(n18932), .Z(n18925) );
  XNOR U19819 ( .A(n18924), .B(n18925), .Z(n18926) );
  XNOR U19820 ( .A(n18927), .B(n18926), .Z(n19065) );
  XNOR U19821 ( .A(n19065), .B(sreg[362]), .Z(n19067) );
  NAND U19822 ( .A(n18919), .B(sreg[361]), .Z(n18923) );
  OR U19823 ( .A(n18921), .B(n18920), .Z(n18922) );
  AND U19824 ( .A(n18923), .B(n18922), .Z(n19066) );
  XOR U19825 ( .A(n19067), .B(n19066), .Z(c[362]) );
  NANDN U19826 ( .A(n18925), .B(n18924), .Z(n18929) );
  NAND U19827 ( .A(n18927), .B(n18926), .Z(n18928) );
  NAND U19828 ( .A(n18929), .B(n18928), .Z(n19073) );
  NANDN U19829 ( .A(n18931), .B(n18930), .Z(n18935) );
  NAND U19830 ( .A(n18933), .B(n18932), .Z(n18934) );
  NAND U19831 ( .A(n18935), .B(n18934), .Z(n19071) );
  NANDN U19832 ( .A(n18941), .B(n18940), .Z(n18945) );
  NANDN U19833 ( .A(n18943), .B(n18942), .Z(n18944) );
  NAND U19834 ( .A(n18945), .B(n18944), .Z(n19087) );
  NANDN U19835 ( .A(n18951), .B(n18950), .Z(n18955) );
  NAND U19836 ( .A(n18953), .B(n18952), .Z(n18954) );
  NAND U19837 ( .A(n18955), .B(n18954), .Z(n19144) );
  NANDN U19838 ( .A(n18957), .B(n18956), .Z(n18961) );
  NAND U19839 ( .A(n18959), .B(n18958), .Z(n18960) );
  AND U19840 ( .A(n18961), .B(n18960), .Z(n19145) );
  XNOR U19841 ( .A(n19144), .B(n19145), .Z(n19146) );
  XOR U19842 ( .A(b[9]), .B(n22518), .Z(n19168) );
  NANDN U19843 ( .A(n19168), .B(n36925), .Z(n18964) );
  NANDN U19844 ( .A(n18962), .B(n36926), .Z(n18963) );
  NAND U19845 ( .A(n18964), .B(n18963), .Z(n19110) );
  XNOR U19846 ( .A(b[15]), .B(a[125]), .Z(n19171) );
  OR U19847 ( .A(n19171), .B(n37665), .Z(n18967) );
  NANDN U19848 ( .A(n18965), .B(n37604), .Z(n18966) );
  AND U19849 ( .A(n18967), .B(n18966), .Z(n19108) );
  XNOR U19850 ( .A(b[21]), .B(a[119]), .Z(n19174) );
  NANDN U19851 ( .A(n19174), .B(n38101), .Z(n18970) );
  NANDN U19852 ( .A(n18968), .B(n38102), .Z(n18969) );
  AND U19853 ( .A(n18970), .B(n18969), .Z(n19109) );
  XOR U19854 ( .A(n19110), .B(n19111), .Z(n19099) );
  XOR U19855 ( .A(b[11]), .B(n22221), .Z(n19177) );
  OR U19856 ( .A(n19177), .B(n37311), .Z(n18973) );
  NANDN U19857 ( .A(n18971), .B(n37218), .Z(n18972) );
  NAND U19858 ( .A(n18973), .B(n18972), .Z(n19097) );
  XOR U19859 ( .A(n1053), .B(a[127]), .Z(n19180) );
  NANDN U19860 ( .A(n19180), .B(n37424), .Z(n18976) );
  NANDN U19861 ( .A(n18974), .B(n37425), .Z(n18975) );
  NAND U19862 ( .A(n18976), .B(n18975), .Z(n19096) );
  XOR U19863 ( .A(n19099), .B(n19098), .Z(n19093) );
  NANDN U19864 ( .A(n1049), .B(a[139]), .Z(n18977) );
  XNOR U19865 ( .A(b[1]), .B(n18977), .Z(n18979) );
  NANDN U19866 ( .A(b[0]), .B(a[138]), .Z(n18978) );
  AND U19867 ( .A(n18979), .B(n18978), .Z(n19117) );
  ANDN U19868 ( .B(b[31]), .A(n18980), .Z(n19114) );
  NANDN U19869 ( .A(n18981), .B(n38490), .Z(n18983) );
  XNOR U19870 ( .A(n1058), .B(a[111]), .Z(n19186) );
  NANDN U19871 ( .A(n1048), .B(n19186), .Z(n18982) );
  NAND U19872 ( .A(n18983), .B(n18982), .Z(n19115) );
  XOR U19873 ( .A(n19114), .B(n19115), .Z(n19116) );
  XNOR U19874 ( .A(n19117), .B(n19116), .Z(n19090) );
  NANDN U19875 ( .A(n18984), .B(n38205), .Z(n18986) );
  XNOR U19876 ( .A(b[23]), .B(a[117]), .Z(n19189) );
  OR U19877 ( .A(n19189), .B(n38268), .Z(n18985) );
  NAND U19878 ( .A(n18986), .B(n18985), .Z(n19159) );
  XOR U19879 ( .A(b[7]), .B(a[133]), .Z(n19192) );
  NAND U19880 ( .A(n19192), .B(n36701), .Z(n18989) );
  NAND U19881 ( .A(n18987), .B(n36702), .Z(n18988) );
  NAND U19882 ( .A(n18989), .B(n18988), .Z(n19156) );
  XOR U19883 ( .A(b[25]), .B(a[115]), .Z(n19195) );
  NAND U19884 ( .A(n19195), .B(n38325), .Z(n18992) );
  NAND U19885 ( .A(n18990), .B(n38326), .Z(n18991) );
  AND U19886 ( .A(n18992), .B(n18991), .Z(n19157) );
  XNOR U19887 ( .A(n19156), .B(n19157), .Z(n19158) );
  XNOR U19888 ( .A(n19159), .B(n19158), .Z(n19091) );
  XOR U19889 ( .A(n19093), .B(n19092), .Z(n19147) );
  XNOR U19890 ( .A(n19146), .B(n19147), .Z(n19084) );
  XOR U19891 ( .A(n19085), .B(n19084), .Z(n19086) );
  XOR U19892 ( .A(n19087), .B(n19086), .Z(n19199) );
  XNOR U19893 ( .A(n19198), .B(n19199), .Z(n19201) );
  NANDN U19894 ( .A(n18994), .B(n18993), .Z(n18998) );
  NAND U19895 ( .A(n18996), .B(n18995), .Z(n18997) );
  NAND U19896 ( .A(n18998), .B(n18997), .Z(n19153) );
  XNOR U19897 ( .A(b[19]), .B(a[121]), .Z(n19120) );
  NANDN U19898 ( .A(n19120), .B(n37934), .Z(n19001) );
  NANDN U19899 ( .A(n18999), .B(n37935), .Z(n19000) );
  NAND U19900 ( .A(n19001), .B(n19000), .Z(n19165) );
  XNOR U19901 ( .A(b[27]), .B(a[113]), .Z(n19123) );
  NANDN U19902 ( .A(n19123), .B(n38423), .Z(n19004) );
  NAND U19903 ( .A(n19002), .B(n38424), .Z(n19003) );
  NAND U19904 ( .A(n19004), .B(n19003), .Z(n19162) );
  XNOR U19905 ( .A(b[5]), .B(a[135]), .Z(n19126) );
  NANDN U19906 ( .A(n19126), .B(n36587), .Z(n19007) );
  NANDN U19907 ( .A(n19005), .B(n36588), .Z(n19006) );
  AND U19908 ( .A(n19007), .B(n19006), .Z(n19163) );
  XNOR U19909 ( .A(n19162), .B(n19163), .Z(n19164) );
  XNOR U19910 ( .A(n19165), .B(n19164), .Z(n19150) );
  NAND U19911 ( .A(n19008), .B(n37762), .Z(n19010) );
  XOR U19912 ( .A(b[17]), .B(a[123]), .Z(n19129) );
  NAND U19913 ( .A(n19129), .B(n37764), .Z(n19009) );
  NAND U19914 ( .A(n19010), .B(n19009), .Z(n19104) );
  XNOR U19915 ( .A(b[31]), .B(a[109]), .Z(n19132) );
  NANDN U19916 ( .A(n19132), .B(n38552), .Z(n19013) );
  NANDN U19917 ( .A(n19011), .B(n38553), .Z(n19012) );
  AND U19918 ( .A(n19013), .B(n19012), .Z(n19102) );
  OR U19919 ( .A(n19014), .B(n36105), .Z(n19016) );
  XOR U19920 ( .A(b[3]), .B(n23393), .Z(n19135) );
  NANDN U19921 ( .A(n19135), .B(n36107), .Z(n19015) );
  AND U19922 ( .A(n19016), .B(n19015), .Z(n19103) );
  XOR U19923 ( .A(n19104), .B(n19105), .Z(n19151) );
  XOR U19924 ( .A(n19150), .B(n19151), .Z(n19152) );
  XNOR U19925 ( .A(n19153), .B(n19152), .Z(n19080) );
  NANDN U19926 ( .A(n19018), .B(n19017), .Z(n19022) );
  OR U19927 ( .A(n19020), .B(n19019), .Z(n19021) );
  NAND U19928 ( .A(n19022), .B(n19021), .Z(n19081) );
  XNOR U19929 ( .A(n19080), .B(n19081), .Z(n19082) );
  NANDN U19930 ( .A(n19024), .B(n19023), .Z(n19028) );
  NAND U19931 ( .A(n19026), .B(n19025), .Z(n19027) );
  NAND U19932 ( .A(n19028), .B(n19027), .Z(n19141) );
  NANDN U19933 ( .A(n19030), .B(n19029), .Z(n19034) );
  NAND U19934 ( .A(n19032), .B(n19031), .Z(n19033) );
  NAND U19935 ( .A(n19034), .B(n19033), .Z(n19138) );
  OR U19936 ( .A(n19036), .B(n19035), .Z(n19040) );
  NANDN U19937 ( .A(n19038), .B(n19037), .Z(n19039) );
  NAND U19938 ( .A(n19040), .B(n19039), .Z(n19139) );
  XNOR U19939 ( .A(n19138), .B(n19139), .Z(n19140) );
  XOR U19940 ( .A(n19141), .B(n19140), .Z(n19083) );
  XNOR U19941 ( .A(n19082), .B(n19083), .Z(n19200) );
  XOR U19942 ( .A(n19201), .B(n19200), .Z(n19205) );
  NANDN U19943 ( .A(n19042), .B(n19041), .Z(n19046) );
  NAND U19944 ( .A(n19044), .B(n19043), .Z(n19045) );
  NAND U19945 ( .A(n19046), .B(n19045), .Z(n19202) );
  NANDN U19946 ( .A(n19048), .B(n19047), .Z(n19052) );
  NAND U19947 ( .A(n19050), .B(n19049), .Z(n19051) );
  NAND U19948 ( .A(n19052), .B(n19051), .Z(n19203) );
  XNOR U19949 ( .A(n19202), .B(n19203), .Z(n19204) );
  XNOR U19950 ( .A(n19205), .B(n19204), .Z(n19077) );
  NANDN U19951 ( .A(n19054), .B(n19053), .Z(n19058) );
  NANDN U19952 ( .A(n19056), .B(n19055), .Z(n19057) );
  NAND U19953 ( .A(n19058), .B(n19057), .Z(n19075) );
  OR U19954 ( .A(n19060), .B(n19059), .Z(n19064) );
  OR U19955 ( .A(n19062), .B(n19061), .Z(n19063) );
  AND U19956 ( .A(n19064), .B(n19063), .Z(n19074) );
  XNOR U19957 ( .A(n19075), .B(n19074), .Z(n19076) );
  XNOR U19958 ( .A(n19077), .B(n19076), .Z(n19070) );
  XOR U19959 ( .A(n19071), .B(n19070), .Z(n19072) );
  XNOR U19960 ( .A(n19073), .B(n19072), .Z(n19208) );
  XNOR U19961 ( .A(n19208), .B(sreg[363]), .Z(n19210) );
  NAND U19962 ( .A(n19065), .B(sreg[362]), .Z(n19069) );
  OR U19963 ( .A(n19067), .B(n19066), .Z(n19068) );
  AND U19964 ( .A(n19069), .B(n19068), .Z(n19209) );
  XOR U19965 ( .A(n19210), .B(n19209), .Z(c[363]) );
  NANDN U19966 ( .A(n19075), .B(n19074), .Z(n19079) );
  NANDN U19967 ( .A(n19077), .B(n19076), .Z(n19078) );
  NAND U19968 ( .A(n19079), .B(n19078), .Z(n19214) );
  NAND U19969 ( .A(n19085), .B(n19084), .Z(n19089) );
  NAND U19970 ( .A(n19087), .B(n19086), .Z(n19088) );
  NAND U19971 ( .A(n19089), .B(n19088), .Z(n19232) );
  XNOR U19972 ( .A(n19231), .B(n19232), .Z(n19233) );
  OR U19973 ( .A(n19091), .B(n19090), .Z(n19095) );
  NANDN U19974 ( .A(n19093), .B(n19092), .Z(n19094) );
  NAND U19975 ( .A(n19095), .B(n19094), .Z(n19348) );
  OR U19976 ( .A(n19097), .B(n19096), .Z(n19101) );
  NAND U19977 ( .A(n19099), .B(n19098), .Z(n19100) );
  NAND U19978 ( .A(n19101), .B(n19100), .Z(n19287) );
  OR U19979 ( .A(n19103), .B(n19102), .Z(n19107) );
  NANDN U19980 ( .A(n19105), .B(n19104), .Z(n19106) );
  NAND U19981 ( .A(n19107), .B(n19106), .Z(n19286) );
  OR U19982 ( .A(n19109), .B(n19108), .Z(n19113) );
  NANDN U19983 ( .A(n19111), .B(n19110), .Z(n19112) );
  NAND U19984 ( .A(n19113), .B(n19112), .Z(n19285) );
  XOR U19985 ( .A(n19287), .B(n19288), .Z(n19346) );
  OR U19986 ( .A(n19115), .B(n19114), .Z(n19119) );
  NANDN U19987 ( .A(n19117), .B(n19116), .Z(n19118) );
  NAND U19988 ( .A(n19119), .B(n19118), .Z(n19299) );
  XNOR U19989 ( .A(b[19]), .B(a[122]), .Z(n19243) );
  NANDN U19990 ( .A(n19243), .B(n37934), .Z(n19122) );
  NANDN U19991 ( .A(n19120), .B(n37935), .Z(n19121) );
  NAND U19992 ( .A(n19122), .B(n19121), .Z(n19312) );
  XOR U19993 ( .A(b[27]), .B(a[114]), .Z(n19246) );
  NAND U19994 ( .A(n38423), .B(n19246), .Z(n19125) );
  NANDN U19995 ( .A(n19123), .B(n38424), .Z(n19124) );
  NAND U19996 ( .A(n19125), .B(n19124), .Z(n19309) );
  XNOR U19997 ( .A(b[5]), .B(a[136]), .Z(n19249) );
  NANDN U19998 ( .A(n19249), .B(n36587), .Z(n19128) );
  NANDN U19999 ( .A(n19126), .B(n36588), .Z(n19127) );
  AND U20000 ( .A(n19128), .B(n19127), .Z(n19310) );
  XNOR U20001 ( .A(n19309), .B(n19310), .Z(n19311) );
  XNOR U20002 ( .A(n19312), .B(n19311), .Z(n19298) );
  NAND U20003 ( .A(n19129), .B(n37762), .Z(n19131) );
  XOR U20004 ( .A(b[17]), .B(a[124]), .Z(n19252) );
  NAND U20005 ( .A(n19252), .B(n37764), .Z(n19130) );
  NAND U20006 ( .A(n19131), .B(n19130), .Z(n19270) );
  XNOR U20007 ( .A(b[31]), .B(a[110]), .Z(n19255) );
  NANDN U20008 ( .A(n19255), .B(n38552), .Z(n19134) );
  NANDN U20009 ( .A(n19132), .B(n38553), .Z(n19133) );
  NAND U20010 ( .A(n19134), .B(n19133), .Z(n19267) );
  OR U20011 ( .A(n19135), .B(n36105), .Z(n19137) );
  XNOR U20012 ( .A(b[3]), .B(a[138]), .Z(n19258) );
  NANDN U20013 ( .A(n19258), .B(n36107), .Z(n19136) );
  AND U20014 ( .A(n19137), .B(n19136), .Z(n19268) );
  XNOR U20015 ( .A(n19267), .B(n19268), .Z(n19269) );
  XOR U20016 ( .A(n19270), .B(n19269), .Z(n19297) );
  XOR U20017 ( .A(n19298), .B(n19297), .Z(n19300) );
  XOR U20018 ( .A(n19299), .B(n19300), .Z(n19345) );
  XOR U20019 ( .A(n19346), .B(n19345), .Z(n19347) );
  XNOR U20020 ( .A(n19348), .B(n19347), .Z(n19228) );
  NANDN U20021 ( .A(n19139), .B(n19138), .Z(n19143) );
  NANDN U20022 ( .A(n19141), .B(n19140), .Z(n19142) );
  NAND U20023 ( .A(n19143), .B(n19142), .Z(n19225) );
  NANDN U20024 ( .A(n19145), .B(n19144), .Z(n19149) );
  NANDN U20025 ( .A(n19147), .B(n19146), .Z(n19148) );
  NAND U20026 ( .A(n19149), .B(n19148), .Z(n19354) );
  OR U20027 ( .A(n19151), .B(n19150), .Z(n19155) );
  NAND U20028 ( .A(n19153), .B(n19152), .Z(n19154) );
  NAND U20029 ( .A(n19155), .B(n19154), .Z(n19351) );
  NANDN U20030 ( .A(n19157), .B(n19156), .Z(n19161) );
  NAND U20031 ( .A(n19159), .B(n19158), .Z(n19160) );
  NAND U20032 ( .A(n19161), .B(n19160), .Z(n19291) );
  NANDN U20033 ( .A(n19163), .B(n19162), .Z(n19167) );
  NAND U20034 ( .A(n19165), .B(n19164), .Z(n19166) );
  AND U20035 ( .A(n19167), .B(n19166), .Z(n19292) );
  XNOR U20036 ( .A(n19291), .B(n19292), .Z(n19293) );
  XNOR U20037 ( .A(b[9]), .B(a[132]), .Z(n19315) );
  NANDN U20038 ( .A(n19315), .B(n36925), .Z(n19170) );
  NANDN U20039 ( .A(n19168), .B(n36926), .Z(n19169) );
  NAND U20040 ( .A(n19170), .B(n19169), .Z(n19275) );
  XNOR U20041 ( .A(b[15]), .B(a[126]), .Z(n19318) );
  OR U20042 ( .A(n19318), .B(n37665), .Z(n19173) );
  NANDN U20043 ( .A(n19171), .B(n37604), .Z(n19172) );
  AND U20044 ( .A(n19173), .B(n19172), .Z(n19273) );
  XNOR U20045 ( .A(b[21]), .B(a[120]), .Z(n19321) );
  NANDN U20046 ( .A(n19321), .B(n38101), .Z(n19176) );
  NANDN U20047 ( .A(n19174), .B(n38102), .Z(n19175) );
  AND U20048 ( .A(n19176), .B(n19175), .Z(n19274) );
  XOR U20049 ( .A(n19275), .B(n19276), .Z(n19264) );
  XNOR U20050 ( .A(b[11]), .B(a[130]), .Z(n19324) );
  OR U20051 ( .A(n19324), .B(n37311), .Z(n19179) );
  NANDN U20052 ( .A(n19177), .B(n37218), .Z(n19178) );
  NAND U20053 ( .A(n19179), .B(n19178), .Z(n19262) );
  XOR U20054 ( .A(n1053), .B(a[128]), .Z(n19327) );
  NANDN U20055 ( .A(n19327), .B(n37424), .Z(n19182) );
  NANDN U20056 ( .A(n19180), .B(n37425), .Z(n19181) );
  AND U20057 ( .A(n19182), .B(n19181), .Z(n19261) );
  XNOR U20058 ( .A(n19262), .B(n19261), .Z(n19263) );
  XOR U20059 ( .A(n19264), .B(n19263), .Z(n19281) );
  NANDN U20060 ( .A(n1049), .B(a[140]), .Z(n19183) );
  XNOR U20061 ( .A(b[1]), .B(n19183), .Z(n19185) );
  IV U20062 ( .A(a[139]), .Z(n23668) );
  NANDN U20063 ( .A(n23668), .B(n1049), .Z(n19184) );
  AND U20064 ( .A(n19185), .B(n19184), .Z(n19239) );
  NAND U20065 ( .A(n19186), .B(n38490), .Z(n19188) );
  XNOR U20066 ( .A(n1058), .B(a[112]), .Z(n19330) );
  NANDN U20067 ( .A(n1048), .B(n19330), .Z(n19187) );
  NAND U20068 ( .A(n19188), .B(n19187), .Z(n19237) );
  NANDN U20069 ( .A(n1059), .B(a[108]), .Z(n19238) );
  XNOR U20070 ( .A(n19237), .B(n19238), .Z(n19240) );
  XOR U20071 ( .A(n19239), .B(n19240), .Z(n19279) );
  NANDN U20072 ( .A(n19189), .B(n38205), .Z(n19191) );
  XOR U20073 ( .A(b[23]), .B(n20271), .Z(n19336) );
  OR U20074 ( .A(n19336), .B(n38268), .Z(n19190) );
  NAND U20075 ( .A(n19191), .B(n19190), .Z(n19306) );
  XOR U20076 ( .A(b[7]), .B(a[134]), .Z(n19339) );
  NAND U20077 ( .A(n19339), .B(n36701), .Z(n19194) );
  NAND U20078 ( .A(n19192), .B(n36702), .Z(n19193) );
  NAND U20079 ( .A(n19194), .B(n19193), .Z(n19303) );
  XOR U20080 ( .A(b[25]), .B(a[116]), .Z(n19342) );
  NAND U20081 ( .A(n19342), .B(n38325), .Z(n19197) );
  NAND U20082 ( .A(n19195), .B(n38326), .Z(n19196) );
  AND U20083 ( .A(n19197), .B(n19196), .Z(n19304) );
  XNOR U20084 ( .A(n19303), .B(n19304), .Z(n19305) );
  XNOR U20085 ( .A(n19306), .B(n19305), .Z(n19280) );
  XOR U20086 ( .A(n19279), .B(n19280), .Z(n19282) );
  XNOR U20087 ( .A(n19281), .B(n19282), .Z(n19294) );
  XOR U20088 ( .A(n19293), .B(n19294), .Z(n19352) );
  XNOR U20089 ( .A(n19351), .B(n19352), .Z(n19353) );
  XOR U20090 ( .A(n19354), .B(n19353), .Z(n19226) );
  XNOR U20091 ( .A(n19225), .B(n19226), .Z(n19227) );
  XOR U20092 ( .A(n19228), .B(n19227), .Z(n19234) );
  XOR U20093 ( .A(n19233), .B(n19234), .Z(n19221) );
  NANDN U20094 ( .A(n19203), .B(n19202), .Z(n19207) );
  NANDN U20095 ( .A(n19205), .B(n19204), .Z(n19206) );
  NAND U20096 ( .A(n19207), .B(n19206), .Z(n19220) );
  XNOR U20097 ( .A(n19219), .B(n19220), .Z(n19222) );
  XOR U20098 ( .A(n19221), .B(n19222), .Z(n19213) );
  XOR U20099 ( .A(n19214), .B(n19213), .Z(n19215) );
  XNOR U20100 ( .A(n19216), .B(n19215), .Z(n19357) );
  XNOR U20101 ( .A(n19357), .B(sreg[364]), .Z(n19359) );
  NAND U20102 ( .A(n19208), .B(sreg[363]), .Z(n19212) );
  OR U20103 ( .A(n19210), .B(n19209), .Z(n19211) );
  AND U20104 ( .A(n19212), .B(n19211), .Z(n19358) );
  XOR U20105 ( .A(n19359), .B(n19358), .Z(c[364]) );
  NAND U20106 ( .A(n19214), .B(n19213), .Z(n19218) );
  NAND U20107 ( .A(n19216), .B(n19215), .Z(n19217) );
  NAND U20108 ( .A(n19218), .B(n19217), .Z(n19365) );
  NANDN U20109 ( .A(n19220), .B(n19219), .Z(n19224) );
  NAND U20110 ( .A(n19222), .B(n19221), .Z(n19223) );
  NAND U20111 ( .A(n19224), .B(n19223), .Z(n19363) );
  NANDN U20112 ( .A(n19226), .B(n19225), .Z(n19230) );
  NAND U20113 ( .A(n19228), .B(n19227), .Z(n19229) );
  NAND U20114 ( .A(n19230), .B(n19229), .Z(n19368) );
  NANDN U20115 ( .A(n19232), .B(n19231), .Z(n19236) );
  NAND U20116 ( .A(n19234), .B(n19233), .Z(n19235) );
  AND U20117 ( .A(n19236), .B(n19235), .Z(n19369) );
  XNOR U20118 ( .A(n19368), .B(n19369), .Z(n19370) );
  NANDN U20119 ( .A(n19238), .B(n19237), .Z(n19242) );
  NAND U20120 ( .A(n19240), .B(n19239), .Z(n19241) );
  NAND U20121 ( .A(n19242), .B(n19241), .Z(n19437) );
  XNOR U20122 ( .A(b[19]), .B(a[123]), .Z(n19404) );
  NANDN U20123 ( .A(n19404), .B(n37934), .Z(n19245) );
  NANDN U20124 ( .A(n19243), .B(n37935), .Z(n19244) );
  NAND U20125 ( .A(n19245), .B(n19244), .Z(n19449) );
  XOR U20126 ( .A(b[27]), .B(a[115]), .Z(n19407) );
  NAND U20127 ( .A(n38423), .B(n19407), .Z(n19248) );
  NAND U20128 ( .A(n19246), .B(n38424), .Z(n19247) );
  NAND U20129 ( .A(n19248), .B(n19247), .Z(n19446) );
  XOR U20130 ( .A(b[5]), .B(n23393), .Z(n19410) );
  NANDN U20131 ( .A(n19410), .B(n36587), .Z(n19251) );
  NANDN U20132 ( .A(n19249), .B(n36588), .Z(n19250) );
  AND U20133 ( .A(n19251), .B(n19250), .Z(n19447) );
  XNOR U20134 ( .A(n19446), .B(n19447), .Z(n19448) );
  XNOR U20135 ( .A(n19449), .B(n19448), .Z(n19434) );
  NAND U20136 ( .A(n19252), .B(n37762), .Z(n19254) );
  XOR U20137 ( .A(b[17]), .B(a[125]), .Z(n19413) );
  NAND U20138 ( .A(n19413), .B(n37764), .Z(n19253) );
  NAND U20139 ( .A(n19254), .B(n19253), .Z(n19388) );
  XNOR U20140 ( .A(b[31]), .B(a[111]), .Z(n19416) );
  NANDN U20141 ( .A(n19416), .B(n38552), .Z(n19257) );
  NANDN U20142 ( .A(n19255), .B(n38553), .Z(n19256) );
  AND U20143 ( .A(n19257), .B(n19256), .Z(n19386) );
  OR U20144 ( .A(n19258), .B(n36105), .Z(n19260) );
  XOR U20145 ( .A(b[3]), .B(n23668), .Z(n19419) );
  NANDN U20146 ( .A(n19419), .B(n36107), .Z(n19259) );
  AND U20147 ( .A(n19260), .B(n19259), .Z(n19387) );
  XOR U20148 ( .A(n19388), .B(n19389), .Z(n19435) );
  XOR U20149 ( .A(n19434), .B(n19435), .Z(n19436) );
  XNOR U20150 ( .A(n19437), .B(n19436), .Z(n19482) );
  NANDN U20151 ( .A(n19262), .B(n19261), .Z(n19266) );
  NAND U20152 ( .A(n19264), .B(n19263), .Z(n19265) );
  NAND U20153 ( .A(n19266), .B(n19265), .Z(n19425) );
  NANDN U20154 ( .A(n19268), .B(n19267), .Z(n19272) );
  NAND U20155 ( .A(n19270), .B(n19269), .Z(n19271) );
  NAND U20156 ( .A(n19272), .B(n19271), .Z(n19423) );
  OR U20157 ( .A(n19274), .B(n19273), .Z(n19278) );
  NANDN U20158 ( .A(n19276), .B(n19275), .Z(n19277) );
  NAND U20159 ( .A(n19278), .B(n19277), .Z(n19422) );
  XNOR U20160 ( .A(n19425), .B(n19424), .Z(n19483) );
  XOR U20161 ( .A(n19482), .B(n19483), .Z(n19485) );
  NANDN U20162 ( .A(n19280), .B(n19279), .Z(n19284) );
  OR U20163 ( .A(n19282), .B(n19281), .Z(n19283) );
  NAND U20164 ( .A(n19284), .B(n19283), .Z(n19484) );
  XOR U20165 ( .A(n19485), .B(n19484), .Z(n19502) );
  OR U20166 ( .A(n19286), .B(n19285), .Z(n19290) );
  NANDN U20167 ( .A(n19288), .B(n19287), .Z(n19289) );
  NAND U20168 ( .A(n19290), .B(n19289), .Z(n19501) );
  NANDN U20169 ( .A(n19292), .B(n19291), .Z(n19296) );
  NANDN U20170 ( .A(n19294), .B(n19293), .Z(n19295) );
  NAND U20171 ( .A(n19296), .B(n19295), .Z(n19490) );
  NANDN U20172 ( .A(n19298), .B(n19297), .Z(n19302) );
  OR U20173 ( .A(n19300), .B(n19299), .Z(n19301) );
  NAND U20174 ( .A(n19302), .B(n19301), .Z(n19489) );
  NANDN U20175 ( .A(n19304), .B(n19303), .Z(n19308) );
  NAND U20176 ( .A(n19306), .B(n19305), .Z(n19307) );
  NAND U20177 ( .A(n19308), .B(n19307), .Z(n19428) );
  NANDN U20178 ( .A(n19310), .B(n19309), .Z(n19314) );
  NAND U20179 ( .A(n19312), .B(n19311), .Z(n19313) );
  AND U20180 ( .A(n19314), .B(n19313), .Z(n19429) );
  XNOR U20181 ( .A(n19428), .B(n19429), .Z(n19430) );
  XNOR U20182 ( .A(n1052), .B(a[133]), .Z(n19458) );
  NAND U20183 ( .A(n36925), .B(n19458), .Z(n19317) );
  NANDN U20184 ( .A(n19315), .B(n36926), .Z(n19316) );
  NAND U20185 ( .A(n19317), .B(n19316), .Z(n19394) );
  XNOR U20186 ( .A(b[15]), .B(a[127]), .Z(n19455) );
  OR U20187 ( .A(n19455), .B(n37665), .Z(n19320) );
  NANDN U20188 ( .A(n19318), .B(n37604), .Z(n19319) );
  AND U20189 ( .A(n19320), .B(n19319), .Z(n19392) );
  XNOR U20190 ( .A(n1056), .B(a[121]), .Z(n19452) );
  NAND U20191 ( .A(n19452), .B(n38101), .Z(n19323) );
  NANDN U20192 ( .A(n19321), .B(n38102), .Z(n19322) );
  AND U20193 ( .A(n19323), .B(n19322), .Z(n19393) );
  XOR U20194 ( .A(n19394), .B(n19395), .Z(n19383) );
  XOR U20195 ( .A(b[11]), .B(n22518), .Z(n19461) );
  OR U20196 ( .A(n19461), .B(n37311), .Z(n19326) );
  NANDN U20197 ( .A(n19324), .B(n37218), .Z(n19325) );
  NAND U20198 ( .A(n19326), .B(n19325), .Z(n19381) );
  XOR U20199 ( .A(n1053), .B(a[129]), .Z(n19464) );
  NANDN U20200 ( .A(n19464), .B(n37424), .Z(n19329) );
  NANDN U20201 ( .A(n19327), .B(n37425), .Z(n19328) );
  NAND U20202 ( .A(n19329), .B(n19328), .Z(n19380) );
  XOR U20203 ( .A(n19383), .B(n19382), .Z(n19377) );
  NAND U20204 ( .A(n38490), .B(n19330), .Z(n19332) );
  XOR U20205 ( .A(n1058), .B(n19909), .Z(n19467) );
  NANDN U20206 ( .A(n1048), .B(n19467), .Z(n19331) );
  NAND U20207 ( .A(n19332), .B(n19331), .Z(n19398) );
  NANDN U20208 ( .A(n1059), .B(a[109]), .Z(n19399) );
  XNOR U20209 ( .A(n19398), .B(n19399), .Z(n19401) );
  NANDN U20210 ( .A(n1049), .B(a[141]), .Z(n19333) );
  XNOR U20211 ( .A(b[1]), .B(n19333), .Z(n19335) );
  NANDN U20212 ( .A(b[0]), .B(a[140]), .Z(n19334) );
  AND U20213 ( .A(n19335), .B(n19334), .Z(n19400) );
  XNOR U20214 ( .A(n19401), .B(n19400), .Z(n19375) );
  NANDN U20215 ( .A(n19336), .B(n38205), .Z(n19338) );
  XNOR U20216 ( .A(b[23]), .B(a[119]), .Z(n19473) );
  OR U20217 ( .A(n19473), .B(n38268), .Z(n19337) );
  NAND U20218 ( .A(n19338), .B(n19337), .Z(n19443) );
  XOR U20219 ( .A(b[7]), .B(a[135]), .Z(n19476) );
  NAND U20220 ( .A(n19476), .B(n36701), .Z(n19341) );
  NAND U20221 ( .A(n19339), .B(n36702), .Z(n19340) );
  NAND U20222 ( .A(n19341), .B(n19340), .Z(n19440) );
  XOR U20223 ( .A(b[25]), .B(a[117]), .Z(n19479) );
  NAND U20224 ( .A(n19479), .B(n38325), .Z(n19344) );
  NAND U20225 ( .A(n19342), .B(n38326), .Z(n19343) );
  AND U20226 ( .A(n19344), .B(n19343), .Z(n19441) );
  XNOR U20227 ( .A(n19440), .B(n19441), .Z(n19442) );
  XOR U20228 ( .A(n19443), .B(n19442), .Z(n19374) );
  XOR U20229 ( .A(n19377), .B(n19376), .Z(n19431) );
  XNOR U20230 ( .A(n19430), .B(n19431), .Z(n19488) );
  XNOR U20231 ( .A(n19489), .B(n19488), .Z(n19491) );
  XNOR U20232 ( .A(n19490), .B(n19491), .Z(n19500) );
  XOR U20233 ( .A(n19501), .B(n19500), .Z(n19503) );
  NAND U20234 ( .A(n19346), .B(n19345), .Z(n19350) );
  NAND U20235 ( .A(n19348), .B(n19347), .Z(n19349) );
  NAND U20236 ( .A(n19350), .B(n19349), .Z(n19495) );
  NANDN U20237 ( .A(n19352), .B(n19351), .Z(n19356) );
  NAND U20238 ( .A(n19354), .B(n19353), .Z(n19355) );
  AND U20239 ( .A(n19356), .B(n19355), .Z(n19494) );
  XNOR U20240 ( .A(n19495), .B(n19494), .Z(n19496) );
  XOR U20241 ( .A(n19497), .B(n19496), .Z(n19371) );
  XOR U20242 ( .A(n19370), .B(n19371), .Z(n19362) );
  XOR U20243 ( .A(n19363), .B(n19362), .Z(n19364) );
  XNOR U20244 ( .A(n19365), .B(n19364), .Z(n19506) );
  XNOR U20245 ( .A(n19506), .B(sreg[365]), .Z(n19508) );
  NAND U20246 ( .A(n19357), .B(sreg[364]), .Z(n19361) );
  OR U20247 ( .A(n19359), .B(n19358), .Z(n19360) );
  AND U20248 ( .A(n19361), .B(n19360), .Z(n19507) );
  XOR U20249 ( .A(n19508), .B(n19507), .Z(c[365]) );
  NAND U20250 ( .A(n19363), .B(n19362), .Z(n19367) );
  NAND U20251 ( .A(n19365), .B(n19364), .Z(n19366) );
  NAND U20252 ( .A(n19367), .B(n19366), .Z(n19514) );
  NANDN U20253 ( .A(n19369), .B(n19368), .Z(n19373) );
  NAND U20254 ( .A(n19371), .B(n19370), .Z(n19372) );
  NAND U20255 ( .A(n19373), .B(n19372), .Z(n19512) );
  NANDN U20256 ( .A(n19375), .B(n19374), .Z(n19379) );
  NANDN U20257 ( .A(n19377), .B(n19376), .Z(n19378) );
  NAND U20258 ( .A(n19379), .B(n19378), .Z(n19630) );
  OR U20259 ( .A(n19381), .B(n19380), .Z(n19385) );
  NAND U20260 ( .A(n19383), .B(n19382), .Z(n19384) );
  NAND U20261 ( .A(n19385), .B(n19384), .Z(n19569) );
  OR U20262 ( .A(n19387), .B(n19386), .Z(n19391) );
  NANDN U20263 ( .A(n19389), .B(n19388), .Z(n19390) );
  NAND U20264 ( .A(n19391), .B(n19390), .Z(n19568) );
  OR U20265 ( .A(n19393), .B(n19392), .Z(n19397) );
  NANDN U20266 ( .A(n19395), .B(n19394), .Z(n19396) );
  NAND U20267 ( .A(n19397), .B(n19396), .Z(n19567) );
  XOR U20268 ( .A(n19569), .B(n19570), .Z(n19627) );
  NANDN U20269 ( .A(n19399), .B(n19398), .Z(n19403) );
  NAND U20270 ( .A(n19401), .B(n19400), .Z(n19402) );
  NAND U20271 ( .A(n19403), .B(n19402), .Z(n19582) );
  XNOR U20272 ( .A(b[19]), .B(a[124]), .Z(n19527) );
  NANDN U20273 ( .A(n19527), .B(n37934), .Z(n19406) );
  NANDN U20274 ( .A(n19404), .B(n37935), .Z(n19405) );
  NAND U20275 ( .A(n19406), .B(n19405), .Z(n19594) );
  XOR U20276 ( .A(b[27]), .B(a[116]), .Z(n19530) );
  NAND U20277 ( .A(n38423), .B(n19530), .Z(n19409) );
  NAND U20278 ( .A(n19407), .B(n38424), .Z(n19408) );
  NAND U20279 ( .A(n19409), .B(n19408), .Z(n19591) );
  XNOR U20280 ( .A(b[5]), .B(a[138]), .Z(n19533) );
  NANDN U20281 ( .A(n19533), .B(n36587), .Z(n19412) );
  NANDN U20282 ( .A(n19410), .B(n36588), .Z(n19411) );
  AND U20283 ( .A(n19412), .B(n19411), .Z(n19592) );
  XNOR U20284 ( .A(n19591), .B(n19592), .Z(n19593) );
  XNOR U20285 ( .A(n19594), .B(n19593), .Z(n19580) );
  NAND U20286 ( .A(n19413), .B(n37762), .Z(n19415) );
  XOR U20287 ( .A(b[17]), .B(a[126]), .Z(n19536) );
  NAND U20288 ( .A(n19536), .B(n37764), .Z(n19414) );
  NAND U20289 ( .A(n19415), .B(n19414), .Z(n19554) );
  XNOR U20290 ( .A(b[31]), .B(a[112]), .Z(n19539) );
  NANDN U20291 ( .A(n19539), .B(n38552), .Z(n19418) );
  NANDN U20292 ( .A(n19416), .B(n38553), .Z(n19417) );
  NAND U20293 ( .A(n19418), .B(n19417), .Z(n19551) );
  OR U20294 ( .A(n19419), .B(n36105), .Z(n19421) );
  XNOR U20295 ( .A(b[3]), .B(a[140]), .Z(n19542) );
  NANDN U20296 ( .A(n19542), .B(n36107), .Z(n19420) );
  AND U20297 ( .A(n19421), .B(n19420), .Z(n19552) );
  XNOR U20298 ( .A(n19551), .B(n19552), .Z(n19553) );
  XOR U20299 ( .A(n19554), .B(n19553), .Z(n19579) );
  XNOR U20300 ( .A(n19580), .B(n19579), .Z(n19581) );
  XNOR U20301 ( .A(n19582), .B(n19581), .Z(n19628) );
  XNOR U20302 ( .A(n19627), .B(n19628), .Z(n19629) );
  XNOR U20303 ( .A(n19630), .B(n19629), .Z(n19648) );
  OR U20304 ( .A(n19423), .B(n19422), .Z(n19427) );
  NAND U20305 ( .A(n19425), .B(n19424), .Z(n19426) );
  NAND U20306 ( .A(n19427), .B(n19426), .Z(n19646) );
  NANDN U20307 ( .A(n19429), .B(n19428), .Z(n19433) );
  NANDN U20308 ( .A(n19431), .B(n19430), .Z(n19432) );
  NAND U20309 ( .A(n19433), .B(n19432), .Z(n19635) );
  OR U20310 ( .A(n19435), .B(n19434), .Z(n19439) );
  NAND U20311 ( .A(n19437), .B(n19436), .Z(n19438) );
  NAND U20312 ( .A(n19439), .B(n19438), .Z(n19634) );
  NANDN U20313 ( .A(n19441), .B(n19440), .Z(n19445) );
  NAND U20314 ( .A(n19443), .B(n19442), .Z(n19444) );
  NAND U20315 ( .A(n19445), .B(n19444), .Z(n19573) );
  NANDN U20316 ( .A(n19447), .B(n19446), .Z(n19451) );
  NAND U20317 ( .A(n19449), .B(n19448), .Z(n19450) );
  AND U20318 ( .A(n19451), .B(n19450), .Z(n19574) );
  XNOR U20319 ( .A(n19573), .B(n19574), .Z(n19575) );
  XOR U20320 ( .A(n1056), .B(a[122]), .Z(n19603) );
  NANDN U20321 ( .A(n19603), .B(n38101), .Z(n19454) );
  NAND U20322 ( .A(n38102), .B(n19452), .Z(n19453) );
  NAND U20323 ( .A(n19454), .B(n19453), .Z(n19563) );
  XNOR U20324 ( .A(b[15]), .B(a[128]), .Z(n19600) );
  OR U20325 ( .A(n19600), .B(n37665), .Z(n19457) );
  NANDN U20326 ( .A(n19455), .B(n37604), .Z(n19456) );
  AND U20327 ( .A(n19457), .B(n19456), .Z(n19564) );
  XNOR U20328 ( .A(n19563), .B(n19564), .Z(n19566) );
  XOR U20329 ( .A(n1052), .B(a[134]), .Z(n19597) );
  NANDN U20330 ( .A(n19597), .B(n36925), .Z(n19460) );
  NAND U20331 ( .A(n36926), .B(n19458), .Z(n19459) );
  NAND U20332 ( .A(n19460), .B(n19459), .Z(n19565) );
  XNOR U20333 ( .A(n19566), .B(n19565), .Z(n19559) );
  XNOR U20334 ( .A(b[11]), .B(a[132]), .Z(n19606) );
  OR U20335 ( .A(n19606), .B(n37311), .Z(n19463) );
  NANDN U20336 ( .A(n19461), .B(n37218), .Z(n19462) );
  NAND U20337 ( .A(n19463), .B(n19462), .Z(n19558) );
  XOR U20338 ( .A(n1053), .B(a[130]), .Z(n19609) );
  NANDN U20339 ( .A(n19609), .B(n37424), .Z(n19466) );
  NANDN U20340 ( .A(n19464), .B(n37425), .Z(n19465) );
  NAND U20341 ( .A(n19466), .B(n19465), .Z(n19557) );
  XNOR U20342 ( .A(n19558), .B(n19557), .Z(n19560) );
  XNOR U20343 ( .A(n19559), .B(n19560), .Z(n19548) );
  NAND U20344 ( .A(n38490), .B(n19467), .Z(n19469) );
  XNOR U20345 ( .A(n1058), .B(a[114]), .Z(n19615) );
  NANDN U20346 ( .A(n1048), .B(n19615), .Z(n19468) );
  NAND U20347 ( .A(n19469), .B(n19468), .Z(n19521) );
  NANDN U20348 ( .A(n1059), .B(a[110]), .Z(n19522) );
  XNOR U20349 ( .A(n19521), .B(n19522), .Z(n19524) );
  NANDN U20350 ( .A(n1049), .B(a[142]), .Z(n19470) );
  XNOR U20351 ( .A(b[1]), .B(n19470), .Z(n19472) );
  IV U20352 ( .A(a[141]), .Z(n23961) );
  NANDN U20353 ( .A(n23961), .B(n1049), .Z(n19471) );
  AND U20354 ( .A(n19472), .B(n19471), .Z(n19523) );
  XNOR U20355 ( .A(n19524), .B(n19523), .Z(n19546) );
  NANDN U20356 ( .A(n19473), .B(n38205), .Z(n19475) );
  XNOR U20357 ( .A(b[23]), .B(a[120]), .Z(n19618) );
  OR U20358 ( .A(n19618), .B(n38268), .Z(n19474) );
  NAND U20359 ( .A(n19475), .B(n19474), .Z(n19588) );
  XOR U20360 ( .A(b[7]), .B(a[136]), .Z(n19621) );
  NAND U20361 ( .A(n19621), .B(n36701), .Z(n19478) );
  NAND U20362 ( .A(n19476), .B(n36702), .Z(n19477) );
  NAND U20363 ( .A(n19478), .B(n19477), .Z(n19585) );
  XNOR U20364 ( .A(b[25]), .B(a[118]), .Z(n19624) );
  NANDN U20365 ( .A(n19624), .B(n38325), .Z(n19481) );
  NAND U20366 ( .A(n19479), .B(n38326), .Z(n19480) );
  AND U20367 ( .A(n19481), .B(n19480), .Z(n19586) );
  XNOR U20368 ( .A(n19585), .B(n19586), .Z(n19587) );
  XOR U20369 ( .A(n19588), .B(n19587), .Z(n19545) );
  XOR U20370 ( .A(n19548), .B(n19547), .Z(n19576) );
  XNOR U20371 ( .A(n19575), .B(n19576), .Z(n19633) );
  XNOR U20372 ( .A(n19634), .B(n19633), .Z(n19636) );
  XNOR U20373 ( .A(n19635), .B(n19636), .Z(n19645) );
  XNOR U20374 ( .A(n19646), .B(n19645), .Z(n19647) );
  XOR U20375 ( .A(n19648), .B(n19647), .Z(n19642) );
  NANDN U20376 ( .A(n19483), .B(n19482), .Z(n19487) );
  OR U20377 ( .A(n19485), .B(n19484), .Z(n19486) );
  NAND U20378 ( .A(n19487), .B(n19486), .Z(n19639) );
  NAND U20379 ( .A(n19489), .B(n19488), .Z(n19493) );
  NANDN U20380 ( .A(n19491), .B(n19490), .Z(n19492) );
  NAND U20381 ( .A(n19493), .B(n19492), .Z(n19640) );
  XNOR U20382 ( .A(n19639), .B(n19640), .Z(n19641) );
  XNOR U20383 ( .A(n19642), .B(n19641), .Z(n19518) );
  NANDN U20384 ( .A(n19495), .B(n19494), .Z(n19499) );
  NAND U20385 ( .A(n19497), .B(n19496), .Z(n19498) );
  NAND U20386 ( .A(n19499), .B(n19498), .Z(n19515) );
  NANDN U20387 ( .A(n19501), .B(n19500), .Z(n19505) );
  OR U20388 ( .A(n19503), .B(n19502), .Z(n19504) );
  NAND U20389 ( .A(n19505), .B(n19504), .Z(n19516) );
  XNOR U20390 ( .A(n19515), .B(n19516), .Z(n19517) );
  XNOR U20391 ( .A(n19518), .B(n19517), .Z(n19511) );
  XOR U20392 ( .A(n19512), .B(n19511), .Z(n19513) );
  XNOR U20393 ( .A(n19514), .B(n19513), .Z(n19651) );
  XNOR U20394 ( .A(n19651), .B(sreg[366]), .Z(n19653) );
  NAND U20395 ( .A(n19506), .B(sreg[365]), .Z(n19510) );
  OR U20396 ( .A(n19508), .B(n19507), .Z(n19509) );
  AND U20397 ( .A(n19510), .B(n19509), .Z(n19652) );
  XOR U20398 ( .A(n19653), .B(n19652), .Z(c[366]) );
  NANDN U20399 ( .A(n19516), .B(n19515), .Z(n19520) );
  NANDN U20400 ( .A(n19518), .B(n19517), .Z(n19519) );
  NAND U20401 ( .A(n19520), .B(n19519), .Z(n19657) );
  NANDN U20402 ( .A(n19522), .B(n19521), .Z(n19526) );
  NAND U20403 ( .A(n19524), .B(n19523), .Z(n19525) );
  NAND U20404 ( .A(n19526), .B(n19525), .Z(n19727) );
  XNOR U20405 ( .A(b[19]), .B(a[125]), .Z(n19674) );
  NANDN U20406 ( .A(n19674), .B(n37934), .Z(n19529) );
  NANDN U20407 ( .A(n19527), .B(n37935), .Z(n19528) );
  NAND U20408 ( .A(n19529), .B(n19528), .Z(n19737) );
  XOR U20409 ( .A(b[27]), .B(a[117]), .Z(n19677) );
  NAND U20410 ( .A(n38423), .B(n19677), .Z(n19532) );
  NAND U20411 ( .A(n19530), .B(n38424), .Z(n19531) );
  NAND U20412 ( .A(n19532), .B(n19531), .Z(n19734) );
  XOR U20413 ( .A(b[5]), .B(n23668), .Z(n19680) );
  NANDN U20414 ( .A(n19680), .B(n36587), .Z(n19535) );
  NANDN U20415 ( .A(n19533), .B(n36588), .Z(n19534) );
  AND U20416 ( .A(n19535), .B(n19534), .Z(n19735) );
  XNOR U20417 ( .A(n19734), .B(n19735), .Z(n19736) );
  XNOR U20418 ( .A(n19737), .B(n19736), .Z(n19725) );
  NAND U20419 ( .A(n19536), .B(n37762), .Z(n19538) );
  XOR U20420 ( .A(b[17]), .B(a[127]), .Z(n19683) );
  NAND U20421 ( .A(n19683), .B(n37764), .Z(n19537) );
  NAND U20422 ( .A(n19538), .B(n19537), .Z(n19701) );
  XOR U20423 ( .A(b[31]), .B(n19909), .Z(n19686) );
  NANDN U20424 ( .A(n19686), .B(n38552), .Z(n19541) );
  NANDN U20425 ( .A(n19539), .B(n38553), .Z(n19540) );
  NAND U20426 ( .A(n19541), .B(n19540), .Z(n19698) );
  OR U20427 ( .A(n19542), .B(n36105), .Z(n19544) );
  XOR U20428 ( .A(b[3]), .B(n23961), .Z(n19689) );
  NANDN U20429 ( .A(n19689), .B(n36107), .Z(n19543) );
  AND U20430 ( .A(n19544), .B(n19543), .Z(n19699) );
  XNOR U20431 ( .A(n19698), .B(n19699), .Z(n19700) );
  XOR U20432 ( .A(n19701), .B(n19700), .Z(n19724) );
  XNOR U20433 ( .A(n19725), .B(n19724), .Z(n19726) );
  XNOR U20434 ( .A(n19727), .B(n19726), .Z(n19776) );
  NANDN U20435 ( .A(n19546), .B(n19545), .Z(n19550) );
  NANDN U20436 ( .A(n19548), .B(n19547), .Z(n19549) );
  NAND U20437 ( .A(n19550), .B(n19549), .Z(n19777) );
  XNOR U20438 ( .A(n19776), .B(n19777), .Z(n19778) );
  NANDN U20439 ( .A(n19552), .B(n19551), .Z(n19556) );
  NAND U20440 ( .A(n19554), .B(n19553), .Z(n19555) );
  NAND U20441 ( .A(n19556), .B(n19555), .Z(n19717) );
  OR U20442 ( .A(n19558), .B(n19557), .Z(n19562) );
  NANDN U20443 ( .A(n19560), .B(n19559), .Z(n19561) );
  NAND U20444 ( .A(n19562), .B(n19561), .Z(n19715) );
  XNOR U20445 ( .A(n19715), .B(n19714), .Z(n19716) );
  XOR U20446 ( .A(n19717), .B(n19716), .Z(n19779) );
  XOR U20447 ( .A(n19778), .B(n19779), .Z(n19789) );
  OR U20448 ( .A(n19568), .B(n19567), .Z(n19572) );
  NANDN U20449 ( .A(n19570), .B(n19569), .Z(n19571) );
  NAND U20450 ( .A(n19572), .B(n19571), .Z(n19787) );
  NANDN U20451 ( .A(n19574), .B(n19573), .Z(n19578) );
  NANDN U20452 ( .A(n19576), .B(n19575), .Z(n19577) );
  NAND U20453 ( .A(n19578), .B(n19577), .Z(n19772) );
  NANDN U20454 ( .A(n19580), .B(n19579), .Z(n19584) );
  NAND U20455 ( .A(n19582), .B(n19581), .Z(n19583) );
  NAND U20456 ( .A(n19584), .B(n19583), .Z(n19771) );
  NANDN U20457 ( .A(n19586), .B(n19585), .Z(n19590) );
  NAND U20458 ( .A(n19588), .B(n19587), .Z(n19589) );
  NAND U20459 ( .A(n19590), .B(n19589), .Z(n19718) );
  NANDN U20460 ( .A(n19592), .B(n19591), .Z(n19596) );
  NAND U20461 ( .A(n19594), .B(n19593), .Z(n19595) );
  AND U20462 ( .A(n19596), .B(n19595), .Z(n19719) );
  XNOR U20463 ( .A(n19718), .B(n19719), .Z(n19720) );
  XNOR U20464 ( .A(b[9]), .B(a[135]), .Z(n19740) );
  NANDN U20465 ( .A(n19740), .B(n36925), .Z(n19599) );
  NANDN U20466 ( .A(n19597), .B(n36926), .Z(n19598) );
  NAND U20467 ( .A(n19599), .B(n19598), .Z(n19706) );
  XNOR U20468 ( .A(n1054), .B(a[129]), .Z(n19743) );
  NANDN U20469 ( .A(n37665), .B(n19743), .Z(n19602) );
  NANDN U20470 ( .A(n19600), .B(n37604), .Z(n19601) );
  NAND U20471 ( .A(n19602), .B(n19601), .Z(n19704) );
  XNOR U20472 ( .A(b[21]), .B(a[123]), .Z(n19746) );
  NANDN U20473 ( .A(n19746), .B(n38101), .Z(n19605) );
  NANDN U20474 ( .A(n19603), .B(n38102), .Z(n19604) );
  NAND U20475 ( .A(n19605), .B(n19604), .Z(n19705) );
  XNOR U20476 ( .A(n19704), .B(n19705), .Z(n19707) );
  XOR U20477 ( .A(n19706), .B(n19707), .Z(n19695) );
  XNOR U20478 ( .A(b[11]), .B(a[133]), .Z(n19749) );
  OR U20479 ( .A(n19749), .B(n37311), .Z(n19608) );
  NANDN U20480 ( .A(n19606), .B(n37218), .Z(n19607) );
  NAND U20481 ( .A(n19608), .B(n19607), .Z(n19693) );
  XOR U20482 ( .A(n1053), .B(a[131]), .Z(n19752) );
  NANDN U20483 ( .A(n19752), .B(n37424), .Z(n19611) );
  NANDN U20484 ( .A(n19609), .B(n37425), .Z(n19610) );
  AND U20485 ( .A(n19611), .B(n19610), .Z(n19692) );
  XNOR U20486 ( .A(n19693), .B(n19692), .Z(n19694) );
  XNOR U20487 ( .A(n19695), .B(n19694), .Z(n19711) );
  NANDN U20488 ( .A(n1049), .B(a[143]), .Z(n19612) );
  XNOR U20489 ( .A(b[1]), .B(n19612), .Z(n19614) );
  IV U20490 ( .A(a[142]), .Z(n24120) );
  NANDN U20491 ( .A(n24120), .B(n1049), .Z(n19613) );
  AND U20492 ( .A(n19614), .B(n19613), .Z(n19670) );
  NAND U20493 ( .A(n38490), .B(n19615), .Z(n19617) );
  XNOR U20494 ( .A(n1058), .B(a[115]), .Z(n19755) );
  NANDN U20495 ( .A(n1048), .B(n19755), .Z(n19616) );
  NAND U20496 ( .A(n19617), .B(n19616), .Z(n19668) );
  NANDN U20497 ( .A(n1059), .B(a[111]), .Z(n19669) );
  XNOR U20498 ( .A(n19668), .B(n19669), .Z(n19671) );
  XNOR U20499 ( .A(n19670), .B(n19671), .Z(n19709) );
  NANDN U20500 ( .A(n19618), .B(n38205), .Z(n19620) );
  XNOR U20501 ( .A(b[23]), .B(a[121]), .Z(n19761) );
  OR U20502 ( .A(n19761), .B(n38268), .Z(n19619) );
  NAND U20503 ( .A(n19620), .B(n19619), .Z(n19731) );
  XNOR U20504 ( .A(b[7]), .B(a[137]), .Z(n19764) );
  NANDN U20505 ( .A(n19764), .B(n36701), .Z(n19623) );
  NAND U20506 ( .A(n19621), .B(n36702), .Z(n19622) );
  NAND U20507 ( .A(n19623), .B(n19622), .Z(n19728) );
  XOR U20508 ( .A(b[25]), .B(a[119]), .Z(n19767) );
  NAND U20509 ( .A(n19767), .B(n38325), .Z(n19626) );
  NANDN U20510 ( .A(n19624), .B(n38326), .Z(n19625) );
  AND U20511 ( .A(n19626), .B(n19625), .Z(n19729) );
  XNOR U20512 ( .A(n19728), .B(n19729), .Z(n19730) );
  XOR U20513 ( .A(n19731), .B(n19730), .Z(n19708) );
  XOR U20514 ( .A(n19711), .B(n19710), .Z(n19721) );
  XOR U20515 ( .A(n19720), .B(n19721), .Z(n19770) );
  XNOR U20516 ( .A(n19771), .B(n19770), .Z(n19773) );
  XNOR U20517 ( .A(n19772), .B(n19773), .Z(n19786) );
  XOR U20518 ( .A(n19787), .B(n19786), .Z(n19788) );
  XNOR U20519 ( .A(n19789), .B(n19788), .Z(n19783) );
  NANDN U20520 ( .A(n19628), .B(n19627), .Z(n19632) );
  NAND U20521 ( .A(n19630), .B(n19629), .Z(n19631) );
  NAND U20522 ( .A(n19632), .B(n19631), .Z(n19781) );
  NAND U20523 ( .A(n19634), .B(n19633), .Z(n19638) );
  NANDN U20524 ( .A(n19636), .B(n19635), .Z(n19637) );
  AND U20525 ( .A(n19638), .B(n19637), .Z(n19780) );
  XNOR U20526 ( .A(n19781), .B(n19780), .Z(n19782) );
  XOR U20527 ( .A(n19783), .B(n19782), .Z(n19664) );
  NANDN U20528 ( .A(n19640), .B(n19639), .Z(n19644) );
  NAND U20529 ( .A(n19642), .B(n19641), .Z(n19643) );
  NAND U20530 ( .A(n19644), .B(n19643), .Z(n19662) );
  NANDN U20531 ( .A(n19646), .B(n19645), .Z(n19650) );
  NANDN U20532 ( .A(n19648), .B(n19647), .Z(n19649) );
  NAND U20533 ( .A(n19650), .B(n19649), .Z(n19663) );
  XNOR U20534 ( .A(n19662), .B(n19663), .Z(n19665) );
  XOR U20535 ( .A(n19664), .B(n19665), .Z(n19656) );
  XOR U20536 ( .A(n19657), .B(n19656), .Z(n19658) );
  XNOR U20537 ( .A(n19659), .B(n19658), .Z(n19792) );
  XNOR U20538 ( .A(n19792), .B(sreg[367]), .Z(n19794) );
  NAND U20539 ( .A(n19651), .B(sreg[366]), .Z(n19655) );
  OR U20540 ( .A(n19653), .B(n19652), .Z(n19654) );
  AND U20541 ( .A(n19655), .B(n19654), .Z(n19793) );
  XOR U20542 ( .A(n19794), .B(n19793), .Z(c[367]) );
  NAND U20543 ( .A(n19657), .B(n19656), .Z(n19661) );
  NAND U20544 ( .A(n19659), .B(n19658), .Z(n19660) );
  NAND U20545 ( .A(n19661), .B(n19660), .Z(n19800) );
  NANDN U20546 ( .A(n19663), .B(n19662), .Z(n19667) );
  NAND U20547 ( .A(n19665), .B(n19664), .Z(n19666) );
  NAND U20548 ( .A(n19667), .B(n19666), .Z(n19798) );
  NANDN U20549 ( .A(n19669), .B(n19668), .Z(n19673) );
  NAND U20550 ( .A(n19671), .B(n19670), .Z(n19672) );
  NAND U20551 ( .A(n19673), .B(n19672), .Z(n19878) );
  XNOR U20552 ( .A(b[19]), .B(a[126]), .Z(n19823) );
  NANDN U20553 ( .A(n19823), .B(n37934), .Z(n19676) );
  NANDN U20554 ( .A(n19674), .B(n37935), .Z(n19675) );
  NAND U20555 ( .A(n19676), .B(n19675), .Z(n19888) );
  XNOR U20556 ( .A(b[27]), .B(a[118]), .Z(n19826) );
  NANDN U20557 ( .A(n19826), .B(n38423), .Z(n19679) );
  NAND U20558 ( .A(n19677), .B(n38424), .Z(n19678) );
  NAND U20559 ( .A(n19679), .B(n19678), .Z(n19885) );
  XNOR U20560 ( .A(b[5]), .B(a[140]), .Z(n19829) );
  NANDN U20561 ( .A(n19829), .B(n36587), .Z(n19682) );
  NANDN U20562 ( .A(n19680), .B(n36588), .Z(n19681) );
  AND U20563 ( .A(n19682), .B(n19681), .Z(n19886) );
  XNOR U20564 ( .A(n19885), .B(n19886), .Z(n19887) );
  XNOR U20565 ( .A(n19888), .B(n19887), .Z(n19876) );
  NAND U20566 ( .A(n19683), .B(n37762), .Z(n19685) );
  XOR U20567 ( .A(b[17]), .B(a[128]), .Z(n19832) );
  NAND U20568 ( .A(n19832), .B(n37764), .Z(n19684) );
  NAND U20569 ( .A(n19685), .B(n19684), .Z(n19850) );
  XNOR U20570 ( .A(b[31]), .B(a[114]), .Z(n19835) );
  NANDN U20571 ( .A(n19835), .B(n38552), .Z(n19688) );
  NANDN U20572 ( .A(n19686), .B(n38553), .Z(n19687) );
  NAND U20573 ( .A(n19688), .B(n19687), .Z(n19847) );
  OR U20574 ( .A(n19689), .B(n36105), .Z(n19691) );
  XOR U20575 ( .A(b[3]), .B(n24120), .Z(n19838) );
  NANDN U20576 ( .A(n19838), .B(n36107), .Z(n19690) );
  AND U20577 ( .A(n19691), .B(n19690), .Z(n19848) );
  XNOR U20578 ( .A(n19847), .B(n19848), .Z(n19849) );
  XOR U20579 ( .A(n19850), .B(n19849), .Z(n19875) );
  XNOR U20580 ( .A(n19876), .B(n19875), .Z(n19877) );
  XNOR U20581 ( .A(n19878), .B(n19877), .Z(n19814) );
  NANDN U20582 ( .A(n19693), .B(n19692), .Z(n19697) );
  NAND U20583 ( .A(n19695), .B(n19694), .Z(n19696) );
  NAND U20584 ( .A(n19697), .B(n19696), .Z(n19867) );
  NANDN U20585 ( .A(n19699), .B(n19698), .Z(n19703) );
  NAND U20586 ( .A(n19701), .B(n19700), .Z(n19702) );
  NAND U20587 ( .A(n19703), .B(n19702), .Z(n19866) );
  XNOR U20588 ( .A(n19866), .B(n19865), .Z(n19868) );
  XOR U20589 ( .A(n19867), .B(n19868), .Z(n19813) );
  XOR U20590 ( .A(n19814), .B(n19813), .Z(n19815) );
  NANDN U20591 ( .A(n19709), .B(n19708), .Z(n19713) );
  NAND U20592 ( .A(n19711), .B(n19710), .Z(n19712) );
  AND U20593 ( .A(n19713), .B(n19712), .Z(n19816) );
  XNOR U20594 ( .A(n19815), .B(n19816), .Z(n19925) );
  NANDN U20595 ( .A(n19719), .B(n19718), .Z(n19723) );
  NAND U20596 ( .A(n19721), .B(n19720), .Z(n19722) );
  NAND U20597 ( .A(n19723), .B(n19722), .Z(n19810) );
  NANDN U20598 ( .A(n19729), .B(n19728), .Z(n19733) );
  NAND U20599 ( .A(n19731), .B(n19730), .Z(n19732) );
  NAND U20600 ( .A(n19733), .B(n19732), .Z(n19869) );
  NANDN U20601 ( .A(n19735), .B(n19734), .Z(n19739) );
  NAND U20602 ( .A(n19737), .B(n19736), .Z(n19738) );
  AND U20603 ( .A(n19739), .B(n19738), .Z(n19870) );
  XNOR U20604 ( .A(n19869), .B(n19870), .Z(n19871) );
  XNOR U20605 ( .A(b[9]), .B(a[136]), .Z(n19891) );
  NANDN U20606 ( .A(n19891), .B(n36925), .Z(n19742) );
  NANDN U20607 ( .A(n19740), .B(n36926), .Z(n19741) );
  NAND U20608 ( .A(n19742), .B(n19741), .Z(n19861) );
  XNOR U20609 ( .A(b[15]), .B(a[130]), .Z(n19894) );
  OR U20610 ( .A(n19894), .B(n37665), .Z(n19745) );
  NAND U20611 ( .A(n19743), .B(n37604), .Z(n19744) );
  AND U20612 ( .A(n19745), .B(n19744), .Z(n19859) );
  XNOR U20613 ( .A(b[21]), .B(a[124]), .Z(n19897) );
  NANDN U20614 ( .A(n19897), .B(n38101), .Z(n19748) );
  NANDN U20615 ( .A(n19746), .B(n38102), .Z(n19747) );
  AND U20616 ( .A(n19748), .B(n19747), .Z(n19860) );
  XOR U20617 ( .A(n19861), .B(n19862), .Z(n19856) );
  XNOR U20618 ( .A(b[11]), .B(a[134]), .Z(n19900) );
  OR U20619 ( .A(n19900), .B(n37311), .Z(n19751) );
  NANDN U20620 ( .A(n19749), .B(n37218), .Z(n19750) );
  NAND U20621 ( .A(n19751), .B(n19750), .Z(n19854) );
  XOR U20622 ( .A(n1053), .B(a[132]), .Z(n19903) );
  NANDN U20623 ( .A(n19903), .B(n37424), .Z(n19754) );
  NANDN U20624 ( .A(n19752), .B(n37425), .Z(n19753) );
  NAND U20625 ( .A(n19754), .B(n19753), .Z(n19853) );
  XOR U20626 ( .A(n19856), .B(n19855), .Z(n19843) );
  NAND U20627 ( .A(n38490), .B(n19755), .Z(n19757) );
  XNOR U20628 ( .A(b[29]), .B(a[116]), .Z(n19910) );
  OR U20629 ( .A(n19910), .B(n1048), .Z(n19756) );
  NAND U20630 ( .A(n19757), .B(n19756), .Z(n19817) );
  NANDN U20631 ( .A(n1059), .B(a[112]), .Z(n19818) );
  XNOR U20632 ( .A(n19817), .B(n19818), .Z(n19820) );
  NANDN U20633 ( .A(n1049), .B(a[144]), .Z(n19758) );
  XNOR U20634 ( .A(b[1]), .B(n19758), .Z(n19760) );
  NANDN U20635 ( .A(b[0]), .B(a[143]), .Z(n19759) );
  AND U20636 ( .A(n19760), .B(n19759), .Z(n19819) );
  XOR U20637 ( .A(n19820), .B(n19819), .Z(n19841) );
  NANDN U20638 ( .A(n19761), .B(n38205), .Z(n19763) );
  XNOR U20639 ( .A(b[23]), .B(a[122]), .Z(n19913) );
  OR U20640 ( .A(n19913), .B(n38268), .Z(n19762) );
  NAND U20641 ( .A(n19763), .B(n19762), .Z(n19882) );
  XOR U20642 ( .A(b[7]), .B(a[138]), .Z(n19916) );
  NAND U20643 ( .A(n19916), .B(n36701), .Z(n19766) );
  NANDN U20644 ( .A(n19764), .B(n36702), .Z(n19765) );
  NAND U20645 ( .A(n19766), .B(n19765), .Z(n19879) );
  XOR U20646 ( .A(b[25]), .B(a[120]), .Z(n19919) );
  NAND U20647 ( .A(n19919), .B(n38325), .Z(n19769) );
  NAND U20648 ( .A(n19767), .B(n38326), .Z(n19768) );
  AND U20649 ( .A(n19769), .B(n19768), .Z(n19880) );
  XNOR U20650 ( .A(n19879), .B(n19880), .Z(n19881) );
  XNOR U20651 ( .A(n19882), .B(n19881), .Z(n19842) );
  XOR U20652 ( .A(n19841), .B(n19842), .Z(n19844) );
  XNOR U20653 ( .A(n19843), .B(n19844), .Z(n19872) );
  XOR U20654 ( .A(n19871), .B(n19872), .Z(n19808) );
  XNOR U20655 ( .A(n19807), .B(n19808), .Z(n19809) );
  XOR U20656 ( .A(n19810), .B(n19809), .Z(n19923) );
  XNOR U20657 ( .A(n19922), .B(n19923), .Z(n19924) );
  XNOR U20658 ( .A(n19925), .B(n19924), .Z(n19929) );
  NAND U20659 ( .A(n19771), .B(n19770), .Z(n19775) );
  NANDN U20660 ( .A(n19773), .B(n19772), .Z(n19774) );
  NAND U20661 ( .A(n19775), .B(n19774), .Z(n19926) );
  XNOR U20662 ( .A(n19926), .B(n19927), .Z(n19928) );
  XNOR U20663 ( .A(n19929), .B(n19928), .Z(n19804) );
  NANDN U20664 ( .A(n19781), .B(n19780), .Z(n19785) );
  NAND U20665 ( .A(n19783), .B(n19782), .Z(n19784) );
  NAND U20666 ( .A(n19785), .B(n19784), .Z(n19801) );
  NANDN U20667 ( .A(n19787), .B(n19786), .Z(n19791) );
  OR U20668 ( .A(n19789), .B(n19788), .Z(n19790) );
  NAND U20669 ( .A(n19791), .B(n19790), .Z(n19802) );
  XNOR U20670 ( .A(n19801), .B(n19802), .Z(n19803) );
  XNOR U20671 ( .A(n19804), .B(n19803), .Z(n19797) );
  XOR U20672 ( .A(n19798), .B(n19797), .Z(n19799) );
  XNOR U20673 ( .A(n19800), .B(n19799), .Z(n19932) );
  XNOR U20674 ( .A(n19932), .B(sreg[368]), .Z(n19934) );
  NAND U20675 ( .A(n19792), .B(sreg[367]), .Z(n19796) );
  OR U20676 ( .A(n19794), .B(n19793), .Z(n19795) );
  AND U20677 ( .A(n19796), .B(n19795), .Z(n19933) );
  XOR U20678 ( .A(n19934), .B(n19933), .Z(c[368]) );
  NANDN U20679 ( .A(n19802), .B(n19801), .Z(n19806) );
  NANDN U20680 ( .A(n19804), .B(n19803), .Z(n19805) );
  NAND U20681 ( .A(n19806), .B(n19805), .Z(n19937) );
  NANDN U20682 ( .A(n19808), .B(n19807), .Z(n19812) );
  NAND U20683 ( .A(n19810), .B(n19809), .Z(n19811) );
  NAND U20684 ( .A(n19812), .B(n19811), .Z(n20069) );
  XNOR U20685 ( .A(n20069), .B(n20070), .Z(n20071) );
  NANDN U20686 ( .A(n19818), .B(n19817), .Z(n19822) );
  NAND U20687 ( .A(n19820), .B(n19819), .Z(n19821) );
  NAND U20688 ( .A(n19822), .B(n19821), .Z(n20006) );
  XNOR U20689 ( .A(b[19]), .B(a[127]), .Z(n19979) );
  NANDN U20690 ( .A(n19979), .B(n37934), .Z(n19825) );
  NANDN U20691 ( .A(n19823), .B(n37935), .Z(n19824) );
  NAND U20692 ( .A(n19825), .B(n19824), .Z(n20018) );
  XOR U20693 ( .A(b[27]), .B(a[119]), .Z(n19982) );
  NAND U20694 ( .A(n38423), .B(n19982), .Z(n19828) );
  NANDN U20695 ( .A(n19826), .B(n38424), .Z(n19827) );
  NAND U20696 ( .A(n19828), .B(n19827), .Z(n20015) );
  XOR U20697 ( .A(b[5]), .B(n23961), .Z(n19985) );
  NANDN U20698 ( .A(n19985), .B(n36587), .Z(n19831) );
  NANDN U20699 ( .A(n19829), .B(n36588), .Z(n19830) );
  AND U20700 ( .A(n19831), .B(n19830), .Z(n20016) );
  XNOR U20701 ( .A(n20015), .B(n20016), .Z(n20017) );
  XNOR U20702 ( .A(n20018), .B(n20017), .Z(n20003) );
  NAND U20703 ( .A(n19832), .B(n37762), .Z(n19834) );
  XNOR U20704 ( .A(b[17]), .B(a[129]), .Z(n19988) );
  NANDN U20705 ( .A(n19988), .B(n37764), .Z(n19833) );
  NAND U20706 ( .A(n19834), .B(n19833), .Z(n19963) );
  XNOR U20707 ( .A(b[31]), .B(a[115]), .Z(n19991) );
  NANDN U20708 ( .A(n19991), .B(n38552), .Z(n19837) );
  NANDN U20709 ( .A(n19835), .B(n38553), .Z(n19836) );
  AND U20710 ( .A(n19837), .B(n19836), .Z(n19961) );
  OR U20711 ( .A(n19838), .B(n36105), .Z(n19840) );
  XNOR U20712 ( .A(b[3]), .B(a[143]), .Z(n19994) );
  NANDN U20713 ( .A(n19994), .B(n36107), .Z(n19839) );
  AND U20714 ( .A(n19840), .B(n19839), .Z(n19962) );
  XOR U20715 ( .A(n19963), .B(n19964), .Z(n20004) );
  XOR U20716 ( .A(n20003), .B(n20004), .Z(n20005) );
  XNOR U20717 ( .A(n20006), .B(n20005), .Z(n20057) );
  NANDN U20718 ( .A(n19842), .B(n19841), .Z(n19846) );
  OR U20719 ( .A(n19844), .B(n19843), .Z(n19845) );
  NAND U20720 ( .A(n19846), .B(n19845), .Z(n20058) );
  XNOR U20721 ( .A(n20057), .B(n20058), .Z(n20059) );
  NANDN U20722 ( .A(n19848), .B(n19847), .Z(n19852) );
  NAND U20723 ( .A(n19850), .B(n19849), .Z(n19851) );
  NAND U20724 ( .A(n19852), .B(n19851), .Z(n20054) );
  OR U20725 ( .A(n19854), .B(n19853), .Z(n19858) );
  NAND U20726 ( .A(n19856), .B(n19855), .Z(n19857) );
  AND U20727 ( .A(n19858), .B(n19857), .Z(n20051) );
  OR U20728 ( .A(n19860), .B(n19859), .Z(n19864) );
  NANDN U20729 ( .A(n19862), .B(n19861), .Z(n19863) );
  NAND U20730 ( .A(n19864), .B(n19863), .Z(n20052) );
  XOR U20731 ( .A(n20054), .B(n20053), .Z(n20060) );
  XNOR U20732 ( .A(n20059), .B(n20060), .Z(n20077) );
  NANDN U20733 ( .A(n19870), .B(n19869), .Z(n19874) );
  NANDN U20734 ( .A(n19872), .B(n19871), .Z(n19873) );
  NAND U20735 ( .A(n19874), .B(n19873), .Z(n20066) );
  NANDN U20736 ( .A(n19880), .B(n19879), .Z(n19884) );
  NAND U20737 ( .A(n19882), .B(n19881), .Z(n19883) );
  NAND U20738 ( .A(n19884), .B(n19883), .Z(n19997) );
  NANDN U20739 ( .A(n19886), .B(n19885), .Z(n19890) );
  NAND U20740 ( .A(n19888), .B(n19887), .Z(n19889) );
  AND U20741 ( .A(n19890), .B(n19889), .Z(n19998) );
  XNOR U20742 ( .A(n19997), .B(n19998), .Z(n19999) );
  XOR U20743 ( .A(n1052), .B(n23393), .Z(n20021) );
  NAND U20744 ( .A(n36925), .B(n20021), .Z(n19893) );
  NANDN U20745 ( .A(n19891), .B(n36926), .Z(n19892) );
  NAND U20746 ( .A(n19893), .B(n19892), .Z(n19969) );
  XOR U20747 ( .A(b[15]), .B(n22518), .Z(n20024) );
  OR U20748 ( .A(n20024), .B(n37665), .Z(n19896) );
  NANDN U20749 ( .A(n19894), .B(n37604), .Z(n19895) );
  AND U20750 ( .A(n19896), .B(n19895), .Z(n19967) );
  XNOR U20751 ( .A(n1056), .B(a[125]), .Z(n20027) );
  NAND U20752 ( .A(n20027), .B(n38101), .Z(n19899) );
  NANDN U20753 ( .A(n19897), .B(n38102), .Z(n19898) );
  AND U20754 ( .A(n19899), .B(n19898), .Z(n19968) );
  XOR U20755 ( .A(n19969), .B(n19970), .Z(n19958) );
  XNOR U20756 ( .A(b[11]), .B(a[135]), .Z(n20030) );
  OR U20757 ( .A(n20030), .B(n37311), .Z(n19902) );
  NANDN U20758 ( .A(n19900), .B(n37218), .Z(n19901) );
  NAND U20759 ( .A(n19902), .B(n19901), .Z(n19956) );
  XOR U20760 ( .A(n1053), .B(a[133]), .Z(n20033) );
  NANDN U20761 ( .A(n20033), .B(n37424), .Z(n19905) );
  NANDN U20762 ( .A(n19903), .B(n37425), .Z(n19904) );
  NAND U20763 ( .A(n19905), .B(n19904), .Z(n19955) );
  XOR U20764 ( .A(n19958), .B(n19957), .Z(n19952) );
  NANDN U20765 ( .A(n1049), .B(a[145]), .Z(n19906) );
  XNOR U20766 ( .A(b[1]), .B(n19906), .Z(n19908) );
  NANDN U20767 ( .A(b[0]), .B(a[144]), .Z(n19907) );
  AND U20768 ( .A(n19908), .B(n19907), .Z(n19976) );
  ANDN U20769 ( .B(b[31]), .A(n19909), .Z(n19973) );
  NANDN U20770 ( .A(n19910), .B(n38490), .Z(n19912) );
  XNOR U20771 ( .A(n1058), .B(a[117]), .Z(n20039) );
  NANDN U20772 ( .A(n1048), .B(n20039), .Z(n19911) );
  NAND U20773 ( .A(n19912), .B(n19911), .Z(n19974) );
  XOR U20774 ( .A(n19973), .B(n19974), .Z(n19975) );
  XNOR U20775 ( .A(n19976), .B(n19975), .Z(n19949) );
  NANDN U20776 ( .A(n19913), .B(n38205), .Z(n19915) );
  XNOR U20777 ( .A(b[23]), .B(a[123]), .Z(n20042) );
  OR U20778 ( .A(n20042), .B(n38268), .Z(n19914) );
  NAND U20779 ( .A(n19915), .B(n19914), .Z(n20012) );
  XNOR U20780 ( .A(b[7]), .B(a[139]), .Z(n20045) );
  NANDN U20781 ( .A(n20045), .B(n36701), .Z(n19918) );
  NAND U20782 ( .A(n19916), .B(n36702), .Z(n19917) );
  NAND U20783 ( .A(n19918), .B(n19917), .Z(n20009) );
  XOR U20784 ( .A(b[25]), .B(a[121]), .Z(n20048) );
  NAND U20785 ( .A(n20048), .B(n38325), .Z(n19921) );
  NAND U20786 ( .A(n19919), .B(n38326), .Z(n19920) );
  AND U20787 ( .A(n19921), .B(n19920), .Z(n20010) );
  XNOR U20788 ( .A(n20009), .B(n20010), .Z(n20011) );
  XNOR U20789 ( .A(n20012), .B(n20011), .Z(n19950) );
  XOR U20790 ( .A(n19952), .B(n19951), .Z(n20000) );
  XNOR U20791 ( .A(n19999), .B(n20000), .Z(n20063) );
  XOR U20792 ( .A(n20064), .B(n20063), .Z(n20065) );
  XNOR U20793 ( .A(n20066), .B(n20065), .Z(n20075) );
  XNOR U20794 ( .A(n20076), .B(n20075), .Z(n20078) );
  XNOR U20795 ( .A(n20077), .B(n20078), .Z(n20072) );
  XOR U20796 ( .A(n20071), .B(n20072), .Z(n19946) );
  NANDN U20797 ( .A(n19927), .B(n19926), .Z(n19931) );
  NANDN U20798 ( .A(n19929), .B(n19928), .Z(n19930) );
  NAND U20799 ( .A(n19931), .B(n19930), .Z(n19944) );
  XNOR U20800 ( .A(n19943), .B(n19944), .Z(n19945) );
  XNOR U20801 ( .A(n19946), .B(n19945), .Z(n19938) );
  XNOR U20802 ( .A(n19937), .B(n19938), .Z(n19939) );
  XNOR U20803 ( .A(n19940), .B(n19939), .Z(n20081) );
  XNOR U20804 ( .A(n20081), .B(sreg[369]), .Z(n20083) );
  NAND U20805 ( .A(n19932), .B(sreg[368]), .Z(n19936) );
  OR U20806 ( .A(n19934), .B(n19933), .Z(n19935) );
  AND U20807 ( .A(n19936), .B(n19935), .Z(n20082) );
  XOR U20808 ( .A(n20083), .B(n20082), .Z(c[369]) );
  NANDN U20809 ( .A(n19938), .B(n19937), .Z(n19942) );
  NAND U20810 ( .A(n19940), .B(n19939), .Z(n19941) );
  NAND U20811 ( .A(n19942), .B(n19941), .Z(n20089) );
  NANDN U20812 ( .A(n19944), .B(n19943), .Z(n19948) );
  NAND U20813 ( .A(n19946), .B(n19945), .Z(n19947) );
  NAND U20814 ( .A(n19948), .B(n19947), .Z(n20087) );
  OR U20815 ( .A(n19950), .B(n19949), .Z(n19954) );
  NANDN U20816 ( .A(n19952), .B(n19951), .Z(n19953) );
  NAND U20817 ( .A(n19954), .B(n19953), .Z(n20217) );
  OR U20818 ( .A(n19956), .B(n19955), .Z(n19960) );
  NAND U20819 ( .A(n19958), .B(n19957), .Z(n19959) );
  NAND U20820 ( .A(n19960), .B(n19959), .Z(n20156) );
  OR U20821 ( .A(n19962), .B(n19961), .Z(n19966) );
  NANDN U20822 ( .A(n19964), .B(n19963), .Z(n19965) );
  NAND U20823 ( .A(n19966), .B(n19965), .Z(n20155) );
  OR U20824 ( .A(n19968), .B(n19967), .Z(n19972) );
  NANDN U20825 ( .A(n19970), .B(n19969), .Z(n19971) );
  NAND U20826 ( .A(n19972), .B(n19971), .Z(n20154) );
  XOR U20827 ( .A(n20156), .B(n20157), .Z(n20215) );
  OR U20828 ( .A(n19974), .B(n19973), .Z(n19978) );
  NANDN U20829 ( .A(n19976), .B(n19975), .Z(n19977) );
  NAND U20830 ( .A(n19978), .B(n19977), .Z(n20168) );
  XNOR U20831 ( .A(b[19]), .B(a[128]), .Z(n20114) );
  NANDN U20832 ( .A(n20114), .B(n37934), .Z(n19981) );
  NANDN U20833 ( .A(n19979), .B(n37935), .Z(n19980) );
  NAND U20834 ( .A(n19981), .B(n19980), .Z(n20181) );
  XOR U20835 ( .A(b[27]), .B(a[120]), .Z(n20117) );
  NAND U20836 ( .A(n38423), .B(n20117), .Z(n19984) );
  NAND U20837 ( .A(n19982), .B(n38424), .Z(n19983) );
  NAND U20838 ( .A(n19984), .B(n19983), .Z(n20178) );
  XOR U20839 ( .A(b[5]), .B(n24120), .Z(n20120) );
  NANDN U20840 ( .A(n20120), .B(n36587), .Z(n19987) );
  NANDN U20841 ( .A(n19985), .B(n36588), .Z(n19986) );
  AND U20842 ( .A(n19987), .B(n19986), .Z(n20179) );
  XNOR U20843 ( .A(n20178), .B(n20179), .Z(n20180) );
  XNOR U20844 ( .A(n20181), .B(n20180), .Z(n20167) );
  NANDN U20845 ( .A(n19988), .B(n37762), .Z(n19990) );
  XOR U20846 ( .A(b[17]), .B(a[130]), .Z(n20123) );
  NAND U20847 ( .A(n20123), .B(n37764), .Z(n19989) );
  NAND U20848 ( .A(n19990), .B(n19989), .Z(n20141) );
  XNOR U20849 ( .A(b[31]), .B(a[116]), .Z(n20126) );
  NANDN U20850 ( .A(n20126), .B(n38552), .Z(n19993) );
  NANDN U20851 ( .A(n19991), .B(n38553), .Z(n19992) );
  NAND U20852 ( .A(n19993), .B(n19992), .Z(n20138) );
  OR U20853 ( .A(n19994), .B(n36105), .Z(n19996) );
  XNOR U20854 ( .A(b[3]), .B(a[144]), .Z(n20129) );
  NANDN U20855 ( .A(n20129), .B(n36107), .Z(n19995) );
  AND U20856 ( .A(n19996), .B(n19995), .Z(n20139) );
  XNOR U20857 ( .A(n20138), .B(n20139), .Z(n20140) );
  XOR U20858 ( .A(n20141), .B(n20140), .Z(n20166) );
  XOR U20859 ( .A(n20167), .B(n20166), .Z(n20169) );
  XOR U20860 ( .A(n20168), .B(n20169), .Z(n20214) );
  XOR U20861 ( .A(n20215), .B(n20214), .Z(n20216) );
  XNOR U20862 ( .A(n20217), .B(n20216), .Z(n20105) );
  NANDN U20863 ( .A(n19998), .B(n19997), .Z(n20002) );
  NANDN U20864 ( .A(n20000), .B(n19999), .Z(n20001) );
  NAND U20865 ( .A(n20002), .B(n20001), .Z(n20222) );
  OR U20866 ( .A(n20004), .B(n20003), .Z(n20008) );
  NAND U20867 ( .A(n20006), .B(n20005), .Z(n20007) );
  NAND U20868 ( .A(n20008), .B(n20007), .Z(n20221) );
  NANDN U20869 ( .A(n20010), .B(n20009), .Z(n20014) );
  NAND U20870 ( .A(n20012), .B(n20011), .Z(n20013) );
  NAND U20871 ( .A(n20014), .B(n20013), .Z(n20160) );
  NANDN U20872 ( .A(n20016), .B(n20015), .Z(n20020) );
  NAND U20873 ( .A(n20018), .B(n20017), .Z(n20019) );
  AND U20874 ( .A(n20020), .B(n20019), .Z(n20161) );
  XNOR U20875 ( .A(n20160), .B(n20161), .Z(n20162) );
  XNOR U20876 ( .A(b[9]), .B(a[138]), .Z(n20184) );
  NANDN U20877 ( .A(n20184), .B(n36925), .Z(n20023) );
  NAND U20878 ( .A(n36926), .B(n20021), .Z(n20022) );
  NAND U20879 ( .A(n20023), .B(n20022), .Z(n20146) );
  XNOR U20880 ( .A(n1054), .B(a[132]), .Z(n20187) );
  NANDN U20881 ( .A(n37665), .B(n20187), .Z(n20026) );
  NANDN U20882 ( .A(n20024), .B(n37604), .Z(n20025) );
  NAND U20883 ( .A(n20026), .B(n20025), .Z(n20144) );
  XNOR U20884 ( .A(b[21]), .B(a[126]), .Z(n20190) );
  NANDN U20885 ( .A(n20190), .B(n38101), .Z(n20029) );
  NAND U20886 ( .A(n38102), .B(n20027), .Z(n20028) );
  NAND U20887 ( .A(n20029), .B(n20028), .Z(n20145) );
  XNOR U20888 ( .A(n20144), .B(n20145), .Z(n20147) );
  XOR U20889 ( .A(n20146), .B(n20147), .Z(n20135) );
  XNOR U20890 ( .A(b[11]), .B(a[136]), .Z(n20193) );
  OR U20891 ( .A(n20193), .B(n37311), .Z(n20032) );
  NANDN U20892 ( .A(n20030), .B(n37218), .Z(n20031) );
  NAND U20893 ( .A(n20032), .B(n20031), .Z(n20133) );
  XOR U20894 ( .A(n1053), .B(a[134]), .Z(n20196) );
  NANDN U20895 ( .A(n20196), .B(n37424), .Z(n20035) );
  NANDN U20896 ( .A(n20033), .B(n37425), .Z(n20034) );
  AND U20897 ( .A(n20035), .B(n20034), .Z(n20132) );
  XNOR U20898 ( .A(n20133), .B(n20132), .Z(n20134) );
  XNOR U20899 ( .A(n20135), .B(n20134), .Z(n20151) );
  NANDN U20900 ( .A(n1049), .B(a[146]), .Z(n20036) );
  XNOR U20901 ( .A(b[1]), .B(n20036), .Z(n20038) );
  IV U20902 ( .A(a[145]), .Z(n24554) );
  NANDN U20903 ( .A(n24554), .B(n1049), .Z(n20037) );
  AND U20904 ( .A(n20038), .B(n20037), .Z(n20110) );
  NAND U20905 ( .A(n20039), .B(n38490), .Z(n20041) );
  XOR U20906 ( .A(n1058), .B(n20271), .Z(n20199) );
  NANDN U20907 ( .A(n1048), .B(n20199), .Z(n20040) );
  NAND U20908 ( .A(n20041), .B(n20040), .Z(n20108) );
  NANDN U20909 ( .A(n1059), .B(a[114]), .Z(n20109) );
  XNOR U20910 ( .A(n20108), .B(n20109), .Z(n20111) );
  XNOR U20911 ( .A(n20110), .B(n20111), .Z(n20149) );
  NANDN U20912 ( .A(n20042), .B(n38205), .Z(n20044) );
  XNOR U20913 ( .A(b[23]), .B(a[124]), .Z(n20205) );
  OR U20914 ( .A(n20205), .B(n38268), .Z(n20043) );
  NAND U20915 ( .A(n20044), .B(n20043), .Z(n20175) );
  XOR U20916 ( .A(b[7]), .B(a[140]), .Z(n20208) );
  NAND U20917 ( .A(n20208), .B(n36701), .Z(n20047) );
  NANDN U20918 ( .A(n20045), .B(n36702), .Z(n20046) );
  NAND U20919 ( .A(n20047), .B(n20046), .Z(n20172) );
  XOR U20920 ( .A(b[25]), .B(a[122]), .Z(n20211) );
  NAND U20921 ( .A(n20211), .B(n38325), .Z(n20050) );
  NAND U20922 ( .A(n20048), .B(n38326), .Z(n20049) );
  AND U20923 ( .A(n20050), .B(n20049), .Z(n20173) );
  XNOR U20924 ( .A(n20172), .B(n20173), .Z(n20174) );
  XOR U20925 ( .A(n20175), .B(n20174), .Z(n20148) );
  XOR U20926 ( .A(n20151), .B(n20150), .Z(n20163) );
  XOR U20927 ( .A(n20162), .B(n20163), .Z(n20220) );
  XNOR U20928 ( .A(n20221), .B(n20220), .Z(n20223) );
  XNOR U20929 ( .A(n20222), .B(n20223), .Z(n20102) );
  OR U20930 ( .A(n20052), .B(n20051), .Z(n20056) );
  NANDN U20931 ( .A(n20054), .B(n20053), .Z(n20055) );
  AND U20932 ( .A(n20056), .B(n20055), .Z(n20103) );
  XNOR U20933 ( .A(n20102), .B(n20103), .Z(n20104) );
  XNOR U20934 ( .A(n20105), .B(n20104), .Z(n20099) );
  NANDN U20935 ( .A(n20058), .B(n20057), .Z(n20062) );
  NANDN U20936 ( .A(n20060), .B(n20059), .Z(n20061) );
  NAND U20937 ( .A(n20062), .B(n20061), .Z(n20096) );
  NAND U20938 ( .A(n20064), .B(n20063), .Z(n20068) );
  NAND U20939 ( .A(n20066), .B(n20065), .Z(n20067) );
  NAND U20940 ( .A(n20068), .B(n20067), .Z(n20097) );
  XNOR U20941 ( .A(n20096), .B(n20097), .Z(n20098) );
  XNOR U20942 ( .A(n20099), .B(n20098), .Z(n20093) );
  NANDN U20943 ( .A(n20070), .B(n20069), .Z(n20074) );
  NANDN U20944 ( .A(n20072), .B(n20071), .Z(n20073) );
  NAND U20945 ( .A(n20074), .B(n20073), .Z(n20091) );
  OR U20946 ( .A(n20076), .B(n20075), .Z(n20080) );
  OR U20947 ( .A(n20078), .B(n20077), .Z(n20079) );
  AND U20948 ( .A(n20080), .B(n20079), .Z(n20090) );
  XNOR U20949 ( .A(n20091), .B(n20090), .Z(n20092) );
  XNOR U20950 ( .A(n20093), .B(n20092), .Z(n20086) );
  XOR U20951 ( .A(n20087), .B(n20086), .Z(n20088) );
  XNOR U20952 ( .A(n20089), .B(n20088), .Z(n20226) );
  XNOR U20953 ( .A(n20226), .B(sreg[370]), .Z(n20228) );
  NAND U20954 ( .A(n20081), .B(sreg[369]), .Z(n20085) );
  OR U20955 ( .A(n20083), .B(n20082), .Z(n20084) );
  AND U20956 ( .A(n20085), .B(n20084), .Z(n20227) );
  XOR U20957 ( .A(n20228), .B(n20227), .Z(c[370]) );
  NANDN U20958 ( .A(n20091), .B(n20090), .Z(n20095) );
  NANDN U20959 ( .A(n20093), .B(n20092), .Z(n20094) );
  NAND U20960 ( .A(n20095), .B(n20094), .Z(n20232) );
  NANDN U20961 ( .A(n20097), .B(n20096), .Z(n20101) );
  NAND U20962 ( .A(n20099), .B(n20098), .Z(n20100) );
  NAND U20963 ( .A(n20101), .B(n20100), .Z(n20237) );
  NAND U20964 ( .A(n20103), .B(n20102), .Z(n20107) );
  OR U20965 ( .A(n20105), .B(n20104), .Z(n20106) );
  NAND U20966 ( .A(n20107), .B(n20106), .Z(n20238) );
  XNOR U20967 ( .A(n20237), .B(n20238), .Z(n20239) );
  NANDN U20968 ( .A(n20109), .B(n20108), .Z(n20113) );
  NAND U20969 ( .A(n20111), .B(n20110), .Z(n20112) );
  NAND U20970 ( .A(n20113), .B(n20112), .Z(n20315) );
  XOR U20971 ( .A(b[19]), .B(n22221), .Z(n20259) );
  NANDN U20972 ( .A(n20259), .B(n37934), .Z(n20116) );
  NANDN U20973 ( .A(n20114), .B(n37935), .Z(n20115) );
  NAND U20974 ( .A(n20116), .B(n20115), .Z(n20325) );
  XOR U20975 ( .A(b[27]), .B(a[121]), .Z(n20262) );
  NAND U20976 ( .A(n38423), .B(n20262), .Z(n20119) );
  NAND U20977 ( .A(n20117), .B(n38424), .Z(n20118) );
  NAND U20978 ( .A(n20119), .B(n20118), .Z(n20322) );
  XNOR U20979 ( .A(b[5]), .B(a[143]), .Z(n20265) );
  NANDN U20980 ( .A(n20265), .B(n36587), .Z(n20122) );
  NANDN U20981 ( .A(n20120), .B(n36588), .Z(n20121) );
  AND U20982 ( .A(n20122), .B(n20121), .Z(n20323) );
  XNOR U20983 ( .A(n20322), .B(n20323), .Z(n20324) );
  XNOR U20984 ( .A(n20325), .B(n20324), .Z(n20313) );
  NAND U20985 ( .A(n20123), .B(n37762), .Z(n20125) );
  XNOR U20986 ( .A(b[17]), .B(a[131]), .Z(n20268) );
  NANDN U20987 ( .A(n20268), .B(n37764), .Z(n20124) );
  NAND U20988 ( .A(n20125), .B(n20124), .Z(n20287) );
  XNOR U20989 ( .A(b[31]), .B(a[117]), .Z(n20272) );
  NANDN U20990 ( .A(n20272), .B(n38552), .Z(n20128) );
  NANDN U20991 ( .A(n20126), .B(n38553), .Z(n20127) );
  NAND U20992 ( .A(n20128), .B(n20127), .Z(n20284) );
  OR U20993 ( .A(n20129), .B(n36105), .Z(n20131) );
  XOR U20994 ( .A(b[3]), .B(n24554), .Z(n20275) );
  NANDN U20995 ( .A(n20275), .B(n36107), .Z(n20130) );
  AND U20996 ( .A(n20131), .B(n20130), .Z(n20285) );
  XNOR U20997 ( .A(n20284), .B(n20285), .Z(n20286) );
  XOR U20998 ( .A(n20287), .B(n20286), .Z(n20312) );
  XNOR U20999 ( .A(n20313), .B(n20312), .Z(n20314) );
  XNOR U21000 ( .A(n20315), .B(n20314), .Z(n20250) );
  NANDN U21001 ( .A(n20133), .B(n20132), .Z(n20137) );
  NAND U21002 ( .A(n20135), .B(n20134), .Z(n20136) );
  NAND U21003 ( .A(n20137), .B(n20136), .Z(n20304) );
  NANDN U21004 ( .A(n20139), .B(n20138), .Z(n20143) );
  NAND U21005 ( .A(n20141), .B(n20140), .Z(n20142) );
  NAND U21006 ( .A(n20143), .B(n20142), .Z(n20303) );
  XNOR U21007 ( .A(n20303), .B(n20302), .Z(n20305) );
  XOR U21008 ( .A(n20304), .B(n20305), .Z(n20249) );
  XOR U21009 ( .A(n20250), .B(n20249), .Z(n20251) );
  NANDN U21010 ( .A(n20149), .B(n20148), .Z(n20153) );
  NAND U21011 ( .A(n20151), .B(n20150), .Z(n20152) );
  NAND U21012 ( .A(n20153), .B(n20152), .Z(n20252) );
  XNOR U21013 ( .A(n20251), .B(n20252), .Z(n20366) );
  OR U21014 ( .A(n20155), .B(n20154), .Z(n20159) );
  NANDN U21015 ( .A(n20157), .B(n20156), .Z(n20158) );
  NAND U21016 ( .A(n20159), .B(n20158), .Z(n20365) );
  NANDN U21017 ( .A(n20161), .B(n20160), .Z(n20165) );
  NAND U21018 ( .A(n20163), .B(n20162), .Z(n20164) );
  NAND U21019 ( .A(n20165), .B(n20164), .Z(n20245) );
  NANDN U21020 ( .A(n20167), .B(n20166), .Z(n20171) );
  OR U21021 ( .A(n20169), .B(n20168), .Z(n20170) );
  NAND U21022 ( .A(n20171), .B(n20170), .Z(n20244) );
  NANDN U21023 ( .A(n20173), .B(n20172), .Z(n20177) );
  NAND U21024 ( .A(n20175), .B(n20174), .Z(n20176) );
  NAND U21025 ( .A(n20177), .B(n20176), .Z(n20306) );
  NANDN U21026 ( .A(n20179), .B(n20178), .Z(n20183) );
  NAND U21027 ( .A(n20181), .B(n20180), .Z(n20182) );
  AND U21028 ( .A(n20183), .B(n20182), .Z(n20307) );
  XNOR U21029 ( .A(n20306), .B(n20307), .Z(n20308) );
  XOR U21030 ( .A(b[9]), .B(n23668), .Z(n20328) );
  NANDN U21031 ( .A(n20328), .B(n36925), .Z(n20186) );
  NANDN U21032 ( .A(n20184), .B(n36926), .Z(n20185) );
  NAND U21033 ( .A(n20186), .B(n20185), .Z(n20292) );
  XNOR U21034 ( .A(b[15]), .B(a[133]), .Z(n20331) );
  OR U21035 ( .A(n20331), .B(n37665), .Z(n20189) );
  NAND U21036 ( .A(n20187), .B(n37604), .Z(n20188) );
  AND U21037 ( .A(n20189), .B(n20188), .Z(n20290) );
  XNOR U21038 ( .A(b[21]), .B(a[127]), .Z(n20334) );
  NANDN U21039 ( .A(n20334), .B(n38101), .Z(n20192) );
  NANDN U21040 ( .A(n20190), .B(n38102), .Z(n20191) );
  AND U21041 ( .A(n20192), .B(n20191), .Z(n20291) );
  XOR U21042 ( .A(n20292), .B(n20293), .Z(n20281) );
  XOR U21043 ( .A(b[11]), .B(n23393), .Z(n20337) );
  OR U21044 ( .A(n20337), .B(n37311), .Z(n20195) );
  NANDN U21045 ( .A(n20193), .B(n37218), .Z(n20194) );
  NAND U21046 ( .A(n20195), .B(n20194), .Z(n20279) );
  XOR U21047 ( .A(n1053), .B(a[135]), .Z(n20340) );
  NANDN U21048 ( .A(n20340), .B(n37424), .Z(n20198) );
  NANDN U21049 ( .A(n20196), .B(n37425), .Z(n20197) );
  AND U21050 ( .A(n20198), .B(n20197), .Z(n20278) );
  XNOR U21051 ( .A(n20279), .B(n20278), .Z(n20280) );
  XOR U21052 ( .A(n20281), .B(n20280), .Z(n20298) );
  NAND U21053 ( .A(n38490), .B(n20199), .Z(n20201) );
  XNOR U21054 ( .A(n1058), .B(a[119]), .Z(n20346) );
  NANDN U21055 ( .A(n1048), .B(n20346), .Z(n20200) );
  NAND U21056 ( .A(n20201), .B(n20200), .Z(n20253) );
  NANDN U21057 ( .A(n1059), .B(a[115]), .Z(n20254) );
  XNOR U21058 ( .A(n20253), .B(n20254), .Z(n20256) );
  NANDN U21059 ( .A(n1049), .B(a[147]), .Z(n20202) );
  XNOR U21060 ( .A(b[1]), .B(n20202), .Z(n20204) );
  NANDN U21061 ( .A(b[0]), .B(a[146]), .Z(n20203) );
  AND U21062 ( .A(n20204), .B(n20203), .Z(n20255) );
  XOR U21063 ( .A(n20256), .B(n20255), .Z(n20296) );
  NANDN U21064 ( .A(n20205), .B(n38205), .Z(n20207) );
  XNOR U21065 ( .A(b[23]), .B(a[125]), .Z(n20349) );
  OR U21066 ( .A(n20349), .B(n38268), .Z(n20206) );
  NAND U21067 ( .A(n20207), .B(n20206), .Z(n20319) );
  XNOR U21068 ( .A(b[7]), .B(a[141]), .Z(n20352) );
  NANDN U21069 ( .A(n20352), .B(n36701), .Z(n20210) );
  NAND U21070 ( .A(n20208), .B(n36702), .Z(n20209) );
  NAND U21071 ( .A(n20210), .B(n20209), .Z(n20316) );
  XOR U21072 ( .A(b[25]), .B(a[123]), .Z(n20355) );
  NAND U21073 ( .A(n20355), .B(n38325), .Z(n20213) );
  NAND U21074 ( .A(n20211), .B(n38326), .Z(n20212) );
  AND U21075 ( .A(n20213), .B(n20212), .Z(n20317) );
  XNOR U21076 ( .A(n20316), .B(n20317), .Z(n20318) );
  XNOR U21077 ( .A(n20319), .B(n20318), .Z(n20297) );
  XOR U21078 ( .A(n20296), .B(n20297), .Z(n20299) );
  XNOR U21079 ( .A(n20298), .B(n20299), .Z(n20309) );
  XNOR U21080 ( .A(n20308), .B(n20309), .Z(n20243) );
  XNOR U21081 ( .A(n20244), .B(n20243), .Z(n20246) );
  XNOR U21082 ( .A(n20245), .B(n20246), .Z(n20364) );
  XOR U21083 ( .A(n20365), .B(n20364), .Z(n20367) );
  NAND U21084 ( .A(n20215), .B(n20214), .Z(n20219) );
  NAND U21085 ( .A(n20217), .B(n20216), .Z(n20218) );
  NAND U21086 ( .A(n20219), .B(n20218), .Z(n20359) );
  NAND U21087 ( .A(n20221), .B(n20220), .Z(n20225) );
  NANDN U21088 ( .A(n20223), .B(n20222), .Z(n20224) );
  AND U21089 ( .A(n20225), .B(n20224), .Z(n20358) );
  XNOR U21090 ( .A(n20359), .B(n20358), .Z(n20360) );
  XOR U21091 ( .A(n20361), .B(n20360), .Z(n20240) );
  XOR U21092 ( .A(n20239), .B(n20240), .Z(n20231) );
  XOR U21093 ( .A(n20232), .B(n20231), .Z(n20233) );
  XNOR U21094 ( .A(n20234), .B(n20233), .Z(n20370) );
  XNOR U21095 ( .A(n20370), .B(sreg[371]), .Z(n20372) );
  NAND U21096 ( .A(n20226), .B(sreg[370]), .Z(n20230) );
  OR U21097 ( .A(n20228), .B(n20227), .Z(n20229) );
  AND U21098 ( .A(n20230), .B(n20229), .Z(n20371) );
  XOR U21099 ( .A(n20372), .B(n20371), .Z(c[371]) );
  NAND U21100 ( .A(n20232), .B(n20231), .Z(n20236) );
  NAND U21101 ( .A(n20234), .B(n20233), .Z(n20235) );
  NAND U21102 ( .A(n20236), .B(n20235), .Z(n20378) );
  NANDN U21103 ( .A(n20238), .B(n20237), .Z(n20242) );
  NAND U21104 ( .A(n20240), .B(n20239), .Z(n20241) );
  NAND U21105 ( .A(n20242), .B(n20241), .Z(n20375) );
  NAND U21106 ( .A(n20244), .B(n20243), .Z(n20248) );
  NANDN U21107 ( .A(n20246), .B(n20245), .Z(n20247) );
  NAND U21108 ( .A(n20248), .B(n20247), .Z(n20387) );
  XNOR U21109 ( .A(n20387), .B(n20388), .Z(n20389) );
  NANDN U21110 ( .A(n20254), .B(n20253), .Z(n20258) );
  NAND U21111 ( .A(n20256), .B(n20255), .Z(n20257) );
  NAND U21112 ( .A(n20258), .B(n20257), .Z(n20462) );
  XNOR U21113 ( .A(b[19]), .B(a[130]), .Z(n20405) );
  NANDN U21114 ( .A(n20405), .B(n37934), .Z(n20261) );
  NANDN U21115 ( .A(n20259), .B(n37935), .Z(n20260) );
  NAND U21116 ( .A(n20261), .B(n20260), .Z(n20472) );
  XOR U21117 ( .A(b[27]), .B(a[122]), .Z(n20408) );
  NAND U21118 ( .A(n38423), .B(n20408), .Z(n20264) );
  NAND U21119 ( .A(n20262), .B(n38424), .Z(n20263) );
  NAND U21120 ( .A(n20264), .B(n20263), .Z(n20469) );
  XNOR U21121 ( .A(b[5]), .B(a[144]), .Z(n20411) );
  NANDN U21122 ( .A(n20411), .B(n36587), .Z(n20267) );
  NANDN U21123 ( .A(n20265), .B(n36588), .Z(n20266) );
  AND U21124 ( .A(n20267), .B(n20266), .Z(n20470) );
  XNOR U21125 ( .A(n20469), .B(n20470), .Z(n20471) );
  XNOR U21126 ( .A(n20472), .B(n20471), .Z(n20460) );
  NANDN U21127 ( .A(n20268), .B(n37762), .Z(n20270) );
  XOR U21128 ( .A(b[17]), .B(a[132]), .Z(n20414) );
  NAND U21129 ( .A(n20414), .B(n37764), .Z(n20269) );
  NAND U21130 ( .A(n20270), .B(n20269), .Z(n20432) );
  XOR U21131 ( .A(b[31]), .B(n20271), .Z(n20417) );
  NANDN U21132 ( .A(n20417), .B(n38552), .Z(n20274) );
  NANDN U21133 ( .A(n20272), .B(n38553), .Z(n20273) );
  NAND U21134 ( .A(n20274), .B(n20273), .Z(n20429) );
  OR U21135 ( .A(n20275), .B(n36105), .Z(n20277) );
  XNOR U21136 ( .A(b[3]), .B(a[146]), .Z(n20420) );
  NANDN U21137 ( .A(n20420), .B(n36107), .Z(n20276) );
  AND U21138 ( .A(n20277), .B(n20276), .Z(n20430) );
  XNOR U21139 ( .A(n20429), .B(n20430), .Z(n20431) );
  XOR U21140 ( .A(n20432), .B(n20431), .Z(n20459) );
  XNOR U21141 ( .A(n20460), .B(n20459), .Z(n20461) );
  XNOR U21142 ( .A(n20462), .B(n20461), .Z(n20505) );
  NANDN U21143 ( .A(n20279), .B(n20278), .Z(n20283) );
  NAND U21144 ( .A(n20281), .B(n20280), .Z(n20282) );
  NAND U21145 ( .A(n20283), .B(n20282), .Z(n20450) );
  NANDN U21146 ( .A(n20285), .B(n20284), .Z(n20289) );
  NAND U21147 ( .A(n20287), .B(n20286), .Z(n20288) );
  NAND U21148 ( .A(n20289), .B(n20288), .Z(n20448) );
  OR U21149 ( .A(n20291), .B(n20290), .Z(n20295) );
  NANDN U21150 ( .A(n20293), .B(n20292), .Z(n20294) );
  NAND U21151 ( .A(n20295), .B(n20294), .Z(n20447) );
  XNOR U21152 ( .A(n20450), .B(n20449), .Z(n20506) );
  XNOR U21153 ( .A(n20505), .B(n20506), .Z(n20507) );
  NANDN U21154 ( .A(n20297), .B(n20296), .Z(n20301) );
  OR U21155 ( .A(n20299), .B(n20298), .Z(n20300) );
  AND U21156 ( .A(n20301), .B(n20300), .Z(n20508) );
  XOR U21157 ( .A(n20507), .B(n20508), .Z(n20395) );
  NANDN U21158 ( .A(n20307), .B(n20306), .Z(n20311) );
  NANDN U21159 ( .A(n20309), .B(n20308), .Z(n20310) );
  NAND U21160 ( .A(n20311), .B(n20310), .Z(n20514) );
  NANDN U21161 ( .A(n20317), .B(n20316), .Z(n20321) );
  NAND U21162 ( .A(n20319), .B(n20318), .Z(n20320) );
  NAND U21163 ( .A(n20321), .B(n20320), .Z(n20453) );
  NANDN U21164 ( .A(n20323), .B(n20322), .Z(n20327) );
  NAND U21165 ( .A(n20325), .B(n20324), .Z(n20326) );
  AND U21166 ( .A(n20327), .B(n20326), .Z(n20454) );
  XNOR U21167 ( .A(n20453), .B(n20454), .Z(n20455) );
  XNOR U21168 ( .A(b[9]), .B(a[140]), .Z(n20475) );
  NANDN U21169 ( .A(n20475), .B(n36925), .Z(n20330) );
  NANDN U21170 ( .A(n20328), .B(n36926), .Z(n20329) );
  NAND U21171 ( .A(n20330), .B(n20329), .Z(n20437) );
  XNOR U21172 ( .A(b[15]), .B(a[134]), .Z(n20478) );
  OR U21173 ( .A(n20478), .B(n37665), .Z(n20333) );
  NANDN U21174 ( .A(n20331), .B(n37604), .Z(n20332) );
  AND U21175 ( .A(n20333), .B(n20332), .Z(n20435) );
  XNOR U21176 ( .A(b[21]), .B(a[128]), .Z(n20481) );
  NANDN U21177 ( .A(n20481), .B(n38101), .Z(n20336) );
  NANDN U21178 ( .A(n20334), .B(n38102), .Z(n20335) );
  AND U21179 ( .A(n20336), .B(n20335), .Z(n20436) );
  XOR U21180 ( .A(n20437), .B(n20438), .Z(n20426) );
  XNOR U21181 ( .A(b[11]), .B(a[138]), .Z(n20484) );
  OR U21182 ( .A(n20484), .B(n37311), .Z(n20339) );
  NANDN U21183 ( .A(n20337), .B(n37218), .Z(n20338) );
  NAND U21184 ( .A(n20339), .B(n20338), .Z(n20424) );
  XOR U21185 ( .A(n1053), .B(a[136]), .Z(n20487) );
  NANDN U21186 ( .A(n20487), .B(n37424), .Z(n20342) );
  NANDN U21187 ( .A(n20340), .B(n37425), .Z(n20341) );
  AND U21188 ( .A(n20342), .B(n20341), .Z(n20423) );
  XNOR U21189 ( .A(n20424), .B(n20423), .Z(n20425) );
  XOR U21190 ( .A(n20426), .B(n20425), .Z(n20443) );
  NANDN U21191 ( .A(n1049), .B(a[148]), .Z(n20343) );
  XNOR U21192 ( .A(b[1]), .B(n20343), .Z(n20345) );
  NANDN U21193 ( .A(b[0]), .B(a[147]), .Z(n20344) );
  AND U21194 ( .A(n20345), .B(n20344), .Z(n20401) );
  NAND U21195 ( .A(n38490), .B(n20346), .Z(n20348) );
  XNOR U21196 ( .A(n1058), .B(a[120]), .Z(n20493) );
  NANDN U21197 ( .A(n1048), .B(n20493), .Z(n20347) );
  NAND U21198 ( .A(n20348), .B(n20347), .Z(n20399) );
  NANDN U21199 ( .A(n1059), .B(a[116]), .Z(n20400) );
  XNOR U21200 ( .A(n20399), .B(n20400), .Z(n20402) );
  XOR U21201 ( .A(n20401), .B(n20402), .Z(n20441) );
  NANDN U21202 ( .A(n20349), .B(n38205), .Z(n20351) );
  XNOR U21203 ( .A(b[23]), .B(a[126]), .Z(n20496) );
  OR U21204 ( .A(n20496), .B(n38268), .Z(n20350) );
  NAND U21205 ( .A(n20351), .B(n20350), .Z(n20466) );
  XNOR U21206 ( .A(b[7]), .B(a[142]), .Z(n20499) );
  NANDN U21207 ( .A(n20499), .B(n36701), .Z(n20354) );
  NANDN U21208 ( .A(n20352), .B(n36702), .Z(n20353) );
  NAND U21209 ( .A(n20354), .B(n20353), .Z(n20463) );
  XOR U21210 ( .A(b[25]), .B(a[124]), .Z(n20502) );
  NAND U21211 ( .A(n20502), .B(n38325), .Z(n20357) );
  NAND U21212 ( .A(n20355), .B(n38326), .Z(n20356) );
  AND U21213 ( .A(n20357), .B(n20356), .Z(n20464) );
  XNOR U21214 ( .A(n20463), .B(n20464), .Z(n20465) );
  XNOR U21215 ( .A(n20466), .B(n20465), .Z(n20442) );
  XOR U21216 ( .A(n20441), .B(n20442), .Z(n20444) );
  XNOR U21217 ( .A(n20443), .B(n20444), .Z(n20456) );
  XOR U21218 ( .A(n20455), .B(n20456), .Z(n20512) );
  XNOR U21219 ( .A(n20511), .B(n20512), .Z(n20513) );
  XNOR U21220 ( .A(n20514), .B(n20513), .Z(n20393) );
  XNOR U21221 ( .A(n20394), .B(n20393), .Z(n20396) );
  XNOR U21222 ( .A(n20395), .B(n20396), .Z(n20390) );
  XOR U21223 ( .A(n20389), .B(n20390), .Z(n20384) );
  NANDN U21224 ( .A(n20359), .B(n20358), .Z(n20363) );
  NAND U21225 ( .A(n20361), .B(n20360), .Z(n20362) );
  NAND U21226 ( .A(n20363), .B(n20362), .Z(n20381) );
  NANDN U21227 ( .A(n20365), .B(n20364), .Z(n20369) );
  OR U21228 ( .A(n20367), .B(n20366), .Z(n20368) );
  NAND U21229 ( .A(n20369), .B(n20368), .Z(n20382) );
  XNOR U21230 ( .A(n20381), .B(n20382), .Z(n20383) );
  XNOR U21231 ( .A(n20384), .B(n20383), .Z(n20376) );
  XNOR U21232 ( .A(n20375), .B(n20376), .Z(n20377) );
  XNOR U21233 ( .A(n20378), .B(n20377), .Z(n20517) );
  XNOR U21234 ( .A(n20517), .B(sreg[372]), .Z(n20519) );
  NAND U21235 ( .A(n20370), .B(sreg[371]), .Z(n20374) );
  OR U21236 ( .A(n20372), .B(n20371), .Z(n20373) );
  AND U21237 ( .A(n20374), .B(n20373), .Z(n20518) );
  XOR U21238 ( .A(n20519), .B(n20518), .Z(c[372]) );
  NANDN U21239 ( .A(n20376), .B(n20375), .Z(n20380) );
  NAND U21240 ( .A(n20378), .B(n20377), .Z(n20379) );
  NAND U21241 ( .A(n20380), .B(n20379), .Z(n20525) );
  NANDN U21242 ( .A(n20382), .B(n20381), .Z(n20386) );
  NAND U21243 ( .A(n20384), .B(n20383), .Z(n20385) );
  NAND U21244 ( .A(n20386), .B(n20385), .Z(n20523) );
  NANDN U21245 ( .A(n20388), .B(n20387), .Z(n20392) );
  NANDN U21246 ( .A(n20390), .B(n20389), .Z(n20391) );
  NAND U21247 ( .A(n20392), .B(n20391), .Z(n20529) );
  OR U21248 ( .A(n20394), .B(n20393), .Z(n20398) );
  OR U21249 ( .A(n20396), .B(n20395), .Z(n20397) );
  AND U21250 ( .A(n20398), .B(n20397), .Z(n20528) );
  XNOR U21251 ( .A(n20529), .B(n20528), .Z(n20530) );
  NANDN U21252 ( .A(n20400), .B(n20399), .Z(n20404) );
  NAND U21253 ( .A(n20402), .B(n20401), .Z(n20403) );
  NAND U21254 ( .A(n20404), .B(n20403), .Z(n20609) );
  XOR U21255 ( .A(b[19]), .B(n22518), .Z(n20552) );
  NANDN U21256 ( .A(n20552), .B(n37934), .Z(n20407) );
  NANDN U21257 ( .A(n20405), .B(n37935), .Z(n20406) );
  NAND U21258 ( .A(n20407), .B(n20406), .Z(n20619) );
  XOR U21259 ( .A(b[27]), .B(a[123]), .Z(n20555) );
  NAND U21260 ( .A(n38423), .B(n20555), .Z(n20410) );
  NAND U21261 ( .A(n20408), .B(n38424), .Z(n20409) );
  NAND U21262 ( .A(n20410), .B(n20409), .Z(n20616) );
  XOR U21263 ( .A(b[5]), .B(n24554), .Z(n20558) );
  NANDN U21264 ( .A(n20558), .B(n36587), .Z(n20413) );
  NANDN U21265 ( .A(n20411), .B(n36588), .Z(n20412) );
  AND U21266 ( .A(n20413), .B(n20412), .Z(n20617) );
  XNOR U21267 ( .A(n20616), .B(n20617), .Z(n20618) );
  XNOR U21268 ( .A(n20619), .B(n20618), .Z(n20607) );
  NAND U21269 ( .A(n20414), .B(n37762), .Z(n20416) );
  XOR U21270 ( .A(b[17]), .B(a[133]), .Z(n20561) );
  NAND U21271 ( .A(n20561), .B(n37764), .Z(n20415) );
  NAND U21272 ( .A(n20416), .B(n20415), .Z(n20579) );
  XNOR U21273 ( .A(b[31]), .B(a[119]), .Z(n20564) );
  NANDN U21274 ( .A(n20564), .B(n38552), .Z(n20419) );
  NANDN U21275 ( .A(n20417), .B(n38553), .Z(n20418) );
  NAND U21276 ( .A(n20419), .B(n20418), .Z(n20576) );
  OR U21277 ( .A(n20420), .B(n36105), .Z(n20422) );
  XNOR U21278 ( .A(b[3]), .B(a[147]), .Z(n20567) );
  NANDN U21279 ( .A(n20567), .B(n36107), .Z(n20421) );
  AND U21280 ( .A(n20422), .B(n20421), .Z(n20577) );
  XNOR U21281 ( .A(n20576), .B(n20577), .Z(n20578) );
  XOR U21282 ( .A(n20579), .B(n20578), .Z(n20606) );
  XNOR U21283 ( .A(n20607), .B(n20606), .Z(n20608) );
  XNOR U21284 ( .A(n20609), .B(n20608), .Z(n20652) );
  NANDN U21285 ( .A(n20424), .B(n20423), .Z(n20428) );
  NAND U21286 ( .A(n20426), .B(n20425), .Z(n20427) );
  NAND U21287 ( .A(n20428), .B(n20427), .Z(n20597) );
  NANDN U21288 ( .A(n20430), .B(n20429), .Z(n20434) );
  NAND U21289 ( .A(n20432), .B(n20431), .Z(n20433) );
  NAND U21290 ( .A(n20434), .B(n20433), .Z(n20595) );
  OR U21291 ( .A(n20436), .B(n20435), .Z(n20440) );
  NANDN U21292 ( .A(n20438), .B(n20437), .Z(n20439) );
  NAND U21293 ( .A(n20440), .B(n20439), .Z(n20594) );
  XNOR U21294 ( .A(n20597), .B(n20596), .Z(n20653) );
  XOR U21295 ( .A(n20652), .B(n20653), .Z(n20655) );
  NANDN U21296 ( .A(n20442), .B(n20441), .Z(n20446) );
  OR U21297 ( .A(n20444), .B(n20443), .Z(n20445) );
  NAND U21298 ( .A(n20446), .B(n20445), .Z(n20654) );
  XOR U21299 ( .A(n20655), .B(n20654), .Z(n20542) );
  OR U21300 ( .A(n20448), .B(n20447), .Z(n20452) );
  NAND U21301 ( .A(n20450), .B(n20449), .Z(n20451) );
  NAND U21302 ( .A(n20452), .B(n20451), .Z(n20541) );
  NANDN U21303 ( .A(n20454), .B(n20453), .Z(n20458) );
  NANDN U21304 ( .A(n20456), .B(n20455), .Z(n20457) );
  NAND U21305 ( .A(n20458), .B(n20457), .Z(n20660) );
  NANDN U21306 ( .A(n20464), .B(n20463), .Z(n20468) );
  NAND U21307 ( .A(n20466), .B(n20465), .Z(n20467) );
  NAND U21308 ( .A(n20468), .B(n20467), .Z(n20600) );
  NANDN U21309 ( .A(n20470), .B(n20469), .Z(n20474) );
  NAND U21310 ( .A(n20472), .B(n20471), .Z(n20473) );
  AND U21311 ( .A(n20474), .B(n20473), .Z(n20601) );
  XNOR U21312 ( .A(n20600), .B(n20601), .Z(n20602) );
  XOR U21313 ( .A(n1052), .B(n23961), .Z(n20622) );
  NAND U21314 ( .A(n36925), .B(n20622), .Z(n20477) );
  NANDN U21315 ( .A(n20475), .B(n36926), .Z(n20476) );
  NAND U21316 ( .A(n20477), .B(n20476), .Z(n20584) );
  XNOR U21317 ( .A(b[15]), .B(a[135]), .Z(n20625) );
  OR U21318 ( .A(n20625), .B(n37665), .Z(n20480) );
  NANDN U21319 ( .A(n20478), .B(n37604), .Z(n20479) );
  AND U21320 ( .A(n20480), .B(n20479), .Z(n20582) );
  XOR U21321 ( .A(n1056), .B(n22221), .Z(n20628) );
  NAND U21322 ( .A(n20628), .B(n38101), .Z(n20483) );
  NANDN U21323 ( .A(n20481), .B(n38102), .Z(n20482) );
  AND U21324 ( .A(n20483), .B(n20482), .Z(n20583) );
  XOR U21325 ( .A(n20584), .B(n20585), .Z(n20573) );
  XOR U21326 ( .A(b[11]), .B(n23668), .Z(n20631) );
  OR U21327 ( .A(n20631), .B(n37311), .Z(n20486) );
  NANDN U21328 ( .A(n20484), .B(n37218), .Z(n20485) );
  NAND U21329 ( .A(n20486), .B(n20485), .Z(n20571) );
  XOR U21330 ( .A(n1053), .B(a[137]), .Z(n20634) );
  NANDN U21331 ( .A(n20634), .B(n37424), .Z(n20489) );
  NANDN U21332 ( .A(n20487), .B(n37425), .Z(n20488) );
  AND U21333 ( .A(n20489), .B(n20488), .Z(n20570) );
  XNOR U21334 ( .A(n20571), .B(n20570), .Z(n20572) );
  XOR U21335 ( .A(n20573), .B(n20572), .Z(n20590) );
  NANDN U21336 ( .A(n1049), .B(a[149]), .Z(n20490) );
  XNOR U21337 ( .A(b[1]), .B(n20490), .Z(n20492) );
  NANDN U21338 ( .A(b[0]), .B(a[148]), .Z(n20491) );
  AND U21339 ( .A(n20492), .B(n20491), .Z(n20548) );
  NAND U21340 ( .A(n38490), .B(n20493), .Z(n20495) );
  XNOR U21341 ( .A(n1058), .B(a[121]), .Z(n20640) );
  NANDN U21342 ( .A(n1048), .B(n20640), .Z(n20494) );
  NAND U21343 ( .A(n20495), .B(n20494), .Z(n20546) );
  NANDN U21344 ( .A(n1059), .B(a[117]), .Z(n20547) );
  XNOR U21345 ( .A(n20546), .B(n20547), .Z(n20549) );
  XOR U21346 ( .A(n20548), .B(n20549), .Z(n20588) );
  NANDN U21347 ( .A(n20496), .B(n38205), .Z(n20498) );
  XNOR U21348 ( .A(b[23]), .B(a[127]), .Z(n20643) );
  OR U21349 ( .A(n20643), .B(n38268), .Z(n20497) );
  NAND U21350 ( .A(n20498), .B(n20497), .Z(n20613) );
  XOR U21351 ( .A(b[7]), .B(a[143]), .Z(n20646) );
  NAND U21352 ( .A(n20646), .B(n36701), .Z(n20501) );
  NANDN U21353 ( .A(n20499), .B(n36702), .Z(n20500) );
  NAND U21354 ( .A(n20501), .B(n20500), .Z(n20610) );
  XOR U21355 ( .A(b[25]), .B(a[125]), .Z(n20649) );
  NAND U21356 ( .A(n20649), .B(n38325), .Z(n20504) );
  NAND U21357 ( .A(n20502), .B(n38326), .Z(n20503) );
  AND U21358 ( .A(n20504), .B(n20503), .Z(n20611) );
  XNOR U21359 ( .A(n20610), .B(n20611), .Z(n20612) );
  XNOR U21360 ( .A(n20613), .B(n20612), .Z(n20589) );
  XOR U21361 ( .A(n20588), .B(n20589), .Z(n20591) );
  XNOR U21362 ( .A(n20590), .B(n20591), .Z(n20603) );
  XNOR U21363 ( .A(n20602), .B(n20603), .Z(n20658) );
  XNOR U21364 ( .A(n20659), .B(n20658), .Z(n20661) );
  XNOR U21365 ( .A(n20660), .B(n20661), .Z(n20540) );
  XOR U21366 ( .A(n20541), .B(n20540), .Z(n20543) );
  NANDN U21367 ( .A(n20506), .B(n20505), .Z(n20510) );
  NAND U21368 ( .A(n20508), .B(n20507), .Z(n20509) );
  NAND U21369 ( .A(n20510), .B(n20509), .Z(n20534) );
  NANDN U21370 ( .A(n20512), .B(n20511), .Z(n20516) );
  NAND U21371 ( .A(n20514), .B(n20513), .Z(n20515) );
  NAND U21372 ( .A(n20516), .B(n20515), .Z(n20535) );
  XNOR U21373 ( .A(n20534), .B(n20535), .Z(n20536) );
  XOR U21374 ( .A(n20537), .B(n20536), .Z(n20531) );
  XOR U21375 ( .A(n20530), .B(n20531), .Z(n20522) );
  XOR U21376 ( .A(n20523), .B(n20522), .Z(n20524) );
  XNOR U21377 ( .A(n20525), .B(n20524), .Z(n20664) );
  XNOR U21378 ( .A(n20664), .B(sreg[373]), .Z(n20666) );
  NAND U21379 ( .A(n20517), .B(sreg[372]), .Z(n20521) );
  OR U21380 ( .A(n20519), .B(n20518), .Z(n20520) );
  AND U21381 ( .A(n20521), .B(n20520), .Z(n20665) );
  XOR U21382 ( .A(n20666), .B(n20665), .Z(c[373]) );
  NAND U21383 ( .A(n20523), .B(n20522), .Z(n20527) );
  NAND U21384 ( .A(n20525), .B(n20524), .Z(n20526) );
  NAND U21385 ( .A(n20527), .B(n20526), .Z(n20672) );
  NANDN U21386 ( .A(n20529), .B(n20528), .Z(n20533) );
  NAND U21387 ( .A(n20531), .B(n20530), .Z(n20532) );
  NAND U21388 ( .A(n20533), .B(n20532), .Z(n20670) );
  NANDN U21389 ( .A(n20535), .B(n20534), .Z(n20539) );
  NAND U21390 ( .A(n20537), .B(n20536), .Z(n20538) );
  NAND U21391 ( .A(n20539), .B(n20538), .Z(n20675) );
  NANDN U21392 ( .A(n20541), .B(n20540), .Z(n20545) );
  OR U21393 ( .A(n20543), .B(n20542), .Z(n20544) );
  NAND U21394 ( .A(n20545), .B(n20544), .Z(n20676) );
  XNOR U21395 ( .A(n20675), .B(n20676), .Z(n20677) );
  NANDN U21396 ( .A(n20547), .B(n20546), .Z(n20551) );
  NAND U21397 ( .A(n20549), .B(n20548), .Z(n20550) );
  NAND U21398 ( .A(n20551), .B(n20550), .Z(n20742) );
  XNOR U21399 ( .A(b[19]), .B(a[132]), .Z(n20687) );
  NANDN U21400 ( .A(n20687), .B(n37934), .Z(n20554) );
  NANDN U21401 ( .A(n20552), .B(n37935), .Z(n20553) );
  NAND U21402 ( .A(n20554), .B(n20553), .Z(n20752) );
  XOR U21403 ( .A(b[27]), .B(a[124]), .Z(n20690) );
  NAND U21404 ( .A(n38423), .B(n20690), .Z(n20557) );
  NAND U21405 ( .A(n20555), .B(n38424), .Z(n20556) );
  NAND U21406 ( .A(n20557), .B(n20556), .Z(n20749) );
  XNOR U21407 ( .A(b[5]), .B(a[146]), .Z(n20693) );
  NANDN U21408 ( .A(n20693), .B(n36587), .Z(n20560) );
  NANDN U21409 ( .A(n20558), .B(n36588), .Z(n20559) );
  AND U21410 ( .A(n20560), .B(n20559), .Z(n20750) );
  XNOR U21411 ( .A(n20749), .B(n20750), .Z(n20751) );
  XNOR U21412 ( .A(n20752), .B(n20751), .Z(n20740) );
  NAND U21413 ( .A(n20561), .B(n37762), .Z(n20563) );
  XOR U21414 ( .A(b[17]), .B(a[134]), .Z(n20696) );
  NAND U21415 ( .A(n20696), .B(n37764), .Z(n20562) );
  NAND U21416 ( .A(n20563), .B(n20562), .Z(n20714) );
  XNOR U21417 ( .A(b[31]), .B(a[120]), .Z(n20699) );
  NANDN U21418 ( .A(n20699), .B(n38552), .Z(n20566) );
  NANDN U21419 ( .A(n20564), .B(n38553), .Z(n20565) );
  NAND U21420 ( .A(n20566), .B(n20565), .Z(n20711) );
  OR U21421 ( .A(n20567), .B(n36105), .Z(n20569) );
  XNOR U21422 ( .A(b[3]), .B(a[148]), .Z(n20702) );
  NANDN U21423 ( .A(n20702), .B(n36107), .Z(n20568) );
  AND U21424 ( .A(n20569), .B(n20568), .Z(n20712) );
  XNOR U21425 ( .A(n20711), .B(n20712), .Z(n20713) );
  XOR U21426 ( .A(n20714), .B(n20713), .Z(n20739) );
  XNOR U21427 ( .A(n20740), .B(n20739), .Z(n20741) );
  XNOR U21428 ( .A(n20742), .B(n20741), .Z(n20785) );
  NANDN U21429 ( .A(n20571), .B(n20570), .Z(n20575) );
  NAND U21430 ( .A(n20573), .B(n20572), .Z(n20574) );
  NAND U21431 ( .A(n20575), .B(n20574), .Z(n20730) );
  NANDN U21432 ( .A(n20577), .B(n20576), .Z(n20581) );
  NAND U21433 ( .A(n20579), .B(n20578), .Z(n20580) );
  NAND U21434 ( .A(n20581), .B(n20580), .Z(n20728) );
  OR U21435 ( .A(n20583), .B(n20582), .Z(n20587) );
  NANDN U21436 ( .A(n20585), .B(n20584), .Z(n20586) );
  NAND U21437 ( .A(n20587), .B(n20586), .Z(n20727) );
  XNOR U21438 ( .A(n20730), .B(n20729), .Z(n20786) );
  XOR U21439 ( .A(n20785), .B(n20786), .Z(n20788) );
  NANDN U21440 ( .A(n20589), .B(n20588), .Z(n20593) );
  OR U21441 ( .A(n20591), .B(n20590), .Z(n20592) );
  NAND U21442 ( .A(n20593), .B(n20592), .Z(n20787) );
  XOR U21443 ( .A(n20788), .B(n20787), .Z(n20805) );
  OR U21444 ( .A(n20595), .B(n20594), .Z(n20599) );
  NAND U21445 ( .A(n20597), .B(n20596), .Z(n20598) );
  NAND U21446 ( .A(n20599), .B(n20598), .Z(n20804) );
  NANDN U21447 ( .A(n20601), .B(n20600), .Z(n20605) );
  NANDN U21448 ( .A(n20603), .B(n20602), .Z(n20604) );
  NAND U21449 ( .A(n20605), .B(n20604), .Z(n20793) );
  NANDN U21450 ( .A(n20611), .B(n20610), .Z(n20615) );
  NAND U21451 ( .A(n20613), .B(n20612), .Z(n20614) );
  NAND U21452 ( .A(n20615), .B(n20614), .Z(n20733) );
  NANDN U21453 ( .A(n20617), .B(n20616), .Z(n20621) );
  NAND U21454 ( .A(n20619), .B(n20618), .Z(n20620) );
  AND U21455 ( .A(n20621), .B(n20620), .Z(n20734) );
  XNOR U21456 ( .A(n20733), .B(n20734), .Z(n20735) );
  XOR U21457 ( .A(b[9]), .B(n24120), .Z(n20755) );
  NANDN U21458 ( .A(n20755), .B(n36925), .Z(n20624) );
  NAND U21459 ( .A(n36926), .B(n20622), .Z(n20623) );
  NAND U21460 ( .A(n20624), .B(n20623), .Z(n20719) );
  XNOR U21461 ( .A(n1054), .B(a[136]), .Z(n20758) );
  NANDN U21462 ( .A(n37665), .B(n20758), .Z(n20627) );
  NANDN U21463 ( .A(n20625), .B(n37604), .Z(n20626) );
  NAND U21464 ( .A(n20627), .B(n20626), .Z(n20717) );
  XNOR U21465 ( .A(b[21]), .B(a[130]), .Z(n20761) );
  NANDN U21466 ( .A(n20761), .B(n38101), .Z(n20630) );
  NAND U21467 ( .A(n38102), .B(n20628), .Z(n20629) );
  NAND U21468 ( .A(n20630), .B(n20629), .Z(n20718) );
  XNOR U21469 ( .A(n20717), .B(n20718), .Z(n20720) );
  XOR U21470 ( .A(n20719), .B(n20720), .Z(n20708) );
  XNOR U21471 ( .A(b[11]), .B(a[140]), .Z(n20764) );
  OR U21472 ( .A(n20764), .B(n37311), .Z(n20633) );
  NANDN U21473 ( .A(n20631), .B(n37218), .Z(n20632) );
  NAND U21474 ( .A(n20633), .B(n20632), .Z(n20706) );
  XOR U21475 ( .A(n1053), .B(a[138]), .Z(n20767) );
  NANDN U21476 ( .A(n20767), .B(n37424), .Z(n20636) );
  NANDN U21477 ( .A(n20634), .B(n37425), .Z(n20635) );
  AND U21478 ( .A(n20636), .B(n20635), .Z(n20705) );
  XNOR U21479 ( .A(n20706), .B(n20705), .Z(n20707) );
  XNOR U21480 ( .A(n20708), .B(n20707), .Z(n20724) );
  NANDN U21481 ( .A(n1049), .B(a[150]), .Z(n20637) );
  XNOR U21482 ( .A(b[1]), .B(n20637), .Z(n20639) );
  NANDN U21483 ( .A(b[0]), .B(a[149]), .Z(n20638) );
  AND U21484 ( .A(n20639), .B(n20638), .Z(n20683) );
  NAND U21485 ( .A(n38490), .B(n20640), .Z(n20642) );
  XNOR U21486 ( .A(n1058), .B(a[122]), .Z(n20773) );
  NANDN U21487 ( .A(n1048), .B(n20773), .Z(n20641) );
  NAND U21488 ( .A(n20642), .B(n20641), .Z(n20681) );
  NANDN U21489 ( .A(n1059), .B(a[118]), .Z(n20682) );
  XNOR U21490 ( .A(n20681), .B(n20682), .Z(n20684) );
  XNOR U21491 ( .A(n20683), .B(n20684), .Z(n20722) );
  NANDN U21492 ( .A(n20643), .B(n38205), .Z(n20645) );
  XNOR U21493 ( .A(b[23]), .B(a[128]), .Z(n20776) );
  OR U21494 ( .A(n20776), .B(n38268), .Z(n20644) );
  NAND U21495 ( .A(n20645), .B(n20644), .Z(n20746) );
  XOR U21496 ( .A(b[7]), .B(a[144]), .Z(n20779) );
  NAND U21497 ( .A(n20779), .B(n36701), .Z(n20648) );
  NAND U21498 ( .A(n20646), .B(n36702), .Z(n20647) );
  NAND U21499 ( .A(n20648), .B(n20647), .Z(n20743) );
  XOR U21500 ( .A(b[25]), .B(a[126]), .Z(n20782) );
  NAND U21501 ( .A(n20782), .B(n38325), .Z(n20651) );
  NAND U21502 ( .A(n20649), .B(n38326), .Z(n20650) );
  AND U21503 ( .A(n20651), .B(n20650), .Z(n20744) );
  XNOR U21504 ( .A(n20743), .B(n20744), .Z(n20745) );
  XOR U21505 ( .A(n20746), .B(n20745), .Z(n20721) );
  XOR U21506 ( .A(n20724), .B(n20723), .Z(n20736) );
  XOR U21507 ( .A(n20735), .B(n20736), .Z(n20791) );
  XNOR U21508 ( .A(n20792), .B(n20791), .Z(n20794) );
  XNOR U21509 ( .A(n20793), .B(n20794), .Z(n20803) );
  XOR U21510 ( .A(n20804), .B(n20803), .Z(n20806) );
  NANDN U21511 ( .A(n20653), .B(n20652), .Z(n20657) );
  OR U21512 ( .A(n20655), .B(n20654), .Z(n20656) );
  NAND U21513 ( .A(n20657), .B(n20656), .Z(n20797) );
  NAND U21514 ( .A(n20659), .B(n20658), .Z(n20663) );
  NANDN U21515 ( .A(n20661), .B(n20660), .Z(n20662) );
  NAND U21516 ( .A(n20663), .B(n20662), .Z(n20798) );
  XNOR U21517 ( .A(n20797), .B(n20798), .Z(n20799) );
  XOR U21518 ( .A(n20800), .B(n20799), .Z(n20678) );
  XOR U21519 ( .A(n20677), .B(n20678), .Z(n20669) );
  XOR U21520 ( .A(n20670), .B(n20669), .Z(n20671) );
  XNOR U21521 ( .A(n20672), .B(n20671), .Z(n20809) );
  XNOR U21522 ( .A(n20809), .B(sreg[374]), .Z(n20811) );
  NAND U21523 ( .A(n20664), .B(sreg[373]), .Z(n20668) );
  OR U21524 ( .A(n20666), .B(n20665), .Z(n20667) );
  AND U21525 ( .A(n20668), .B(n20667), .Z(n20810) );
  XOR U21526 ( .A(n20811), .B(n20810), .Z(c[374]) );
  NAND U21527 ( .A(n20670), .B(n20669), .Z(n20674) );
  NAND U21528 ( .A(n20672), .B(n20671), .Z(n20673) );
  NAND U21529 ( .A(n20674), .B(n20673), .Z(n20817) );
  NANDN U21530 ( .A(n20676), .B(n20675), .Z(n20680) );
  NAND U21531 ( .A(n20678), .B(n20677), .Z(n20679) );
  NAND U21532 ( .A(n20680), .B(n20679), .Z(n20815) );
  NANDN U21533 ( .A(n20682), .B(n20681), .Z(n20686) );
  NAND U21534 ( .A(n20684), .B(n20683), .Z(n20685) );
  NAND U21535 ( .A(n20686), .B(n20685), .Z(n20897) );
  XNOR U21536 ( .A(b[19]), .B(a[133]), .Z(n20842) );
  NANDN U21537 ( .A(n20842), .B(n37934), .Z(n20689) );
  NANDN U21538 ( .A(n20687), .B(n37935), .Z(n20688) );
  NAND U21539 ( .A(n20689), .B(n20688), .Z(n20907) );
  XOR U21540 ( .A(b[27]), .B(a[125]), .Z(n20845) );
  NAND U21541 ( .A(n38423), .B(n20845), .Z(n20692) );
  NAND U21542 ( .A(n20690), .B(n38424), .Z(n20691) );
  NAND U21543 ( .A(n20692), .B(n20691), .Z(n20904) );
  XNOR U21544 ( .A(b[5]), .B(a[147]), .Z(n20848) );
  NANDN U21545 ( .A(n20848), .B(n36587), .Z(n20695) );
  NANDN U21546 ( .A(n20693), .B(n36588), .Z(n20694) );
  AND U21547 ( .A(n20695), .B(n20694), .Z(n20905) );
  XNOR U21548 ( .A(n20904), .B(n20905), .Z(n20906) );
  XNOR U21549 ( .A(n20907), .B(n20906), .Z(n20895) );
  NAND U21550 ( .A(n20696), .B(n37762), .Z(n20698) );
  XOR U21551 ( .A(b[17]), .B(a[135]), .Z(n20851) );
  NAND U21552 ( .A(n20851), .B(n37764), .Z(n20697) );
  NAND U21553 ( .A(n20698), .B(n20697), .Z(n20869) );
  XNOR U21554 ( .A(b[31]), .B(a[121]), .Z(n20854) );
  NANDN U21555 ( .A(n20854), .B(n38552), .Z(n20701) );
  NANDN U21556 ( .A(n20699), .B(n38553), .Z(n20700) );
  NAND U21557 ( .A(n20701), .B(n20700), .Z(n20866) );
  OR U21558 ( .A(n20702), .B(n36105), .Z(n20704) );
  XNOR U21559 ( .A(b[3]), .B(a[149]), .Z(n20857) );
  NANDN U21560 ( .A(n20857), .B(n36107), .Z(n20703) );
  AND U21561 ( .A(n20704), .B(n20703), .Z(n20867) );
  XNOR U21562 ( .A(n20866), .B(n20867), .Z(n20868) );
  XOR U21563 ( .A(n20869), .B(n20868), .Z(n20894) );
  XNOR U21564 ( .A(n20895), .B(n20894), .Z(n20896) );
  XNOR U21565 ( .A(n20897), .B(n20896), .Z(n20833) );
  NANDN U21566 ( .A(n20706), .B(n20705), .Z(n20710) );
  NAND U21567 ( .A(n20708), .B(n20707), .Z(n20709) );
  NAND U21568 ( .A(n20710), .B(n20709), .Z(n20886) );
  NANDN U21569 ( .A(n20712), .B(n20711), .Z(n20716) );
  NAND U21570 ( .A(n20714), .B(n20713), .Z(n20715) );
  NAND U21571 ( .A(n20716), .B(n20715), .Z(n20885) );
  XNOR U21572 ( .A(n20885), .B(n20884), .Z(n20887) );
  XOR U21573 ( .A(n20886), .B(n20887), .Z(n20832) );
  XOR U21574 ( .A(n20833), .B(n20832), .Z(n20834) );
  NANDN U21575 ( .A(n20722), .B(n20721), .Z(n20726) );
  NAND U21576 ( .A(n20724), .B(n20723), .Z(n20725) );
  NAND U21577 ( .A(n20726), .B(n20725), .Z(n20835) );
  XNOR U21578 ( .A(n20834), .B(n20835), .Z(n20948) );
  OR U21579 ( .A(n20728), .B(n20727), .Z(n20732) );
  NAND U21580 ( .A(n20730), .B(n20729), .Z(n20731) );
  NAND U21581 ( .A(n20732), .B(n20731), .Z(n20947) );
  NANDN U21582 ( .A(n20734), .B(n20733), .Z(n20738) );
  NAND U21583 ( .A(n20736), .B(n20735), .Z(n20737) );
  NAND U21584 ( .A(n20738), .B(n20737), .Z(n20828) );
  NANDN U21585 ( .A(n20744), .B(n20743), .Z(n20748) );
  NAND U21586 ( .A(n20746), .B(n20745), .Z(n20747) );
  NAND U21587 ( .A(n20748), .B(n20747), .Z(n20888) );
  NANDN U21588 ( .A(n20750), .B(n20749), .Z(n20754) );
  NAND U21589 ( .A(n20752), .B(n20751), .Z(n20753) );
  AND U21590 ( .A(n20754), .B(n20753), .Z(n20889) );
  XNOR U21591 ( .A(n20888), .B(n20889), .Z(n20890) );
  XNOR U21592 ( .A(b[9]), .B(a[143]), .Z(n20910) );
  NANDN U21593 ( .A(n20910), .B(n36925), .Z(n20757) );
  NANDN U21594 ( .A(n20755), .B(n36926), .Z(n20756) );
  NAND U21595 ( .A(n20757), .B(n20756), .Z(n20874) );
  XOR U21596 ( .A(b[15]), .B(n23393), .Z(n20913) );
  OR U21597 ( .A(n20913), .B(n37665), .Z(n20760) );
  NAND U21598 ( .A(n20758), .B(n37604), .Z(n20759) );
  AND U21599 ( .A(n20760), .B(n20759), .Z(n20872) );
  XOR U21600 ( .A(b[21]), .B(n22518), .Z(n20916) );
  NANDN U21601 ( .A(n20916), .B(n38101), .Z(n20763) );
  NANDN U21602 ( .A(n20761), .B(n38102), .Z(n20762) );
  AND U21603 ( .A(n20763), .B(n20762), .Z(n20873) );
  XOR U21604 ( .A(n20874), .B(n20875), .Z(n20863) );
  XOR U21605 ( .A(b[11]), .B(n23961), .Z(n20919) );
  OR U21606 ( .A(n20919), .B(n37311), .Z(n20766) );
  NANDN U21607 ( .A(n20764), .B(n37218), .Z(n20765) );
  NAND U21608 ( .A(n20766), .B(n20765), .Z(n20861) );
  XOR U21609 ( .A(n1053), .B(a[139]), .Z(n20922) );
  NANDN U21610 ( .A(n20922), .B(n37424), .Z(n20769) );
  NANDN U21611 ( .A(n20767), .B(n37425), .Z(n20768) );
  AND U21612 ( .A(n20769), .B(n20768), .Z(n20860) );
  XNOR U21613 ( .A(n20861), .B(n20860), .Z(n20862) );
  XOR U21614 ( .A(n20863), .B(n20862), .Z(n20880) );
  NANDN U21615 ( .A(n1049), .B(a[151]), .Z(n20770) );
  XNOR U21616 ( .A(b[1]), .B(n20770), .Z(n20772) );
  NANDN U21617 ( .A(b[0]), .B(a[150]), .Z(n20771) );
  AND U21618 ( .A(n20772), .B(n20771), .Z(n20838) );
  NAND U21619 ( .A(n38490), .B(n20773), .Z(n20775) );
  XNOR U21620 ( .A(n1058), .B(a[123]), .Z(n20928) );
  NANDN U21621 ( .A(n1048), .B(n20928), .Z(n20774) );
  NAND U21622 ( .A(n20775), .B(n20774), .Z(n20836) );
  NANDN U21623 ( .A(n1059), .B(a[119]), .Z(n20837) );
  XNOR U21624 ( .A(n20836), .B(n20837), .Z(n20839) );
  XOR U21625 ( .A(n20838), .B(n20839), .Z(n20878) );
  NANDN U21626 ( .A(n20776), .B(n38205), .Z(n20778) );
  XOR U21627 ( .A(b[23]), .B(n22221), .Z(n20931) );
  OR U21628 ( .A(n20931), .B(n38268), .Z(n20777) );
  NAND U21629 ( .A(n20778), .B(n20777), .Z(n20901) );
  XNOR U21630 ( .A(b[7]), .B(a[145]), .Z(n20934) );
  NANDN U21631 ( .A(n20934), .B(n36701), .Z(n20781) );
  NAND U21632 ( .A(n20779), .B(n36702), .Z(n20780) );
  NAND U21633 ( .A(n20781), .B(n20780), .Z(n20898) );
  XOR U21634 ( .A(b[25]), .B(a[127]), .Z(n20937) );
  NAND U21635 ( .A(n20937), .B(n38325), .Z(n20784) );
  NAND U21636 ( .A(n20782), .B(n38326), .Z(n20783) );
  AND U21637 ( .A(n20784), .B(n20783), .Z(n20899) );
  XNOR U21638 ( .A(n20898), .B(n20899), .Z(n20900) );
  XNOR U21639 ( .A(n20901), .B(n20900), .Z(n20879) );
  XOR U21640 ( .A(n20878), .B(n20879), .Z(n20881) );
  XNOR U21641 ( .A(n20880), .B(n20881), .Z(n20891) );
  XNOR U21642 ( .A(n20890), .B(n20891), .Z(n20826) );
  XNOR U21643 ( .A(n20827), .B(n20826), .Z(n20829) );
  XNOR U21644 ( .A(n20828), .B(n20829), .Z(n20946) );
  XOR U21645 ( .A(n20947), .B(n20946), .Z(n20949) );
  NANDN U21646 ( .A(n20786), .B(n20785), .Z(n20790) );
  OR U21647 ( .A(n20788), .B(n20787), .Z(n20789) );
  NAND U21648 ( .A(n20790), .B(n20789), .Z(n20940) );
  NAND U21649 ( .A(n20792), .B(n20791), .Z(n20796) );
  NANDN U21650 ( .A(n20794), .B(n20793), .Z(n20795) );
  NAND U21651 ( .A(n20796), .B(n20795), .Z(n20941) );
  XNOR U21652 ( .A(n20940), .B(n20941), .Z(n20942) );
  XOR U21653 ( .A(n20943), .B(n20942), .Z(n20822) );
  NANDN U21654 ( .A(n20798), .B(n20797), .Z(n20802) );
  NAND U21655 ( .A(n20800), .B(n20799), .Z(n20801) );
  NAND U21656 ( .A(n20802), .B(n20801), .Z(n20820) );
  NANDN U21657 ( .A(n20804), .B(n20803), .Z(n20808) );
  OR U21658 ( .A(n20806), .B(n20805), .Z(n20807) );
  NAND U21659 ( .A(n20808), .B(n20807), .Z(n20821) );
  XNOR U21660 ( .A(n20820), .B(n20821), .Z(n20823) );
  XOR U21661 ( .A(n20822), .B(n20823), .Z(n20814) );
  XOR U21662 ( .A(n20815), .B(n20814), .Z(n20816) );
  XNOR U21663 ( .A(n20817), .B(n20816), .Z(n20952) );
  XNOR U21664 ( .A(n20952), .B(sreg[375]), .Z(n20954) );
  NAND U21665 ( .A(n20809), .B(sreg[374]), .Z(n20813) );
  OR U21666 ( .A(n20811), .B(n20810), .Z(n20812) );
  AND U21667 ( .A(n20813), .B(n20812), .Z(n20953) );
  XOR U21668 ( .A(n20954), .B(n20953), .Z(c[375]) );
  NAND U21669 ( .A(n20815), .B(n20814), .Z(n20819) );
  NAND U21670 ( .A(n20817), .B(n20816), .Z(n20818) );
  NAND U21671 ( .A(n20819), .B(n20818), .Z(n20960) );
  NANDN U21672 ( .A(n20821), .B(n20820), .Z(n20825) );
  NAND U21673 ( .A(n20823), .B(n20822), .Z(n20824) );
  NAND U21674 ( .A(n20825), .B(n20824), .Z(n20957) );
  NAND U21675 ( .A(n20827), .B(n20826), .Z(n20831) );
  NANDN U21676 ( .A(n20829), .B(n20828), .Z(n20830) );
  NAND U21677 ( .A(n20831), .B(n20830), .Z(n20969) );
  XNOR U21678 ( .A(n20969), .B(n20970), .Z(n20971) );
  NANDN U21679 ( .A(n20837), .B(n20836), .Z(n20841) );
  NAND U21680 ( .A(n20839), .B(n20838), .Z(n20840) );
  NAND U21681 ( .A(n20841), .B(n20840), .Z(n21044) );
  XNOR U21682 ( .A(b[19]), .B(a[134]), .Z(n20987) );
  NANDN U21683 ( .A(n20987), .B(n37934), .Z(n20844) );
  NANDN U21684 ( .A(n20842), .B(n37935), .Z(n20843) );
  NAND U21685 ( .A(n20844), .B(n20843), .Z(n21054) );
  XOR U21686 ( .A(b[27]), .B(a[126]), .Z(n20990) );
  NAND U21687 ( .A(n38423), .B(n20990), .Z(n20847) );
  NAND U21688 ( .A(n20845), .B(n38424), .Z(n20846) );
  NAND U21689 ( .A(n20847), .B(n20846), .Z(n21051) );
  XNOR U21690 ( .A(b[5]), .B(a[148]), .Z(n20993) );
  NANDN U21691 ( .A(n20993), .B(n36587), .Z(n20850) );
  NANDN U21692 ( .A(n20848), .B(n36588), .Z(n20849) );
  AND U21693 ( .A(n20850), .B(n20849), .Z(n21052) );
  XNOR U21694 ( .A(n21051), .B(n21052), .Z(n21053) );
  XNOR U21695 ( .A(n21054), .B(n21053), .Z(n21042) );
  NAND U21696 ( .A(n20851), .B(n37762), .Z(n20853) );
  XOR U21697 ( .A(b[17]), .B(a[136]), .Z(n20996) );
  NAND U21698 ( .A(n20996), .B(n37764), .Z(n20852) );
  NAND U21699 ( .A(n20853), .B(n20852), .Z(n21014) );
  XNOR U21700 ( .A(b[31]), .B(a[122]), .Z(n20999) );
  NANDN U21701 ( .A(n20999), .B(n38552), .Z(n20856) );
  NANDN U21702 ( .A(n20854), .B(n38553), .Z(n20855) );
  NAND U21703 ( .A(n20856), .B(n20855), .Z(n21011) );
  OR U21704 ( .A(n20857), .B(n36105), .Z(n20859) );
  XNOR U21705 ( .A(b[3]), .B(a[150]), .Z(n21002) );
  NANDN U21706 ( .A(n21002), .B(n36107), .Z(n20858) );
  AND U21707 ( .A(n20859), .B(n20858), .Z(n21012) );
  XNOR U21708 ( .A(n21011), .B(n21012), .Z(n21013) );
  XOR U21709 ( .A(n21014), .B(n21013), .Z(n21041) );
  XNOR U21710 ( .A(n21042), .B(n21041), .Z(n21043) );
  XNOR U21711 ( .A(n21044), .B(n21043), .Z(n21087) );
  NANDN U21712 ( .A(n20861), .B(n20860), .Z(n20865) );
  NAND U21713 ( .A(n20863), .B(n20862), .Z(n20864) );
  NAND U21714 ( .A(n20865), .B(n20864), .Z(n21032) );
  NANDN U21715 ( .A(n20867), .B(n20866), .Z(n20871) );
  NAND U21716 ( .A(n20869), .B(n20868), .Z(n20870) );
  NAND U21717 ( .A(n20871), .B(n20870), .Z(n21030) );
  OR U21718 ( .A(n20873), .B(n20872), .Z(n20877) );
  NANDN U21719 ( .A(n20875), .B(n20874), .Z(n20876) );
  NAND U21720 ( .A(n20877), .B(n20876), .Z(n21029) );
  XNOR U21721 ( .A(n21032), .B(n21031), .Z(n21088) );
  XNOR U21722 ( .A(n21087), .B(n21088), .Z(n21089) );
  NANDN U21723 ( .A(n20879), .B(n20878), .Z(n20883) );
  OR U21724 ( .A(n20881), .B(n20880), .Z(n20882) );
  AND U21725 ( .A(n20883), .B(n20882), .Z(n21090) );
  XOR U21726 ( .A(n21089), .B(n21090), .Z(n20977) );
  NANDN U21727 ( .A(n20889), .B(n20888), .Z(n20893) );
  NANDN U21728 ( .A(n20891), .B(n20890), .Z(n20892) );
  NAND U21729 ( .A(n20893), .B(n20892), .Z(n21096) );
  NANDN U21730 ( .A(n20899), .B(n20898), .Z(n20903) );
  NAND U21731 ( .A(n20901), .B(n20900), .Z(n20902) );
  NAND U21732 ( .A(n20903), .B(n20902), .Z(n21035) );
  NANDN U21733 ( .A(n20905), .B(n20904), .Z(n20909) );
  NAND U21734 ( .A(n20907), .B(n20906), .Z(n20908) );
  AND U21735 ( .A(n20909), .B(n20908), .Z(n21036) );
  XNOR U21736 ( .A(n21035), .B(n21036), .Z(n21037) );
  XNOR U21737 ( .A(b[9]), .B(a[144]), .Z(n21057) );
  NANDN U21738 ( .A(n21057), .B(n36925), .Z(n20912) );
  NANDN U21739 ( .A(n20910), .B(n36926), .Z(n20911) );
  NAND U21740 ( .A(n20912), .B(n20911), .Z(n21019) );
  XNOR U21741 ( .A(b[15]), .B(a[138]), .Z(n21060) );
  OR U21742 ( .A(n21060), .B(n37665), .Z(n20915) );
  NANDN U21743 ( .A(n20913), .B(n37604), .Z(n20914) );
  AND U21744 ( .A(n20915), .B(n20914), .Z(n21017) );
  XNOR U21745 ( .A(b[21]), .B(a[132]), .Z(n21063) );
  NANDN U21746 ( .A(n21063), .B(n38101), .Z(n20918) );
  NANDN U21747 ( .A(n20916), .B(n38102), .Z(n20917) );
  AND U21748 ( .A(n20918), .B(n20917), .Z(n21018) );
  XOR U21749 ( .A(n21019), .B(n21020), .Z(n21008) );
  XOR U21750 ( .A(b[11]), .B(n24120), .Z(n21066) );
  OR U21751 ( .A(n21066), .B(n37311), .Z(n20921) );
  NANDN U21752 ( .A(n20919), .B(n37218), .Z(n20920) );
  NAND U21753 ( .A(n20921), .B(n20920), .Z(n21006) );
  XOR U21754 ( .A(n1053), .B(a[140]), .Z(n21069) );
  NANDN U21755 ( .A(n21069), .B(n37424), .Z(n20924) );
  NANDN U21756 ( .A(n20922), .B(n37425), .Z(n20923) );
  AND U21757 ( .A(n20924), .B(n20923), .Z(n21005) );
  XNOR U21758 ( .A(n21006), .B(n21005), .Z(n21007) );
  XOR U21759 ( .A(n21008), .B(n21007), .Z(n21025) );
  ANDN U21760 ( .B(a[152]), .A(n1049), .Z(n20925) );
  XOR U21761 ( .A(b[1]), .B(n20925), .Z(n20927) );
  IV U21762 ( .A(a[151]), .Z(n25435) );
  NANDN U21763 ( .A(n25435), .B(n1049), .Z(n20926) );
  NAND U21764 ( .A(n20927), .B(n20926), .Z(n20984) );
  NAND U21765 ( .A(n38490), .B(n20928), .Z(n20930) );
  XNOR U21766 ( .A(n1058), .B(a[124]), .Z(n21075) );
  NANDN U21767 ( .A(n1048), .B(n21075), .Z(n20929) );
  NAND U21768 ( .A(n20930), .B(n20929), .Z(n20981) );
  NANDN U21769 ( .A(n1059), .B(a[120]), .Z(n20982) );
  XNOR U21770 ( .A(n20981), .B(n20982), .Z(n20983) );
  XNOR U21771 ( .A(n20984), .B(n20983), .Z(n21023) );
  NANDN U21772 ( .A(n20931), .B(n38205), .Z(n20933) );
  XNOR U21773 ( .A(b[23]), .B(a[130]), .Z(n21078) );
  OR U21774 ( .A(n21078), .B(n38268), .Z(n20932) );
  NAND U21775 ( .A(n20933), .B(n20932), .Z(n21048) );
  XOR U21776 ( .A(b[7]), .B(a[146]), .Z(n21081) );
  NAND U21777 ( .A(n21081), .B(n36701), .Z(n20936) );
  NANDN U21778 ( .A(n20934), .B(n36702), .Z(n20935) );
  NAND U21779 ( .A(n20936), .B(n20935), .Z(n21045) );
  XOR U21780 ( .A(b[25]), .B(a[128]), .Z(n21084) );
  NAND U21781 ( .A(n21084), .B(n38325), .Z(n20939) );
  NAND U21782 ( .A(n20937), .B(n38326), .Z(n20938) );
  AND U21783 ( .A(n20939), .B(n20938), .Z(n21046) );
  XNOR U21784 ( .A(n21045), .B(n21046), .Z(n21047) );
  XNOR U21785 ( .A(n21048), .B(n21047), .Z(n21024) );
  XOR U21786 ( .A(n21023), .B(n21024), .Z(n21026) );
  XNOR U21787 ( .A(n21025), .B(n21026), .Z(n21038) );
  XOR U21788 ( .A(n21037), .B(n21038), .Z(n21094) );
  XNOR U21789 ( .A(n21093), .B(n21094), .Z(n21095) );
  XNOR U21790 ( .A(n21096), .B(n21095), .Z(n20975) );
  XNOR U21791 ( .A(n20976), .B(n20975), .Z(n20978) );
  XNOR U21792 ( .A(n20977), .B(n20978), .Z(n20972) );
  XOR U21793 ( .A(n20971), .B(n20972), .Z(n20966) );
  NANDN U21794 ( .A(n20941), .B(n20940), .Z(n20945) );
  NAND U21795 ( .A(n20943), .B(n20942), .Z(n20944) );
  NAND U21796 ( .A(n20945), .B(n20944), .Z(n20963) );
  NANDN U21797 ( .A(n20947), .B(n20946), .Z(n20951) );
  OR U21798 ( .A(n20949), .B(n20948), .Z(n20950) );
  NAND U21799 ( .A(n20951), .B(n20950), .Z(n20964) );
  XNOR U21800 ( .A(n20963), .B(n20964), .Z(n20965) );
  XNOR U21801 ( .A(n20966), .B(n20965), .Z(n20958) );
  XNOR U21802 ( .A(n20957), .B(n20958), .Z(n20959) );
  XNOR U21803 ( .A(n20960), .B(n20959), .Z(n21099) );
  XNOR U21804 ( .A(n21099), .B(sreg[376]), .Z(n21101) );
  NAND U21805 ( .A(n20952), .B(sreg[375]), .Z(n20956) );
  OR U21806 ( .A(n20954), .B(n20953), .Z(n20955) );
  AND U21807 ( .A(n20956), .B(n20955), .Z(n21100) );
  XOR U21808 ( .A(n21101), .B(n21100), .Z(c[376]) );
  NANDN U21809 ( .A(n20958), .B(n20957), .Z(n20962) );
  NAND U21810 ( .A(n20960), .B(n20959), .Z(n20961) );
  NAND U21811 ( .A(n20962), .B(n20961), .Z(n21107) );
  NANDN U21812 ( .A(n20964), .B(n20963), .Z(n20968) );
  NAND U21813 ( .A(n20966), .B(n20965), .Z(n20967) );
  NAND U21814 ( .A(n20968), .B(n20967), .Z(n21105) );
  NANDN U21815 ( .A(n20970), .B(n20969), .Z(n20974) );
  NANDN U21816 ( .A(n20972), .B(n20971), .Z(n20973) );
  NAND U21817 ( .A(n20974), .B(n20973), .Z(n21111) );
  OR U21818 ( .A(n20976), .B(n20975), .Z(n20980) );
  OR U21819 ( .A(n20978), .B(n20977), .Z(n20979) );
  AND U21820 ( .A(n20980), .B(n20979), .Z(n21110) );
  XNOR U21821 ( .A(n21111), .B(n21110), .Z(n21112) );
  NANDN U21822 ( .A(n20982), .B(n20981), .Z(n20986) );
  NANDN U21823 ( .A(n20984), .B(n20983), .Z(n20985) );
  NAND U21824 ( .A(n20986), .B(n20985), .Z(n21179) );
  XNOR U21825 ( .A(b[19]), .B(a[135]), .Z(n21122) );
  NANDN U21826 ( .A(n21122), .B(n37934), .Z(n20989) );
  NANDN U21827 ( .A(n20987), .B(n37935), .Z(n20988) );
  NAND U21828 ( .A(n20989), .B(n20988), .Z(n21189) );
  XOR U21829 ( .A(b[27]), .B(a[127]), .Z(n21125) );
  NAND U21830 ( .A(n38423), .B(n21125), .Z(n20992) );
  NAND U21831 ( .A(n20990), .B(n38424), .Z(n20991) );
  NAND U21832 ( .A(n20992), .B(n20991), .Z(n21186) );
  XNOR U21833 ( .A(b[5]), .B(a[149]), .Z(n21128) );
  NANDN U21834 ( .A(n21128), .B(n36587), .Z(n20995) );
  NANDN U21835 ( .A(n20993), .B(n36588), .Z(n20994) );
  AND U21836 ( .A(n20995), .B(n20994), .Z(n21187) );
  XNOR U21837 ( .A(n21186), .B(n21187), .Z(n21188) );
  XNOR U21838 ( .A(n21189), .B(n21188), .Z(n21177) );
  NAND U21839 ( .A(n20996), .B(n37762), .Z(n20998) );
  XNOR U21840 ( .A(b[17]), .B(a[137]), .Z(n21131) );
  NANDN U21841 ( .A(n21131), .B(n37764), .Z(n20997) );
  NAND U21842 ( .A(n20998), .B(n20997), .Z(n21149) );
  XNOR U21843 ( .A(b[31]), .B(a[123]), .Z(n21134) );
  NANDN U21844 ( .A(n21134), .B(n38552), .Z(n21001) );
  NANDN U21845 ( .A(n20999), .B(n38553), .Z(n21000) );
  NAND U21846 ( .A(n21001), .B(n21000), .Z(n21146) );
  OR U21847 ( .A(n21002), .B(n36105), .Z(n21004) );
  XOR U21848 ( .A(b[3]), .B(n25435), .Z(n21137) );
  NANDN U21849 ( .A(n21137), .B(n36107), .Z(n21003) );
  AND U21850 ( .A(n21004), .B(n21003), .Z(n21147) );
  XNOR U21851 ( .A(n21146), .B(n21147), .Z(n21148) );
  XOR U21852 ( .A(n21149), .B(n21148), .Z(n21176) );
  XNOR U21853 ( .A(n21177), .B(n21176), .Z(n21178) );
  XNOR U21854 ( .A(n21179), .B(n21178), .Z(n21222) );
  NANDN U21855 ( .A(n21006), .B(n21005), .Z(n21010) );
  NAND U21856 ( .A(n21008), .B(n21007), .Z(n21009) );
  NAND U21857 ( .A(n21010), .B(n21009), .Z(n21167) );
  NANDN U21858 ( .A(n21012), .B(n21011), .Z(n21016) );
  NAND U21859 ( .A(n21014), .B(n21013), .Z(n21015) );
  NAND U21860 ( .A(n21016), .B(n21015), .Z(n21165) );
  OR U21861 ( .A(n21018), .B(n21017), .Z(n21022) );
  NANDN U21862 ( .A(n21020), .B(n21019), .Z(n21021) );
  NAND U21863 ( .A(n21022), .B(n21021), .Z(n21164) );
  XNOR U21864 ( .A(n21167), .B(n21166), .Z(n21223) );
  XOR U21865 ( .A(n21222), .B(n21223), .Z(n21225) );
  NANDN U21866 ( .A(n21024), .B(n21023), .Z(n21028) );
  OR U21867 ( .A(n21026), .B(n21025), .Z(n21027) );
  NAND U21868 ( .A(n21028), .B(n21027), .Z(n21224) );
  XOR U21869 ( .A(n21225), .B(n21224), .Z(n21242) );
  OR U21870 ( .A(n21030), .B(n21029), .Z(n21034) );
  NAND U21871 ( .A(n21032), .B(n21031), .Z(n21033) );
  NAND U21872 ( .A(n21034), .B(n21033), .Z(n21241) );
  NANDN U21873 ( .A(n21036), .B(n21035), .Z(n21040) );
  NANDN U21874 ( .A(n21038), .B(n21037), .Z(n21039) );
  NAND U21875 ( .A(n21040), .B(n21039), .Z(n21230) );
  NANDN U21876 ( .A(n21046), .B(n21045), .Z(n21050) );
  NAND U21877 ( .A(n21048), .B(n21047), .Z(n21049) );
  NAND U21878 ( .A(n21050), .B(n21049), .Z(n21170) );
  NANDN U21879 ( .A(n21052), .B(n21051), .Z(n21056) );
  NAND U21880 ( .A(n21054), .B(n21053), .Z(n21055) );
  AND U21881 ( .A(n21056), .B(n21055), .Z(n21171) );
  XNOR U21882 ( .A(n21170), .B(n21171), .Z(n21172) );
  XOR U21883 ( .A(n1052), .B(n24554), .Z(n21192) );
  NAND U21884 ( .A(n36925), .B(n21192), .Z(n21059) );
  NANDN U21885 ( .A(n21057), .B(n36926), .Z(n21058) );
  NAND U21886 ( .A(n21059), .B(n21058), .Z(n21154) );
  XOR U21887 ( .A(b[15]), .B(n23668), .Z(n21195) );
  OR U21888 ( .A(n21195), .B(n37665), .Z(n21062) );
  NANDN U21889 ( .A(n21060), .B(n37604), .Z(n21061) );
  AND U21890 ( .A(n21062), .B(n21061), .Z(n21152) );
  XNOR U21891 ( .A(n1056), .B(a[133]), .Z(n21198) );
  NAND U21892 ( .A(n21198), .B(n38101), .Z(n21065) );
  NANDN U21893 ( .A(n21063), .B(n38102), .Z(n21064) );
  AND U21894 ( .A(n21065), .B(n21064), .Z(n21153) );
  XOR U21895 ( .A(n21154), .B(n21155), .Z(n21143) );
  XNOR U21896 ( .A(b[11]), .B(a[143]), .Z(n21201) );
  OR U21897 ( .A(n21201), .B(n37311), .Z(n21068) );
  NANDN U21898 ( .A(n21066), .B(n37218), .Z(n21067) );
  NAND U21899 ( .A(n21068), .B(n21067), .Z(n21141) );
  XOR U21900 ( .A(n1053), .B(a[141]), .Z(n21204) );
  NANDN U21901 ( .A(n21204), .B(n37424), .Z(n21071) );
  NANDN U21902 ( .A(n21069), .B(n37425), .Z(n21070) );
  AND U21903 ( .A(n21071), .B(n21070), .Z(n21140) );
  XNOR U21904 ( .A(n21141), .B(n21140), .Z(n21142) );
  XOR U21905 ( .A(n21143), .B(n21142), .Z(n21160) );
  NANDN U21906 ( .A(n1049), .B(a[153]), .Z(n21072) );
  XNOR U21907 ( .A(b[1]), .B(n21072), .Z(n21074) );
  IV U21908 ( .A(a[152]), .Z(n25213) );
  NANDN U21909 ( .A(n25213), .B(n1049), .Z(n21073) );
  AND U21910 ( .A(n21074), .B(n21073), .Z(n21118) );
  NAND U21911 ( .A(n38490), .B(n21075), .Z(n21077) );
  XNOR U21912 ( .A(n1058), .B(a[125]), .Z(n21210) );
  NANDN U21913 ( .A(n1048), .B(n21210), .Z(n21076) );
  NAND U21914 ( .A(n21077), .B(n21076), .Z(n21116) );
  NANDN U21915 ( .A(n1059), .B(a[121]), .Z(n21117) );
  XNOR U21916 ( .A(n21116), .B(n21117), .Z(n21119) );
  XOR U21917 ( .A(n21118), .B(n21119), .Z(n21158) );
  NANDN U21918 ( .A(n21078), .B(n38205), .Z(n21080) );
  XOR U21919 ( .A(b[23]), .B(n22518), .Z(n21213) );
  OR U21920 ( .A(n21213), .B(n38268), .Z(n21079) );
  NAND U21921 ( .A(n21080), .B(n21079), .Z(n21183) );
  XOR U21922 ( .A(b[7]), .B(a[147]), .Z(n21216) );
  NAND U21923 ( .A(n21216), .B(n36701), .Z(n21083) );
  NAND U21924 ( .A(n21081), .B(n36702), .Z(n21082) );
  NAND U21925 ( .A(n21083), .B(n21082), .Z(n21180) );
  XNOR U21926 ( .A(b[25]), .B(a[129]), .Z(n21219) );
  NANDN U21927 ( .A(n21219), .B(n38325), .Z(n21086) );
  NAND U21928 ( .A(n21084), .B(n38326), .Z(n21085) );
  AND U21929 ( .A(n21086), .B(n21085), .Z(n21181) );
  XNOR U21930 ( .A(n21180), .B(n21181), .Z(n21182) );
  XNOR U21931 ( .A(n21183), .B(n21182), .Z(n21159) );
  XOR U21932 ( .A(n21158), .B(n21159), .Z(n21161) );
  XNOR U21933 ( .A(n21160), .B(n21161), .Z(n21173) );
  XNOR U21934 ( .A(n21172), .B(n21173), .Z(n21228) );
  XNOR U21935 ( .A(n21229), .B(n21228), .Z(n21231) );
  XNOR U21936 ( .A(n21230), .B(n21231), .Z(n21240) );
  XOR U21937 ( .A(n21241), .B(n21240), .Z(n21243) );
  NANDN U21938 ( .A(n21088), .B(n21087), .Z(n21092) );
  NAND U21939 ( .A(n21090), .B(n21089), .Z(n21091) );
  NAND U21940 ( .A(n21092), .B(n21091), .Z(n21234) );
  NANDN U21941 ( .A(n21094), .B(n21093), .Z(n21098) );
  NAND U21942 ( .A(n21096), .B(n21095), .Z(n21097) );
  NAND U21943 ( .A(n21098), .B(n21097), .Z(n21235) );
  XNOR U21944 ( .A(n21234), .B(n21235), .Z(n21236) );
  XOR U21945 ( .A(n21237), .B(n21236), .Z(n21113) );
  XOR U21946 ( .A(n21112), .B(n21113), .Z(n21104) );
  XOR U21947 ( .A(n21105), .B(n21104), .Z(n21106) );
  XNOR U21948 ( .A(n21107), .B(n21106), .Z(n21246) );
  XNOR U21949 ( .A(n21246), .B(sreg[377]), .Z(n21248) );
  NAND U21950 ( .A(n21099), .B(sreg[376]), .Z(n21103) );
  OR U21951 ( .A(n21101), .B(n21100), .Z(n21102) );
  AND U21952 ( .A(n21103), .B(n21102), .Z(n21247) );
  XOR U21953 ( .A(n21248), .B(n21247), .Z(c[377]) );
  NAND U21954 ( .A(n21105), .B(n21104), .Z(n21109) );
  NAND U21955 ( .A(n21107), .B(n21106), .Z(n21108) );
  NAND U21956 ( .A(n21109), .B(n21108), .Z(n21254) );
  NANDN U21957 ( .A(n21111), .B(n21110), .Z(n21115) );
  NAND U21958 ( .A(n21113), .B(n21112), .Z(n21114) );
  NAND U21959 ( .A(n21115), .B(n21114), .Z(n21252) );
  NANDN U21960 ( .A(n21117), .B(n21116), .Z(n21121) );
  NAND U21961 ( .A(n21119), .B(n21118), .Z(n21120) );
  NAND U21962 ( .A(n21121), .B(n21120), .Z(n21324) );
  XNOR U21963 ( .A(b[19]), .B(a[136]), .Z(n21269) );
  NANDN U21964 ( .A(n21269), .B(n37934), .Z(n21124) );
  NANDN U21965 ( .A(n21122), .B(n37935), .Z(n21123) );
  NAND U21966 ( .A(n21124), .B(n21123), .Z(n21334) );
  XOR U21967 ( .A(b[27]), .B(a[128]), .Z(n21272) );
  NAND U21968 ( .A(n38423), .B(n21272), .Z(n21127) );
  NAND U21969 ( .A(n21125), .B(n38424), .Z(n21126) );
  NAND U21970 ( .A(n21127), .B(n21126), .Z(n21331) );
  XNOR U21971 ( .A(b[5]), .B(a[150]), .Z(n21275) );
  NANDN U21972 ( .A(n21275), .B(n36587), .Z(n21130) );
  NANDN U21973 ( .A(n21128), .B(n36588), .Z(n21129) );
  AND U21974 ( .A(n21130), .B(n21129), .Z(n21332) );
  XNOR U21975 ( .A(n21331), .B(n21332), .Z(n21333) );
  XNOR U21976 ( .A(n21334), .B(n21333), .Z(n21322) );
  NANDN U21977 ( .A(n21131), .B(n37762), .Z(n21133) );
  XOR U21978 ( .A(b[17]), .B(a[138]), .Z(n21278) );
  NAND U21979 ( .A(n21278), .B(n37764), .Z(n21132) );
  NAND U21980 ( .A(n21133), .B(n21132), .Z(n21296) );
  XNOR U21981 ( .A(b[31]), .B(a[124]), .Z(n21281) );
  NANDN U21982 ( .A(n21281), .B(n38552), .Z(n21136) );
  NANDN U21983 ( .A(n21134), .B(n38553), .Z(n21135) );
  NAND U21984 ( .A(n21136), .B(n21135), .Z(n21293) );
  OR U21985 ( .A(n21137), .B(n36105), .Z(n21139) );
  XOR U21986 ( .A(b[3]), .B(n25213), .Z(n21284) );
  NANDN U21987 ( .A(n21284), .B(n36107), .Z(n21138) );
  AND U21988 ( .A(n21139), .B(n21138), .Z(n21294) );
  XNOR U21989 ( .A(n21293), .B(n21294), .Z(n21295) );
  XOR U21990 ( .A(n21296), .B(n21295), .Z(n21321) );
  XNOR U21991 ( .A(n21322), .B(n21321), .Z(n21323) );
  XNOR U21992 ( .A(n21324), .B(n21323), .Z(n21367) );
  NANDN U21993 ( .A(n21141), .B(n21140), .Z(n21145) );
  NAND U21994 ( .A(n21143), .B(n21142), .Z(n21144) );
  NAND U21995 ( .A(n21145), .B(n21144), .Z(n21312) );
  NANDN U21996 ( .A(n21147), .B(n21146), .Z(n21151) );
  NAND U21997 ( .A(n21149), .B(n21148), .Z(n21150) );
  NAND U21998 ( .A(n21151), .B(n21150), .Z(n21310) );
  OR U21999 ( .A(n21153), .B(n21152), .Z(n21157) );
  NANDN U22000 ( .A(n21155), .B(n21154), .Z(n21156) );
  NAND U22001 ( .A(n21157), .B(n21156), .Z(n21309) );
  XNOR U22002 ( .A(n21312), .B(n21311), .Z(n21368) );
  XOR U22003 ( .A(n21367), .B(n21368), .Z(n21370) );
  NANDN U22004 ( .A(n21159), .B(n21158), .Z(n21163) );
  OR U22005 ( .A(n21161), .B(n21160), .Z(n21162) );
  NAND U22006 ( .A(n21163), .B(n21162), .Z(n21369) );
  XOR U22007 ( .A(n21370), .B(n21369), .Z(n21387) );
  OR U22008 ( .A(n21165), .B(n21164), .Z(n21169) );
  NAND U22009 ( .A(n21167), .B(n21166), .Z(n21168) );
  NAND U22010 ( .A(n21169), .B(n21168), .Z(n21386) );
  NANDN U22011 ( .A(n21171), .B(n21170), .Z(n21175) );
  NANDN U22012 ( .A(n21173), .B(n21172), .Z(n21174) );
  NAND U22013 ( .A(n21175), .B(n21174), .Z(n21375) );
  NANDN U22014 ( .A(n21181), .B(n21180), .Z(n21185) );
  NAND U22015 ( .A(n21183), .B(n21182), .Z(n21184) );
  NAND U22016 ( .A(n21185), .B(n21184), .Z(n21315) );
  NANDN U22017 ( .A(n21187), .B(n21186), .Z(n21191) );
  NAND U22018 ( .A(n21189), .B(n21188), .Z(n21190) );
  AND U22019 ( .A(n21191), .B(n21190), .Z(n21316) );
  XNOR U22020 ( .A(n21315), .B(n21316), .Z(n21317) );
  XNOR U22021 ( .A(b[9]), .B(a[146]), .Z(n21337) );
  NANDN U22022 ( .A(n21337), .B(n36925), .Z(n21194) );
  NAND U22023 ( .A(n36926), .B(n21192), .Z(n21193) );
  NAND U22024 ( .A(n21194), .B(n21193), .Z(n21301) );
  XNOR U22025 ( .A(n1054), .B(a[140]), .Z(n21340) );
  NANDN U22026 ( .A(n37665), .B(n21340), .Z(n21197) );
  NANDN U22027 ( .A(n21195), .B(n37604), .Z(n21196) );
  NAND U22028 ( .A(n21197), .B(n21196), .Z(n21299) );
  XNOR U22029 ( .A(b[21]), .B(a[134]), .Z(n21343) );
  NANDN U22030 ( .A(n21343), .B(n38101), .Z(n21200) );
  NAND U22031 ( .A(n38102), .B(n21198), .Z(n21199) );
  NAND U22032 ( .A(n21200), .B(n21199), .Z(n21300) );
  XNOR U22033 ( .A(n21299), .B(n21300), .Z(n21302) );
  XOR U22034 ( .A(n21301), .B(n21302), .Z(n21290) );
  XNOR U22035 ( .A(b[11]), .B(a[144]), .Z(n21346) );
  OR U22036 ( .A(n21346), .B(n37311), .Z(n21203) );
  NANDN U22037 ( .A(n21201), .B(n37218), .Z(n21202) );
  NAND U22038 ( .A(n21203), .B(n21202), .Z(n21288) );
  XOR U22039 ( .A(n1053), .B(a[142]), .Z(n21349) );
  NANDN U22040 ( .A(n21349), .B(n37424), .Z(n21206) );
  NANDN U22041 ( .A(n21204), .B(n37425), .Z(n21205) );
  AND U22042 ( .A(n21206), .B(n21205), .Z(n21287) );
  XNOR U22043 ( .A(n21288), .B(n21287), .Z(n21289) );
  XNOR U22044 ( .A(n21290), .B(n21289), .Z(n21306) );
  NANDN U22045 ( .A(n1049), .B(a[154]), .Z(n21207) );
  XNOR U22046 ( .A(b[1]), .B(n21207), .Z(n21209) );
  NANDN U22047 ( .A(b[0]), .B(a[153]), .Z(n21208) );
  AND U22048 ( .A(n21209), .B(n21208), .Z(n21265) );
  NAND U22049 ( .A(n38490), .B(n21210), .Z(n21212) );
  XNOR U22050 ( .A(n1058), .B(a[126]), .Z(n21355) );
  NANDN U22051 ( .A(n1048), .B(n21355), .Z(n21211) );
  NAND U22052 ( .A(n21212), .B(n21211), .Z(n21263) );
  NANDN U22053 ( .A(n1059), .B(a[122]), .Z(n21264) );
  XNOR U22054 ( .A(n21263), .B(n21264), .Z(n21266) );
  XNOR U22055 ( .A(n21265), .B(n21266), .Z(n21304) );
  NANDN U22056 ( .A(n21213), .B(n38205), .Z(n21215) );
  XNOR U22057 ( .A(b[23]), .B(a[132]), .Z(n21358) );
  OR U22058 ( .A(n21358), .B(n38268), .Z(n21214) );
  NAND U22059 ( .A(n21215), .B(n21214), .Z(n21328) );
  XOR U22060 ( .A(b[7]), .B(a[148]), .Z(n21361) );
  NAND U22061 ( .A(n21361), .B(n36701), .Z(n21218) );
  NAND U22062 ( .A(n21216), .B(n36702), .Z(n21217) );
  NAND U22063 ( .A(n21218), .B(n21217), .Z(n21325) );
  XOR U22064 ( .A(b[25]), .B(a[130]), .Z(n21364) );
  NAND U22065 ( .A(n21364), .B(n38325), .Z(n21221) );
  NANDN U22066 ( .A(n21219), .B(n38326), .Z(n21220) );
  AND U22067 ( .A(n21221), .B(n21220), .Z(n21326) );
  XNOR U22068 ( .A(n21325), .B(n21326), .Z(n21327) );
  XOR U22069 ( .A(n21328), .B(n21327), .Z(n21303) );
  XOR U22070 ( .A(n21306), .B(n21305), .Z(n21318) );
  XOR U22071 ( .A(n21317), .B(n21318), .Z(n21373) );
  XNOR U22072 ( .A(n21374), .B(n21373), .Z(n21376) );
  XNOR U22073 ( .A(n21375), .B(n21376), .Z(n21385) );
  XOR U22074 ( .A(n21386), .B(n21385), .Z(n21388) );
  NANDN U22075 ( .A(n21223), .B(n21222), .Z(n21227) );
  OR U22076 ( .A(n21225), .B(n21224), .Z(n21226) );
  NAND U22077 ( .A(n21227), .B(n21226), .Z(n21379) );
  NAND U22078 ( .A(n21229), .B(n21228), .Z(n21233) );
  NANDN U22079 ( .A(n21231), .B(n21230), .Z(n21232) );
  NAND U22080 ( .A(n21233), .B(n21232), .Z(n21380) );
  XNOR U22081 ( .A(n21379), .B(n21380), .Z(n21381) );
  XOR U22082 ( .A(n21382), .B(n21381), .Z(n21259) );
  NANDN U22083 ( .A(n21235), .B(n21234), .Z(n21239) );
  NAND U22084 ( .A(n21237), .B(n21236), .Z(n21238) );
  NAND U22085 ( .A(n21239), .B(n21238), .Z(n21257) );
  NANDN U22086 ( .A(n21241), .B(n21240), .Z(n21245) );
  OR U22087 ( .A(n21243), .B(n21242), .Z(n21244) );
  NAND U22088 ( .A(n21245), .B(n21244), .Z(n21258) );
  XNOR U22089 ( .A(n21257), .B(n21258), .Z(n21260) );
  XOR U22090 ( .A(n21259), .B(n21260), .Z(n21251) );
  XOR U22091 ( .A(n21252), .B(n21251), .Z(n21253) );
  XNOR U22092 ( .A(n21254), .B(n21253), .Z(n21391) );
  XNOR U22093 ( .A(n21391), .B(sreg[378]), .Z(n21393) );
  NAND U22094 ( .A(n21246), .B(sreg[377]), .Z(n21250) );
  OR U22095 ( .A(n21248), .B(n21247), .Z(n21249) );
  AND U22096 ( .A(n21250), .B(n21249), .Z(n21392) );
  XOR U22097 ( .A(n21393), .B(n21392), .Z(c[378]) );
  NAND U22098 ( .A(n21252), .B(n21251), .Z(n21256) );
  NAND U22099 ( .A(n21254), .B(n21253), .Z(n21255) );
  NAND U22100 ( .A(n21256), .B(n21255), .Z(n21399) );
  NANDN U22101 ( .A(n21258), .B(n21257), .Z(n21262) );
  NAND U22102 ( .A(n21260), .B(n21259), .Z(n21261) );
  NAND U22103 ( .A(n21262), .B(n21261), .Z(n21397) );
  NANDN U22104 ( .A(n21264), .B(n21263), .Z(n21268) );
  NAND U22105 ( .A(n21266), .B(n21265), .Z(n21267) );
  NAND U22106 ( .A(n21268), .B(n21267), .Z(n21479) );
  XOR U22107 ( .A(b[19]), .B(n23393), .Z(n21424) );
  NANDN U22108 ( .A(n21424), .B(n37934), .Z(n21271) );
  NANDN U22109 ( .A(n21269), .B(n37935), .Z(n21270) );
  NAND U22110 ( .A(n21271), .B(n21270), .Z(n21489) );
  XNOR U22111 ( .A(b[27]), .B(a[129]), .Z(n21427) );
  NANDN U22112 ( .A(n21427), .B(n38423), .Z(n21274) );
  NAND U22113 ( .A(n21272), .B(n38424), .Z(n21273) );
  NAND U22114 ( .A(n21274), .B(n21273), .Z(n21486) );
  XOR U22115 ( .A(b[5]), .B(n25435), .Z(n21430) );
  NANDN U22116 ( .A(n21430), .B(n36587), .Z(n21277) );
  NANDN U22117 ( .A(n21275), .B(n36588), .Z(n21276) );
  AND U22118 ( .A(n21277), .B(n21276), .Z(n21487) );
  XNOR U22119 ( .A(n21486), .B(n21487), .Z(n21488) );
  XNOR U22120 ( .A(n21489), .B(n21488), .Z(n21477) );
  NAND U22121 ( .A(n21278), .B(n37762), .Z(n21280) );
  XNOR U22122 ( .A(b[17]), .B(a[139]), .Z(n21433) );
  NANDN U22123 ( .A(n21433), .B(n37764), .Z(n21279) );
  NAND U22124 ( .A(n21280), .B(n21279), .Z(n21451) );
  XNOR U22125 ( .A(b[31]), .B(a[125]), .Z(n21436) );
  NANDN U22126 ( .A(n21436), .B(n38552), .Z(n21283) );
  NANDN U22127 ( .A(n21281), .B(n38553), .Z(n21282) );
  NAND U22128 ( .A(n21283), .B(n21282), .Z(n21448) );
  OR U22129 ( .A(n21284), .B(n36105), .Z(n21286) );
  XNOR U22130 ( .A(b[3]), .B(a[153]), .Z(n21439) );
  NANDN U22131 ( .A(n21439), .B(n36107), .Z(n21285) );
  AND U22132 ( .A(n21286), .B(n21285), .Z(n21449) );
  XNOR U22133 ( .A(n21448), .B(n21449), .Z(n21450) );
  XOR U22134 ( .A(n21451), .B(n21450), .Z(n21476) );
  XNOR U22135 ( .A(n21477), .B(n21476), .Z(n21478) );
  XNOR U22136 ( .A(n21479), .B(n21478), .Z(n21415) );
  NANDN U22137 ( .A(n21288), .B(n21287), .Z(n21292) );
  NAND U22138 ( .A(n21290), .B(n21289), .Z(n21291) );
  NAND U22139 ( .A(n21292), .B(n21291), .Z(n21468) );
  NANDN U22140 ( .A(n21294), .B(n21293), .Z(n21298) );
  NAND U22141 ( .A(n21296), .B(n21295), .Z(n21297) );
  NAND U22142 ( .A(n21298), .B(n21297), .Z(n21467) );
  XNOR U22143 ( .A(n21467), .B(n21466), .Z(n21469) );
  XOR U22144 ( .A(n21468), .B(n21469), .Z(n21414) );
  XOR U22145 ( .A(n21415), .B(n21414), .Z(n21416) );
  NANDN U22146 ( .A(n21304), .B(n21303), .Z(n21308) );
  NAND U22147 ( .A(n21306), .B(n21305), .Z(n21307) );
  NAND U22148 ( .A(n21308), .B(n21307), .Z(n21417) );
  XNOR U22149 ( .A(n21416), .B(n21417), .Z(n21530) );
  OR U22150 ( .A(n21310), .B(n21309), .Z(n21314) );
  NAND U22151 ( .A(n21312), .B(n21311), .Z(n21313) );
  NAND U22152 ( .A(n21314), .B(n21313), .Z(n21529) );
  NANDN U22153 ( .A(n21316), .B(n21315), .Z(n21320) );
  NAND U22154 ( .A(n21318), .B(n21317), .Z(n21319) );
  NAND U22155 ( .A(n21320), .B(n21319), .Z(n21410) );
  NANDN U22156 ( .A(n21326), .B(n21325), .Z(n21330) );
  NAND U22157 ( .A(n21328), .B(n21327), .Z(n21329) );
  NAND U22158 ( .A(n21330), .B(n21329), .Z(n21470) );
  NANDN U22159 ( .A(n21332), .B(n21331), .Z(n21336) );
  NAND U22160 ( .A(n21334), .B(n21333), .Z(n21335) );
  AND U22161 ( .A(n21336), .B(n21335), .Z(n21471) );
  XNOR U22162 ( .A(n21470), .B(n21471), .Z(n21472) );
  XNOR U22163 ( .A(b[9]), .B(a[147]), .Z(n21492) );
  NANDN U22164 ( .A(n21492), .B(n36925), .Z(n21339) );
  NANDN U22165 ( .A(n21337), .B(n36926), .Z(n21338) );
  NAND U22166 ( .A(n21339), .B(n21338), .Z(n21456) );
  XOR U22167 ( .A(b[15]), .B(n23961), .Z(n21495) );
  OR U22168 ( .A(n21495), .B(n37665), .Z(n21342) );
  NAND U22169 ( .A(n21340), .B(n37604), .Z(n21341) );
  AND U22170 ( .A(n21342), .B(n21341), .Z(n21454) );
  XNOR U22171 ( .A(b[21]), .B(a[135]), .Z(n21498) );
  NANDN U22172 ( .A(n21498), .B(n38101), .Z(n21345) );
  NANDN U22173 ( .A(n21343), .B(n38102), .Z(n21344) );
  AND U22174 ( .A(n21345), .B(n21344), .Z(n21455) );
  XOR U22175 ( .A(n21456), .B(n21457), .Z(n21445) );
  XOR U22176 ( .A(b[11]), .B(n24554), .Z(n21501) );
  OR U22177 ( .A(n21501), .B(n37311), .Z(n21348) );
  NANDN U22178 ( .A(n21346), .B(n37218), .Z(n21347) );
  NAND U22179 ( .A(n21348), .B(n21347), .Z(n21443) );
  XOR U22180 ( .A(n1053), .B(a[143]), .Z(n21504) );
  NANDN U22181 ( .A(n21504), .B(n37424), .Z(n21351) );
  NANDN U22182 ( .A(n21349), .B(n37425), .Z(n21350) );
  AND U22183 ( .A(n21351), .B(n21350), .Z(n21442) );
  XNOR U22184 ( .A(n21443), .B(n21442), .Z(n21444) );
  XOR U22185 ( .A(n21445), .B(n21444), .Z(n21462) );
  NANDN U22186 ( .A(n1049), .B(a[155]), .Z(n21352) );
  XNOR U22187 ( .A(b[1]), .B(n21352), .Z(n21354) );
  IV U22188 ( .A(a[154]), .Z(n25862) );
  NANDN U22189 ( .A(n25862), .B(n1049), .Z(n21353) );
  AND U22190 ( .A(n21354), .B(n21353), .Z(n21420) );
  NAND U22191 ( .A(n38490), .B(n21355), .Z(n21357) );
  XNOR U22192 ( .A(n1058), .B(a[127]), .Z(n21507) );
  NANDN U22193 ( .A(n1048), .B(n21507), .Z(n21356) );
  NAND U22194 ( .A(n21357), .B(n21356), .Z(n21418) );
  NANDN U22195 ( .A(n1059), .B(a[123]), .Z(n21419) );
  XNOR U22196 ( .A(n21418), .B(n21419), .Z(n21421) );
  XOR U22197 ( .A(n21420), .B(n21421), .Z(n21460) );
  NANDN U22198 ( .A(n21358), .B(n38205), .Z(n21360) );
  XNOR U22199 ( .A(b[23]), .B(a[133]), .Z(n21513) );
  OR U22200 ( .A(n21513), .B(n38268), .Z(n21359) );
  NAND U22201 ( .A(n21360), .B(n21359), .Z(n21483) );
  XOR U22202 ( .A(b[7]), .B(a[149]), .Z(n21516) );
  NAND U22203 ( .A(n21516), .B(n36701), .Z(n21363) );
  NAND U22204 ( .A(n21361), .B(n36702), .Z(n21362) );
  NAND U22205 ( .A(n21363), .B(n21362), .Z(n21480) );
  XNOR U22206 ( .A(b[25]), .B(a[131]), .Z(n21519) );
  NANDN U22207 ( .A(n21519), .B(n38325), .Z(n21366) );
  NAND U22208 ( .A(n21364), .B(n38326), .Z(n21365) );
  AND U22209 ( .A(n21366), .B(n21365), .Z(n21481) );
  XNOR U22210 ( .A(n21480), .B(n21481), .Z(n21482) );
  XNOR U22211 ( .A(n21483), .B(n21482), .Z(n21461) );
  XOR U22212 ( .A(n21460), .B(n21461), .Z(n21463) );
  XNOR U22213 ( .A(n21462), .B(n21463), .Z(n21473) );
  XNOR U22214 ( .A(n21472), .B(n21473), .Z(n21408) );
  XNOR U22215 ( .A(n21409), .B(n21408), .Z(n21411) );
  XNOR U22216 ( .A(n21410), .B(n21411), .Z(n21528) );
  XOR U22217 ( .A(n21529), .B(n21528), .Z(n21531) );
  NANDN U22218 ( .A(n21368), .B(n21367), .Z(n21372) );
  OR U22219 ( .A(n21370), .B(n21369), .Z(n21371) );
  NAND U22220 ( .A(n21372), .B(n21371), .Z(n21522) );
  NAND U22221 ( .A(n21374), .B(n21373), .Z(n21378) );
  NANDN U22222 ( .A(n21376), .B(n21375), .Z(n21377) );
  NAND U22223 ( .A(n21378), .B(n21377), .Z(n21523) );
  XNOR U22224 ( .A(n21522), .B(n21523), .Z(n21524) );
  XOR U22225 ( .A(n21525), .B(n21524), .Z(n21404) );
  NANDN U22226 ( .A(n21380), .B(n21379), .Z(n21384) );
  NAND U22227 ( .A(n21382), .B(n21381), .Z(n21383) );
  NAND U22228 ( .A(n21384), .B(n21383), .Z(n21402) );
  NANDN U22229 ( .A(n21386), .B(n21385), .Z(n21390) );
  OR U22230 ( .A(n21388), .B(n21387), .Z(n21389) );
  NAND U22231 ( .A(n21390), .B(n21389), .Z(n21403) );
  XNOR U22232 ( .A(n21402), .B(n21403), .Z(n21405) );
  XOR U22233 ( .A(n21404), .B(n21405), .Z(n21396) );
  XOR U22234 ( .A(n21397), .B(n21396), .Z(n21398) );
  XNOR U22235 ( .A(n21399), .B(n21398), .Z(n21534) );
  XNOR U22236 ( .A(n21534), .B(sreg[379]), .Z(n21536) );
  NAND U22237 ( .A(n21391), .B(sreg[378]), .Z(n21395) );
  OR U22238 ( .A(n21393), .B(n21392), .Z(n21394) );
  AND U22239 ( .A(n21395), .B(n21394), .Z(n21535) );
  XOR U22240 ( .A(n21536), .B(n21535), .Z(c[379]) );
  NAND U22241 ( .A(n21397), .B(n21396), .Z(n21401) );
  NAND U22242 ( .A(n21399), .B(n21398), .Z(n21400) );
  NAND U22243 ( .A(n21401), .B(n21400), .Z(n21542) );
  NANDN U22244 ( .A(n21403), .B(n21402), .Z(n21407) );
  NAND U22245 ( .A(n21405), .B(n21404), .Z(n21406) );
  NAND U22246 ( .A(n21407), .B(n21406), .Z(n21539) );
  NAND U22247 ( .A(n21409), .B(n21408), .Z(n21413) );
  NANDN U22248 ( .A(n21411), .B(n21410), .Z(n21412) );
  NAND U22249 ( .A(n21413), .B(n21412), .Z(n21551) );
  XNOR U22250 ( .A(n21551), .B(n21552), .Z(n21553) );
  NANDN U22251 ( .A(n21419), .B(n21418), .Z(n21423) );
  NAND U22252 ( .A(n21421), .B(n21420), .Z(n21422) );
  NAND U22253 ( .A(n21423), .B(n21422), .Z(n21626) );
  XNOR U22254 ( .A(b[19]), .B(a[138]), .Z(n21569) );
  NANDN U22255 ( .A(n21569), .B(n37934), .Z(n21426) );
  NANDN U22256 ( .A(n21424), .B(n37935), .Z(n21425) );
  NAND U22257 ( .A(n21426), .B(n21425), .Z(n21636) );
  XOR U22258 ( .A(b[27]), .B(a[130]), .Z(n21572) );
  NAND U22259 ( .A(n38423), .B(n21572), .Z(n21429) );
  NANDN U22260 ( .A(n21427), .B(n38424), .Z(n21428) );
  NAND U22261 ( .A(n21429), .B(n21428), .Z(n21633) );
  XOR U22262 ( .A(b[5]), .B(n25213), .Z(n21575) );
  NANDN U22263 ( .A(n21575), .B(n36587), .Z(n21432) );
  NANDN U22264 ( .A(n21430), .B(n36588), .Z(n21431) );
  AND U22265 ( .A(n21432), .B(n21431), .Z(n21634) );
  XNOR U22266 ( .A(n21633), .B(n21634), .Z(n21635) );
  XNOR U22267 ( .A(n21636), .B(n21635), .Z(n21624) );
  NANDN U22268 ( .A(n21433), .B(n37762), .Z(n21435) );
  XOR U22269 ( .A(b[17]), .B(a[140]), .Z(n21578) );
  NAND U22270 ( .A(n21578), .B(n37764), .Z(n21434) );
  NAND U22271 ( .A(n21435), .B(n21434), .Z(n21596) );
  XNOR U22272 ( .A(b[31]), .B(a[126]), .Z(n21581) );
  NANDN U22273 ( .A(n21581), .B(n38552), .Z(n21438) );
  NANDN U22274 ( .A(n21436), .B(n38553), .Z(n21437) );
  NAND U22275 ( .A(n21438), .B(n21437), .Z(n21593) );
  OR U22276 ( .A(n21439), .B(n36105), .Z(n21441) );
  XOR U22277 ( .A(b[3]), .B(n25862), .Z(n21584) );
  NANDN U22278 ( .A(n21584), .B(n36107), .Z(n21440) );
  AND U22279 ( .A(n21441), .B(n21440), .Z(n21594) );
  XNOR U22280 ( .A(n21593), .B(n21594), .Z(n21595) );
  XOR U22281 ( .A(n21596), .B(n21595), .Z(n21623) );
  XNOR U22282 ( .A(n21624), .B(n21623), .Z(n21625) );
  XNOR U22283 ( .A(n21626), .B(n21625), .Z(n21669) );
  NANDN U22284 ( .A(n21443), .B(n21442), .Z(n21447) );
  NAND U22285 ( .A(n21445), .B(n21444), .Z(n21446) );
  NAND U22286 ( .A(n21447), .B(n21446), .Z(n21614) );
  NANDN U22287 ( .A(n21449), .B(n21448), .Z(n21453) );
  NAND U22288 ( .A(n21451), .B(n21450), .Z(n21452) );
  NAND U22289 ( .A(n21453), .B(n21452), .Z(n21612) );
  OR U22290 ( .A(n21455), .B(n21454), .Z(n21459) );
  NANDN U22291 ( .A(n21457), .B(n21456), .Z(n21458) );
  NAND U22292 ( .A(n21459), .B(n21458), .Z(n21611) );
  XNOR U22293 ( .A(n21614), .B(n21613), .Z(n21670) );
  XNOR U22294 ( .A(n21669), .B(n21670), .Z(n21671) );
  NANDN U22295 ( .A(n21461), .B(n21460), .Z(n21465) );
  OR U22296 ( .A(n21463), .B(n21462), .Z(n21464) );
  AND U22297 ( .A(n21465), .B(n21464), .Z(n21672) );
  XOR U22298 ( .A(n21671), .B(n21672), .Z(n21559) );
  NANDN U22299 ( .A(n21471), .B(n21470), .Z(n21475) );
  NANDN U22300 ( .A(n21473), .B(n21472), .Z(n21474) );
  NAND U22301 ( .A(n21475), .B(n21474), .Z(n21678) );
  NANDN U22302 ( .A(n21481), .B(n21480), .Z(n21485) );
  NAND U22303 ( .A(n21483), .B(n21482), .Z(n21484) );
  NAND U22304 ( .A(n21485), .B(n21484), .Z(n21617) );
  NANDN U22305 ( .A(n21487), .B(n21486), .Z(n21491) );
  NAND U22306 ( .A(n21489), .B(n21488), .Z(n21490) );
  AND U22307 ( .A(n21491), .B(n21490), .Z(n21618) );
  XNOR U22308 ( .A(n21617), .B(n21618), .Z(n21619) );
  XNOR U22309 ( .A(n1052), .B(a[148]), .Z(n21639) );
  NAND U22310 ( .A(n36925), .B(n21639), .Z(n21494) );
  NANDN U22311 ( .A(n21492), .B(n36926), .Z(n21493) );
  NAND U22312 ( .A(n21494), .B(n21493), .Z(n21601) );
  XOR U22313 ( .A(b[15]), .B(n24120), .Z(n21642) );
  OR U22314 ( .A(n21642), .B(n37665), .Z(n21497) );
  NANDN U22315 ( .A(n21495), .B(n37604), .Z(n21496) );
  AND U22316 ( .A(n21497), .B(n21496), .Z(n21599) );
  XNOR U22317 ( .A(n1056), .B(a[136]), .Z(n21645) );
  NAND U22318 ( .A(n21645), .B(n38101), .Z(n21500) );
  NANDN U22319 ( .A(n21498), .B(n38102), .Z(n21499) );
  AND U22320 ( .A(n21500), .B(n21499), .Z(n21600) );
  XOR U22321 ( .A(n21601), .B(n21602), .Z(n21590) );
  XNOR U22322 ( .A(b[11]), .B(a[146]), .Z(n21648) );
  OR U22323 ( .A(n21648), .B(n37311), .Z(n21503) );
  NANDN U22324 ( .A(n21501), .B(n37218), .Z(n21502) );
  NAND U22325 ( .A(n21503), .B(n21502), .Z(n21588) );
  XOR U22326 ( .A(n1053), .B(a[144]), .Z(n21651) );
  NANDN U22327 ( .A(n21651), .B(n37424), .Z(n21506) );
  NANDN U22328 ( .A(n21504), .B(n37425), .Z(n21505) );
  AND U22329 ( .A(n21506), .B(n21505), .Z(n21587) );
  XNOR U22330 ( .A(n21588), .B(n21587), .Z(n21589) );
  XOR U22331 ( .A(n21590), .B(n21589), .Z(n21607) );
  NAND U22332 ( .A(n38490), .B(n21507), .Z(n21509) );
  XNOR U22333 ( .A(n1058), .B(a[128]), .Z(n21657) );
  NANDN U22334 ( .A(n1048), .B(n21657), .Z(n21508) );
  NAND U22335 ( .A(n21509), .B(n21508), .Z(n21563) );
  NANDN U22336 ( .A(n1059), .B(a[124]), .Z(n21564) );
  XNOR U22337 ( .A(n21563), .B(n21564), .Z(n21566) );
  NANDN U22338 ( .A(n1049), .B(a[156]), .Z(n21510) );
  XNOR U22339 ( .A(b[1]), .B(n21510), .Z(n21512) );
  NANDN U22340 ( .A(b[0]), .B(a[155]), .Z(n21511) );
  AND U22341 ( .A(n21512), .B(n21511), .Z(n21565) );
  XOR U22342 ( .A(n21566), .B(n21565), .Z(n21605) );
  NANDN U22343 ( .A(n21513), .B(n38205), .Z(n21515) );
  XNOR U22344 ( .A(b[23]), .B(a[134]), .Z(n21660) );
  OR U22345 ( .A(n21660), .B(n38268), .Z(n21514) );
  NAND U22346 ( .A(n21515), .B(n21514), .Z(n21630) );
  XOR U22347 ( .A(b[7]), .B(a[150]), .Z(n21663) );
  NAND U22348 ( .A(n21663), .B(n36701), .Z(n21518) );
  NAND U22349 ( .A(n21516), .B(n36702), .Z(n21517) );
  NAND U22350 ( .A(n21518), .B(n21517), .Z(n21627) );
  XOR U22351 ( .A(b[25]), .B(a[132]), .Z(n21666) );
  NAND U22352 ( .A(n21666), .B(n38325), .Z(n21521) );
  NANDN U22353 ( .A(n21519), .B(n38326), .Z(n21520) );
  AND U22354 ( .A(n21521), .B(n21520), .Z(n21628) );
  XNOR U22355 ( .A(n21627), .B(n21628), .Z(n21629) );
  XNOR U22356 ( .A(n21630), .B(n21629), .Z(n21606) );
  XOR U22357 ( .A(n21605), .B(n21606), .Z(n21608) );
  XNOR U22358 ( .A(n21607), .B(n21608), .Z(n21620) );
  XOR U22359 ( .A(n21619), .B(n21620), .Z(n21676) );
  XNOR U22360 ( .A(n21675), .B(n21676), .Z(n21677) );
  XNOR U22361 ( .A(n21678), .B(n21677), .Z(n21557) );
  XNOR U22362 ( .A(n21558), .B(n21557), .Z(n21560) );
  XNOR U22363 ( .A(n21559), .B(n21560), .Z(n21554) );
  XOR U22364 ( .A(n21553), .B(n21554), .Z(n21548) );
  NANDN U22365 ( .A(n21523), .B(n21522), .Z(n21527) );
  NAND U22366 ( .A(n21525), .B(n21524), .Z(n21526) );
  NAND U22367 ( .A(n21527), .B(n21526), .Z(n21545) );
  NANDN U22368 ( .A(n21529), .B(n21528), .Z(n21533) );
  OR U22369 ( .A(n21531), .B(n21530), .Z(n21532) );
  NAND U22370 ( .A(n21533), .B(n21532), .Z(n21546) );
  XNOR U22371 ( .A(n21545), .B(n21546), .Z(n21547) );
  XNOR U22372 ( .A(n21548), .B(n21547), .Z(n21540) );
  XNOR U22373 ( .A(n21539), .B(n21540), .Z(n21541) );
  XNOR U22374 ( .A(n21542), .B(n21541), .Z(n21681) );
  XNOR U22375 ( .A(n21681), .B(sreg[380]), .Z(n21683) );
  NAND U22376 ( .A(n21534), .B(sreg[379]), .Z(n21538) );
  OR U22377 ( .A(n21536), .B(n21535), .Z(n21537) );
  AND U22378 ( .A(n21538), .B(n21537), .Z(n21682) );
  XOR U22379 ( .A(n21683), .B(n21682), .Z(c[380]) );
  NANDN U22380 ( .A(n21540), .B(n21539), .Z(n21544) );
  NAND U22381 ( .A(n21542), .B(n21541), .Z(n21543) );
  NAND U22382 ( .A(n21544), .B(n21543), .Z(n21689) );
  NANDN U22383 ( .A(n21546), .B(n21545), .Z(n21550) );
  NAND U22384 ( .A(n21548), .B(n21547), .Z(n21549) );
  NAND U22385 ( .A(n21550), .B(n21549), .Z(n21687) );
  NANDN U22386 ( .A(n21552), .B(n21551), .Z(n21556) );
  NANDN U22387 ( .A(n21554), .B(n21553), .Z(n21555) );
  NAND U22388 ( .A(n21556), .B(n21555), .Z(n21693) );
  OR U22389 ( .A(n21558), .B(n21557), .Z(n21562) );
  OR U22390 ( .A(n21560), .B(n21559), .Z(n21561) );
  AND U22391 ( .A(n21562), .B(n21561), .Z(n21692) );
  XNOR U22392 ( .A(n21693), .B(n21692), .Z(n21694) );
  NANDN U22393 ( .A(n21564), .B(n21563), .Z(n21568) );
  NAND U22394 ( .A(n21566), .B(n21565), .Z(n21567) );
  NAND U22395 ( .A(n21568), .B(n21567), .Z(n21759) );
  XOR U22396 ( .A(b[19]), .B(n23668), .Z(n21704) );
  NANDN U22397 ( .A(n21704), .B(n37934), .Z(n21571) );
  NANDN U22398 ( .A(n21569), .B(n37935), .Z(n21570) );
  NAND U22399 ( .A(n21571), .B(n21570), .Z(n21769) );
  XNOR U22400 ( .A(b[27]), .B(a[131]), .Z(n21707) );
  NANDN U22401 ( .A(n21707), .B(n38423), .Z(n21574) );
  NAND U22402 ( .A(n21572), .B(n38424), .Z(n21573) );
  NAND U22403 ( .A(n21574), .B(n21573), .Z(n21766) );
  XNOR U22404 ( .A(b[5]), .B(a[153]), .Z(n21710) );
  NANDN U22405 ( .A(n21710), .B(n36587), .Z(n21577) );
  NANDN U22406 ( .A(n21575), .B(n36588), .Z(n21576) );
  AND U22407 ( .A(n21577), .B(n21576), .Z(n21767) );
  XNOR U22408 ( .A(n21766), .B(n21767), .Z(n21768) );
  XNOR U22409 ( .A(n21769), .B(n21768), .Z(n21757) );
  NAND U22410 ( .A(n21578), .B(n37762), .Z(n21580) );
  XNOR U22411 ( .A(b[17]), .B(a[141]), .Z(n21713) );
  NANDN U22412 ( .A(n21713), .B(n37764), .Z(n21579) );
  NAND U22413 ( .A(n21580), .B(n21579), .Z(n21731) );
  XNOR U22414 ( .A(b[31]), .B(a[127]), .Z(n21716) );
  NANDN U22415 ( .A(n21716), .B(n38552), .Z(n21583) );
  NANDN U22416 ( .A(n21581), .B(n38553), .Z(n21582) );
  NAND U22417 ( .A(n21583), .B(n21582), .Z(n21728) );
  OR U22418 ( .A(n21584), .B(n36105), .Z(n21586) );
  XNOR U22419 ( .A(b[3]), .B(a[155]), .Z(n21719) );
  NANDN U22420 ( .A(n21719), .B(n36107), .Z(n21585) );
  AND U22421 ( .A(n21586), .B(n21585), .Z(n21729) );
  XNOR U22422 ( .A(n21728), .B(n21729), .Z(n21730) );
  XOR U22423 ( .A(n21731), .B(n21730), .Z(n21756) );
  XNOR U22424 ( .A(n21757), .B(n21756), .Z(n21758) );
  XNOR U22425 ( .A(n21759), .B(n21758), .Z(n21802) );
  NANDN U22426 ( .A(n21588), .B(n21587), .Z(n21592) );
  NAND U22427 ( .A(n21590), .B(n21589), .Z(n21591) );
  NAND U22428 ( .A(n21592), .B(n21591), .Z(n21747) );
  NANDN U22429 ( .A(n21594), .B(n21593), .Z(n21598) );
  NAND U22430 ( .A(n21596), .B(n21595), .Z(n21597) );
  NAND U22431 ( .A(n21598), .B(n21597), .Z(n21745) );
  OR U22432 ( .A(n21600), .B(n21599), .Z(n21604) );
  NANDN U22433 ( .A(n21602), .B(n21601), .Z(n21603) );
  NAND U22434 ( .A(n21604), .B(n21603), .Z(n21744) );
  XNOR U22435 ( .A(n21747), .B(n21746), .Z(n21803) );
  XOR U22436 ( .A(n21802), .B(n21803), .Z(n21805) );
  NANDN U22437 ( .A(n21606), .B(n21605), .Z(n21610) );
  OR U22438 ( .A(n21608), .B(n21607), .Z(n21609) );
  NAND U22439 ( .A(n21610), .B(n21609), .Z(n21804) );
  XOR U22440 ( .A(n21805), .B(n21804), .Z(n21822) );
  OR U22441 ( .A(n21612), .B(n21611), .Z(n21616) );
  NAND U22442 ( .A(n21614), .B(n21613), .Z(n21615) );
  NAND U22443 ( .A(n21616), .B(n21615), .Z(n21821) );
  NANDN U22444 ( .A(n21618), .B(n21617), .Z(n21622) );
  NANDN U22445 ( .A(n21620), .B(n21619), .Z(n21621) );
  NAND U22446 ( .A(n21622), .B(n21621), .Z(n21810) );
  NANDN U22447 ( .A(n21628), .B(n21627), .Z(n21632) );
  NAND U22448 ( .A(n21630), .B(n21629), .Z(n21631) );
  NAND U22449 ( .A(n21632), .B(n21631), .Z(n21750) );
  NANDN U22450 ( .A(n21634), .B(n21633), .Z(n21638) );
  NAND U22451 ( .A(n21636), .B(n21635), .Z(n21637) );
  AND U22452 ( .A(n21638), .B(n21637), .Z(n21751) );
  XNOR U22453 ( .A(n21750), .B(n21751), .Z(n21752) );
  XOR U22454 ( .A(n1052), .B(a[149]), .Z(n21778) );
  NANDN U22455 ( .A(n21778), .B(n36925), .Z(n21641) );
  NAND U22456 ( .A(n36926), .B(n21639), .Z(n21640) );
  NAND U22457 ( .A(n21641), .B(n21640), .Z(n21736) );
  XNOR U22458 ( .A(n1054), .B(a[143]), .Z(n21775) );
  NANDN U22459 ( .A(n37665), .B(n21775), .Z(n21644) );
  NANDN U22460 ( .A(n21642), .B(n37604), .Z(n21643) );
  NAND U22461 ( .A(n21644), .B(n21643), .Z(n21734) );
  XOR U22462 ( .A(n1056), .B(a[137]), .Z(n21772) );
  NANDN U22463 ( .A(n21772), .B(n38101), .Z(n21647) );
  NAND U22464 ( .A(n38102), .B(n21645), .Z(n21646) );
  NAND U22465 ( .A(n21647), .B(n21646), .Z(n21735) );
  XNOR U22466 ( .A(n21734), .B(n21735), .Z(n21737) );
  XOR U22467 ( .A(n21736), .B(n21737), .Z(n21725) );
  XNOR U22468 ( .A(b[11]), .B(a[147]), .Z(n21781) );
  OR U22469 ( .A(n21781), .B(n37311), .Z(n21650) );
  NANDN U22470 ( .A(n21648), .B(n37218), .Z(n21649) );
  NAND U22471 ( .A(n21650), .B(n21649), .Z(n21723) );
  XOR U22472 ( .A(n1053), .B(a[145]), .Z(n21784) );
  NANDN U22473 ( .A(n21784), .B(n37424), .Z(n21653) );
  NANDN U22474 ( .A(n21651), .B(n37425), .Z(n21652) );
  AND U22475 ( .A(n21653), .B(n21652), .Z(n21722) );
  XNOR U22476 ( .A(n21723), .B(n21722), .Z(n21724) );
  XNOR U22477 ( .A(n21725), .B(n21724), .Z(n21741) );
  NANDN U22478 ( .A(n1049), .B(a[157]), .Z(n21654) );
  XNOR U22479 ( .A(b[1]), .B(n21654), .Z(n21656) );
  NANDN U22480 ( .A(b[0]), .B(a[156]), .Z(n21655) );
  AND U22481 ( .A(n21656), .B(n21655), .Z(n21700) );
  NAND U22482 ( .A(n38490), .B(n21657), .Z(n21659) );
  XOR U22483 ( .A(n1058), .B(n22221), .Z(n21790) );
  NANDN U22484 ( .A(n1048), .B(n21790), .Z(n21658) );
  NAND U22485 ( .A(n21659), .B(n21658), .Z(n21698) );
  NANDN U22486 ( .A(n1059), .B(a[125]), .Z(n21699) );
  XNOR U22487 ( .A(n21698), .B(n21699), .Z(n21701) );
  XNOR U22488 ( .A(n21700), .B(n21701), .Z(n21739) );
  NANDN U22489 ( .A(n21660), .B(n38205), .Z(n21662) );
  XNOR U22490 ( .A(b[23]), .B(a[135]), .Z(n21793) );
  OR U22491 ( .A(n21793), .B(n38268), .Z(n21661) );
  NAND U22492 ( .A(n21662), .B(n21661), .Z(n21763) );
  XNOR U22493 ( .A(b[7]), .B(a[151]), .Z(n21796) );
  NANDN U22494 ( .A(n21796), .B(n36701), .Z(n21665) );
  NAND U22495 ( .A(n21663), .B(n36702), .Z(n21664) );
  NAND U22496 ( .A(n21665), .B(n21664), .Z(n21760) );
  XOR U22497 ( .A(b[25]), .B(a[133]), .Z(n21799) );
  NAND U22498 ( .A(n21799), .B(n38325), .Z(n21668) );
  NAND U22499 ( .A(n21666), .B(n38326), .Z(n21667) );
  AND U22500 ( .A(n21668), .B(n21667), .Z(n21761) );
  XNOR U22501 ( .A(n21760), .B(n21761), .Z(n21762) );
  XOR U22502 ( .A(n21763), .B(n21762), .Z(n21738) );
  XOR U22503 ( .A(n21741), .B(n21740), .Z(n21753) );
  XOR U22504 ( .A(n21752), .B(n21753), .Z(n21808) );
  XNOR U22505 ( .A(n21809), .B(n21808), .Z(n21811) );
  XNOR U22506 ( .A(n21810), .B(n21811), .Z(n21820) );
  XOR U22507 ( .A(n21821), .B(n21820), .Z(n21823) );
  NANDN U22508 ( .A(n21670), .B(n21669), .Z(n21674) );
  NAND U22509 ( .A(n21672), .B(n21671), .Z(n21673) );
  NAND U22510 ( .A(n21674), .B(n21673), .Z(n21814) );
  NANDN U22511 ( .A(n21676), .B(n21675), .Z(n21680) );
  NAND U22512 ( .A(n21678), .B(n21677), .Z(n21679) );
  NAND U22513 ( .A(n21680), .B(n21679), .Z(n21815) );
  XNOR U22514 ( .A(n21814), .B(n21815), .Z(n21816) );
  XOR U22515 ( .A(n21817), .B(n21816), .Z(n21695) );
  XOR U22516 ( .A(n21694), .B(n21695), .Z(n21686) );
  XOR U22517 ( .A(n21687), .B(n21686), .Z(n21688) );
  XNOR U22518 ( .A(n21689), .B(n21688), .Z(n21826) );
  XNOR U22519 ( .A(n21826), .B(sreg[381]), .Z(n21828) );
  NAND U22520 ( .A(n21681), .B(sreg[380]), .Z(n21685) );
  OR U22521 ( .A(n21683), .B(n21682), .Z(n21684) );
  AND U22522 ( .A(n21685), .B(n21684), .Z(n21827) );
  XOR U22523 ( .A(n21828), .B(n21827), .Z(c[381]) );
  NAND U22524 ( .A(n21687), .B(n21686), .Z(n21691) );
  NAND U22525 ( .A(n21689), .B(n21688), .Z(n21690) );
  NAND U22526 ( .A(n21691), .B(n21690), .Z(n21834) );
  NANDN U22527 ( .A(n21693), .B(n21692), .Z(n21697) );
  NAND U22528 ( .A(n21695), .B(n21694), .Z(n21696) );
  NAND U22529 ( .A(n21697), .B(n21696), .Z(n21832) );
  NANDN U22530 ( .A(n21699), .B(n21698), .Z(n21703) );
  NAND U22531 ( .A(n21701), .B(n21700), .Z(n21702) );
  NAND U22532 ( .A(n21703), .B(n21702), .Z(n21912) );
  XNOR U22533 ( .A(b[19]), .B(a[140]), .Z(n21859) );
  NANDN U22534 ( .A(n21859), .B(n37934), .Z(n21706) );
  NANDN U22535 ( .A(n21704), .B(n37935), .Z(n21705) );
  NAND U22536 ( .A(n21706), .B(n21705), .Z(n21922) );
  XOR U22537 ( .A(b[27]), .B(a[132]), .Z(n21862) );
  NAND U22538 ( .A(n38423), .B(n21862), .Z(n21709) );
  NANDN U22539 ( .A(n21707), .B(n38424), .Z(n21708) );
  NAND U22540 ( .A(n21709), .B(n21708), .Z(n21919) );
  XOR U22541 ( .A(b[5]), .B(n25862), .Z(n21865) );
  NANDN U22542 ( .A(n21865), .B(n36587), .Z(n21712) );
  NANDN U22543 ( .A(n21710), .B(n36588), .Z(n21711) );
  AND U22544 ( .A(n21712), .B(n21711), .Z(n21920) );
  XNOR U22545 ( .A(n21919), .B(n21920), .Z(n21921) );
  XNOR U22546 ( .A(n21922), .B(n21921), .Z(n21910) );
  NANDN U22547 ( .A(n21713), .B(n37762), .Z(n21715) );
  XNOR U22548 ( .A(b[17]), .B(a[142]), .Z(n21868) );
  NANDN U22549 ( .A(n21868), .B(n37764), .Z(n21714) );
  NAND U22550 ( .A(n21715), .B(n21714), .Z(n21886) );
  XNOR U22551 ( .A(b[31]), .B(a[128]), .Z(n21871) );
  NANDN U22552 ( .A(n21871), .B(n38552), .Z(n21718) );
  NANDN U22553 ( .A(n21716), .B(n38553), .Z(n21717) );
  NAND U22554 ( .A(n21718), .B(n21717), .Z(n21883) );
  OR U22555 ( .A(n21719), .B(n36105), .Z(n21721) );
  XNOR U22556 ( .A(b[3]), .B(a[156]), .Z(n21874) );
  NANDN U22557 ( .A(n21874), .B(n36107), .Z(n21720) );
  AND U22558 ( .A(n21721), .B(n21720), .Z(n21884) );
  XNOR U22559 ( .A(n21883), .B(n21884), .Z(n21885) );
  XOR U22560 ( .A(n21886), .B(n21885), .Z(n21909) );
  XNOR U22561 ( .A(n21910), .B(n21909), .Z(n21911) );
  XNOR U22562 ( .A(n21912), .B(n21911), .Z(n21850) );
  NANDN U22563 ( .A(n21723), .B(n21722), .Z(n21727) );
  NAND U22564 ( .A(n21725), .B(n21724), .Z(n21726) );
  NAND U22565 ( .A(n21727), .B(n21726), .Z(n21901) );
  NANDN U22566 ( .A(n21729), .B(n21728), .Z(n21733) );
  NAND U22567 ( .A(n21731), .B(n21730), .Z(n21732) );
  NAND U22568 ( .A(n21733), .B(n21732), .Z(n21900) );
  XNOR U22569 ( .A(n21900), .B(n21899), .Z(n21902) );
  XOR U22570 ( .A(n21901), .B(n21902), .Z(n21849) );
  XOR U22571 ( .A(n21850), .B(n21849), .Z(n21851) );
  NANDN U22572 ( .A(n21739), .B(n21738), .Z(n21743) );
  NAND U22573 ( .A(n21741), .B(n21740), .Z(n21742) );
  NAND U22574 ( .A(n21743), .B(n21742), .Z(n21852) );
  XNOR U22575 ( .A(n21851), .B(n21852), .Z(n21963) );
  OR U22576 ( .A(n21745), .B(n21744), .Z(n21749) );
  NAND U22577 ( .A(n21747), .B(n21746), .Z(n21748) );
  NAND U22578 ( .A(n21749), .B(n21748), .Z(n21962) );
  NANDN U22579 ( .A(n21751), .B(n21750), .Z(n21755) );
  NAND U22580 ( .A(n21753), .B(n21752), .Z(n21754) );
  NAND U22581 ( .A(n21755), .B(n21754), .Z(n21845) );
  NANDN U22582 ( .A(n21761), .B(n21760), .Z(n21765) );
  NAND U22583 ( .A(n21763), .B(n21762), .Z(n21764) );
  NAND U22584 ( .A(n21765), .B(n21764), .Z(n21903) );
  NANDN U22585 ( .A(n21767), .B(n21766), .Z(n21771) );
  NAND U22586 ( .A(n21769), .B(n21768), .Z(n21770) );
  AND U22587 ( .A(n21771), .B(n21770), .Z(n21904) );
  XNOR U22588 ( .A(n21903), .B(n21904), .Z(n21905) );
  XNOR U22589 ( .A(b[21]), .B(a[138]), .Z(n21931) );
  NANDN U22590 ( .A(n21931), .B(n38101), .Z(n21774) );
  NANDN U22591 ( .A(n21772), .B(n38102), .Z(n21773) );
  NAND U22592 ( .A(n21774), .B(n21773), .Z(n21895) );
  XNOR U22593 ( .A(b[15]), .B(a[144]), .Z(n21928) );
  OR U22594 ( .A(n21928), .B(n37665), .Z(n21777) );
  NAND U22595 ( .A(n21775), .B(n37604), .Z(n21776) );
  AND U22596 ( .A(n21777), .B(n21776), .Z(n21896) );
  XNOR U22597 ( .A(n21895), .B(n21896), .Z(n21898) );
  XNOR U22598 ( .A(b[9]), .B(a[150]), .Z(n21925) );
  NANDN U22599 ( .A(n21925), .B(n36925), .Z(n21780) );
  NANDN U22600 ( .A(n21778), .B(n36926), .Z(n21779) );
  NAND U22601 ( .A(n21780), .B(n21779), .Z(n21897) );
  XNOR U22602 ( .A(n21898), .B(n21897), .Z(n21891) );
  XNOR U22603 ( .A(b[11]), .B(a[148]), .Z(n21934) );
  OR U22604 ( .A(n21934), .B(n37311), .Z(n21783) );
  NANDN U22605 ( .A(n21781), .B(n37218), .Z(n21782) );
  NAND U22606 ( .A(n21783), .B(n21782), .Z(n21890) );
  XOR U22607 ( .A(n1053), .B(a[146]), .Z(n21937) );
  NANDN U22608 ( .A(n21937), .B(n37424), .Z(n21786) );
  NANDN U22609 ( .A(n21784), .B(n37425), .Z(n21785) );
  NAND U22610 ( .A(n21786), .B(n21785), .Z(n21889) );
  XNOR U22611 ( .A(n21890), .B(n21889), .Z(n21892) );
  XNOR U22612 ( .A(n21891), .B(n21892), .Z(n21880) );
  NANDN U22613 ( .A(n1049), .B(a[158]), .Z(n21787) );
  XNOR U22614 ( .A(b[1]), .B(n21787), .Z(n21789) );
  NANDN U22615 ( .A(b[0]), .B(a[157]), .Z(n21788) );
  AND U22616 ( .A(n21789), .B(n21788), .Z(n21855) );
  NAND U22617 ( .A(n38490), .B(n21790), .Z(n21792) );
  XNOR U22618 ( .A(n1058), .B(a[130]), .Z(n21943) );
  NANDN U22619 ( .A(n1048), .B(n21943), .Z(n21791) );
  NAND U22620 ( .A(n21792), .B(n21791), .Z(n21853) );
  NANDN U22621 ( .A(n1059), .B(a[126]), .Z(n21854) );
  XNOR U22622 ( .A(n21853), .B(n21854), .Z(n21856) );
  XNOR U22623 ( .A(n21855), .B(n21856), .Z(n21878) );
  NANDN U22624 ( .A(n21793), .B(n38205), .Z(n21795) );
  XNOR U22625 ( .A(b[23]), .B(a[136]), .Z(n21946) );
  OR U22626 ( .A(n21946), .B(n38268), .Z(n21794) );
  NAND U22627 ( .A(n21795), .B(n21794), .Z(n21916) );
  XNOR U22628 ( .A(b[7]), .B(a[152]), .Z(n21949) );
  NANDN U22629 ( .A(n21949), .B(n36701), .Z(n21798) );
  NANDN U22630 ( .A(n21796), .B(n36702), .Z(n21797) );
  NAND U22631 ( .A(n21798), .B(n21797), .Z(n21913) );
  XOR U22632 ( .A(b[25]), .B(a[134]), .Z(n21952) );
  NAND U22633 ( .A(n21952), .B(n38325), .Z(n21801) );
  NAND U22634 ( .A(n21799), .B(n38326), .Z(n21800) );
  AND U22635 ( .A(n21801), .B(n21800), .Z(n21914) );
  XNOR U22636 ( .A(n21913), .B(n21914), .Z(n21915) );
  XOR U22637 ( .A(n21916), .B(n21915), .Z(n21877) );
  XOR U22638 ( .A(n21880), .B(n21879), .Z(n21906) );
  XNOR U22639 ( .A(n21905), .B(n21906), .Z(n21843) );
  XNOR U22640 ( .A(n21844), .B(n21843), .Z(n21846) );
  XNOR U22641 ( .A(n21845), .B(n21846), .Z(n21961) );
  XOR U22642 ( .A(n21962), .B(n21961), .Z(n21964) );
  NANDN U22643 ( .A(n21803), .B(n21802), .Z(n21807) );
  OR U22644 ( .A(n21805), .B(n21804), .Z(n21806) );
  NAND U22645 ( .A(n21807), .B(n21806), .Z(n21955) );
  NAND U22646 ( .A(n21809), .B(n21808), .Z(n21813) );
  NANDN U22647 ( .A(n21811), .B(n21810), .Z(n21812) );
  NAND U22648 ( .A(n21813), .B(n21812), .Z(n21956) );
  XNOR U22649 ( .A(n21955), .B(n21956), .Z(n21957) );
  XOR U22650 ( .A(n21958), .B(n21957), .Z(n21839) );
  NANDN U22651 ( .A(n21815), .B(n21814), .Z(n21819) );
  NAND U22652 ( .A(n21817), .B(n21816), .Z(n21818) );
  NAND U22653 ( .A(n21819), .B(n21818), .Z(n21837) );
  NANDN U22654 ( .A(n21821), .B(n21820), .Z(n21825) );
  OR U22655 ( .A(n21823), .B(n21822), .Z(n21824) );
  NAND U22656 ( .A(n21825), .B(n21824), .Z(n21838) );
  XNOR U22657 ( .A(n21837), .B(n21838), .Z(n21840) );
  XOR U22658 ( .A(n21839), .B(n21840), .Z(n21831) );
  XOR U22659 ( .A(n21832), .B(n21831), .Z(n21833) );
  XNOR U22660 ( .A(n21834), .B(n21833), .Z(n21967) );
  XNOR U22661 ( .A(n21967), .B(sreg[382]), .Z(n21969) );
  NAND U22662 ( .A(n21826), .B(sreg[381]), .Z(n21830) );
  OR U22663 ( .A(n21828), .B(n21827), .Z(n21829) );
  AND U22664 ( .A(n21830), .B(n21829), .Z(n21968) );
  XOR U22665 ( .A(n21969), .B(n21968), .Z(c[382]) );
  NAND U22666 ( .A(n21832), .B(n21831), .Z(n21836) );
  NAND U22667 ( .A(n21834), .B(n21833), .Z(n21835) );
  NAND U22668 ( .A(n21836), .B(n21835), .Z(n21975) );
  NANDN U22669 ( .A(n21838), .B(n21837), .Z(n21842) );
  NAND U22670 ( .A(n21840), .B(n21839), .Z(n21841) );
  NAND U22671 ( .A(n21842), .B(n21841), .Z(n21972) );
  NAND U22672 ( .A(n21844), .B(n21843), .Z(n21848) );
  NANDN U22673 ( .A(n21846), .B(n21845), .Z(n21847) );
  NAND U22674 ( .A(n21848), .B(n21847), .Z(n22100) );
  XNOR U22675 ( .A(n22100), .B(n22101), .Z(n22102) );
  NANDN U22676 ( .A(n21854), .B(n21853), .Z(n21858) );
  NAND U22677 ( .A(n21856), .B(n21855), .Z(n21857) );
  NAND U22678 ( .A(n21858), .B(n21857), .Z(n22045) );
  XOR U22679 ( .A(b[19]), .B(n23961), .Z(n21990) );
  NANDN U22680 ( .A(n21990), .B(n37934), .Z(n21861) );
  NANDN U22681 ( .A(n21859), .B(n37935), .Z(n21860) );
  NAND U22682 ( .A(n21861), .B(n21860), .Z(n22055) );
  XOR U22683 ( .A(b[27]), .B(a[133]), .Z(n21993) );
  NAND U22684 ( .A(n38423), .B(n21993), .Z(n21864) );
  NAND U22685 ( .A(n21862), .B(n38424), .Z(n21863) );
  NAND U22686 ( .A(n21864), .B(n21863), .Z(n22052) );
  XNOR U22687 ( .A(b[5]), .B(a[155]), .Z(n21996) );
  NANDN U22688 ( .A(n21996), .B(n36587), .Z(n21867) );
  NANDN U22689 ( .A(n21865), .B(n36588), .Z(n21866) );
  AND U22690 ( .A(n21867), .B(n21866), .Z(n22053) );
  XNOR U22691 ( .A(n22052), .B(n22053), .Z(n22054) );
  XNOR U22692 ( .A(n22055), .B(n22054), .Z(n22043) );
  NANDN U22693 ( .A(n21868), .B(n37762), .Z(n21870) );
  XOR U22694 ( .A(b[17]), .B(a[143]), .Z(n21999) );
  NAND U22695 ( .A(n21999), .B(n37764), .Z(n21869) );
  NAND U22696 ( .A(n21870), .B(n21869), .Z(n22017) );
  XOR U22697 ( .A(b[31]), .B(n22221), .Z(n22002) );
  NANDN U22698 ( .A(n22002), .B(n38552), .Z(n21873) );
  NANDN U22699 ( .A(n21871), .B(n38553), .Z(n21872) );
  NAND U22700 ( .A(n21873), .B(n21872), .Z(n22014) );
  OR U22701 ( .A(n21874), .B(n36105), .Z(n21876) );
  XNOR U22702 ( .A(b[3]), .B(a[157]), .Z(n22005) );
  NANDN U22703 ( .A(n22005), .B(n36107), .Z(n21875) );
  AND U22704 ( .A(n21876), .B(n21875), .Z(n22015) );
  XNOR U22705 ( .A(n22014), .B(n22015), .Z(n22016) );
  XOR U22706 ( .A(n22017), .B(n22016), .Z(n22042) );
  XNOR U22707 ( .A(n22043), .B(n22042), .Z(n22044) );
  XNOR U22708 ( .A(n22045), .B(n22044), .Z(n22094) );
  NANDN U22709 ( .A(n21878), .B(n21877), .Z(n21882) );
  NANDN U22710 ( .A(n21880), .B(n21879), .Z(n21881) );
  NAND U22711 ( .A(n21882), .B(n21881), .Z(n22095) );
  XNOR U22712 ( .A(n22094), .B(n22095), .Z(n22096) );
  NANDN U22713 ( .A(n21884), .B(n21883), .Z(n21888) );
  NAND U22714 ( .A(n21886), .B(n21885), .Z(n21887) );
  NAND U22715 ( .A(n21888), .B(n21887), .Z(n22035) );
  OR U22716 ( .A(n21890), .B(n21889), .Z(n21894) );
  NANDN U22717 ( .A(n21892), .B(n21891), .Z(n21893) );
  NAND U22718 ( .A(n21894), .B(n21893), .Z(n22033) );
  XNOR U22719 ( .A(n22033), .B(n22032), .Z(n22034) );
  XOR U22720 ( .A(n22035), .B(n22034), .Z(n22097) );
  XOR U22721 ( .A(n22096), .B(n22097), .Z(n22108) );
  NANDN U22722 ( .A(n21904), .B(n21903), .Z(n21908) );
  NANDN U22723 ( .A(n21906), .B(n21905), .Z(n21907) );
  NAND U22724 ( .A(n21908), .B(n21907), .Z(n22091) );
  NANDN U22725 ( .A(n21914), .B(n21913), .Z(n21918) );
  NAND U22726 ( .A(n21916), .B(n21915), .Z(n21917) );
  NAND U22727 ( .A(n21918), .B(n21917), .Z(n22036) );
  NANDN U22728 ( .A(n21920), .B(n21919), .Z(n21924) );
  NAND U22729 ( .A(n21922), .B(n21921), .Z(n21923) );
  AND U22730 ( .A(n21924), .B(n21923), .Z(n22037) );
  XNOR U22731 ( .A(n22036), .B(n22037), .Z(n22038) );
  XOR U22732 ( .A(b[9]), .B(n25435), .Z(n22058) );
  NANDN U22733 ( .A(n22058), .B(n36925), .Z(n21927) );
  NANDN U22734 ( .A(n21925), .B(n36926), .Z(n21926) );
  NAND U22735 ( .A(n21927), .B(n21926), .Z(n22022) );
  XOR U22736 ( .A(b[15]), .B(n24554), .Z(n22061) );
  OR U22737 ( .A(n22061), .B(n37665), .Z(n21930) );
  NANDN U22738 ( .A(n21928), .B(n37604), .Z(n21929) );
  AND U22739 ( .A(n21930), .B(n21929), .Z(n22020) );
  XOR U22740 ( .A(b[21]), .B(n23668), .Z(n22064) );
  NANDN U22741 ( .A(n22064), .B(n38101), .Z(n21933) );
  NANDN U22742 ( .A(n21931), .B(n38102), .Z(n21932) );
  AND U22743 ( .A(n21933), .B(n21932), .Z(n22021) );
  XOR U22744 ( .A(n22022), .B(n22023), .Z(n22011) );
  XNOR U22745 ( .A(b[11]), .B(a[149]), .Z(n22067) );
  OR U22746 ( .A(n22067), .B(n37311), .Z(n21936) );
  NANDN U22747 ( .A(n21934), .B(n37218), .Z(n21935) );
  NAND U22748 ( .A(n21936), .B(n21935), .Z(n22009) );
  XOR U22749 ( .A(n1053), .B(a[147]), .Z(n22070) );
  NANDN U22750 ( .A(n22070), .B(n37424), .Z(n21939) );
  NANDN U22751 ( .A(n21937), .B(n37425), .Z(n21938) );
  AND U22752 ( .A(n21939), .B(n21938), .Z(n22008) );
  XNOR U22753 ( .A(n22009), .B(n22008), .Z(n22010) );
  XOR U22754 ( .A(n22011), .B(n22010), .Z(n22028) );
  NANDN U22755 ( .A(n1049), .B(a[159]), .Z(n21940) );
  XNOR U22756 ( .A(b[1]), .B(n21940), .Z(n21942) );
  NANDN U22757 ( .A(b[0]), .B(a[158]), .Z(n21941) );
  AND U22758 ( .A(n21942), .B(n21941), .Z(n21986) );
  NAND U22759 ( .A(n38490), .B(n21943), .Z(n21945) );
  XOR U22760 ( .A(n1058), .B(n22518), .Z(n22076) );
  NANDN U22761 ( .A(n1048), .B(n22076), .Z(n21944) );
  NAND U22762 ( .A(n21945), .B(n21944), .Z(n21984) );
  NANDN U22763 ( .A(n1059), .B(a[127]), .Z(n21985) );
  XNOR U22764 ( .A(n21984), .B(n21985), .Z(n21987) );
  XOR U22765 ( .A(n21986), .B(n21987), .Z(n22026) );
  NANDN U22766 ( .A(n21946), .B(n38205), .Z(n21948) );
  XOR U22767 ( .A(b[23]), .B(n23393), .Z(n22079) );
  OR U22768 ( .A(n22079), .B(n38268), .Z(n21947) );
  NAND U22769 ( .A(n21948), .B(n21947), .Z(n22049) );
  XOR U22770 ( .A(b[7]), .B(a[153]), .Z(n22082) );
  NAND U22771 ( .A(n22082), .B(n36701), .Z(n21951) );
  NANDN U22772 ( .A(n21949), .B(n36702), .Z(n21950) );
  NAND U22773 ( .A(n21951), .B(n21950), .Z(n22046) );
  XOR U22774 ( .A(b[25]), .B(a[135]), .Z(n22085) );
  NAND U22775 ( .A(n22085), .B(n38325), .Z(n21954) );
  NAND U22776 ( .A(n21952), .B(n38326), .Z(n21953) );
  AND U22777 ( .A(n21954), .B(n21953), .Z(n22047) );
  XNOR U22778 ( .A(n22046), .B(n22047), .Z(n22048) );
  XNOR U22779 ( .A(n22049), .B(n22048), .Z(n22027) );
  XOR U22780 ( .A(n22026), .B(n22027), .Z(n22029) );
  XNOR U22781 ( .A(n22028), .B(n22029), .Z(n22039) );
  XOR U22782 ( .A(n22038), .B(n22039), .Z(n22089) );
  XNOR U22783 ( .A(n22088), .B(n22089), .Z(n22090) );
  XNOR U22784 ( .A(n22091), .B(n22090), .Z(n22106) );
  XNOR U22785 ( .A(n22107), .B(n22106), .Z(n22109) );
  XNOR U22786 ( .A(n22108), .B(n22109), .Z(n22103) );
  XOR U22787 ( .A(n22102), .B(n22103), .Z(n21981) );
  NANDN U22788 ( .A(n21956), .B(n21955), .Z(n21960) );
  NAND U22789 ( .A(n21958), .B(n21957), .Z(n21959) );
  NAND U22790 ( .A(n21960), .B(n21959), .Z(n21978) );
  NANDN U22791 ( .A(n21962), .B(n21961), .Z(n21966) );
  OR U22792 ( .A(n21964), .B(n21963), .Z(n21965) );
  NAND U22793 ( .A(n21966), .B(n21965), .Z(n21979) );
  XNOR U22794 ( .A(n21978), .B(n21979), .Z(n21980) );
  XNOR U22795 ( .A(n21981), .B(n21980), .Z(n21973) );
  XNOR U22796 ( .A(n21972), .B(n21973), .Z(n21974) );
  XNOR U22797 ( .A(n21975), .B(n21974), .Z(n22112) );
  XNOR U22798 ( .A(n22112), .B(sreg[383]), .Z(n22114) );
  NAND U22799 ( .A(n21967), .B(sreg[382]), .Z(n21971) );
  OR U22800 ( .A(n21969), .B(n21968), .Z(n21970) );
  AND U22801 ( .A(n21971), .B(n21970), .Z(n22113) );
  XOR U22802 ( .A(n22114), .B(n22113), .Z(c[383]) );
  NANDN U22803 ( .A(n21973), .B(n21972), .Z(n21977) );
  NAND U22804 ( .A(n21975), .B(n21974), .Z(n21976) );
  NAND U22805 ( .A(n21977), .B(n21976), .Z(n22120) );
  NANDN U22806 ( .A(n21979), .B(n21978), .Z(n21983) );
  NAND U22807 ( .A(n21981), .B(n21980), .Z(n21982) );
  NAND U22808 ( .A(n21983), .B(n21982), .Z(n22118) );
  NANDN U22809 ( .A(n21985), .B(n21984), .Z(n21989) );
  NAND U22810 ( .A(n21987), .B(n21986), .Z(n21988) );
  NAND U22811 ( .A(n21989), .B(n21988), .Z(n22190) );
  XOR U22812 ( .A(b[19]), .B(n24120), .Z(n22133) );
  NANDN U22813 ( .A(n22133), .B(n37934), .Z(n21992) );
  NANDN U22814 ( .A(n21990), .B(n37935), .Z(n21991) );
  NAND U22815 ( .A(n21992), .B(n21991), .Z(n22200) );
  XOR U22816 ( .A(b[27]), .B(a[134]), .Z(n22136) );
  NAND U22817 ( .A(n38423), .B(n22136), .Z(n21995) );
  NAND U22818 ( .A(n21993), .B(n38424), .Z(n21994) );
  NAND U22819 ( .A(n21995), .B(n21994), .Z(n22197) );
  XNOR U22820 ( .A(b[5]), .B(a[156]), .Z(n22139) );
  NANDN U22821 ( .A(n22139), .B(n36587), .Z(n21998) );
  NANDN U22822 ( .A(n21996), .B(n36588), .Z(n21997) );
  AND U22823 ( .A(n21998), .B(n21997), .Z(n22198) );
  XNOR U22824 ( .A(n22197), .B(n22198), .Z(n22199) );
  XNOR U22825 ( .A(n22200), .B(n22199), .Z(n22188) );
  NAND U22826 ( .A(n21999), .B(n37762), .Z(n22001) );
  XOR U22827 ( .A(b[17]), .B(a[144]), .Z(n22142) );
  NAND U22828 ( .A(n22142), .B(n37764), .Z(n22000) );
  NAND U22829 ( .A(n22001), .B(n22000), .Z(n22160) );
  XNOR U22830 ( .A(b[31]), .B(a[130]), .Z(n22145) );
  NANDN U22831 ( .A(n22145), .B(n38552), .Z(n22004) );
  NANDN U22832 ( .A(n22002), .B(n38553), .Z(n22003) );
  NAND U22833 ( .A(n22004), .B(n22003), .Z(n22157) );
  OR U22834 ( .A(n22005), .B(n36105), .Z(n22007) );
  XNOR U22835 ( .A(b[3]), .B(a[158]), .Z(n22148) );
  NANDN U22836 ( .A(n22148), .B(n36107), .Z(n22006) );
  AND U22837 ( .A(n22007), .B(n22006), .Z(n22158) );
  XNOR U22838 ( .A(n22157), .B(n22158), .Z(n22159) );
  XOR U22839 ( .A(n22160), .B(n22159), .Z(n22187) );
  XNOR U22840 ( .A(n22188), .B(n22187), .Z(n22189) );
  XNOR U22841 ( .A(n22190), .B(n22189), .Z(n22234) );
  NANDN U22842 ( .A(n22009), .B(n22008), .Z(n22013) );
  NAND U22843 ( .A(n22011), .B(n22010), .Z(n22012) );
  NAND U22844 ( .A(n22013), .B(n22012), .Z(n22178) );
  NANDN U22845 ( .A(n22015), .B(n22014), .Z(n22019) );
  NAND U22846 ( .A(n22017), .B(n22016), .Z(n22018) );
  NAND U22847 ( .A(n22019), .B(n22018), .Z(n22176) );
  OR U22848 ( .A(n22021), .B(n22020), .Z(n22025) );
  NANDN U22849 ( .A(n22023), .B(n22022), .Z(n22024) );
  NAND U22850 ( .A(n22025), .B(n22024), .Z(n22175) );
  XNOR U22851 ( .A(n22178), .B(n22177), .Z(n22235) );
  XNOR U22852 ( .A(n22234), .B(n22235), .Z(n22236) );
  NANDN U22853 ( .A(n22027), .B(n22026), .Z(n22031) );
  OR U22854 ( .A(n22029), .B(n22028), .Z(n22030) );
  AND U22855 ( .A(n22031), .B(n22030), .Z(n22237) );
  XNOR U22856 ( .A(n22236), .B(n22237), .Z(n22249) );
  NANDN U22857 ( .A(n22037), .B(n22036), .Z(n22041) );
  NANDN U22858 ( .A(n22039), .B(n22038), .Z(n22040) );
  NAND U22859 ( .A(n22041), .B(n22040), .Z(n22243) );
  NANDN U22860 ( .A(n22047), .B(n22046), .Z(n22051) );
  NAND U22861 ( .A(n22049), .B(n22048), .Z(n22050) );
  NAND U22862 ( .A(n22051), .B(n22050), .Z(n22181) );
  NANDN U22863 ( .A(n22053), .B(n22052), .Z(n22057) );
  NAND U22864 ( .A(n22055), .B(n22054), .Z(n22056) );
  AND U22865 ( .A(n22057), .B(n22056), .Z(n22182) );
  XNOR U22866 ( .A(n22181), .B(n22182), .Z(n22183) );
  XOR U22867 ( .A(b[9]), .B(n25213), .Z(n22203) );
  NANDN U22868 ( .A(n22203), .B(n36925), .Z(n22060) );
  NANDN U22869 ( .A(n22058), .B(n36926), .Z(n22059) );
  NAND U22870 ( .A(n22060), .B(n22059), .Z(n22165) );
  XNOR U22871 ( .A(b[15]), .B(a[146]), .Z(n22206) );
  OR U22872 ( .A(n22206), .B(n37665), .Z(n22063) );
  NANDN U22873 ( .A(n22061), .B(n37604), .Z(n22062) );
  AND U22874 ( .A(n22063), .B(n22062), .Z(n22163) );
  XNOR U22875 ( .A(b[21]), .B(a[140]), .Z(n22209) );
  NANDN U22876 ( .A(n22209), .B(n38101), .Z(n22066) );
  NANDN U22877 ( .A(n22064), .B(n38102), .Z(n22065) );
  AND U22878 ( .A(n22066), .B(n22065), .Z(n22164) );
  XOR U22879 ( .A(n22165), .B(n22166), .Z(n22154) );
  XNOR U22880 ( .A(b[11]), .B(a[150]), .Z(n22212) );
  OR U22881 ( .A(n22212), .B(n37311), .Z(n22069) );
  NANDN U22882 ( .A(n22067), .B(n37218), .Z(n22068) );
  NAND U22883 ( .A(n22069), .B(n22068), .Z(n22152) );
  XOR U22884 ( .A(n1053), .B(a[148]), .Z(n22215) );
  NANDN U22885 ( .A(n22215), .B(n37424), .Z(n22072) );
  NANDN U22886 ( .A(n22070), .B(n37425), .Z(n22071) );
  AND U22887 ( .A(n22072), .B(n22071), .Z(n22151) );
  XNOR U22888 ( .A(n22152), .B(n22151), .Z(n22153) );
  XOR U22889 ( .A(n22154), .B(n22153), .Z(n22171) );
  NANDN U22890 ( .A(n1049), .B(a[160]), .Z(n22073) );
  XNOR U22891 ( .A(b[1]), .B(n22073), .Z(n22075) );
  NANDN U22892 ( .A(b[0]), .B(a[159]), .Z(n22074) );
  AND U22893 ( .A(n22075), .B(n22074), .Z(n22129) );
  NAND U22894 ( .A(n38490), .B(n22076), .Z(n22078) );
  XNOR U22895 ( .A(b[29]), .B(a[132]), .Z(n22222) );
  OR U22896 ( .A(n22222), .B(n1048), .Z(n22077) );
  NAND U22897 ( .A(n22078), .B(n22077), .Z(n22127) );
  NANDN U22898 ( .A(n1059), .B(a[128]), .Z(n22128) );
  XNOR U22899 ( .A(n22127), .B(n22128), .Z(n22130) );
  XOR U22900 ( .A(n22129), .B(n22130), .Z(n22169) );
  NANDN U22901 ( .A(n22079), .B(n38205), .Z(n22081) );
  XNOR U22902 ( .A(b[23]), .B(a[138]), .Z(n22225) );
  OR U22903 ( .A(n22225), .B(n38268), .Z(n22080) );
  NAND U22904 ( .A(n22081), .B(n22080), .Z(n22194) );
  XNOR U22905 ( .A(b[7]), .B(a[154]), .Z(n22228) );
  NANDN U22906 ( .A(n22228), .B(n36701), .Z(n22084) );
  NAND U22907 ( .A(n22082), .B(n36702), .Z(n22083) );
  NAND U22908 ( .A(n22084), .B(n22083), .Z(n22191) );
  XOR U22909 ( .A(b[25]), .B(a[136]), .Z(n22231) );
  NAND U22910 ( .A(n22231), .B(n38325), .Z(n22087) );
  NAND U22911 ( .A(n22085), .B(n38326), .Z(n22086) );
  AND U22912 ( .A(n22087), .B(n22086), .Z(n22192) );
  XNOR U22913 ( .A(n22191), .B(n22192), .Z(n22193) );
  XNOR U22914 ( .A(n22194), .B(n22193), .Z(n22170) );
  XOR U22915 ( .A(n22169), .B(n22170), .Z(n22172) );
  XNOR U22916 ( .A(n22171), .B(n22172), .Z(n22184) );
  XOR U22917 ( .A(n22183), .B(n22184), .Z(n22241) );
  XNOR U22918 ( .A(n22240), .B(n22241), .Z(n22242) );
  XOR U22919 ( .A(n22243), .B(n22242), .Z(n22247) );
  XNOR U22920 ( .A(n22246), .B(n22247), .Z(n22248) );
  XNOR U22921 ( .A(n22249), .B(n22248), .Z(n22253) );
  NANDN U22922 ( .A(n22089), .B(n22088), .Z(n22093) );
  NAND U22923 ( .A(n22091), .B(n22090), .Z(n22092) );
  NAND U22924 ( .A(n22093), .B(n22092), .Z(n22250) );
  NANDN U22925 ( .A(n22095), .B(n22094), .Z(n22099) );
  NAND U22926 ( .A(n22097), .B(n22096), .Z(n22098) );
  NAND U22927 ( .A(n22099), .B(n22098), .Z(n22251) );
  XNOR U22928 ( .A(n22250), .B(n22251), .Z(n22252) );
  XNOR U22929 ( .A(n22253), .B(n22252), .Z(n22124) );
  NANDN U22930 ( .A(n22101), .B(n22100), .Z(n22105) );
  NANDN U22931 ( .A(n22103), .B(n22102), .Z(n22104) );
  NAND U22932 ( .A(n22105), .B(n22104), .Z(n22122) );
  OR U22933 ( .A(n22107), .B(n22106), .Z(n22111) );
  OR U22934 ( .A(n22109), .B(n22108), .Z(n22110) );
  AND U22935 ( .A(n22111), .B(n22110), .Z(n22121) );
  XNOR U22936 ( .A(n22122), .B(n22121), .Z(n22123) );
  XNOR U22937 ( .A(n22124), .B(n22123), .Z(n22117) );
  XOR U22938 ( .A(n22118), .B(n22117), .Z(n22119) );
  XNOR U22939 ( .A(n22120), .B(n22119), .Z(n22256) );
  XNOR U22940 ( .A(n22256), .B(sreg[384]), .Z(n22258) );
  NAND U22941 ( .A(n22112), .B(sreg[383]), .Z(n22116) );
  OR U22942 ( .A(n22114), .B(n22113), .Z(n22115) );
  AND U22943 ( .A(n22116), .B(n22115), .Z(n22257) );
  XOR U22944 ( .A(n22258), .B(n22257), .Z(c[384]) );
  NANDN U22945 ( .A(n22122), .B(n22121), .Z(n22126) );
  NANDN U22946 ( .A(n22124), .B(n22123), .Z(n22125) );
  NAND U22947 ( .A(n22126), .B(n22125), .Z(n22262) );
  NANDN U22948 ( .A(n22128), .B(n22127), .Z(n22132) );
  NAND U22949 ( .A(n22130), .B(n22129), .Z(n22131) );
  NAND U22950 ( .A(n22132), .B(n22131), .Z(n22348) );
  XNOR U22951 ( .A(b[19]), .B(a[143]), .Z(n22315) );
  NANDN U22952 ( .A(n22315), .B(n37934), .Z(n22135) );
  NANDN U22953 ( .A(n22133), .B(n37935), .Z(n22134) );
  NAND U22954 ( .A(n22135), .B(n22134), .Z(n22384) );
  XOR U22955 ( .A(b[27]), .B(a[135]), .Z(n22318) );
  NAND U22956 ( .A(n38423), .B(n22318), .Z(n22138) );
  NAND U22957 ( .A(n22136), .B(n38424), .Z(n22137) );
  NAND U22958 ( .A(n22138), .B(n22137), .Z(n22381) );
  XNOR U22959 ( .A(b[5]), .B(a[157]), .Z(n22321) );
  NANDN U22960 ( .A(n22321), .B(n36587), .Z(n22141) );
  NANDN U22961 ( .A(n22139), .B(n36588), .Z(n22140) );
  AND U22962 ( .A(n22141), .B(n22140), .Z(n22382) );
  XNOR U22963 ( .A(n22381), .B(n22382), .Z(n22383) );
  XNOR U22964 ( .A(n22384), .B(n22383), .Z(n22345) );
  NAND U22965 ( .A(n22142), .B(n37762), .Z(n22144) );
  XNOR U22966 ( .A(b[17]), .B(a[145]), .Z(n22324) );
  NANDN U22967 ( .A(n22324), .B(n37764), .Z(n22143) );
  NAND U22968 ( .A(n22144), .B(n22143), .Z(n22299) );
  XOR U22969 ( .A(b[31]), .B(n22518), .Z(n22327) );
  NANDN U22970 ( .A(n22327), .B(n38552), .Z(n22147) );
  NANDN U22971 ( .A(n22145), .B(n38553), .Z(n22146) );
  AND U22972 ( .A(n22147), .B(n22146), .Z(n22297) );
  OR U22973 ( .A(n22148), .B(n36105), .Z(n22150) );
  XNOR U22974 ( .A(b[3]), .B(a[159]), .Z(n22330) );
  NANDN U22975 ( .A(n22330), .B(n36107), .Z(n22149) );
  AND U22976 ( .A(n22150), .B(n22149), .Z(n22298) );
  XOR U22977 ( .A(n22299), .B(n22300), .Z(n22346) );
  XOR U22978 ( .A(n22345), .B(n22346), .Z(n22347) );
  XNOR U22979 ( .A(n22348), .B(n22347), .Z(n22393) );
  NANDN U22980 ( .A(n22152), .B(n22151), .Z(n22156) );
  NAND U22981 ( .A(n22154), .B(n22153), .Z(n22155) );
  NAND U22982 ( .A(n22156), .B(n22155), .Z(n22336) );
  NANDN U22983 ( .A(n22158), .B(n22157), .Z(n22162) );
  NAND U22984 ( .A(n22160), .B(n22159), .Z(n22161) );
  NAND U22985 ( .A(n22162), .B(n22161), .Z(n22334) );
  OR U22986 ( .A(n22164), .B(n22163), .Z(n22168) );
  NANDN U22987 ( .A(n22166), .B(n22165), .Z(n22167) );
  NAND U22988 ( .A(n22168), .B(n22167), .Z(n22333) );
  XNOR U22989 ( .A(n22336), .B(n22335), .Z(n22394) );
  XOR U22990 ( .A(n22393), .B(n22394), .Z(n22396) );
  NANDN U22991 ( .A(n22170), .B(n22169), .Z(n22174) );
  OR U22992 ( .A(n22172), .B(n22171), .Z(n22173) );
  NAND U22993 ( .A(n22174), .B(n22173), .Z(n22395) );
  XOR U22994 ( .A(n22396), .B(n22395), .Z(n22281) );
  OR U22995 ( .A(n22176), .B(n22175), .Z(n22180) );
  NAND U22996 ( .A(n22178), .B(n22177), .Z(n22179) );
  NAND U22997 ( .A(n22180), .B(n22179), .Z(n22280) );
  NANDN U22998 ( .A(n22182), .B(n22181), .Z(n22186) );
  NANDN U22999 ( .A(n22184), .B(n22183), .Z(n22185) );
  NAND U23000 ( .A(n22186), .B(n22185), .Z(n22401) );
  NANDN U23001 ( .A(n22192), .B(n22191), .Z(n22196) );
  NAND U23002 ( .A(n22194), .B(n22193), .Z(n22195) );
  NAND U23003 ( .A(n22196), .B(n22195), .Z(n22339) );
  NANDN U23004 ( .A(n22198), .B(n22197), .Z(n22202) );
  NAND U23005 ( .A(n22200), .B(n22199), .Z(n22201) );
  AND U23006 ( .A(n22202), .B(n22201), .Z(n22340) );
  XNOR U23007 ( .A(n22339), .B(n22340), .Z(n22341) );
  XNOR U23008 ( .A(b[9]), .B(a[153]), .Z(n22351) );
  NANDN U23009 ( .A(n22351), .B(n36925), .Z(n22205) );
  NANDN U23010 ( .A(n22203), .B(n36926), .Z(n22204) );
  NAND U23011 ( .A(n22205), .B(n22204), .Z(n22305) );
  XNOR U23012 ( .A(b[15]), .B(a[147]), .Z(n22354) );
  OR U23013 ( .A(n22354), .B(n37665), .Z(n22208) );
  NANDN U23014 ( .A(n22206), .B(n37604), .Z(n22207) );
  AND U23015 ( .A(n22208), .B(n22207), .Z(n22303) );
  XOR U23016 ( .A(b[21]), .B(n23961), .Z(n22357) );
  NANDN U23017 ( .A(n22357), .B(n38101), .Z(n22211) );
  NANDN U23018 ( .A(n22209), .B(n38102), .Z(n22210) );
  AND U23019 ( .A(n22211), .B(n22210), .Z(n22304) );
  XOR U23020 ( .A(n22305), .B(n22306), .Z(n22294) );
  XOR U23021 ( .A(b[11]), .B(n25435), .Z(n22360) );
  OR U23022 ( .A(n22360), .B(n37311), .Z(n22214) );
  NANDN U23023 ( .A(n22212), .B(n37218), .Z(n22213) );
  NAND U23024 ( .A(n22214), .B(n22213), .Z(n22292) );
  XOR U23025 ( .A(n1053), .B(a[149]), .Z(n22363) );
  NANDN U23026 ( .A(n22363), .B(n37424), .Z(n22217) );
  NANDN U23027 ( .A(n22215), .B(n37425), .Z(n22216) );
  NAND U23028 ( .A(n22217), .B(n22216), .Z(n22291) );
  XOR U23029 ( .A(n22294), .B(n22293), .Z(n22288) );
  NANDN U23030 ( .A(n1049), .B(a[161]), .Z(n22218) );
  XNOR U23031 ( .A(b[1]), .B(n22218), .Z(n22220) );
  NANDN U23032 ( .A(b[0]), .B(a[160]), .Z(n22219) );
  AND U23033 ( .A(n22220), .B(n22219), .Z(n22312) );
  ANDN U23034 ( .B(b[31]), .A(n22221), .Z(n22309) );
  NANDN U23035 ( .A(n22222), .B(n38490), .Z(n22224) );
  XNOR U23036 ( .A(n1058), .B(a[133]), .Z(n22369) );
  NANDN U23037 ( .A(n1048), .B(n22369), .Z(n22223) );
  NAND U23038 ( .A(n22224), .B(n22223), .Z(n22310) );
  XOR U23039 ( .A(n22309), .B(n22310), .Z(n22311) );
  XNOR U23040 ( .A(n22312), .B(n22311), .Z(n22285) );
  NANDN U23041 ( .A(n22225), .B(n38205), .Z(n22227) );
  XOR U23042 ( .A(b[23]), .B(n23668), .Z(n22372) );
  OR U23043 ( .A(n22372), .B(n38268), .Z(n22226) );
  NAND U23044 ( .A(n22227), .B(n22226), .Z(n22390) );
  XOR U23045 ( .A(b[7]), .B(a[155]), .Z(n22375) );
  NAND U23046 ( .A(n22375), .B(n36701), .Z(n22230) );
  NANDN U23047 ( .A(n22228), .B(n36702), .Z(n22229) );
  NAND U23048 ( .A(n22230), .B(n22229), .Z(n22387) );
  XNOR U23049 ( .A(b[25]), .B(a[137]), .Z(n22378) );
  NANDN U23050 ( .A(n22378), .B(n38325), .Z(n22233) );
  NAND U23051 ( .A(n22231), .B(n38326), .Z(n22232) );
  AND U23052 ( .A(n22233), .B(n22232), .Z(n22388) );
  XNOR U23053 ( .A(n22387), .B(n22388), .Z(n22389) );
  XNOR U23054 ( .A(n22390), .B(n22389), .Z(n22286) );
  XOR U23055 ( .A(n22288), .B(n22287), .Z(n22342) );
  XNOR U23056 ( .A(n22341), .B(n22342), .Z(n22399) );
  XNOR U23057 ( .A(n22400), .B(n22399), .Z(n22402) );
  XNOR U23058 ( .A(n22401), .B(n22402), .Z(n22279) );
  XOR U23059 ( .A(n22280), .B(n22279), .Z(n22282) );
  NANDN U23060 ( .A(n22235), .B(n22234), .Z(n22239) );
  NAND U23061 ( .A(n22237), .B(n22236), .Z(n22238) );
  NAND U23062 ( .A(n22239), .B(n22238), .Z(n22273) );
  NANDN U23063 ( .A(n22241), .B(n22240), .Z(n22245) );
  NAND U23064 ( .A(n22243), .B(n22242), .Z(n22244) );
  NAND U23065 ( .A(n22245), .B(n22244), .Z(n22274) );
  XNOR U23066 ( .A(n22273), .B(n22274), .Z(n22275) );
  XOR U23067 ( .A(n22276), .B(n22275), .Z(n22269) );
  NANDN U23068 ( .A(n22251), .B(n22250), .Z(n22255) );
  NANDN U23069 ( .A(n22253), .B(n22252), .Z(n22254) );
  NAND U23070 ( .A(n22255), .B(n22254), .Z(n22268) );
  XNOR U23071 ( .A(n22267), .B(n22268), .Z(n22270) );
  XOR U23072 ( .A(n22269), .B(n22270), .Z(n22261) );
  XOR U23073 ( .A(n22262), .B(n22261), .Z(n22263) );
  XNOR U23074 ( .A(n22264), .B(n22263), .Z(n22405) );
  XNOR U23075 ( .A(n22405), .B(sreg[385]), .Z(n22407) );
  NAND U23076 ( .A(n22256), .B(sreg[384]), .Z(n22260) );
  OR U23077 ( .A(n22258), .B(n22257), .Z(n22259) );
  AND U23078 ( .A(n22260), .B(n22259), .Z(n22406) );
  XOR U23079 ( .A(n22407), .B(n22406), .Z(c[385]) );
  NAND U23080 ( .A(n22262), .B(n22261), .Z(n22266) );
  NAND U23081 ( .A(n22264), .B(n22263), .Z(n22265) );
  NAND U23082 ( .A(n22266), .B(n22265), .Z(n22413) );
  NANDN U23083 ( .A(n22268), .B(n22267), .Z(n22272) );
  NAND U23084 ( .A(n22270), .B(n22269), .Z(n22271) );
  NAND U23085 ( .A(n22272), .B(n22271), .Z(n22411) );
  NANDN U23086 ( .A(n22274), .B(n22273), .Z(n22278) );
  NAND U23087 ( .A(n22276), .B(n22275), .Z(n22277) );
  NAND U23088 ( .A(n22278), .B(n22277), .Z(n22416) );
  NANDN U23089 ( .A(n22280), .B(n22279), .Z(n22284) );
  OR U23090 ( .A(n22282), .B(n22281), .Z(n22283) );
  NAND U23091 ( .A(n22284), .B(n22283), .Z(n22417) );
  XNOR U23092 ( .A(n22416), .B(n22417), .Z(n22418) );
  OR U23093 ( .A(n22286), .B(n22285), .Z(n22290) );
  NANDN U23094 ( .A(n22288), .B(n22287), .Z(n22289) );
  NAND U23095 ( .A(n22290), .B(n22289), .Z(n22534) );
  OR U23096 ( .A(n22292), .B(n22291), .Z(n22296) );
  NAND U23097 ( .A(n22294), .B(n22293), .Z(n22295) );
  NAND U23098 ( .A(n22296), .B(n22295), .Z(n22472) );
  OR U23099 ( .A(n22298), .B(n22297), .Z(n22302) );
  NANDN U23100 ( .A(n22300), .B(n22299), .Z(n22301) );
  NAND U23101 ( .A(n22302), .B(n22301), .Z(n22471) );
  OR U23102 ( .A(n22304), .B(n22303), .Z(n22308) );
  NANDN U23103 ( .A(n22306), .B(n22305), .Z(n22307) );
  NAND U23104 ( .A(n22308), .B(n22307), .Z(n22470) );
  XOR U23105 ( .A(n22472), .B(n22473), .Z(n22532) );
  OR U23106 ( .A(n22310), .B(n22309), .Z(n22314) );
  NANDN U23107 ( .A(n22312), .B(n22311), .Z(n22313) );
  NAND U23108 ( .A(n22314), .B(n22313), .Z(n22485) );
  XNOR U23109 ( .A(b[19]), .B(a[144]), .Z(n22452) );
  NANDN U23110 ( .A(n22452), .B(n37934), .Z(n22317) );
  NANDN U23111 ( .A(n22315), .B(n37935), .Z(n22316) );
  NAND U23112 ( .A(n22317), .B(n22316), .Z(n22497) );
  XOR U23113 ( .A(b[27]), .B(a[136]), .Z(n22455) );
  NAND U23114 ( .A(n38423), .B(n22455), .Z(n22320) );
  NAND U23115 ( .A(n22318), .B(n38424), .Z(n22319) );
  NAND U23116 ( .A(n22320), .B(n22319), .Z(n22494) );
  XNOR U23117 ( .A(b[5]), .B(a[158]), .Z(n22458) );
  NANDN U23118 ( .A(n22458), .B(n36587), .Z(n22323) );
  NANDN U23119 ( .A(n22321), .B(n36588), .Z(n22322) );
  AND U23120 ( .A(n22323), .B(n22322), .Z(n22495) );
  XNOR U23121 ( .A(n22494), .B(n22495), .Z(n22496) );
  XNOR U23122 ( .A(n22497), .B(n22496), .Z(n22482) );
  NANDN U23123 ( .A(n22324), .B(n37762), .Z(n22326) );
  XOR U23124 ( .A(b[17]), .B(a[146]), .Z(n22461) );
  NAND U23125 ( .A(n22461), .B(n37764), .Z(n22325) );
  NAND U23126 ( .A(n22326), .B(n22325), .Z(n22436) );
  XNOR U23127 ( .A(b[31]), .B(a[132]), .Z(n22464) );
  NANDN U23128 ( .A(n22464), .B(n38552), .Z(n22329) );
  NANDN U23129 ( .A(n22327), .B(n38553), .Z(n22328) );
  AND U23130 ( .A(n22329), .B(n22328), .Z(n22434) );
  OR U23131 ( .A(n22330), .B(n36105), .Z(n22332) );
  XNOR U23132 ( .A(b[3]), .B(a[160]), .Z(n22467) );
  NANDN U23133 ( .A(n22467), .B(n36107), .Z(n22331) );
  AND U23134 ( .A(n22332), .B(n22331), .Z(n22435) );
  XOR U23135 ( .A(n22436), .B(n22437), .Z(n22483) );
  XOR U23136 ( .A(n22482), .B(n22483), .Z(n22484) );
  XNOR U23137 ( .A(n22485), .B(n22484), .Z(n22531) );
  XOR U23138 ( .A(n22532), .B(n22531), .Z(n22533) );
  XNOR U23139 ( .A(n22534), .B(n22533), .Z(n22550) );
  OR U23140 ( .A(n22334), .B(n22333), .Z(n22338) );
  NAND U23141 ( .A(n22336), .B(n22335), .Z(n22337) );
  NAND U23142 ( .A(n22338), .B(n22337), .Z(n22548) );
  NANDN U23143 ( .A(n22340), .B(n22339), .Z(n22344) );
  NANDN U23144 ( .A(n22342), .B(n22341), .Z(n22343) );
  NAND U23145 ( .A(n22344), .B(n22343), .Z(n22538) );
  OR U23146 ( .A(n22346), .B(n22345), .Z(n22350) );
  NAND U23147 ( .A(n22348), .B(n22347), .Z(n22349) );
  NAND U23148 ( .A(n22350), .B(n22349), .Z(n22535) );
  XOR U23149 ( .A(b[9]), .B(n25862), .Z(n22500) );
  NANDN U23150 ( .A(n22500), .B(n36925), .Z(n22353) );
  NANDN U23151 ( .A(n22351), .B(n36926), .Z(n22352) );
  NAND U23152 ( .A(n22353), .B(n22352), .Z(n22442) );
  XNOR U23153 ( .A(b[15]), .B(a[148]), .Z(n22503) );
  OR U23154 ( .A(n22503), .B(n37665), .Z(n22356) );
  NANDN U23155 ( .A(n22354), .B(n37604), .Z(n22355) );
  AND U23156 ( .A(n22356), .B(n22355), .Z(n22440) );
  XOR U23157 ( .A(b[21]), .B(n24120), .Z(n22506) );
  NANDN U23158 ( .A(n22506), .B(n38101), .Z(n22359) );
  NANDN U23159 ( .A(n22357), .B(n38102), .Z(n22358) );
  AND U23160 ( .A(n22359), .B(n22358), .Z(n22441) );
  XOR U23161 ( .A(n22442), .B(n22443), .Z(n22431) );
  XOR U23162 ( .A(b[11]), .B(n25213), .Z(n22509) );
  OR U23163 ( .A(n22509), .B(n37311), .Z(n22362) );
  NANDN U23164 ( .A(n22360), .B(n37218), .Z(n22361) );
  NAND U23165 ( .A(n22362), .B(n22361), .Z(n22429) );
  XOR U23166 ( .A(n1053), .B(a[150]), .Z(n22512) );
  NANDN U23167 ( .A(n22512), .B(n37424), .Z(n22365) );
  NANDN U23168 ( .A(n22363), .B(n37425), .Z(n22364) );
  NAND U23169 ( .A(n22365), .B(n22364), .Z(n22428) );
  XOR U23170 ( .A(n22431), .B(n22430), .Z(n22425) );
  NANDN U23171 ( .A(n1049), .B(a[162]), .Z(n22366) );
  XNOR U23172 ( .A(b[1]), .B(n22366), .Z(n22368) );
  IV U23173 ( .A(a[161]), .Z(n26869) );
  NANDN U23174 ( .A(n26869), .B(n1049), .Z(n22367) );
  AND U23175 ( .A(n22368), .B(n22367), .Z(n22448) );
  NAND U23176 ( .A(n22369), .B(n38490), .Z(n22371) );
  XNOR U23177 ( .A(b[29]), .B(a[134]), .Z(n22519) );
  OR U23178 ( .A(n22519), .B(n1048), .Z(n22370) );
  NAND U23179 ( .A(n22371), .B(n22370), .Z(n22446) );
  NANDN U23180 ( .A(n1059), .B(a[130]), .Z(n22447) );
  XNOR U23181 ( .A(n22446), .B(n22447), .Z(n22449) );
  XNOR U23182 ( .A(n22448), .B(n22449), .Z(n22423) );
  NANDN U23183 ( .A(n22372), .B(n38205), .Z(n22374) );
  XNOR U23184 ( .A(b[23]), .B(a[140]), .Z(n22522) );
  OR U23185 ( .A(n22522), .B(n38268), .Z(n22373) );
  NAND U23186 ( .A(n22374), .B(n22373), .Z(n22491) );
  XOR U23187 ( .A(b[7]), .B(a[156]), .Z(n22525) );
  NAND U23188 ( .A(n22525), .B(n36701), .Z(n22377) );
  NAND U23189 ( .A(n22375), .B(n36702), .Z(n22376) );
  NAND U23190 ( .A(n22377), .B(n22376), .Z(n22488) );
  XOR U23191 ( .A(b[25]), .B(a[138]), .Z(n22528) );
  NAND U23192 ( .A(n22528), .B(n38325), .Z(n22380) );
  NANDN U23193 ( .A(n22378), .B(n38326), .Z(n22379) );
  AND U23194 ( .A(n22380), .B(n22379), .Z(n22489) );
  XNOR U23195 ( .A(n22488), .B(n22489), .Z(n22490) );
  XOR U23196 ( .A(n22491), .B(n22490), .Z(n22422) );
  XNOR U23197 ( .A(n22425), .B(n22424), .Z(n22479) );
  NANDN U23198 ( .A(n22382), .B(n22381), .Z(n22386) );
  NAND U23199 ( .A(n22384), .B(n22383), .Z(n22385) );
  NAND U23200 ( .A(n22386), .B(n22385), .Z(n22477) );
  NANDN U23201 ( .A(n22388), .B(n22387), .Z(n22392) );
  NAND U23202 ( .A(n22390), .B(n22389), .Z(n22391) );
  AND U23203 ( .A(n22392), .B(n22391), .Z(n22476) );
  XNOR U23204 ( .A(n22477), .B(n22476), .Z(n22478) );
  XNOR U23205 ( .A(n22479), .B(n22478), .Z(n22536) );
  XNOR U23206 ( .A(n22535), .B(n22536), .Z(n22537) );
  XOR U23207 ( .A(n22538), .B(n22537), .Z(n22547) );
  XNOR U23208 ( .A(n22548), .B(n22547), .Z(n22549) );
  XOR U23209 ( .A(n22550), .B(n22549), .Z(n22544) );
  NANDN U23210 ( .A(n22394), .B(n22393), .Z(n22398) );
  OR U23211 ( .A(n22396), .B(n22395), .Z(n22397) );
  NAND U23212 ( .A(n22398), .B(n22397), .Z(n22541) );
  NAND U23213 ( .A(n22400), .B(n22399), .Z(n22404) );
  NANDN U23214 ( .A(n22402), .B(n22401), .Z(n22403) );
  NAND U23215 ( .A(n22404), .B(n22403), .Z(n22542) );
  XNOR U23216 ( .A(n22541), .B(n22542), .Z(n22543) );
  XOR U23217 ( .A(n22544), .B(n22543), .Z(n22419) );
  XOR U23218 ( .A(n22418), .B(n22419), .Z(n22410) );
  XOR U23219 ( .A(n22411), .B(n22410), .Z(n22412) );
  XNOR U23220 ( .A(n22413), .B(n22412), .Z(n22553) );
  XNOR U23221 ( .A(n22553), .B(sreg[386]), .Z(n22555) );
  NAND U23222 ( .A(n22405), .B(sreg[385]), .Z(n22409) );
  OR U23223 ( .A(n22407), .B(n22406), .Z(n22408) );
  AND U23224 ( .A(n22409), .B(n22408), .Z(n22554) );
  XOR U23225 ( .A(n22555), .B(n22554), .Z(c[386]) );
  NAND U23226 ( .A(n22411), .B(n22410), .Z(n22415) );
  NAND U23227 ( .A(n22413), .B(n22412), .Z(n22414) );
  NAND U23228 ( .A(n22415), .B(n22414), .Z(n22561) );
  NANDN U23229 ( .A(n22417), .B(n22416), .Z(n22421) );
  NAND U23230 ( .A(n22419), .B(n22418), .Z(n22420) );
  NAND U23231 ( .A(n22421), .B(n22420), .Z(n22559) );
  NANDN U23232 ( .A(n22423), .B(n22422), .Z(n22427) );
  NANDN U23233 ( .A(n22425), .B(n22424), .Z(n22426) );
  NAND U23234 ( .A(n22427), .B(n22426), .Z(n22691) );
  OR U23235 ( .A(n22429), .B(n22428), .Z(n22433) );
  NAND U23236 ( .A(n22431), .B(n22430), .Z(n22432) );
  NAND U23237 ( .A(n22433), .B(n22432), .Z(n22630) );
  OR U23238 ( .A(n22435), .B(n22434), .Z(n22439) );
  NANDN U23239 ( .A(n22437), .B(n22436), .Z(n22438) );
  NAND U23240 ( .A(n22439), .B(n22438), .Z(n22629) );
  OR U23241 ( .A(n22441), .B(n22440), .Z(n22445) );
  NANDN U23242 ( .A(n22443), .B(n22442), .Z(n22444) );
  NAND U23243 ( .A(n22445), .B(n22444), .Z(n22628) );
  XOR U23244 ( .A(n22630), .B(n22631), .Z(n22688) );
  NANDN U23245 ( .A(n22447), .B(n22446), .Z(n22451) );
  NAND U23246 ( .A(n22449), .B(n22448), .Z(n22450) );
  NAND U23247 ( .A(n22451), .B(n22450), .Z(n22643) );
  XOR U23248 ( .A(b[19]), .B(n24554), .Z(n22610) );
  NANDN U23249 ( .A(n22610), .B(n37934), .Z(n22454) );
  NANDN U23250 ( .A(n22452), .B(n37935), .Z(n22453) );
  NAND U23251 ( .A(n22454), .B(n22453), .Z(n22655) );
  XNOR U23252 ( .A(b[27]), .B(a[137]), .Z(n22613) );
  NANDN U23253 ( .A(n22613), .B(n38423), .Z(n22457) );
  NAND U23254 ( .A(n22455), .B(n38424), .Z(n22456) );
  NAND U23255 ( .A(n22457), .B(n22456), .Z(n22652) );
  XNOR U23256 ( .A(b[5]), .B(a[159]), .Z(n22616) );
  NANDN U23257 ( .A(n22616), .B(n36587), .Z(n22460) );
  NANDN U23258 ( .A(n22458), .B(n36588), .Z(n22459) );
  AND U23259 ( .A(n22460), .B(n22459), .Z(n22653) );
  XNOR U23260 ( .A(n22652), .B(n22653), .Z(n22654) );
  XNOR U23261 ( .A(n22655), .B(n22654), .Z(n22640) );
  NAND U23262 ( .A(n22461), .B(n37762), .Z(n22463) );
  XOR U23263 ( .A(b[17]), .B(a[147]), .Z(n22619) );
  NAND U23264 ( .A(n22619), .B(n37764), .Z(n22462) );
  NAND U23265 ( .A(n22463), .B(n22462), .Z(n22594) );
  XNOR U23266 ( .A(b[31]), .B(a[133]), .Z(n22622) );
  NANDN U23267 ( .A(n22622), .B(n38552), .Z(n22466) );
  NANDN U23268 ( .A(n22464), .B(n38553), .Z(n22465) );
  AND U23269 ( .A(n22466), .B(n22465), .Z(n22592) );
  OR U23270 ( .A(n22467), .B(n36105), .Z(n22469) );
  XOR U23271 ( .A(b[3]), .B(n26869), .Z(n22625) );
  NANDN U23272 ( .A(n22625), .B(n36107), .Z(n22468) );
  AND U23273 ( .A(n22469), .B(n22468), .Z(n22593) );
  XOR U23274 ( .A(n22594), .B(n22595), .Z(n22641) );
  XOR U23275 ( .A(n22640), .B(n22641), .Z(n22642) );
  XNOR U23276 ( .A(n22643), .B(n22642), .Z(n22689) );
  XNOR U23277 ( .A(n22688), .B(n22689), .Z(n22690) );
  XNOR U23278 ( .A(n22691), .B(n22690), .Z(n22577) );
  OR U23279 ( .A(n22471), .B(n22470), .Z(n22475) );
  NANDN U23280 ( .A(n22473), .B(n22472), .Z(n22474) );
  NAND U23281 ( .A(n22475), .B(n22474), .Z(n22575) );
  NANDN U23282 ( .A(n22477), .B(n22476), .Z(n22481) );
  NANDN U23283 ( .A(n22479), .B(n22478), .Z(n22480) );
  NAND U23284 ( .A(n22481), .B(n22480), .Z(n22697) );
  OR U23285 ( .A(n22483), .B(n22482), .Z(n22487) );
  NANDN U23286 ( .A(n22485), .B(n22484), .Z(n22486) );
  NAND U23287 ( .A(n22487), .B(n22486), .Z(n22695) );
  NANDN U23288 ( .A(n22489), .B(n22488), .Z(n22493) );
  NAND U23289 ( .A(n22491), .B(n22490), .Z(n22492) );
  NAND U23290 ( .A(n22493), .B(n22492), .Z(n22634) );
  NANDN U23291 ( .A(n22495), .B(n22494), .Z(n22499) );
  NAND U23292 ( .A(n22497), .B(n22496), .Z(n22498) );
  AND U23293 ( .A(n22499), .B(n22498), .Z(n22635) );
  XNOR U23294 ( .A(n22634), .B(n22635), .Z(n22636) );
  XNOR U23295 ( .A(b[9]), .B(a[155]), .Z(n22658) );
  NANDN U23296 ( .A(n22658), .B(n36925), .Z(n22502) );
  NANDN U23297 ( .A(n22500), .B(n36926), .Z(n22501) );
  NAND U23298 ( .A(n22502), .B(n22501), .Z(n22600) );
  XNOR U23299 ( .A(b[15]), .B(a[149]), .Z(n22661) );
  OR U23300 ( .A(n22661), .B(n37665), .Z(n22505) );
  NANDN U23301 ( .A(n22503), .B(n37604), .Z(n22504) );
  AND U23302 ( .A(n22505), .B(n22504), .Z(n22598) );
  XNOR U23303 ( .A(b[21]), .B(a[143]), .Z(n22664) );
  NANDN U23304 ( .A(n22664), .B(n38101), .Z(n22508) );
  NANDN U23305 ( .A(n22506), .B(n38102), .Z(n22507) );
  AND U23306 ( .A(n22508), .B(n22507), .Z(n22599) );
  XOR U23307 ( .A(n22600), .B(n22601), .Z(n22589) );
  XNOR U23308 ( .A(b[11]), .B(a[153]), .Z(n22667) );
  OR U23309 ( .A(n22667), .B(n37311), .Z(n22511) );
  NANDN U23310 ( .A(n22509), .B(n37218), .Z(n22510) );
  NAND U23311 ( .A(n22511), .B(n22510), .Z(n22587) );
  XOR U23312 ( .A(n1053), .B(a[151]), .Z(n22670) );
  NANDN U23313 ( .A(n22670), .B(n37424), .Z(n22514) );
  NANDN U23314 ( .A(n22512), .B(n37425), .Z(n22513) );
  NAND U23315 ( .A(n22514), .B(n22513), .Z(n22586) );
  XOR U23316 ( .A(n22589), .B(n22588), .Z(n22583) );
  NANDN U23317 ( .A(n1049), .B(a[163]), .Z(n22515) );
  XNOR U23318 ( .A(b[1]), .B(n22515), .Z(n22517) );
  NANDN U23319 ( .A(b[0]), .B(a[162]), .Z(n22516) );
  AND U23320 ( .A(n22517), .B(n22516), .Z(n22607) );
  ANDN U23321 ( .B(b[31]), .A(n22518), .Z(n22604) );
  NANDN U23322 ( .A(n22519), .B(n38490), .Z(n22521) );
  XNOR U23323 ( .A(n1058), .B(a[135]), .Z(n22676) );
  NANDN U23324 ( .A(n1048), .B(n22676), .Z(n22520) );
  NAND U23325 ( .A(n22521), .B(n22520), .Z(n22605) );
  XOR U23326 ( .A(n22604), .B(n22605), .Z(n22606) );
  XNOR U23327 ( .A(n22607), .B(n22606), .Z(n22580) );
  NANDN U23328 ( .A(n22522), .B(n38205), .Z(n22524) );
  XOR U23329 ( .A(b[23]), .B(n23961), .Z(n22679) );
  OR U23330 ( .A(n22679), .B(n38268), .Z(n22523) );
  NAND U23331 ( .A(n22524), .B(n22523), .Z(n22649) );
  XOR U23332 ( .A(b[7]), .B(a[157]), .Z(n22682) );
  NAND U23333 ( .A(n22682), .B(n36701), .Z(n22527) );
  NAND U23334 ( .A(n22525), .B(n36702), .Z(n22526) );
  NAND U23335 ( .A(n22527), .B(n22526), .Z(n22646) );
  XNOR U23336 ( .A(b[25]), .B(a[139]), .Z(n22685) );
  NANDN U23337 ( .A(n22685), .B(n38325), .Z(n22530) );
  NAND U23338 ( .A(n22528), .B(n38326), .Z(n22529) );
  AND U23339 ( .A(n22530), .B(n22529), .Z(n22647) );
  XNOR U23340 ( .A(n22646), .B(n22647), .Z(n22648) );
  XNOR U23341 ( .A(n22649), .B(n22648), .Z(n22581) );
  XOR U23342 ( .A(n22583), .B(n22582), .Z(n22637) );
  XNOR U23343 ( .A(n22636), .B(n22637), .Z(n22694) );
  XOR U23344 ( .A(n22695), .B(n22694), .Z(n22696) );
  XNOR U23345 ( .A(n22697), .B(n22696), .Z(n22574) );
  XNOR U23346 ( .A(n22575), .B(n22574), .Z(n22576) );
  XOR U23347 ( .A(n22577), .B(n22576), .Z(n22571) );
  NANDN U23348 ( .A(n22536), .B(n22535), .Z(n22540) );
  NAND U23349 ( .A(n22538), .B(n22537), .Z(n22539) );
  AND U23350 ( .A(n22540), .B(n22539), .Z(n22568) );
  XNOR U23351 ( .A(n22569), .B(n22568), .Z(n22570) );
  XNOR U23352 ( .A(n22571), .B(n22570), .Z(n22565) );
  NANDN U23353 ( .A(n22542), .B(n22541), .Z(n22546) );
  NAND U23354 ( .A(n22544), .B(n22543), .Z(n22545) );
  NAND U23355 ( .A(n22546), .B(n22545), .Z(n22562) );
  NANDN U23356 ( .A(n22548), .B(n22547), .Z(n22552) );
  NANDN U23357 ( .A(n22550), .B(n22549), .Z(n22551) );
  NAND U23358 ( .A(n22552), .B(n22551), .Z(n22563) );
  XNOR U23359 ( .A(n22562), .B(n22563), .Z(n22564) );
  XNOR U23360 ( .A(n22565), .B(n22564), .Z(n22558) );
  XOR U23361 ( .A(n22559), .B(n22558), .Z(n22560) );
  XNOR U23362 ( .A(n22561), .B(n22560), .Z(n22700) );
  XNOR U23363 ( .A(n22700), .B(sreg[387]), .Z(n22702) );
  NAND U23364 ( .A(n22553), .B(sreg[386]), .Z(n22557) );
  OR U23365 ( .A(n22555), .B(n22554), .Z(n22556) );
  AND U23366 ( .A(n22557), .B(n22556), .Z(n22701) );
  XOR U23367 ( .A(n22702), .B(n22701), .Z(c[387]) );
  NANDN U23368 ( .A(n22563), .B(n22562), .Z(n22567) );
  NANDN U23369 ( .A(n22565), .B(n22564), .Z(n22566) );
  NAND U23370 ( .A(n22567), .B(n22566), .Z(n22706) );
  NANDN U23371 ( .A(n22569), .B(n22568), .Z(n22573) );
  NAND U23372 ( .A(n22571), .B(n22570), .Z(n22572) );
  NAND U23373 ( .A(n22573), .B(n22572), .Z(n22711) );
  NANDN U23374 ( .A(n22575), .B(n22574), .Z(n22579) );
  NANDN U23375 ( .A(n22577), .B(n22576), .Z(n22578) );
  NAND U23376 ( .A(n22579), .B(n22578), .Z(n22712) );
  XNOR U23377 ( .A(n22711), .B(n22712), .Z(n22713) );
  OR U23378 ( .A(n22581), .B(n22580), .Z(n22585) );
  NANDN U23379 ( .A(n22583), .B(n22582), .Z(n22584) );
  NAND U23380 ( .A(n22585), .B(n22584), .Z(n22840) );
  OR U23381 ( .A(n22587), .B(n22586), .Z(n22591) );
  NAND U23382 ( .A(n22589), .B(n22588), .Z(n22590) );
  NAND U23383 ( .A(n22591), .B(n22590), .Z(n22779) );
  OR U23384 ( .A(n22593), .B(n22592), .Z(n22597) );
  NANDN U23385 ( .A(n22595), .B(n22594), .Z(n22596) );
  NAND U23386 ( .A(n22597), .B(n22596), .Z(n22778) );
  OR U23387 ( .A(n22599), .B(n22598), .Z(n22603) );
  NANDN U23388 ( .A(n22601), .B(n22600), .Z(n22602) );
  NAND U23389 ( .A(n22603), .B(n22602), .Z(n22777) );
  XOR U23390 ( .A(n22779), .B(n22780), .Z(n22838) );
  OR U23391 ( .A(n22605), .B(n22604), .Z(n22609) );
  NANDN U23392 ( .A(n22607), .B(n22606), .Z(n22608) );
  NAND U23393 ( .A(n22609), .B(n22608), .Z(n22791) );
  XNOR U23394 ( .A(b[19]), .B(a[146]), .Z(n22735) );
  NANDN U23395 ( .A(n22735), .B(n37934), .Z(n22612) );
  NANDN U23396 ( .A(n22610), .B(n37935), .Z(n22611) );
  NAND U23397 ( .A(n22612), .B(n22611), .Z(n22804) );
  XOR U23398 ( .A(b[27]), .B(a[138]), .Z(n22738) );
  NAND U23399 ( .A(n38423), .B(n22738), .Z(n22615) );
  NANDN U23400 ( .A(n22613), .B(n38424), .Z(n22614) );
  NAND U23401 ( .A(n22615), .B(n22614), .Z(n22801) );
  XNOR U23402 ( .A(b[5]), .B(a[160]), .Z(n22741) );
  NANDN U23403 ( .A(n22741), .B(n36587), .Z(n22618) );
  NANDN U23404 ( .A(n22616), .B(n36588), .Z(n22617) );
  AND U23405 ( .A(n22618), .B(n22617), .Z(n22802) );
  XNOR U23406 ( .A(n22801), .B(n22802), .Z(n22803) );
  XNOR U23407 ( .A(n22804), .B(n22803), .Z(n22790) );
  NAND U23408 ( .A(n22619), .B(n37762), .Z(n22621) );
  XOR U23409 ( .A(b[17]), .B(a[148]), .Z(n22744) );
  NAND U23410 ( .A(n22744), .B(n37764), .Z(n22620) );
  NAND U23411 ( .A(n22621), .B(n22620), .Z(n22762) );
  XNOR U23412 ( .A(b[31]), .B(a[134]), .Z(n22747) );
  NANDN U23413 ( .A(n22747), .B(n38552), .Z(n22624) );
  NANDN U23414 ( .A(n22622), .B(n38553), .Z(n22623) );
  NAND U23415 ( .A(n22624), .B(n22623), .Z(n22759) );
  OR U23416 ( .A(n22625), .B(n36105), .Z(n22627) );
  XNOR U23417 ( .A(b[3]), .B(a[162]), .Z(n22750) );
  NANDN U23418 ( .A(n22750), .B(n36107), .Z(n22626) );
  AND U23419 ( .A(n22627), .B(n22626), .Z(n22760) );
  XNOR U23420 ( .A(n22759), .B(n22760), .Z(n22761) );
  XOR U23421 ( .A(n22762), .B(n22761), .Z(n22789) );
  XOR U23422 ( .A(n22790), .B(n22789), .Z(n22792) );
  XOR U23423 ( .A(n22791), .B(n22792), .Z(n22837) );
  XOR U23424 ( .A(n22838), .B(n22837), .Z(n22839) );
  XNOR U23425 ( .A(n22840), .B(n22839), .Z(n22726) );
  OR U23426 ( .A(n22629), .B(n22628), .Z(n22633) );
  NANDN U23427 ( .A(n22631), .B(n22630), .Z(n22632) );
  NAND U23428 ( .A(n22633), .B(n22632), .Z(n22724) );
  NANDN U23429 ( .A(n22635), .B(n22634), .Z(n22639) );
  NANDN U23430 ( .A(n22637), .B(n22636), .Z(n22638) );
  NAND U23431 ( .A(n22639), .B(n22638), .Z(n22845) );
  OR U23432 ( .A(n22641), .B(n22640), .Z(n22645) );
  NAND U23433 ( .A(n22643), .B(n22642), .Z(n22644) );
  NAND U23434 ( .A(n22645), .B(n22644), .Z(n22844) );
  NANDN U23435 ( .A(n22647), .B(n22646), .Z(n22651) );
  NAND U23436 ( .A(n22649), .B(n22648), .Z(n22650) );
  NAND U23437 ( .A(n22651), .B(n22650), .Z(n22783) );
  NANDN U23438 ( .A(n22653), .B(n22652), .Z(n22657) );
  NAND U23439 ( .A(n22655), .B(n22654), .Z(n22656) );
  AND U23440 ( .A(n22657), .B(n22656), .Z(n22784) );
  XNOR U23441 ( .A(n22783), .B(n22784), .Z(n22785) );
  XNOR U23442 ( .A(n1052), .B(a[156]), .Z(n22807) );
  NAND U23443 ( .A(n36925), .B(n22807), .Z(n22660) );
  NANDN U23444 ( .A(n22658), .B(n36926), .Z(n22659) );
  NAND U23445 ( .A(n22660), .B(n22659), .Z(n22767) );
  XNOR U23446 ( .A(b[15]), .B(a[150]), .Z(n22810) );
  OR U23447 ( .A(n22810), .B(n37665), .Z(n22663) );
  NANDN U23448 ( .A(n22661), .B(n37604), .Z(n22662) );
  AND U23449 ( .A(n22663), .B(n22662), .Z(n22765) );
  XNOR U23450 ( .A(n1056), .B(a[144]), .Z(n22813) );
  NAND U23451 ( .A(n22813), .B(n38101), .Z(n22666) );
  NANDN U23452 ( .A(n22664), .B(n38102), .Z(n22665) );
  AND U23453 ( .A(n22666), .B(n22665), .Z(n22766) );
  XOR U23454 ( .A(n22767), .B(n22768), .Z(n22756) );
  XOR U23455 ( .A(b[11]), .B(n25862), .Z(n22816) );
  OR U23456 ( .A(n22816), .B(n37311), .Z(n22669) );
  NANDN U23457 ( .A(n22667), .B(n37218), .Z(n22668) );
  NAND U23458 ( .A(n22669), .B(n22668), .Z(n22754) );
  XOR U23459 ( .A(n1053), .B(a[152]), .Z(n22819) );
  NANDN U23460 ( .A(n22819), .B(n37424), .Z(n22672) );
  NANDN U23461 ( .A(n22670), .B(n37425), .Z(n22671) );
  AND U23462 ( .A(n22672), .B(n22671), .Z(n22753) );
  XNOR U23463 ( .A(n22754), .B(n22753), .Z(n22755) );
  XOR U23464 ( .A(n22756), .B(n22755), .Z(n22773) );
  NANDN U23465 ( .A(n1049), .B(a[164]), .Z(n22673) );
  XNOR U23466 ( .A(b[1]), .B(n22673), .Z(n22675) );
  IV U23467 ( .A(a[163]), .Z(n27178) );
  NANDN U23468 ( .A(n27178), .B(n1049), .Z(n22674) );
  AND U23469 ( .A(n22675), .B(n22674), .Z(n22731) );
  NAND U23470 ( .A(n22676), .B(n38490), .Z(n22678) );
  XNOR U23471 ( .A(n1058), .B(a[136]), .Z(n22825) );
  NANDN U23472 ( .A(n1048), .B(n22825), .Z(n22677) );
  NAND U23473 ( .A(n22678), .B(n22677), .Z(n22729) );
  NANDN U23474 ( .A(n1059), .B(a[132]), .Z(n22730) );
  XNOR U23475 ( .A(n22729), .B(n22730), .Z(n22732) );
  XOR U23476 ( .A(n22731), .B(n22732), .Z(n22771) );
  NANDN U23477 ( .A(n22679), .B(n38205), .Z(n22681) );
  XOR U23478 ( .A(b[23]), .B(n24120), .Z(n22828) );
  OR U23479 ( .A(n22828), .B(n38268), .Z(n22680) );
  NAND U23480 ( .A(n22681), .B(n22680), .Z(n22798) );
  XOR U23481 ( .A(b[7]), .B(a[158]), .Z(n22831) );
  NAND U23482 ( .A(n22831), .B(n36701), .Z(n22684) );
  NAND U23483 ( .A(n22682), .B(n36702), .Z(n22683) );
  NAND U23484 ( .A(n22684), .B(n22683), .Z(n22795) );
  XOR U23485 ( .A(b[25]), .B(a[140]), .Z(n22834) );
  NAND U23486 ( .A(n22834), .B(n38325), .Z(n22687) );
  NANDN U23487 ( .A(n22685), .B(n38326), .Z(n22686) );
  AND U23488 ( .A(n22687), .B(n22686), .Z(n22796) );
  XNOR U23489 ( .A(n22795), .B(n22796), .Z(n22797) );
  XNOR U23490 ( .A(n22798), .B(n22797), .Z(n22772) );
  XOR U23491 ( .A(n22771), .B(n22772), .Z(n22774) );
  XNOR U23492 ( .A(n22773), .B(n22774), .Z(n22786) );
  XNOR U23493 ( .A(n22785), .B(n22786), .Z(n22843) );
  XNOR U23494 ( .A(n22844), .B(n22843), .Z(n22846) );
  XNOR U23495 ( .A(n22845), .B(n22846), .Z(n22723) );
  XNOR U23496 ( .A(n22724), .B(n22723), .Z(n22725) );
  XOR U23497 ( .A(n22726), .B(n22725), .Z(n22720) );
  NANDN U23498 ( .A(n22689), .B(n22688), .Z(n22693) );
  NAND U23499 ( .A(n22691), .B(n22690), .Z(n22692) );
  NAND U23500 ( .A(n22693), .B(n22692), .Z(n22718) );
  NAND U23501 ( .A(n22695), .B(n22694), .Z(n22699) );
  NANDN U23502 ( .A(n22697), .B(n22696), .Z(n22698) );
  AND U23503 ( .A(n22699), .B(n22698), .Z(n22717) );
  XNOR U23504 ( .A(n22718), .B(n22717), .Z(n22719) );
  XOR U23505 ( .A(n22720), .B(n22719), .Z(n22714) );
  XOR U23506 ( .A(n22713), .B(n22714), .Z(n22705) );
  XOR U23507 ( .A(n22706), .B(n22705), .Z(n22707) );
  XNOR U23508 ( .A(n22708), .B(n22707), .Z(n22849) );
  XNOR U23509 ( .A(n22849), .B(sreg[388]), .Z(n22851) );
  NAND U23510 ( .A(n22700), .B(sreg[387]), .Z(n22704) );
  OR U23511 ( .A(n22702), .B(n22701), .Z(n22703) );
  AND U23512 ( .A(n22704), .B(n22703), .Z(n22850) );
  XOR U23513 ( .A(n22851), .B(n22850), .Z(c[388]) );
  NAND U23514 ( .A(n22706), .B(n22705), .Z(n22710) );
  NAND U23515 ( .A(n22708), .B(n22707), .Z(n22709) );
  NAND U23516 ( .A(n22710), .B(n22709), .Z(n22857) );
  NANDN U23517 ( .A(n22712), .B(n22711), .Z(n22716) );
  NAND U23518 ( .A(n22714), .B(n22713), .Z(n22715) );
  NAND U23519 ( .A(n22716), .B(n22715), .Z(n22855) );
  NANDN U23520 ( .A(n22718), .B(n22717), .Z(n22722) );
  NAND U23521 ( .A(n22720), .B(n22719), .Z(n22721) );
  NAND U23522 ( .A(n22722), .B(n22721), .Z(n22860) );
  NANDN U23523 ( .A(n22724), .B(n22723), .Z(n22728) );
  NANDN U23524 ( .A(n22726), .B(n22725), .Z(n22727) );
  NAND U23525 ( .A(n22728), .B(n22727), .Z(n22861) );
  XNOR U23526 ( .A(n22860), .B(n22861), .Z(n22862) );
  NANDN U23527 ( .A(n22730), .B(n22729), .Z(n22734) );
  NAND U23528 ( .A(n22732), .B(n22731), .Z(n22733) );
  NAND U23529 ( .A(n22734), .B(n22733), .Z(n22939) );
  XNOR U23530 ( .A(b[19]), .B(a[147]), .Z(n22884) );
  NANDN U23531 ( .A(n22884), .B(n37934), .Z(n22737) );
  NANDN U23532 ( .A(n22735), .B(n37935), .Z(n22736) );
  NAND U23533 ( .A(n22737), .B(n22736), .Z(n22949) );
  XNOR U23534 ( .A(b[27]), .B(a[139]), .Z(n22887) );
  NANDN U23535 ( .A(n22887), .B(n38423), .Z(n22740) );
  NAND U23536 ( .A(n22738), .B(n38424), .Z(n22739) );
  NAND U23537 ( .A(n22740), .B(n22739), .Z(n22946) );
  XOR U23538 ( .A(b[5]), .B(n26869), .Z(n22890) );
  NANDN U23539 ( .A(n22890), .B(n36587), .Z(n22743) );
  NANDN U23540 ( .A(n22741), .B(n36588), .Z(n22742) );
  AND U23541 ( .A(n22743), .B(n22742), .Z(n22947) );
  XNOR U23542 ( .A(n22946), .B(n22947), .Z(n22948) );
  XNOR U23543 ( .A(n22949), .B(n22948), .Z(n22937) );
  NAND U23544 ( .A(n22744), .B(n37762), .Z(n22746) );
  XOR U23545 ( .A(b[17]), .B(a[149]), .Z(n22893) );
  NAND U23546 ( .A(n22893), .B(n37764), .Z(n22745) );
  NAND U23547 ( .A(n22746), .B(n22745), .Z(n22911) );
  XNOR U23548 ( .A(b[31]), .B(a[135]), .Z(n22896) );
  NANDN U23549 ( .A(n22896), .B(n38552), .Z(n22749) );
  NANDN U23550 ( .A(n22747), .B(n38553), .Z(n22748) );
  NAND U23551 ( .A(n22749), .B(n22748), .Z(n22908) );
  OR U23552 ( .A(n22750), .B(n36105), .Z(n22752) );
  XOR U23553 ( .A(b[3]), .B(n27178), .Z(n22899) );
  NANDN U23554 ( .A(n22899), .B(n36107), .Z(n22751) );
  AND U23555 ( .A(n22752), .B(n22751), .Z(n22909) );
  XNOR U23556 ( .A(n22908), .B(n22909), .Z(n22910) );
  XOR U23557 ( .A(n22911), .B(n22910), .Z(n22936) );
  XNOR U23558 ( .A(n22937), .B(n22936), .Z(n22938) );
  XNOR U23559 ( .A(n22939), .B(n22938), .Z(n22982) );
  NANDN U23560 ( .A(n22754), .B(n22753), .Z(n22758) );
  NAND U23561 ( .A(n22756), .B(n22755), .Z(n22757) );
  NAND U23562 ( .A(n22758), .B(n22757), .Z(n22927) );
  NANDN U23563 ( .A(n22760), .B(n22759), .Z(n22764) );
  NAND U23564 ( .A(n22762), .B(n22761), .Z(n22763) );
  NAND U23565 ( .A(n22764), .B(n22763), .Z(n22925) );
  OR U23566 ( .A(n22766), .B(n22765), .Z(n22770) );
  NANDN U23567 ( .A(n22768), .B(n22767), .Z(n22769) );
  NAND U23568 ( .A(n22770), .B(n22769), .Z(n22924) );
  XNOR U23569 ( .A(n22927), .B(n22926), .Z(n22983) );
  XOR U23570 ( .A(n22982), .B(n22983), .Z(n22985) );
  NANDN U23571 ( .A(n22772), .B(n22771), .Z(n22776) );
  OR U23572 ( .A(n22774), .B(n22773), .Z(n22775) );
  NAND U23573 ( .A(n22776), .B(n22775), .Z(n22984) );
  XOR U23574 ( .A(n22985), .B(n22984), .Z(n22874) );
  OR U23575 ( .A(n22778), .B(n22777), .Z(n22782) );
  NANDN U23576 ( .A(n22780), .B(n22779), .Z(n22781) );
  NAND U23577 ( .A(n22782), .B(n22781), .Z(n22873) );
  NANDN U23578 ( .A(n22784), .B(n22783), .Z(n22788) );
  NANDN U23579 ( .A(n22786), .B(n22785), .Z(n22787) );
  NAND U23580 ( .A(n22788), .B(n22787), .Z(n22990) );
  NANDN U23581 ( .A(n22790), .B(n22789), .Z(n22794) );
  OR U23582 ( .A(n22792), .B(n22791), .Z(n22793) );
  NAND U23583 ( .A(n22794), .B(n22793), .Z(n22989) );
  NANDN U23584 ( .A(n22796), .B(n22795), .Z(n22800) );
  NAND U23585 ( .A(n22798), .B(n22797), .Z(n22799) );
  NAND U23586 ( .A(n22800), .B(n22799), .Z(n22930) );
  NANDN U23587 ( .A(n22802), .B(n22801), .Z(n22806) );
  NAND U23588 ( .A(n22804), .B(n22803), .Z(n22805) );
  AND U23589 ( .A(n22806), .B(n22805), .Z(n22931) );
  XNOR U23590 ( .A(n22930), .B(n22931), .Z(n22932) );
  XOR U23591 ( .A(n1052), .B(a[157]), .Z(n22958) );
  NANDN U23592 ( .A(n22958), .B(n36925), .Z(n22809) );
  NAND U23593 ( .A(n36926), .B(n22807), .Z(n22808) );
  NAND U23594 ( .A(n22809), .B(n22808), .Z(n22916) );
  XNOR U23595 ( .A(n1054), .B(a[151]), .Z(n22955) );
  NANDN U23596 ( .A(n37665), .B(n22955), .Z(n22812) );
  NANDN U23597 ( .A(n22810), .B(n37604), .Z(n22811) );
  NAND U23598 ( .A(n22812), .B(n22811), .Z(n22914) );
  XOR U23599 ( .A(n1056), .B(a[145]), .Z(n22952) );
  NANDN U23600 ( .A(n22952), .B(n38101), .Z(n22815) );
  NAND U23601 ( .A(n38102), .B(n22813), .Z(n22814) );
  NAND U23602 ( .A(n22815), .B(n22814), .Z(n22915) );
  XNOR U23603 ( .A(n22914), .B(n22915), .Z(n22917) );
  XOR U23604 ( .A(n22916), .B(n22917), .Z(n22905) );
  XNOR U23605 ( .A(b[11]), .B(a[155]), .Z(n22961) );
  OR U23606 ( .A(n22961), .B(n37311), .Z(n22818) );
  NANDN U23607 ( .A(n22816), .B(n37218), .Z(n22817) );
  NAND U23608 ( .A(n22818), .B(n22817), .Z(n22903) );
  XOR U23609 ( .A(n1053), .B(a[153]), .Z(n22964) );
  NANDN U23610 ( .A(n22964), .B(n37424), .Z(n22821) );
  NANDN U23611 ( .A(n22819), .B(n37425), .Z(n22820) );
  AND U23612 ( .A(n22821), .B(n22820), .Z(n22902) );
  XNOR U23613 ( .A(n22903), .B(n22902), .Z(n22904) );
  XNOR U23614 ( .A(n22905), .B(n22904), .Z(n22921) );
  NANDN U23615 ( .A(n1049), .B(a[165]), .Z(n22822) );
  XNOR U23616 ( .A(b[1]), .B(n22822), .Z(n22824) );
  NANDN U23617 ( .A(b[0]), .B(a[164]), .Z(n22823) );
  AND U23618 ( .A(n22824), .B(n22823), .Z(n22880) );
  NAND U23619 ( .A(n38490), .B(n22825), .Z(n22827) );
  XOR U23620 ( .A(n1058), .B(n23393), .Z(n22967) );
  NANDN U23621 ( .A(n1048), .B(n22967), .Z(n22826) );
  NAND U23622 ( .A(n22827), .B(n22826), .Z(n22878) );
  NANDN U23623 ( .A(n1059), .B(a[133]), .Z(n22879) );
  XNOR U23624 ( .A(n22878), .B(n22879), .Z(n22881) );
  XNOR U23625 ( .A(n22880), .B(n22881), .Z(n22919) );
  NANDN U23626 ( .A(n22828), .B(n38205), .Z(n22830) );
  XNOR U23627 ( .A(b[23]), .B(a[143]), .Z(n22973) );
  OR U23628 ( .A(n22973), .B(n38268), .Z(n22829) );
  NAND U23629 ( .A(n22830), .B(n22829), .Z(n22943) );
  XOR U23630 ( .A(b[7]), .B(a[159]), .Z(n22976) );
  NAND U23631 ( .A(n22976), .B(n36701), .Z(n22833) );
  NAND U23632 ( .A(n22831), .B(n36702), .Z(n22832) );
  NAND U23633 ( .A(n22833), .B(n22832), .Z(n22940) );
  XNOR U23634 ( .A(b[25]), .B(a[141]), .Z(n22979) );
  NANDN U23635 ( .A(n22979), .B(n38325), .Z(n22836) );
  NAND U23636 ( .A(n22834), .B(n38326), .Z(n22835) );
  AND U23637 ( .A(n22836), .B(n22835), .Z(n22941) );
  XNOR U23638 ( .A(n22940), .B(n22941), .Z(n22942) );
  XOR U23639 ( .A(n22943), .B(n22942), .Z(n22918) );
  XOR U23640 ( .A(n22921), .B(n22920), .Z(n22933) );
  XOR U23641 ( .A(n22932), .B(n22933), .Z(n22988) );
  XNOR U23642 ( .A(n22989), .B(n22988), .Z(n22991) );
  XNOR U23643 ( .A(n22990), .B(n22991), .Z(n22872) );
  XOR U23644 ( .A(n22873), .B(n22872), .Z(n22875) );
  NAND U23645 ( .A(n22838), .B(n22837), .Z(n22842) );
  NAND U23646 ( .A(n22840), .B(n22839), .Z(n22841) );
  NAND U23647 ( .A(n22842), .B(n22841), .Z(n22867) );
  NAND U23648 ( .A(n22844), .B(n22843), .Z(n22848) );
  NANDN U23649 ( .A(n22846), .B(n22845), .Z(n22847) );
  AND U23650 ( .A(n22848), .B(n22847), .Z(n22866) );
  XNOR U23651 ( .A(n22867), .B(n22866), .Z(n22868) );
  XOR U23652 ( .A(n22869), .B(n22868), .Z(n22863) );
  XOR U23653 ( .A(n22862), .B(n22863), .Z(n22854) );
  XOR U23654 ( .A(n22855), .B(n22854), .Z(n22856) );
  XNOR U23655 ( .A(n22857), .B(n22856), .Z(n22994) );
  XNOR U23656 ( .A(n22994), .B(sreg[389]), .Z(n22996) );
  NAND U23657 ( .A(n22849), .B(sreg[388]), .Z(n22853) );
  OR U23658 ( .A(n22851), .B(n22850), .Z(n22852) );
  AND U23659 ( .A(n22853), .B(n22852), .Z(n22995) );
  XOR U23660 ( .A(n22996), .B(n22995), .Z(c[389]) );
  NAND U23661 ( .A(n22855), .B(n22854), .Z(n22859) );
  NAND U23662 ( .A(n22857), .B(n22856), .Z(n22858) );
  NAND U23663 ( .A(n22859), .B(n22858), .Z(n23002) );
  NANDN U23664 ( .A(n22861), .B(n22860), .Z(n22865) );
  NAND U23665 ( .A(n22863), .B(n22862), .Z(n22864) );
  NAND U23666 ( .A(n22865), .B(n22864), .Z(n23000) );
  NANDN U23667 ( .A(n22867), .B(n22866), .Z(n22871) );
  NAND U23668 ( .A(n22869), .B(n22868), .Z(n22870) );
  NAND U23669 ( .A(n22871), .B(n22870), .Z(n23005) );
  NANDN U23670 ( .A(n22873), .B(n22872), .Z(n22877) );
  OR U23671 ( .A(n22875), .B(n22874), .Z(n22876) );
  NAND U23672 ( .A(n22877), .B(n22876), .Z(n23006) );
  XNOR U23673 ( .A(n23005), .B(n23006), .Z(n23007) );
  NANDN U23674 ( .A(n22879), .B(n22878), .Z(n22883) );
  NAND U23675 ( .A(n22881), .B(n22880), .Z(n22882) );
  NAND U23676 ( .A(n22883), .B(n22882), .Z(n23080) );
  XNOR U23677 ( .A(b[19]), .B(a[148]), .Z(n23027) );
  NANDN U23678 ( .A(n23027), .B(n37934), .Z(n22886) );
  NANDN U23679 ( .A(n22884), .B(n37935), .Z(n22885) );
  NAND U23680 ( .A(n22886), .B(n22885), .Z(n23090) );
  XOR U23681 ( .A(b[27]), .B(a[140]), .Z(n23030) );
  NAND U23682 ( .A(n38423), .B(n23030), .Z(n22889) );
  NANDN U23683 ( .A(n22887), .B(n38424), .Z(n22888) );
  NAND U23684 ( .A(n22889), .B(n22888), .Z(n23087) );
  XNOR U23685 ( .A(b[5]), .B(a[162]), .Z(n23033) );
  NANDN U23686 ( .A(n23033), .B(n36587), .Z(n22892) );
  NANDN U23687 ( .A(n22890), .B(n36588), .Z(n22891) );
  AND U23688 ( .A(n22892), .B(n22891), .Z(n23088) );
  XNOR U23689 ( .A(n23087), .B(n23088), .Z(n23089) );
  XNOR U23690 ( .A(n23090), .B(n23089), .Z(n23078) );
  NAND U23691 ( .A(n22893), .B(n37762), .Z(n22895) );
  XOR U23692 ( .A(b[17]), .B(a[150]), .Z(n23036) );
  NAND U23693 ( .A(n23036), .B(n37764), .Z(n22894) );
  NAND U23694 ( .A(n22895), .B(n22894), .Z(n23054) );
  XNOR U23695 ( .A(b[31]), .B(a[136]), .Z(n23039) );
  NANDN U23696 ( .A(n23039), .B(n38552), .Z(n22898) );
  NANDN U23697 ( .A(n22896), .B(n38553), .Z(n22897) );
  NAND U23698 ( .A(n22898), .B(n22897), .Z(n23051) );
  OR U23699 ( .A(n22899), .B(n36105), .Z(n22901) );
  XNOR U23700 ( .A(b[3]), .B(a[164]), .Z(n23042) );
  NANDN U23701 ( .A(n23042), .B(n36107), .Z(n22900) );
  AND U23702 ( .A(n22901), .B(n22900), .Z(n23052) );
  XNOR U23703 ( .A(n23051), .B(n23052), .Z(n23053) );
  XOR U23704 ( .A(n23054), .B(n23053), .Z(n23077) );
  XNOR U23705 ( .A(n23078), .B(n23077), .Z(n23079) );
  XNOR U23706 ( .A(n23080), .B(n23079), .Z(n23018) );
  NANDN U23707 ( .A(n22903), .B(n22902), .Z(n22907) );
  NAND U23708 ( .A(n22905), .B(n22904), .Z(n22906) );
  NAND U23709 ( .A(n22907), .B(n22906), .Z(n23069) );
  NANDN U23710 ( .A(n22909), .B(n22908), .Z(n22913) );
  NAND U23711 ( .A(n22911), .B(n22910), .Z(n22912) );
  NAND U23712 ( .A(n22913), .B(n22912), .Z(n23068) );
  XNOR U23713 ( .A(n23068), .B(n23067), .Z(n23070) );
  XOR U23714 ( .A(n23069), .B(n23070), .Z(n23017) );
  XOR U23715 ( .A(n23018), .B(n23017), .Z(n23019) );
  NANDN U23716 ( .A(n22919), .B(n22918), .Z(n22923) );
  NAND U23717 ( .A(n22921), .B(n22920), .Z(n22922) );
  NAND U23718 ( .A(n22923), .B(n22922), .Z(n23020) );
  XNOR U23719 ( .A(n23019), .B(n23020), .Z(n23131) );
  OR U23720 ( .A(n22925), .B(n22924), .Z(n22929) );
  NAND U23721 ( .A(n22927), .B(n22926), .Z(n22928) );
  NAND U23722 ( .A(n22929), .B(n22928), .Z(n23130) );
  NANDN U23723 ( .A(n22931), .B(n22930), .Z(n22935) );
  NAND U23724 ( .A(n22933), .B(n22932), .Z(n22934) );
  NAND U23725 ( .A(n22935), .B(n22934), .Z(n23013) );
  NANDN U23726 ( .A(n22941), .B(n22940), .Z(n22945) );
  NAND U23727 ( .A(n22943), .B(n22942), .Z(n22944) );
  NAND U23728 ( .A(n22945), .B(n22944), .Z(n23071) );
  NANDN U23729 ( .A(n22947), .B(n22946), .Z(n22951) );
  NAND U23730 ( .A(n22949), .B(n22948), .Z(n22950) );
  AND U23731 ( .A(n22951), .B(n22950), .Z(n23072) );
  XNOR U23732 ( .A(n23071), .B(n23072), .Z(n23073) );
  XOR U23733 ( .A(n1056), .B(a[146]), .Z(n23099) );
  NANDN U23734 ( .A(n23099), .B(n38101), .Z(n22954) );
  NANDN U23735 ( .A(n22952), .B(n38102), .Z(n22953) );
  NAND U23736 ( .A(n22954), .B(n22953), .Z(n23063) );
  XOR U23737 ( .A(b[15]), .B(n25213), .Z(n23096) );
  OR U23738 ( .A(n23096), .B(n37665), .Z(n22957) );
  NAND U23739 ( .A(n22955), .B(n37604), .Z(n22956) );
  AND U23740 ( .A(n22957), .B(n22956), .Z(n23064) );
  XNOR U23741 ( .A(n23063), .B(n23064), .Z(n23066) );
  XOR U23742 ( .A(n1052), .B(a[158]), .Z(n23093) );
  NANDN U23743 ( .A(n23093), .B(n36925), .Z(n22960) );
  NANDN U23744 ( .A(n22958), .B(n36926), .Z(n22959) );
  NAND U23745 ( .A(n22960), .B(n22959), .Z(n23065) );
  XNOR U23746 ( .A(n23066), .B(n23065), .Z(n23059) );
  XNOR U23747 ( .A(b[11]), .B(a[156]), .Z(n23102) );
  OR U23748 ( .A(n23102), .B(n37311), .Z(n22963) );
  NANDN U23749 ( .A(n22961), .B(n37218), .Z(n22962) );
  NAND U23750 ( .A(n22963), .B(n22962), .Z(n23058) );
  XOR U23751 ( .A(n1053), .B(a[154]), .Z(n23105) );
  NANDN U23752 ( .A(n23105), .B(n37424), .Z(n22966) );
  NANDN U23753 ( .A(n22964), .B(n37425), .Z(n22965) );
  NAND U23754 ( .A(n22966), .B(n22965), .Z(n23057) );
  XNOR U23755 ( .A(n23058), .B(n23057), .Z(n23060) );
  XNOR U23756 ( .A(n23059), .B(n23060), .Z(n23048) );
  NAND U23757 ( .A(n38490), .B(n22967), .Z(n22969) );
  XNOR U23758 ( .A(n1058), .B(a[138]), .Z(n23111) );
  NANDN U23759 ( .A(n1048), .B(n23111), .Z(n22968) );
  NAND U23760 ( .A(n22969), .B(n22968), .Z(n23021) );
  NANDN U23761 ( .A(n1059), .B(a[134]), .Z(n23022) );
  XNOR U23762 ( .A(n23021), .B(n23022), .Z(n23024) );
  NANDN U23763 ( .A(n1049), .B(a[166]), .Z(n22970) );
  XNOR U23764 ( .A(b[1]), .B(n22970), .Z(n22972) );
  NANDN U23765 ( .A(b[0]), .B(a[165]), .Z(n22971) );
  AND U23766 ( .A(n22972), .B(n22971), .Z(n23023) );
  XNOR U23767 ( .A(n23024), .B(n23023), .Z(n23046) );
  NANDN U23768 ( .A(n22973), .B(n38205), .Z(n22975) );
  XNOR U23769 ( .A(b[23]), .B(a[144]), .Z(n23114) );
  OR U23770 ( .A(n23114), .B(n38268), .Z(n22974) );
  NAND U23771 ( .A(n22975), .B(n22974), .Z(n23084) );
  XOR U23772 ( .A(b[7]), .B(a[160]), .Z(n23117) );
  NAND U23773 ( .A(n23117), .B(n36701), .Z(n22978) );
  NAND U23774 ( .A(n22976), .B(n36702), .Z(n22977) );
  NAND U23775 ( .A(n22978), .B(n22977), .Z(n23081) );
  XNOR U23776 ( .A(b[25]), .B(a[142]), .Z(n23120) );
  NANDN U23777 ( .A(n23120), .B(n38325), .Z(n22981) );
  NANDN U23778 ( .A(n22979), .B(n38326), .Z(n22980) );
  AND U23779 ( .A(n22981), .B(n22980), .Z(n23082) );
  XNOR U23780 ( .A(n23081), .B(n23082), .Z(n23083) );
  XOR U23781 ( .A(n23084), .B(n23083), .Z(n23045) );
  XOR U23782 ( .A(n23048), .B(n23047), .Z(n23074) );
  XNOR U23783 ( .A(n23073), .B(n23074), .Z(n23011) );
  XNOR U23784 ( .A(n23012), .B(n23011), .Z(n23014) );
  XNOR U23785 ( .A(n23013), .B(n23014), .Z(n23129) );
  XOR U23786 ( .A(n23130), .B(n23129), .Z(n23132) );
  NANDN U23787 ( .A(n22983), .B(n22982), .Z(n22987) );
  OR U23788 ( .A(n22985), .B(n22984), .Z(n22986) );
  NAND U23789 ( .A(n22987), .B(n22986), .Z(n23123) );
  NAND U23790 ( .A(n22989), .B(n22988), .Z(n22993) );
  NANDN U23791 ( .A(n22991), .B(n22990), .Z(n22992) );
  NAND U23792 ( .A(n22993), .B(n22992), .Z(n23124) );
  XNOR U23793 ( .A(n23123), .B(n23124), .Z(n23125) );
  XOR U23794 ( .A(n23126), .B(n23125), .Z(n23008) );
  XOR U23795 ( .A(n23007), .B(n23008), .Z(n22999) );
  XOR U23796 ( .A(n23000), .B(n22999), .Z(n23001) );
  XNOR U23797 ( .A(n23002), .B(n23001), .Z(n23135) );
  XNOR U23798 ( .A(n23135), .B(sreg[390]), .Z(n23137) );
  NAND U23799 ( .A(n22994), .B(sreg[389]), .Z(n22998) );
  OR U23800 ( .A(n22996), .B(n22995), .Z(n22997) );
  AND U23801 ( .A(n22998), .B(n22997), .Z(n23136) );
  XOR U23802 ( .A(n23137), .B(n23136), .Z(c[390]) );
  NAND U23803 ( .A(n23000), .B(n22999), .Z(n23004) );
  NAND U23804 ( .A(n23002), .B(n23001), .Z(n23003) );
  NAND U23805 ( .A(n23004), .B(n23003), .Z(n23143) );
  NANDN U23806 ( .A(n23006), .B(n23005), .Z(n23010) );
  NAND U23807 ( .A(n23008), .B(n23007), .Z(n23009) );
  NAND U23808 ( .A(n23010), .B(n23009), .Z(n23140) );
  NAND U23809 ( .A(n23012), .B(n23011), .Z(n23016) );
  NANDN U23810 ( .A(n23014), .B(n23013), .Z(n23015) );
  NAND U23811 ( .A(n23016), .B(n23015), .Z(n23266) );
  XNOR U23812 ( .A(n23266), .B(n23267), .Z(n23268) );
  NANDN U23813 ( .A(n23022), .B(n23021), .Z(n23026) );
  NAND U23814 ( .A(n23024), .B(n23023), .Z(n23025) );
  NAND U23815 ( .A(n23026), .B(n23025), .Z(n23211) );
  XNOR U23816 ( .A(b[19]), .B(a[149]), .Z(n23158) );
  NANDN U23817 ( .A(n23158), .B(n37934), .Z(n23029) );
  NANDN U23818 ( .A(n23027), .B(n37935), .Z(n23028) );
  NAND U23819 ( .A(n23029), .B(n23028), .Z(n23221) );
  XNOR U23820 ( .A(b[27]), .B(a[141]), .Z(n23161) );
  NANDN U23821 ( .A(n23161), .B(n38423), .Z(n23032) );
  NAND U23822 ( .A(n23030), .B(n38424), .Z(n23031) );
  NAND U23823 ( .A(n23032), .B(n23031), .Z(n23218) );
  XOR U23824 ( .A(b[5]), .B(n27178), .Z(n23164) );
  NANDN U23825 ( .A(n23164), .B(n36587), .Z(n23035) );
  NANDN U23826 ( .A(n23033), .B(n36588), .Z(n23034) );
  AND U23827 ( .A(n23035), .B(n23034), .Z(n23219) );
  XNOR U23828 ( .A(n23218), .B(n23219), .Z(n23220) );
  XNOR U23829 ( .A(n23221), .B(n23220), .Z(n23209) );
  NAND U23830 ( .A(n23036), .B(n37762), .Z(n23038) );
  XNOR U23831 ( .A(b[17]), .B(a[151]), .Z(n23167) );
  NANDN U23832 ( .A(n23167), .B(n37764), .Z(n23037) );
  NAND U23833 ( .A(n23038), .B(n23037), .Z(n23185) );
  XOR U23834 ( .A(b[31]), .B(n23393), .Z(n23170) );
  NANDN U23835 ( .A(n23170), .B(n38552), .Z(n23041) );
  NANDN U23836 ( .A(n23039), .B(n38553), .Z(n23040) );
  NAND U23837 ( .A(n23041), .B(n23040), .Z(n23182) );
  OR U23838 ( .A(n23042), .B(n36105), .Z(n23044) );
  XNOR U23839 ( .A(b[3]), .B(a[165]), .Z(n23173) );
  NANDN U23840 ( .A(n23173), .B(n36107), .Z(n23043) );
  AND U23841 ( .A(n23044), .B(n23043), .Z(n23183) );
  XNOR U23842 ( .A(n23182), .B(n23183), .Z(n23184) );
  XOR U23843 ( .A(n23185), .B(n23184), .Z(n23208) );
  XNOR U23844 ( .A(n23209), .B(n23208), .Z(n23210) );
  XNOR U23845 ( .A(n23211), .B(n23210), .Z(n23260) );
  NANDN U23846 ( .A(n23046), .B(n23045), .Z(n23050) );
  NANDN U23847 ( .A(n23048), .B(n23047), .Z(n23049) );
  NAND U23848 ( .A(n23050), .B(n23049), .Z(n23261) );
  XNOR U23849 ( .A(n23260), .B(n23261), .Z(n23262) );
  NANDN U23850 ( .A(n23052), .B(n23051), .Z(n23056) );
  NAND U23851 ( .A(n23054), .B(n23053), .Z(n23055) );
  NAND U23852 ( .A(n23056), .B(n23055), .Z(n23201) );
  OR U23853 ( .A(n23058), .B(n23057), .Z(n23062) );
  NANDN U23854 ( .A(n23060), .B(n23059), .Z(n23061) );
  NAND U23855 ( .A(n23062), .B(n23061), .Z(n23199) );
  XNOR U23856 ( .A(n23199), .B(n23198), .Z(n23200) );
  XOR U23857 ( .A(n23201), .B(n23200), .Z(n23263) );
  XOR U23858 ( .A(n23262), .B(n23263), .Z(n23274) );
  NANDN U23859 ( .A(n23072), .B(n23071), .Z(n23076) );
  NANDN U23860 ( .A(n23074), .B(n23073), .Z(n23075) );
  NAND U23861 ( .A(n23076), .B(n23075), .Z(n23257) );
  NANDN U23862 ( .A(n23082), .B(n23081), .Z(n23086) );
  NAND U23863 ( .A(n23084), .B(n23083), .Z(n23085) );
  NAND U23864 ( .A(n23086), .B(n23085), .Z(n23202) );
  NANDN U23865 ( .A(n23088), .B(n23087), .Z(n23092) );
  NAND U23866 ( .A(n23090), .B(n23089), .Z(n23091) );
  AND U23867 ( .A(n23092), .B(n23091), .Z(n23203) );
  XNOR U23868 ( .A(n23202), .B(n23203), .Z(n23204) );
  XOR U23869 ( .A(n1052), .B(a[159]), .Z(n23230) );
  NANDN U23870 ( .A(n23230), .B(n36925), .Z(n23095) );
  NANDN U23871 ( .A(n23093), .B(n36926), .Z(n23094) );
  NAND U23872 ( .A(n23095), .B(n23094), .Z(n23190) );
  XNOR U23873 ( .A(n1054), .B(a[153]), .Z(n23227) );
  NANDN U23874 ( .A(n37665), .B(n23227), .Z(n23098) );
  NANDN U23875 ( .A(n23096), .B(n37604), .Z(n23097) );
  NAND U23876 ( .A(n23098), .B(n23097), .Z(n23188) );
  XOR U23877 ( .A(n1056), .B(a[147]), .Z(n23224) );
  NANDN U23878 ( .A(n23224), .B(n38101), .Z(n23101) );
  NANDN U23879 ( .A(n23099), .B(n38102), .Z(n23100) );
  NAND U23880 ( .A(n23101), .B(n23100), .Z(n23189) );
  XNOR U23881 ( .A(n23188), .B(n23189), .Z(n23191) );
  XOR U23882 ( .A(n23190), .B(n23191), .Z(n23179) );
  XNOR U23883 ( .A(b[11]), .B(a[157]), .Z(n23233) );
  OR U23884 ( .A(n23233), .B(n37311), .Z(n23104) );
  NANDN U23885 ( .A(n23102), .B(n37218), .Z(n23103) );
  NAND U23886 ( .A(n23104), .B(n23103), .Z(n23177) );
  XOR U23887 ( .A(n1053), .B(a[155]), .Z(n23236) );
  NANDN U23888 ( .A(n23236), .B(n37424), .Z(n23107) );
  NANDN U23889 ( .A(n23105), .B(n37425), .Z(n23106) );
  AND U23890 ( .A(n23107), .B(n23106), .Z(n23176) );
  XNOR U23891 ( .A(n23177), .B(n23176), .Z(n23178) );
  XNOR U23892 ( .A(n23179), .B(n23178), .Z(n23195) );
  NANDN U23893 ( .A(n1049), .B(a[167]), .Z(n23108) );
  XNOR U23894 ( .A(b[1]), .B(n23108), .Z(n23110) );
  NANDN U23895 ( .A(b[0]), .B(a[166]), .Z(n23109) );
  AND U23896 ( .A(n23110), .B(n23109), .Z(n23154) );
  NAND U23897 ( .A(n38490), .B(n23111), .Z(n23113) );
  XOR U23898 ( .A(n1058), .B(n23668), .Z(n23242) );
  NANDN U23899 ( .A(n1048), .B(n23242), .Z(n23112) );
  NAND U23900 ( .A(n23113), .B(n23112), .Z(n23152) );
  NANDN U23901 ( .A(n1059), .B(a[135]), .Z(n23153) );
  XNOR U23902 ( .A(n23152), .B(n23153), .Z(n23155) );
  XNOR U23903 ( .A(n23154), .B(n23155), .Z(n23193) );
  NANDN U23904 ( .A(n23114), .B(n38205), .Z(n23116) );
  XOR U23905 ( .A(b[23]), .B(n24554), .Z(n23245) );
  OR U23906 ( .A(n23245), .B(n38268), .Z(n23115) );
  NAND U23907 ( .A(n23116), .B(n23115), .Z(n23215) );
  XNOR U23908 ( .A(b[7]), .B(a[161]), .Z(n23248) );
  NANDN U23909 ( .A(n23248), .B(n36701), .Z(n23119) );
  NAND U23910 ( .A(n23117), .B(n36702), .Z(n23118) );
  NAND U23911 ( .A(n23119), .B(n23118), .Z(n23212) );
  XOR U23912 ( .A(b[25]), .B(a[143]), .Z(n23251) );
  NAND U23913 ( .A(n23251), .B(n38325), .Z(n23122) );
  NANDN U23914 ( .A(n23120), .B(n38326), .Z(n23121) );
  AND U23915 ( .A(n23122), .B(n23121), .Z(n23213) );
  XNOR U23916 ( .A(n23212), .B(n23213), .Z(n23214) );
  XOR U23917 ( .A(n23215), .B(n23214), .Z(n23192) );
  XOR U23918 ( .A(n23195), .B(n23194), .Z(n23205) );
  XOR U23919 ( .A(n23204), .B(n23205), .Z(n23254) );
  XOR U23920 ( .A(n23255), .B(n23254), .Z(n23256) );
  XNOR U23921 ( .A(n23257), .B(n23256), .Z(n23272) );
  XNOR U23922 ( .A(n23273), .B(n23272), .Z(n23275) );
  XNOR U23923 ( .A(n23274), .B(n23275), .Z(n23269) );
  XOR U23924 ( .A(n23268), .B(n23269), .Z(n23149) );
  NANDN U23925 ( .A(n23124), .B(n23123), .Z(n23128) );
  NAND U23926 ( .A(n23126), .B(n23125), .Z(n23127) );
  NAND U23927 ( .A(n23128), .B(n23127), .Z(n23146) );
  NANDN U23928 ( .A(n23130), .B(n23129), .Z(n23134) );
  OR U23929 ( .A(n23132), .B(n23131), .Z(n23133) );
  NAND U23930 ( .A(n23134), .B(n23133), .Z(n23147) );
  XNOR U23931 ( .A(n23146), .B(n23147), .Z(n23148) );
  XNOR U23932 ( .A(n23149), .B(n23148), .Z(n23141) );
  XNOR U23933 ( .A(n23140), .B(n23141), .Z(n23142) );
  XNOR U23934 ( .A(n23143), .B(n23142), .Z(n23278) );
  XNOR U23935 ( .A(n23278), .B(sreg[391]), .Z(n23280) );
  NAND U23936 ( .A(n23135), .B(sreg[390]), .Z(n23139) );
  OR U23937 ( .A(n23137), .B(n23136), .Z(n23138) );
  AND U23938 ( .A(n23139), .B(n23138), .Z(n23279) );
  XOR U23939 ( .A(n23280), .B(n23279), .Z(c[391]) );
  NANDN U23940 ( .A(n23141), .B(n23140), .Z(n23145) );
  NAND U23941 ( .A(n23143), .B(n23142), .Z(n23144) );
  NAND U23942 ( .A(n23145), .B(n23144), .Z(n23286) );
  NANDN U23943 ( .A(n23147), .B(n23146), .Z(n23151) );
  NAND U23944 ( .A(n23149), .B(n23148), .Z(n23150) );
  NAND U23945 ( .A(n23151), .B(n23150), .Z(n23284) );
  NANDN U23946 ( .A(n23153), .B(n23152), .Z(n23157) );
  NAND U23947 ( .A(n23155), .B(n23154), .Z(n23156) );
  NAND U23948 ( .A(n23157), .B(n23156), .Z(n23362) );
  XNOR U23949 ( .A(b[19]), .B(a[150]), .Z(n23309) );
  NANDN U23950 ( .A(n23309), .B(n37934), .Z(n23160) );
  NANDN U23951 ( .A(n23158), .B(n37935), .Z(n23159) );
  NAND U23952 ( .A(n23160), .B(n23159), .Z(n23372) );
  XNOR U23953 ( .A(b[27]), .B(a[142]), .Z(n23312) );
  NANDN U23954 ( .A(n23312), .B(n38423), .Z(n23163) );
  NANDN U23955 ( .A(n23161), .B(n38424), .Z(n23162) );
  NAND U23956 ( .A(n23163), .B(n23162), .Z(n23369) );
  XNOR U23957 ( .A(b[5]), .B(a[164]), .Z(n23315) );
  NANDN U23958 ( .A(n23315), .B(n36587), .Z(n23166) );
  NANDN U23959 ( .A(n23164), .B(n36588), .Z(n23165) );
  AND U23960 ( .A(n23166), .B(n23165), .Z(n23370) );
  XNOR U23961 ( .A(n23369), .B(n23370), .Z(n23371) );
  XNOR U23962 ( .A(n23372), .B(n23371), .Z(n23360) );
  NANDN U23963 ( .A(n23167), .B(n37762), .Z(n23169) );
  XNOR U23964 ( .A(b[17]), .B(a[152]), .Z(n23318) );
  NANDN U23965 ( .A(n23318), .B(n37764), .Z(n23168) );
  NAND U23966 ( .A(n23169), .B(n23168), .Z(n23336) );
  XNOR U23967 ( .A(b[31]), .B(a[138]), .Z(n23321) );
  NANDN U23968 ( .A(n23321), .B(n38552), .Z(n23172) );
  NANDN U23969 ( .A(n23170), .B(n38553), .Z(n23171) );
  NAND U23970 ( .A(n23172), .B(n23171), .Z(n23333) );
  OR U23971 ( .A(n23173), .B(n36105), .Z(n23175) );
  XNOR U23972 ( .A(b[3]), .B(a[166]), .Z(n23324) );
  NANDN U23973 ( .A(n23324), .B(n36107), .Z(n23174) );
  AND U23974 ( .A(n23175), .B(n23174), .Z(n23334) );
  XNOR U23975 ( .A(n23333), .B(n23334), .Z(n23335) );
  XOR U23976 ( .A(n23336), .B(n23335), .Z(n23359) );
  XNOR U23977 ( .A(n23360), .B(n23359), .Z(n23361) );
  XNOR U23978 ( .A(n23362), .B(n23361), .Z(n23300) );
  NANDN U23979 ( .A(n23177), .B(n23176), .Z(n23181) );
  NAND U23980 ( .A(n23179), .B(n23178), .Z(n23180) );
  NAND U23981 ( .A(n23181), .B(n23180), .Z(n23351) );
  NANDN U23982 ( .A(n23183), .B(n23182), .Z(n23187) );
  NAND U23983 ( .A(n23185), .B(n23184), .Z(n23186) );
  NAND U23984 ( .A(n23187), .B(n23186), .Z(n23350) );
  XNOR U23985 ( .A(n23350), .B(n23349), .Z(n23352) );
  XOR U23986 ( .A(n23351), .B(n23352), .Z(n23299) );
  XOR U23987 ( .A(n23300), .B(n23299), .Z(n23301) );
  NANDN U23988 ( .A(n23193), .B(n23192), .Z(n23197) );
  NAND U23989 ( .A(n23195), .B(n23194), .Z(n23196) );
  AND U23990 ( .A(n23197), .B(n23196), .Z(n23302) );
  XNOR U23991 ( .A(n23301), .B(n23302), .Z(n23409) );
  NANDN U23992 ( .A(n23203), .B(n23202), .Z(n23207) );
  NAND U23993 ( .A(n23205), .B(n23204), .Z(n23206) );
  NAND U23994 ( .A(n23207), .B(n23206), .Z(n23296) );
  NANDN U23995 ( .A(n23213), .B(n23212), .Z(n23217) );
  NAND U23996 ( .A(n23215), .B(n23214), .Z(n23216) );
  NAND U23997 ( .A(n23217), .B(n23216), .Z(n23353) );
  NANDN U23998 ( .A(n23219), .B(n23218), .Z(n23223) );
  NAND U23999 ( .A(n23221), .B(n23220), .Z(n23222) );
  AND U24000 ( .A(n23223), .B(n23222), .Z(n23354) );
  XNOR U24001 ( .A(n23353), .B(n23354), .Z(n23355) );
  XOR U24002 ( .A(n1056), .B(a[148]), .Z(n23375) );
  NANDN U24003 ( .A(n23375), .B(n38101), .Z(n23226) );
  NANDN U24004 ( .A(n23224), .B(n38102), .Z(n23225) );
  NAND U24005 ( .A(n23226), .B(n23225), .Z(n23345) );
  XOR U24006 ( .A(b[15]), .B(n25862), .Z(n23378) );
  OR U24007 ( .A(n23378), .B(n37665), .Z(n23229) );
  NAND U24008 ( .A(n23227), .B(n37604), .Z(n23228) );
  AND U24009 ( .A(n23229), .B(n23228), .Z(n23346) );
  XNOR U24010 ( .A(n23345), .B(n23346), .Z(n23348) );
  XOR U24011 ( .A(n1052), .B(a[160]), .Z(n23381) );
  NANDN U24012 ( .A(n23381), .B(n36925), .Z(n23232) );
  NANDN U24013 ( .A(n23230), .B(n36926), .Z(n23231) );
  NAND U24014 ( .A(n23232), .B(n23231), .Z(n23347) );
  XNOR U24015 ( .A(n23348), .B(n23347), .Z(n23341) );
  XNOR U24016 ( .A(b[11]), .B(a[158]), .Z(n23384) );
  OR U24017 ( .A(n23384), .B(n37311), .Z(n23235) );
  NANDN U24018 ( .A(n23233), .B(n37218), .Z(n23234) );
  NAND U24019 ( .A(n23235), .B(n23234), .Z(n23340) );
  XOR U24020 ( .A(n1053), .B(a[156]), .Z(n23387) );
  NANDN U24021 ( .A(n23387), .B(n37424), .Z(n23238) );
  NANDN U24022 ( .A(n23236), .B(n37425), .Z(n23237) );
  NAND U24023 ( .A(n23238), .B(n23237), .Z(n23339) );
  XNOR U24024 ( .A(n23340), .B(n23339), .Z(n23342) );
  XNOR U24025 ( .A(n23341), .B(n23342), .Z(n23330) );
  NANDN U24026 ( .A(n1049), .B(a[168]), .Z(n23239) );
  XNOR U24027 ( .A(b[1]), .B(n23239), .Z(n23241) );
  NANDN U24028 ( .A(b[0]), .B(a[167]), .Z(n23240) );
  AND U24029 ( .A(n23241), .B(n23240), .Z(n23305) );
  NAND U24030 ( .A(n38490), .B(n23242), .Z(n23244) );
  XNOR U24031 ( .A(b[29]), .B(a[140]), .Z(n23394) );
  OR U24032 ( .A(n23394), .B(n1048), .Z(n23243) );
  NAND U24033 ( .A(n23244), .B(n23243), .Z(n23303) );
  NANDN U24034 ( .A(n1059), .B(a[136]), .Z(n23304) );
  XNOR U24035 ( .A(n23303), .B(n23304), .Z(n23306) );
  XNOR U24036 ( .A(n23305), .B(n23306), .Z(n23328) );
  NANDN U24037 ( .A(n23245), .B(n38205), .Z(n23247) );
  XNOR U24038 ( .A(b[23]), .B(a[146]), .Z(n23397) );
  OR U24039 ( .A(n23397), .B(n38268), .Z(n23246) );
  NAND U24040 ( .A(n23247), .B(n23246), .Z(n23366) );
  XOR U24041 ( .A(b[7]), .B(a[162]), .Z(n23400) );
  NAND U24042 ( .A(n23400), .B(n36701), .Z(n23250) );
  NANDN U24043 ( .A(n23248), .B(n36702), .Z(n23249) );
  NAND U24044 ( .A(n23250), .B(n23249), .Z(n23363) );
  XOR U24045 ( .A(b[25]), .B(a[144]), .Z(n23403) );
  NAND U24046 ( .A(n23403), .B(n38325), .Z(n23253) );
  NAND U24047 ( .A(n23251), .B(n38326), .Z(n23252) );
  AND U24048 ( .A(n23253), .B(n23252), .Z(n23364) );
  XNOR U24049 ( .A(n23363), .B(n23364), .Z(n23365) );
  XOR U24050 ( .A(n23366), .B(n23365), .Z(n23327) );
  XOR U24051 ( .A(n23330), .B(n23329), .Z(n23356) );
  XNOR U24052 ( .A(n23355), .B(n23356), .Z(n23293) );
  XOR U24053 ( .A(n23294), .B(n23293), .Z(n23295) );
  XOR U24054 ( .A(n23296), .B(n23295), .Z(n23407) );
  XNOR U24055 ( .A(n23406), .B(n23407), .Z(n23408) );
  XNOR U24056 ( .A(n23409), .B(n23408), .Z(n23413) );
  NAND U24057 ( .A(n23255), .B(n23254), .Z(n23259) );
  NAND U24058 ( .A(n23257), .B(n23256), .Z(n23258) );
  NAND U24059 ( .A(n23259), .B(n23258), .Z(n23410) );
  NANDN U24060 ( .A(n23261), .B(n23260), .Z(n23265) );
  NAND U24061 ( .A(n23263), .B(n23262), .Z(n23264) );
  NAND U24062 ( .A(n23265), .B(n23264), .Z(n23411) );
  XNOR U24063 ( .A(n23410), .B(n23411), .Z(n23412) );
  XNOR U24064 ( .A(n23413), .B(n23412), .Z(n23290) );
  NANDN U24065 ( .A(n23267), .B(n23266), .Z(n23271) );
  NANDN U24066 ( .A(n23269), .B(n23268), .Z(n23270) );
  NAND U24067 ( .A(n23271), .B(n23270), .Z(n23288) );
  OR U24068 ( .A(n23273), .B(n23272), .Z(n23277) );
  OR U24069 ( .A(n23275), .B(n23274), .Z(n23276) );
  AND U24070 ( .A(n23277), .B(n23276), .Z(n23287) );
  XNOR U24071 ( .A(n23288), .B(n23287), .Z(n23289) );
  XNOR U24072 ( .A(n23290), .B(n23289), .Z(n23283) );
  XOR U24073 ( .A(n23284), .B(n23283), .Z(n23285) );
  XNOR U24074 ( .A(n23286), .B(n23285), .Z(n23416) );
  XNOR U24075 ( .A(n23416), .B(sreg[392]), .Z(n23418) );
  NAND U24076 ( .A(n23278), .B(sreg[391]), .Z(n23282) );
  OR U24077 ( .A(n23280), .B(n23279), .Z(n23281) );
  AND U24078 ( .A(n23282), .B(n23281), .Z(n23417) );
  XOR U24079 ( .A(n23418), .B(n23417), .Z(c[392]) );
  NANDN U24080 ( .A(n23288), .B(n23287), .Z(n23292) );
  NANDN U24081 ( .A(n23290), .B(n23289), .Z(n23291) );
  NAND U24082 ( .A(n23292), .B(n23291), .Z(n23421) );
  NAND U24083 ( .A(n23294), .B(n23293), .Z(n23298) );
  NAND U24084 ( .A(n23296), .B(n23295), .Z(n23297) );
  NAND U24085 ( .A(n23298), .B(n23297), .Z(n23547) );
  XNOR U24086 ( .A(n23547), .B(n23548), .Z(n23549) );
  NANDN U24087 ( .A(n23304), .B(n23303), .Z(n23308) );
  NAND U24088 ( .A(n23306), .B(n23305), .Z(n23307) );
  NAND U24089 ( .A(n23308), .B(n23307), .Z(n23446) );
  XOR U24090 ( .A(b[19]), .B(n25435), .Z(n23495) );
  NANDN U24091 ( .A(n23495), .B(n37934), .Z(n23311) );
  NANDN U24092 ( .A(n23309), .B(n37935), .Z(n23310) );
  NAND U24093 ( .A(n23311), .B(n23310), .Z(n23456) );
  XOR U24094 ( .A(b[27]), .B(a[143]), .Z(n23498) );
  NAND U24095 ( .A(n38423), .B(n23498), .Z(n23314) );
  NANDN U24096 ( .A(n23312), .B(n38424), .Z(n23313) );
  NAND U24097 ( .A(n23314), .B(n23313), .Z(n23453) );
  XNOR U24098 ( .A(b[5]), .B(a[165]), .Z(n23501) );
  NANDN U24099 ( .A(n23501), .B(n36587), .Z(n23317) );
  NANDN U24100 ( .A(n23315), .B(n36588), .Z(n23316) );
  AND U24101 ( .A(n23317), .B(n23316), .Z(n23454) );
  XNOR U24102 ( .A(n23453), .B(n23454), .Z(n23455) );
  XNOR U24103 ( .A(n23456), .B(n23455), .Z(n23444) );
  NANDN U24104 ( .A(n23318), .B(n37762), .Z(n23320) );
  XOR U24105 ( .A(b[17]), .B(a[153]), .Z(n23504) );
  NAND U24106 ( .A(n23504), .B(n37764), .Z(n23319) );
  NAND U24107 ( .A(n23320), .B(n23319), .Z(n23522) );
  XOR U24108 ( .A(b[31]), .B(n23668), .Z(n23507) );
  NANDN U24109 ( .A(n23507), .B(n38552), .Z(n23323) );
  NANDN U24110 ( .A(n23321), .B(n38553), .Z(n23322) );
  NAND U24111 ( .A(n23323), .B(n23322), .Z(n23519) );
  OR U24112 ( .A(n23324), .B(n36105), .Z(n23326) );
  XNOR U24113 ( .A(b[3]), .B(a[167]), .Z(n23510) );
  NANDN U24114 ( .A(n23510), .B(n36107), .Z(n23325) );
  AND U24115 ( .A(n23326), .B(n23325), .Z(n23520) );
  XNOR U24116 ( .A(n23519), .B(n23520), .Z(n23521) );
  XOR U24117 ( .A(n23522), .B(n23521), .Z(n23443) );
  XNOR U24118 ( .A(n23444), .B(n23443), .Z(n23445) );
  XNOR U24119 ( .A(n23446), .B(n23445), .Z(n23541) );
  NANDN U24120 ( .A(n23328), .B(n23327), .Z(n23332) );
  NANDN U24121 ( .A(n23330), .B(n23329), .Z(n23331) );
  NAND U24122 ( .A(n23332), .B(n23331), .Z(n23542) );
  XNOR U24123 ( .A(n23541), .B(n23542), .Z(n23543) );
  NANDN U24124 ( .A(n23334), .B(n23333), .Z(n23338) );
  NAND U24125 ( .A(n23336), .B(n23335), .Z(n23337) );
  NAND U24126 ( .A(n23338), .B(n23337), .Z(n23436) );
  OR U24127 ( .A(n23340), .B(n23339), .Z(n23344) );
  NANDN U24128 ( .A(n23342), .B(n23341), .Z(n23343) );
  NAND U24129 ( .A(n23344), .B(n23343), .Z(n23434) );
  XNOR U24130 ( .A(n23434), .B(n23433), .Z(n23435) );
  XOR U24131 ( .A(n23436), .B(n23435), .Z(n23544) );
  XOR U24132 ( .A(n23543), .B(n23544), .Z(n23555) );
  NANDN U24133 ( .A(n23354), .B(n23353), .Z(n23358) );
  NANDN U24134 ( .A(n23356), .B(n23355), .Z(n23357) );
  NAND U24135 ( .A(n23358), .B(n23357), .Z(n23538) );
  NANDN U24136 ( .A(n23364), .B(n23363), .Z(n23368) );
  NAND U24137 ( .A(n23366), .B(n23365), .Z(n23367) );
  NAND U24138 ( .A(n23368), .B(n23367), .Z(n23437) );
  NANDN U24139 ( .A(n23370), .B(n23369), .Z(n23374) );
  NAND U24140 ( .A(n23372), .B(n23371), .Z(n23373) );
  AND U24141 ( .A(n23374), .B(n23373), .Z(n23438) );
  XNOR U24142 ( .A(n23437), .B(n23438), .Z(n23439) );
  XNOR U24143 ( .A(b[21]), .B(a[149]), .Z(n23465) );
  NANDN U24144 ( .A(n23465), .B(n38101), .Z(n23377) );
  NANDN U24145 ( .A(n23375), .B(n38102), .Z(n23376) );
  NAND U24146 ( .A(n23377), .B(n23376), .Z(n23531) );
  XNOR U24147 ( .A(b[15]), .B(a[155]), .Z(n23462) );
  OR U24148 ( .A(n23462), .B(n37665), .Z(n23380) );
  NANDN U24149 ( .A(n23378), .B(n37604), .Z(n23379) );
  AND U24150 ( .A(n23380), .B(n23379), .Z(n23532) );
  XNOR U24151 ( .A(n23531), .B(n23532), .Z(n23534) );
  XOR U24152 ( .A(b[9]), .B(n26869), .Z(n23459) );
  NANDN U24153 ( .A(n23459), .B(n36925), .Z(n23383) );
  NANDN U24154 ( .A(n23381), .B(n36926), .Z(n23382) );
  NAND U24155 ( .A(n23383), .B(n23382), .Z(n23533) );
  XNOR U24156 ( .A(n23534), .B(n23533), .Z(n23527) );
  XNOR U24157 ( .A(b[11]), .B(a[159]), .Z(n23468) );
  OR U24158 ( .A(n23468), .B(n37311), .Z(n23386) );
  NANDN U24159 ( .A(n23384), .B(n37218), .Z(n23385) );
  NAND U24160 ( .A(n23386), .B(n23385), .Z(n23526) );
  XOR U24161 ( .A(n1053), .B(a[157]), .Z(n23471) );
  NANDN U24162 ( .A(n23471), .B(n37424), .Z(n23389) );
  NANDN U24163 ( .A(n23387), .B(n37425), .Z(n23388) );
  NAND U24164 ( .A(n23389), .B(n23388), .Z(n23525) );
  XNOR U24165 ( .A(n23526), .B(n23525), .Z(n23528) );
  XNOR U24166 ( .A(n23527), .B(n23528), .Z(n23516) );
  NANDN U24167 ( .A(n1049), .B(a[169]), .Z(n23390) );
  XNOR U24168 ( .A(b[1]), .B(n23390), .Z(n23392) );
  NANDN U24169 ( .A(b[0]), .B(a[168]), .Z(n23391) );
  AND U24170 ( .A(n23392), .B(n23391), .Z(n23492) );
  ANDN U24171 ( .B(b[31]), .A(n23393), .Z(n23489) );
  NANDN U24172 ( .A(n23394), .B(n38490), .Z(n23396) );
  XNOR U24173 ( .A(n1058), .B(a[141]), .Z(n23477) );
  NANDN U24174 ( .A(n1048), .B(n23477), .Z(n23395) );
  NAND U24175 ( .A(n23396), .B(n23395), .Z(n23490) );
  XOR U24176 ( .A(n23489), .B(n23490), .Z(n23491) );
  XNOR U24177 ( .A(n23492), .B(n23491), .Z(n23513) );
  NANDN U24178 ( .A(n23397), .B(n38205), .Z(n23399) );
  XNOR U24179 ( .A(b[23]), .B(a[147]), .Z(n23480) );
  OR U24180 ( .A(n23480), .B(n38268), .Z(n23398) );
  NAND U24181 ( .A(n23399), .B(n23398), .Z(n23450) );
  XNOR U24182 ( .A(b[7]), .B(a[163]), .Z(n23483) );
  NANDN U24183 ( .A(n23483), .B(n36701), .Z(n23402) );
  NAND U24184 ( .A(n23400), .B(n36702), .Z(n23401) );
  NAND U24185 ( .A(n23402), .B(n23401), .Z(n23447) );
  XNOR U24186 ( .A(b[25]), .B(a[145]), .Z(n23486) );
  NANDN U24187 ( .A(n23486), .B(n38325), .Z(n23405) );
  NAND U24188 ( .A(n23403), .B(n38326), .Z(n23404) );
  AND U24189 ( .A(n23405), .B(n23404), .Z(n23448) );
  XNOR U24190 ( .A(n23447), .B(n23448), .Z(n23449) );
  XNOR U24191 ( .A(n23450), .B(n23449), .Z(n23514) );
  XOR U24192 ( .A(n23516), .B(n23515), .Z(n23440) );
  XNOR U24193 ( .A(n23439), .B(n23440), .Z(n23535) );
  XOR U24194 ( .A(n23536), .B(n23535), .Z(n23537) );
  XNOR U24195 ( .A(n23538), .B(n23537), .Z(n23553) );
  XNOR U24196 ( .A(n23554), .B(n23553), .Z(n23556) );
  XNOR U24197 ( .A(n23555), .B(n23556), .Z(n23550) );
  XOR U24198 ( .A(n23549), .B(n23550), .Z(n23430) );
  NANDN U24199 ( .A(n23411), .B(n23410), .Z(n23415) );
  NANDN U24200 ( .A(n23413), .B(n23412), .Z(n23414) );
  NAND U24201 ( .A(n23415), .B(n23414), .Z(n23428) );
  XNOR U24202 ( .A(n23427), .B(n23428), .Z(n23429) );
  XNOR U24203 ( .A(n23430), .B(n23429), .Z(n23422) );
  XNOR U24204 ( .A(n23421), .B(n23422), .Z(n23423) );
  XNOR U24205 ( .A(n23424), .B(n23423), .Z(n23559) );
  XNOR U24206 ( .A(n23559), .B(sreg[393]), .Z(n23561) );
  NAND U24207 ( .A(n23416), .B(sreg[392]), .Z(n23420) );
  OR U24208 ( .A(n23418), .B(n23417), .Z(n23419) );
  AND U24209 ( .A(n23420), .B(n23419), .Z(n23560) );
  XOR U24210 ( .A(n23561), .B(n23560), .Z(c[393]) );
  NANDN U24211 ( .A(n23422), .B(n23421), .Z(n23426) );
  NAND U24212 ( .A(n23424), .B(n23423), .Z(n23425) );
  NAND U24213 ( .A(n23426), .B(n23425), .Z(n23567) );
  NANDN U24214 ( .A(n23428), .B(n23427), .Z(n23432) );
  NAND U24215 ( .A(n23430), .B(n23429), .Z(n23431) );
  NAND U24216 ( .A(n23432), .B(n23431), .Z(n23565) );
  NANDN U24217 ( .A(n23438), .B(n23437), .Z(n23442) );
  NANDN U24218 ( .A(n23440), .B(n23439), .Z(n23441) );
  NAND U24219 ( .A(n23442), .B(n23441), .Z(n23684) );
  NANDN U24220 ( .A(n23448), .B(n23447), .Z(n23452) );
  NAND U24221 ( .A(n23450), .B(n23449), .Z(n23451) );
  NAND U24222 ( .A(n23452), .B(n23451), .Z(n23626) );
  NANDN U24223 ( .A(n23454), .B(n23453), .Z(n23458) );
  NAND U24224 ( .A(n23456), .B(n23455), .Z(n23457) );
  AND U24225 ( .A(n23458), .B(n23457), .Z(n23627) );
  XNOR U24226 ( .A(n23626), .B(n23627), .Z(n23628) );
  XNOR U24227 ( .A(b[9]), .B(a[162]), .Z(n23650) );
  NANDN U24228 ( .A(n23650), .B(n36925), .Z(n23461) );
  NANDN U24229 ( .A(n23459), .B(n36926), .Z(n23460) );
  NAND U24230 ( .A(n23461), .B(n23460), .Z(n23612) );
  XNOR U24231 ( .A(b[15]), .B(a[156]), .Z(n23653) );
  OR U24232 ( .A(n23653), .B(n37665), .Z(n23464) );
  NANDN U24233 ( .A(n23462), .B(n37604), .Z(n23463) );
  AND U24234 ( .A(n23464), .B(n23463), .Z(n23610) );
  XNOR U24235 ( .A(b[21]), .B(a[150]), .Z(n23656) );
  NANDN U24236 ( .A(n23656), .B(n38101), .Z(n23467) );
  NANDN U24237 ( .A(n23465), .B(n38102), .Z(n23466) );
  AND U24238 ( .A(n23467), .B(n23466), .Z(n23611) );
  XOR U24239 ( .A(n23612), .B(n23613), .Z(n23601) );
  XNOR U24240 ( .A(b[11]), .B(a[160]), .Z(n23659) );
  OR U24241 ( .A(n23659), .B(n37311), .Z(n23470) );
  NANDN U24242 ( .A(n23468), .B(n37218), .Z(n23469) );
  NAND U24243 ( .A(n23470), .B(n23469), .Z(n23599) );
  XOR U24244 ( .A(n1053), .B(a[158]), .Z(n23662) );
  NANDN U24245 ( .A(n23662), .B(n37424), .Z(n23473) );
  NANDN U24246 ( .A(n23471), .B(n37425), .Z(n23472) );
  AND U24247 ( .A(n23473), .B(n23472), .Z(n23598) );
  XNOR U24248 ( .A(n23599), .B(n23598), .Z(n23600) );
  XOR U24249 ( .A(n23601), .B(n23600), .Z(n23618) );
  NANDN U24250 ( .A(n1049), .B(a[170]), .Z(n23474) );
  XNOR U24251 ( .A(b[1]), .B(n23474), .Z(n23476) );
  NANDN U24252 ( .A(b[0]), .B(a[169]), .Z(n23475) );
  AND U24253 ( .A(n23476), .B(n23475), .Z(n23576) );
  NAND U24254 ( .A(n23477), .B(n38490), .Z(n23479) );
  XOR U24255 ( .A(b[29]), .B(n24120), .Z(n23669) );
  OR U24256 ( .A(n23669), .B(n1048), .Z(n23478) );
  NAND U24257 ( .A(n23479), .B(n23478), .Z(n23574) );
  NANDN U24258 ( .A(n1059), .B(a[138]), .Z(n23575) );
  XNOR U24259 ( .A(n23574), .B(n23575), .Z(n23577) );
  XOR U24260 ( .A(n23576), .B(n23577), .Z(n23616) );
  NANDN U24261 ( .A(n23480), .B(n38205), .Z(n23482) );
  XNOR U24262 ( .A(b[23]), .B(a[148]), .Z(n23672) );
  OR U24263 ( .A(n23672), .B(n38268), .Z(n23481) );
  NAND U24264 ( .A(n23482), .B(n23481), .Z(n23641) );
  XOR U24265 ( .A(b[7]), .B(a[164]), .Z(n23675) );
  NAND U24266 ( .A(n23675), .B(n36701), .Z(n23485) );
  NANDN U24267 ( .A(n23483), .B(n36702), .Z(n23484) );
  NAND U24268 ( .A(n23485), .B(n23484), .Z(n23638) );
  XOR U24269 ( .A(b[25]), .B(a[146]), .Z(n23678) );
  NAND U24270 ( .A(n23678), .B(n38325), .Z(n23488) );
  NANDN U24271 ( .A(n23486), .B(n38326), .Z(n23487) );
  AND U24272 ( .A(n23488), .B(n23487), .Z(n23639) );
  XNOR U24273 ( .A(n23638), .B(n23639), .Z(n23640) );
  XNOR U24274 ( .A(n23641), .B(n23640), .Z(n23617) );
  XOR U24275 ( .A(n23616), .B(n23617), .Z(n23619) );
  XNOR U24276 ( .A(n23618), .B(n23619), .Z(n23629) );
  XOR U24277 ( .A(n23628), .B(n23629), .Z(n23682) );
  XNOR U24278 ( .A(n23681), .B(n23682), .Z(n23683) );
  XOR U24279 ( .A(n23684), .B(n23683), .Z(n23694) );
  XNOR U24280 ( .A(n23693), .B(n23694), .Z(n23696) );
  OR U24281 ( .A(n23490), .B(n23489), .Z(n23494) );
  NANDN U24282 ( .A(n23492), .B(n23491), .Z(n23493) );
  NAND U24283 ( .A(n23494), .B(n23493), .Z(n23634) );
  XOR U24284 ( .A(b[19]), .B(n25213), .Z(n23580) );
  NANDN U24285 ( .A(n23580), .B(n37934), .Z(n23497) );
  NANDN U24286 ( .A(n23495), .B(n37935), .Z(n23496) );
  NAND U24287 ( .A(n23497), .B(n23496), .Z(n23647) );
  XOR U24288 ( .A(b[27]), .B(a[144]), .Z(n23583) );
  NAND U24289 ( .A(n38423), .B(n23583), .Z(n23500) );
  NAND U24290 ( .A(n23498), .B(n38424), .Z(n23499) );
  NAND U24291 ( .A(n23500), .B(n23499), .Z(n23644) );
  XNOR U24292 ( .A(b[5]), .B(a[166]), .Z(n23586) );
  NANDN U24293 ( .A(n23586), .B(n36587), .Z(n23503) );
  NANDN U24294 ( .A(n23501), .B(n36588), .Z(n23502) );
  AND U24295 ( .A(n23503), .B(n23502), .Z(n23645) );
  XNOR U24296 ( .A(n23644), .B(n23645), .Z(n23646) );
  XNOR U24297 ( .A(n23647), .B(n23646), .Z(n23633) );
  NAND U24298 ( .A(n23504), .B(n37762), .Z(n23506) );
  XNOR U24299 ( .A(b[17]), .B(a[154]), .Z(n23589) );
  NANDN U24300 ( .A(n23589), .B(n37764), .Z(n23505) );
  NAND U24301 ( .A(n23506), .B(n23505), .Z(n23607) );
  XNOR U24302 ( .A(b[31]), .B(a[140]), .Z(n23592) );
  NANDN U24303 ( .A(n23592), .B(n38552), .Z(n23509) );
  NANDN U24304 ( .A(n23507), .B(n38553), .Z(n23508) );
  NAND U24305 ( .A(n23509), .B(n23508), .Z(n23604) );
  OR U24306 ( .A(n23510), .B(n36105), .Z(n23512) );
  XNOR U24307 ( .A(b[3]), .B(a[168]), .Z(n23595) );
  NANDN U24308 ( .A(n23595), .B(n36107), .Z(n23511) );
  AND U24309 ( .A(n23512), .B(n23511), .Z(n23605) );
  XNOR U24310 ( .A(n23604), .B(n23605), .Z(n23606) );
  XOR U24311 ( .A(n23607), .B(n23606), .Z(n23632) );
  XOR U24312 ( .A(n23633), .B(n23632), .Z(n23635) );
  XNOR U24313 ( .A(n23634), .B(n23635), .Z(n23687) );
  OR U24314 ( .A(n23514), .B(n23513), .Z(n23518) );
  NANDN U24315 ( .A(n23516), .B(n23515), .Z(n23517) );
  NAND U24316 ( .A(n23518), .B(n23517), .Z(n23688) );
  XNOR U24317 ( .A(n23687), .B(n23688), .Z(n23689) );
  NANDN U24318 ( .A(n23520), .B(n23519), .Z(n23524) );
  NAND U24319 ( .A(n23522), .B(n23521), .Z(n23523) );
  NAND U24320 ( .A(n23524), .B(n23523), .Z(n23625) );
  OR U24321 ( .A(n23526), .B(n23525), .Z(n23530) );
  NANDN U24322 ( .A(n23528), .B(n23527), .Z(n23529) );
  NAND U24323 ( .A(n23530), .B(n23529), .Z(n23623) );
  XNOR U24324 ( .A(n23623), .B(n23622), .Z(n23624) );
  XOR U24325 ( .A(n23625), .B(n23624), .Z(n23690) );
  XOR U24326 ( .A(n23689), .B(n23690), .Z(n23695) );
  XOR U24327 ( .A(n23696), .B(n23695), .Z(n23700) );
  NAND U24328 ( .A(n23536), .B(n23535), .Z(n23540) );
  NAND U24329 ( .A(n23538), .B(n23537), .Z(n23539) );
  NAND U24330 ( .A(n23540), .B(n23539), .Z(n23697) );
  NANDN U24331 ( .A(n23542), .B(n23541), .Z(n23546) );
  NAND U24332 ( .A(n23544), .B(n23543), .Z(n23545) );
  NAND U24333 ( .A(n23546), .B(n23545), .Z(n23698) );
  XNOR U24334 ( .A(n23697), .B(n23698), .Z(n23699) );
  XNOR U24335 ( .A(n23700), .B(n23699), .Z(n23571) );
  NANDN U24336 ( .A(n23548), .B(n23547), .Z(n23552) );
  NANDN U24337 ( .A(n23550), .B(n23549), .Z(n23551) );
  NAND U24338 ( .A(n23552), .B(n23551), .Z(n23569) );
  OR U24339 ( .A(n23554), .B(n23553), .Z(n23558) );
  OR U24340 ( .A(n23556), .B(n23555), .Z(n23557) );
  AND U24341 ( .A(n23558), .B(n23557), .Z(n23568) );
  XNOR U24342 ( .A(n23569), .B(n23568), .Z(n23570) );
  XNOR U24343 ( .A(n23571), .B(n23570), .Z(n23564) );
  XOR U24344 ( .A(n23565), .B(n23564), .Z(n23566) );
  XNOR U24345 ( .A(n23567), .B(n23566), .Z(n23703) );
  XNOR U24346 ( .A(n23703), .B(sreg[394]), .Z(n23705) );
  NAND U24347 ( .A(n23559), .B(sreg[393]), .Z(n23563) );
  OR U24348 ( .A(n23561), .B(n23560), .Z(n23562) );
  AND U24349 ( .A(n23563), .B(n23562), .Z(n23704) );
  XOR U24350 ( .A(n23705), .B(n23704), .Z(c[394]) );
  NANDN U24351 ( .A(n23569), .B(n23568), .Z(n23573) );
  NANDN U24352 ( .A(n23571), .B(n23570), .Z(n23572) );
  NAND U24353 ( .A(n23573), .B(n23572), .Z(n23709) );
  NANDN U24354 ( .A(n23575), .B(n23574), .Z(n23579) );
  NAND U24355 ( .A(n23577), .B(n23576), .Z(n23578) );
  NAND U24356 ( .A(n23579), .B(n23578), .Z(n23791) );
  XNOR U24357 ( .A(b[19]), .B(a[153]), .Z(n23758) );
  NANDN U24358 ( .A(n23758), .B(n37934), .Z(n23582) );
  NANDN U24359 ( .A(n23580), .B(n37935), .Z(n23581) );
  NAND U24360 ( .A(n23582), .B(n23581), .Z(n23803) );
  XNOR U24361 ( .A(b[27]), .B(a[145]), .Z(n23761) );
  NANDN U24362 ( .A(n23761), .B(n38423), .Z(n23585) );
  NAND U24363 ( .A(n23583), .B(n38424), .Z(n23584) );
  NAND U24364 ( .A(n23585), .B(n23584), .Z(n23800) );
  XNOR U24365 ( .A(b[5]), .B(a[167]), .Z(n23764) );
  NANDN U24366 ( .A(n23764), .B(n36587), .Z(n23588) );
  NANDN U24367 ( .A(n23586), .B(n36588), .Z(n23587) );
  AND U24368 ( .A(n23588), .B(n23587), .Z(n23801) );
  XNOR U24369 ( .A(n23800), .B(n23801), .Z(n23802) );
  XNOR U24370 ( .A(n23803), .B(n23802), .Z(n23788) );
  NANDN U24371 ( .A(n23589), .B(n37762), .Z(n23591) );
  XOR U24372 ( .A(b[17]), .B(a[155]), .Z(n23767) );
  NAND U24373 ( .A(n23767), .B(n37764), .Z(n23590) );
  NAND U24374 ( .A(n23591), .B(n23590), .Z(n23742) );
  XOR U24375 ( .A(b[31]), .B(n23961), .Z(n23770) );
  NANDN U24376 ( .A(n23770), .B(n38552), .Z(n23594) );
  NANDN U24377 ( .A(n23592), .B(n38553), .Z(n23593) );
  AND U24378 ( .A(n23594), .B(n23593), .Z(n23740) );
  OR U24379 ( .A(n23595), .B(n36105), .Z(n23597) );
  XNOR U24380 ( .A(b[3]), .B(a[169]), .Z(n23773) );
  NANDN U24381 ( .A(n23773), .B(n36107), .Z(n23596) );
  AND U24382 ( .A(n23597), .B(n23596), .Z(n23741) );
  XOR U24383 ( .A(n23742), .B(n23743), .Z(n23789) );
  XOR U24384 ( .A(n23788), .B(n23789), .Z(n23790) );
  XNOR U24385 ( .A(n23791), .B(n23790), .Z(n23836) );
  NANDN U24386 ( .A(n23599), .B(n23598), .Z(n23603) );
  NAND U24387 ( .A(n23601), .B(n23600), .Z(n23602) );
  NAND U24388 ( .A(n23603), .B(n23602), .Z(n23779) );
  NANDN U24389 ( .A(n23605), .B(n23604), .Z(n23609) );
  NAND U24390 ( .A(n23607), .B(n23606), .Z(n23608) );
  NAND U24391 ( .A(n23609), .B(n23608), .Z(n23777) );
  OR U24392 ( .A(n23611), .B(n23610), .Z(n23615) );
  NANDN U24393 ( .A(n23613), .B(n23612), .Z(n23614) );
  NAND U24394 ( .A(n23615), .B(n23614), .Z(n23776) );
  XNOR U24395 ( .A(n23779), .B(n23778), .Z(n23837) );
  XNOR U24396 ( .A(n23836), .B(n23837), .Z(n23838) );
  NANDN U24397 ( .A(n23617), .B(n23616), .Z(n23621) );
  OR U24398 ( .A(n23619), .B(n23618), .Z(n23620) );
  AND U24399 ( .A(n23621), .B(n23620), .Z(n23839) );
  XNOR U24400 ( .A(n23838), .B(n23839), .Z(n23721) );
  NANDN U24401 ( .A(n23627), .B(n23626), .Z(n23631) );
  NANDN U24402 ( .A(n23629), .B(n23628), .Z(n23630) );
  NAND U24403 ( .A(n23631), .B(n23630), .Z(n23845) );
  NANDN U24404 ( .A(n23633), .B(n23632), .Z(n23637) );
  OR U24405 ( .A(n23635), .B(n23634), .Z(n23636) );
  NAND U24406 ( .A(n23637), .B(n23636), .Z(n23843) );
  NANDN U24407 ( .A(n23639), .B(n23638), .Z(n23643) );
  NAND U24408 ( .A(n23641), .B(n23640), .Z(n23642) );
  NAND U24409 ( .A(n23643), .B(n23642), .Z(n23782) );
  NANDN U24410 ( .A(n23645), .B(n23644), .Z(n23649) );
  NAND U24411 ( .A(n23647), .B(n23646), .Z(n23648) );
  AND U24412 ( .A(n23649), .B(n23648), .Z(n23783) );
  XNOR U24413 ( .A(n23782), .B(n23783), .Z(n23784) );
  XOR U24414 ( .A(b[9]), .B(n27178), .Z(n23806) );
  NANDN U24415 ( .A(n23806), .B(n36925), .Z(n23652) );
  NANDN U24416 ( .A(n23650), .B(n36926), .Z(n23651) );
  NAND U24417 ( .A(n23652), .B(n23651), .Z(n23748) );
  XNOR U24418 ( .A(b[15]), .B(a[157]), .Z(n23809) );
  OR U24419 ( .A(n23809), .B(n37665), .Z(n23655) );
  NANDN U24420 ( .A(n23653), .B(n37604), .Z(n23654) );
  AND U24421 ( .A(n23655), .B(n23654), .Z(n23746) );
  XOR U24422 ( .A(b[21]), .B(n25435), .Z(n23812) );
  NANDN U24423 ( .A(n23812), .B(n38101), .Z(n23658) );
  NANDN U24424 ( .A(n23656), .B(n38102), .Z(n23657) );
  AND U24425 ( .A(n23658), .B(n23657), .Z(n23747) );
  XOR U24426 ( .A(n23748), .B(n23749), .Z(n23737) );
  XOR U24427 ( .A(b[11]), .B(n26869), .Z(n23815) );
  OR U24428 ( .A(n23815), .B(n37311), .Z(n23661) );
  NANDN U24429 ( .A(n23659), .B(n37218), .Z(n23660) );
  NAND U24430 ( .A(n23661), .B(n23660), .Z(n23735) );
  XOR U24431 ( .A(n1053), .B(a[159]), .Z(n23818) );
  NANDN U24432 ( .A(n23818), .B(n37424), .Z(n23664) );
  NANDN U24433 ( .A(n23662), .B(n37425), .Z(n23663) );
  NAND U24434 ( .A(n23664), .B(n23663), .Z(n23734) );
  XOR U24435 ( .A(n23737), .B(n23736), .Z(n23731) );
  NANDN U24436 ( .A(n1049), .B(a[171]), .Z(n23665) );
  XNOR U24437 ( .A(b[1]), .B(n23665), .Z(n23667) );
  NANDN U24438 ( .A(b[0]), .B(a[170]), .Z(n23666) );
  AND U24439 ( .A(n23667), .B(n23666), .Z(n23755) );
  ANDN U24440 ( .B(b[31]), .A(n23668), .Z(n23752) );
  NANDN U24441 ( .A(n23669), .B(n38490), .Z(n23671) );
  XNOR U24442 ( .A(n1058), .B(a[143]), .Z(n23821) );
  NANDN U24443 ( .A(n1048), .B(n23821), .Z(n23670) );
  NAND U24444 ( .A(n23671), .B(n23670), .Z(n23753) );
  XOR U24445 ( .A(n23752), .B(n23753), .Z(n23754) );
  XNOR U24446 ( .A(n23755), .B(n23754), .Z(n23728) );
  NANDN U24447 ( .A(n23672), .B(n38205), .Z(n23674) );
  XNOR U24448 ( .A(b[23]), .B(a[149]), .Z(n23827) );
  OR U24449 ( .A(n23827), .B(n38268), .Z(n23673) );
  NAND U24450 ( .A(n23674), .B(n23673), .Z(n23797) );
  XOR U24451 ( .A(b[7]), .B(a[165]), .Z(n23830) );
  NAND U24452 ( .A(n23830), .B(n36701), .Z(n23677) );
  NAND U24453 ( .A(n23675), .B(n36702), .Z(n23676) );
  NAND U24454 ( .A(n23677), .B(n23676), .Z(n23794) );
  XOR U24455 ( .A(b[25]), .B(a[147]), .Z(n23833) );
  NAND U24456 ( .A(n23833), .B(n38325), .Z(n23680) );
  NAND U24457 ( .A(n23678), .B(n38326), .Z(n23679) );
  AND U24458 ( .A(n23680), .B(n23679), .Z(n23795) );
  XNOR U24459 ( .A(n23794), .B(n23795), .Z(n23796) );
  XNOR U24460 ( .A(n23797), .B(n23796), .Z(n23729) );
  XOR U24461 ( .A(n23731), .B(n23730), .Z(n23785) );
  XNOR U24462 ( .A(n23784), .B(n23785), .Z(n23842) );
  XOR U24463 ( .A(n23843), .B(n23842), .Z(n23844) );
  XOR U24464 ( .A(n23845), .B(n23844), .Z(n23719) );
  XNOR U24465 ( .A(n23718), .B(n23719), .Z(n23720) );
  XNOR U24466 ( .A(n23721), .B(n23720), .Z(n23725) );
  NANDN U24467 ( .A(n23682), .B(n23681), .Z(n23686) );
  NAND U24468 ( .A(n23684), .B(n23683), .Z(n23685) );
  NAND U24469 ( .A(n23686), .B(n23685), .Z(n23722) );
  NANDN U24470 ( .A(n23688), .B(n23687), .Z(n23692) );
  NAND U24471 ( .A(n23690), .B(n23689), .Z(n23691) );
  NAND U24472 ( .A(n23692), .B(n23691), .Z(n23723) );
  XNOR U24473 ( .A(n23722), .B(n23723), .Z(n23724) );
  XNOR U24474 ( .A(n23725), .B(n23724), .Z(n23715) );
  NANDN U24475 ( .A(n23698), .B(n23697), .Z(n23702) );
  NANDN U24476 ( .A(n23700), .B(n23699), .Z(n23701) );
  NAND U24477 ( .A(n23702), .B(n23701), .Z(n23713) );
  XNOR U24478 ( .A(n23712), .B(n23713), .Z(n23714) );
  XNOR U24479 ( .A(n23715), .B(n23714), .Z(n23708) );
  XOR U24480 ( .A(n23709), .B(n23708), .Z(n23710) );
  XNOR U24481 ( .A(n23711), .B(n23710), .Z(n23848) );
  XNOR U24482 ( .A(n23848), .B(sreg[395]), .Z(n23850) );
  NAND U24483 ( .A(n23703), .B(sreg[394]), .Z(n23707) );
  OR U24484 ( .A(n23705), .B(n23704), .Z(n23706) );
  AND U24485 ( .A(n23707), .B(n23706), .Z(n23849) );
  XOR U24486 ( .A(n23850), .B(n23849), .Z(c[395]) );
  NANDN U24487 ( .A(n23713), .B(n23712), .Z(n23717) );
  NANDN U24488 ( .A(n23715), .B(n23714), .Z(n23716) );
  NAND U24489 ( .A(n23717), .B(n23716), .Z(n23854) );
  NANDN U24490 ( .A(n23723), .B(n23722), .Z(n23727) );
  NANDN U24491 ( .A(n23725), .B(n23724), .Z(n23726) );
  NAND U24492 ( .A(n23727), .B(n23726), .Z(n23860) );
  XNOR U24493 ( .A(n23859), .B(n23860), .Z(n23861) );
  OR U24494 ( .A(n23729), .B(n23728), .Z(n23733) );
  NANDN U24495 ( .A(n23731), .B(n23730), .Z(n23732) );
  NAND U24496 ( .A(n23733), .B(n23732), .Z(n23977) );
  OR U24497 ( .A(n23735), .B(n23734), .Z(n23739) );
  NAND U24498 ( .A(n23737), .B(n23736), .Z(n23738) );
  NAND U24499 ( .A(n23739), .B(n23738), .Z(n23915) );
  OR U24500 ( .A(n23741), .B(n23740), .Z(n23745) );
  NANDN U24501 ( .A(n23743), .B(n23742), .Z(n23744) );
  NAND U24502 ( .A(n23745), .B(n23744), .Z(n23914) );
  OR U24503 ( .A(n23747), .B(n23746), .Z(n23751) );
  NANDN U24504 ( .A(n23749), .B(n23748), .Z(n23750) );
  NAND U24505 ( .A(n23751), .B(n23750), .Z(n23913) );
  XOR U24506 ( .A(n23915), .B(n23916), .Z(n23975) );
  OR U24507 ( .A(n23753), .B(n23752), .Z(n23757) );
  NANDN U24508 ( .A(n23755), .B(n23754), .Z(n23756) );
  NAND U24509 ( .A(n23757), .B(n23756), .Z(n23927) );
  XOR U24510 ( .A(b[19]), .B(n25862), .Z(n23871) );
  NANDN U24511 ( .A(n23871), .B(n37934), .Z(n23760) );
  NANDN U24512 ( .A(n23758), .B(n37935), .Z(n23759) );
  NAND U24513 ( .A(n23760), .B(n23759), .Z(n23940) );
  XOR U24514 ( .A(b[27]), .B(a[146]), .Z(n23874) );
  NAND U24515 ( .A(n38423), .B(n23874), .Z(n23763) );
  NANDN U24516 ( .A(n23761), .B(n38424), .Z(n23762) );
  NAND U24517 ( .A(n23763), .B(n23762), .Z(n23937) );
  XNOR U24518 ( .A(b[5]), .B(a[168]), .Z(n23877) );
  NANDN U24519 ( .A(n23877), .B(n36587), .Z(n23766) );
  NANDN U24520 ( .A(n23764), .B(n36588), .Z(n23765) );
  AND U24521 ( .A(n23766), .B(n23765), .Z(n23938) );
  XNOR U24522 ( .A(n23937), .B(n23938), .Z(n23939) );
  XNOR U24523 ( .A(n23940), .B(n23939), .Z(n23926) );
  NAND U24524 ( .A(n23767), .B(n37762), .Z(n23769) );
  XOR U24525 ( .A(b[17]), .B(a[156]), .Z(n23880) );
  NAND U24526 ( .A(n23880), .B(n37764), .Z(n23768) );
  NAND U24527 ( .A(n23769), .B(n23768), .Z(n23898) );
  XOR U24528 ( .A(b[31]), .B(n24120), .Z(n23883) );
  NANDN U24529 ( .A(n23883), .B(n38552), .Z(n23772) );
  NANDN U24530 ( .A(n23770), .B(n38553), .Z(n23771) );
  NAND U24531 ( .A(n23772), .B(n23771), .Z(n23895) );
  OR U24532 ( .A(n23773), .B(n36105), .Z(n23775) );
  XNOR U24533 ( .A(b[3]), .B(a[170]), .Z(n23886) );
  NANDN U24534 ( .A(n23886), .B(n36107), .Z(n23774) );
  AND U24535 ( .A(n23775), .B(n23774), .Z(n23896) );
  XNOR U24536 ( .A(n23895), .B(n23896), .Z(n23897) );
  XOR U24537 ( .A(n23898), .B(n23897), .Z(n23925) );
  XOR U24538 ( .A(n23926), .B(n23925), .Z(n23928) );
  XOR U24539 ( .A(n23927), .B(n23928), .Z(n23974) );
  XOR U24540 ( .A(n23975), .B(n23974), .Z(n23976) );
  XNOR U24541 ( .A(n23977), .B(n23976), .Z(n23995) );
  OR U24542 ( .A(n23777), .B(n23776), .Z(n23781) );
  NAND U24543 ( .A(n23779), .B(n23778), .Z(n23780) );
  NAND U24544 ( .A(n23781), .B(n23780), .Z(n23993) );
  NANDN U24545 ( .A(n23783), .B(n23782), .Z(n23787) );
  NANDN U24546 ( .A(n23785), .B(n23784), .Z(n23786) );
  NAND U24547 ( .A(n23787), .B(n23786), .Z(n23982) );
  OR U24548 ( .A(n23789), .B(n23788), .Z(n23793) );
  NAND U24549 ( .A(n23791), .B(n23790), .Z(n23792) );
  NAND U24550 ( .A(n23793), .B(n23792), .Z(n23981) );
  NANDN U24551 ( .A(n23795), .B(n23794), .Z(n23799) );
  NAND U24552 ( .A(n23797), .B(n23796), .Z(n23798) );
  NAND U24553 ( .A(n23799), .B(n23798), .Z(n23919) );
  NANDN U24554 ( .A(n23801), .B(n23800), .Z(n23805) );
  NAND U24555 ( .A(n23803), .B(n23802), .Z(n23804) );
  AND U24556 ( .A(n23805), .B(n23804), .Z(n23920) );
  XNOR U24557 ( .A(n23919), .B(n23920), .Z(n23921) );
  XNOR U24558 ( .A(b[9]), .B(a[164]), .Z(n23943) );
  NANDN U24559 ( .A(n23943), .B(n36925), .Z(n23808) );
  NANDN U24560 ( .A(n23806), .B(n36926), .Z(n23807) );
  NAND U24561 ( .A(n23808), .B(n23807), .Z(n23903) );
  XNOR U24562 ( .A(b[15]), .B(a[158]), .Z(n23946) );
  OR U24563 ( .A(n23946), .B(n37665), .Z(n23811) );
  NANDN U24564 ( .A(n23809), .B(n37604), .Z(n23810) );
  AND U24565 ( .A(n23811), .B(n23810), .Z(n23901) );
  XOR U24566 ( .A(b[21]), .B(n25213), .Z(n23949) );
  NANDN U24567 ( .A(n23949), .B(n38101), .Z(n23814) );
  NANDN U24568 ( .A(n23812), .B(n38102), .Z(n23813) );
  AND U24569 ( .A(n23814), .B(n23813), .Z(n23902) );
  XOR U24570 ( .A(n23903), .B(n23904), .Z(n23892) );
  XNOR U24571 ( .A(b[11]), .B(a[162]), .Z(n23952) );
  OR U24572 ( .A(n23952), .B(n37311), .Z(n23817) );
  NANDN U24573 ( .A(n23815), .B(n37218), .Z(n23816) );
  NAND U24574 ( .A(n23817), .B(n23816), .Z(n23890) );
  XOR U24575 ( .A(n1053), .B(a[160]), .Z(n23955) );
  NANDN U24576 ( .A(n23955), .B(n37424), .Z(n23820) );
  NANDN U24577 ( .A(n23818), .B(n37425), .Z(n23819) );
  AND U24578 ( .A(n23820), .B(n23819), .Z(n23889) );
  XNOR U24579 ( .A(n23890), .B(n23889), .Z(n23891) );
  XOR U24580 ( .A(n23892), .B(n23891), .Z(n23909) );
  NAND U24581 ( .A(n23821), .B(n38490), .Z(n23823) );
  XNOR U24582 ( .A(b[29]), .B(a[144]), .Z(n23962) );
  OR U24583 ( .A(n23962), .B(n1048), .Z(n23822) );
  NAND U24584 ( .A(n23823), .B(n23822), .Z(n23865) );
  NANDN U24585 ( .A(n1059), .B(a[140]), .Z(n23866) );
  XNOR U24586 ( .A(n23865), .B(n23866), .Z(n23868) );
  NANDN U24587 ( .A(n1049), .B(a[172]), .Z(n23824) );
  XNOR U24588 ( .A(b[1]), .B(n23824), .Z(n23826) );
  NANDN U24589 ( .A(b[0]), .B(a[171]), .Z(n23825) );
  AND U24590 ( .A(n23826), .B(n23825), .Z(n23867) );
  XOR U24591 ( .A(n23868), .B(n23867), .Z(n23907) );
  NANDN U24592 ( .A(n23827), .B(n38205), .Z(n23829) );
  XNOR U24593 ( .A(b[23]), .B(a[150]), .Z(n23965) );
  OR U24594 ( .A(n23965), .B(n38268), .Z(n23828) );
  NAND U24595 ( .A(n23829), .B(n23828), .Z(n23934) );
  XOR U24596 ( .A(b[7]), .B(a[166]), .Z(n23968) );
  NAND U24597 ( .A(n23968), .B(n36701), .Z(n23832) );
  NAND U24598 ( .A(n23830), .B(n36702), .Z(n23831) );
  NAND U24599 ( .A(n23832), .B(n23831), .Z(n23931) );
  XOR U24600 ( .A(b[25]), .B(a[148]), .Z(n23971) );
  NAND U24601 ( .A(n23971), .B(n38325), .Z(n23835) );
  NAND U24602 ( .A(n23833), .B(n38326), .Z(n23834) );
  AND U24603 ( .A(n23835), .B(n23834), .Z(n23932) );
  XNOR U24604 ( .A(n23931), .B(n23932), .Z(n23933) );
  XNOR U24605 ( .A(n23934), .B(n23933), .Z(n23908) );
  XOR U24606 ( .A(n23907), .B(n23908), .Z(n23910) );
  XNOR U24607 ( .A(n23909), .B(n23910), .Z(n23922) );
  XNOR U24608 ( .A(n23921), .B(n23922), .Z(n23980) );
  XNOR U24609 ( .A(n23981), .B(n23980), .Z(n23983) );
  XNOR U24610 ( .A(n23982), .B(n23983), .Z(n23992) );
  XNOR U24611 ( .A(n23993), .B(n23992), .Z(n23994) );
  XOR U24612 ( .A(n23995), .B(n23994), .Z(n23989) );
  NANDN U24613 ( .A(n23837), .B(n23836), .Z(n23841) );
  NAND U24614 ( .A(n23839), .B(n23838), .Z(n23840) );
  NAND U24615 ( .A(n23841), .B(n23840), .Z(n23986) );
  NAND U24616 ( .A(n23843), .B(n23842), .Z(n23847) );
  NAND U24617 ( .A(n23845), .B(n23844), .Z(n23846) );
  NAND U24618 ( .A(n23847), .B(n23846), .Z(n23987) );
  XNOR U24619 ( .A(n23986), .B(n23987), .Z(n23988) );
  XOR U24620 ( .A(n23989), .B(n23988), .Z(n23862) );
  XOR U24621 ( .A(n23861), .B(n23862), .Z(n23853) );
  XOR U24622 ( .A(n23854), .B(n23853), .Z(n23855) );
  XNOR U24623 ( .A(n23856), .B(n23855), .Z(n23998) );
  XNOR U24624 ( .A(n23998), .B(sreg[396]), .Z(n24000) );
  NAND U24625 ( .A(n23848), .B(sreg[395]), .Z(n23852) );
  OR U24626 ( .A(n23850), .B(n23849), .Z(n23851) );
  AND U24627 ( .A(n23852), .B(n23851), .Z(n23999) );
  XOR U24628 ( .A(n24000), .B(n23999), .Z(c[396]) );
  NAND U24629 ( .A(n23854), .B(n23853), .Z(n23858) );
  NAND U24630 ( .A(n23856), .B(n23855), .Z(n23857) );
  NAND U24631 ( .A(n23858), .B(n23857), .Z(n24006) );
  NANDN U24632 ( .A(n23860), .B(n23859), .Z(n23864) );
  NAND U24633 ( .A(n23862), .B(n23861), .Z(n23863) );
  NAND U24634 ( .A(n23864), .B(n23863), .Z(n24004) );
  NANDN U24635 ( .A(n23866), .B(n23865), .Z(n23870) );
  NAND U24636 ( .A(n23868), .B(n23867), .Z(n23869) );
  NAND U24637 ( .A(n23870), .B(n23869), .Z(n24090) );
  XNOR U24638 ( .A(b[19]), .B(a[155]), .Z(n24057) );
  NANDN U24639 ( .A(n24057), .B(n37934), .Z(n23873) );
  NANDN U24640 ( .A(n23871), .B(n37935), .Z(n23872) );
  NAND U24641 ( .A(n23873), .B(n23872), .Z(n24102) );
  XOR U24642 ( .A(b[27]), .B(a[147]), .Z(n24060) );
  NAND U24643 ( .A(n38423), .B(n24060), .Z(n23876) );
  NAND U24644 ( .A(n23874), .B(n38424), .Z(n23875) );
  NAND U24645 ( .A(n23876), .B(n23875), .Z(n24099) );
  XNOR U24646 ( .A(b[5]), .B(a[169]), .Z(n24063) );
  NANDN U24647 ( .A(n24063), .B(n36587), .Z(n23879) );
  NANDN U24648 ( .A(n23877), .B(n36588), .Z(n23878) );
  AND U24649 ( .A(n23879), .B(n23878), .Z(n24100) );
  XNOR U24650 ( .A(n24099), .B(n24100), .Z(n24101) );
  XNOR U24651 ( .A(n24102), .B(n24101), .Z(n24087) );
  NAND U24652 ( .A(n23880), .B(n37762), .Z(n23882) );
  XOR U24653 ( .A(b[17]), .B(a[157]), .Z(n24066) );
  NAND U24654 ( .A(n24066), .B(n37764), .Z(n23881) );
  NAND U24655 ( .A(n23882), .B(n23881), .Z(n24041) );
  XNOR U24656 ( .A(b[31]), .B(a[143]), .Z(n24069) );
  NANDN U24657 ( .A(n24069), .B(n38552), .Z(n23885) );
  NANDN U24658 ( .A(n23883), .B(n38553), .Z(n23884) );
  AND U24659 ( .A(n23885), .B(n23884), .Z(n24039) );
  OR U24660 ( .A(n23886), .B(n36105), .Z(n23888) );
  XNOR U24661 ( .A(b[3]), .B(a[171]), .Z(n24072) );
  NANDN U24662 ( .A(n24072), .B(n36107), .Z(n23887) );
  AND U24663 ( .A(n23888), .B(n23887), .Z(n24040) );
  XOR U24664 ( .A(n24041), .B(n24042), .Z(n24088) );
  XOR U24665 ( .A(n24087), .B(n24088), .Z(n24089) );
  XNOR U24666 ( .A(n24090), .B(n24089), .Z(n24136) );
  NANDN U24667 ( .A(n23890), .B(n23889), .Z(n23894) );
  NAND U24668 ( .A(n23892), .B(n23891), .Z(n23893) );
  NAND U24669 ( .A(n23894), .B(n23893), .Z(n24078) );
  NANDN U24670 ( .A(n23896), .B(n23895), .Z(n23900) );
  NAND U24671 ( .A(n23898), .B(n23897), .Z(n23899) );
  NAND U24672 ( .A(n23900), .B(n23899), .Z(n24076) );
  OR U24673 ( .A(n23902), .B(n23901), .Z(n23906) );
  NANDN U24674 ( .A(n23904), .B(n23903), .Z(n23905) );
  NAND U24675 ( .A(n23906), .B(n23905), .Z(n24075) );
  XNOR U24676 ( .A(n24078), .B(n24077), .Z(n24137) );
  XOR U24677 ( .A(n24136), .B(n24137), .Z(n24139) );
  NANDN U24678 ( .A(n23908), .B(n23907), .Z(n23912) );
  OR U24679 ( .A(n23910), .B(n23909), .Z(n23911) );
  NAND U24680 ( .A(n23912), .B(n23911), .Z(n24138) );
  XOR U24681 ( .A(n24139), .B(n24138), .Z(n24023) );
  OR U24682 ( .A(n23914), .B(n23913), .Z(n23918) );
  NANDN U24683 ( .A(n23916), .B(n23915), .Z(n23917) );
  NAND U24684 ( .A(n23918), .B(n23917), .Z(n24022) );
  NANDN U24685 ( .A(n23920), .B(n23919), .Z(n23924) );
  NANDN U24686 ( .A(n23922), .B(n23921), .Z(n23923) );
  NAND U24687 ( .A(n23924), .B(n23923), .Z(n24144) );
  NANDN U24688 ( .A(n23926), .B(n23925), .Z(n23930) );
  OR U24689 ( .A(n23928), .B(n23927), .Z(n23929) );
  NAND U24690 ( .A(n23930), .B(n23929), .Z(n24143) );
  NANDN U24691 ( .A(n23932), .B(n23931), .Z(n23936) );
  NAND U24692 ( .A(n23934), .B(n23933), .Z(n23935) );
  NAND U24693 ( .A(n23936), .B(n23935), .Z(n24081) );
  NANDN U24694 ( .A(n23938), .B(n23937), .Z(n23942) );
  NAND U24695 ( .A(n23940), .B(n23939), .Z(n23941) );
  AND U24696 ( .A(n23942), .B(n23941), .Z(n24082) );
  XNOR U24697 ( .A(n24081), .B(n24082), .Z(n24083) );
  XNOR U24698 ( .A(n1052), .B(a[165]), .Z(n24111) );
  NAND U24699 ( .A(n36925), .B(n24111), .Z(n23945) );
  NANDN U24700 ( .A(n23943), .B(n36926), .Z(n23944) );
  NAND U24701 ( .A(n23945), .B(n23944), .Z(n24047) );
  XNOR U24702 ( .A(b[15]), .B(a[159]), .Z(n24108) );
  OR U24703 ( .A(n24108), .B(n37665), .Z(n23948) );
  NANDN U24704 ( .A(n23946), .B(n37604), .Z(n23947) );
  AND U24705 ( .A(n23948), .B(n23947), .Z(n24045) );
  XNOR U24706 ( .A(n1056), .B(a[153]), .Z(n24105) );
  NAND U24707 ( .A(n24105), .B(n38101), .Z(n23951) );
  NANDN U24708 ( .A(n23949), .B(n38102), .Z(n23950) );
  AND U24709 ( .A(n23951), .B(n23950), .Z(n24046) );
  XOR U24710 ( .A(n24047), .B(n24048), .Z(n24036) );
  XOR U24711 ( .A(b[11]), .B(n27178), .Z(n24114) );
  OR U24712 ( .A(n24114), .B(n37311), .Z(n23954) );
  NANDN U24713 ( .A(n23952), .B(n37218), .Z(n23953) );
  NAND U24714 ( .A(n23954), .B(n23953), .Z(n24034) );
  XOR U24715 ( .A(n1053), .B(a[161]), .Z(n24117) );
  NANDN U24716 ( .A(n24117), .B(n37424), .Z(n23957) );
  NANDN U24717 ( .A(n23955), .B(n37425), .Z(n23956) );
  NAND U24718 ( .A(n23957), .B(n23956), .Z(n24033) );
  XOR U24719 ( .A(n24036), .B(n24035), .Z(n24030) );
  NANDN U24720 ( .A(n1049), .B(a[173]), .Z(n23958) );
  XNOR U24721 ( .A(b[1]), .B(n23958), .Z(n23960) );
  NANDN U24722 ( .A(b[0]), .B(a[172]), .Z(n23959) );
  AND U24723 ( .A(n23960), .B(n23959), .Z(n24054) );
  ANDN U24724 ( .B(b[31]), .A(n23961), .Z(n24051) );
  NANDN U24725 ( .A(n23962), .B(n38490), .Z(n23964) );
  XOR U24726 ( .A(b[29]), .B(n24554), .Z(n24121) );
  OR U24727 ( .A(n24121), .B(n1048), .Z(n23963) );
  NAND U24728 ( .A(n23964), .B(n23963), .Z(n24052) );
  XOR U24729 ( .A(n24051), .B(n24052), .Z(n24053) );
  XNOR U24730 ( .A(n24054), .B(n24053), .Z(n24027) );
  NANDN U24731 ( .A(n23965), .B(n38205), .Z(n23967) );
  XOR U24732 ( .A(b[23]), .B(n25435), .Z(n24127) );
  OR U24733 ( .A(n24127), .B(n38268), .Z(n23966) );
  NAND U24734 ( .A(n23967), .B(n23966), .Z(n24096) );
  XOR U24735 ( .A(b[7]), .B(a[167]), .Z(n24130) );
  NAND U24736 ( .A(n24130), .B(n36701), .Z(n23970) );
  NAND U24737 ( .A(n23968), .B(n36702), .Z(n23969) );
  NAND U24738 ( .A(n23970), .B(n23969), .Z(n24093) );
  XOR U24739 ( .A(b[25]), .B(a[149]), .Z(n24133) );
  NAND U24740 ( .A(n24133), .B(n38325), .Z(n23973) );
  NAND U24741 ( .A(n23971), .B(n38326), .Z(n23972) );
  AND U24742 ( .A(n23973), .B(n23972), .Z(n24094) );
  XNOR U24743 ( .A(n24093), .B(n24094), .Z(n24095) );
  XNOR U24744 ( .A(n24096), .B(n24095), .Z(n24028) );
  XOR U24745 ( .A(n24030), .B(n24029), .Z(n24084) );
  XNOR U24746 ( .A(n24083), .B(n24084), .Z(n24142) );
  XNOR U24747 ( .A(n24143), .B(n24142), .Z(n24145) );
  XNOR U24748 ( .A(n24144), .B(n24145), .Z(n24021) );
  XOR U24749 ( .A(n24022), .B(n24021), .Z(n24024) );
  NAND U24750 ( .A(n23975), .B(n23974), .Z(n23979) );
  NAND U24751 ( .A(n23977), .B(n23976), .Z(n23978) );
  NAND U24752 ( .A(n23979), .B(n23978), .Z(n24016) );
  NAND U24753 ( .A(n23981), .B(n23980), .Z(n23985) );
  NANDN U24754 ( .A(n23983), .B(n23982), .Z(n23984) );
  AND U24755 ( .A(n23985), .B(n23984), .Z(n24015) );
  XNOR U24756 ( .A(n24016), .B(n24015), .Z(n24017) );
  XOR U24757 ( .A(n24018), .B(n24017), .Z(n24011) );
  NANDN U24758 ( .A(n23987), .B(n23986), .Z(n23991) );
  NAND U24759 ( .A(n23989), .B(n23988), .Z(n23990) );
  NAND U24760 ( .A(n23991), .B(n23990), .Z(n24009) );
  NANDN U24761 ( .A(n23993), .B(n23992), .Z(n23997) );
  NANDN U24762 ( .A(n23995), .B(n23994), .Z(n23996) );
  NAND U24763 ( .A(n23997), .B(n23996), .Z(n24010) );
  XNOR U24764 ( .A(n24009), .B(n24010), .Z(n24012) );
  XOR U24765 ( .A(n24011), .B(n24012), .Z(n24003) );
  XOR U24766 ( .A(n24004), .B(n24003), .Z(n24005) );
  XNOR U24767 ( .A(n24006), .B(n24005), .Z(n24148) );
  XNOR U24768 ( .A(n24148), .B(sreg[397]), .Z(n24150) );
  NAND U24769 ( .A(n23998), .B(sreg[396]), .Z(n24002) );
  OR U24770 ( .A(n24000), .B(n23999), .Z(n24001) );
  AND U24771 ( .A(n24002), .B(n24001), .Z(n24149) );
  XOR U24772 ( .A(n24150), .B(n24149), .Z(c[397]) );
  NAND U24773 ( .A(n24004), .B(n24003), .Z(n24008) );
  NAND U24774 ( .A(n24006), .B(n24005), .Z(n24007) );
  NAND U24775 ( .A(n24008), .B(n24007), .Z(n24156) );
  NANDN U24776 ( .A(n24010), .B(n24009), .Z(n24014) );
  NAND U24777 ( .A(n24012), .B(n24011), .Z(n24013) );
  NAND U24778 ( .A(n24014), .B(n24013), .Z(n24154) );
  NANDN U24779 ( .A(n24016), .B(n24015), .Z(n24020) );
  NAND U24780 ( .A(n24018), .B(n24017), .Z(n24019) );
  NAND U24781 ( .A(n24020), .B(n24019), .Z(n24159) );
  NANDN U24782 ( .A(n24022), .B(n24021), .Z(n24026) );
  OR U24783 ( .A(n24024), .B(n24023), .Z(n24025) );
  NAND U24784 ( .A(n24026), .B(n24025), .Z(n24160) );
  XNOR U24785 ( .A(n24159), .B(n24160), .Z(n24161) );
  OR U24786 ( .A(n24028), .B(n24027), .Z(n24032) );
  NANDN U24787 ( .A(n24030), .B(n24029), .Z(n24031) );
  NAND U24788 ( .A(n24032), .B(n24031), .Z(n24274) );
  OR U24789 ( .A(n24034), .B(n24033), .Z(n24038) );
  NAND U24790 ( .A(n24036), .B(n24035), .Z(n24037) );
  NAND U24791 ( .A(n24038), .B(n24037), .Z(n24213) );
  OR U24792 ( .A(n24040), .B(n24039), .Z(n24044) );
  NANDN U24793 ( .A(n24042), .B(n24041), .Z(n24043) );
  NAND U24794 ( .A(n24044), .B(n24043), .Z(n24212) );
  OR U24795 ( .A(n24046), .B(n24045), .Z(n24050) );
  NANDN U24796 ( .A(n24048), .B(n24047), .Z(n24049) );
  NAND U24797 ( .A(n24050), .B(n24049), .Z(n24211) );
  XOR U24798 ( .A(n24213), .B(n24214), .Z(n24272) );
  OR U24799 ( .A(n24052), .B(n24051), .Z(n24056) );
  NANDN U24800 ( .A(n24054), .B(n24053), .Z(n24055) );
  NAND U24801 ( .A(n24056), .B(n24055), .Z(n24225) );
  XNOR U24802 ( .A(b[19]), .B(a[156]), .Z(n24171) );
  NANDN U24803 ( .A(n24171), .B(n37934), .Z(n24059) );
  NANDN U24804 ( .A(n24057), .B(n37935), .Z(n24058) );
  NAND U24805 ( .A(n24059), .B(n24058), .Z(n24238) );
  XOR U24806 ( .A(b[27]), .B(a[148]), .Z(n24174) );
  NAND U24807 ( .A(n38423), .B(n24174), .Z(n24062) );
  NAND U24808 ( .A(n24060), .B(n38424), .Z(n24061) );
  NAND U24809 ( .A(n24062), .B(n24061), .Z(n24235) );
  XNOR U24810 ( .A(b[5]), .B(a[170]), .Z(n24177) );
  NANDN U24811 ( .A(n24177), .B(n36587), .Z(n24065) );
  NANDN U24812 ( .A(n24063), .B(n36588), .Z(n24064) );
  AND U24813 ( .A(n24065), .B(n24064), .Z(n24236) );
  XNOR U24814 ( .A(n24235), .B(n24236), .Z(n24237) );
  XNOR U24815 ( .A(n24238), .B(n24237), .Z(n24224) );
  NAND U24816 ( .A(n24066), .B(n37762), .Z(n24068) );
  XOR U24817 ( .A(b[17]), .B(a[158]), .Z(n24180) );
  NAND U24818 ( .A(n24180), .B(n37764), .Z(n24067) );
  NAND U24819 ( .A(n24068), .B(n24067), .Z(n24198) );
  XNOR U24820 ( .A(b[31]), .B(a[144]), .Z(n24183) );
  NANDN U24821 ( .A(n24183), .B(n38552), .Z(n24071) );
  NANDN U24822 ( .A(n24069), .B(n38553), .Z(n24070) );
  NAND U24823 ( .A(n24071), .B(n24070), .Z(n24195) );
  OR U24824 ( .A(n24072), .B(n36105), .Z(n24074) );
  XNOR U24825 ( .A(b[3]), .B(a[172]), .Z(n24186) );
  NANDN U24826 ( .A(n24186), .B(n36107), .Z(n24073) );
  AND U24827 ( .A(n24074), .B(n24073), .Z(n24196) );
  XNOR U24828 ( .A(n24195), .B(n24196), .Z(n24197) );
  XOR U24829 ( .A(n24198), .B(n24197), .Z(n24223) );
  XOR U24830 ( .A(n24224), .B(n24223), .Z(n24226) );
  XOR U24831 ( .A(n24225), .B(n24226), .Z(n24271) );
  XOR U24832 ( .A(n24272), .B(n24271), .Z(n24273) );
  XNOR U24833 ( .A(n24274), .B(n24273), .Z(n24292) );
  OR U24834 ( .A(n24076), .B(n24075), .Z(n24080) );
  NAND U24835 ( .A(n24078), .B(n24077), .Z(n24079) );
  NAND U24836 ( .A(n24080), .B(n24079), .Z(n24290) );
  NANDN U24837 ( .A(n24082), .B(n24081), .Z(n24086) );
  NANDN U24838 ( .A(n24084), .B(n24083), .Z(n24085) );
  NAND U24839 ( .A(n24086), .B(n24085), .Z(n24279) );
  OR U24840 ( .A(n24088), .B(n24087), .Z(n24092) );
  NAND U24841 ( .A(n24090), .B(n24089), .Z(n24091) );
  NAND U24842 ( .A(n24092), .B(n24091), .Z(n24278) );
  NANDN U24843 ( .A(n24094), .B(n24093), .Z(n24098) );
  NAND U24844 ( .A(n24096), .B(n24095), .Z(n24097) );
  NAND U24845 ( .A(n24098), .B(n24097), .Z(n24217) );
  NANDN U24846 ( .A(n24100), .B(n24099), .Z(n24104) );
  NAND U24847 ( .A(n24102), .B(n24101), .Z(n24103) );
  AND U24848 ( .A(n24104), .B(n24103), .Z(n24218) );
  XNOR U24849 ( .A(n24217), .B(n24218), .Z(n24219) );
  XOR U24850 ( .A(n1056), .B(a[154]), .Z(n24247) );
  NANDN U24851 ( .A(n24247), .B(n38101), .Z(n24107) );
  NAND U24852 ( .A(n38102), .B(n24105), .Z(n24106) );
  NAND U24853 ( .A(n24107), .B(n24106), .Z(n24207) );
  XNOR U24854 ( .A(b[15]), .B(a[160]), .Z(n24244) );
  OR U24855 ( .A(n24244), .B(n37665), .Z(n24110) );
  NANDN U24856 ( .A(n24108), .B(n37604), .Z(n24109) );
  AND U24857 ( .A(n24110), .B(n24109), .Z(n24208) );
  XNOR U24858 ( .A(n24207), .B(n24208), .Z(n24210) );
  XOR U24859 ( .A(n1052), .B(a[166]), .Z(n24241) );
  NANDN U24860 ( .A(n24241), .B(n36925), .Z(n24113) );
  NAND U24861 ( .A(n36926), .B(n24111), .Z(n24112) );
  NAND U24862 ( .A(n24113), .B(n24112), .Z(n24209) );
  XNOR U24863 ( .A(n24210), .B(n24209), .Z(n24203) );
  XNOR U24864 ( .A(b[11]), .B(a[164]), .Z(n24250) );
  OR U24865 ( .A(n24250), .B(n37311), .Z(n24116) );
  NANDN U24866 ( .A(n24114), .B(n37218), .Z(n24115) );
  NAND U24867 ( .A(n24116), .B(n24115), .Z(n24202) );
  XOR U24868 ( .A(n1053), .B(a[162]), .Z(n24253) );
  NANDN U24869 ( .A(n24253), .B(n37424), .Z(n24119) );
  NANDN U24870 ( .A(n24117), .B(n37425), .Z(n24118) );
  NAND U24871 ( .A(n24119), .B(n24118), .Z(n24201) );
  XNOR U24872 ( .A(n24202), .B(n24201), .Z(n24204) );
  XNOR U24873 ( .A(n24203), .B(n24204), .Z(n24192) );
  ANDN U24874 ( .B(b[31]), .A(n24120), .Z(n24165) );
  NANDN U24875 ( .A(n24121), .B(n38490), .Z(n24123) );
  XNOR U24876 ( .A(n1058), .B(a[146]), .Z(n24259) );
  NANDN U24877 ( .A(n1048), .B(n24259), .Z(n24122) );
  NAND U24878 ( .A(n24123), .B(n24122), .Z(n24166) );
  XOR U24879 ( .A(n24165), .B(n24166), .Z(n24167) );
  NANDN U24880 ( .A(n1049), .B(a[174]), .Z(n24124) );
  XNOR U24881 ( .A(b[1]), .B(n24124), .Z(n24126) );
  NANDN U24882 ( .A(b[0]), .B(a[173]), .Z(n24125) );
  AND U24883 ( .A(n24126), .B(n24125), .Z(n24168) );
  XNOR U24884 ( .A(n24167), .B(n24168), .Z(n24189) );
  NANDN U24885 ( .A(n24127), .B(n38205), .Z(n24129) );
  XOR U24886 ( .A(b[23]), .B(n25213), .Z(n24262) );
  OR U24887 ( .A(n24262), .B(n38268), .Z(n24128) );
  NAND U24888 ( .A(n24129), .B(n24128), .Z(n24232) );
  XOR U24889 ( .A(b[7]), .B(a[168]), .Z(n24265) );
  NAND U24890 ( .A(n24265), .B(n36701), .Z(n24132) );
  NAND U24891 ( .A(n24130), .B(n36702), .Z(n24131) );
  NAND U24892 ( .A(n24132), .B(n24131), .Z(n24229) );
  XOR U24893 ( .A(b[25]), .B(a[150]), .Z(n24268) );
  NAND U24894 ( .A(n24268), .B(n38325), .Z(n24135) );
  NAND U24895 ( .A(n24133), .B(n38326), .Z(n24134) );
  AND U24896 ( .A(n24135), .B(n24134), .Z(n24230) );
  XNOR U24897 ( .A(n24229), .B(n24230), .Z(n24231) );
  XNOR U24898 ( .A(n24232), .B(n24231), .Z(n24190) );
  XOR U24899 ( .A(n24192), .B(n24191), .Z(n24220) );
  XNOR U24900 ( .A(n24219), .B(n24220), .Z(n24277) );
  XNOR U24901 ( .A(n24278), .B(n24277), .Z(n24280) );
  XNOR U24902 ( .A(n24279), .B(n24280), .Z(n24289) );
  XNOR U24903 ( .A(n24290), .B(n24289), .Z(n24291) );
  XOR U24904 ( .A(n24292), .B(n24291), .Z(n24286) );
  NANDN U24905 ( .A(n24137), .B(n24136), .Z(n24141) );
  OR U24906 ( .A(n24139), .B(n24138), .Z(n24140) );
  NAND U24907 ( .A(n24141), .B(n24140), .Z(n24283) );
  NAND U24908 ( .A(n24143), .B(n24142), .Z(n24147) );
  NANDN U24909 ( .A(n24145), .B(n24144), .Z(n24146) );
  NAND U24910 ( .A(n24147), .B(n24146), .Z(n24284) );
  XNOR U24911 ( .A(n24283), .B(n24284), .Z(n24285) );
  XOR U24912 ( .A(n24286), .B(n24285), .Z(n24162) );
  XOR U24913 ( .A(n24161), .B(n24162), .Z(n24153) );
  XOR U24914 ( .A(n24154), .B(n24153), .Z(n24155) );
  XNOR U24915 ( .A(n24156), .B(n24155), .Z(n24295) );
  XNOR U24916 ( .A(n24295), .B(sreg[398]), .Z(n24297) );
  NAND U24917 ( .A(n24148), .B(sreg[397]), .Z(n24152) );
  OR U24918 ( .A(n24150), .B(n24149), .Z(n24151) );
  AND U24919 ( .A(n24152), .B(n24151), .Z(n24296) );
  XOR U24920 ( .A(n24297), .B(n24296), .Z(c[398]) );
  NAND U24921 ( .A(n24154), .B(n24153), .Z(n24158) );
  NAND U24922 ( .A(n24156), .B(n24155), .Z(n24157) );
  NAND U24923 ( .A(n24158), .B(n24157), .Z(n24303) );
  NANDN U24924 ( .A(n24160), .B(n24159), .Z(n24164) );
  NAND U24925 ( .A(n24162), .B(n24161), .Z(n24163) );
  NAND U24926 ( .A(n24164), .B(n24163), .Z(n24301) );
  OR U24927 ( .A(n24166), .B(n24165), .Z(n24170) );
  NANDN U24928 ( .A(n24168), .B(n24167), .Z(n24169) );
  NAND U24929 ( .A(n24170), .B(n24169), .Z(n24370) );
  XNOR U24930 ( .A(b[19]), .B(a[157]), .Z(n24318) );
  NANDN U24931 ( .A(n24318), .B(n37934), .Z(n24173) );
  NANDN U24932 ( .A(n24171), .B(n37935), .Z(n24172) );
  NAND U24933 ( .A(n24173), .B(n24172), .Z(n24383) );
  XOR U24934 ( .A(b[27]), .B(a[149]), .Z(n24321) );
  NAND U24935 ( .A(n38423), .B(n24321), .Z(n24176) );
  NAND U24936 ( .A(n24174), .B(n38424), .Z(n24175) );
  NAND U24937 ( .A(n24176), .B(n24175), .Z(n24380) );
  XNOR U24938 ( .A(b[5]), .B(a[171]), .Z(n24324) );
  NANDN U24939 ( .A(n24324), .B(n36587), .Z(n24179) );
  NANDN U24940 ( .A(n24177), .B(n36588), .Z(n24178) );
  AND U24941 ( .A(n24179), .B(n24178), .Z(n24381) );
  XNOR U24942 ( .A(n24380), .B(n24381), .Z(n24382) );
  XNOR U24943 ( .A(n24383), .B(n24382), .Z(n24369) );
  NAND U24944 ( .A(n24180), .B(n37762), .Z(n24182) );
  XOR U24945 ( .A(b[17]), .B(a[159]), .Z(n24327) );
  NAND U24946 ( .A(n24327), .B(n37764), .Z(n24181) );
  NAND U24947 ( .A(n24182), .B(n24181), .Z(n24345) );
  XOR U24948 ( .A(b[31]), .B(n24554), .Z(n24330) );
  NANDN U24949 ( .A(n24330), .B(n38552), .Z(n24185) );
  NANDN U24950 ( .A(n24183), .B(n38553), .Z(n24184) );
  NAND U24951 ( .A(n24185), .B(n24184), .Z(n24342) );
  OR U24952 ( .A(n24186), .B(n36105), .Z(n24188) );
  XNOR U24953 ( .A(b[3]), .B(a[173]), .Z(n24333) );
  NANDN U24954 ( .A(n24333), .B(n36107), .Z(n24187) );
  AND U24955 ( .A(n24188), .B(n24187), .Z(n24343) );
  XNOR U24956 ( .A(n24342), .B(n24343), .Z(n24344) );
  XOR U24957 ( .A(n24345), .B(n24344), .Z(n24368) );
  XOR U24958 ( .A(n24369), .B(n24368), .Z(n24371) );
  XNOR U24959 ( .A(n24370), .B(n24371), .Z(n24422) );
  OR U24960 ( .A(n24190), .B(n24189), .Z(n24194) );
  NANDN U24961 ( .A(n24192), .B(n24191), .Z(n24193) );
  NAND U24962 ( .A(n24194), .B(n24193), .Z(n24423) );
  XNOR U24963 ( .A(n24422), .B(n24423), .Z(n24424) );
  NANDN U24964 ( .A(n24196), .B(n24195), .Z(n24200) );
  NAND U24965 ( .A(n24198), .B(n24197), .Z(n24199) );
  NAND U24966 ( .A(n24200), .B(n24199), .Z(n24361) );
  OR U24967 ( .A(n24202), .B(n24201), .Z(n24206) );
  NANDN U24968 ( .A(n24204), .B(n24203), .Z(n24205) );
  NAND U24969 ( .A(n24206), .B(n24205), .Z(n24359) );
  XNOR U24970 ( .A(n24359), .B(n24358), .Z(n24360) );
  XOR U24971 ( .A(n24361), .B(n24360), .Z(n24425) );
  XOR U24972 ( .A(n24424), .B(n24425), .Z(n24437) );
  OR U24973 ( .A(n24212), .B(n24211), .Z(n24216) );
  NANDN U24974 ( .A(n24214), .B(n24213), .Z(n24215) );
  NAND U24975 ( .A(n24216), .B(n24215), .Z(n24435) );
  NANDN U24976 ( .A(n24218), .B(n24217), .Z(n24222) );
  NANDN U24977 ( .A(n24220), .B(n24219), .Z(n24221) );
  NAND U24978 ( .A(n24222), .B(n24221), .Z(n24418) );
  NANDN U24979 ( .A(n24224), .B(n24223), .Z(n24228) );
  OR U24980 ( .A(n24226), .B(n24225), .Z(n24227) );
  NAND U24981 ( .A(n24228), .B(n24227), .Z(n24417) );
  NANDN U24982 ( .A(n24230), .B(n24229), .Z(n24234) );
  NAND U24983 ( .A(n24232), .B(n24231), .Z(n24233) );
  NAND U24984 ( .A(n24234), .B(n24233), .Z(n24362) );
  NANDN U24985 ( .A(n24236), .B(n24235), .Z(n24240) );
  NAND U24986 ( .A(n24238), .B(n24237), .Z(n24239) );
  AND U24987 ( .A(n24240), .B(n24239), .Z(n24363) );
  XNOR U24988 ( .A(n24362), .B(n24363), .Z(n24364) );
  XNOR U24989 ( .A(b[9]), .B(a[167]), .Z(n24386) );
  NANDN U24990 ( .A(n24386), .B(n36925), .Z(n24243) );
  NANDN U24991 ( .A(n24241), .B(n36926), .Z(n24242) );
  NAND U24992 ( .A(n24243), .B(n24242), .Z(n24350) );
  XNOR U24993 ( .A(n1054), .B(a[161]), .Z(n24389) );
  NANDN U24994 ( .A(n37665), .B(n24389), .Z(n24246) );
  NANDN U24995 ( .A(n24244), .B(n37604), .Z(n24245) );
  NAND U24996 ( .A(n24246), .B(n24245), .Z(n24348) );
  XNOR U24997 ( .A(b[21]), .B(a[155]), .Z(n24392) );
  NANDN U24998 ( .A(n24392), .B(n38101), .Z(n24249) );
  NANDN U24999 ( .A(n24247), .B(n38102), .Z(n24248) );
  NAND U25000 ( .A(n24249), .B(n24248), .Z(n24349) );
  XNOR U25001 ( .A(n24348), .B(n24349), .Z(n24351) );
  XOR U25002 ( .A(n24350), .B(n24351), .Z(n24339) );
  XNOR U25003 ( .A(b[11]), .B(a[165]), .Z(n24395) );
  OR U25004 ( .A(n24395), .B(n37311), .Z(n24252) );
  NANDN U25005 ( .A(n24250), .B(n37218), .Z(n24251) );
  NAND U25006 ( .A(n24252), .B(n24251), .Z(n24337) );
  XOR U25007 ( .A(n1053), .B(a[163]), .Z(n24398) );
  NANDN U25008 ( .A(n24398), .B(n37424), .Z(n24255) );
  NANDN U25009 ( .A(n24253), .B(n37425), .Z(n24254) );
  AND U25010 ( .A(n24255), .B(n24254), .Z(n24336) );
  XNOR U25011 ( .A(n24337), .B(n24336), .Z(n24338) );
  XNOR U25012 ( .A(n24339), .B(n24338), .Z(n24355) );
  NANDN U25013 ( .A(n1049), .B(a[175]), .Z(n24256) );
  XNOR U25014 ( .A(b[1]), .B(n24256), .Z(n24258) );
  NANDN U25015 ( .A(b[0]), .B(a[174]), .Z(n24257) );
  AND U25016 ( .A(n24258), .B(n24257), .Z(n24314) );
  NAND U25017 ( .A(n24259), .B(n38490), .Z(n24261) );
  XNOR U25018 ( .A(n1058), .B(a[147]), .Z(n24404) );
  NANDN U25019 ( .A(n1048), .B(n24404), .Z(n24260) );
  NAND U25020 ( .A(n24261), .B(n24260), .Z(n24312) );
  NANDN U25021 ( .A(n1059), .B(a[143]), .Z(n24313) );
  XNOR U25022 ( .A(n24312), .B(n24313), .Z(n24315) );
  XNOR U25023 ( .A(n24314), .B(n24315), .Z(n24353) );
  NANDN U25024 ( .A(n24262), .B(n38205), .Z(n24264) );
  XNOR U25025 ( .A(b[23]), .B(a[153]), .Z(n24407) );
  OR U25026 ( .A(n24407), .B(n38268), .Z(n24263) );
  NAND U25027 ( .A(n24264), .B(n24263), .Z(n24377) );
  XOR U25028 ( .A(b[7]), .B(a[169]), .Z(n24410) );
  NAND U25029 ( .A(n24410), .B(n36701), .Z(n24267) );
  NAND U25030 ( .A(n24265), .B(n36702), .Z(n24266) );
  NAND U25031 ( .A(n24267), .B(n24266), .Z(n24374) );
  XNOR U25032 ( .A(b[25]), .B(a[151]), .Z(n24413) );
  NANDN U25033 ( .A(n24413), .B(n38325), .Z(n24270) );
  NAND U25034 ( .A(n24268), .B(n38326), .Z(n24269) );
  AND U25035 ( .A(n24270), .B(n24269), .Z(n24375) );
  XNOR U25036 ( .A(n24374), .B(n24375), .Z(n24376) );
  XOR U25037 ( .A(n24377), .B(n24376), .Z(n24352) );
  XOR U25038 ( .A(n24355), .B(n24354), .Z(n24365) );
  XOR U25039 ( .A(n24364), .B(n24365), .Z(n24416) );
  XNOR U25040 ( .A(n24417), .B(n24416), .Z(n24419) );
  XNOR U25041 ( .A(n24418), .B(n24419), .Z(n24434) );
  XOR U25042 ( .A(n24435), .B(n24434), .Z(n24436) );
  XNOR U25043 ( .A(n24437), .B(n24436), .Z(n24431) );
  NAND U25044 ( .A(n24272), .B(n24271), .Z(n24276) );
  NAND U25045 ( .A(n24274), .B(n24273), .Z(n24275) );
  NAND U25046 ( .A(n24276), .B(n24275), .Z(n24429) );
  NAND U25047 ( .A(n24278), .B(n24277), .Z(n24282) );
  NANDN U25048 ( .A(n24280), .B(n24279), .Z(n24281) );
  AND U25049 ( .A(n24282), .B(n24281), .Z(n24428) );
  XNOR U25050 ( .A(n24429), .B(n24428), .Z(n24430) );
  XOR U25051 ( .A(n24431), .B(n24430), .Z(n24308) );
  NANDN U25052 ( .A(n24284), .B(n24283), .Z(n24288) );
  NAND U25053 ( .A(n24286), .B(n24285), .Z(n24287) );
  NAND U25054 ( .A(n24288), .B(n24287), .Z(n24306) );
  NANDN U25055 ( .A(n24290), .B(n24289), .Z(n24294) );
  NANDN U25056 ( .A(n24292), .B(n24291), .Z(n24293) );
  NAND U25057 ( .A(n24294), .B(n24293), .Z(n24307) );
  XNOR U25058 ( .A(n24306), .B(n24307), .Z(n24309) );
  XOR U25059 ( .A(n24308), .B(n24309), .Z(n24300) );
  XOR U25060 ( .A(n24301), .B(n24300), .Z(n24302) );
  XNOR U25061 ( .A(n24303), .B(n24302), .Z(n24440) );
  XNOR U25062 ( .A(n24440), .B(sreg[399]), .Z(n24442) );
  NAND U25063 ( .A(n24295), .B(sreg[398]), .Z(n24299) );
  OR U25064 ( .A(n24297), .B(n24296), .Z(n24298) );
  AND U25065 ( .A(n24299), .B(n24298), .Z(n24441) );
  XOR U25066 ( .A(n24442), .B(n24441), .Z(c[399]) );
  NAND U25067 ( .A(n24301), .B(n24300), .Z(n24305) );
  NAND U25068 ( .A(n24303), .B(n24302), .Z(n24304) );
  NAND U25069 ( .A(n24305), .B(n24304), .Z(n24448) );
  NANDN U25070 ( .A(n24307), .B(n24306), .Z(n24311) );
  NAND U25071 ( .A(n24309), .B(n24308), .Z(n24310) );
  NAND U25072 ( .A(n24311), .B(n24310), .Z(n24446) );
  NANDN U25073 ( .A(n24313), .B(n24312), .Z(n24317) );
  NAND U25074 ( .A(n24315), .B(n24314), .Z(n24316) );
  NAND U25075 ( .A(n24317), .B(n24316), .Z(n24526) );
  XNOR U25076 ( .A(b[19]), .B(a[158]), .Z(n24471) );
  NANDN U25077 ( .A(n24471), .B(n37934), .Z(n24320) );
  NANDN U25078 ( .A(n24318), .B(n37935), .Z(n24319) );
  NAND U25079 ( .A(n24320), .B(n24319), .Z(n24536) );
  XOR U25080 ( .A(b[27]), .B(a[150]), .Z(n24474) );
  NAND U25081 ( .A(n38423), .B(n24474), .Z(n24323) );
  NAND U25082 ( .A(n24321), .B(n38424), .Z(n24322) );
  NAND U25083 ( .A(n24323), .B(n24322), .Z(n24533) );
  XNOR U25084 ( .A(b[5]), .B(a[172]), .Z(n24477) );
  NANDN U25085 ( .A(n24477), .B(n36587), .Z(n24326) );
  NANDN U25086 ( .A(n24324), .B(n36588), .Z(n24325) );
  AND U25087 ( .A(n24326), .B(n24325), .Z(n24534) );
  XNOR U25088 ( .A(n24533), .B(n24534), .Z(n24535) );
  XNOR U25089 ( .A(n24536), .B(n24535), .Z(n24524) );
  NAND U25090 ( .A(n24327), .B(n37762), .Z(n24329) );
  XOR U25091 ( .A(b[17]), .B(a[160]), .Z(n24480) );
  NAND U25092 ( .A(n24480), .B(n37764), .Z(n24328) );
  NAND U25093 ( .A(n24329), .B(n24328), .Z(n24498) );
  XNOR U25094 ( .A(b[31]), .B(a[146]), .Z(n24483) );
  NANDN U25095 ( .A(n24483), .B(n38552), .Z(n24332) );
  NANDN U25096 ( .A(n24330), .B(n38553), .Z(n24331) );
  NAND U25097 ( .A(n24332), .B(n24331), .Z(n24495) );
  OR U25098 ( .A(n24333), .B(n36105), .Z(n24335) );
  XNOR U25099 ( .A(b[3]), .B(a[174]), .Z(n24486) );
  NANDN U25100 ( .A(n24486), .B(n36107), .Z(n24334) );
  AND U25101 ( .A(n24335), .B(n24334), .Z(n24496) );
  XNOR U25102 ( .A(n24495), .B(n24496), .Z(n24497) );
  XOR U25103 ( .A(n24498), .B(n24497), .Z(n24523) );
  XNOR U25104 ( .A(n24524), .B(n24523), .Z(n24525) );
  XNOR U25105 ( .A(n24526), .B(n24525), .Z(n24462) );
  NANDN U25106 ( .A(n24337), .B(n24336), .Z(n24341) );
  NAND U25107 ( .A(n24339), .B(n24338), .Z(n24340) );
  NAND U25108 ( .A(n24341), .B(n24340), .Z(n24515) );
  NANDN U25109 ( .A(n24343), .B(n24342), .Z(n24347) );
  NAND U25110 ( .A(n24345), .B(n24344), .Z(n24346) );
  NAND U25111 ( .A(n24347), .B(n24346), .Z(n24514) );
  XNOR U25112 ( .A(n24514), .B(n24513), .Z(n24516) );
  XOR U25113 ( .A(n24515), .B(n24516), .Z(n24461) );
  XOR U25114 ( .A(n24462), .B(n24461), .Z(n24463) );
  NANDN U25115 ( .A(n24353), .B(n24352), .Z(n24357) );
  NAND U25116 ( .A(n24355), .B(n24354), .Z(n24356) );
  AND U25117 ( .A(n24357), .B(n24356), .Z(n24464) );
  XNOR U25118 ( .A(n24463), .B(n24464), .Z(n24573) );
  NANDN U25119 ( .A(n24363), .B(n24362), .Z(n24367) );
  NAND U25120 ( .A(n24365), .B(n24364), .Z(n24366) );
  NAND U25121 ( .A(n24367), .B(n24366), .Z(n24458) );
  NANDN U25122 ( .A(n24369), .B(n24368), .Z(n24373) );
  OR U25123 ( .A(n24371), .B(n24370), .Z(n24372) );
  NAND U25124 ( .A(n24373), .B(n24372), .Z(n24455) );
  NANDN U25125 ( .A(n24375), .B(n24374), .Z(n24379) );
  NAND U25126 ( .A(n24377), .B(n24376), .Z(n24378) );
  NAND U25127 ( .A(n24379), .B(n24378), .Z(n24517) );
  NANDN U25128 ( .A(n24381), .B(n24380), .Z(n24385) );
  NAND U25129 ( .A(n24383), .B(n24382), .Z(n24384) );
  AND U25130 ( .A(n24385), .B(n24384), .Z(n24518) );
  XNOR U25131 ( .A(n24517), .B(n24518), .Z(n24519) );
  XNOR U25132 ( .A(b[9]), .B(a[168]), .Z(n24539) );
  NANDN U25133 ( .A(n24539), .B(n36925), .Z(n24388) );
  NANDN U25134 ( .A(n24386), .B(n36926), .Z(n24387) );
  NAND U25135 ( .A(n24388), .B(n24387), .Z(n24509) );
  XNOR U25136 ( .A(b[15]), .B(a[162]), .Z(n24542) );
  OR U25137 ( .A(n24542), .B(n37665), .Z(n24391) );
  NAND U25138 ( .A(n24389), .B(n37604), .Z(n24390) );
  AND U25139 ( .A(n24391), .B(n24390), .Z(n24507) );
  XNOR U25140 ( .A(b[21]), .B(a[156]), .Z(n24545) );
  NANDN U25141 ( .A(n24545), .B(n38101), .Z(n24394) );
  NANDN U25142 ( .A(n24392), .B(n38102), .Z(n24393) );
  AND U25143 ( .A(n24394), .B(n24393), .Z(n24508) );
  XOR U25144 ( .A(n24509), .B(n24510), .Z(n24504) );
  XNOR U25145 ( .A(b[11]), .B(a[166]), .Z(n24548) );
  OR U25146 ( .A(n24548), .B(n37311), .Z(n24397) );
  NANDN U25147 ( .A(n24395), .B(n37218), .Z(n24396) );
  NAND U25148 ( .A(n24397), .B(n24396), .Z(n24502) );
  XOR U25149 ( .A(n1053), .B(a[164]), .Z(n24551) );
  NANDN U25150 ( .A(n24551), .B(n37424), .Z(n24400) );
  NANDN U25151 ( .A(n24398), .B(n37425), .Z(n24399) );
  AND U25152 ( .A(n24400), .B(n24399), .Z(n24501) );
  XNOR U25153 ( .A(n24502), .B(n24501), .Z(n24503) );
  XOR U25154 ( .A(n24504), .B(n24503), .Z(n24491) );
  NANDN U25155 ( .A(n1049), .B(a[176]), .Z(n24401) );
  XNOR U25156 ( .A(b[1]), .B(n24401), .Z(n24403) );
  NANDN U25157 ( .A(b[0]), .B(a[175]), .Z(n24402) );
  AND U25158 ( .A(n24403), .B(n24402), .Z(n24467) );
  NAND U25159 ( .A(n38490), .B(n24404), .Z(n24406) );
  XNOR U25160 ( .A(b[29]), .B(a[148]), .Z(n24555) );
  OR U25161 ( .A(n24555), .B(n1048), .Z(n24405) );
  NAND U25162 ( .A(n24406), .B(n24405), .Z(n24465) );
  NANDN U25163 ( .A(n1059), .B(a[144]), .Z(n24466) );
  XNOR U25164 ( .A(n24465), .B(n24466), .Z(n24468) );
  XOR U25165 ( .A(n24467), .B(n24468), .Z(n24489) );
  NANDN U25166 ( .A(n24407), .B(n38205), .Z(n24409) );
  XOR U25167 ( .A(b[23]), .B(n25862), .Z(n24561) );
  OR U25168 ( .A(n24561), .B(n38268), .Z(n24408) );
  NAND U25169 ( .A(n24409), .B(n24408), .Z(n24530) );
  XOR U25170 ( .A(b[7]), .B(a[170]), .Z(n24564) );
  NAND U25171 ( .A(n24564), .B(n36701), .Z(n24412) );
  NAND U25172 ( .A(n24410), .B(n36702), .Z(n24411) );
  NAND U25173 ( .A(n24412), .B(n24411), .Z(n24527) );
  XNOR U25174 ( .A(b[25]), .B(a[152]), .Z(n24567) );
  NANDN U25175 ( .A(n24567), .B(n38325), .Z(n24415) );
  NANDN U25176 ( .A(n24413), .B(n38326), .Z(n24414) );
  AND U25177 ( .A(n24415), .B(n24414), .Z(n24528) );
  XNOR U25178 ( .A(n24527), .B(n24528), .Z(n24529) );
  XNOR U25179 ( .A(n24530), .B(n24529), .Z(n24490) );
  XOR U25180 ( .A(n24489), .B(n24490), .Z(n24492) );
  XNOR U25181 ( .A(n24491), .B(n24492), .Z(n24520) );
  XOR U25182 ( .A(n24519), .B(n24520), .Z(n24456) );
  XNOR U25183 ( .A(n24455), .B(n24456), .Z(n24457) );
  XOR U25184 ( .A(n24458), .B(n24457), .Z(n24571) );
  XNOR U25185 ( .A(n24570), .B(n24571), .Z(n24572) );
  XNOR U25186 ( .A(n24573), .B(n24572), .Z(n24577) );
  NAND U25187 ( .A(n24417), .B(n24416), .Z(n24421) );
  NANDN U25188 ( .A(n24419), .B(n24418), .Z(n24420) );
  NAND U25189 ( .A(n24421), .B(n24420), .Z(n24574) );
  NANDN U25190 ( .A(n24423), .B(n24422), .Z(n24427) );
  NAND U25191 ( .A(n24425), .B(n24424), .Z(n24426) );
  NAND U25192 ( .A(n24427), .B(n24426), .Z(n24575) );
  XNOR U25193 ( .A(n24574), .B(n24575), .Z(n24576) );
  XNOR U25194 ( .A(n24577), .B(n24576), .Z(n24452) );
  NANDN U25195 ( .A(n24429), .B(n24428), .Z(n24433) );
  NAND U25196 ( .A(n24431), .B(n24430), .Z(n24432) );
  NAND U25197 ( .A(n24433), .B(n24432), .Z(n24449) );
  NANDN U25198 ( .A(n24435), .B(n24434), .Z(n24439) );
  OR U25199 ( .A(n24437), .B(n24436), .Z(n24438) );
  NAND U25200 ( .A(n24439), .B(n24438), .Z(n24450) );
  XNOR U25201 ( .A(n24449), .B(n24450), .Z(n24451) );
  XNOR U25202 ( .A(n24452), .B(n24451), .Z(n24445) );
  XOR U25203 ( .A(n24446), .B(n24445), .Z(n24447) );
  XNOR U25204 ( .A(n24448), .B(n24447), .Z(n24580) );
  XNOR U25205 ( .A(n24580), .B(sreg[400]), .Z(n24582) );
  NAND U25206 ( .A(n24440), .B(sreg[399]), .Z(n24444) );
  OR U25207 ( .A(n24442), .B(n24441), .Z(n24443) );
  AND U25208 ( .A(n24444), .B(n24443), .Z(n24581) );
  XOR U25209 ( .A(n24582), .B(n24581), .Z(c[400]) );
  NANDN U25210 ( .A(n24450), .B(n24449), .Z(n24454) );
  NANDN U25211 ( .A(n24452), .B(n24451), .Z(n24453) );
  NAND U25212 ( .A(n24454), .B(n24453), .Z(n24585) );
  NANDN U25213 ( .A(n24456), .B(n24455), .Z(n24460) );
  NAND U25214 ( .A(n24458), .B(n24457), .Z(n24459) );
  NAND U25215 ( .A(n24460), .B(n24459), .Z(n24717) );
  XNOR U25216 ( .A(n24717), .B(n24718), .Z(n24719) );
  NANDN U25217 ( .A(n24466), .B(n24465), .Z(n24470) );
  NAND U25218 ( .A(n24468), .B(n24467), .Z(n24469) );
  NAND U25219 ( .A(n24470), .B(n24469), .Z(n24672) );
  XNOR U25220 ( .A(b[19]), .B(a[159]), .Z(n24639) );
  NANDN U25221 ( .A(n24639), .B(n37934), .Z(n24473) );
  NANDN U25222 ( .A(n24471), .B(n37935), .Z(n24472) );
  NAND U25223 ( .A(n24473), .B(n24472), .Z(n24684) );
  XNOR U25224 ( .A(b[27]), .B(a[151]), .Z(n24642) );
  NANDN U25225 ( .A(n24642), .B(n38423), .Z(n24476) );
  NAND U25226 ( .A(n24474), .B(n38424), .Z(n24475) );
  NAND U25227 ( .A(n24476), .B(n24475), .Z(n24681) );
  XNOR U25228 ( .A(b[5]), .B(a[173]), .Z(n24645) );
  NANDN U25229 ( .A(n24645), .B(n36587), .Z(n24479) );
  NANDN U25230 ( .A(n24477), .B(n36588), .Z(n24478) );
  AND U25231 ( .A(n24479), .B(n24478), .Z(n24682) );
  XNOR U25232 ( .A(n24681), .B(n24682), .Z(n24683) );
  XNOR U25233 ( .A(n24684), .B(n24683), .Z(n24669) );
  NAND U25234 ( .A(n24480), .B(n37762), .Z(n24482) );
  XNOR U25235 ( .A(b[17]), .B(a[161]), .Z(n24648) );
  NANDN U25236 ( .A(n24648), .B(n37764), .Z(n24481) );
  NAND U25237 ( .A(n24482), .B(n24481), .Z(n24623) );
  XNOR U25238 ( .A(b[31]), .B(a[147]), .Z(n24651) );
  NANDN U25239 ( .A(n24651), .B(n38552), .Z(n24485) );
  NANDN U25240 ( .A(n24483), .B(n38553), .Z(n24484) );
  AND U25241 ( .A(n24485), .B(n24484), .Z(n24621) );
  OR U25242 ( .A(n24486), .B(n36105), .Z(n24488) );
  XNOR U25243 ( .A(b[3]), .B(a[175]), .Z(n24654) );
  NANDN U25244 ( .A(n24654), .B(n36107), .Z(n24487) );
  AND U25245 ( .A(n24488), .B(n24487), .Z(n24622) );
  XOR U25246 ( .A(n24623), .B(n24624), .Z(n24670) );
  XOR U25247 ( .A(n24669), .B(n24670), .Z(n24671) );
  XNOR U25248 ( .A(n24672), .B(n24671), .Z(n24597) );
  NANDN U25249 ( .A(n24490), .B(n24489), .Z(n24494) );
  OR U25250 ( .A(n24492), .B(n24491), .Z(n24493) );
  NAND U25251 ( .A(n24494), .B(n24493), .Z(n24598) );
  XNOR U25252 ( .A(n24597), .B(n24598), .Z(n24599) );
  NANDN U25253 ( .A(n24496), .B(n24495), .Z(n24500) );
  NAND U25254 ( .A(n24498), .B(n24497), .Z(n24499) );
  NAND U25255 ( .A(n24500), .B(n24499), .Z(n24660) );
  NANDN U25256 ( .A(n24502), .B(n24501), .Z(n24506) );
  NAND U25257 ( .A(n24504), .B(n24503), .Z(n24505) );
  NAND U25258 ( .A(n24506), .B(n24505), .Z(n24657) );
  OR U25259 ( .A(n24508), .B(n24507), .Z(n24512) );
  NANDN U25260 ( .A(n24510), .B(n24509), .Z(n24511) );
  NAND U25261 ( .A(n24512), .B(n24511), .Z(n24658) );
  XNOR U25262 ( .A(n24657), .B(n24658), .Z(n24659) );
  XOR U25263 ( .A(n24660), .B(n24659), .Z(n24600) );
  XNOR U25264 ( .A(n24599), .B(n24600), .Z(n24725) );
  NANDN U25265 ( .A(n24518), .B(n24517), .Z(n24522) );
  NANDN U25266 ( .A(n24520), .B(n24519), .Z(n24521) );
  NAND U25267 ( .A(n24522), .B(n24521), .Z(n24606) );
  NANDN U25268 ( .A(n24528), .B(n24527), .Z(n24532) );
  NAND U25269 ( .A(n24530), .B(n24529), .Z(n24531) );
  NAND U25270 ( .A(n24532), .B(n24531), .Z(n24663) );
  NANDN U25271 ( .A(n24534), .B(n24533), .Z(n24538) );
  NAND U25272 ( .A(n24536), .B(n24535), .Z(n24537) );
  AND U25273 ( .A(n24538), .B(n24537), .Z(n24664) );
  XNOR U25274 ( .A(n24663), .B(n24664), .Z(n24665) );
  XNOR U25275 ( .A(b[9]), .B(a[169]), .Z(n24687) );
  NANDN U25276 ( .A(n24687), .B(n36925), .Z(n24541) );
  NANDN U25277 ( .A(n24539), .B(n36926), .Z(n24540) );
  NAND U25278 ( .A(n24541), .B(n24540), .Z(n24629) );
  XOR U25279 ( .A(b[15]), .B(n27178), .Z(n24690) );
  OR U25280 ( .A(n24690), .B(n37665), .Z(n24544) );
  NANDN U25281 ( .A(n24542), .B(n37604), .Z(n24543) );
  AND U25282 ( .A(n24544), .B(n24543), .Z(n24627) );
  XNOR U25283 ( .A(b[21]), .B(a[157]), .Z(n24693) );
  NANDN U25284 ( .A(n24693), .B(n38101), .Z(n24547) );
  NANDN U25285 ( .A(n24545), .B(n38102), .Z(n24546) );
  AND U25286 ( .A(n24547), .B(n24546), .Z(n24628) );
  XOR U25287 ( .A(n24629), .B(n24630), .Z(n24618) );
  XNOR U25288 ( .A(b[11]), .B(a[167]), .Z(n24696) );
  OR U25289 ( .A(n24696), .B(n37311), .Z(n24550) );
  NANDN U25290 ( .A(n24548), .B(n37218), .Z(n24549) );
  NAND U25291 ( .A(n24550), .B(n24549), .Z(n24616) );
  XOR U25292 ( .A(n1053), .B(a[165]), .Z(n24699) );
  NANDN U25293 ( .A(n24699), .B(n37424), .Z(n24553) );
  NANDN U25294 ( .A(n24551), .B(n37425), .Z(n24552) );
  NAND U25295 ( .A(n24553), .B(n24552), .Z(n24615) );
  XOR U25296 ( .A(n24618), .B(n24617), .Z(n24612) );
  ANDN U25297 ( .B(b[31]), .A(n24554), .Z(n24633) );
  NANDN U25298 ( .A(n24555), .B(n38490), .Z(n24557) );
  XNOR U25299 ( .A(n1058), .B(a[149]), .Z(n24705) );
  NANDN U25300 ( .A(n1048), .B(n24705), .Z(n24556) );
  NAND U25301 ( .A(n24557), .B(n24556), .Z(n24634) );
  XOR U25302 ( .A(n24633), .B(n24634), .Z(n24635) );
  NANDN U25303 ( .A(n1049), .B(a[177]), .Z(n24558) );
  XNOR U25304 ( .A(b[1]), .B(n24558), .Z(n24560) );
  NANDN U25305 ( .A(b[0]), .B(a[176]), .Z(n24559) );
  AND U25306 ( .A(n24560), .B(n24559), .Z(n24636) );
  XNOR U25307 ( .A(n24635), .B(n24636), .Z(n24609) );
  NANDN U25308 ( .A(n24561), .B(n38205), .Z(n24563) );
  XNOR U25309 ( .A(b[23]), .B(a[155]), .Z(n24708) );
  OR U25310 ( .A(n24708), .B(n38268), .Z(n24562) );
  NAND U25311 ( .A(n24563), .B(n24562), .Z(n24678) );
  XOR U25312 ( .A(b[7]), .B(a[171]), .Z(n24711) );
  NAND U25313 ( .A(n24711), .B(n36701), .Z(n24566) );
  NAND U25314 ( .A(n24564), .B(n36702), .Z(n24565) );
  NAND U25315 ( .A(n24566), .B(n24565), .Z(n24675) );
  XOR U25316 ( .A(b[25]), .B(a[153]), .Z(n24714) );
  NAND U25317 ( .A(n24714), .B(n38325), .Z(n24569) );
  NANDN U25318 ( .A(n24567), .B(n38326), .Z(n24568) );
  AND U25319 ( .A(n24569), .B(n24568), .Z(n24676) );
  XNOR U25320 ( .A(n24675), .B(n24676), .Z(n24677) );
  XNOR U25321 ( .A(n24678), .B(n24677), .Z(n24610) );
  XOR U25322 ( .A(n24612), .B(n24611), .Z(n24666) );
  XNOR U25323 ( .A(n24665), .B(n24666), .Z(n24603) );
  XOR U25324 ( .A(n24604), .B(n24603), .Z(n24605) );
  XNOR U25325 ( .A(n24606), .B(n24605), .Z(n24723) );
  XNOR U25326 ( .A(n24724), .B(n24723), .Z(n24726) );
  XNOR U25327 ( .A(n24725), .B(n24726), .Z(n24720) );
  XOR U25328 ( .A(n24719), .B(n24720), .Z(n24594) );
  NANDN U25329 ( .A(n24575), .B(n24574), .Z(n24579) );
  NANDN U25330 ( .A(n24577), .B(n24576), .Z(n24578) );
  NAND U25331 ( .A(n24579), .B(n24578), .Z(n24592) );
  XNOR U25332 ( .A(n24591), .B(n24592), .Z(n24593) );
  XNOR U25333 ( .A(n24594), .B(n24593), .Z(n24586) );
  XNOR U25334 ( .A(n24585), .B(n24586), .Z(n24587) );
  XNOR U25335 ( .A(n24588), .B(n24587), .Z(n24729) );
  XNOR U25336 ( .A(n24729), .B(sreg[401]), .Z(n24731) );
  NAND U25337 ( .A(n24580), .B(sreg[400]), .Z(n24584) );
  OR U25338 ( .A(n24582), .B(n24581), .Z(n24583) );
  AND U25339 ( .A(n24584), .B(n24583), .Z(n24730) );
  XOR U25340 ( .A(n24731), .B(n24730), .Z(c[401]) );
  NANDN U25341 ( .A(n24586), .B(n24585), .Z(n24590) );
  NAND U25342 ( .A(n24588), .B(n24587), .Z(n24589) );
  NAND U25343 ( .A(n24590), .B(n24589), .Z(n24737) );
  NANDN U25344 ( .A(n24592), .B(n24591), .Z(n24596) );
  NAND U25345 ( .A(n24594), .B(n24593), .Z(n24595) );
  NAND U25346 ( .A(n24596), .B(n24595), .Z(n24735) );
  NANDN U25347 ( .A(n24598), .B(n24597), .Z(n24602) );
  NANDN U25348 ( .A(n24600), .B(n24599), .Z(n24601) );
  NAND U25349 ( .A(n24602), .B(n24601), .Z(n24870) );
  NAND U25350 ( .A(n24604), .B(n24603), .Z(n24608) );
  NAND U25351 ( .A(n24606), .B(n24605), .Z(n24607) );
  NAND U25352 ( .A(n24608), .B(n24607), .Z(n24871) );
  XNOR U25353 ( .A(n24870), .B(n24871), .Z(n24872) );
  OR U25354 ( .A(n24610), .B(n24609), .Z(n24614) );
  NANDN U25355 ( .A(n24612), .B(n24611), .Z(n24613) );
  NAND U25356 ( .A(n24614), .B(n24613), .Z(n24857) );
  OR U25357 ( .A(n24616), .B(n24615), .Z(n24620) );
  NAND U25358 ( .A(n24618), .B(n24617), .Z(n24619) );
  NAND U25359 ( .A(n24620), .B(n24619), .Z(n24796) );
  OR U25360 ( .A(n24622), .B(n24621), .Z(n24626) );
  NANDN U25361 ( .A(n24624), .B(n24623), .Z(n24625) );
  NAND U25362 ( .A(n24626), .B(n24625), .Z(n24795) );
  OR U25363 ( .A(n24628), .B(n24627), .Z(n24632) );
  NANDN U25364 ( .A(n24630), .B(n24629), .Z(n24631) );
  NAND U25365 ( .A(n24632), .B(n24631), .Z(n24794) );
  XOR U25366 ( .A(n24796), .B(n24797), .Z(n24855) );
  OR U25367 ( .A(n24634), .B(n24633), .Z(n24638) );
  NANDN U25368 ( .A(n24636), .B(n24635), .Z(n24637) );
  NAND U25369 ( .A(n24638), .B(n24637), .Z(n24809) );
  XNOR U25370 ( .A(b[19]), .B(a[160]), .Z(n24776) );
  NANDN U25371 ( .A(n24776), .B(n37934), .Z(n24641) );
  NANDN U25372 ( .A(n24639), .B(n37935), .Z(n24640) );
  NAND U25373 ( .A(n24641), .B(n24640), .Z(n24821) );
  XNOR U25374 ( .A(b[27]), .B(a[152]), .Z(n24779) );
  NANDN U25375 ( .A(n24779), .B(n38423), .Z(n24644) );
  NANDN U25376 ( .A(n24642), .B(n38424), .Z(n24643) );
  NAND U25377 ( .A(n24644), .B(n24643), .Z(n24818) );
  XNOR U25378 ( .A(b[5]), .B(a[174]), .Z(n24782) );
  NANDN U25379 ( .A(n24782), .B(n36587), .Z(n24647) );
  NANDN U25380 ( .A(n24645), .B(n36588), .Z(n24646) );
  AND U25381 ( .A(n24647), .B(n24646), .Z(n24819) );
  XNOR U25382 ( .A(n24818), .B(n24819), .Z(n24820) );
  XNOR U25383 ( .A(n24821), .B(n24820), .Z(n24806) );
  NANDN U25384 ( .A(n24648), .B(n37762), .Z(n24650) );
  XOR U25385 ( .A(b[17]), .B(a[162]), .Z(n24785) );
  NAND U25386 ( .A(n24785), .B(n37764), .Z(n24649) );
  NAND U25387 ( .A(n24650), .B(n24649), .Z(n24760) );
  XNOR U25388 ( .A(b[31]), .B(a[148]), .Z(n24788) );
  NANDN U25389 ( .A(n24788), .B(n38552), .Z(n24653) );
  NANDN U25390 ( .A(n24651), .B(n38553), .Z(n24652) );
  AND U25391 ( .A(n24653), .B(n24652), .Z(n24758) );
  OR U25392 ( .A(n24654), .B(n36105), .Z(n24656) );
  XNOR U25393 ( .A(b[3]), .B(a[176]), .Z(n24791) );
  NANDN U25394 ( .A(n24791), .B(n36107), .Z(n24655) );
  AND U25395 ( .A(n24656), .B(n24655), .Z(n24759) );
  XOR U25396 ( .A(n24760), .B(n24761), .Z(n24807) );
  XOR U25397 ( .A(n24806), .B(n24807), .Z(n24808) );
  XNOR U25398 ( .A(n24809), .B(n24808), .Z(n24854) );
  XOR U25399 ( .A(n24855), .B(n24854), .Z(n24856) );
  XNOR U25400 ( .A(n24857), .B(n24856), .Z(n24867) );
  NANDN U25401 ( .A(n24658), .B(n24657), .Z(n24662) );
  NANDN U25402 ( .A(n24660), .B(n24659), .Z(n24661) );
  NAND U25403 ( .A(n24662), .B(n24661), .Z(n24864) );
  NANDN U25404 ( .A(n24664), .B(n24663), .Z(n24668) );
  NANDN U25405 ( .A(n24666), .B(n24665), .Z(n24667) );
  NAND U25406 ( .A(n24668), .B(n24667), .Z(n24861) );
  OR U25407 ( .A(n24670), .B(n24669), .Z(n24674) );
  NAND U25408 ( .A(n24672), .B(n24671), .Z(n24673) );
  NAND U25409 ( .A(n24674), .B(n24673), .Z(n24859) );
  NANDN U25410 ( .A(n24676), .B(n24675), .Z(n24680) );
  NAND U25411 ( .A(n24678), .B(n24677), .Z(n24679) );
  NAND U25412 ( .A(n24680), .B(n24679), .Z(n24800) );
  NANDN U25413 ( .A(n24682), .B(n24681), .Z(n24686) );
  NAND U25414 ( .A(n24684), .B(n24683), .Z(n24685) );
  AND U25415 ( .A(n24686), .B(n24685), .Z(n24801) );
  XNOR U25416 ( .A(n24800), .B(n24801), .Z(n24802) );
  XNOR U25417 ( .A(b[9]), .B(a[170]), .Z(n24824) );
  NANDN U25418 ( .A(n24824), .B(n36925), .Z(n24689) );
  NANDN U25419 ( .A(n24687), .B(n36926), .Z(n24688) );
  NAND U25420 ( .A(n24689), .B(n24688), .Z(n24766) );
  XNOR U25421 ( .A(b[15]), .B(a[164]), .Z(n24827) );
  OR U25422 ( .A(n24827), .B(n37665), .Z(n24692) );
  NANDN U25423 ( .A(n24690), .B(n37604), .Z(n24691) );
  AND U25424 ( .A(n24692), .B(n24691), .Z(n24764) );
  XNOR U25425 ( .A(b[21]), .B(a[158]), .Z(n24830) );
  NANDN U25426 ( .A(n24830), .B(n38101), .Z(n24695) );
  NANDN U25427 ( .A(n24693), .B(n38102), .Z(n24694) );
  AND U25428 ( .A(n24695), .B(n24694), .Z(n24765) );
  XOR U25429 ( .A(n24766), .B(n24767), .Z(n24755) );
  XNOR U25430 ( .A(b[11]), .B(a[168]), .Z(n24833) );
  OR U25431 ( .A(n24833), .B(n37311), .Z(n24698) );
  NANDN U25432 ( .A(n24696), .B(n37218), .Z(n24697) );
  NAND U25433 ( .A(n24698), .B(n24697), .Z(n24753) );
  XOR U25434 ( .A(n1053), .B(a[166]), .Z(n24836) );
  NANDN U25435 ( .A(n24836), .B(n37424), .Z(n24701) );
  NANDN U25436 ( .A(n24699), .B(n37425), .Z(n24700) );
  NAND U25437 ( .A(n24701), .B(n24700), .Z(n24752) );
  XOR U25438 ( .A(n24755), .B(n24754), .Z(n24749) );
  NANDN U25439 ( .A(n1049), .B(a[178]), .Z(n24702) );
  XNOR U25440 ( .A(b[1]), .B(n24702), .Z(n24704) );
  NANDN U25441 ( .A(b[0]), .B(a[177]), .Z(n24703) );
  AND U25442 ( .A(n24704), .B(n24703), .Z(n24772) );
  NAND U25443 ( .A(n24705), .B(n38490), .Z(n24707) );
  XNOR U25444 ( .A(n1058), .B(a[150]), .Z(n24839) );
  NANDN U25445 ( .A(n1048), .B(n24839), .Z(n24706) );
  NAND U25446 ( .A(n24707), .B(n24706), .Z(n24770) );
  NANDN U25447 ( .A(n1059), .B(a[146]), .Z(n24771) );
  XNOR U25448 ( .A(n24770), .B(n24771), .Z(n24773) );
  XNOR U25449 ( .A(n24772), .B(n24773), .Z(n24747) );
  NANDN U25450 ( .A(n24708), .B(n38205), .Z(n24710) );
  XNOR U25451 ( .A(b[23]), .B(a[156]), .Z(n24845) );
  OR U25452 ( .A(n24845), .B(n38268), .Z(n24709) );
  NAND U25453 ( .A(n24710), .B(n24709), .Z(n24815) );
  XOR U25454 ( .A(b[7]), .B(a[172]), .Z(n24848) );
  NAND U25455 ( .A(n24848), .B(n36701), .Z(n24713) );
  NAND U25456 ( .A(n24711), .B(n36702), .Z(n24712) );
  NAND U25457 ( .A(n24713), .B(n24712), .Z(n24812) );
  XNOR U25458 ( .A(b[25]), .B(a[154]), .Z(n24851) );
  NANDN U25459 ( .A(n24851), .B(n38325), .Z(n24716) );
  NAND U25460 ( .A(n24714), .B(n38326), .Z(n24715) );
  AND U25461 ( .A(n24716), .B(n24715), .Z(n24813) );
  XNOR U25462 ( .A(n24812), .B(n24813), .Z(n24814) );
  XOR U25463 ( .A(n24815), .B(n24814), .Z(n24746) );
  XOR U25464 ( .A(n24749), .B(n24748), .Z(n24803) );
  XNOR U25465 ( .A(n24802), .B(n24803), .Z(n24858) );
  XOR U25466 ( .A(n24859), .B(n24858), .Z(n24860) );
  XOR U25467 ( .A(n24861), .B(n24860), .Z(n24865) );
  XNOR U25468 ( .A(n24864), .B(n24865), .Z(n24866) );
  XOR U25469 ( .A(n24867), .B(n24866), .Z(n24873) );
  XOR U25470 ( .A(n24872), .B(n24873), .Z(n24742) );
  NANDN U25471 ( .A(n24718), .B(n24717), .Z(n24722) );
  NANDN U25472 ( .A(n24720), .B(n24719), .Z(n24721) );
  NAND U25473 ( .A(n24722), .B(n24721), .Z(n24741) );
  OR U25474 ( .A(n24724), .B(n24723), .Z(n24728) );
  OR U25475 ( .A(n24726), .B(n24725), .Z(n24727) );
  AND U25476 ( .A(n24728), .B(n24727), .Z(n24740) );
  XNOR U25477 ( .A(n24741), .B(n24740), .Z(n24743) );
  XOR U25478 ( .A(n24742), .B(n24743), .Z(n24734) );
  XOR U25479 ( .A(n24735), .B(n24734), .Z(n24736) );
  XNOR U25480 ( .A(n24737), .B(n24736), .Z(n24876) );
  XNOR U25481 ( .A(n24876), .B(sreg[402]), .Z(n24878) );
  NAND U25482 ( .A(n24729), .B(sreg[401]), .Z(n24733) );
  OR U25483 ( .A(n24731), .B(n24730), .Z(n24732) );
  AND U25484 ( .A(n24733), .B(n24732), .Z(n24877) );
  XOR U25485 ( .A(n24878), .B(n24877), .Z(c[402]) );
  NAND U25486 ( .A(n24735), .B(n24734), .Z(n24739) );
  NAND U25487 ( .A(n24737), .B(n24736), .Z(n24738) );
  NAND U25488 ( .A(n24739), .B(n24738), .Z(n24884) );
  NANDN U25489 ( .A(n24741), .B(n24740), .Z(n24745) );
  NAND U25490 ( .A(n24743), .B(n24742), .Z(n24744) );
  NAND U25491 ( .A(n24745), .B(n24744), .Z(n24882) );
  NANDN U25492 ( .A(n24747), .B(n24746), .Z(n24751) );
  NANDN U25493 ( .A(n24749), .B(n24748), .Z(n24750) );
  NAND U25494 ( .A(n24751), .B(n24750), .Z(n25002) );
  OR U25495 ( .A(n24753), .B(n24752), .Z(n24757) );
  NAND U25496 ( .A(n24755), .B(n24754), .Z(n24756) );
  NAND U25497 ( .A(n24757), .B(n24756), .Z(n24941) );
  OR U25498 ( .A(n24759), .B(n24758), .Z(n24763) );
  NANDN U25499 ( .A(n24761), .B(n24760), .Z(n24762) );
  NAND U25500 ( .A(n24763), .B(n24762), .Z(n24940) );
  OR U25501 ( .A(n24765), .B(n24764), .Z(n24769) );
  NANDN U25502 ( .A(n24767), .B(n24766), .Z(n24768) );
  NAND U25503 ( .A(n24769), .B(n24768), .Z(n24939) );
  XOR U25504 ( .A(n24941), .B(n24942), .Z(n24999) );
  NANDN U25505 ( .A(n24771), .B(n24770), .Z(n24775) );
  NAND U25506 ( .A(n24773), .B(n24772), .Z(n24774) );
  NAND U25507 ( .A(n24775), .B(n24774), .Z(n24954) );
  XOR U25508 ( .A(b[19]), .B(n26869), .Z(n24897) );
  NANDN U25509 ( .A(n24897), .B(n37934), .Z(n24778) );
  NANDN U25510 ( .A(n24776), .B(n37935), .Z(n24777) );
  NAND U25511 ( .A(n24778), .B(n24777), .Z(n24966) );
  XOR U25512 ( .A(b[27]), .B(a[153]), .Z(n24900) );
  NAND U25513 ( .A(n38423), .B(n24900), .Z(n24781) );
  NANDN U25514 ( .A(n24779), .B(n38424), .Z(n24780) );
  NAND U25515 ( .A(n24781), .B(n24780), .Z(n24963) );
  XNOR U25516 ( .A(b[5]), .B(a[175]), .Z(n24903) );
  NANDN U25517 ( .A(n24903), .B(n36587), .Z(n24784) );
  NANDN U25518 ( .A(n24782), .B(n36588), .Z(n24783) );
  AND U25519 ( .A(n24784), .B(n24783), .Z(n24964) );
  XNOR U25520 ( .A(n24963), .B(n24964), .Z(n24965) );
  XNOR U25521 ( .A(n24966), .B(n24965), .Z(n24952) );
  NAND U25522 ( .A(n24785), .B(n37762), .Z(n24787) );
  XNOR U25523 ( .A(b[17]), .B(a[163]), .Z(n24906) );
  NANDN U25524 ( .A(n24906), .B(n37764), .Z(n24786) );
  NAND U25525 ( .A(n24787), .B(n24786), .Z(n24924) );
  XNOR U25526 ( .A(b[31]), .B(a[149]), .Z(n24909) );
  NANDN U25527 ( .A(n24909), .B(n38552), .Z(n24790) );
  NANDN U25528 ( .A(n24788), .B(n38553), .Z(n24789) );
  NAND U25529 ( .A(n24790), .B(n24789), .Z(n24921) );
  OR U25530 ( .A(n24791), .B(n36105), .Z(n24793) );
  XNOR U25531 ( .A(b[3]), .B(a[177]), .Z(n24912) );
  NANDN U25532 ( .A(n24912), .B(n36107), .Z(n24792) );
  AND U25533 ( .A(n24793), .B(n24792), .Z(n24922) );
  XNOR U25534 ( .A(n24921), .B(n24922), .Z(n24923) );
  XOR U25535 ( .A(n24924), .B(n24923), .Z(n24951) );
  XNOR U25536 ( .A(n24952), .B(n24951), .Z(n24953) );
  XNOR U25537 ( .A(n24954), .B(n24953), .Z(n25000) );
  XNOR U25538 ( .A(n24999), .B(n25000), .Z(n25001) );
  XNOR U25539 ( .A(n25002), .B(n25001), .Z(n25020) );
  OR U25540 ( .A(n24795), .B(n24794), .Z(n24799) );
  NANDN U25541 ( .A(n24797), .B(n24796), .Z(n24798) );
  NAND U25542 ( .A(n24799), .B(n24798), .Z(n25018) );
  NANDN U25543 ( .A(n24801), .B(n24800), .Z(n24805) );
  NANDN U25544 ( .A(n24803), .B(n24802), .Z(n24804) );
  NAND U25545 ( .A(n24805), .B(n24804), .Z(n25007) );
  OR U25546 ( .A(n24807), .B(n24806), .Z(n24811) );
  NANDN U25547 ( .A(n24809), .B(n24808), .Z(n24810) );
  NAND U25548 ( .A(n24811), .B(n24810), .Z(n25006) );
  NANDN U25549 ( .A(n24813), .B(n24812), .Z(n24817) );
  NAND U25550 ( .A(n24815), .B(n24814), .Z(n24816) );
  NAND U25551 ( .A(n24817), .B(n24816), .Z(n24945) );
  NANDN U25552 ( .A(n24819), .B(n24818), .Z(n24823) );
  NAND U25553 ( .A(n24821), .B(n24820), .Z(n24822) );
  AND U25554 ( .A(n24823), .B(n24822), .Z(n24946) );
  XNOR U25555 ( .A(n24945), .B(n24946), .Z(n24947) );
  XNOR U25556 ( .A(n1052), .B(a[171]), .Z(n24969) );
  NAND U25557 ( .A(n36925), .B(n24969), .Z(n24826) );
  NANDN U25558 ( .A(n24824), .B(n36926), .Z(n24825) );
  NAND U25559 ( .A(n24826), .B(n24825), .Z(n24929) );
  XNOR U25560 ( .A(b[15]), .B(a[165]), .Z(n24972) );
  OR U25561 ( .A(n24972), .B(n37665), .Z(n24829) );
  NANDN U25562 ( .A(n24827), .B(n37604), .Z(n24828) );
  AND U25563 ( .A(n24829), .B(n24828), .Z(n24927) );
  XNOR U25564 ( .A(n1056), .B(a[159]), .Z(n24975) );
  NAND U25565 ( .A(n24975), .B(n38101), .Z(n24832) );
  NANDN U25566 ( .A(n24830), .B(n38102), .Z(n24831) );
  AND U25567 ( .A(n24832), .B(n24831), .Z(n24928) );
  XOR U25568 ( .A(n24929), .B(n24930), .Z(n24918) );
  XNOR U25569 ( .A(b[11]), .B(a[169]), .Z(n24978) );
  OR U25570 ( .A(n24978), .B(n37311), .Z(n24835) );
  NANDN U25571 ( .A(n24833), .B(n37218), .Z(n24834) );
  NAND U25572 ( .A(n24835), .B(n24834), .Z(n24916) );
  XOR U25573 ( .A(n1053), .B(a[167]), .Z(n24981) );
  NANDN U25574 ( .A(n24981), .B(n37424), .Z(n24838) );
  NANDN U25575 ( .A(n24836), .B(n37425), .Z(n24837) );
  AND U25576 ( .A(n24838), .B(n24837), .Z(n24915) );
  XNOR U25577 ( .A(n24916), .B(n24915), .Z(n24917) );
  XOR U25578 ( .A(n24918), .B(n24917), .Z(n24935) );
  NAND U25579 ( .A(n38490), .B(n24839), .Z(n24841) );
  XOR U25580 ( .A(n1058), .B(n25435), .Z(n24987) );
  NANDN U25581 ( .A(n1048), .B(n24987), .Z(n24840) );
  NAND U25582 ( .A(n24841), .B(n24840), .Z(n24891) );
  NANDN U25583 ( .A(n1059), .B(a[147]), .Z(n24892) );
  XNOR U25584 ( .A(n24891), .B(n24892), .Z(n24894) );
  NANDN U25585 ( .A(n1049), .B(a[179]), .Z(n24842) );
  XNOR U25586 ( .A(b[1]), .B(n24842), .Z(n24844) );
  NANDN U25587 ( .A(b[0]), .B(a[178]), .Z(n24843) );
  AND U25588 ( .A(n24844), .B(n24843), .Z(n24893) );
  XOR U25589 ( .A(n24894), .B(n24893), .Z(n24933) );
  NANDN U25590 ( .A(n24845), .B(n38205), .Z(n24847) );
  XNOR U25591 ( .A(b[23]), .B(a[157]), .Z(n24990) );
  OR U25592 ( .A(n24990), .B(n38268), .Z(n24846) );
  NAND U25593 ( .A(n24847), .B(n24846), .Z(n24960) );
  XOR U25594 ( .A(b[7]), .B(a[173]), .Z(n24993) );
  NAND U25595 ( .A(n24993), .B(n36701), .Z(n24850) );
  NAND U25596 ( .A(n24848), .B(n36702), .Z(n24849) );
  NAND U25597 ( .A(n24850), .B(n24849), .Z(n24957) );
  XOR U25598 ( .A(b[25]), .B(a[155]), .Z(n24996) );
  NAND U25599 ( .A(n24996), .B(n38325), .Z(n24853) );
  NANDN U25600 ( .A(n24851), .B(n38326), .Z(n24852) );
  AND U25601 ( .A(n24853), .B(n24852), .Z(n24958) );
  XNOR U25602 ( .A(n24957), .B(n24958), .Z(n24959) );
  XNOR U25603 ( .A(n24960), .B(n24959), .Z(n24934) );
  XOR U25604 ( .A(n24933), .B(n24934), .Z(n24936) );
  XNOR U25605 ( .A(n24935), .B(n24936), .Z(n24948) );
  XNOR U25606 ( .A(n24947), .B(n24948), .Z(n25005) );
  XNOR U25607 ( .A(n25006), .B(n25005), .Z(n25008) );
  XNOR U25608 ( .A(n25007), .B(n25008), .Z(n25017) );
  XNOR U25609 ( .A(n25018), .B(n25017), .Z(n25019) );
  XOR U25610 ( .A(n25020), .B(n25019), .Z(n25014) );
  NAND U25611 ( .A(n24859), .B(n24858), .Z(n24863) );
  NAND U25612 ( .A(n24861), .B(n24860), .Z(n24862) );
  AND U25613 ( .A(n24863), .B(n24862), .Z(n25011) );
  XNOR U25614 ( .A(n25012), .B(n25011), .Z(n25013) );
  XNOR U25615 ( .A(n25014), .B(n25013), .Z(n24888) );
  NANDN U25616 ( .A(n24865), .B(n24864), .Z(n24869) );
  NAND U25617 ( .A(n24867), .B(n24866), .Z(n24868) );
  NAND U25618 ( .A(n24869), .B(n24868), .Z(n24885) );
  NANDN U25619 ( .A(n24871), .B(n24870), .Z(n24875) );
  NAND U25620 ( .A(n24873), .B(n24872), .Z(n24874) );
  AND U25621 ( .A(n24875), .B(n24874), .Z(n24886) );
  XNOR U25622 ( .A(n24885), .B(n24886), .Z(n24887) );
  XNOR U25623 ( .A(n24888), .B(n24887), .Z(n24881) );
  XOR U25624 ( .A(n24882), .B(n24881), .Z(n24883) );
  XNOR U25625 ( .A(n24884), .B(n24883), .Z(n25023) );
  XNOR U25626 ( .A(n25023), .B(sreg[403]), .Z(n25025) );
  NAND U25627 ( .A(n24876), .B(sreg[402]), .Z(n24880) );
  OR U25628 ( .A(n24878), .B(n24877), .Z(n24879) );
  AND U25629 ( .A(n24880), .B(n24879), .Z(n25024) );
  XOR U25630 ( .A(n25025), .B(n25024), .Z(c[403]) );
  NANDN U25631 ( .A(n24886), .B(n24885), .Z(n24890) );
  NANDN U25632 ( .A(n24888), .B(n24887), .Z(n24889) );
  NAND U25633 ( .A(n24890), .B(n24889), .Z(n25029) );
  NANDN U25634 ( .A(n24892), .B(n24891), .Z(n24896) );
  NAND U25635 ( .A(n24894), .B(n24893), .Z(n24895) );
  NAND U25636 ( .A(n24896), .B(n24895), .Z(n25101) );
  XNOR U25637 ( .A(b[19]), .B(a[162]), .Z(n25046) );
  NANDN U25638 ( .A(n25046), .B(n37934), .Z(n24899) );
  NANDN U25639 ( .A(n24897), .B(n37935), .Z(n24898) );
  NAND U25640 ( .A(n24899), .B(n24898), .Z(n25111) );
  XNOR U25641 ( .A(b[27]), .B(a[154]), .Z(n25049) );
  NANDN U25642 ( .A(n25049), .B(n38423), .Z(n24902) );
  NAND U25643 ( .A(n24900), .B(n38424), .Z(n24901) );
  NAND U25644 ( .A(n24902), .B(n24901), .Z(n25108) );
  XNOR U25645 ( .A(b[5]), .B(a[176]), .Z(n25052) );
  NANDN U25646 ( .A(n25052), .B(n36587), .Z(n24905) );
  NANDN U25647 ( .A(n24903), .B(n36588), .Z(n24904) );
  AND U25648 ( .A(n24905), .B(n24904), .Z(n25109) );
  XNOR U25649 ( .A(n25108), .B(n25109), .Z(n25110) );
  XNOR U25650 ( .A(n25111), .B(n25110), .Z(n25099) );
  NANDN U25651 ( .A(n24906), .B(n37762), .Z(n24908) );
  XOR U25652 ( .A(b[17]), .B(a[164]), .Z(n25055) );
  NAND U25653 ( .A(n25055), .B(n37764), .Z(n24907) );
  NAND U25654 ( .A(n24908), .B(n24907), .Z(n25073) );
  XNOR U25655 ( .A(b[31]), .B(a[150]), .Z(n25058) );
  NANDN U25656 ( .A(n25058), .B(n38552), .Z(n24911) );
  NANDN U25657 ( .A(n24909), .B(n38553), .Z(n24910) );
  NAND U25658 ( .A(n24911), .B(n24910), .Z(n25070) );
  OR U25659 ( .A(n24912), .B(n36105), .Z(n24914) );
  XNOR U25660 ( .A(b[3]), .B(a[178]), .Z(n25061) );
  NANDN U25661 ( .A(n25061), .B(n36107), .Z(n24913) );
  AND U25662 ( .A(n24914), .B(n24913), .Z(n25071) );
  XNOR U25663 ( .A(n25070), .B(n25071), .Z(n25072) );
  XOR U25664 ( .A(n25073), .B(n25072), .Z(n25098) );
  XNOR U25665 ( .A(n25099), .B(n25098), .Z(n25100) );
  XNOR U25666 ( .A(n25101), .B(n25100), .Z(n25144) );
  NANDN U25667 ( .A(n24916), .B(n24915), .Z(n24920) );
  NAND U25668 ( .A(n24918), .B(n24917), .Z(n24919) );
  NAND U25669 ( .A(n24920), .B(n24919), .Z(n25089) );
  NANDN U25670 ( .A(n24922), .B(n24921), .Z(n24926) );
  NAND U25671 ( .A(n24924), .B(n24923), .Z(n24925) );
  NAND U25672 ( .A(n24926), .B(n24925), .Z(n25087) );
  OR U25673 ( .A(n24928), .B(n24927), .Z(n24932) );
  NANDN U25674 ( .A(n24930), .B(n24929), .Z(n24931) );
  NAND U25675 ( .A(n24932), .B(n24931), .Z(n25086) );
  XNOR U25676 ( .A(n25089), .B(n25088), .Z(n25145) );
  XOR U25677 ( .A(n25144), .B(n25145), .Z(n25147) );
  NANDN U25678 ( .A(n24934), .B(n24933), .Z(n24938) );
  OR U25679 ( .A(n24936), .B(n24935), .Z(n24937) );
  NAND U25680 ( .A(n24938), .B(n24937), .Z(n25146) );
  XOR U25681 ( .A(n25147), .B(n25146), .Z(n25164) );
  OR U25682 ( .A(n24940), .B(n24939), .Z(n24944) );
  NANDN U25683 ( .A(n24942), .B(n24941), .Z(n24943) );
  NAND U25684 ( .A(n24944), .B(n24943), .Z(n25163) );
  NANDN U25685 ( .A(n24946), .B(n24945), .Z(n24950) );
  NANDN U25686 ( .A(n24948), .B(n24947), .Z(n24949) );
  NAND U25687 ( .A(n24950), .B(n24949), .Z(n25152) );
  NANDN U25688 ( .A(n24952), .B(n24951), .Z(n24956) );
  NAND U25689 ( .A(n24954), .B(n24953), .Z(n24955) );
  NAND U25690 ( .A(n24956), .B(n24955), .Z(n25151) );
  NANDN U25691 ( .A(n24958), .B(n24957), .Z(n24962) );
  NAND U25692 ( .A(n24960), .B(n24959), .Z(n24961) );
  NAND U25693 ( .A(n24962), .B(n24961), .Z(n25092) );
  NANDN U25694 ( .A(n24964), .B(n24963), .Z(n24968) );
  NAND U25695 ( .A(n24966), .B(n24965), .Z(n24967) );
  AND U25696 ( .A(n24968), .B(n24967), .Z(n25093) );
  XNOR U25697 ( .A(n25092), .B(n25093), .Z(n25094) );
  XNOR U25698 ( .A(b[9]), .B(a[172]), .Z(n25114) );
  NANDN U25699 ( .A(n25114), .B(n36925), .Z(n24971) );
  NAND U25700 ( .A(n36926), .B(n24969), .Z(n24970) );
  NAND U25701 ( .A(n24971), .B(n24970), .Z(n25078) );
  XNOR U25702 ( .A(n1054), .B(a[166]), .Z(n25117) );
  NANDN U25703 ( .A(n37665), .B(n25117), .Z(n24974) );
  NANDN U25704 ( .A(n24972), .B(n37604), .Z(n24973) );
  NAND U25705 ( .A(n24974), .B(n24973), .Z(n25076) );
  XNOR U25706 ( .A(b[21]), .B(a[160]), .Z(n25120) );
  NANDN U25707 ( .A(n25120), .B(n38101), .Z(n24977) );
  NAND U25708 ( .A(n38102), .B(n24975), .Z(n24976) );
  NAND U25709 ( .A(n24977), .B(n24976), .Z(n25077) );
  XNOR U25710 ( .A(n25076), .B(n25077), .Z(n25079) );
  XOR U25711 ( .A(n25078), .B(n25079), .Z(n25067) );
  XNOR U25712 ( .A(b[11]), .B(a[170]), .Z(n25123) );
  OR U25713 ( .A(n25123), .B(n37311), .Z(n24980) );
  NANDN U25714 ( .A(n24978), .B(n37218), .Z(n24979) );
  NAND U25715 ( .A(n24980), .B(n24979), .Z(n25065) );
  XOR U25716 ( .A(n1053), .B(a[168]), .Z(n25126) );
  NANDN U25717 ( .A(n25126), .B(n37424), .Z(n24983) );
  NANDN U25718 ( .A(n24981), .B(n37425), .Z(n24982) );
  AND U25719 ( .A(n24983), .B(n24982), .Z(n25064) );
  XNOR U25720 ( .A(n25065), .B(n25064), .Z(n25066) );
  XNOR U25721 ( .A(n25067), .B(n25066), .Z(n25083) );
  NANDN U25722 ( .A(n1049), .B(a[180]), .Z(n24984) );
  XNOR U25723 ( .A(b[1]), .B(n24984), .Z(n24986) );
  NANDN U25724 ( .A(b[0]), .B(a[179]), .Z(n24985) );
  AND U25725 ( .A(n24986), .B(n24985), .Z(n25042) );
  NAND U25726 ( .A(n38490), .B(n24987), .Z(n24989) );
  XOR U25727 ( .A(n1058), .B(n25213), .Z(n25129) );
  NANDN U25728 ( .A(n1048), .B(n25129), .Z(n24988) );
  NAND U25729 ( .A(n24989), .B(n24988), .Z(n25040) );
  NANDN U25730 ( .A(n1059), .B(a[148]), .Z(n25041) );
  XNOR U25731 ( .A(n25040), .B(n25041), .Z(n25043) );
  XNOR U25732 ( .A(n25042), .B(n25043), .Z(n25081) );
  NANDN U25733 ( .A(n24990), .B(n38205), .Z(n24992) );
  XNOR U25734 ( .A(b[23]), .B(a[158]), .Z(n25135) );
  OR U25735 ( .A(n25135), .B(n38268), .Z(n24991) );
  NAND U25736 ( .A(n24992), .B(n24991), .Z(n25105) );
  XOR U25737 ( .A(b[7]), .B(a[174]), .Z(n25138) );
  NAND U25738 ( .A(n25138), .B(n36701), .Z(n24995) );
  NAND U25739 ( .A(n24993), .B(n36702), .Z(n24994) );
  NAND U25740 ( .A(n24995), .B(n24994), .Z(n25102) );
  XOR U25741 ( .A(b[25]), .B(a[156]), .Z(n25141) );
  NAND U25742 ( .A(n25141), .B(n38325), .Z(n24998) );
  NAND U25743 ( .A(n24996), .B(n38326), .Z(n24997) );
  AND U25744 ( .A(n24998), .B(n24997), .Z(n25103) );
  XNOR U25745 ( .A(n25102), .B(n25103), .Z(n25104) );
  XOR U25746 ( .A(n25105), .B(n25104), .Z(n25080) );
  XOR U25747 ( .A(n25083), .B(n25082), .Z(n25095) );
  XOR U25748 ( .A(n25094), .B(n25095), .Z(n25150) );
  XNOR U25749 ( .A(n25151), .B(n25150), .Z(n25153) );
  XNOR U25750 ( .A(n25152), .B(n25153), .Z(n25162) );
  XOR U25751 ( .A(n25163), .B(n25162), .Z(n25165) );
  NANDN U25752 ( .A(n25000), .B(n24999), .Z(n25004) );
  NAND U25753 ( .A(n25002), .B(n25001), .Z(n25003) );
  NAND U25754 ( .A(n25004), .B(n25003), .Z(n25157) );
  NAND U25755 ( .A(n25006), .B(n25005), .Z(n25010) );
  NANDN U25756 ( .A(n25008), .B(n25007), .Z(n25009) );
  AND U25757 ( .A(n25010), .B(n25009), .Z(n25156) );
  XNOR U25758 ( .A(n25157), .B(n25156), .Z(n25158) );
  XOR U25759 ( .A(n25159), .B(n25158), .Z(n25036) );
  NANDN U25760 ( .A(n25012), .B(n25011), .Z(n25016) );
  NAND U25761 ( .A(n25014), .B(n25013), .Z(n25015) );
  NAND U25762 ( .A(n25016), .B(n25015), .Z(n25034) );
  NANDN U25763 ( .A(n25018), .B(n25017), .Z(n25022) );
  NANDN U25764 ( .A(n25020), .B(n25019), .Z(n25021) );
  NAND U25765 ( .A(n25022), .B(n25021), .Z(n25035) );
  XNOR U25766 ( .A(n25034), .B(n25035), .Z(n25037) );
  XOR U25767 ( .A(n25036), .B(n25037), .Z(n25028) );
  XOR U25768 ( .A(n25029), .B(n25028), .Z(n25030) );
  XNOR U25769 ( .A(n25031), .B(n25030), .Z(n25168) );
  XNOR U25770 ( .A(n25168), .B(sreg[404]), .Z(n25170) );
  NAND U25771 ( .A(n25023), .B(sreg[403]), .Z(n25027) );
  OR U25772 ( .A(n25025), .B(n25024), .Z(n25026) );
  AND U25773 ( .A(n25027), .B(n25026), .Z(n25169) );
  XOR U25774 ( .A(n25170), .B(n25169), .Z(c[404]) );
  NAND U25775 ( .A(n25029), .B(n25028), .Z(n25033) );
  NAND U25776 ( .A(n25031), .B(n25030), .Z(n25032) );
  NAND U25777 ( .A(n25033), .B(n25032), .Z(n25176) );
  NANDN U25778 ( .A(n25035), .B(n25034), .Z(n25039) );
  NAND U25779 ( .A(n25037), .B(n25036), .Z(n25038) );
  NAND U25780 ( .A(n25039), .B(n25038), .Z(n25174) );
  NANDN U25781 ( .A(n25041), .B(n25040), .Z(n25045) );
  NAND U25782 ( .A(n25043), .B(n25042), .Z(n25044) );
  NAND U25783 ( .A(n25045), .B(n25044), .Z(n25257) );
  XOR U25784 ( .A(b[19]), .B(n27178), .Z(n25201) );
  NANDN U25785 ( .A(n25201), .B(n37934), .Z(n25048) );
  NANDN U25786 ( .A(n25046), .B(n37935), .Z(n25047) );
  NAND U25787 ( .A(n25048), .B(n25047), .Z(n25267) );
  XOR U25788 ( .A(b[27]), .B(a[155]), .Z(n25204) );
  NAND U25789 ( .A(n38423), .B(n25204), .Z(n25051) );
  NANDN U25790 ( .A(n25049), .B(n38424), .Z(n25050) );
  NAND U25791 ( .A(n25051), .B(n25050), .Z(n25264) );
  XNOR U25792 ( .A(b[5]), .B(a[177]), .Z(n25207) );
  NANDN U25793 ( .A(n25207), .B(n36587), .Z(n25054) );
  NANDN U25794 ( .A(n25052), .B(n36588), .Z(n25053) );
  AND U25795 ( .A(n25054), .B(n25053), .Z(n25265) );
  XNOR U25796 ( .A(n25264), .B(n25265), .Z(n25266) );
  XNOR U25797 ( .A(n25267), .B(n25266), .Z(n25255) );
  NAND U25798 ( .A(n25055), .B(n37762), .Z(n25057) );
  XOR U25799 ( .A(b[17]), .B(a[165]), .Z(n25210) );
  NAND U25800 ( .A(n25210), .B(n37764), .Z(n25056) );
  NAND U25801 ( .A(n25057), .B(n25056), .Z(n25229) );
  XOR U25802 ( .A(b[31]), .B(n25435), .Z(n25214) );
  NANDN U25803 ( .A(n25214), .B(n38552), .Z(n25060) );
  NANDN U25804 ( .A(n25058), .B(n38553), .Z(n25059) );
  NAND U25805 ( .A(n25060), .B(n25059), .Z(n25226) );
  OR U25806 ( .A(n25061), .B(n36105), .Z(n25063) );
  XNOR U25807 ( .A(b[3]), .B(a[179]), .Z(n25217) );
  NANDN U25808 ( .A(n25217), .B(n36107), .Z(n25062) );
  AND U25809 ( .A(n25063), .B(n25062), .Z(n25227) );
  XNOR U25810 ( .A(n25226), .B(n25227), .Z(n25228) );
  XOR U25811 ( .A(n25229), .B(n25228), .Z(n25254) );
  XNOR U25812 ( .A(n25255), .B(n25254), .Z(n25256) );
  XNOR U25813 ( .A(n25257), .B(n25256), .Z(n25192) );
  NANDN U25814 ( .A(n25065), .B(n25064), .Z(n25069) );
  NAND U25815 ( .A(n25067), .B(n25066), .Z(n25068) );
  NAND U25816 ( .A(n25069), .B(n25068), .Z(n25246) );
  NANDN U25817 ( .A(n25071), .B(n25070), .Z(n25075) );
  NAND U25818 ( .A(n25073), .B(n25072), .Z(n25074) );
  NAND U25819 ( .A(n25075), .B(n25074), .Z(n25245) );
  XNOR U25820 ( .A(n25245), .B(n25244), .Z(n25247) );
  XOR U25821 ( .A(n25246), .B(n25247), .Z(n25191) );
  XOR U25822 ( .A(n25192), .B(n25191), .Z(n25193) );
  NANDN U25823 ( .A(n25081), .B(n25080), .Z(n25085) );
  NAND U25824 ( .A(n25083), .B(n25082), .Z(n25084) );
  NAND U25825 ( .A(n25085), .B(n25084), .Z(n25194) );
  XNOR U25826 ( .A(n25193), .B(n25194), .Z(n25308) );
  OR U25827 ( .A(n25087), .B(n25086), .Z(n25091) );
  NAND U25828 ( .A(n25089), .B(n25088), .Z(n25090) );
  NAND U25829 ( .A(n25091), .B(n25090), .Z(n25307) );
  NANDN U25830 ( .A(n25093), .B(n25092), .Z(n25097) );
  NAND U25831 ( .A(n25095), .B(n25094), .Z(n25096) );
  NAND U25832 ( .A(n25097), .B(n25096), .Z(n25187) );
  NANDN U25833 ( .A(n25103), .B(n25102), .Z(n25107) );
  NAND U25834 ( .A(n25105), .B(n25104), .Z(n25106) );
  NAND U25835 ( .A(n25107), .B(n25106), .Z(n25248) );
  NANDN U25836 ( .A(n25109), .B(n25108), .Z(n25113) );
  NAND U25837 ( .A(n25111), .B(n25110), .Z(n25112) );
  AND U25838 ( .A(n25113), .B(n25112), .Z(n25249) );
  XNOR U25839 ( .A(n25248), .B(n25249), .Z(n25250) );
  XNOR U25840 ( .A(b[9]), .B(a[173]), .Z(n25270) );
  NANDN U25841 ( .A(n25270), .B(n36925), .Z(n25116) );
  NANDN U25842 ( .A(n25114), .B(n36926), .Z(n25115) );
  NAND U25843 ( .A(n25116), .B(n25115), .Z(n25234) );
  XNOR U25844 ( .A(b[15]), .B(a[167]), .Z(n25273) );
  OR U25845 ( .A(n25273), .B(n37665), .Z(n25119) );
  NAND U25846 ( .A(n25117), .B(n37604), .Z(n25118) );
  AND U25847 ( .A(n25119), .B(n25118), .Z(n25232) );
  XOR U25848 ( .A(b[21]), .B(n26869), .Z(n25276) );
  NANDN U25849 ( .A(n25276), .B(n38101), .Z(n25122) );
  NANDN U25850 ( .A(n25120), .B(n38102), .Z(n25121) );
  AND U25851 ( .A(n25122), .B(n25121), .Z(n25233) );
  XOR U25852 ( .A(n25234), .B(n25235), .Z(n25223) );
  XNOR U25853 ( .A(b[11]), .B(a[171]), .Z(n25279) );
  OR U25854 ( .A(n25279), .B(n37311), .Z(n25125) );
  NANDN U25855 ( .A(n25123), .B(n37218), .Z(n25124) );
  NAND U25856 ( .A(n25125), .B(n25124), .Z(n25221) );
  XOR U25857 ( .A(n1053), .B(a[169]), .Z(n25282) );
  NANDN U25858 ( .A(n25282), .B(n37424), .Z(n25128) );
  NANDN U25859 ( .A(n25126), .B(n37425), .Z(n25127) );
  AND U25860 ( .A(n25128), .B(n25127), .Z(n25220) );
  XNOR U25861 ( .A(n25221), .B(n25220), .Z(n25222) );
  XOR U25862 ( .A(n25223), .B(n25222), .Z(n25240) );
  NAND U25863 ( .A(n38490), .B(n25129), .Z(n25131) );
  XNOR U25864 ( .A(n1058), .B(a[153]), .Z(n25288) );
  NANDN U25865 ( .A(n1048), .B(n25288), .Z(n25130) );
  NAND U25866 ( .A(n25131), .B(n25130), .Z(n25195) );
  NANDN U25867 ( .A(n1059), .B(a[149]), .Z(n25196) );
  XNOR U25868 ( .A(n25195), .B(n25196), .Z(n25198) );
  NANDN U25869 ( .A(n1049), .B(a[181]), .Z(n25132) );
  XNOR U25870 ( .A(b[1]), .B(n25132), .Z(n25134) );
  NANDN U25871 ( .A(b[0]), .B(a[180]), .Z(n25133) );
  AND U25872 ( .A(n25134), .B(n25133), .Z(n25197) );
  XOR U25873 ( .A(n25198), .B(n25197), .Z(n25238) );
  NANDN U25874 ( .A(n25135), .B(n38205), .Z(n25137) );
  XNOR U25875 ( .A(b[23]), .B(a[159]), .Z(n25291) );
  OR U25876 ( .A(n25291), .B(n38268), .Z(n25136) );
  NAND U25877 ( .A(n25137), .B(n25136), .Z(n25261) );
  XOR U25878 ( .A(b[7]), .B(a[175]), .Z(n25294) );
  NAND U25879 ( .A(n25294), .B(n36701), .Z(n25140) );
  NAND U25880 ( .A(n25138), .B(n36702), .Z(n25139) );
  NAND U25881 ( .A(n25140), .B(n25139), .Z(n25258) );
  XOR U25882 ( .A(b[25]), .B(a[157]), .Z(n25297) );
  NAND U25883 ( .A(n25297), .B(n38325), .Z(n25143) );
  NAND U25884 ( .A(n25141), .B(n38326), .Z(n25142) );
  AND U25885 ( .A(n25143), .B(n25142), .Z(n25259) );
  XNOR U25886 ( .A(n25258), .B(n25259), .Z(n25260) );
  XNOR U25887 ( .A(n25261), .B(n25260), .Z(n25239) );
  XOR U25888 ( .A(n25238), .B(n25239), .Z(n25241) );
  XNOR U25889 ( .A(n25240), .B(n25241), .Z(n25251) );
  XNOR U25890 ( .A(n25250), .B(n25251), .Z(n25185) );
  XNOR U25891 ( .A(n25186), .B(n25185), .Z(n25188) );
  XNOR U25892 ( .A(n25187), .B(n25188), .Z(n25306) );
  XOR U25893 ( .A(n25307), .B(n25306), .Z(n25309) );
  NANDN U25894 ( .A(n25145), .B(n25144), .Z(n25149) );
  OR U25895 ( .A(n25147), .B(n25146), .Z(n25148) );
  NAND U25896 ( .A(n25149), .B(n25148), .Z(n25300) );
  NAND U25897 ( .A(n25151), .B(n25150), .Z(n25155) );
  NANDN U25898 ( .A(n25153), .B(n25152), .Z(n25154) );
  NAND U25899 ( .A(n25155), .B(n25154), .Z(n25301) );
  XNOR U25900 ( .A(n25300), .B(n25301), .Z(n25302) );
  XOR U25901 ( .A(n25303), .B(n25302), .Z(n25181) );
  NANDN U25902 ( .A(n25157), .B(n25156), .Z(n25161) );
  NAND U25903 ( .A(n25159), .B(n25158), .Z(n25160) );
  NAND U25904 ( .A(n25161), .B(n25160), .Z(n25179) );
  NANDN U25905 ( .A(n25163), .B(n25162), .Z(n25167) );
  OR U25906 ( .A(n25165), .B(n25164), .Z(n25166) );
  NAND U25907 ( .A(n25167), .B(n25166), .Z(n25180) );
  XNOR U25908 ( .A(n25179), .B(n25180), .Z(n25182) );
  XOR U25909 ( .A(n25181), .B(n25182), .Z(n25173) );
  XOR U25910 ( .A(n25174), .B(n25173), .Z(n25175) );
  XNOR U25911 ( .A(n25176), .B(n25175), .Z(n25312) );
  XNOR U25912 ( .A(n25312), .B(sreg[405]), .Z(n25314) );
  NAND U25913 ( .A(n25168), .B(sreg[404]), .Z(n25172) );
  OR U25914 ( .A(n25170), .B(n25169), .Z(n25171) );
  AND U25915 ( .A(n25172), .B(n25171), .Z(n25313) );
  XOR U25916 ( .A(n25314), .B(n25313), .Z(c[405]) );
  NAND U25917 ( .A(n25174), .B(n25173), .Z(n25178) );
  NAND U25918 ( .A(n25176), .B(n25175), .Z(n25177) );
  NAND U25919 ( .A(n25178), .B(n25177), .Z(n25320) );
  NANDN U25920 ( .A(n25180), .B(n25179), .Z(n25184) );
  NAND U25921 ( .A(n25182), .B(n25181), .Z(n25183) );
  NAND U25922 ( .A(n25184), .B(n25183), .Z(n25317) );
  NAND U25923 ( .A(n25186), .B(n25185), .Z(n25190) );
  NANDN U25924 ( .A(n25188), .B(n25187), .Z(n25189) );
  NAND U25925 ( .A(n25190), .B(n25189), .Z(n25329) );
  XNOR U25926 ( .A(n25329), .B(n25330), .Z(n25331) );
  NANDN U25927 ( .A(n25196), .B(n25195), .Z(n25200) );
  NAND U25928 ( .A(n25198), .B(n25197), .Z(n25199) );
  NAND U25929 ( .A(n25200), .B(n25199), .Z(n25404) );
  XNOR U25930 ( .A(b[19]), .B(a[164]), .Z(n25347) );
  NANDN U25931 ( .A(n25347), .B(n37934), .Z(n25203) );
  NANDN U25932 ( .A(n25201), .B(n37935), .Z(n25202) );
  NAND U25933 ( .A(n25203), .B(n25202), .Z(n25414) );
  XOR U25934 ( .A(b[27]), .B(a[156]), .Z(n25350) );
  NAND U25935 ( .A(n38423), .B(n25350), .Z(n25206) );
  NAND U25936 ( .A(n25204), .B(n38424), .Z(n25205) );
  NAND U25937 ( .A(n25206), .B(n25205), .Z(n25411) );
  XNOR U25938 ( .A(b[5]), .B(a[178]), .Z(n25353) );
  NANDN U25939 ( .A(n25353), .B(n36587), .Z(n25209) );
  NANDN U25940 ( .A(n25207), .B(n36588), .Z(n25208) );
  AND U25941 ( .A(n25209), .B(n25208), .Z(n25412) );
  XNOR U25942 ( .A(n25411), .B(n25412), .Z(n25413) );
  XNOR U25943 ( .A(n25414), .B(n25413), .Z(n25402) );
  NAND U25944 ( .A(n25210), .B(n37762), .Z(n25212) );
  XOR U25945 ( .A(b[17]), .B(a[166]), .Z(n25356) );
  NAND U25946 ( .A(n25356), .B(n37764), .Z(n25211) );
  NAND U25947 ( .A(n25212), .B(n25211), .Z(n25374) );
  XOR U25948 ( .A(b[31]), .B(n25213), .Z(n25359) );
  NANDN U25949 ( .A(n25359), .B(n38552), .Z(n25216) );
  NANDN U25950 ( .A(n25214), .B(n38553), .Z(n25215) );
  NAND U25951 ( .A(n25216), .B(n25215), .Z(n25371) );
  OR U25952 ( .A(n25217), .B(n36105), .Z(n25219) );
  XNOR U25953 ( .A(b[3]), .B(a[180]), .Z(n25362) );
  NANDN U25954 ( .A(n25362), .B(n36107), .Z(n25218) );
  AND U25955 ( .A(n25219), .B(n25218), .Z(n25372) );
  XNOR U25956 ( .A(n25371), .B(n25372), .Z(n25373) );
  XOR U25957 ( .A(n25374), .B(n25373), .Z(n25401) );
  XNOR U25958 ( .A(n25402), .B(n25401), .Z(n25403) );
  XNOR U25959 ( .A(n25404), .B(n25403), .Z(n25448) );
  NANDN U25960 ( .A(n25221), .B(n25220), .Z(n25225) );
  NAND U25961 ( .A(n25223), .B(n25222), .Z(n25224) );
  NAND U25962 ( .A(n25225), .B(n25224), .Z(n25392) );
  NANDN U25963 ( .A(n25227), .B(n25226), .Z(n25231) );
  NAND U25964 ( .A(n25229), .B(n25228), .Z(n25230) );
  NAND U25965 ( .A(n25231), .B(n25230), .Z(n25390) );
  OR U25966 ( .A(n25233), .B(n25232), .Z(n25237) );
  NANDN U25967 ( .A(n25235), .B(n25234), .Z(n25236) );
  NAND U25968 ( .A(n25237), .B(n25236), .Z(n25389) );
  XNOR U25969 ( .A(n25392), .B(n25391), .Z(n25449) );
  XNOR U25970 ( .A(n25448), .B(n25449), .Z(n25450) );
  NANDN U25971 ( .A(n25239), .B(n25238), .Z(n25243) );
  OR U25972 ( .A(n25241), .B(n25240), .Z(n25242) );
  AND U25973 ( .A(n25243), .B(n25242), .Z(n25451) );
  XOR U25974 ( .A(n25450), .B(n25451), .Z(n25337) );
  NANDN U25975 ( .A(n25249), .B(n25248), .Z(n25253) );
  NANDN U25976 ( .A(n25251), .B(n25250), .Z(n25252) );
  NAND U25977 ( .A(n25253), .B(n25252), .Z(n25457) );
  NANDN U25978 ( .A(n25259), .B(n25258), .Z(n25263) );
  NAND U25979 ( .A(n25261), .B(n25260), .Z(n25262) );
  NAND U25980 ( .A(n25263), .B(n25262), .Z(n25395) );
  NANDN U25981 ( .A(n25265), .B(n25264), .Z(n25269) );
  NAND U25982 ( .A(n25267), .B(n25266), .Z(n25268) );
  AND U25983 ( .A(n25269), .B(n25268), .Z(n25396) );
  XNOR U25984 ( .A(n25395), .B(n25396), .Z(n25397) );
  XNOR U25985 ( .A(b[9]), .B(a[174]), .Z(n25417) );
  NANDN U25986 ( .A(n25417), .B(n36925), .Z(n25272) );
  NANDN U25987 ( .A(n25270), .B(n36926), .Z(n25271) );
  NAND U25988 ( .A(n25272), .B(n25271), .Z(n25379) );
  XNOR U25989 ( .A(b[15]), .B(a[168]), .Z(n25420) );
  OR U25990 ( .A(n25420), .B(n37665), .Z(n25275) );
  NANDN U25991 ( .A(n25273), .B(n37604), .Z(n25274) );
  AND U25992 ( .A(n25275), .B(n25274), .Z(n25377) );
  XNOR U25993 ( .A(b[21]), .B(a[162]), .Z(n25423) );
  NANDN U25994 ( .A(n25423), .B(n38101), .Z(n25278) );
  NANDN U25995 ( .A(n25276), .B(n38102), .Z(n25277) );
  AND U25996 ( .A(n25278), .B(n25277), .Z(n25378) );
  XOR U25997 ( .A(n25379), .B(n25380), .Z(n25368) );
  XNOR U25998 ( .A(b[11]), .B(a[172]), .Z(n25426) );
  OR U25999 ( .A(n25426), .B(n37311), .Z(n25281) );
  NANDN U26000 ( .A(n25279), .B(n37218), .Z(n25280) );
  NAND U26001 ( .A(n25281), .B(n25280), .Z(n25366) );
  XOR U26002 ( .A(n1053), .B(a[170]), .Z(n25429) );
  NANDN U26003 ( .A(n25429), .B(n37424), .Z(n25284) );
  NANDN U26004 ( .A(n25282), .B(n37425), .Z(n25283) );
  AND U26005 ( .A(n25284), .B(n25283), .Z(n25365) );
  XNOR U26006 ( .A(n25366), .B(n25365), .Z(n25367) );
  XOR U26007 ( .A(n25368), .B(n25367), .Z(n25385) );
  NANDN U26008 ( .A(n1049), .B(a[182]), .Z(n25285) );
  XNOR U26009 ( .A(b[1]), .B(n25285), .Z(n25287) );
  NANDN U26010 ( .A(b[0]), .B(a[181]), .Z(n25286) );
  AND U26011 ( .A(n25287), .B(n25286), .Z(n25343) );
  NAND U26012 ( .A(n38490), .B(n25288), .Z(n25290) );
  XOR U26013 ( .A(b[29]), .B(n25862), .Z(n25436) );
  OR U26014 ( .A(n25436), .B(n1048), .Z(n25289) );
  NAND U26015 ( .A(n25290), .B(n25289), .Z(n25341) );
  NANDN U26016 ( .A(n1059), .B(a[150]), .Z(n25342) );
  XNOR U26017 ( .A(n25341), .B(n25342), .Z(n25344) );
  XOR U26018 ( .A(n25343), .B(n25344), .Z(n25383) );
  NANDN U26019 ( .A(n25291), .B(n38205), .Z(n25293) );
  XNOR U26020 ( .A(b[23]), .B(a[160]), .Z(n25439) );
  OR U26021 ( .A(n25439), .B(n38268), .Z(n25292) );
  NAND U26022 ( .A(n25293), .B(n25292), .Z(n25408) );
  XOR U26023 ( .A(b[7]), .B(a[176]), .Z(n25442) );
  NAND U26024 ( .A(n25442), .B(n36701), .Z(n25296) );
  NAND U26025 ( .A(n25294), .B(n36702), .Z(n25295) );
  NAND U26026 ( .A(n25296), .B(n25295), .Z(n25405) );
  XOR U26027 ( .A(b[25]), .B(a[158]), .Z(n25445) );
  NAND U26028 ( .A(n25445), .B(n38325), .Z(n25299) );
  NAND U26029 ( .A(n25297), .B(n38326), .Z(n25298) );
  AND U26030 ( .A(n25299), .B(n25298), .Z(n25406) );
  XNOR U26031 ( .A(n25405), .B(n25406), .Z(n25407) );
  XNOR U26032 ( .A(n25408), .B(n25407), .Z(n25384) );
  XOR U26033 ( .A(n25383), .B(n25384), .Z(n25386) );
  XNOR U26034 ( .A(n25385), .B(n25386), .Z(n25398) );
  XOR U26035 ( .A(n25397), .B(n25398), .Z(n25455) );
  XNOR U26036 ( .A(n25454), .B(n25455), .Z(n25456) );
  XNOR U26037 ( .A(n25457), .B(n25456), .Z(n25335) );
  XNOR U26038 ( .A(n25336), .B(n25335), .Z(n25338) );
  XNOR U26039 ( .A(n25337), .B(n25338), .Z(n25332) );
  XOR U26040 ( .A(n25331), .B(n25332), .Z(n25326) );
  NANDN U26041 ( .A(n25301), .B(n25300), .Z(n25305) );
  NAND U26042 ( .A(n25303), .B(n25302), .Z(n25304) );
  NAND U26043 ( .A(n25305), .B(n25304), .Z(n25323) );
  NANDN U26044 ( .A(n25307), .B(n25306), .Z(n25311) );
  OR U26045 ( .A(n25309), .B(n25308), .Z(n25310) );
  NAND U26046 ( .A(n25311), .B(n25310), .Z(n25324) );
  XNOR U26047 ( .A(n25323), .B(n25324), .Z(n25325) );
  XNOR U26048 ( .A(n25326), .B(n25325), .Z(n25318) );
  XNOR U26049 ( .A(n25317), .B(n25318), .Z(n25319) );
  XNOR U26050 ( .A(n25320), .B(n25319), .Z(n25460) );
  XNOR U26051 ( .A(n25460), .B(sreg[406]), .Z(n25462) );
  NAND U26052 ( .A(n25312), .B(sreg[405]), .Z(n25316) );
  OR U26053 ( .A(n25314), .B(n25313), .Z(n25315) );
  AND U26054 ( .A(n25316), .B(n25315), .Z(n25461) );
  XOR U26055 ( .A(n25462), .B(n25461), .Z(c[406]) );
  NANDN U26056 ( .A(n25318), .B(n25317), .Z(n25322) );
  NAND U26057 ( .A(n25320), .B(n25319), .Z(n25321) );
  NAND U26058 ( .A(n25322), .B(n25321), .Z(n25468) );
  NANDN U26059 ( .A(n25324), .B(n25323), .Z(n25328) );
  NAND U26060 ( .A(n25326), .B(n25325), .Z(n25327) );
  NAND U26061 ( .A(n25328), .B(n25327), .Z(n25466) );
  NANDN U26062 ( .A(n25330), .B(n25329), .Z(n25334) );
  NANDN U26063 ( .A(n25332), .B(n25331), .Z(n25333) );
  NAND U26064 ( .A(n25334), .B(n25333), .Z(n25472) );
  OR U26065 ( .A(n25336), .B(n25335), .Z(n25340) );
  OR U26066 ( .A(n25338), .B(n25337), .Z(n25339) );
  AND U26067 ( .A(n25340), .B(n25339), .Z(n25471) );
  XNOR U26068 ( .A(n25472), .B(n25471), .Z(n25473) );
  NANDN U26069 ( .A(n25342), .B(n25341), .Z(n25346) );
  NAND U26070 ( .A(n25344), .B(n25343), .Z(n25345) );
  NAND U26071 ( .A(n25346), .B(n25345), .Z(n25552) );
  XNOR U26072 ( .A(b[19]), .B(a[165]), .Z(n25519) );
  NANDN U26073 ( .A(n25519), .B(n37934), .Z(n25349) );
  NANDN U26074 ( .A(n25347), .B(n37935), .Z(n25348) );
  NAND U26075 ( .A(n25349), .B(n25348), .Z(n25564) );
  XOR U26076 ( .A(b[27]), .B(a[157]), .Z(n25522) );
  NAND U26077 ( .A(n38423), .B(n25522), .Z(n25352) );
  NAND U26078 ( .A(n25350), .B(n38424), .Z(n25351) );
  NAND U26079 ( .A(n25352), .B(n25351), .Z(n25561) );
  XNOR U26080 ( .A(b[5]), .B(a[179]), .Z(n25525) );
  NANDN U26081 ( .A(n25525), .B(n36587), .Z(n25355) );
  NANDN U26082 ( .A(n25353), .B(n36588), .Z(n25354) );
  AND U26083 ( .A(n25355), .B(n25354), .Z(n25562) );
  XNOR U26084 ( .A(n25561), .B(n25562), .Z(n25563) );
  XNOR U26085 ( .A(n25564), .B(n25563), .Z(n25549) );
  NAND U26086 ( .A(n25356), .B(n37762), .Z(n25358) );
  XOR U26087 ( .A(b[17]), .B(a[167]), .Z(n25528) );
  NAND U26088 ( .A(n25528), .B(n37764), .Z(n25357) );
  NAND U26089 ( .A(n25358), .B(n25357), .Z(n25503) );
  XNOR U26090 ( .A(b[31]), .B(a[153]), .Z(n25531) );
  NANDN U26091 ( .A(n25531), .B(n38552), .Z(n25361) );
  NANDN U26092 ( .A(n25359), .B(n38553), .Z(n25360) );
  AND U26093 ( .A(n25361), .B(n25360), .Z(n25501) );
  OR U26094 ( .A(n25362), .B(n36105), .Z(n25364) );
  XNOR U26095 ( .A(b[3]), .B(a[181]), .Z(n25534) );
  NANDN U26096 ( .A(n25534), .B(n36107), .Z(n25363) );
  AND U26097 ( .A(n25364), .B(n25363), .Z(n25502) );
  XOR U26098 ( .A(n25503), .B(n25504), .Z(n25550) );
  XOR U26099 ( .A(n25549), .B(n25550), .Z(n25551) );
  XNOR U26100 ( .A(n25552), .B(n25551), .Z(n25597) );
  NANDN U26101 ( .A(n25366), .B(n25365), .Z(n25370) );
  NAND U26102 ( .A(n25368), .B(n25367), .Z(n25369) );
  NAND U26103 ( .A(n25370), .B(n25369), .Z(n25540) );
  NANDN U26104 ( .A(n25372), .B(n25371), .Z(n25376) );
  NAND U26105 ( .A(n25374), .B(n25373), .Z(n25375) );
  NAND U26106 ( .A(n25376), .B(n25375), .Z(n25538) );
  OR U26107 ( .A(n25378), .B(n25377), .Z(n25382) );
  NANDN U26108 ( .A(n25380), .B(n25379), .Z(n25381) );
  NAND U26109 ( .A(n25382), .B(n25381), .Z(n25537) );
  XNOR U26110 ( .A(n25540), .B(n25539), .Z(n25598) );
  XOR U26111 ( .A(n25597), .B(n25598), .Z(n25600) );
  NANDN U26112 ( .A(n25384), .B(n25383), .Z(n25388) );
  OR U26113 ( .A(n25386), .B(n25385), .Z(n25387) );
  NAND U26114 ( .A(n25388), .B(n25387), .Z(n25599) );
  XOR U26115 ( .A(n25600), .B(n25599), .Z(n25485) );
  OR U26116 ( .A(n25390), .B(n25389), .Z(n25394) );
  NAND U26117 ( .A(n25392), .B(n25391), .Z(n25393) );
  NAND U26118 ( .A(n25394), .B(n25393), .Z(n25484) );
  NANDN U26119 ( .A(n25396), .B(n25395), .Z(n25400) );
  NANDN U26120 ( .A(n25398), .B(n25397), .Z(n25399) );
  NAND U26121 ( .A(n25400), .B(n25399), .Z(n25605) );
  NANDN U26122 ( .A(n25406), .B(n25405), .Z(n25410) );
  NAND U26123 ( .A(n25408), .B(n25407), .Z(n25409) );
  NAND U26124 ( .A(n25410), .B(n25409), .Z(n25543) );
  NANDN U26125 ( .A(n25412), .B(n25411), .Z(n25416) );
  NAND U26126 ( .A(n25414), .B(n25413), .Z(n25415) );
  AND U26127 ( .A(n25416), .B(n25415), .Z(n25544) );
  XNOR U26128 ( .A(n25543), .B(n25544), .Z(n25545) );
  XNOR U26129 ( .A(n1052), .B(a[175]), .Z(n25573) );
  NAND U26130 ( .A(n36925), .B(n25573), .Z(n25419) );
  NANDN U26131 ( .A(n25417), .B(n36926), .Z(n25418) );
  NAND U26132 ( .A(n25419), .B(n25418), .Z(n25509) );
  XNOR U26133 ( .A(b[15]), .B(a[169]), .Z(n25570) );
  OR U26134 ( .A(n25570), .B(n37665), .Z(n25422) );
  NANDN U26135 ( .A(n25420), .B(n37604), .Z(n25421) );
  AND U26136 ( .A(n25422), .B(n25421), .Z(n25507) );
  XOR U26137 ( .A(n1056), .B(n27178), .Z(n25567) );
  NAND U26138 ( .A(n25567), .B(n38101), .Z(n25425) );
  NANDN U26139 ( .A(n25423), .B(n38102), .Z(n25424) );
  AND U26140 ( .A(n25425), .B(n25424), .Z(n25508) );
  XOR U26141 ( .A(n25509), .B(n25510), .Z(n25498) );
  XNOR U26142 ( .A(b[11]), .B(a[173]), .Z(n25576) );
  OR U26143 ( .A(n25576), .B(n37311), .Z(n25428) );
  NANDN U26144 ( .A(n25426), .B(n37218), .Z(n25427) );
  NAND U26145 ( .A(n25428), .B(n25427), .Z(n25496) );
  XOR U26146 ( .A(n1053), .B(a[171]), .Z(n25579) );
  NANDN U26147 ( .A(n25579), .B(n37424), .Z(n25431) );
  NANDN U26148 ( .A(n25429), .B(n37425), .Z(n25430) );
  NAND U26149 ( .A(n25431), .B(n25430), .Z(n25495) );
  XOR U26150 ( .A(n25498), .B(n25497), .Z(n25492) );
  NANDN U26151 ( .A(n1049), .B(a[183]), .Z(n25432) );
  XNOR U26152 ( .A(b[1]), .B(n25432), .Z(n25434) );
  NANDN U26153 ( .A(b[0]), .B(a[182]), .Z(n25433) );
  AND U26154 ( .A(n25434), .B(n25433), .Z(n25516) );
  ANDN U26155 ( .B(b[31]), .A(n25435), .Z(n25513) );
  NANDN U26156 ( .A(n25436), .B(n38490), .Z(n25438) );
  XNOR U26157 ( .A(n1058), .B(a[155]), .Z(n25585) );
  NANDN U26158 ( .A(n1048), .B(n25585), .Z(n25437) );
  NAND U26159 ( .A(n25438), .B(n25437), .Z(n25514) );
  XOR U26160 ( .A(n25513), .B(n25514), .Z(n25515) );
  XNOR U26161 ( .A(n25516), .B(n25515), .Z(n25489) );
  NANDN U26162 ( .A(n25439), .B(n38205), .Z(n25441) );
  XOR U26163 ( .A(b[23]), .B(n26869), .Z(n25588) );
  OR U26164 ( .A(n25588), .B(n38268), .Z(n25440) );
  NAND U26165 ( .A(n25441), .B(n25440), .Z(n25558) );
  XOR U26166 ( .A(b[7]), .B(a[177]), .Z(n25591) );
  NAND U26167 ( .A(n25591), .B(n36701), .Z(n25444) );
  NAND U26168 ( .A(n25442), .B(n36702), .Z(n25443) );
  NAND U26169 ( .A(n25444), .B(n25443), .Z(n25555) );
  XOR U26170 ( .A(b[25]), .B(a[159]), .Z(n25594) );
  NAND U26171 ( .A(n25594), .B(n38325), .Z(n25447) );
  NAND U26172 ( .A(n25445), .B(n38326), .Z(n25446) );
  AND U26173 ( .A(n25447), .B(n25446), .Z(n25556) );
  XNOR U26174 ( .A(n25555), .B(n25556), .Z(n25557) );
  XNOR U26175 ( .A(n25558), .B(n25557), .Z(n25490) );
  XOR U26176 ( .A(n25492), .B(n25491), .Z(n25546) );
  XNOR U26177 ( .A(n25545), .B(n25546), .Z(n25603) );
  XNOR U26178 ( .A(n25604), .B(n25603), .Z(n25606) );
  XNOR U26179 ( .A(n25605), .B(n25606), .Z(n25483) );
  XOR U26180 ( .A(n25484), .B(n25483), .Z(n25486) );
  NANDN U26181 ( .A(n25449), .B(n25448), .Z(n25453) );
  NAND U26182 ( .A(n25451), .B(n25450), .Z(n25452) );
  NAND U26183 ( .A(n25453), .B(n25452), .Z(n25477) );
  NANDN U26184 ( .A(n25455), .B(n25454), .Z(n25459) );
  NAND U26185 ( .A(n25457), .B(n25456), .Z(n25458) );
  NAND U26186 ( .A(n25459), .B(n25458), .Z(n25478) );
  XNOR U26187 ( .A(n25477), .B(n25478), .Z(n25479) );
  XOR U26188 ( .A(n25480), .B(n25479), .Z(n25474) );
  XOR U26189 ( .A(n25473), .B(n25474), .Z(n25465) );
  XOR U26190 ( .A(n25466), .B(n25465), .Z(n25467) );
  XNOR U26191 ( .A(n25468), .B(n25467), .Z(n25609) );
  XNOR U26192 ( .A(n25609), .B(sreg[407]), .Z(n25611) );
  NAND U26193 ( .A(n25460), .B(sreg[406]), .Z(n25464) );
  OR U26194 ( .A(n25462), .B(n25461), .Z(n25463) );
  AND U26195 ( .A(n25464), .B(n25463), .Z(n25610) );
  XOR U26196 ( .A(n25611), .B(n25610), .Z(c[407]) );
  NAND U26197 ( .A(n25466), .B(n25465), .Z(n25470) );
  NAND U26198 ( .A(n25468), .B(n25467), .Z(n25469) );
  NAND U26199 ( .A(n25470), .B(n25469), .Z(n25617) );
  NANDN U26200 ( .A(n25472), .B(n25471), .Z(n25476) );
  NAND U26201 ( .A(n25474), .B(n25473), .Z(n25475) );
  NAND U26202 ( .A(n25476), .B(n25475), .Z(n25615) );
  NANDN U26203 ( .A(n25478), .B(n25477), .Z(n25482) );
  NAND U26204 ( .A(n25480), .B(n25479), .Z(n25481) );
  NAND U26205 ( .A(n25482), .B(n25481), .Z(n25620) );
  NANDN U26206 ( .A(n25484), .B(n25483), .Z(n25488) );
  OR U26207 ( .A(n25486), .B(n25485), .Z(n25487) );
  NAND U26208 ( .A(n25488), .B(n25487), .Z(n25621) );
  XNOR U26209 ( .A(n25620), .B(n25621), .Z(n25622) );
  OR U26210 ( .A(n25490), .B(n25489), .Z(n25494) );
  NANDN U26211 ( .A(n25492), .B(n25491), .Z(n25493) );
  NAND U26212 ( .A(n25494), .B(n25493), .Z(n25747) );
  OR U26213 ( .A(n25496), .B(n25495), .Z(n25500) );
  NAND U26214 ( .A(n25498), .B(n25497), .Z(n25499) );
  NAND U26215 ( .A(n25500), .B(n25499), .Z(n25686) );
  OR U26216 ( .A(n25502), .B(n25501), .Z(n25506) );
  NANDN U26217 ( .A(n25504), .B(n25503), .Z(n25505) );
  NAND U26218 ( .A(n25506), .B(n25505), .Z(n25685) );
  OR U26219 ( .A(n25508), .B(n25507), .Z(n25512) );
  NANDN U26220 ( .A(n25510), .B(n25509), .Z(n25511) );
  NAND U26221 ( .A(n25512), .B(n25511), .Z(n25684) );
  XOR U26222 ( .A(n25686), .B(n25687), .Z(n25745) );
  OR U26223 ( .A(n25514), .B(n25513), .Z(n25518) );
  NANDN U26224 ( .A(n25516), .B(n25515), .Z(n25517) );
  NAND U26225 ( .A(n25518), .B(n25517), .Z(n25698) );
  XNOR U26226 ( .A(b[19]), .B(a[166]), .Z(n25644) );
  NANDN U26227 ( .A(n25644), .B(n37934), .Z(n25521) );
  NANDN U26228 ( .A(n25519), .B(n37935), .Z(n25520) );
  NAND U26229 ( .A(n25521), .B(n25520), .Z(n25711) );
  XOR U26230 ( .A(b[27]), .B(a[158]), .Z(n25647) );
  NAND U26231 ( .A(n38423), .B(n25647), .Z(n25524) );
  NAND U26232 ( .A(n25522), .B(n38424), .Z(n25523) );
  NAND U26233 ( .A(n25524), .B(n25523), .Z(n25708) );
  XNOR U26234 ( .A(b[5]), .B(a[180]), .Z(n25650) );
  NANDN U26235 ( .A(n25650), .B(n36587), .Z(n25527) );
  NANDN U26236 ( .A(n25525), .B(n36588), .Z(n25526) );
  AND U26237 ( .A(n25527), .B(n25526), .Z(n25709) );
  XNOR U26238 ( .A(n25708), .B(n25709), .Z(n25710) );
  XNOR U26239 ( .A(n25711), .B(n25710), .Z(n25697) );
  NAND U26240 ( .A(n25528), .B(n37762), .Z(n25530) );
  XOR U26241 ( .A(b[17]), .B(a[168]), .Z(n25653) );
  NAND U26242 ( .A(n25653), .B(n37764), .Z(n25529) );
  NAND U26243 ( .A(n25530), .B(n25529), .Z(n25671) );
  XOR U26244 ( .A(b[31]), .B(n25862), .Z(n25656) );
  NANDN U26245 ( .A(n25656), .B(n38552), .Z(n25533) );
  NANDN U26246 ( .A(n25531), .B(n38553), .Z(n25532) );
  NAND U26247 ( .A(n25533), .B(n25532), .Z(n25668) );
  OR U26248 ( .A(n25534), .B(n36105), .Z(n25536) );
  XNOR U26249 ( .A(b[3]), .B(a[182]), .Z(n25659) );
  NANDN U26250 ( .A(n25659), .B(n36107), .Z(n25535) );
  AND U26251 ( .A(n25536), .B(n25535), .Z(n25669) );
  XNOR U26252 ( .A(n25668), .B(n25669), .Z(n25670) );
  XOR U26253 ( .A(n25671), .B(n25670), .Z(n25696) );
  XOR U26254 ( .A(n25697), .B(n25696), .Z(n25699) );
  XOR U26255 ( .A(n25698), .B(n25699), .Z(n25744) );
  XOR U26256 ( .A(n25745), .B(n25744), .Z(n25746) );
  XNOR U26257 ( .A(n25747), .B(n25746), .Z(n25635) );
  OR U26258 ( .A(n25538), .B(n25537), .Z(n25542) );
  NAND U26259 ( .A(n25540), .B(n25539), .Z(n25541) );
  NAND U26260 ( .A(n25542), .B(n25541), .Z(n25633) );
  NANDN U26261 ( .A(n25544), .B(n25543), .Z(n25548) );
  NANDN U26262 ( .A(n25546), .B(n25545), .Z(n25547) );
  NAND U26263 ( .A(n25548), .B(n25547), .Z(n25752) );
  OR U26264 ( .A(n25550), .B(n25549), .Z(n25554) );
  NAND U26265 ( .A(n25552), .B(n25551), .Z(n25553) );
  NAND U26266 ( .A(n25554), .B(n25553), .Z(n25751) );
  NANDN U26267 ( .A(n25556), .B(n25555), .Z(n25560) );
  NAND U26268 ( .A(n25558), .B(n25557), .Z(n25559) );
  NAND U26269 ( .A(n25560), .B(n25559), .Z(n25690) );
  NANDN U26270 ( .A(n25562), .B(n25561), .Z(n25566) );
  NAND U26271 ( .A(n25564), .B(n25563), .Z(n25565) );
  AND U26272 ( .A(n25566), .B(n25565), .Z(n25691) );
  XNOR U26273 ( .A(n25690), .B(n25691), .Z(n25692) );
  XNOR U26274 ( .A(b[21]), .B(a[164]), .Z(n25720) );
  NANDN U26275 ( .A(n25720), .B(n38101), .Z(n25569) );
  NAND U26276 ( .A(n38102), .B(n25567), .Z(n25568) );
  NAND U26277 ( .A(n25569), .B(n25568), .Z(n25680) );
  XNOR U26278 ( .A(b[15]), .B(a[170]), .Z(n25717) );
  OR U26279 ( .A(n25717), .B(n37665), .Z(n25572) );
  NANDN U26280 ( .A(n25570), .B(n37604), .Z(n25571) );
  AND U26281 ( .A(n25572), .B(n25571), .Z(n25681) );
  XNOR U26282 ( .A(n25680), .B(n25681), .Z(n25683) );
  XNOR U26283 ( .A(b[9]), .B(a[176]), .Z(n25714) );
  NANDN U26284 ( .A(n25714), .B(n36925), .Z(n25575) );
  NAND U26285 ( .A(n36926), .B(n25573), .Z(n25574) );
  NAND U26286 ( .A(n25575), .B(n25574), .Z(n25682) );
  XNOR U26287 ( .A(n25683), .B(n25682), .Z(n25676) );
  XNOR U26288 ( .A(b[11]), .B(a[174]), .Z(n25723) );
  OR U26289 ( .A(n25723), .B(n37311), .Z(n25578) );
  NANDN U26290 ( .A(n25576), .B(n37218), .Z(n25577) );
  NAND U26291 ( .A(n25578), .B(n25577), .Z(n25675) );
  XOR U26292 ( .A(n1053), .B(a[172]), .Z(n25726) );
  NANDN U26293 ( .A(n25726), .B(n37424), .Z(n25581) );
  NANDN U26294 ( .A(n25579), .B(n37425), .Z(n25580) );
  NAND U26295 ( .A(n25581), .B(n25580), .Z(n25674) );
  XNOR U26296 ( .A(n25675), .B(n25674), .Z(n25677) );
  XNOR U26297 ( .A(n25676), .B(n25677), .Z(n25665) );
  NANDN U26298 ( .A(n1049), .B(a[184]), .Z(n25582) );
  XNOR U26299 ( .A(b[1]), .B(n25582), .Z(n25584) );
  NANDN U26300 ( .A(b[0]), .B(a[183]), .Z(n25583) );
  AND U26301 ( .A(n25584), .B(n25583), .Z(n25640) );
  NAND U26302 ( .A(n25585), .B(n38490), .Z(n25587) );
  XNOR U26303 ( .A(n1058), .B(a[156]), .Z(n25732) );
  NANDN U26304 ( .A(n1048), .B(n25732), .Z(n25586) );
  NAND U26305 ( .A(n25587), .B(n25586), .Z(n25638) );
  NANDN U26306 ( .A(n1059), .B(a[152]), .Z(n25639) );
  XNOR U26307 ( .A(n25638), .B(n25639), .Z(n25641) );
  XNOR U26308 ( .A(n25640), .B(n25641), .Z(n25663) );
  NANDN U26309 ( .A(n25588), .B(n38205), .Z(n25590) );
  XNOR U26310 ( .A(b[23]), .B(a[162]), .Z(n25735) );
  OR U26311 ( .A(n25735), .B(n38268), .Z(n25589) );
  NAND U26312 ( .A(n25590), .B(n25589), .Z(n25705) );
  XOR U26313 ( .A(b[7]), .B(a[178]), .Z(n25738) );
  NAND U26314 ( .A(n25738), .B(n36701), .Z(n25593) );
  NAND U26315 ( .A(n25591), .B(n36702), .Z(n25592) );
  NAND U26316 ( .A(n25593), .B(n25592), .Z(n25702) );
  XOR U26317 ( .A(b[25]), .B(a[160]), .Z(n25741) );
  NAND U26318 ( .A(n25741), .B(n38325), .Z(n25596) );
  NAND U26319 ( .A(n25594), .B(n38326), .Z(n25595) );
  AND U26320 ( .A(n25596), .B(n25595), .Z(n25703) );
  XNOR U26321 ( .A(n25702), .B(n25703), .Z(n25704) );
  XOR U26322 ( .A(n25705), .B(n25704), .Z(n25662) );
  XOR U26323 ( .A(n25665), .B(n25664), .Z(n25693) );
  XNOR U26324 ( .A(n25692), .B(n25693), .Z(n25750) );
  XNOR U26325 ( .A(n25751), .B(n25750), .Z(n25753) );
  XNOR U26326 ( .A(n25752), .B(n25753), .Z(n25632) );
  XNOR U26327 ( .A(n25633), .B(n25632), .Z(n25634) );
  XOR U26328 ( .A(n25635), .B(n25634), .Z(n25629) );
  NANDN U26329 ( .A(n25598), .B(n25597), .Z(n25602) );
  OR U26330 ( .A(n25600), .B(n25599), .Z(n25601) );
  NAND U26331 ( .A(n25602), .B(n25601), .Z(n25626) );
  NAND U26332 ( .A(n25604), .B(n25603), .Z(n25608) );
  NANDN U26333 ( .A(n25606), .B(n25605), .Z(n25607) );
  NAND U26334 ( .A(n25608), .B(n25607), .Z(n25627) );
  XNOR U26335 ( .A(n25626), .B(n25627), .Z(n25628) );
  XOR U26336 ( .A(n25629), .B(n25628), .Z(n25623) );
  XOR U26337 ( .A(n25622), .B(n25623), .Z(n25614) );
  XOR U26338 ( .A(n25615), .B(n25614), .Z(n25616) );
  XNOR U26339 ( .A(n25617), .B(n25616), .Z(n25756) );
  XNOR U26340 ( .A(n25756), .B(sreg[408]), .Z(n25758) );
  NAND U26341 ( .A(n25609), .B(sreg[407]), .Z(n25613) );
  OR U26342 ( .A(n25611), .B(n25610), .Z(n25612) );
  AND U26343 ( .A(n25613), .B(n25612), .Z(n25757) );
  XOR U26344 ( .A(n25758), .B(n25757), .Z(c[408]) );
  NAND U26345 ( .A(n25615), .B(n25614), .Z(n25619) );
  NAND U26346 ( .A(n25617), .B(n25616), .Z(n25618) );
  NAND U26347 ( .A(n25619), .B(n25618), .Z(n25764) );
  NANDN U26348 ( .A(n25621), .B(n25620), .Z(n25625) );
  NAND U26349 ( .A(n25623), .B(n25622), .Z(n25624) );
  NAND U26350 ( .A(n25625), .B(n25624), .Z(n25762) );
  NANDN U26351 ( .A(n25627), .B(n25626), .Z(n25631) );
  NAND U26352 ( .A(n25629), .B(n25628), .Z(n25630) );
  NAND U26353 ( .A(n25631), .B(n25630), .Z(n25767) );
  NANDN U26354 ( .A(n25633), .B(n25632), .Z(n25637) );
  NANDN U26355 ( .A(n25635), .B(n25634), .Z(n25636) );
  NAND U26356 ( .A(n25637), .B(n25636), .Z(n25768) );
  XNOR U26357 ( .A(n25767), .B(n25768), .Z(n25769) );
  NANDN U26358 ( .A(n25639), .B(n25638), .Z(n25643) );
  NAND U26359 ( .A(n25641), .B(n25640), .Z(n25642) );
  NAND U26360 ( .A(n25643), .B(n25642), .Z(n25834) );
  XNOR U26361 ( .A(b[19]), .B(a[167]), .Z(n25779) );
  NANDN U26362 ( .A(n25779), .B(n37934), .Z(n25646) );
  NANDN U26363 ( .A(n25644), .B(n37935), .Z(n25645) );
  NAND U26364 ( .A(n25646), .B(n25645), .Z(n25844) );
  XOR U26365 ( .A(b[27]), .B(a[159]), .Z(n25782) );
  NAND U26366 ( .A(n38423), .B(n25782), .Z(n25649) );
  NAND U26367 ( .A(n25647), .B(n38424), .Z(n25648) );
  NAND U26368 ( .A(n25649), .B(n25648), .Z(n25841) );
  XNOR U26369 ( .A(b[5]), .B(a[181]), .Z(n25785) );
  NANDN U26370 ( .A(n25785), .B(n36587), .Z(n25652) );
  NANDN U26371 ( .A(n25650), .B(n36588), .Z(n25651) );
  AND U26372 ( .A(n25652), .B(n25651), .Z(n25842) );
  XNOR U26373 ( .A(n25841), .B(n25842), .Z(n25843) );
  XNOR U26374 ( .A(n25844), .B(n25843), .Z(n25832) );
  NAND U26375 ( .A(n25653), .B(n37762), .Z(n25655) );
  XOR U26376 ( .A(b[17]), .B(a[169]), .Z(n25788) );
  NAND U26377 ( .A(n25788), .B(n37764), .Z(n25654) );
  NAND U26378 ( .A(n25655), .B(n25654), .Z(n25806) );
  XNOR U26379 ( .A(b[31]), .B(a[155]), .Z(n25791) );
  NANDN U26380 ( .A(n25791), .B(n38552), .Z(n25658) );
  NANDN U26381 ( .A(n25656), .B(n38553), .Z(n25657) );
  NAND U26382 ( .A(n25658), .B(n25657), .Z(n25803) );
  OR U26383 ( .A(n25659), .B(n36105), .Z(n25661) );
  XNOR U26384 ( .A(b[3]), .B(a[183]), .Z(n25794) );
  NANDN U26385 ( .A(n25794), .B(n36107), .Z(n25660) );
  AND U26386 ( .A(n25661), .B(n25660), .Z(n25804) );
  XNOR U26387 ( .A(n25803), .B(n25804), .Z(n25805) );
  XOR U26388 ( .A(n25806), .B(n25805), .Z(n25831) );
  XNOR U26389 ( .A(n25832), .B(n25831), .Z(n25833) );
  XNOR U26390 ( .A(n25834), .B(n25833), .Z(n25884) );
  NANDN U26391 ( .A(n25663), .B(n25662), .Z(n25667) );
  NANDN U26392 ( .A(n25665), .B(n25664), .Z(n25666) );
  NAND U26393 ( .A(n25667), .B(n25666), .Z(n25885) );
  XNOR U26394 ( .A(n25884), .B(n25885), .Z(n25886) );
  NANDN U26395 ( .A(n25669), .B(n25668), .Z(n25673) );
  NAND U26396 ( .A(n25671), .B(n25670), .Z(n25672) );
  NAND U26397 ( .A(n25673), .B(n25672), .Z(n25824) );
  OR U26398 ( .A(n25675), .B(n25674), .Z(n25679) );
  NANDN U26399 ( .A(n25677), .B(n25676), .Z(n25678) );
  NAND U26400 ( .A(n25679), .B(n25678), .Z(n25822) );
  XNOR U26401 ( .A(n25822), .B(n25821), .Z(n25823) );
  XOR U26402 ( .A(n25824), .B(n25823), .Z(n25887) );
  XOR U26403 ( .A(n25886), .B(n25887), .Z(n25897) );
  OR U26404 ( .A(n25685), .B(n25684), .Z(n25689) );
  NANDN U26405 ( .A(n25687), .B(n25686), .Z(n25688) );
  NAND U26406 ( .A(n25689), .B(n25688), .Z(n25895) );
  NANDN U26407 ( .A(n25691), .B(n25690), .Z(n25695) );
  NANDN U26408 ( .A(n25693), .B(n25692), .Z(n25694) );
  NAND U26409 ( .A(n25695), .B(n25694), .Z(n25880) );
  NANDN U26410 ( .A(n25697), .B(n25696), .Z(n25701) );
  OR U26411 ( .A(n25699), .B(n25698), .Z(n25700) );
  NAND U26412 ( .A(n25701), .B(n25700), .Z(n25879) );
  NANDN U26413 ( .A(n25703), .B(n25702), .Z(n25707) );
  NAND U26414 ( .A(n25705), .B(n25704), .Z(n25706) );
  NAND U26415 ( .A(n25707), .B(n25706), .Z(n25825) );
  NANDN U26416 ( .A(n25709), .B(n25708), .Z(n25713) );
  NAND U26417 ( .A(n25711), .B(n25710), .Z(n25712) );
  AND U26418 ( .A(n25713), .B(n25712), .Z(n25826) );
  XNOR U26419 ( .A(n25825), .B(n25826), .Z(n25827) );
  XNOR U26420 ( .A(b[9]), .B(a[177]), .Z(n25847) );
  NANDN U26421 ( .A(n25847), .B(n36925), .Z(n25716) );
  NANDN U26422 ( .A(n25714), .B(n36926), .Z(n25715) );
  NAND U26423 ( .A(n25716), .B(n25715), .Z(n25811) );
  XNOR U26424 ( .A(b[15]), .B(a[171]), .Z(n25850) );
  OR U26425 ( .A(n25850), .B(n37665), .Z(n25719) );
  NANDN U26426 ( .A(n25717), .B(n37604), .Z(n25718) );
  AND U26427 ( .A(n25719), .B(n25718), .Z(n25809) );
  XNOR U26428 ( .A(b[21]), .B(a[165]), .Z(n25853) );
  NANDN U26429 ( .A(n25853), .B(n38101), .Z(n25722) );
  NANDN U26430 ( .A(n25720), .B(n38102), .Z(n25721) );
  AND U26431 ( .A(n25722), .B(n25721), .Z(n25810) );
  XOR U26432 ( .A(n25811), .B(n25812), .Z(n25800) );
  XNOR U26433 ( .A(b[11]), .B(a[175]), .Z(n25856) );
  OR U26434 ( .A(n25856), .B(n37311), .Z(n25725) );
  NANDN U26435 ( .A(n25723), .B(n37218), .Z(n25724) );
  NAND U26436 ( .A(n25725), .B(n25724), .Z(n25798) );
  XOR U26437 ( .A(n1053), .B(a[173]), .Z(n25859) );
  NANDN U26438 ( .A(n25859), .B(n37424), .Z(n25728) );
  NANDN U26439 ( .A(n25726), .B(n37425), .Z(n25727) );
  AND U26440 ( .A(n25728), .B(n25727), .Z(n25797) );
  XNOR U26441 ( .A(n25798), .B(n25797), .Z(n25799) );
  XOR U26442 ( .A(n25800), .B(n25799), .Z(n25817) );
  NANDN U26443 ( .A(n1049), .B(a[185]), .Z(n25729) );
  XNOR U26444 ( .A(b[1]), .B(n25729), .Z(n25731) );
  NANDN U26445 ( .A(b[0]), .B(a[184]), .Z(n25730) );
  AND U26446 ( .A(n25731), .B(n25730), .Z(n25775) );
  NAND U26447 ( .A(n38490), .B(n25732), .Z(n25734) );
  XNOR U26448 ( .A(b[29]), .B(a[157]), .Z(n25863) );
  OR U26449 ( .A(n25863), .B(n1048), .Z(n25733) );
  NAND U26450 ( .A(n25734), .B(n25733), .Z(n25773) );
  NANDN U26451 ( .A(n1059), .B(a[153]), .Z(n25774) );
  XNOR U26452 ( .A(n25773), .B(n25774), .Z(n25776) );
  XOR U26453 ( .A(n25775), .B(n25776), .Z(n25815) );
  NANDN U26454 ( .A(n25735), .B(n38205), .Z(n25737) );
  XOR U26455 ( .A(b[23]), .B(n27178), .Z(n25869) );
  OR U26456 ( .A(n25869), .B(n38268), .Z(n25736) );
  NAND U26457 ( .A(n25737), .B(n25736), .Z(n25838) );
  XOR U26458 ( .A(b[7]), .B(a[179]), .Z(n25872) );
  NAND U26459 ( .A(n25872), .B(n36701), .Z(n25740) );
  NAND U26460 ( .A(n25738), .B(n36702), .Z(n25739) );
  NAND U26461 ( .A(n25740), .B(n25739), .Z(n25835) );
  XNOR U26462 ( .A(b[25]), .B(a[161]), .Z(n25875) );
  NANDN U26463 ( .A(n25875), .B(n38325), .Z(n25743) );
  NAND U26464 ( .A(n25741), .B(n38326), .Z(n25742) );
  AND U26465 ( .A(n25743), .B(n25742), .Z(n25836) );
  XNOR U26466 ( .A(n25835), .B(n25836), .Z(n25837) );
  XNOR U26467 ( .A(n25838), .B(n25837), .Z(n25816) );
  XOR U26468 ( .A(n25815), .B(n25816), .Z(n25818) );
  XNOR U26469 ( .A(n25817), .B(n25818), .Z(n25828) );
  XNOR U26470 ( .A(n25827), .B(n25828), .Z(n25878) );
  XNOR U26471 ( .A(n25879), .B(n25878), .Z(n25881) );
  XNOR U26472 ( .A(n25880), .B(n25881), .Z(n25894) );
  XOR U26473 ( .A(n25895), .B(n25894), .Z(n25896) );
  XNOR U26474 ( .A(n25897), .B(n25896), .Z(n25891) );
  NAND U26475 ( .A(n25745), .B(n25744), .Z(n25749) );
  NAND U26476 ( .A(n25747), .B(n25746), .Z(n25748) );
  NAND U26477 ( .A(n25749), .B(n25748), .Z(n25889) );
  NAND U26478 ( .A(n25751), .B(n25750), .Z(n25755) );
  NANDN U26479 ( .A(n25753), .B(n25752), .Z(n25754) );
  AND U26480 ( .A(n25755), .B(n25754), .Z(n25888) );
  XNOR U26481 ( .A(n25889), .B(n25888), .Z(n25890) );
  XOR U26482 ( .A(n25891), .B(n25890), .Z(n25770) );
  XOR U26483 ( .A(n25769), .B(n25770), .Z(n25761) );
  XOR U26484 ( .A(n25762), .B(n25761), .Z(n25763) );
  XNOR U26485 ( .A(n25764), .B(n25763), .Z(n25900) );
  XNOR U26486 ( .A(n25900), .B(sreg[409]), .Z(n25902) );
  NAND U26487 ( .A(n25756), .B(sreg[408]), .Z(n25760) );
  OR U26488 ( .A(n25758), .B(n25757), .Z(n25759) );
  AND U26489 ( .A(n25760), .B(n25759), .Z(n25901) );
  XOR U26490 ( .A(n25902), .B(n25901), .Z(c[409]) );
  NAND U26491 ( .A(n25762), .B(n25761), .Z(n25766) );
  NAND U26492 ( .A(n25764), .B(n25763), .Z(n25765) );
  NAND U26493 ( .A(n25766), .B(n25765), .Z(n25908) );
  NANDN U26494 ( .A(n25768), .B(n25767), .Z(n25772) );
  NAND U26495 ( .A(n25770), .B(n25769), .Z(n25771) );
  NAND U26496 ( .A(n25772), .B(n25771), .Z(n25906) );
  NANDN U26497 ( .A(n25774), .B(n25773), .Z(n25778) );
  NAND U26498 ( .A(n25776), .B(n25775), .Z(n25777) );
  NAND U26499 ( .A(n25778), .B(n25777), .Z(n25988) );
  XNOR U26500 ( .A(b[19]), .B(a[168]), .Z(n25955) );
  NANDN U26501 ( .A(n25955), .B(n37934), .Z(n25781) );
  NANDN U26502 ( .A(n25779), .B(n37935), .Z(n25780) );
  NAND U26503 ( .A(n25781), .B(n25780), .Z(n26024) );
  XOR U26504 ( .A(b[27]), .B(a[160]), .Z(n25958) );
  NAND U26505 ( .A(n38423), .B(n25958), .Z(n25784) );
  NAND U26506 ( .A(n25782), .B(n38424), .Z(n25783) );
  NAND U26507 ( .A(n25784), .B(n25783), .Z(n26021) );
  XNOR U26508 ( .A(b[5]), .B(a[182]), .Z(n25961) );
  NANDN U26509 ( .A(n25961), .B(n36587), .Z(n25787) );
  NANDN U26510 ( .A(n25785), .B(n36588), .Z(n25786) );
  AND U26511 ( .A(n25787), .B(n25786), .Z(n26022) );
  XNOR U26512 ( .A(n26021), .B(n26022), .Z(n26023) );
  XNOR U26513 ( .A(n26024), .B(n26023), .Z(n25985) );
  NAND U26514 ( .A(n25788), .B(n37762), .Z(n25790) );
  XOR U26515 ( .A(b[17]), .B(a[170]), .Z(n25964) );
  NAND U26516 ( .A(n25964), .B(n37764), .Z(n25789) );
  NAND U26517 ( .A(n25790), .B(n25789), .Z(n25939) );
  XNOR U26518 ( .A(b[31]), .B(a[156]), .Z(n25967) );
  NANDN U26519 ( .A(n25967), .B(n38552), .Z(n25793) );
  NANDN U26520 ( .A(n25791), .B(n38553), .Z(n25792) );
  AND U26521 ( .A(n25793), .B(n25792), .Z(n25937) );
  OR U26522 ( .A(n25794), .B(n36105), .Z(n25796) );
  XNOR U26523 ( .A(b[3]), .B(a[184]), .Z(n25970) );
  NANDN U26524 ( .A(n25970), .B(n36107), .Z(n25795) );
  AND U26525 ( .A(n25796), .B(n25795), .Z(n25938) );
  XOR U26526 ( .A(n25939), .B(n25940), .Z(n25986) );
  XOR U26527 ( .A(n25985), .B(n25986), .Z(n25987) );
  XNOR U26528 ( .A(n25988), .B(n25987), .Z(n26033) );
  NANDN U26529 ( .A(n25798), .B(n25797), .Z(n25802) );
  NAND U26530 ( .A(n25800), .B(n25799), .Z(n25801) );
  NAND U26531 ( .A(n25802), .B(n25801), .Z(n25976) );
  NANDN U26532 ( .A(n25804), .B(n25803), .Z(n25808) );
  NAND U26533 ( .A(n25806), .B(n25805), .Z(n25807) );
  NAND U26534 ( .A(n25808), .B(n25807), .Z(n25974) );
  OR U26535 ( .A(n25810), .B(n25809), .Z(n25814) );
  NANDN U26536 ( .A(n25812), .B(n25811), .Z(n25813) );
  NAND U26537 ( .A(n25814), .B(n25813), .Z(n25973) );
  XNOR U26538 ( .A(n25976), .B(n25975), .Z(n26034) );
  XNOR U26539 ( .A(n26033), .B(n26034), .Z(n26035) );
  NANDN U26540 ( .A(n25816), .B(n25815), .Z(n25820) );
  OR U26541 ( .A(n25818), .B(n25817), .Z(n25819) );
  AND U26542 ( .A(n25820), .B(n25819), .Z(n26036) );
  XNOR U26543 ( .A(n26035), .B(n26036), .Z(n25918) );
  NANDN U26544 ( .A(n25826), .B(n25825), .Z(n25830) );
  NANDN U26545 ( .A(n25828), .B(n25827), .Z(n25829) );
  NAND U26546 ( .A(n25830), .B(n25829), .Z(n26042) );
  NANDN U26547 ( .A(n25836), .B(n25835), .Z(n25840) );
  NAND U26548 ( .A(n25838), .B(n25837), .Z(n25839) );
  NAND U26549 ( .A(n25840), .B(n25839), .Z(n25979) );
  NANDN U26550 ( .A(n25842), .B(n25841), .Z(n25846) );
  NAND U26551 ( .A(n25844), .B(n25843), .Z(n25845) );
  AND U26552 ( .A(n25846), .B(n25845), .Z(n25980) );
  XNOR U26553 ( .A(n25979), .B(n25980), .Z(n25981) );
  XNOR U26554 ( .A(b[9]), .B(a[178]), .Z(n25991) );
  NANDN U26555 ( .A(n25991), .B(n36925), .Z(n25849) );
  NANDN U26556 ( .A(n25847), .B(n36926), .Z(n25848) );
  NAND U26557 ( .A(n25849), .B(n25848), .Z(n25945) );
  XNOR U26558 ( .A(b[15]), .B(a[172]), .Z(n25994) );
  OR U26559 ( .A(n25994), .B(n37665), .Z(n25852) );
  NANDN U26560 ( .A(n25850), .B(n37604), .Z(n25851) );
  AND U26561 ( .A(n25852), .B(n25851), .Z(n25943) );
  XNOR U26562 ( .A(b[21]), .B(a[166]), .Z(n25997) );
  NANDN U26563 ( .A(n25997), .B(n38101), .Z(n25855) );
  NANDN U26564 ( .A(n25853), .B(n38102), .Z(n25854) );
  AND U26565 ( .A(n25855), .B(n25854), .Z(n25944) );
  XOR U26566 ( .A(n25945), .B(n25946), .Z(n25934) );
  XNOR U26567 ( .A(b[11]), .B(a[176]), .Z(n26000) );
  OR U26568 ( .A(n26000), .B(n37311), .Z(n25858) );
  NANDN U26569 ( .A(n25856), .B(n37218), .Z(n25857) );
  NAND U26570 ( .A(n25858), .B(n25857), .Z(n25932) );
  XOR U26571 ( .A(n1053), .B(a[174]), .Z(n26003) );
  NANDN U26572 ( .A(n26003), .B(n37424), .Z(n25861) );
  NANDN U26573 ( .A(n25859), .B(n37425), .Z(n25860) );
  NAND U26574 ( .A(n25861), .B(n25860), .Z(n25931) );
  XOR U26575 ( .A(n25934), .B(n25933), .Z(n25928) );
  ANDN U26576 ( .B(b[31]), .A(n25862), .Z(n25949) );
  NANDN U26577 ( .A(n25863), .B(n38490), .Z(n25865) );
  XNOR U26578 ( .A(n1058), .B(a[158]), .Z(n26009) );
  NANDN U26579 ( .A(n1048), .B(n26009), .Z(n25864) );
  NAND U26580 ( .A(n25865), .B(n25864), .Z(n25950) );
  XOR U26581 ( .A(n25949), .B(n25950), .Z(n25951) );
  NANDN U26582 ( .A(n1049), .B(a[186]), .Z(n25866) );
  XNOR U26583 ( .A(b[1]), .B(n25866), .Z(n25868) );
  NANDN U26584 ( .A(b[0]), .B(a[185]), .Z(n25867) );
  AND U26585 ( .A(n25868), .B(n25867), .Z(n25952) );
  XNOR U26586 ( .A(n25951), .B(n25952), .Z(n25925) );
  NANDN U26587 ( .A(n25869), .B(n38205), .Z(n25871) );
  XNOR U26588 ( .A(b[23]), .B(a[164]), .Z(n26012) );
  OR U26589 ( .A(n26012), .B(n38268), .Z(n25870) );
  NAND U26590 ( .A(n25871), .B(n25870), .Z(n26030) );
  XOR U26591 ( .A(b[7]), .B(a[180]), .Z(n26015) );
  NAND U26592 ( .A(n26015), .B(n36701), .Z(n25874) );
  NAND U26593 ( .A(n25872), .B(n36702), .Z(n25873) );
  NAND U26594 ( .A(n25874), .B(n25873), .Z(n26027) );
  XOR U26595 ( .A(b[25]), .B(a[162]), .Z(n26018) );
  NAND U26596 ( .A(n26018), .B(n38325), .Z(n25877) );
  NANDN U26597 ( .A(n25875), .B(n38326), .Z(n25876) );
  AND U26598 ( .A(n25877), .B(n25876), .Z(n26028) );
  XNOR U26599 ( .A(n26027), .B(n26028), .Z(n26029) );
  XNOR U26600 ( .A(n26030), .B(n26029), .Z(n25926) );
  XOR U26601 ( .A(n25928), .B(n25927), .Z(n25982) );
  XNOR U26602 ( .A(n25981), .B(n25982), .Z(n26039) );
  XOR U26603 ( .A(n26040), .B(n26039), .Z(n26041) );
  XOR U26604 ( .A(n26042), .B(n26041), .Z(n25916) );
  XNOR U26605 ( .A(n25915), .B(n25916), .Z(n25917) );
  XNOR U26606 ( .A(n25918), .B(n25917), .Z(n25922) );
  NAND U26607 ( .A(n25879), .B(n25878), .Z(n25883) );
  NANDN U26608 ( .A(n25881), .B(n25880), .Z(n25882) );
  NAND U26609 ( .A(n25883), .B(n25882), .Z(n25919) );
  XNOR U26610 ( .A(n25919), .B(n25920), .Z(n25921) );
  XNOR U26611 ( .A(n25922), .B(n25921), .Z(n25912) );
  NANDN U26612 ( .A(n25889), .B(n25888), .Z(n25893) );
  NAND U26613 ( .A(n25891), .B(n25890), .Z(n25892) );
  NAND U26614 ( .A(n25893), .B(n25892), .Z(n25909) );
  NANDN U26615 ( .A(n25895), .B(n25894), .Z(n25899) );
  OR U26616 ( .A(n25897), .B(n25896), .Z(n25898) );
  NAND U26617 ( .A(n25899), .B(n25898), .Z(n25910) );
  XNOR U26618 ( .A(n25909), .B(n25910), .Z(n25911) );
  XNOR U26619 ( .A(n25912), .B(n25911), .Z(n25905) );
  XOR U26620 ( .A(n25906), .B(n25905), .Z(n25907) );
  XNOR U26621 ( .A(n25908), .B(n25907), .Z(n26045) );
  XNOR U26622 ( .A(n26045), .B(sreg[410]), .Z(n26047) );
  NAND U26623 ( .A(n25900), .B(sreg[409]), .Z(n25904) );
  OR U26624 ( .A(n25902), .B(n25901), .Z(n25903) );
  AND U26625 ( .A(n25904), .B(n25903), .Z(n26046) );
  XOR U26626 ( .A(n26047), .B(n26046), .Z(c[410]) );
  NANDN U26627 ( .A(n25910), .B(n25909), .Z(n25914) );
  NANDN U26628 ( .A(n25912), .B(n25911), .Z(n25913) );
  NAND U26629 ( .A(n25914), .B(n25913), .Z(n26051) );
  NANDN U26630 ( .A(n25920), .B(n25919), .Z(n25924) );
  NANDN U26631 ( .A(n25922), .B(n25921), .Z(n25923) );
  NAND U26632 ( .A(n25924), .B(n25923), .Z(n26057) );
  XNOR U26633 ( .A(n26056), .B(n26057), .Z(n26058) );
  OR U26634 ( .A(n25926), .B(n25925), .Z(n25930) );
  NANDN U26635 ( .A(n25928), .B(n25927), .Z(n25929) );
  NAND U26636 ( .A(n25930), .B(n25929), .Z(n26173) );
  OR U26637 ( .A(n25932), .B(n25931), .Z(n25936) );
  NAND U26638 ( .A(n25934), .B(n25933), .Z(n25935) );
  NAND U26639 ( .A(n25936), .B(n25935), .Z(n26112) );
  OR U26640 ( .A(n25938), .B(n25937), .Z(n25942) );
  NANDN U26641 ( .A(n25940), .B(n25939), .Z(n25941) );
  NAND U26642 ( .A(n25942), .B(n25941), .Z(n26111) );
  OR U26643 ( .A(n25944), .B(n25943), .Z(n25948) );
  NANDN U26644 ( .A(n25946), .B(n25945), .Z(n25947) );
  NAND U26645 ( .A(n25948), .B(n25947), .Z(n26110) );
  XOR U26646 ( .A(n26112), .B(n26113), .Z(n26171) );
  OR U26647 ( .A(n25950), .B(n25949), .Z(n25954) );
  NANDN U26648 ( .A(n25952), .B(n25951), .Z(n25953) );
  NAND U26649 ( .A(n25954), .B(n25953), .Z(n26125) );
  XNOR U26650 ( .A(b[19]), .B(a[169]), .Z(n26092) );
  NANDN U26651 ( .A(n26092), .B(n37934), .Z(n25957) );
  NANDN U26652 ( .A(n25955), .B(n37935), .Z(n25956) );
  NAND U26653 ( .A(n25957), .B(n25956), .Z(n26137) );
  XNOR U26654 ( .A(b[27]), .B(a[161]), .Z(n26095) );
  NANDN U26655 ( .A(n26095), .B(n38423), .Z(n25960) );
  NAND U26656 ( .A(n25958), .B(n38424), .Z(n25959) );
  NAND U26657 ( .A(n25960), .B(n25959), .Z(n26134) );
  XNOR U26658 ( .A(b[5]), .B(a[183]), .Z(n26098) );
  NANDN U26659 ( .A(n26098), .B(n36587), .Z(n25963) );
  NANDN U26660 ( .A(n25961), .B(n36588), .Z(n25962) );
  AND U26661 ( .A(n25963), .B(n25962), .Z(n26135) );
  XNOR U26662 ( .A(n26134), .B(n26135), .Z(n26136) );
  XNOR U26663 ( .A(n26137), .B(n26136), .Z(n26122) );
  NAND U26664 ( .A(n25964), .B(n37762), .Z(n25966) );
  XOR U26665 ( .A(b[17]), .B(a[171]), .Z(n26101) );
  NAND U26666 ( .A(n26101), .B(n37764), .Z(n25965) );
  NAND U26667 ( .A(n25966), .B(n25965), .Z(n26076) );
  XNOR U26668 ( .A(b[31]), .B(a[157]), .Z(n26104) );
  NANDN U26669 ( .A(n26104), .B(n38552), .Z(n25969) );
  NANDN U26670 ( .A(n25967), .B(n38553), .Z(n25968) );
  AND U26671 ( .A(n25969), .B(n25968), .Z(n26074) );
  OR U26672 ( .A(n25970), .B(n36105), .Z(n25972) );
  XNOR U26673 ( .A(b[3]), .B(a[185]), .Z(n26107) );
  NANDN U26674 ( .A(n26107), .B(n36107), .Z(n25971) );
  AND U26675 ( .A(n25972), .B(n25971), .Z(n26075) );
  XOR U26676 ( .A(n26076), .B(n26077), .Z(n26123) );
  XOR U26677 ( .A(n26122), .B(n26123), .Z(n26124) );
  XNOR U26678 ( .A(n26125), .B(n26124), .Z(n26170) );
  XOR U26679 ( .A(n26171), .B(n26170), .Z(n26172) );
  XNOR U26680 ( .A(n26173), .B(n26172), .Z(n26189) );
  OR U26681 ( .A(n25974), .B(n25973), .Z(n25978) );
  NAND U26682 ( .A(n25976), .B(n25975), .Z(n25977) );
  NAND U26683 ( .A(n25978), .B(n25977), .Z(n26187) );
  NANDN U26684 ( .A(n25980), .B(n25979), .Z(n25984) );
  NANDN U26685 ( .A(n25982), .B(n25981), .Z(n25983) );
  NAND U26686 ( .A(n25984), .B(n25983), .Z(n26177) );
  OR U26687 ( .A(n25986), .B(n25985), .Z(n25990) );
  NAND U26688 ( .A(n25988), .B(n25987), .Z(n25989) );
  NAND U26689 ( .A(n25990), .B(n25989), .Z(n26174) );
  XNOR U26690 ( .A(n1052), .B(a[179]), .Z(n26140) );
  NAND U26691 ( .A(n36925), .B(n26140), .Z(n25993) );
  NANDN U26692 ( .A(n25991), .B(n36926), .Z(n25992) );
  NAND U26693 ( .A(n25993), .B(n25992), .Z(n26082) );
  XNOR U26694 ( .A(b[15]), .B(a[173]), .Z(n26143) );
  OR U26695 ( .A(n26143), .B(n37665), .Z(n25996) );
  NANDN U26696 ( .A(n25994), .B(n37604), .Z(n25995) );
  AND U26697 ( .A(n25996), .B(n25995), .Z(n26080) );
  XNOR U26698 ( .A(n1056), .B(a[167]), .Z(n26146) );
  NAND U26699 ( .A(n26146), .B(n38101), .Z(n25999) );
  NANDN U26700 ( .A(n25997), .B(n38102), .Z(n25998) );
  AND U26701 ( .A(n25999), .B(n25998), .Z(n26081) );
  XOR U26702 ( .A(n26082), .B(n26083), .Z(n26071) );
  XNOR U26703 ( .A(b[11]), .B(a[177]), .Z(n26149) );
  OR U26704 ( .A(n26149), .B(n37311), .Z(n26002) );
  NANDN U26705 ( .A(n26000), .B(n37218), .Z(n26001) );
  NAND U26706 ( .A(n26002), .B(n26001), .Z(n26069) );
  XOR U26707 ( .A(n1053), .B(a[175]), .Z(n26152) );
  NANDN U26708 ( .A(n26152), .B(n37424), .Z(n26005) );
  NANDN U26709 ( .A(n26003), .B(n37425), .Z(n26004) );
  NAND U26710 ( .A(n26005), .B(n26004), .Z(n26068) );
  XOR U26711 ( .A(n26071), .B(n26070), .Z(n26065) );
  NANDN U26712 ( .A(n1049), .B(a[187]), .Z(n26006) );
  XNOR U26713 ( .A(b[1]), .B(n26006), .Z(n26008) );
  NANDN U26714 ( .A(b[0]), .B(a[186]), .Z(n26007) );
  AND U26715 ( .A(n26008), .B(n26007), .Z(n26088) );
  NAND U26716 ( .A(n26009), .B(n38490), .Z(n26011) );
  XNOR U26717 ( .A(n1058), .B(a[159]), .Z(n26158) );
  NANDN U26718 ( .A(n1048), .B(n26158), .Z(n26010) );
  NAND U26719 ( .A(n26011), .B(n26010), .Z(n26086) );
  NANDN U26720 ( .A(n1059), .B(a[155]), .Z(n26087) );
  XNOR U26721 ( .A(n26086), .B(n26087), .Z(n26089) );
  XNOR U26722 ( .A(n26088), .B(n26089), .Z(n26063) );
  NANDN U26723 ( .A(n26012), .B(n38205), .Z(n26014) );
  XNOR U26724 ( .A(b[23]), .B(a[165]), .Z(n26161) );
  OR U26725 ( .A(n26161), .B(n38268), .Z(n26013) );
  NAND U26726 ( .A(n26014), .B(n26013), .Z(n26131) );
  XOR U26727 ( .A(b[7]), .B(a[181]), .Z(n26164) );
  NAND U26728 ( .A(n26164), .B(n36701), .Z(n26017) );
  NAND U26729 ( .A(n26015), .B(n36702), .Z(n26016) );
  NAND U26730 ( .A(n26017), .B(n26016), .Z(n26128) );
  XNOR U26731 ( .A(b[25]), .B(a[163]), .Z(n26167) );
  NANDN U26732 ( .A(n26167), .B(n38325), .Z(n26020) );
  NAND U26733 ( .A(n26018), .B(n38326), .Z(n26019) );
  AND U26734 ( .A(n26020), .B(n26019), .Z(n26129) );
  XNOR U26735 ( .A(n26128), .B(n26129), .Z(n26130) );
  XOR U26736 ( .A(n26131), .B(n26130), .Z(n26062) );
  XNOR U26737 ( .A(n26065), .B(n26064), .Z(n26119) );
  NANDN U26738 ( .A(n26022), .B(n26021), .Z(n26026) );
  NAND U26739 ( .A(n26024), .B(n26023), .Z(n26025) );
  NAND U26740 ( .A(n26026), .B(n26025), .Z(n26117) );
  NANDN U26741 ( .A(n26028), .B(n26027), .Z(n26032) );
  NAND U26742 ( .A(n26030), .B(n26029), .Z(n26031) );
  AND U26743 ( .A(n26032), .B(n26031), .Z(n26116) );
  XNOR U26744 ( .A(n26117), .B(n26116), .Z(n26118) );
  XNOR U26745 ( .A(n26119), .B(n26118), .Z(n26175) );
  XNOR U26746 ( .A(n26174), .B(n26175), .Z(n26176) );
  XOR U26747 ( .A(n26177), .B(n26176), .Z(n26186) );
  XNOR U26748 ( .A(n26187), .B(n26186), .Z(n26188) );
  XOR U26749 ( .A(n26189), .B(n26188), .Z(n26183) );
  NANDN U26750 ( .A(n26034), .B(n26033), .Z(n26038) );
  NAND U26751 ( .A(n26036), .B(n26035), .Z(n26037) );
  NAND U26752 ( .A(n26038), .B(n26037), .Z(n26180) );
  NAND U26753 ( .A(n26040), .B(n26039), .Z(n26044) );
  NAND U26754 ( .A(n26042), .B(n26041), .Z(n26043) );
  NAND U26755 ( .A(n26044), .B(n26043), .Z(n26181) );
  XNOR U26756 ( .A(n26180), .B(n26181), .Z(n26182) );
  XOR U26757 ( .A(n26183), .B(n26182), .Z(n26059) );
  XOR U26758 ( .A(n26058), .B(n26059), .Z(n26050) );
  XOR U26759 ( .A(n26051), .B(n26050), .Z(n26052) );
  XNOR U26760 ( .A(n26053), .B(n26052), .Z(n26192) );
  XNOR U26761 ( .A(n26192), .B(sreg[411]), .Z(n26194) );
  NAND U26762 ( .A(n26045), .B(sreg[410]), .Z(n26049) );
  OR U26763 ( .A(n26047), .B(n26046), .Z(n26048) );
  AND U26764 ( .A(n26049), .B(n26048), .Z(n26193) );
  XOR U26765 ( .A(n26194), .B(n26193), .Z(c[411]) );
  NAND U26766 ( .A(n26051), .B(n26050), .Z(n26055) );
  NAND U26767 ( .A(n26053), .B(n26052), .Z(n26054) );
  NAND U26768 ( .A(n26055), .B(n26054), .Z(n26200) );
  NANDN U26769 ( .A(n26057), .B(n26056), .Z(n26061) );
  NAND U26770 ( .A(n26059), .B(n26058), .Z(n26060) );
  NAND U26771 ( .A(n26061), .B(n26060), .Z(n26198) );
  NANDN U26772 ( .A(n26063), .B(n26062), .Z(n26067) );
  NANDN U26773 ( .A(n26065), .B(n26064), .Z(n26066) );
  NAND U26774 ( .A(n26067), .B(n26066), .Z(n26328) );
  OR U26775 ( .A(n26069), .B(n26068), .Z(n26073) );
  NAND U26776 ( .A(n26071), .B(n26070), .Z(n26072) );
  NAND U26777 ( .A(n26073), .B(n26072), .Z(n26267) );
  OR U26778 ( .A(n26075), .B(n26074), .Z(n26079) );
  NANDN U26779 ( .A(n26077), .B(n26076), .Z(n26078) );
  NAND U26780 ( .A(n26079), .B(n26078), .Z(n26266) );
  OR U26781 ( .A(n26081), .B(n26080), .Z(n26085) );
  NANDN U26782 ( .A(n26083), .B(n26082), .Z(n26084) );
  NAND U26783 ( .A(n26085), .B(n26084), .Z(n26265) );
  XOR U26784 ( .A(n26267), .B(n26268), .Z(n26325) );
  NANDN U26785 ( .A(n26087), .B(n26086), .Z(n26091) );
  NAND U26786 ( .A(n26089), .B(n26088), .Z(n26090) );
  NAND U26787 ( .A(n26091), .B(n26090), .Z(n26280) );
  XNOR U26788 ( .A(b[19]), .B(a[170]), .Z(n26225) );
  NANDN U26789 ( .A(n26225), .B(n37934), .Z(n26094) );
  NANDN U26790 ( .A(n26092), .B(n37935), .Z(n26093) );
  NAND U26791 ( .A(n26094), .B(n26093), .Z(n26292) );
  XOR U26792 ( .A(b[27]), .B(a[162]), .Z(n26228) );
  NAND U26793 ( .A(n38423), .B(n26228), .Z(n26097) );
  NANDN U26794 ( .A(n26095), .B(n38424), .Z(n26096) );
  NAND U26795 ( .A(n26097), .B(n26096), .Z(n26289) );
  XNOR U26796 ( .A(b[5]), .B(a[184]), .Z(n26231) );
  NANDN U26797 ( .A(n26231), .B(n36587), .Z(n26100) );
  NANDN U26798 ( .A(n26098), .B(n36588), .Z(n26099) );
  AND U26799 ( .A(n26100), .B(n26099), .Z(n26290) );
  XNOR U26800 ( .A(n26289), .B(n26290), .Z(n26291) );
  XNOR U26801 ( .A(n26292), .B(n26291), .Z(n26278) );
  NAND U26802 ( .A(n26101), .B(n37762), .Z(n26103) );
  XOR U26803 ( .A(b[17]), .B(a[172]), .Z(n26234) );
  NAND U26804 ( .A(n26234), .B(n37764), .Z(n26102) );
  NAND U26805 ( .A(n26103), .B(n26102), .Z(n26252) );
  XNOR U26806 ( .A(b[31]), .B(a[158]), .Z(n26237) );
  NANDN U26807 ( .A(n26237), .B(n38552), .Z(n26106) );
  NANDN U26808 ( .A(n26104), .B(n38553), .Z(n26105) );
  NAND U26809 ( .A(n26106), .B(n26105), .Z(n26249) );
  OR U26810 ( .A(n26107), .B(n36105), .Z(n26109) );
  XNOR U26811 ( .A(b[3]), .B(a[186]), .Z(n26240) );
  NANDN U26812 ( .A(n26240), .B(n36107), .Z(n26108) );
  AND U26813 ( .A(n26109), .B(n26108), .Z(n26250) );
  XNOR U26814 ( .A(n26249), .B(n26250), .Z(n26251) );
  XOR U26815 ( .A(n26252), .B(n26251), .Z(n26277) );
  XNOR U26816 ( .A(n26278), .B(n26277), .Z(n26279) );
  XNOR U26817 ( .A(n26280), .B(n26279), .Z(n26326) );
  XNOR U26818 ( .A(n26325), .B(n26326), .Z(n26327) );
  XNOR U26819 ( .A(n26328), .B(n26327), .Z(n26216) );
  OR U26820 ( .A(n26111), .B(n26110), .Z(n26115) );
  NANDN U26821 ( .A(n26113), .B(n26112), .Z(n26114) );
  NAND U26822 ( .A(n26115), .B(n26114), .Z(n26214) );
  NANDN U26823 ( .A(n26117), .B(n26116), .Z(n26121) );
  NANDN U26824 ( .A(n26119), .B(n26118), .Z(n26120) );
  NAND U26825 ( .A(n26121), .B(n26120), .Z(n26334) );
  OR U26826 ( .A(n26123), .B(n26122), .Z(n26127) );
  NANDN U26827 ( .A(n26125), .B(n26124), .Z(n26126) );
  NAND U26828 ( .A(n26127), .B(n26126), .Z(n26332) );
  NANDN U26829 ( .A(n26129), .B(n26128), .Z(n26133) );
  NAND U26830 ( .A(n26131), .B(n26130), .Z(n26132) );
  NAND U26831 ( .A(n26133), .B(n26132), .Z(n26271) );
  NANDN U26832 ( .A(n26135), .B(n26134), .Z(n26139) );
  NAND U26833 ( .A(n26137), .B(n26136), .Z(n26138) );
  AND U26834 ( .A(n26139), .B(n26138), .Z(n26272) );
  XNOR U26835 ( .A(n26271), .B(n26272), .Z(n26273) );
  XOR U26836 ( .A(n1052), .B(a[180]), .Z(n26301) );
  NANDN U26837 ( .A(n26301), .B(n36925), .Z(n26142) );
  NAND U26838 ( .A(n36926), .B(n26140), .Z(n26141) );
  NAND U26839 ( .A(n26142), .B(n26141), .Z(n26257) );
  XNOR U26840 ( .A(n1054), .B(a[174]), .Z(n26298) );
  NANDN U26841 ( .A(n37665), .B(n26298), .Z(n26145) );
  NANDN U26842 ( .A(n26143), .B(n37604), .Z(n26144) );
  NAND U26843 ( .A(n26145), .B(n26144), .Z(n26255) );
  XOR U26844 ( .A(n1056), .B(a[168]), .Z(n26295) );
  NANDN U26845 ( .A(n26295), .B(n38101), .Z(n26148) );
  NAND U26846 ( .A(n38102), .B(n26146), .Z(n26147) );
  NAND U26847 ( .A(n26148), .B(n26147), .Z(n26256) );
  XNOR U26848 ( .A(n26255), .B(n26256), .Z(n26258) );
  XOR U26849 ( .A(n26257), .B(n26258), .Z(n26246) );
  XNOR U26850 ( .A(b[11]), .B(a[178]), .Z(n26304) );
  OR U26851 ( .A(n26304), .B(n37311), .Z(n26151) );
  NANDN U26852 ( .A(n26149), .B(n37218), .Z(n26150) );
  NAND U26853 ( .A(n26151), .B(n26150), .Z(n26244) );
  XOR U26854 ( .A(n1053), .B(a[176]), .Z(n26307) );
  NANDN U26855 ( .A(n26307), .B(n37424), .Z(n26154) );
  NANDN U26856 ( .A(n26152), .B(n37425), .Z(n26153) );
  AND U26857 ( .A(n26154), .B(n26153), .Z(n26243) );
  XNOR U26858 ( .A(n26244), .B(n26243), .Z(n26245) );
  XNOR U26859 ( .A(n26246), .B(n26245), .Z(n26262) );
  NANDN U26860 ( .A(n1049), .B(a[188]), .Z(n26155) );
  XNOR U26861 ( .A(b[1]), .B(n26155), .Z(n26157) );
  NANDN U26862 ( .A(b[0]), .B(a[187]), .Z(n26156) );
  AND U26863 ( .A(n26157), .B(n26156), .Z(n26221) );
  NAND U26864 ( .A(n38490), .B(n26158), .Z(n26160) );
  XNOR U26865 ( .A(n1058), .B(a[160]), .Z(n26310) );
  NANDN U26866 ( .A(n1048), .B(n26310), .Z(n26159) );
  NAND U26867 ( .A(n26160), .B(n26159), .Z(n26219) );
  NANDN U26868 ( .A(n1059), .B(a[156]), .Z(n26220) );
  XNOR U26869 ( .A(n26219), .B(n26220), .Z(n26222) );
  XNOR U26870 ( .A(n26221), .B(n26222), .Z(n26260) );
  NANDN U26871 ( .A(n26161), .B(n38205), .Z(n26163) );
  XNOR U26872 ( .A(b[23]), .B(a[166]), .Z(n26316) );
  OR U26873 ( .A(n26316), .B(n38268), .Z(n26162) );
  NAND U26874 ( .A(n26163), .B(n26162), .Z(n26286) );
  XOR U26875 ( .A(b[7]), .B(a[182]), .Z(n26319) );
  NAND U26876 ( .A(n26319), .B(n36701), .Z(n26166) );
  NAND U26877 ( .A(n26164), .B(n36702), .Z(n26165) );
  NAND U26878 ( .A(n26166), .B(n26165), .Z(n26283) );
  XOR U26879 ( .A(b[25]), .B(a[164]), .Z(n26322) );
  NAND U26880 ( .A(n26322), .B(n38325), .Z(n26169) );
  NANDN U26881 ( .A(n26167), .B(n38326), .Z(n26168) );
  AND U26882 ( .A(n26169), .B(n26168), .Z(n26284) );
  XNOR U26883 ( .A(n26283), .B(n26284), .Z(n26285) );
  XOR U26884 ( .A(n26286), .B(n26285), .Z(n26259) );
  XOR U26885 ( .A(n26262), .B(n26261), .Z(n26274) );
  XOR U26886 ( .A(n26273), .B(n26274), .Z(n26331) );
  XOR U26887 ( .A(n26332), .B(n26331), .Z(n26333) );
  XNOR U26888 ( .A(n26334), .B(n26333), .Z(n26213) );
  XNOR U26889 ( .A(n26214), .B(n26213), .Z(n26215) );
  XOR U26890 ( .A(n26216), .B(n26215), .Z(n26210) );
  NANDN U26891 ( .A(n26175), .B(n26174), .Z(n26179) );
  NAND U26892 ( .A(n26177), .B(n26176), .Z(n26178) );
  AND U26893 ( .A(n26179), .B(n26178), .Z(n26207) );
  XNOR U26894 ( .A(n26208), .B(n26207), .Z(n26209) );
  XNOR U26895 ( .A(n26210), .B(n26209), .Z(n26204) );
  NANDN U26896 ( .A(n26181), .B(n26180), .Z(n26185) );
  NAND U26897 ( .A(n26183), .B(n26182), .Z(n26184) );
  NAND U26898 ( .A(n26185), .B(n26184), .Z(n26201) );
  NANDN U26899 ( .A(n26187), .B(n26186), .Z(n26191) );
  NANDN U26900 ( .A(n26189), .B(n26188), .Z(n26190) );
  NAND U26901 ( .A(n26191), .B(n26190), .Z(n26202) );
  XNOR U26902 ( .A(n26201), .B(n26202), .Z(n26203) );
  XNOR U26903 ( .A(n26204), .B(n26203), .Z(n26197) );
  XOR U26904 ( .A(n26198), .B(n26197), .Z(n26199) );
  XNOR U26905 ( .A(n26200), .B(n26199), .Z(n26337) );
  XNOR U26906 ( .A(n26337), .B(sreg[412]), .Z(n26339) );
  NAND U26907 ( .A(n26192), .B(sreg[411]), .Z(n26196) );
  OR U26908 ( .A(n26194), .B(n26193), .Z(n26195) );
  AND U26909 ( .A(n26196), .B(n26195), .Z(n26338) );
  XOR U26910 ( .A(n26339), .B(n26338), .Z(c[412]) );
  NANDN U26911 ( .A(n26202), .B(n26201), .Z(n26206) );
  NANDN U26912 ( .A(n26204), .B(n26203), .Z(n26205) );
  NAND U26913 ( .A(n26206), .B(n26205), .Z(n26343) );
  NANDN U26914 ( .A(n26208), .B(n26207), .Z(n26212) );
  NAND U26915 ( .A(n26210), .B(n26209), .Z(n26211) );
  NAND U26916 ( .A(n26212), .B(n26211), .Z(n26348) );
  NANDN U26917 ( .A(n26214), .B(n26213), .Z(n26218) );
  NANDN U26918 ( .A(n26216), .B(n26215), .Z(n26217) );
  NAND U26919 ( .A(n26218), .B(n26217), .Z(n26349) );
  XNOR U26920 ( .A(n26348), .B(n26349), .Z(n26350) );
  NANDN U26921 ( .A(n26220), .B(n26219), .Z(n26224) );
  NAND U26922 ( .A(n26222), .B(n26221), .Z(n26223) );
  NAND U26923 ( .A(n26224), .B(n26223), .Z(n26423) );
  XNOR U26924 ( .A(b[19]), .B(a[171]), .Z(n26370) );
  NANDN U26925 ( .A(n26370), .B(n37934), .Z(n26227) );
  NANDN U26926 ( .A(n26225), .B(n37935), .Z(n26226) );
  NAND U26927 ( .A(n26227), .B(n26226), .Z(n26433) );
  XNOR U26928 ( .A(b[27]), .B(a[163]), .Z(n26373) );
  NANDN U26929 ( .A(n26373), .B(n38423), .Z(n26230) );
  NAND U26930 ( .A(n26228), .B(n38424), .Z(n26229) );
  NAND U26931 ( .A(n26230), .B(n26229), .Z(n26430) );
  XNOR U26932 ( .A(b[5]), .B(a[185]), .Z(n26376) );
  NANDN U26933 ( .A(n26376), .B(n36587), .Z(n26233) );
  NANDN U26934 ( .A(n26231), .B(n36588), .Z(n26232) );
  AND U26935 ( .A(n26233), .B(n26232), .Z(n26431) );
  XNOR U26936 ( .A(n26430), .B(n26431), .Z(n26432) );
  XNOR U26937 ( .A(n26433), .B(n26432), .Z(n26421) );
  NAND U26938 ( .A(n26234), .B(n37762), .Z(n26236) );
  XOR U26939 ( .A(b[17]), .B(a[173]), .Z(n26379) );
  NAND U26940 ( .A(n26379), .B(n37764), .Z(n26235) );
  NAND U26941 ( .A(n26236), .B(n26235), .Z(n26397) );
  XNOR U26942 ( .A(b[31]), .B(a[159]), .Z(n26382) );
  NANDN U26943 ( .A(n26382), .B(n38552), .Z(n26239) );
  NANDN U26944 ( .A(n26237), .B(n38553), .Z(n26238) );
  NAND U26945 ( .A(n26239), .B(n26238), .Z(n26394) );
  OR U26946 ( .A(n26240), .B(n36105), .Z(n26242) );
  XNOR U26947 ( .A(b[3]), .B(a[187]), .Z(n26385) );
  NANDN U26948 ( .A(n26385), .B(n36107), .Z(n26241) );
  AND U26949 ( .A(n26242), .B(n26241), .Z(n26395) );
  XNOR U26950 ( .A(n26394), .B(n26395), .Z(n26396) );
  XOR U26951 ( .A(n26397), .B(n26396), .Z(n26420) );
  XNOR U26952 ( .A(n26421), .B(n26420), .Z(n26422) );
  XNOR U26953 ( .A(n26423), .B(n26422), .Z(n26361) );
  NANDN U26954 ( .A(n26244), .B(n26243), .Z(n26248) );
  NAND U26955 ( .A(n26246), .B(n26245), .Z(n26247) );
  NAND U26956 ( .A(n26248), .B(n26247), .Z(n26412) );
  NANDN U26957 ( .A(n26250), .B(n26249), .Z(n26254) );
  NAND U26958 ( .A(n26252), .B(n26251), .Z(n26253) );
  NAND U26959 ( .A(n26254), .B(n26253), .Z(n26411) );
  XNOR U26960 ( .A(n26411), .B(n26410), .Z(n26413) );
  XOR U26961 ( .A(n26412), .B(n26413), .Z(n26360) );
  XOR U26962 ( .A(n26361), .B(n26360), .Z(n26362) );
  NANDN U26963 ( .A(n26260), .B(n26259), .Z(n26264) );
  NAND U26964 ( .A(n26262), .B(n26261), .Z(n26263) );
  NAND U26965 ( .A(n26264), .B(n26263), .Z(n26363) );
  XNOR U26966 ( .A(n26362), .B(n26363), .Z(n26474) );
  OR U26967 ( .A(n26266), .B(n26265), .Z(n26270) );
  NANDN U26968 ( .A(n26268), .B(n26267), .Z(n26269) );
  NAND U26969 ( .A(n26270), .B(n26269), .Z(n26473) );
  NANDN U26970 ( .A(n26272), .B(n26271), .Z(n26276) );
  NAND U26971 ( .A(n26274), .B(n26273), .Z(n26275) );
  NAND U26972 ( .A(n26276), .B(n26275), .Z(n26356) );
  NANDN U26973 ( .A(n26278), .B(n26277), .Z(n26282) );
  NAND U26974 ( .A(n26280), .B(n26279), .Z(n26281) );
  NAND U26975 ( .A(n26282), .B(n26281), .Z(n26355) );
  NANDN U26976 ( .A(n26284), .B(n26283), .Z(n26288) );
  NAND U26977 ( .A(n26286), .B(n26285), .Z(n26287) );
  NAND U26978 ( .A(n26288), .B(n26287), .Z(n26414) );
  NANDN U26979 ( .A(n26290), .B(n26289), .Z(n26294) );
  NAND U26980 ( .A(n26292), .B(n26291), .Z(n26293) );
  AND U26981 ( .A(n26294), .B(n26293), .Z(n26415) );
  XNOR U26982 ( .A(n26414), .B(n26415), .Z(n26416) );
  XOR U26983 ( .A(n1056), .B(a[169]), .Z(n26436) );
  NANDN U26984 ( .A(n26436), .B(n38101), .Z(n26297) );
  NANDN U26985 ( .A(n26295), .B(n38102), .Z(n26296) );
  NAND U26986 ( .A(n26297), .B(n26296), .Z(n26406) );
  XNOR U26987 ( .A(b[15]), .B(a[175]), .Z(n26439) );
  OR U26988 ( .A(n26439), .B(n37665), .Z(n26300) );
  NAND U26989 ( .A(n26298), .B(n37604), .Z(n26299) );
  AND U26990 ( .A(n26300), .B(n26299), .Z(n26407) );
  XNOR U26991 ( .A(n26406), .B(n26407), .Z(n26409) );
  XOR U26992 ( .A(n1052), .B(a[181]), .Z(n26442) );
  NANDN U26993 ( .A(n26442), .B(n36925), .Z(n26303) );
  NANDN U26994 ( .A(n26301), .B(n36926), .Z(n26302) );
  NAND U26995 ( .A(n26303), .B(n26302), .Z(n26408) );
  XNOR U26996 ( .A(n26409), .B(n26408), .Z(n26402) );
  XNOR U26997 ( .A(b[11]), .B(a[179]), .Z(n26445) );
  OR U26998 ( .A(n26445), .B(n37311), .Z(n26306) );
  NANDN U26999 ( .A(n26304), .B(n37218), .Z(n26305) );
  NAND U27000 ( .A(n26306), .B(n26305), .Z(n26401) );
  XOR U27001 ( .A(n1053), .B(a[177]), .Z(n26448) );
  NANDN U27002 ( .A(n26448), .B(n37424), .Z(n26309) );
  NANDN U27003 ( .A(n26307), .B(n37425), .Z(n26308) );
  NAND U27004 ( .A(n26309), .B(n26308), .Z(n26400) );
  XNOR U27005 ( .A(n26401), .B(n26400), .Z(n26403) );
  XNOR U27006 ( .A(n26402), .B(n26403), .Z(n26391) );
  NAND U27007 ( .A(n38490), .B(n26310), .Z(n26312) );
  XOR U27008 ( .A(n1058), .B(n26869), .Z(n26454) );
  NANDN U27009 ( .A(n1048), .B(n26454), .Z(n26311) );
  NAND U27010 ( .A(n26312), .B(n26311), .Z(n26364) );
  NANDN U27011 ( .A(n1059), .B(a[157]), .Z(n26365) );
  XNOR U27012 ( .A(n26364), .B(n26365), .Z(n26367) );
  NANDN U27013 ( .A(n1049), .B(a[189]), .Z(n26313) );
  XNOR U27014 ( .A(b[1]), .B(n26313), .Z(n26315) );
  NANDN U27015 ( .A(b[0]), .B(a[188]), .Z(n26314) );
  AND U27016 ( .A(n26315), .B(n26314), .Z(n26366) );
  XNOR U27017 ( .A(n26367), .B(n26366), .Z(n26389) );
  NANDN U27018 ( .A(n26316), .B(n38205), .Z(n26318) );
  XNOR U27019 ( .A(b[23]), .B(a[167]), .Z(n26457) );
  OR U27020 ( .A(n26457), .B(n38268), .Z(n26317) );
  NAND U27021 ( .A(n26318), .B(n26317), .Z(n26427) );
  XOR U27022 ( .A(b[7]), .B(a[183]), .Z(n26460) );
  NAND U27023 ( .A(n26460), .B(n36701), .Z(n26321) );
  NAND U27024 ( .A(n26319), .B(n36702), .Z(n26320) );
  NAND U27025 ( .A(n26321), .B(n26320), .Z(n26424) );
  XOR U27026 ( .A(b[25]), .B(a[165]), .Z(n26463) );
  NAND U27027 ( .A(n26463), .B(n38325), .Z(n26324) );
  NAND U27028 ( .A(n26322), .B(n38326), .Z(n26323) );
  AND U27029 ( .A(n26324), .B(n26323), .Z(n26425) );
  XNOR U27030 ( .A(n26424), .B(n26425), .Z(n26426) );
  XOR U27031 ( .A(n26427), .B(n26426), .Z(n26388) );
  XOR U27032 ( .A(n26391), .B(n26390), .Z(n26417) );
  XNOR U27033 ( .A(n26416), .B(n26417), .Z(n26354) );
  XNOR U27034 ( .A(n26355), .B(n26354), .Z(n26357) );
  XNOR U27035 ( .A(n26356), .B(n26357), .Z(n26472) );
  XOR U27036 ( .A(n26473), .B(n26472), .Z(n26475) );
  NANDN U27037 ( .A(n26326), .B(n26325), .Z(n26330) );
  NAND U27038 ( .A(n26328), .B(n26327), .Z(n26329) );
  NAND U27039 ( .A(n26330), .B(n26329), .Z(n26467) );
  NAND U27040 ( .A(n26332), .B(n26331), .Z(n26336) );
  NANDN U27041 ( .A(n26334), .B(n26333), .Z(n26335) );
  AND U27042 ( .A(n26336), .B(n26335), .Z(n26466) );
  XNOR U27043 ( .A(n26467), .B(n26466), .Z(n26468) );
  XOR U27044 ( .A(n26469), .B(n26468), .Z(n26351) );
  XOR U27045 ( .A(n26350), .B(n26351), .Z(n26342) );
  XOR U27046 ( .A(n26343), .B(n26342), .Z(n26344) );
  XNOR U27047 ( .A(n26345), .B(n26344), .Z(n26478) );
  XNOR U27048 ( .A(n26478), .B(sreg[413]), .Z(n26480) );
  NAND U27049 ( .A(n26337), .B(sreg[412]), .Z(n26341) );
  OR U27050 ( .A(n26339), .B(n26338), .Z(n26340) );
  AND U27051 ( .A(n26341), .B(n26340), .Z(n26479) );
  XOR U27052 ( .A(n26480), .B(n26479), .Z(c[413]) );
  NAND U27053 ( .A(n26343), .B(n26342), .Z(n26347) );
  NAND U27054 ( .A(n26345), .B(n26344), .Z(n26346) );
  NAND U27055 ( .A(n26347), .B(n26346), .Z(n26486) );
  NANDN U27056 ( .A(n26349), .B(n26348), .Z(n26353) );
  NAND U27057 ( .A(n26351), .B(n26350), .Z(n26352) );
  NAND U27058 ( .A(n26353), .B(n26352), .Z(n26483) );
  NAND U27059 ( .A(n26355), .B(n26354), .Z(n26359) );
  NANDN U27060 ( .A(n26357), .B(n26356), .Z(n26358) );
  NAND U27061 ( .A(n26359), .B(n26358), .Z(n26609) );
  XNOR U27062 ( .A(n26609), .B(n26610), .Z(n26611) );
  NANDN U27063 ( .A(n26365), .B(n26364), .Z(n26369) );
  NAND U27064 ( .A(n26367), .B(n26366), .Z(n26368) );
  NAND U27065 ( .A(n26369), .B(n26368), .Z(n26508) );
  XNOR U27066 ( .A(b[19]), .B(a[172]), .Z(n26557) );
  NANDN U27067 ( .A(n26557), .B(n37934), .Z(n26372) );
  NANDN U27068 ( .A(n26370), .B(n37935), .Z(n26371) );
  NAND U27069 ( .A(n26372), .B(n26371), .Z(n26542) );
  XOR U27070 ( .A(b[27]), .B(a[164]), .Z(n26560) );
  NAND U27071 ( .A(n38423), .B(n26560), .Z(n26375) );
  NANDN U27072 ( .A(n26373), .B(n38424), .Z(n26374) );
  NAND U27073 ( .A(n26375), .B(n26374), .Z(n26539) );
  XNOR U27074 ( .A(b[5]), .B(a[186]), .Z(n26563) );
  NANDN U27075 ( .A(n26563), .B(n36587), .Z(n26378) );
  NANDN U27076 ( .A(n26376), .B(n36588), .Z(n26377) );
  AND U27077 ( .A(n26378), .B(n26377), .Z(n26540) );
  XNOR U27078 ( .A(n26539), .B(n26540), .Z(n26541) );
  XNOR U27079 ( .A(n26542), .B(n26541), .Z(n26506) );
  NAND U27080 ( .A(n26379), .B(n37762), .Z(n26381) );
  XOR U27081 ( .A(b[17]), .B(a[174]), .Z(n26566) );
  NAND U27082 ( .A(n26566), .B(n37764), .Z(n26380) );
  NAND U27083 ( .A(n26381), .B(n26380), .Z(n26584) );
  XNOR U27084 ( .A(b[31]), .B(a[160]), .Z(n26569) );
  NANDN U27085 ( .A(n26569), .B(n38552), .Z(n26384) );
  NANDN U27086 ( .A(n26382), .B(n38553), .Z(n26383) );
  NAND U27087 ( .A(n26384), .B(n26383), .Z(n26581) );
  OR U27088 ( .A(n26385), .B(n36105), .Z(n26387) );
  XNOR U27089 ( .A(b[3]), .B(a[188]), .Z(n26572) );
  NANDN U27090 ( .A(n26572), .B(n36107), .Z(n26386) );
  AND U27091 ( .A(n26387), .B(n26386), .Z(n26582) );
  XNOR U27092 ( .A(n26581), .B(n26582), .Z(n26583) );
  XOR U27093 ( .A(n26584), .B(n26583), .Z(n26505) );
  XNOR U27094 ( .A(n26506), .B(n26505), .Z(n26507) );
  XNOR U27095 ( .A(n26508), .B(n26507), .Z(n26603) );
  NANDN U27096 ( .A(n26389), .B(n26388), .Z(n26393) );
  NANDN U27097 ( .A(n26391), .B(n26390), .Z(n26392) );
  NAND U27098 ( .A(n26393), .B(n26392), .Z(n26604) );
  XNOR U27099 ( .A(n26603), .B(n26604), .Z(n26605) );
  NANDN U27100 ( .A(n26395), .B(n26394), .Z(n26399) );
  NAND U27101 ( .A(n26397), .B(n26396), .Z(n26398) );
  NAND U27102 ( .A(n26399), .B(n26398), .Z(n26498) );
  OR U27103 ( .A(n26401), .B(n26400), .Z(n26405) );
  NANDN U27104 ( .A(n26403), .B(n26402), .Z(n26404) );
  NAND U27105 ( .A(n26405), .B(n26404), .Z(n26496) );
  XNOR U27106 ( .A(n26496), .B(n26495), .Z(n26497) );
  XOR U27107 ( .A(n26498), .B(n26497), .Z(n26606) );
  XOR U27108 ( .A(n26605), .B(n26606), .Z(n26617) );
  NANDN U27109 ( .A(n26415), .B(n26414), .Z(n26419) );
  NANDN U27110 ( .A(n26417), .B(n26416), .Z(n26418) );
  NAND U27111 ( .A(n26419), .B(n26418), .Z(n26600) );
  NANDN U27112 ( .A(n26425), .B(n26424), .Z(n26429) );
  NAND U27113 ( .A(n26427), .B(n26426), .Z(n26428) );
  NAND U27114 ( .A(n26429), .B(n26428), .Z(n26499) );
  NANDN U27115 ( .A(n26431), .B(n26430), .Z(n26435) );
  NAND U27116 ( .A(n26433), .B(n26432), .Z(n26434) );
  AND U27117 ( .A(n26435), .B(n26434), .Z(n26500) );
  XNOR U27118 ( .A(n26499), .B(n26500), .Z(n26501) );
  XNOR U27119 ( .A(b[21]), .B(a[170]), .Z(n26515) );
  NANDN U27120 ( .A(n26515), .B(n38101), .Z(n26438) );
  NANDN U27121 ( .A(n26436), .B(n38102), .Z(n26437) );
  NAND U27122 ( .A(n26438), .B(n26437), .Z(n26593) );
  XNOR U27123 ( .A(b[15]), .B(a[176]), .Z(n26512) );
  OR U27124 ( .A(n26512), .B(n37665), .Z(n26441) );
  NANDN U27125 ( .A(n26439), .B(n37604), .Z(n26440) );
  AND U27126 ( .A(n26441), .B(n26440), .Z(n26594) );
  XNOR U27127 ( .A(n26593), .B(n26594), .Z(n26596) );
  XNOR U27128 ( .A(b[9]), .B(a[182]), .Z(n26509) );
  NANDN U27129 ( .A(n26509), .B(n36925), .Z(n26444) );
  NANDN U27130 ( .A(n26442), .B(n36926), .Z(n26443) );
  NAND U27131 ( .A(n26444), .B(n26443), .Z(n26595) );
  XNOR U27132 ( .A(n26596), .B(n26595), .Z(n26589) );
  XNOR U27133 ( .A(b[11]), .B(a[180]), .Z(n26518) );
  OR U27134 ( .A(n26518), .B(n37311), .Z(n26447) );
  NANDN U27135 ( .A(n26445), .B(n37218), .Z(n26446) );
  NAND U27136 ( .A(n26447), .B(n26446), .Z(n26588) );
  XOR U27137 ( .A(n1053), .B(a[178]), .Z(n26521) );
  NANDN U27138 ( .A(n26521), .B(n37424), .Z(n26450) );
  NANDN U27139 ( .A(n26448), .B(n37425), .Z(n26449) );
  NAND U27140 ( .A(n26450), .B(n26449), .Z(n26587) );
  XNOR U27141 ( .A(n26588), .B(n26587), .Z(n26590) );
  XNOR U27142 ( .A(n26589), .B(n26590), .Z(n26578) );
  NANDN U27143 ( .A(n1049), .B(a[190]), .Z(n26451) );
  XNOR U27144 ( .A(b[1]), .B(n26451), .Z(n26453) );
  IV U27145 ( .A(a[189]), .Z(n30936) );
  NANDN U27146 ( .A(n30936), .B(n1049), .Z(n26452) );
  AND U27147 ( .A(n26453), .B(n26452), .Z(n26553) );
  NAND U27148 ( .A(n38490), .B(n26454), .Z(n26456) );
  XNOR U27149 ( .A(n1058), .B(a[162]), .Z(n26527) );
  NANDN U27150 ( .A(n1048), .B(n26527), .Z(n26455) );
  NAND U27151 ( .A(n26456), .B(n26455), .Z(n26551) );
  NANDN U27152 ( .A(n1059), .B(a[158]), .Z(n26552) );
  XNOR U27153 ( .A(n26551), .B(n26552), .Z(n26554) );
  XNOR U27154 ( .A(n26553), .B(n26554), .Z(n26576) );
  NANDN U27155 ( .A(n26457), .B(n38205), .Z(n26459) );
  XNOR U27156 ( .A(b[23]), .B(a[168]), .Z(n26530) );
  OR U27157 ( .A(n26530), .B(n38268), .Z(n26458) );
  NAND U27158 ( .A(n26459), .B(n26458), .Z(n26548) );
  XOR U27159 ( .A(b[7]), .B(a[184]), .Z(n26533) );
  NAND U27160 ( .A(n26533), .B(n36701), .Z(n26462) );
  NAND U27161 ( .A(n26460), .B(n36702), .Z(n26461) );
  NAND U27162 ( .A(n26462), .B(n26461), .Z(n26545) );
  XOR U27163 ( .A(b[25]), .B(a[166]), .Z(n26536) );
  NAND U27164 ( .A(n26536), .B(n38325), .Z(n26465) );
  NAND U27165 ( .A(n26463), .B(n38326), .Z(n26464) );
  AND U27166 ( .A(n26465), .B(n26464), .Z(n26546) );
  XNOR U27167 ( .A(n26545), .B(n26546), .Z(n26547) );
  XOR U27168 ( .A(n26548), .B(n26547), .Z(n26575) );
  XOR U27169 ( .A(n26578), .B(n26577), .Z(n26502) );
  XNOR U27170 ( .A(n26501), .B(n26502), .Z(n26597) );
  XOR U27171 ( .A(n26598), .B(n26597), .Z(n26599) );
  XNOR U27172 ( .A(n26600), .B(n26599), .Z(n26615) );
  XNOR U27173 ( .A(n26616), .B(n26615), .Z(n26618) );
  XNOR U27174 ( .A(n26617), .B(n26618), .Z(n26612) );
  XOR U27175 ( .A(n26611), .B(n26612), .Z(n26492) );
  NANDN U27176 ( .A(n26467), .B(n26466), .Z(n26471) );
  NAND U27177 ( .A(n26469), .B(n26468), .Z(n26470) );
  NAND U27178 ( .A(n26471), .B(n26470), .Z(n26489) );
  NANDN U27179 ( .A(n26473), .B(n26472), .Z(n26477) );
  OR U27180 ( .A(n26475), .B(n26474), .Z(n26476) );
  NAND U27181 ( .A(n26477), .B(n26476), .Z(n26490) );
  XNOR U27182 ( .A(n26489), .B(n26490), .Z(n26491) );
  XNOR U27183 ( .A(n26492), .B(n26491), .Z(n26484) );
  XNOR U27184 ( .A(n26483), .B(n26484), .Z(n26485) );
  XNOR U27185 ( .A(n26486), .B(n26485), .Z(n26621) );
  XNOR U27186 ( .A(n26621), .B(sreg[414]), .Z(n26623) );
  NAND U27187 ( .A(n26478), .B(sreg[413]), .Z(n26482) );
  OR U27188 ( .A(n26480), .B(n26479), .Z(n26481) );
  AND U27189 ( .A(n26482), .B(n26481), .Z(n26622) );
  XOR U27190 ( .A(n26623), .B(n26622), .Z(c[414]) );
  NANDN U27191 ( .A(n26484), .B(n26483), .Z(n26488) );
  NAND U27192 ( .A(n26486), .B(n26485), .Z(n26487) );
  NAND U27193 ( .A(n26488), .B(n26487), .Z(n26629) );
  NANDN U27194 ( .A(n26490), .B(n26489), .Z(n26494) );
  NAND U27195 ( .A(n26492), .B(n26491), .Z(n26493) );
  NAND U27196 ( .A(n26494), .B(n26493), .Z(n26627) );
  NANDN U27197 ( .A(n26500), .B(n26499), .Z(n26504) );
  NANDN U27198 ( .A(n26502), .B(n26501), .Z(n26503) );
  NAND U27199 ( .A(n26504), .B(n26503), .Z(n26743) );
  XNOR U27200 ( .A(b[9]), .B(a[183]), .Z(n26710) );
  NANDN U27201 ( .A(n26710), .B(n36925), .Z(n26511) );
  NANDN U27202 ( .A(n26509), .B(n36926), .Z(n26510) );
  NAND U27203 ( .A(n26511), .B(n26510), .Z(n26674) );
  XNOR U27204 ( .A(b[15]), .B(a[177]), .Z(n26713) );
  OR U27205 ( .A(n26713), .B(n37665), .Z(n26514) );
  NANDN U27206 ( .A(n26512), .B(n37604), .Z(n26513) );
  AND U27207 ( .A(n26514), .B(n26513), .Z(n26672) );
  XNOR U27208 ( .A(b[21]), .B(a[171]), .Z(n26716) );
  NANDN U27209 ( .A(n26716), .B(n38101), .Z(n26517) );
  NANDN U27210 ( .A(n26515), .B(n38102), .Z(n26516) );
  AND U27211 ( .A(n26517), .B(n26516), .Z(n26673) );
  XOR U27212 ( .A(n26674), .B(n26675), .Z(n26663) );
  XNOR U27213 ( .A(b[11]), .B(a[181]), .Z(n26719) );
  OR U27214 ( .A(n26719), .B(n37311), .Z(n26520) );
  NANDN U27215 ( .A(n26518), .B(n37218), .Z(n26519) );
  NAND U27216 ( .A(n26520), .B(n26519), .Z(n26661) );
  XOR U27217 ( .A(n1053), .B(a[179]), .Z(n26722) );
  NANDN U27218 ( .A(n26722), .B(n37424), .Z(n26523) );
  NANDN U27219 ( .A(n26521), .B(n37425), .Z(n26522) );
  AND U27220 ( .A(n26523), .B(n26522), .Z(n26660) );
  XNOR U27221 ( .A(n26661), .B(n26660), .Z(n26662) );
  XOR U27222 ( .A(n26663), .B(n26662), .Z(n26681) );
  NANDN U27223 ( .A(n1049), .B(a[191]), .Z(n26524) );
  XNOR U27224 ( .A(b[1]), .B(n26524), .Z(n26526) );
  NANDN U27225 ( .A(b[0]), .B(a[190]), .Z(n26525) );
  AND U27226 ( .A(n26526), .B(n26525), .Z(n26638) );
  NAND U27227 ( .A(n38490), .B(n26527), .Z(n26529) );
  XOR U27228 ( .A(n1058), .B(n27178), .Z(n26728) );
  NANDN U27229 ( .A(n1048), .B(n26728), .Z(n26528) );
  NAND U27230 ( .A(n26529), .B(n26528), .Z(n26636) );
  NANDN U27231 ( .A(n1059), .B(a[159]), .Z(n26637) );
  XNOR U27232 ( .A(n26636), .B(n26637), .Z(n26639) );
  XOR U27233 ( .A(n26638), .B(n26639), .Z(n26678) );
  NANDN U27234 ( .A(n26530), .B(n38205), .Z(n26532) );
  XNOR U27235 ( .A(b[23]), .B(a[169]), .Z(n26731) );
  OR U27236 ( .A(n26731), .B(n38268), .Z(n26531) );
  NAND U27237 ( .A(n26532), .B(n26531), .Z(n26701) );
  XOR U27238 ( .A(b[7]), .B(a[185]), .Z(n26734) );
  NAND U27239 ( .A(n26734), .B(n36701), .Z(n26535) );
  NAND U27240 ( .A(n26533), .B(n36702), .Z(n26534) );
  NAND U27241 ( .A(n26535), .B(n26534), .Z(n26698) );
  XOR U27242 ( .A(b[25]), .B(a[167]), .Z(n26737) );
  NAND U27243 ( .A(n26737), .B(n38325), .Z(n26538) );
  NAND U27244 ( .A(n26536), .B(n38326), .Z(n26537) );
  AND U27245 ( .A(n26538), .B(n26537), .Z(n26699) );
  XNOR U27246 ( .A(n26698), .B(n26699), .Z(n26700) );
  XNOR U27247 ( .A(n26701), .B(n26700), .Z(n26679) );
  XNOR U27248 ( .A(n26678), .B(n26679), .Z(n26680) );
  XNOR U27249 ( .A(n26681), .B(n26680), .Z(n26691) );
  NANDN U27250 ( .A(n26540), .B(n26539), .Z(n26544) );
  NAND U27251 ( .A(n26542), .B(n26541), .Z(n26543) );
  NAND U27252 ( .A(n26544), .B(n26543), .Z(n26689) );
  NANDN U27253 ( .A(n26546), .B(n26545), .Z(n26550) );
  NAND U27254 ( .A(n26548), .B(n26547), .Z(n26549) );
  AND U27255 ( .A(n26550), .B(n26549), .Z(n26688) );
  XNOR U27256 ( .A(n26689), .B(n26688), .Z(n26690) );
  XNOR U27257 ( .A(n26691), .B(n26690), .Z(n26741) );
  XNOR U27258 ( .A(n26740), .B(n26741), .Z(n26742) );
  XOR U27259 ( .A(n26743), .B(n26742), .Z(n26751) );
  XNOR U27260 ( .A(n26750), .B(n26751), .Z(n26753) );
  NANDN U27261 ( .A(n26552), .B(n26551), .Z(n26556) );
  NAND U27262 ( .A(n26554), .B(n26553), .Z(n26555) );
  NAND U27263 ( .A(n26556), .B(n26555), .Z(n26697) );
  XNOR U27264 ( .A(b[19]), .B(a[173]), .Z(n26642) );
  NANDN U27265 ( .A(n26642), .B(n37934), .Z(n26559) );
  NANDN U27266 ( .A(n26557), .B(n37935), .Z(n26558) );
  NAND U27267 ( .A(n26559), .B(n26558), .Z(n26707) );
  XOR U27268 ( .A(b[27]), .B(a[165]), .Z(n26645) );
  NAND U27269 ( .A(n38423), .B(n26645), .Z(n26562) );
  NAND U27270 ( .A(n26560), .B(n38424), .Z(n26561) );
  NAND U27271 ( .A(n26562), .B(n26561), .Z(n26704) );
  XNOR U27272 ( .A(b[5]), .B(a[187]), .Z(n26648) );
  NANDN U27273 ( .A(n26648), .B(n36587), .Z(n26565) );
  NANDN U27274 ( .A(n26563), .B(n36588), .Z(n26564) );
  AND U27275 ( .A(n26565), .B(n26564), .Z(n26705) );
  XNOR U27276 ( .A(n26704), .B(n26705), .Z(n26706) );
  XNOR U27277 ( .A(n26707), .B(n26706), .Z(n26695) );
  NAND U27278 ( .A(n26566), .B(n37762), .Z(n26568) );
  XOR U27279 ( .A(b[17]), .B(a[175]), .Z(n26651) );
  NAND U27280 ( .A(n26651), .B(n37764), .Z(n26567) );
  NAND U27281 ( .A(n26568), .B(n26567), .Z(n26669) );
  XOR U27282 ( .A(b[31]), .B(n26869), .Z(n26654) );
  NANDN U27283 ( .A(n26654), .B(n38552), .Z(n26571) );
  NANDN U27284 ( .A(n26569), .B(n38553), .Z(n26570) );
  NAND U27285 ( .A(n26571), .B(n26570), .Z(n26666) );
  OR U27286 ( .A(n26572), .B(n36105), .Z(n26574) );
  XOR U27287 ( .A(b[3]), .B(n30936), .Z(n26657) );
  NANDN U27288 ( .A(n26657), .B(n36107), .Z(n26573) );
  AND U27289 ( .A(n26574), .B(n26573), .Z(n26667) );
  XNOR U27290 ( .A(n26666), .B(n26667), .Z(n26668) );
  XOR U27291 ( .A(n26669), .B(n26668), .Z(n26694) );
  XNOR U27292 ( .A(n26695), .B(n26694), .Z(n26696) );
  XNOR U27293 ( .A(n26697), .B(n26696), .Z(n26746) );
  NANDN U27294 ( .A(n26576), .B(n26575), .Z(n26580) );
  NANDN U27295 ( .A(n26578), .B(n26577), .Z(n26579) );
  NAND U27296 ( .A(n26580), .B(n26579), .Z(n26747) );
  XNOR U27297 ( .A(n26746), .B(n26747), .Z(n26748) );
  NANDN U27298 ( .A(n26582), .B(n26581), .Z(n26586) );
  NAND U27299 ( .A(n26584), .B(n26583), .Z(n26585) );
  NAND U27300 ( .A(n26586), .B(n26585), .Z(n26687) );
  OR U27301 ( .A(n26588), .B(n26587), .Z(n26592) );
  NANDN U27302 ( .A(n26590), .B(n26589), .Z(n26591) );
  NAND U27303 ( .A(n26592), .B(n26591), .Z(n26685) );
  XNOR U27304 ( .A(n26685), .B(n26684), .Z(n26686) );
  XOR U27305 ( .A(n26687), .B(n26686), .Z(n26749) );
  XOR U27306 ( .A(n26748), .B(n26749), .Z(n26752) );
  XOR U27307 ( .A(n26753), .B(n26752), .Z(n26757) );
  NAND U27308 ( .A(n26598), .B(n26597), .Z(n26602) );
  NAND U27309 ( .A(n26600), .B(n26599), .Z(n26601) );
  NAND U27310 ( .A(n26602), .B(n26601), .Z(n26754) );
  NANDN U27311 ( .A(n26604), .B(n26603), .Z(n26608) );
  NAND U27312 ( .A(n26606), .B(n26605), .Z(n26607) );
  NAND U27313 ( .A(n26608), .B(n26607), .Z(n26755) );
  XNOR U27314 ( .A(n26754), .B(n26755), .Z(n26756) );
  XNOR U27315 ( .A(n26757), .B(n26756), .Z(n26633) );
  NANDN U27316 ( .A(n26610), .B(n26609), .Z(n26614) );
  NANDN U27317 ( .A(n26612), .B(n26611), .Z(n26613) );
  NAND U27318 ( .A(n26614), .B(n26613), .Z(n26631) );
  OR U27319 ( .A(n26616), .B(n26615), .Z(n26620) );
  OR U27320 ( .A(n26618), .B(n26617), .Z(n26619) );
  AND U27321 ( .A(n26620), .B(n26619), .Z(n26630) );
  XNOR U27322 ( .A(n26631), .B(n26630), .Z(n26632) );
  XNOR U27323 ( .A(n26633), .B(n26632), .Z(n26626) );
  XOR U27324 ( .A(n26627), .B(n26626), .Z(n26628) );
  XNOR U27325 ( .A(n26629), .B(n26628), .Z(n26760) );
  XNOR U27326 ( .A(n26760), .B(sreg[415]), .Z(n26762) );
  NAND U27327 ( .A(n26621), .B(sreg[414]), .Z(n26625) );
  OR U27328 ( .A(n26623), .B(n26622), .Z(n26624) );
  AND U27329 ( .A(n26625), .B(n26624), .Z(n26761) );
  XOR U27330 ( .A(n26762), .B(n26761), .Z(c[415]) );
  NANDN U27331 ( .A(n26631), .B(n26630), .Z(n26635) );
  NANDN U27332 ( .A(n26633), .B(n26632), .Z(n26634) );
  NAND U27333 ( .A(n26635), .B(n26634), .Z(n26766) );
  NANDN U27334 ( .A(n26637), .B(n26636), .Z(n26641) );
  NAND U27335 ( .A(n26639), .B(n26638), .Z(n26640) );
  NAND U27336 ( .A(n26641), .B(n26640), .Z(n26838) );
  XNOR U27337 ( .A(b[19]), .B(a[174]), .Z(n26781) );
  NANDN U27338 ( .A(n26781), .B(n37934), .Z(n26644) );
  NANDN U27339 ( .A(n26642), .B(n37935), .Z(n26643) );
  NAND U27340 ( .A(n26644), .B(n26643), .Z(n26848) );
  XOR U27341 ( .A(b[27]), .B(a[166]), .Z(n26784) );
  NAND U27342 ( .A(n38423), .B(n26784), .Z(n26647) );
  NAND U27343 ( .A(n26645), .B(n38424), .Z(n26646) );
  NAND U27344 ( .A(n26647), .B(n26646), .Z(n26845) );
  XNOR U27345 ( .A(b[5]), .B(a[188]), .Z(n26787) );
  NANDN U27346 ( .A(n26787), .B(n36587), .Z(n26650) );
  NANDN U27347 ( .A(n26648), .B(n36588), .Z(n26649) );
  AND U27348 ( .A(n26650), .B(n26649), .Z(n26846) );
  XNOR U27349 ( .A(n26845), .B(n26846), .Z(n26847) );
  XNOR U27350 ( .A(n26848), .B(n26847), .Z(n26836) );
  NAND U27351 ( .A(n26651), .B(n37762), .Z(n26653) );
  XOR U27352 ( .A(b[17]), .B(a[176]), .Z(n26790) );
  NAND U27353 ( .A(n26790), .B(n37764), .Z(n26652) );
  NAND U27354 ( .A(n26653), .B(n26652), .Z(n26808) );
  XNOR U27355 ( .A(b[31]), .B(a[162]), .Z(n26793) );
  NANDN U27356 ( .A(n26793), .B(n38552), .Z(n26656) );
  NANDN U27357 ( .A(n26654), .B(n38553), .Z(n26655) );
  NAND U27358 ( .A(n26656), .B(n26655), .Z(n26805) );
  OR U27359 ( .A(n26657), .B(n36105), .Z(n26659) );
  XNOR U27360 ( .A(b[3]), .B(a[190]), .Z(n26796) );
  NANDN U27361 ( .A(n26796), .B(n36107), .Z(n26658) );
  AND U27362 ( .A(n26659), .B(n26658), .Z(n26806) );
  XNOR U27363 ( .A(n26805), .B(n26806), .Z(n26807) );
  XOR U27364 ( .A(n26808), .B(n26807), .Z(n26835) );
  XNOR U27365 ( .A(n26836), .B(n26835), .Z(n26837) );
  XNOR U27366 ( .A(n26838), .B(n26837), .Z(n26882) );
  NANDN U27367 ( .A(n26661), .B(n26660), .Z(n26665) );
  NAND U27368 ( .A(n26663), .B(n26662), .Z(n26664) );
  NAND U27369 ( .A(n26665), .B(n26664), .Z(n26826) );
  NANDN U27370 ( .A(n26667), .B(n26666), .Z(n26671) );
  NAND U27371 ( .A(n26669), .B(n26668), .Z(n26670) );
  NAND U27372 ( .A(n26671), .B(n26670), .Z(n26824) );
  OR U27373 ( .A(n26673), .B(n26672), .Z(n26677) );
  NANDN U27374 ( .A(n26675), .B(n26674), .Z(n26676) );
  NAND U27375 ( .A(n26677), .B(n26676), .Z(n26823) );
  XNOR U27376 ( .A(n26826), .B(n26825), .Z(n26883) );
  XNOR U27377 ( .A(n26882), .B(n26883), .Z(n26884) );
  NANDN U27378 ( .A(n26679), .B(n26678), .Z(n26683) );
  NANDN U27379 ( .A(n26681), .B(n26680), .Z(n26682) );
  AND U27380 ( .A(n26683), .B(n26682), .Z(n26885) );
  XNOR U27381 ( .A(n26884), .B(n26885), .Z(n26897) );
  NANDN U27382 ( .A(n26689), .B(n26688), .Z(n26693) );
  NANDN U27383 ( .A(n26691), .B(n26690), .Z(n26692) );
  NAND U27384 ( .A(n26693), .B(n26692), .Z(n26891) );
  NANDN U27385 ( .A(n26699), .B(n26698), .Z(n26703) );
  NAND U27386 ( .A(n26701), .B(n26700), .Z(n26702) );
  NAND U27387 ( .A(n26703), .B(n26702), .Z(n26829) );
  NANDN U27388 ( .A(n26705), .B(n26704), .Z(n26709) );
  NAND U27389 ( .A(n26707), .B(n26706), .Z(n26708) );
  AND U27390 ( .A(n26709), .B(n26708), .Z(n26830) );
  XNOR U27391 ( .A(n26829), .B(n26830), .Z(n26831) );
  XNOR U27392 ( .A(b[9]), .B(a[184]), .Z(n26851) );
  NANDN U27393 ( .A(n26851), .B(n36925), .Z(n26712) );
  NANDN U27394 ( .A(n26710), .B(n36926), .Z(n26711) );
  NAND U27395 ( .A(n26712), .B(n26711), .Z(n26813) );
  XNOR U27396 ( .A(b[15]), .B(a[178]), .Z(n26854) );
  OR U27397 ( .A(n26854), .B(n37665), .Z(n26715) );
  NANDN U27398 ( .A(n26713), .B(n37604), .Z(n26714) );
  AND U27399 ( .A(n26715), .B(n26714), .Z(n26811) );
  XNOR U27400 ( .A(b[21]), .B(a[172]), .Z(n26857) );
  NANDN U27401 ( .A(n26857), .B(n38101), .Z(n26718) );
  NANDN U27402 ( .A(n26716), .B(n38102), .Z(n26717) );
  AND U27403 ( .A(n26718), .B(n26717), .Z(n26812) );
  XOR U27404 ( .A(n26813), .B(n26814), .Z(n26802) );
  XNOR U27405 ( .A(b[11]), .B(a[182]), .Z(n26860) );
  OR U27406 ( .A(n26860), .B(n37311), .Z(n26721) );
  NANDN U27407 ( .A(n26719), .B(n37218), .Z(n26720) );
  NAND U27408 ( .A(n26721), .B(n26720), .Z(n26800) );
  XOR U27409 ( .A(n1053), .B(a[180]), .Z(n26863) );
  NANDN U27410 ( .A(n26863), .B(n37424), .Z(n26724) );
  NANDN U27411 ( .A(n26722), .B(n37425), .Z(n26723) );
  AND U27412 ( .A(n26724), .B(n26723), .Z(n26799) );
  XNOR U27413 ( .A(n26800), .B(n26799), .Z(n26801) );
  XOR U27414 ( .A(n26802), .B(n26801), .Z(n26819) );
  NANDN U27415 ( .A(n1049), .B(a[192]), .Z(n26725) );
  XNOR U27416 ( .A(b[1]), .B(n26725), .Z(n26727) );
  NANDN U27417 ( .A(b[0]), .B(a[191]), .Z(n26726) );
  AND U27418 ( .A(n26727), .B(n26726), .Z(n26777) );
  NAND U27419 ( .A(n38490), .B(n26728), .Z(n26730) );
  XNOR U27420 ( .A(b[29]), .B(a[164]), .Z(n26870) );
  OR U27421 ( .A(n26870), .B(n1048), .Z(n26729) );
  NAND U27422 ( .A(n26730), .B(n26729), .Z(n26775) );
  NANDN U27423 ( .A(n1059), .B(a[160]), .Z(n26776) );
  XNOR U27424 ( .A(n26775), .B(n26776), .Z(n26778) );
  XOR U27425 ( .A(n26777), .B(n26778), .Z(n26817) );
  NANDN U27426 ( .A(n26731), .B(n38205), .Z(n26733) );
  XNOR U27427 ( .A(b[23]), .B(a[170]), .Z(n26873) );
  OR U27428 ( .A(n26873), .B(n38268), .Z(n26732) );
  NAND U27429 ( .A(n26733), .B(n26732), .Z(n26842) );
  XOR U27430 ( .A(b[7]), .B(a[186]), .Z(n26876) );
  NAND U27431 ( .A(n26876), .B(n36701), .Z(n26736) );
  NAND U27432 ( .A(n26734), .B(n36702), .Z(n26735) );
  NAND U27433 ( .A(n26736), .B(n26735), .Z(n26839) );
  XOR U27434 ( .A(b[25]), .B(a[168]), .Z(n26879) );
  NAND U27435 ( .A(n26879), .B(n38325), .Z(n26739) );
  NAND U27436 ( .A(n26737), .B(n38326), .Z(n26738) );
  AND U27437 ( .A(n26739), .B(n26738), .Z(n26840) );
  XNOR U27438 ( .A(n26839), .B(n26840), .Z(n26841) );
  XNOR U27439 ( .A(n26842), .B(n26841), .Z(n26818) );
  XOR U27440 ( .A(n26817), .B(n26818), .Z(n26820) );
  XNOR U27441 ( .A(n26819), .B(n26820), .Z(n26832) );
  XNOR U27442 ( .A(n26831), .B(n26832), .Z(n26888) );
  XNOR U27443 ( .A(n26889), .B(n26888), .Z(n26890) );
  XOR U27444 ( .A(n26891), .B(n26890), .Z(n26895) );
  XNOR U27445 ( .A(n26894), .B(n26895), .Z(n26896) );
  XNOR U27446 ( .A(n26897), .B(n26896), .Z(n26901) );
  NANDN U27447 ( .A(n26741), .B(n26740), .Z(n26745) );
  NAND U27448 ( .A(n26743), .B(n26742), .Z(n26744) );
  NAND U27449 ( .A(n26745), .B(n26744), .Z(n26898) );
  XNOR U27450 ( .A(n26898), .B(n26899), .Z(n26900) );
  XNOR U27451 ( .A(n26901), .B(n26900), .Z(n26772) );
  NANDN U27452 ( .A(n26755), .B(n26754), .Z(n26759) );
  NANDN U27453 ( .A(n26757), .B(n26756), .Z(n26758) );
  NAND U27454 ( .A(n26759), .B(n26758), .Z(n26770) );
  XNOR U27455 ( .A(n26769), .B(n26770), .Z(n26771) );
  XNOR U27456 ( .A(n26772), .B(n26771), .Z(n26765) );
  XOR U27457 ( .A(n26766), .B(n26765), .Z(n26767) );
  XNOR U27458 ( .A(n26768), .B(n26767), .Z(n26904) );
  XNOR U27459 ( .A(n26904), .B(sreg[416]), .Z(n26906) );
  NAND U27460 ( .A(n26760), .B(sreg[415]), .Z(n26764) );
  OR U27461 ( .A(n26762), .B(n26761), .Z(n26763) );
  AND U27462 ( .A(n26764), .B(n26763), .Z(n26905) );
  XOR U27463 ( .A(n26906), .B(n26905), .Z(c[416]) );
  NANDN U27464 ( .A(n26770), .B(n26769), .Z(n26774) );
  NANDN U27465 ( .A(n26772), .B(n26771), .Z(n26773) );
  NAND U27466 ( .A(n26774), .B(n26773), .Z(n26910) );
  NANDN U27467 ( .A(n26776), .B(n26775), .Z(n26780) );
  NAND U27468 ( .A(n26778), .B(n26777), .Z(n26779) );
  NAND U27469 ( .A(n26780), .B(n26779), .Z(n26996) );
  XNOR U27470 ( .A(b[19]), .B(a[175]), .Z(n26963) );
  NANDN U27471 ( .A(n26963), .B(n37934), .Z(n26783) );
  NANDN U27472 ( .A(n26781), .B(n37935), .Z(n26782) );
  NAND U27473 ( .A(n26783), .B(n26782), .Z(n27008) );
  XOR U27474 ( .A(b[27]), .B(a[167]), .Z(n26966) );
  NAND U27475 ( .A(n38423), .B(n26966), .Z(n26786) );
  NAND U27476 ( .A(n26784), .B(n38424), .Z(n26785) );
  NAND U27477 ( .A(n26786), .B(n26785), .Z(n27005) );
  XOR U27478 ( .A(b[5]), .B(n30936), .Z(n26969) );
  NANDN U27479 ( .A(n26969), .B(n36587), .Z(n26789) );
  NANDN U27480 ( .A(n26787), .B(n36588), .Z(n26788) );
  AND U27481 ( .A(n26789), .B(n26788), .Z(n27006) );
  XNOR U27482 ( .A(n27005), .B(n27006), .Z(n27007) );
  XNOR U27483 ( .A(n27008), .B(n27007), .Z(n26993) );
  NAND U27484 ( .A(n26790), .B(n37762), .Z(n26792) );
  XOR U27485 ( .A(b[17]), .B(a[177]), .Z(n26972) );
  NAND U27486 ( .A(n26972), .B(n37764), .Z(n26791) );
  NAND U27487 ( .A(n26792), .B(n26791), .Z(n26947) );
  XOR U27488 ( .A(b[31]), .B(n27178), .Z(n26975) );
  NANDN U27489 ( .A(n26975), .B(n38552), .Z(n26795) );
  NANDN U27490 ( .A(n26793), .B(n38553), .Z(n26794) );
  AND U27491 ( .A(n26795), .B(n26794), .Z(n26945) );
  OR U27492 ( .A(n26796), .B(n36105), .Z(n26798) );
  XNOR U27493 ( .A(b[3]), .B(a[191]), .Z(n26978) );
  NANDN U27494 ( .A(n26978), .B(n36107), .Z(n26797) );
  AND U27495 ( .A(n26798), .B(n26797), .Z(n26946) );
  XOR U27496 ( .A(n26947), .B(n26948), .Z(n26994) );
  XOR U27497 ( .A(n26993), .B(n26994), .Z(n26995) );
  XNOR U27498 ( .A(n26996), .B(n26995), .Z(n27041) );
  NANDN U27499 ( .A(n26800), .B(n26799), .Z(n26804) );
  NAND U27500 ( .A(n26802), .B(n26801), .Z(n26803) );
  NAND U27501 ( .A(n26804), .B(n26803), .Z(n26984) );
  NANDN U27502 ( .A(n26806), .B(n26805), .Z(n26810) );
  NAND U27503 ( .A(n26808), .B(n26807), .Z(n26809) );
  NAND U27504 ( .A(n26810), .B(n26809), .Z(n26982) );
  OR U27505 ( .A(n26812), .B(n26811), .Z(n26816) );
  NANDN U27506 ( .A(n26814), .B(n26813), .Z(n26815) );
  NAND U27507 ( .A(n26816), .B(n26815), .Z(n26981) );
  XNOR U27508 ( .A(n26984), .B(n26983), .Z(n27042) );
  XOR U27509 ( .A(n27041), .B(n27042), .Z(n27044) );
  NANDN U27510 ( .A(n26818), .B(n26817), .Z(n26822) );
  OR U27511 ( .A(n26820), .B(n26819), .Z(n26821) );
  NAND U27512 ( .A(n26822), .B(n26821), .Z(n27043) );
  XOR U27513 ( .A(n27044), .B(n27043), .Z(n26929) );
  OR U27514 ( .A(n26824), .B(n26823), .Z(n26828) );
  NAND U27515 ( .A(n26826), .B(n26825), .Z(n26827) );
  NAND U27516 ( .A(n26828), .B(n26827), .Z(n26928) );
  NANDN U27517 ( .A(n26830), .B(n26829), .Z(n26834) );
  NANDN U27518 ( .A(n26832), .B(n26831), .Z(n26833) );
  NAND U27519 ( .A(n26834), .B(n26833), .Z(n27049) );
  NANDN U27520 ( .A(n26840), .B(n26839), .Z(n26844) );
  NAND U27521 ( .A(n26842), .B(n26841), .Z(n26843) );
  NAND U27522 ( .A(n26844), .B(n26843), .Z(n26987) );
  NANDN U27523 ( .A(n26846), .B(n26845), .Z(n26850) );
  NAND U27524 ( .A(n26848), .B(n26847), .Z(n26849) );
  AND U27525 ( .A(n26850), .B(n26849), .Z(n26988) );
  XNOR U27526 ( .A(n26987), .B(n26988), .Z(n26989) );
  XNOR U27527 ( .A(b[9]), .B(a[185]), .Z(n27011) );
  NANDN U27528 ( .A(n27011), .B(n36925), .Z(n26853) );
  NANDN U27529 ( .A(n26851), .B(n36926), .Z(n26852) );
  NAND U27530 ( .A(n26853), .B(n26852), .Z(n26953) );
  XNOR U27531 ( .A(b[15]), .B(a[179]), .Z(n27014) );
  OR U27532 ( .A(n27014), .B(n37665), .Z(n26856) );
  NANDN U27533 ( .A(n26854), .B(n37604), .Z(n26855) );
  AND U27534 ( .A(n26856), .B(n26855), .Z(n26951) );
  XNOR U27535 ( .A(b[21]), .B(a[173]), .Z(n27017) );
  NANDN U27536 ( .A(n27017), .B(n38101), .Z(n26859) );
  NANDN U27537 ( .A(n26857), .B(n38102), .Z(n26858) );
  AND U27538 ( .A(n26859), .B(n26858), .Z(n26952) );
  XOR U27539 ( .A(n26953), .B(n26954), .Z(n26942) );
  XNOR U27540 ( .A(b[11]), .B(a[183]), .Z(n27020) );
  OR U27541 ( .A(n27020), .B(n37311), .Z(n26862) );
  NANDN U27542 ( .A(n26860), .B(n37218), .Z(n26861) );
  NAND U27543 ( .A(n26862), .B(n26861), .Z(n26940) );
  XOR U27544 ( .A(n1053), .B(a[181]), .Z(n27023) );
  NANDN U27545 ( .A(n27023), .B(n37424), .Z(n26865) );
  NANDN U27546 ( .A(n26863), .B(n37425), .Z(n26864) );
  NAND U27547 ( .A(n26865), .B(n26864), .Z(n26939) );
  XOR U27548 ( .A(n26942), .B(n26941), .Z(n26936) );
  NANDN U27549 ( .A(n1049), .B(a[193]), .Z(n26866) );
  XNOR U27550 ( .A(b[1]), .B(n26866), .Z(n26868) );
  NANDN U27551 ( .A(b[0]), .B(a[192]), .Z(n26867) );
  AND U27552 ( .A(n26868), .B(n26867), .Z(n26960) );
  ANDN U27553 ( .B(b[31]), .A(n26869), .Z(n26957) );
  NANDN U27554 ( .A(n26870), .B(n38490), .Z(n26872) );
  XNOR U27555 ( .A(n1058), .B(a[165]), .Z(n27029) );
  NANDN U27556 ( .A(n1048), .B(n27029), .Z(n26871) );
  NAND U27557 ( .A(n26872), .B(n26871), .Z(n26958) );
  XOR U27558 ( .A(n26957), .B(n26958), .Z(n26959) );
  XNOR U27559 ( .A(n26960), .B(n26959), .Z(n26933) );
  NANDN U27560 ( .A(n26873), .B(n38205), .Z(n26875) );
  XNOR U27561 ( .A(b[23]), .B(a[171]), .Z(n27032) );
  OR U27562 ( .A(n27032), .B(n38268), .Z(n26874) );
  NAND U27563 ( .A(n26875), .B(n26874), .Z(n27002) );
  XOR U27564 ( .A(b[7]), .B(a[187]), .Z(n27035) );
  NAND U27565 ( .A(n27035), .B(n36701), .Z(n26878) );
  NAND U27566 ( .A(n26876), .B(n36702), .Z(n26877) );
  NAND U27567 ( .A(n26878), .B(n26877), .Z(n26999) );
  XOR U27568 ( .A(b[25]), .B(a[169]), .Z(n27038) );
  NAND U27569 ( .A(n27038), .B(n38325), .Z(n26881) );
  NAND U27570 ( .A(n26879), .B(n38326), .Z(n26880) );
  AND U27571 ( .A(n26881), .B(n26880), .Z(n27000) );
  XNOR U27572 ( .A(n26999), .B(n27000), .Z(n27001) );
  XNOR U27573 ( .A(n27002), .B(n27001), .Z(n26934) );
  XOR U27574 ( .A(n26936), .B(n26935), .Z(n26990) );
  XNOR U27575 ( .A(n26989), .B(n26990), .Z(n27047) );
  XNOR U27576 ( .A(n27048), .B(n27047), .Z(n27050) );
  XNOR U27577 ( .A(n27049), .B(n27050), .Z(n26927) );
  XOR U27578 ( .A(n26928), .B(n26927), .Z(n26930) );
  NANDN U27579 ( .A(n26883), .B(n26882), .Z(n26887) );
  NAND U27580 ( .A(n26885), .B(n26884), .Z(n26886) );
  NAND U27581 ( .A(n26887), .B(n26886), .Z(n26921) );
  NAND U27582 ( .A(n26889), .B(n26888), .Z(n26893) );
  OR U27583 ( .A(n26891), .B(n26890), .Z(n26892) );
  NAND U27584 ( .A(n26893), .B(n26892), .Z(n26922) );
  XNOR U27585 ( .A(n26921), .B(n26922), .Z(n26923) );
  XOR U27586 ( .A(n26924), .B(n26923), .Z(n26917) );
  NANDN U27587 ( .A(n26899), .B(n26898), .Z(n26903) );
  NANDN U27588 ( .A(n26901), .B(n26900), .Z(n26902) );
  NAND U27589 ( .A(n26903), .B(n26902), .Z(n26916) );
  XNOR U27590 ( .A(n26915), .B(n26916), .Z(n26918) );
  XOR U27591 ( .A(n26917), .B(n26918), .Z(n26909) );
  XOR U27592 ( .A(n26910), .B(n26909), .Z(n26911) );
  XNOR U27593 ( .A(n26912), .B(n26911), .Z(n27053) );
  XNOR U27594 ( .A(n27053), .B(sreg[417]), .Z(n27055) );
  NAND U27595 ( .A(n26904), .B(sreg[416]), .Z(n26908) );
  OR U27596 ( .A(n26906), .B(n26905), .Z(n26907) );
  AND U27597 ( .A(n26908), .B(n26907), .Z(n27054) );
  XOR U27598 ( .A(n27055), .B(n27054), .Z(c[417]) );
  NAND U27599 ( .A(n26910), .B(n26909), .Z(n26914) );
  NAND U27600 ( .A(n26912), .B(n26911), .Z(n26913) );
  NAND U27601 ( .A(n26914), .B(n26913), .Z(n27061) );
  NANDN U27602 ( .A(n26916), .B(n26915), .Z(n26920) );
  NAND U27603 ( .A(n26918), .B(n26917), .Z(n26919) );
  NAND U27604 ( .A(n26920), .B(n26919), .Z(n27059) );
  NANDN U27605 ( .A(n26922), .B(n26921), .Z(n26926) );
  NAND U27606 ( .A(n26924), .B(n26923), .Z(n26925) );
  NAND U27607 ( .A(n26926), .B(n26925), .Z(n27064) );
  NANDN U27608 ( .A(n26928), .B(n26927), .Z(n26932) );
  OR U27609 ( .A(n26930), .B(n26929), .Z(n26931) );
  NAND U27610 ( .A(n26932), .B(n26931), .Z(n27065) );
  XNOR U27611 ( .A(n27064), .B(n27065), .Z(n27066) );
  OR U27612 ( .A(n26934), .B(n26933), .Z(n26938) );
  NANDN U27613 ( .A(n26936), .B(n26935), .Z(n26937) );
  NAND U27614 ( .A(n26938), .B(n26937), .Z(n27194) );
  OR U27615 ( .A(n26940), .B(n26939), .Z(n26944) );
  NAND U27616 ( .A(n26942), .B(n26941), .Z(n26943) );
  NAND U27617 ( .A(n26944), .B(n26943), .Z(n27132) );
  OR U27618 ( .A(n26946), .B(n26945), .Z(n26950) );
  NANDN U27619 ( .A(n26948), .B(n26947), .Z(n26949) );
  NAND U27620 ( .A(n26950), .B(n26949), .Z(n27131) );
  OR U27621 ( .A(n26952), .B(n26951), .Z(n26956) );
  NANDN U27622 ( .A(n26954), .B(n26953), .Z(n26955) );
  NAND U27623 ( .A(n26956), .B(n26955), .Z(n27130) );
  XOR U27624 ( .A(n27132), .B(n27133), .Z(n27192) );
  OR U27625 ( .A(n26958), .B(n26957), .Z(n26962) );
  NANDN U27626 ( .A(n26960), .B(n26959), .Z(n26961) );
  NAND U27627 ( .A(n26962), .B(n26961), .Z(n27144) );
  XNOR U27628 ( .A(b[19]), .B(a[176]), .Z(n27088) );
  NANDN U27629 ( .A(n27088), .B(n37934), .Z(n26965) );
  NANDN U27630 ( .A(n26963), .B(n37935), .Z(n26964) );
  NAND U27631 ( .A(n26965), .B(n26964), .Z(n27157) );
  XOR U27632 ( .A(b[27]), .B(a[168]), .Z(n27091) );
  NAND U27633 ( .A(n38423), .B(n27091), .Z(n26968) );
  NAND U27634 ( .A(n26966), .B(n38424), .Z(n26967) );
  NAND U27635 ( .A(n26968), .B(n26967), .Z(n27154) );
  XNOR U27636 ( .A(b[5]), .B(a[190]), .Z(n27094) );
  NANDN U27637 ( .A(n27094), .B(n36587), .Z(n26971) );
  NANDN U27638 ( .A(n26969), .B(n36588), .Z(n26970) );
  AND U27639 ( .A(n26971), .B(n26970), .Z(n27155) );
  XNOR U27640 ( .A(n27154), .B(n27155), .Z(n27156) );
  XNOR U27641 ( .A(n27157), .B(n27156), .Z(n27143) );
  NAND U27642 ( .A(n26972), .B(n37762), .Z(n26974) );
  XOR U27643 ( .A(b[17]), .B(a[178]), .Z(n27097) );
  NAND U27644 ( .A(n27097), .B(n37764), .Z(n26973) );
  NAND U27645 ( .A(n26974), .B(n26973), .Z(n27115) );
  XNOR U27646 ( .A(b[31]), .B(a[164]), .Z(n27100) );
  NANDN U27647 ( .A(n27100), .B(n38552), .Z(n26977) );
  NANDN U27648 ( .A(n26975), .B(n38553), .Z(n26976) );
  NAND U27649 ( .A(n26977), .B(n26976), .Z(n27112) );
  OR U27650 ( .A(n26978), .B(n36105), .Z(n26980) );
  XNOR U27651 ( .A(b[3]), .B(a[192]), .Z(n27103) );
  NANDN U27652 ( .A(n27103), .B(n36107), .Z(n26979) );
  AND U27653 ( .A(n26980), .B(n26979), .Z(n27113) );
  XNOR U27654 ( .A(n27112), .B(n27113), .Z(n27114) );
  XOR U27655 ( .A(n27115), .B(n27114), .Z(n27142) );
  XOR U27656 ( .A(n27143), .B(n27142), .Z(n27145) );
  XOR U27657 ( .A(n27144), .B(n27145), .Z(n27191) );
  XOR U27658 ( .A(n27192), .B(n27191), .Z(n27193) );
  XNOR U27659 ( .A(n27194), .B(n27193), .Z(n27079) );
  OR U27660 ( .A(n26982), .B(n26981), .Z(n26986) );
  NAND U27661 ( .A(n26984), .B(n26983), .Z(n26985) );
  NAND U27662 ( .A(n26986), .B(n26985), .Z(n27077) );
  NANDN U27663 ( .A(n26988), .B(n26987), .Z(n26992) );
  NANDN U27664 ( .A(n26990), .B(n26989), .Z(n26991) );
  NAND U27665 ( .A(n26992), .B(n26991), .Z(n27199) );
  OR U27666 ( .A(n26994), .B(n26993), .Z(n26998) );
  NAND U27667 ( .A(n26996), .B(n26995), .Z(n26997) );
  NAND U27668 ( .A(n26998), .B(n26997), .Z(n27198) );
  NANDN U27669 ( .A(n27000), .B(n26999), .Z(n27004) );
  NAND U27670 ( .A(n27002), .B(n27001), .Z(n27003) );
  NAND U27671 ( .A(n27004), .B(n27003), .Z(n27136) );
  NANDN U27672 ( .A(n27006), .B(n27005), .Z(n27010) );
  NAND U27673 ( .A(n27008), .B(n27007), .Z(n27009) );
  AND U27674 ( .A(n27010), .B(n27009), .Z(n27137) );
  XNOR U27675 ( .A(n27136), .B(n27137), .Z(n27138) );
  XNOR U27676 ( .A(b[9]), .B(a[186]), .Z(n27160) );
  NANDN U27677 ( .A(n27160), .B(n36925), .Z(n27013) );
  NANDN U27678 ( .A(n27011), .B(n36926), .Z(n27012) );
  NAND U27679 ( .A(n27013), .B(n27012), .Z(n27120) );
  XNOR U27680 ( .A(b[15]), .B(a[180]), .Z(n27163) );
  OR U27681 ( .A(n27163), .B(n37665), .Z(n27016) );
  NANDN U27682 ( .A(n27014), .B(n37604), .Z(n27015) );
  AND U27683 ( .A(n27016), .B(n27015), .Z(n27118) );
  XNOR U27684 ( .A(b[21]), .B(a[174]), .Z(n27166) );
  NANDN U27685 ( .A(n27166), .B(n38101), .Z(n27019) );
  NANDN U27686 ( .A(n27017), .B(n38102), .Z(n27018) );
  AND U27687 ( .A(n27019), .B(n27018), .Z(n27119) );
  XOR U27688 ( .A(n27120), .B(n27121), .Z(n27109) );
  XNOR U27689 ( .A(b[11]), .B(a[184]), .Z(n27169) );
  OR U27690 ( .A(n27169), .B(n37311), .Z(n27022) );
  NANDN U27691 ( .A(n27020), .B(n37218), .Z(n27021) );
  NAND U27692 ( .A(n27022), .B(n27021), .Z(n27107) );
  XOR U27693 ( .A(n1053), .B(a[182]), .Z(n27172) );
  NANDN U27694 ( .A(n27172), .B(n37424), .Z(n27025) );
  NANDN U27695 ( .A(n27023), .B(n37425), .Z(n27024) );
  AND U27696 ( .A(n27025), .B(n27024), .Z(n27106) );
  XNOR U27697 ( .A(n27107), .B(n27106), .Z(n27108) );
  XOR U27698 ( .A(n27109), .B(n27108), .Z(n27126) );
  NANDN U27699 ( .A(n1049), .B(a[194]), .Z(n27026) );
  XNOR U27700 ( .A(b[1]), .B(n27026), .Z(n27028) );
  IV U27701 ( .A(a[193]), .Z(n31508) );
  NANDN U27702 ( .A(n31508), .B(n1049), .Z(n27027) );
  AND U27703 ( .A(n27028), .B(n27027), .Z(n27084) );
  NAND U27704 ( .A(n27029), .B(n38490), .Z(n27031) );
  XNOR U27705 ( .A(b[29]), .B(a[166]), .Z(n27179) );
  OR U27706 ( .A(n27179), .B(n1048), .Z(n27030) );
  NAND U27707 ( .A(n27031), .B(n27030), .Z(n27082) );
  NANDN U27708 ( .A(n1059), .B(a[162]), .Z(n27083) );
  XNOR U27709 ( .A(n27082), .B(n27083), .Z(n27085) );
  XOR U27710 ( .A(n27084), .B(n27085), .Z(n27124) );
  NANDN U27711 ( .A(n27032), .B(n38205), .Z(n27034) );
  XNOR U27712 ( .A(b[23]), .B(a[172]), .Z(n27182) );
  OR U27713 ( .A(n27182), .B(n38268), .Z(n27033) );
  NAND U27714 ( .A(n27034), .B(n27033), .Z(n27151) );
  XOR U27715 ( .A(b[7]), .B(a[188]), .Z(n27185) );
  NAND U27716 ( .A(n27185), .B(n36701), .Z(n27037) );
  NAND U27717 ( .A(n27035), .B(n36702), .Z(n27036) );
  NAND U27718 ( .A(n27037), .B(n27036), .Z(n27148) );
  XOR U27719 ( .A(b[25]), .B(a[170]), .Z(n27188) );
  NAND U27720 ( .A(n27188), .B(n38325), .Z(n27040) );
  NAND U27721 ( .A(n27038), .B(n38326), .Z(n27039) );
  AND U27722 ( .A(n27040), .B(n27039), .Z(n27149) );
  XNOR U27723 ( .A(n27148), .B(n27149), .Z(n27150) );
  XNOR U27724 ( .A(n27151), .B(n27150), .Z(n27125) );
  XOR U27725 ( .A(n27124), .B(n27125), .Z(n27127) );
  XNOR U27726 ( .A(n27126), .B(n27127), .Z(n27139) );
  XNOR U27727 ( .A(n27138), .B(n27139), .Z(n27197) );
  XNOR U27728 ( .A(n27198), .B(n27197), .Z(n27200) );
  XNOR U27729 ( .A(n27199), .B(n27200), .Z(n27076) );
  XNOR U27730 ( .A(n27077), .B(n27076), .Z(n27078) );
  XOR U27731 ( .A(n27079), .B(n27078), .Z(n27073) );
  NANDN U27732 ( .A(n27042), .B(n27041), .Z(n27046) );
  OR U27733 ( .A(n27044), .B(n27043), .Z(n27045) );
  NAND U27734 ( .A(n27046), .B(n27045), .Z(n27070) );
  NAND U27735 ( .A(n27048), .B(n27047), .Z(n27052) );
  NANDN U27736 ( .A(n27050), .B(n27049), .Z(n27051) );
  NAND U27737 ( .A(n27052), .B(n27051), .Z(n27071) );
  XNOR U27738 ( .A(n27070), .B(n27071), .Z(n27072) );
  XOR U27739 ( .A(n27073), .B(n27072), .Z(n27067) );
  XOR U27740 ( .A(n27066), .B(n27067), .Z(n27058) );
  XOR U27741 ( .A(n27059), .B(n27058), .Z(n27060) );
  XNOR U27742 ( .A(n27061), .B(n27060), .Z(n27203) );
  XNOR U27743 ( .A(n27203), .B(sreg[418]), .Z(n27205) );
  NAND U27744 ( .A(n27053), .B(sreg[417]), .Z(n27057) );
  OR U27745 ( .A(n27055), .B(n27054), .Z(n27056) );
  AND U27746 ( .A(n27057), .B(n27056), .Z(n27204) );
  XOR U27747 ( .A(n27205), .B(n27204), .Z(c[418]) );
  NAND U27748 ( .A(n27059), .B(n27058), .Z(n27063) );
  NAND U27749 ( .A(n27061), .B(n27060), .Z(n27062) );
  NAND U27750 ( .A(n27063), .B(n27062), .Z(n27211) );
  NANDN U27751 ( .A(n27065), .B(n27064), .Z(n27069) );
  NAND U27752 ( .A(n27067), .B(n27066), .Z(n27068) );
  NAND U27753 ( .A(n27069), .B(n27068), .Z(n27209) );
  NANDN U27754 ( .A(n27071), .B(n27070), .Z(n27075) );
  NAND U27755 ( .A(n27073), .B(n27072), .Z(n27074) );
  NAND U27756 ( .A(n27075), .B(n27074), .Z(n27214) );
  NANDN U27757 ( .A(n27077), .B(n27076), .Z(n27081) );
  NANDN U27758 ( .A(n27079), .B(n27078), .Z(n27080) );
  NAND U27759 ( .A(n27081), .B(n27080), .Z(n27215) );
  XNOR U27760 ( .A(n27214), .B(n27215), .Z(n27216) );
  NANDN U27761 ( .A(n27083), .B(n27082), .Z(n27087) );
  NAND U27762 ( .A(n27085), .B(n27084), .Z(n27086) );
  NAND U27763 ( .A(n27087), .B(n27086), .Z(n27283) );
  XNOR U27764 ( .A(b[19]), .B(a[177]), .Z(n27250) );
  NANDN U27765 ( .A(n27250), .B(n37934), .Z(n27090) );
  NANDN U27766 ( .A(n27088), .B(n37935), .Z(n27089) );
  NAND U27767 ( .A(n27090), .B(n27089), .Z(n27295) );
  XOR U27768 ( .A(b[27]), .B(a[169]), .Z(n27253) );
  NAND U27769 ( .A(n38423), .B(n27253), .Z(n27093) );
  NAND U27770 ( .A(n27091), .B(n38424), .Z(n27092) );
  NAND U27771 ( .A(n27093), .B(n27092), .Z(n27292) );
  XNOR U27772 ( .A(b[5]), .B(a[191]), .Z(n27256) );
  NANDN U27773 ( .A(n27256), .B(n36587), .Z(n27096) );
  NANDN U27774 ( .A(n27094), .B(n36588), .Z(n27095) );
  AND U27775 ( .A(n27096), .B(n27095), .Z(n27293) );
  XNOR U27776 ( .A(n27292), .B(n27293), .Z(n27294) );
  XNOR U27777 ( .A(n27295), .B(n27294), .Z(n27280) );
  NAND U27778 ( .A(n27097), .B(n37762), .Z(n27099) );
  XOR U27779 ( .A(b[17]), .B(a[179]), .Z(n27259) );
  NAND U27780 ( .A(n27259), .B(n37764), .Z(n27098) );
  NAND U27781 ( .A(n27099), .B(n27098), .Z(n27234) );
  XNOR U27782 ( .A(b[31]), .B(a[165]), .Z(n27262) );
  NANDN U27783 ( .A(n27262), .B(n38552), .Z(n27102) );
  NANDN U27784 ( .A(n27100), .B(n38553), .Z(n27101) );
  AND U27785 ( .A(n27102), .B(n27101), .Z(n27232) );
  OR U27786 ( .A(n27103), .B(n36105), .Z(n27105) );
  XOR U27787 ( .A(b[3]), .B(n31508), .Z(n27265) );
  NANDN U27788 ( .A(n27265), .B(n36107), .Z(n27104) );
  AND U27789 ( .A(n27105), .B(n27104), .Z(n27233) );
  XOR U27790 ( .A(n27234), .B(n27235), .Z(n27281) );
  XOR U27791 ( .A(n27280), .B(n27281), .Z(n27282) );
  XNOR U27792 ( .A(n27283), .B(n27282), .Z(n27328) );
  NANDN U27793 ( .A(n27107), .B(n27106), .Z(n27111) );
  NAND U27794 ( .A(n27109), .B(n27108), .Z(n27110) );
  NAND U27795 ( .A(n27111), .B(n27110), .Z(n27271) );
  NANDN U27796 ( .A(n27113), .B(n27112), .Z(n27117) );
  NAND U27797 ( .A(n27115), .B(n27114), .Z(n27116) );
  NAND U27798 ( .A(n27117), .B(n27116), .Z(n27269) );
  OR U27799 ( .A(n27119), .B(n27118), .Z(n27123) );
  NANDN U27800 ( .A(n27121), .B(n27120), .Z(n27122) );
  NAND U27801 ( .A(n27123), .B(n27122), .Z(n27268) );
  XNOR U27802 ( .A(n27271), .B(n27270), .Z(n27329) );
  XOR U27803 ( .A(n27328), .B(n27329), .Z(n27331) );
  NANDN U27804 ( .A(n27125), .B(n27124), .Z(n27129) );
  OR U27805 ( .A(n27127), .B(n27126), .Z(n27128) );
  NAND U27806 ( .A(n27129), .B(n27128), .Z(n27330) );
  XOR U27807 ( .A(n27331), .B(n27330), .Z(n27348) );
  OR U27808 ( .A(n27131), .B(n27130), .Z(n27135) );
  NANDN U27809 ( .A(n27133), .B(n27132), .Z(n27134) );
  NAND U27810 ( .A(n27135), .B(n27134), .Z(n27347) );
  NANDN U27811 ( .A(n27137), .B(n27136), .Z(n27141) );
  NANDN U27812 ( .A(n27139), .B(n27138), .Z(n27140) );
  NAND U27813 ( .A(n27141), .B(n27140), .Z(n27336) );
  NANDN U27814 ( .A(n27143), .B(n27142), .Z(n27147) );
  OR U27815 ( .A(n27145), .B(n27144), .Z(n27146) );
  NAND U27816 ( .A(n27147), .B(n27146), .Z(n27335) );
  NANDN U27817 ( .A(n27149), .B(n27148), .Z(n27153) );
  NAND U27818 ( .A(n27151), .B(n27150), .Z(n27152) );
  NAND U27819 ( .A(n27153), .B(n27152), .Z(n27274) );
  NANDN U27820 ( .A(n27155), .B(n27154), .Z(n27159) );
  NAND U27821 ( .A(n27157), .B(n27156), .Z(n27158) );
  AND U27822 ( .A(n27159), .B(n27158), .Z(n27275) );
  XNOR U27823 ( .A(n27274), .B(n27275), .Z(n27276) );
  XNOR U27824 ( .A(b[9]), .B(a[187]), .Z(n27298) );
  NANDN U27825 ( .A(n27298), .B(n36925), .Z(n27162) );
  NANDN U27826 ( .A(n27160), .B(n36926), .Z(n27161) );
  NAND U27827 ( .A(n27162), .B(n27161), .Z(n27240) );
  XNOR U27828 ( .A(b[15]), .B(a[181]), .Z(n27301) );
  OR U27829 ( .A(n27301), .B(n37665), .Z(n27165) );
  NANDN U27830 ( .A(n27163), .B(n37604), .Z(n27164) );
  AND U27831 ( .A(n27165), .B(n27164), .Z(n27238) );
  XNOR U27832 ( .A(b[21]), .B(a[175]), .Z(n27304) );
  NANDN U27833 ( .A(n27304), .B(n38101), .Z(n27168) );
  NANDN U27834 ( .A(n27166), .B(n38102), .Z(n27167) );
  AND U27835 ( .A(n27168), .B(n27167), .Z(n27239) );
  XOR U27836 ( .A(n27240), .B(n27241), .Z(n27229) );
  XNOR U27837 ( .A(b[11]), .B(a[185]), .Z(n27307) );
  OR U27838 ( .A(n27307), .B(n37311), .Z(n27171) );
  NANDN U27839 ( .A(n27169), .B(n37218), .Z(n27170) );
  NAND U27840 ( .A(n27171), .B(n27170), .Z(n27227) );
  XOR U27841 ( .A(n1053), .B(a[183]), .Z(n27310) );
  NANDN U27842 ( .A(n27310), .B(n37424), .Z(n27174) );
  NANDN U27843 ( .A(n27172), .B(n37425), .Z(n27173) );
  NAND U27844 ( .A(n27174), .B(n27173), .Z(n27226) );
  XOR U27845 ( .A(n27229), .B(n27228), .Z(n27223) );
  ANDN U27846 ( .B(a[195]), .A(n1049), .Z(n27175) );
  XOR U27847 ( .A(b[1]), .B(n27175), .Z(n27177) );
  IV U27848 ( .A(a[194]), .Z(n31644) );
  NANDN U27849 ( .A(n31644), .B(n1049), .Z(n27176) );
  NAND U27850 ( .A(n27177), .B(n27176), .Z(n27247) );
  ANDN U27851 ( .B(b[31]), .A(n27178), .Z(n27244) );
  NANDN U27852 ( .A(n27179), .B(n38490), .Z(n27181) );
  XNOR U27853 ( .A(n1058), .B(a[167]), .Z(n27316) );
  NANDN U27854 ( .A(n1048), .B(n27316), .Z(n27180) );
  NAND U27855 ( .A(n27181), .B(n27180), .Z(n27245) );
  XOR U27856 ( .A(n27244), .B(n27245), .Z(n27246) );
  XNOR U27857 ( .A(n27247), .B(n27246), .Z(n27220) );
  NANDN U27858 ( .A(n27182), .B(n38205), .Z(n27184) );
  XNOR U27859 ( .A(b[23]), .B(a[173]), .Z(n27319) );
  OR U27860 ( .A(n27319), .B(n38268), .Z(n27183) );
  NAND U27861 ( .A(n27184), .B(n27183), .Z(n27289) );
  XNOR U27862 ( .A(b[7]), .B(a[189]), .Z(n27322) );
  NANDN U27863 ( .A(n27322), .B(n36701), .Z(n27187) );
  NAND U27864 ( .A(n27185), .B(n36702), .Z(n27186) );
  NAND U27865 ( .A(n27187), .B(n27186), .Z(n27286) );
  XOR U27866 ( .A(b[25]), .B(a[171]), .Z(n27325) );
  NAND U27867 ( .A(n27325), .B(n38325), .Z(n27190) );
  NAND U27868 ( .A(n27188), .B(n38326), .Z(n27189) );
  AND U27869 ( .A(n27190), .B(n27189), .Z(n27287) );
  XNOR U27870 ( .A(n27286), .B(n27287), .Z(n27288) );
  XNOR U27871 ( .A(n27289), .B(n27288), .Z(n27221) );
  XNOR U27872 ( .A(n27220), .B(n27221), .Z(n27222) );
  XOR U27873 ( .A(n27223), .B(n27222), .Z(n27277) );
  XNOR U27874 ( .A(n27276), .B(n27277), .Z(n27334) );
  XNOR U27875 ( .A(n27335), .B(n27334), .Z(n27337) );
  XNOR U27876 ( .A(n27336), .B(n27337), .Z(n27346) );
  XOR U27877 ( .A(n27347), .B(n27346), .Z(n27349) );
  NAND U27878 ( .A(n27192), .B(n27191), .Z(n27196) );
  NAND U27879 ( .A(n27194), .B(n27193), .Z(n27195) );
  NAND U27880 ( .A(n27196), .B(n27195), .Z(n27341) );
  NAND U27881 ( .A(n27198), .B(n27197), .Z(n27202) );
  NANDN U27882 ( .A(n27200), .B(n27199), .Z(n27201) );
  AND U27883 ( .A(n27202), .B(n27201), .Z(n27340) );
  XNOR U27884 ( .A(n27341), .B(n27340), .Z(n27342) );
  XOR U27885 ( .A(n27343), .B(n27342), .Z(n27217) );
  XOR U27886 ( .A(n27216), .B(n27217), .Z(n27208) );
  XOR U27887 ( .A(n27209), .B(n27208), .Z(n27210) );
  XNOR U27888 ( .A(n27211), .B(n27210), .Z(n27352) );
  XNOR U27889 ( .A(n27352), .B(sreg[419]), .Z(n27354) );
  NAND U27890 ( .A(n27203), .B(sreg[418]), .Z(n27207) );
  OR U27891 ( .A(n27205), .B(n27204), .Z(n27206) );
  AND U27892 ( .A(n27207), .B(n27206), .Z(n27353) );
  XOR U27893 ( .A(n27354), .B(n27353), .Z(c[419]) );
  NAND U27894 ( .A(n27209), .B(n27208), .Z(n27213) );
  NAND U27895 ( .A(n27211), .B(n27210), .Z(n27212) );
  NAND U27896 ( .A(n27213), .B(n27212), .Z(n27360) );
  NANDN U27897 ( .A(n27215), .B(n27214), .Z(n27219) );
  NAND U27898 ( .A(n27217), .B(n27216), .Z(n27218) );
  NAND U27899 ( .A(n27219), .B(n27218), .Z(n27358) );
  NANDN U27900 ( .A(n27221), .B(n27220), .Z(n27225) );
  NANDN U27901 ( .A(n27223), .B(n27222), .Z(n27224) );
  NAND U27902 ( .A(n27225), .B(n27224), .Z(n27478) );
  OR U27903 ( .A(n27227), .B(n27226), .Z(n27231) );
  NAND U27904 ( .A(n27229), .B(n27228), .Z(n27230) );
  NAND U27905 ( .A(n27231), .B(n27230), .Z(n27417) );
  OR U27906 ( .A(n27233), .B(n27232), .Z(n27237) );
  NANDN U27907 ( .A(n27235), .B(n27234), .Z(n27236) );
  NAND U27908 ( .A(n27237), .B(n27236), .Z(n27416) );
  OR U27909 ( .A(n27239), .B(n27238), .Z(n27243) );
  NANDN U27910 ( .A(n27241), .B(n27240), .Z(n27242) );
  NAND U27911 ( .A(n27243), .B(n27242), .Z(n27415) );
  XOR U27912 ( .A(n27417), .B(n27418), .Z(n27476) );
  OR U27913 ( .A(n27245), .B(n27244), .Z(n27249) );
  NAND U27914 ( .A(n27247), .B(n27246), .Z(n27248) );
  NAND U27915 ( .A(n27249), .B(n27248), .Z(n27429) );
  XNOR U27916 ( .A(b[19]), .B(a[178]), .Z(n27373) );
  NANDN U27917 ( .A(n27373), .B(n37934), .Z(n27252) );
  NANDN U27918 ( .A(n27250), .B(n37935), .Z(n27251) );
  NAND U27919 ( .A(n27252), .B(n27251), .Z(n27442) );
  XOR U27920 ( .A(b[27]), .B(a[170]), .Z(n27376) );
  NAND U27921 ( .A(n38423), .B(n27376), .Z(n27255) );
  NAND U27922 ( .A(n27253), .B(n38424), .Z(n27254) );
  NAND U27923 ( .A(n27255), .B(n27254), .Z(n27439) );
  XNOR U27924 ( .A(b[5]), .B(a[192]), .Z(n27379) );
  NANDN U27925 ( .A(n27379), .B(n36587), .Z(n27258) );
  NANDN U27926 ( .A(n27256), .B(n36588), .Z(n27257) );
  AND U27927 ( .A(n27258), .B(n27257), .Z(n27440) );
  XNOR U27928 ( .A(n27439), .B(n27440), .Z(n27441) );
  XNOR U27929 ( .A(n27442), .B(n27441), .Z(n27428) );
  NAND U27930 ( .A(n27259), .B(n37762), .Z(n27261) );
  XOR U27931 ( .A(b[17]), .B(a[180]), .Z(n27382) );
  NAND U27932 ( .A(n27382), .B(n37764), .Z(n27260) );
  NAND U27933 ( .A(n27261), .B(n27260), .Z(n27400) );
  XNOR U27934 ( .A(b[31]), .B(a[166]), .Z(n27385) );
  NANDN U27935 ( .A(n27385), .B(n38552), .Z(n27264) );
  NANDN U27936 ( .A(n27262), .B(n38553), .Z(n27263) );
  NAND U27937 ( .A(n27264), .B(n27263), .Z(n27397) );
  OR U27938 ( .A(n27265), .B(n36105), .Z(n27267) );
  XOR U27939 ( .A(b[3]), .B(n31644), .Z(n27388) );
  NANDN U27940 ( .A(n27388), .B(n36107), .Z(n27266) );
  AND U27941 ( .A(n27267), .B(n27266), .Z(n27398) );
  XNOR U27942 ( .A(n27397), .B(n27398), .Z(n27399) );
  XOR U27943 ( .A(n27400), .B(n27399), .Z(n27427) );
  XOR U27944 ( .A(n27428), .B(n27427), .Z(n27430) );
  XOR U27945 ( .A(n27429), .B(n27430), .Z(n27475) );
  XOR U27946 ( .A(n27476), .B(n27475), .Z(n27477) );
  XNOR U27947 ( .A(n27478), .B(n27477), .Z(n27496) );
  OR U27948 ( .A(n27269), .B(n27268), .Z(n27273) );
  NAND U27949 ( .A(n27271), .B(n27270), .Z(n27272) );
  NAND U27950 ( .A(n27273), .B(n27272), .Z(n27494) );
  NANDN U27951 ( .A(n27275), .B(n27274), .Z(n27279) );
  NANDN U27952 ( .A(n27277), .B(n27276), .Z(n27278) );
  NAND U27953 ( .A(n27279), .B(n27278), .Z(n27483) );
  OR U27954 ( .A(n27281), .B(n27280), .Z(n27285) );
  NAND U27955 ( .A(n27283), .B(n27282), .Z(n27284) );
  NAND U27956 ( .A(n27285), .B(n27284), .Z(n27482) );
  NANDN U27957 ( .A(n27287), .B(n27286), .Z(n27291) );
  NAND U27958 ( .A(n27289), .B(n27288), .Z(n27290) );
  NAND U27959 ( .A(n27291), .B(n27290), .Z(n27421) );
  NANDN U27960 ( .A(n27293), .B(n27292), .Z(n27297) );
  NAND U27961 ( .A(n27295), .B(n27294), .Z(n27296) );
  AND U27962 ( .A(n27297), .B(n27296), .Z(n27422) );
  XNOR U27963 ( .A(n27421), .B(n27422), .Z(n27423) );
  XNOR U27964 ( .A(b[9]), .B(a[188]), .Z(n27445) );
  NANDN U27965 ( .A(n27445), .B(n36925), .Z(n27300) );
  NANDN U27966 ( .A(n27298), .B(n36926), .Z(n27299) );
  NAND U27967 ( .A(n27300), .B(n27299), .Z(n27405) );
  XNOR U27968 ( .A(b[15]), .B(a[182]), .Z(n27448) );
  OR U27969 ( .A(n27448), .B(n37665), .Z(n27303) );
  NANDN U27970 ( .A(n27301), .B(n37604), .Z(n27302) );
  AND U27971 ( .A(n27303), .B(n27302), .Z(n27403) );
  XNOR U27972 ( .A(b[21]), .B(a[176]), .Z(n27451) );
  NANDN U27973 ( .A(n27451), .B(n38101), .Z(n27306) );
  NANDN U27974 ( .A(n27304), .B(n38102), .Z(n27305) );
  AND U27975 ( .A(n27306), .B(n27305), .Z(n27404) );
  XOR U27976 ( .A(n27405), .B(n27406), .Z(n27394) );
  XNOR U27977 ( .A(b[11]), .B(a[186]), .Z(n27454) );
  OR U27978 ( .A(n27454), .B(n37311), .Z(n27309) );
  NANDN U27979 ( .A(n27307), .B(n37218), .Z(n27308) );
  NAND U27980 ( .A(n27309), .B(n27308), .Z(n27392) );
  XOR U27981 ( .A(n1053), .B(a[184]), .Z(n27457) );
  NANDN U27982 ( .A(n27457), .B(n37424), .Z(n27312) );
  NANDN U27983 ( .A(n27310), .B(n37425), .Z(n27311) );
  AND U27984 ( .A(n27312), .B(n27311), .Z(n27391) );
  XNOR U27985 ( .A(n27392), .B(n27391), .Z(n27393) );
  XOR U27986 ( .A(n27394), .B(n27393), .Z(n27411) );
  NANDN U27987 ( .A(n1049), .B(a[196]), .Z(n27313) );
  XNOR U27988 ( .A(b[1]), .B(n27313), .Z(n27315) );
  IV U27989 ( .A(a[195]), .Z(n31434) );
  NANDN U27990 ( .A(n31434), .B(n1049), .Z(n27314) );
  AND U27991 ( .A(n27315), .B(n27314), .Z(n27369) );
  NAND U27992 ( .A(n27316), .B(n38490), .Z(n27318) );
  XNOR U27993 ( .A(n1058), .B(a[168]), .Z(n27460) );
  NANDN U27994 ( .A(n1048), .B(n27460), .Z(n27317) );
  NAND U27995 ( .A(n27318), .B(n27317), .Z(n27367) );
  NANDN U27996 ( .A(n1059), .B(a[164]), .Z(n27368) );
  XNOR U27997 ( .A(n27367), .B(n27368), .Z(n27370) );
  XOR U27998 ( .A(n27369), .B(n27370), .Z(n27409) );
  NANDN U27999 ( .A(n27319), .B(n38205), .Z(n27321) );
  XNOR U28000 ( .A(b[23]), .B(a[174]), .Z(n27466) );
  OR U28001 ( .A(n27466), .B(n38268), .Z(n27320) );
  NAND U28002 ( .A(n27321), .B(n27320), .Z(n27436) );
  XOR U28003 ( .A(b[7]), .B(a[190]), .Z(n27469) );
  NAND U28004 ( .A(n27469), .B(n36701), .Z(n27324) );
  NANDN U28005 ( .A(n27322), .B(n36702), .Z(n27323) );
  NAND U28006 ( .A(n27324), .B(n27323), .Z(n27433) );
  XOR U28007 ( .A(b[25]), .B(a[172]), .Z(n27472) );
  NAND U28008 ( .A(n27472), .B(n38325), .Z(n27327) );
  NAND U28009 ( .A(n27325), .B(n38326), .Z(n27326) );
  AND U28010 ( .A(n27327), .B(n27326), .Z(n27434) );
  XNOR U28011 ( .A(n27433), .B(n27434), .Z(n27435) );
  XNOR U28012 ( .A(n27436), .B(n27435), .Z(n27410) );
  XOR U28013 ( .A(n27409), .B(n27410), .Z(n27412) );
  XNOR U28014 ( .A(n27411), .B(n27412), .Z(n27424) );
  XNOR U28015 ( .A(n27423), .B(n27424), .Z(n27481) );
  XNOR U28016 ( .A(n27482), .B(n27481), .Z(n27484) );
  XNOR U28017 ( .A(n27483), .B(n27484), .Z(n27493) );
  XNOR U28018 ( .A(n27494), .B(n27493), .Z(n27495) );
  XOR U28019 ( .A(n27496), .B(n27495), .Z(n27490) );
  NANDN U28020 ( .A(n27329), .B(n27328), .Z(n27333) );
  OR U28021 ( .A(n27331), .B(n27330), .Z(n27332) );
  NAND U28022 ( .A(n27333), .B(n27332), .Z(n27487) );
  NAND U28023 ( .A(n27335), .B(n27334), .Z(n27339) );
  NANDN U28024 ( .A(n27337), .B(n27336), .Z(n27338) );
  NAND U28025 ( .A(n27339), .B(n27338), .Z(n27488) );
  XNOR U28026 ( .A(n27487), .B(n27488), .Z(n27489) );
  XNOR U28027 ( .A(n27490), .B(n27489), .Z(n27364) );
  NANDN U28028 ( .A(n27341), .B(n27340), .Z(n27345) );
  NAND U28029 ( .A(n27343), .B(n27342), .Z(n27344) );
  NAND U28030 ( .A(n27345), .B(n27344), .Z(n27361) );
  NANDN U28031 ( .A(n27347), .B(n27346), .Z(n27351) );
  OR U28032 ( .A(n27349), .B(n27348), .Z(n27350) );
  NAND U28033 ( .A(n27351), .B(n27350), .Z(n27362) );
  XNOR U28034 ( .A(n27361), .B(n27362), .Z(n27363) );
  XNOR U28035 ( .A(n27364), .B(n27363), .Z(n27357) );
  XOR U28036 ( .A(n27358), .B(n27357), .Z(n27359) );
  XNOR U28037 ( .A(n27360), .B(n27359), .Z(n27499) );
  XNOR U28038 ( .A(n27499), .B(sreg[420]), .Z(n27501) );
  NAND U28039 ( .A(n27352), .B(sreg[419]), .Z(n27356) );
  OR U28040 ( .A(n27354), .B(n27353), .Z(n27355) );
  AND U28041 ( .A(n27356), .B(n27355), .Z(n27500) );
  XOR U28042 ( .A(n27501), .B(n27500), .Z(c[420]) );
  NANDN U28043 ( .A(n27362), .B(n27361), .Z(n27366) );
  NANDN U28044 ( .A(n27364), .B(n27363), .Z(n27365) );
  NAND U28045 ( .A(n27366), .B(n27365), .Z(n27505) );
  NANDN U28046 ( .A(n27368), .B(n27367), .Z(n27372) );
  NAND U28047 ( .A(n27370), .B(n27369), .Z(n27371) );
  NAND U28048 ( .A(n27372), .B(n27371), .Z(n27591) );
  XNOR U28049 ( .A(b[19]), .B(a[179]), .Z(n27534) );
  NANDN U28050 ( .A(n27534), .B(n37934), .Z(n27375) );
  NANDN U28051 ( .A(n27373), .B(n37935), .Z(n27374) );
  NAND U28052 ( .A(n27375), .B(n27374), .Z(n27625) );
  XOR U28053 ( .A(b[27]), .B(a[171]), .Z(n27537) );
  NAND U28054 ( .A(n38423), .B(n27537), .Z(n27378) );
  NAND U28055 ( .A(n27376), .B(n38424), .Z(n27377) );
  NAND U28056 ( .A(n27378), .B(n27377), .Z(n27622) );
  XOR U28057 ( .A(b[5]), .B(n31508), .Z(n27540) );
  NANDN U28058 ( .A(n27540), .B(n36587), .Z(n27381) );
  NANDN U28059 ( .A(n27379), .B(n36588), .Z(n27380) );
  AND U28060 ( .A(n27381), .B(n27380), .Z(n27623) );
  XNOR U28061 ( .A(n27622), .B(n27623), .Z(n27624) );
  XNOR U28062 ( .A(n27625), .B(n27624), .Z(n27589) );
  NAND U28063 ( .A(n27382), .B(n37762), .Z(n27384) );
  XOR U28064 ( .A(b[17]), .B(a[181]), .Z(n27543) );
  NAND U28065 ( .A(n27543), .B(n37764), .Z(n27383) );
  NAND U28066 ( .A(n27384), .B(n27383), .Z(n27561) );
  XNOR U28067 ( .A(b[31]), .B(a[167]), .Z(n27546) );
  NANDN U28068 ( .A(n27546), .B(n38552), .Z(n27387) );
  NANDN U28069 ( .A(n27385), .B(n38553), .Z(n27386) );
  NAND U28070 ( .A(n27387), .B(n27386), .Z(n27558) );
  OR U28071 ( .A(n27388), .B(n36105), .Z(n27390) );
  XOR U28072 ( .A(b[3]), .B(n31434), .Z(n27549) );
  NANDN U28073 ( .A(n27549), .B(n36107), .Z(n27389) );
  AND U28074 ( .A(n27390), .B(n27389), .Z(n27559) );
  XNOR U28075 ( .A(n27558), .B(n27559), .Z(n27560) );
  XOR U28076 ( .A(n27561), .B(n27560), .Z(n27588) );
  XNOR U28077 ( .A(n27589), .B(n27588), .Z(n27590) );
  XNOR U28078 ( .A(n27591), .B(n27590), .Z(n27634) );
  NANDN U28079 ( .A(n27392), .B(n27391), .Z(n27396) );
  NAND U28080 ( .A(n27394), .B(n27393), .Z(n27395) );
  NAND U28081 ( .A(n27396), .B(n27395), .Z(n27579) );
  NANDN U28082 ( .A(n27398), .B(n27397), .Z(n27402) );
  NAND U28083 ( .A(n27400), .B(n27399), .Z(n27401) );
  NAND U28084 ( .A(n27402), .B(n27401), .Z(n27577) );
  OR U28085 ( .A(n27404), .B(n27403), .Z(n27408) );
  NANDN U28086 ( .A(n27406), .B(n27405), .Z(n27407) );
  NAND U28087 ( .A(n27408), .B(n27407), .Z(n27576) );
  XNOR U28088 ( .A(n27579), .B(n27578), .Z(n27635) );
  XOR U28089 ( .A(n27634), .B(n27635), .Z(n27637) );
  NANDN U28090 ( .A(n27410), .B(n27409), .Z(n27414) );
  OR U28091 ( .A(n27412), .B(n27411), .Z(n27413) );
  NAND U28092 ( .A(n27414), .B(n27413), .Z(n27636) );
  XOR U28093 ( .A(n27637), .B(n27636), .Z(n27524) );
  OR U28094 ( .A(n27416), .B(n27415), .Z(n27420) );
  NANDN U28095 ( .A(n27418), .B(n27417), .Z(n27419) );
  NAND U28096 ( .A(n27420), .B(n27419), .Z(n27523) );
  NANDN U28097 ( .A(n27422), .B(n27421), .Z(n27426) );
  NANDN U28098 ( .A(n27424), .B(n27423), .Z(n27425) );
  NAND U28099 ( .A(n27426), .B(n27425), .Z(n27642) );
  NANDN U28100 ( .A(n27428), .B(n27427), .Z(n27432) );
  OR U28101 ( .A(n27430), .B(n27429), .Z(n27431) );
  NAND U28102 ( .A(n27432), .B(n27431), .Z(n27641) );
  NANDN U28103 ( .A(n27434), .B(n27433), .Z(n27438) );
  NAND U28104 ( .A(n27436), .B(n27435), .Z(n27437) );
  NAND U28105 ( .A(n27438), .B(n27437), .Z(n27582) );
  NANDN U28106 ( .A(n27440), .B(n27439), .Z(n27444) );
  NAND U28107 ( .A(n27442), .B(n27441), .Z(n27443) );
  AND U28108 ( .A(n27444), .B(n27443), .Z(n27583) );
  XNOR U28109 ( .A(n27582), .B(n27583), .Z(n27584) );
  XOR U28110 ( .A(b[9]), .B(n30936), .Z(n27592) );
  NANDN U28111 ( .A(n27592), .B(n36925), .Z(n27447) );
  NANDN U28112 ( .A(n27445), .B(n36926), .Z(n27446) );
  NAND U28113 ( .A(n27447), .B(n27446), .Z(n27566) );
  XNOR U28114 ( .A(b[15]), .B(a[183]), .Z(n27595) );
  OR U28115 ( .A(n27595), .B(n37665), .Z(n27450) );
  NANDN U28116 ( .A(n27448), .B(n37604), .Z(n27449) );
  AND U28117 ( .A(n27450), .B(n27449), .Z(n27564) );
  XNOR U28118 ( .A(b[21]), .B(a[177]), .Z(n27598) );
  NANDN U28119 ( .A(n27598), .B(n38101), .Z(n27453) );
  NANDN U28120 ( .A(n27451), .B(n38102), .Z(n27452) );
  AND U28121 ( .A(n27453), .B(n27452), .Z(n27565) );
  XOR U28122 ( .A(n27566), .B(n27567), .Z(n27555) );
  XNOR U28123 ( .A(b[11]), .B(a[187]), .Z(n27601) );
  OR U28124 ( .A(n27601), .B(n37311), .Z(n27456) );
  NANDN U28125 ( .A(n27454), .B(n37218), .Z(n27455) );
  NAND U28126 ( .A(n27456), .B(n27455), .Z(n27553) );
  XOR U28127 ( .A(n1053), .B(a[185]), .Z(n27604) );
  NANDN U28128 ( .A(n27604), .B(n37424), .Z(n27459) );
  NANDN U28129 ( .A(n27457), .B(n37425), .Z(n27458) );
  AND U28130 ( .A(n27459), .B(n27458), .Z(n27552) );
  XNOR U28131 ( .A(n27553), .B(n27552), .Z(n27554) );
  XOR U28132 ( .A(n27555), .B(n27554), .Z(n27572) );
  NAND U28133 ( .A(n38490), .B(n27460), .Z(n27462) );
  XNOR U28134 ( .A(n1058), .B(a[169]), .Z(n27610) );
  NANDN U28135 ( .A(n1048), .B(n27610), .Z(n27461) );
  NAND U28136 ( .A(n27462), .B(n27461), .Z(n27528) );
  NANDN U28137 ( .A(n1059), .B(a[165]), .Z(n27529) );
  XNOR U28138 ( .A(n27528), .B(n27529), .Z(n27531) );
  NANDN U28139 ( .A(n1049), .B(a[197]), .Z(n27463) );
  XNOR U28140 ( .A(b[1]), .B(n27463), .Z(n27465) );
  NANDN U28141 ( .A(b[0]), .B(a[196]), .Z(n27464) );
  AND U28142 ( .A(n27465), .B(n27464), .Z(n27530) );
  XOR U28143 ( .A(n27531), .B(n27530), .Z(n27570) );
  NANDN U28144 ( .A(n27466), .B(n38205), .Z(n27468) );
  XNOR U28145 ( .A(b[23]), .B(a[175]), .Z(n27613) );
  OR U28146 ( .A(n27613), .B(n38268), .Z(n27467) );
  NAND U28147 ( .A(n27468), .B(n27467), .Z(n27631) );
  XOR U28148 ( .A(b[7]), .B(a[191]), .Z(n27616) );
  NAND U28149 ( .A(n27616), .B(n36701), .Z(n27471) );
  NAND U28150 ( .A(n27469), .B(n36702), .Z(n27470) );
  NAND U28151 ( .A(n27471), .B(n27470), .Z(n27628) );
  XOR U28152 ( .A(b[25]), .B(a[173]), .Z(n27619) );
  NAND U28153 ( .A(n27619), .B(n38325), .Z(n27474) );
  NAND U28154 ( .A(n27472), .B(n38326), .Z(n27473) );
  AND U28155 ( .A(n27474), .B(n27473), .Z(n27629) );
  XNOR U28156 ( .A(n27628), .B(n27629), .Z(n27630) );
  XNOR U28157 ( .A(n27631), .B(n27630), .Z(n27571) );
  XOR U28158 ( .A(n27570), .B(n27571), .Z(n27573) );
  XNOR U28159 ( .A(n27572), .B(n27573), .Z(n27585) );
  XNOR U28160 ( .A(n27584), .B(n27585), .Z(n27640) );
  XNOR U28161 ( .A(n27641), .B(n27640), .Z(n27643) );
  XNOR U28162 ( .A(n27642), .B(n27643), .Z(n27522) );
  XOR U28163 ( .A(n27523), .B(n27522), .Z(n27525) );
  NAND U28164 ( .A(n27476), .B(n27475), .Z(n27480) );
  NAND U28165 ( .A(n27478), .B(n27477), .Z(n27479) );
  NAND U28166 ( .A(n27480), .B(n27479), .Z(n27517) );
  NAND U28167 ( .A(n27482), .B(n27481), .Z(n27486) );
  NANDN U28168 ( .A(n27484), .B(n27483), .Z(n27485) );
  AND U28169 ( .A(n27486), .B(n27485), .Z(n27516) );
  XNOR U28170 ( .A(n27517), .B(n27516), .Z(n27518) );
  XOR U28171 ( .A(n27519), .B(n27518), .Z(n27512) );
  NANDN U28172 ( .A(n27488), .B(n27487), .Z(n27492) );
  NAND U28173 ( .A(n27490), .B(n27489), .Z(n27491) );
  NAND U28174 ( .A(n27492), .B(n27491), .Z(n27510) );
  NANDN U28175 ( .A(n27494), .B(n27493), .Z(n27498) );
  NANDN U28176 ( .A(n27496), .B(n27495), .Z(n27497) );
  NAND U28177 ( .A(n27498), .B(n27497), .Z(n27511) );
  XNOR U28178 ( .A(n27510), .B(n27511), .Z(n27513) );
  XOR U28179 ( .A(n27512), .B(n27513), .Z(n27504) );
  XOR U28180 ( .A(n27505), .B(n27504), .Z(n27506) );
  XNOR U28181 ( .A(n27507), .B(n27506), .Z(n27646) );
  XNOR U28182 ( .A(n27646), .B(sreg[421]), .Z(n27648) );
  NAND U28183 ( .A(n27499), .B(sreg[420]), .Z(n27503) );
  OR U28184 ( .A(n27501), .B(n27500), .Z(n27502) );
  AND U28185 ( .A(n27503), .B(n27502), .Z(n27647) );
  XOR U28186 ( .A(n27648), .B(n27647), .Z(c[421]) );
  NAND U28187 ( .A(n27505), .B(n27504), .Z(n27509) );
  NAND U28188 ( .A(n27507), .B(n27506), .Z(n27508) );
  NAND U28189 ( .A(n27509), .B(n27508), .Z(n27654) );
  NANDN U28190 ( .A(n27511), .B(n27510), .Z(n27515) );
  NAND U28191 ( .A(n27513), .B(n27512), .Z(n27514) );
  NAND U28192 ( .A(n27515), .B(n27514), .Z(n27652) );
  NANDN U28193 ( .A(n27517), .B(n27516), .Z(n27521) );
  NAND U28194 ( .A(n27519), .B(n27518), .Z(n27520) );
  NAND U28195 ( .A(n27521), .B(n27520), .Z(n27657) );
  NANDN U28196 ( .A(n27523), .B(n27522), .Z(n27527) );
  OR U28197 ( .A(n27525), .B(n27524), .Z(n27526) );
  NAND U28198 ( .A(n27527), .B(n27526), .Z(n27658) );
  XNOR U28199 ( .A(n27657), .B(n27658), .Z(n27659) );
  NANDN U28200 ( .A(n27529), .B(n27528), .Z(n27533) );
  NAND U28201 ( .A(n27531), .B(n27530), .Z(n27532) );
  NAND U28202 ( .A(n27533), .B(n27532), .Z(n27726) );
  XNOR U28203 ( .A(b[19]), .B(a[180]), .Z(n27693) );
  NANDN U28204 ( .A(n27693), .B(n37934), .Z(n27536) );
  NANDN U28205 ( .A(n27534), .B(n37935), .Z(n27535) );
  NAND U28206 ( .A(n27536), .B(n27535), .Z(n27738) );
  XOR U28207 ( .A(b[27]), .B(a[172]), .Z(n27696) );
  NAND U28208 ( .A(n38423), .B(n27696), .Z(n27539) );
  NAND U28209 ( .A(n27537), .B(n38424), .Z(n27538) );
  NAND U28210 ( .A(n27539), .B(n27538), .Z(n27735) );
  XOR U28211 ( .A(b[5]), .B(n31644), .Z(n27699) );
  NANDN U28212 ( .A(n27699), .B(n36587), .Z(n27542) );
  NANDN U28213 ( .A(n27540), .B(n36588), .Z(n27541) );
  AND U28214 ( .A(n27542), .B(n27541), .Z(n27736) );
  XNOR U28215 ( .A(n27735), .B(n27736), .Z(n27737) );
  XNOR U28216 ( .A(n27738), .B(n27737), .Z(n27723) );
  NAND U28217 ( .A(n27543), .B(n37762), .Z(n27545) );
  XOR U28218 ( .A(b[17]), .B(a[182]), .Z(n27702) );
  NAND U28219 ( .A(n27702), .B(n37764), .Z(n27544) );
  NAND U28220 ( .A(n27545), .B(n27544), .Z(n27677) );
  XNOR U28221 ( .A(b[31]), .B(a[168]), .Z(n27705) );
  NANDN U28222 ( .A(n27705), .B(n38552), .Z(n27548) );
  NANDN U28223 ( .A(n27546), .B(n38553), .Z(n27547) );
  AND U28224 ( .A(n27548), .B(n27547), .Z(n27675) );
  OR U28225 ( .A(n27549), .B(n36105), .Z(n27551) );
  XNOR U28226 ( .A(b[3]), .B(a[196]), .Z(n27708) );
  NANDN U28227 ( .A(n27708), .B(n36107), .Z(n27550) );
  AND U28228 ( .A(n27551), .B(n27550), .Z(n27676) );
  XOR U28229 ( .A(n27677), .B(n27678), .Z(n27724) );
  XOR U28230 ( .A(n27723), .B(n27724), .Z(n27725) );
  XNOR U28231 ( .A(n27726), .B(n27725), .Z(n27771) );
  NANDN U28232 ( .A(n27553), .B(n27552), .Z(n27557) );
  NAND U28233 ( .A(n27555), .B(n27554), .Z(n27556) );
  NAND U28234 ( .A(n27557), .B(n27556), .Z(n27714) );
  NANDN U28235 ( .A(n27559), .B(n27558), .Z(n27563) );
  NAND U28236 ( .A(n27561), .B(n27560), .Z(n27562) );
  NAND U28237 ( .A(n27563), .B(n27562), .Z(n27712) );
  OR U28238 ( .A(n27565), .B(n27564), .Z(n27569) );
  NANDN U28239 ( .A(n27567), .B(n27566), .Z(n27568) );
  NAND U28240 ( .A(n27569), .B(n27568), .Z(n27711) );
  XNOR U28241 ( .A(n27714), .B(n27713), .Z(n27772) );
  XOR U28242 ( .A(n27771), .B(n27772), .Z(n27774) );
  NANDN U28243 ( .A(n27571), .B(n27570), .Z(n27575) );
  OR U28244 ( .A(n27573), .B(n27572), .Z(n27574) );
  NAND U28245 ( .A(n27575), .B(n27574), .Z(n27773) );
  XOR U28246 ( .A(n27774), .B(n27773), .Z(n27791) );
  OR U28247 ( .A(n27577), .B(n27576), .Z(n27581) );
  NAND U28248 ( .A(n27579), .B(n27578), .Z(n27580) );
  NAND U28249 ( .A(n27581), .B(n27580), .Z(n27790) );
  NANDN U28250 ( .A(n27583), .B(n27582), .Z(n27587) );
  NANDN U28251 ( .A(n27585), .B(n27584), .Z(n27586) );
  NAND U28252 ( .A(n27587), .B(n27586), .Z(n27780) );
  XNOR U28253 ( .A(n1052), .B(a[190]), .Z(n27741) );
  NAND U28254 ( .A(n36925), .B(n27741), .Z(n27594) );
  NANDN U28255 ( .A(n27592), .B(n36926), .Z(n27593) );
  NAND U28256 ( .A(n27594), .B(n27593), .Z(n27683) );
  XNOR U28257 ( .A(b[15]), .B(a[184]), .Z(n27744) );
  OR U28258 ( .A(n27744), .B(n37665), .Z(n27597) );
  NANDN U28259 ( .A(n27595), .B(n37604), .Z(n27596) );
  AND U28260 ( .A(n27597), .B(n27596), .Z(n27681) );
  XNOR U28261 ( .A(n1056), .B(a[178]), .Z(n27747) );
  NAND U28262 ( .A(n27747), .B(n38101), .Z(n27600) );
  NANDN U28263 ( .A(n27598), .B(n38102), .Z(n27599) );
  AND U28264 ( .A(n27600), .B(n27599), .Z(n27682) );
  XOR U28265 ( .A(n27683), .B(n27684), .Z(n27672) );
  XNOR U28266 ( .A(b[11]), .B(a[188]), .Z(n27750) );
  OR U28267 ( .A(n27750), .B(n37311), .Z(n27603) );
  NANDN U28268 ( .A(n27601), .B(n37218), .Z(n27602) );
  NAND U28269 ( .A(n27603), .B(n27602), .Z(n27670) );
  XOR U28270 ( .A(n1053), .B(a[186]), .Z(n27753) );
  NANDN U28271 ( .A(n27753), .B(n37424), .Z(n27606) );
  NANDN U28272 ( .A(n27604), .B(n37425), .Z(n27605) );
  NAND U28273 ( .A(n27606), .B(n27605), .Z(n27669) );
  XOR U28274 ( .A(n27672), .B(n27671), .Z(n27666) );
  NANDN U28275 ( .A(n1049), .B(a[198]), .Z(n27607) );
  XNOR U28276 ( .A(b[1]), .B(n27607), .Z(n27609) );
  NANDN U28277 ( .A(b[0]), .B(a[197]), .Z(n27608) );
  AND U28278 ( .A(n27609), .B(n27608), .Z(n27689) );
  NAND U28279 ( .A(n38490), .B(n27610), .Z(n27612) );
  XNOR U28280 ( .A(n1058), .B(a[170]), .Z(n27759) );
  NANDN U28281 ( .A(n1048), .B(n27759), .Z(n27611) );
  NAND U28282 ( .A(n27612), .B(n27611), .Z(n27687) );
  NANDN U28283 ( .A(n1059), .B(a[166]), .Z(n27688) );
  XNOR U28284 ( .A(n27687), .B(n27688), .Z(n27690) );
  XNOR U28285 ( .A(n27689), .B(n27690), .Z(n27664) );
  NANDN U28286 ( .A(n27613), .B(n38205), .Z(n27615) );
  XNOR U28287 ( .A(b[23]), .B(a[176]), .Z(n27762) );
  OR U28288 ( .A(n27762), .B(n38268), .Z(n27614) );
  NAND U28289 ( .A(n27615), .B(n27614), .Z(n27732) );
  XOR U28290 ( .A(b[7]), .B(a[192]), .Z(n27765) );
  NAND U28291 ( .A(n27765), .B(n36701), .Z(n27618) );
  NAND U28292 ( .A(n27616), .B(n36702), .Z(n27617) );
  NAND U28293 ( .A(n27618), .B(n27617), .Z(n27729) );
  XOR U28294 ( .A(b[25]), .B(a[174]), .Z(n27768) );
  NAND U28295 ( .A(n27768), .B(n38325), .Z(n27621) );
  NAND U28296 ( .A(n27619), .B(n38326), .Z(n27620) );
  AND U28297 ( .A(n27621), .B(n27620), .Z(n27730) );
  XNOR U28298 ( .A(n27729), .B(n27730), .Z(n27731) );
  XOR U28299 ( .A(n27732), .B(n27731), .Z(n27663) );
  XNOR U28300 ( .A(n27666), .B(n27665), .Z(n27720) );
  NANDN U28301 ( .A(n27623), .B(n27622), .Z(n27627) );
  NAND U28302 ( .A(n27625), .B(n27624), .Z(n27626) );
  NAND U28303 ( .A(n27627), .B(n27626), .Z(n27718) );
  NANDN U28304 ( .A(n27629), .B(n27628), .Z(n27633) );
  NAND U28305 ( .A(n27631), .B(n27630), .Z(n27632) );
  AND U28306 ( .A(n27633), .B(n27632), .Z(n27717) );
  XNOR U28307 ( .A(n27718), .B(n27717), .Z(n27719) );
  XNOR U28308 ( .A(n27720), .B(n27719), .Z(n27778) );
  XNOR U28309 ( .A(n27777), .B(n27778), .Z(n27779) );
  XOR U28310 ( .A(n27780), .B(n27779), .Z(n27789) );
  XOR U28311 ( .A(n27790), .B(n27789), .Z(n27792) );
  NANDN U28312 ( .A(n27635), .B(n27634), .Z(n27639) );
  OR U28313 ( .A(n27637), .B(n27636), .Z(n27638) );
  NAND U28314 ( .A(n27639), .B(n27638), .Z(n27783) );
  NAND U28315 ( .A(n27641), .B(n27640), .Z(n27645) );
  NANDN U28316 ( .A(n27643), .B(n27642), .Z(n27644) );
  NAND U28317 ( .A(n27645), .B(n27644), .Z(n27784) );
  XNOR U28318 ( .A(n27783), .B(n27784), .Z(n27785) );
  XOR U28319 ( .A(n27786), .B(n27785), .Z(n27660) );
  XOR U28320 ( .A(n27659), .B(n27660), .Z(n27651) );
  XOR U28321 ( .A(n27652), .B(n27651), .Z(n27653) );
  XNOR U28322 ( .A(n27654), .B(n27653), .Z(n27795) );
  XNOR U28323 ( .A(n27795), .B(sreg[422]), .Z(n27797) );
  NAND U28324 ( .A(n27646), .B(sreg[421]), .Z(n27650) );
  OR U28325 ( .A(n27648), .B(n27647), .Z(n27649) );
  AND U28326 ( .A(n27650), .B(n27649), .Z(n27796) );
  XOR U28327 ( .A(n27797), .B(n27796), .Z(c[422]) );
  NAND U28328 ( .A(n27652), .B(n27651), .Z(n27656) );
  NAND U28329 ( .A(n27654), .B(n27653), .Z(n27655) );
  NAND U28330 ( .A(n27656), .B(n27655), .Z(n27803) );
  NANDN U28331 ( .A(n27658), .B(n27657), .Z(n27662) );
  NAND U28332 ( .A(n27660), .B(n27659), .Z(n27661) );
  NAND U28333 ( .A(n27662), .B(n27661), .Z(n27801) );
  NANDN U28334 ( .A(n27664), .B(n27663), .Z(n27668) );
  NANDN U28335 ( .A(n27666), .B(n27665), .Z(n27667) );
  NAND U28336 ( .A(n27668), .B(n27667), .Z(n27919) );
  OR U28337 ( .A(n27670), .B(n27669), .Z(n27674) );
  NAND U28338 ( .A(n27672), .B(n27671), .Z(n27673) );
  NAND U28339 ( .A(n27674), .B(n27673), .Z(n27858) );
  OR U28340 ( .A(n27676), .B(n27675), .Z(n27680) );
  NANDN U28341 ( .A(n27678), .B(n27677), .Z(n27679) );
  NAND U28342 ( .A(n27680), .B(n27679), .Z(n27857) );
  OR U28343 ( .A(n27682), .B(n27681), .Z(n27686) );
  NANDN U28344 ( .A(n27684), .B(n27683), .Z(n27685) );
  NAND U28345 ( .A(n27686), .B(n27685), .Z(n27856) );
  XOR U28346 ( .A(n27858), .B(n27859), .Z(n27916) );
  NANDN U28347 ( .A(n27688), .B(n27687), .Z(n27692) );
  NAND U28348 ( .A(n27690), .B(n27689), .Z(n27691) );
  NAND U28349 ( .A(n27692), .B(n27691), .Z(n27871) );
  XNOR U28350 ( .A(b[19]), .B(a[181]), .Z(n27816) );
  NANDN U28351 ( .A(n27816), .B(n37934), .Z(n27695) );
  NANDN U28352 ( .A(n27693), .B(n37935), .Z(n27694) );
  NAND U28353 ( .A(n27695), .B(n27694), .Z(n27883) );
  XOR U28354 ( .A(b[27]), .B(a[173]), .Z(n27819) );
  NAND U28355 ( .A(n38423), .B(n27819), .Z(n27698) );
  NAND U28356 ( .A(n27696), .B(n38424), .Z(n27697) );
  NAND U28357 ( .A(n27698), .B(n27697), .Z(n27880) );
  XOR U28358 ( .A(b[5]), .B(n31434), .Z(n27822) );
  NANDN U28359 ( .A(n27822), .B(n36587), .Z(n27701) );
  NANDN U28360 ( .A(n27699), .B(n36588), .Z(n27700) );
  AND U28361 ( .A(n27701), .B(n27700), .Z(n27881) );
  XNOR U28362 ( .A(n27880), .B(n27881), .Z(n27882) );
  XNOR U28363 ( .A(n27883), .B(n27882), .Z(n27869) );
  NAND U28364 ( .A(n27702), .B(n37762), .Z(n27704) );
  XOR U28365 ( .A(b[17]), .B(a[183]), .Z(n27825) );
  NAND U28366 ( .A(n27825), .B(n37764), .Z(n27703) );
  NAND U28367 ( .A(n27704), .B(n27703), .Z(n27843) );
  XNOR U28368 ( .A(b[31]), .B(a[169]), .Z(n27828) );
  NANDN U28369 ( .A(n27828), .B(n38552), .Z(n27707) );
  NANDN U28370 ( .A(n27705), .B(n38553), .Z(n27706) );
  NAND U28371 ( .A(n27707), .B(n27706), .Z(n27840) );
  OR U28372 ( .A(n27708), .B(n36105), .Z(n27710) );
  XNOR U28373 ( .A(b[3]), .B(a[197]), .Z(n27831) );
  NANDN U28374 ( .A(n27831), .B(n36107), .Z(n27709) );
  AND U28375 ( .A(n27710), .B(n27709), .Z(n27841) );
  XNOR U28376 ( .A(n27840), .B(n27841), .Z(n27842) );
  XOR U28377 ( .A(n27843), .B(n27842), .Z(n27868) );
  XNOR U28378 ( .A(n27869), .B(n27868), .Z(n27870) );
  XNOR U28379 ( .A(n27871), .B(n27870), .Z(n27917) );
  XNOR U28380 ( .A(n27916), .B(n27917), .Z(n27918) );
  XNOR U28381 ( .A(n27919), .B(n27918), .Z(n27937) );
  OR U28382 ( .A(n27712), .B(n27711), .Z(n27716) );
  NAND U28383 ( .A(n27714), .B(n27713), .Z(n27715) );
  NAND U28384 ( .A(n27716), .B(n27715), .Z(n27935) );
  NANDN U28385 ( .A(n27718), .B(n27717), .Z(n27722) );
  NANDN U28386 ( .A(n27720), .B(n27719), .Z(n27721) );
  NAND U28387 ( .A(n27722), .B(n27721), .Z(n27925) );
  OR U28388 ( .A(n27724), .B(n27723), .Z(n27728) );
  NAND U28389 ( .A(n27726), .B(n27725), .Z(n27727) );
  NAND U28390 ( .A(n27728), .B(n27727), .Z(n27923) );
  NANDN U28391 ( .A(n27730), .B(n27729), .Z(n27734) );
  NAND U28392 ( .A(n27732), .B(n27731), .Z(n27733) );
  NAND U28393 ( .A(n27734), .B(n27733), .Z(n27862) );
  NANDN U28394 ( .A(n27736), .B(n27735), .Z(n27740) );
  NAND U28395 ( .A(n27738), .B(n27737), .Z(n27739) );
  AND U28396 ( .A(n27740), .B(n27739), .Z(n27863) );
  XNOR U28397 ( .A(n27862), .B(n27863), .Z(n27864) );
  XNOR U28398 ( .A(b[9]), .B(a[191]), .Z(n27886) );
  NANDN U28399 ( .A(n27886), .B(n36925), .Z(n27743) );
  NAND U28400 ( .A(n36926), .B(n27741), .Z(n27742) );
  NAND U28401 ( .A(n27743), .B(n27742), .Z(n27848) );
  XNOR U28402 ( .A(n1054), .B(a[185]), .Z(n27889) );
  NANDN U28403 ( .A(n37665), .B(n27889), .Z(n27746) );
  NANDN U28404 ( .A(n27744), .B(n37604), .Z(n27745) );
  NAND U28405 ( .A(n27746), .B(n27745), .Z(n27846) );
  XNOR U28406 ( .A(b[21]), .B(a[179]), .Z(n27892) );
  NANDN U28407 ( .A(n27892), .B(n38101), .Z(n27749) );
  NAND U28408 ( .A(n38102), .B(n27747), .Z(n27748) );
  NAND U28409 ( .A(n27749), .B(n27748), .Z(n27847) );
  XNOR U28410 ( .A(n27846), .B(n27847), .Z(n27849) );
  XOR U28411 ( .A(n27848), .B(n27849), .Z(n27837) );
  XOR U28412 ( .A(b[11]), .B(n30936), .Z(n27895) );
  OR U28413 ( .A(n27895), .B(n37311), .Z(n27752) );
  NANDN U28414 ( .A(n27750), .B(n37218), .Z(n27751) );
  NAND U28415 ( .A(n27752), .B(n27751), .Z(n27835) );
  XOR U28416 ( .A(n1053), .B(a[187]), .Z(n27898) );
  NANDN U28417 ( .A(n27898), .B(n37424), .Z(n27755) );
  NANDN U28418 ( .A(n27753), .B(n37425), .Z(n27754) );
  AND U28419 ( .A(n27755), .B(n27754), .Z(n27834) );
  XNOR U28420 ( .A(n27835), .B(n27834), .Z(n27836) );
  XNOR U28421 ( .A(n27837), .B(n27836), .Z(n27853) );
  NANDN U28422 ( .A(n1049), .B(a[199]), .Z(n27756) );
  XNOR U28423 ( .A(b[1]), .B(n27756), .Z(n27758) );
  IV U28424 ( .A(a[198]), .Z(n32246) );
  NANDN U28425 ( .A(n32246), .B(n1049), .Z(n27757) );
  AND U28426 ( .A(n27758), .B(n27757), .Z(n27812) );
  NAND U28427 ( .A(n38490), .B(n27759), .Z(n27761) );
  XNOR U28428 ( .A(n1058), .B(a[171]), .Z(n27904) );
  NANDN U28429 ( .A(n1048), .B(n27904), .Z(n27760) );
  NAND U28430 ( .A(n27761), .B(n27760), .Z(n27810) );
  NANDN U28431 ( .A(n1059), .B(a[167]), .Z(n27811) );
  XNOR U28432 ( .A(n27810), .B(n27811), .Z(n27813) );
  XNOR U28433 ( .A(n27812), .B(n27813), .Z(n27851) );
  NANDN U28434 ( .A(n27762), .B(n38205), .Z(n27764) );
  XNOR U28435 ( .A(b[23]), .B(a[177]), .Z(n27907) );
  OR U28436 ( .A(n27907), .B(n38268), .Z(n27763) );
  NAND U28437 ( .A(n27764), .B(n27763), .Z(n27877) );
  XNOR U28438 ( .A(b[7]), .B(a[193]), .Z(n27910) );
  NANDN U28439 ( .A(n27910), .B(n36701), .Z(n27767) );
  NAND U28440 ( .A(n27765), .B(n36702), .Z(n27766) );
  NAND U28441 ( .A(n27767), .B(n27766), .Z(n27874) );
  XOR U28442 ( .A(b[25]), .B(a[175]), .Z(n27913) );
  NAND U28443 ( .A(n27913), .B(n38325), .Z(n27770) );
  NAND U28444 ( .A(n27768), .B(n38326), .Z(n27769) );
  AND U28445 ( .A(n27770), .B(n27769), .Z(n27875) );
  XNOR U28446 ( .A(n27874), .B(n27875), .Z(n27876) );
  XOR U28447 ( .A(n27877), .B(n27876), .Z(n27850) );
  XOR U28448 ( .A(n27853), .B(n27852), .Z(n27865) );
  XOR U28449 ( .A(n27864), .B(n27865), .Z(n27922) );
  XOR U28450 ( .A(n27923), .B(n27922), .Z(n27924) );
  XNOR U28451 ( .A(n27925), .B(n27924), .Z(n27934) );
  XNOR U28452 ( .A(n27935), .B(n27934), .Z(n27936) );
  XOR U28453 ( .A(n27937), .B(n27936), .Z(n27931) );
  NANDN U28454 ( .A(n27772), .B(n27771), .Z(n27776) );
  OR U28455 ( .A(n27774), .B(n27773), .Z(n27775) );
  NAND U28456 ( .A(n27776), .B(n27775), .Z(n27928) );
  NANDN U28457 ( .A(n27778), .B(n27777), .Z(n27782) );
  NAND U28458 ( .A(n27780), .B(n27779), .Z(n27781) );
  NAND U28459 ( .A(n27782), .B(n27781), .Z(n27929) );
  XNOR U28460 ( .A(n27928), .B(n27929), .Z(n27930) );
  XNOR U28461 ( .A(n27931), .B(n27930), .Z(n27807) );
  NANDN U28462 ( .A(n27784), .B(n27783), .Z(n27788) );
  NAND U28463 ( .A(n27786), .B(n27785), .Z(n27787) );
  NAND U28464 ( .A(n27788), .B(n27787), .Z(n27804) );
  NANDN U28465 ( .A(n27790), .B(n27789), .Z(n27794) );
  OR U28466 ( .A(n27792), .B(n27791), .Z(n27793) );
  NAND U28467 ( .A(n27794), .B(n27793), .Z(n27805) );
  XNOR U28468 ( .A(n27804), .B(n27805), .Z(n27806) );
  XNOR U28469 ( .A(n27807), .B(n27806), .Z(n27800) );
  XOR U28470 ( .A(n27801), .B(n27800), .Z(n27802) );
  XNOR U28471 ( .A(n27803), .B(n27802), .Z(n27940) );
  XNOR U28472 ( .A(n27940), .B(sreg[423]), .Z(n27942) );
  NAND U28473 ( .A(n27795), .B(sreg[422]), .Z(n27799) );
  OR U28474 ( .A(n27797), .B(n27796), .Z(n27798) );
  AND U28475 ( .A(n27799), .B(n27798), .Z(n27941) );
  XOR U28476 ( .A(n27942), .B(n27941), .Z(c[423]) );
  NANDN U28477 ( .A(n27805), .B(n27804), .Z(n27809) );
  NANDN U28478 ( .A(n27807), .B(n27806), .Z(n27808) );
  NAND U28479 ( .A(n27809), .B(n27808), .Z(n27946) );
  NANDN U28480 ( .A(n27811), .B(n27810), .Z(n27815) );
  NAND U28481 ( .A(n27813), .B(n27812), .Z(n27814) );
  NAND U28482 ( .A(n27815), .B(n27814), .Z(n28028) );
  XNOR U28483 ( .A(b[19]), .B(a[182]), .Z(n27973) );
  NANDN U28484 ( .A(n27973), .B(n37934), .Z(n27818) );
  NANDN U28485 ( .A(n27816), .B(n37935), .Z(n27817) );
  NAND U28486 ( .A(n27818), .B(n27817), .Z(n28038) );
  XOR U28487 ( .A(b[27]), .B(a[174]), .Z(n27976) );
  NAND U28488 ( .A(n38423), .B(n27976), .Z(n27821) );
  NAND U28489 ( .A(n27819), .B(n38424), .Z(n27820) );
  NAND U28490 ( .A(n27821), .B(n27820), .Z(n28035) );
  XNOR U28491 ( .A(b[5]), .B(a[196]), .Z(n27979) );
  NANDN U28492 ( .A(n27979), .B(n36587), .Z(n27824) );
  NANDN U28493 ( .A(n27822), .B(n36588), .Z(n27823) );
  AND U28494 ( .A(n27824), .B(n27823), .Z(n28036) );
  XNOR U28495 ( .A(n28035), .B(n28036), .Z(n28037) );
  XNOR U28496 ( .A(n28038), .B(n28037), .Z(n28026) );
  NAND U28497 ( .A(n27825), .B(n37762), .Z(n27827) );
  XOR U28498 ( .A(b[17]), .B(a[184]), .Z(n27982) );
  NAND U28499 ( .A(n27982), .B(n37764), .Z(n27826) );
  NAND U28500 ( .A(n27827), .B(n27826), .Z(n28000) );
  XNOR U28501 ( .A(b[31]), .B(a[170]), .Z(n27985) );
  NANDN U28502 ( .A(n27985), .B(n38552), .Z(n27830) );
  NANDN U28503 ( .A(n27828), .B(n38553), .Z(n27829) );
  NAND U28504 ( .A(n27830), .B(n27829), .Z(n27997) );
  OR U28505 ( .A(n27831), .B(n36105), .Z(n27833) );
  XOR U28506 ( .A(b[3]), .B(n32246), .Z(n27988) );
  NANDN U28507 ( .A(n27988), .B(n36107), .Z(n27832) );
  AND U28508 ( .A(n27833), .B(n27832), .Z(n27998) );
  XNOR U28509 ( .A(n27997), .B(n27998), .Z(n27999) );
  XOR U28510 ( .A(n28000), .B(n27999), .Z(n28025) );
  XNOR U28511 ( .A(n28026), .B(n28025), .Z(n28027) );
  XNOR U28512 ( .A(n28028), .B(n28027), .Z(n27964) );
  NANDN U28513 ( .A(n27835), .B(n27834), .Z(n27839) );
  NAND U28514 ( .A(n27837), .B(n27836), .Z(n27838) );
  NAND U28515 ( .A(n27839), .B(n27838), .Z(n28017) );
  NANDN U28516 ( .A(n27841), .B(n27840), .Z(n27845) );
  NAND U28517 ( .A(n27843), .B(n27842), .Z(n27844) );
  NAND U28518 ( .A(n27845), .B(n27844), .Z(n28016) );
  XNOR U28519 ( .A(n28016), .B(n28015), .Z(n28018) );
  XOR U28520 ( .A(n28017), .B(n28018), .Z(n27963) );
  XOR U28521 ( .A(n27964), .B(n27963), .Z(n27965) );
  NANDN U28522 ( .A(n27851), .B(n27850), .Z(n27855) );
  NAND U28523 ( .A(n27853), .B(n27852), .Z(n27854) );
  NAND U28524 ( .A(n27855), .B(n27854), .Z(n27966) );
  XNOR U28525 ( .A(n27965), .B(n27966), .Z(n28079) );
  OR U28526 ( .A(n27857), .B(n27856), .Z(n27861) );
  NANDN U28527 ( .A(n27859), .B(n27858), .Z(n27860) );
  NAND U28528 ( .A(n27861), .B(n27860), .Z(n28078) );
  NANDN U28529 ( .A(n27863), .B(n27862), .Z(n27867) );
  NAND U28530 ( .A(n27865), .B(n27864), .Z(n27866) );
  NAND U28531 ( .A(n27867), .B(n27866), .Z(n27959) );
  NANDN U28532 ( .A(n27869), .B(n27868), .Z(n27873) );
  NAND U28533 ( .A(n27871), .B(n27870), .Z(n27872) );
  NAND U28534 ( .A(n27873), .B(n27872), .Z(n27958) );
  NANDN U28535 ( .A(n27875), .B(n27874), .Z(n27879) );
  NAND U28536 ( .A(n27877), .B(n27876), .Z(n27878) );
  NAND U28537 ( .A(n27879), .B(n27878), .Z(n28019) );
  NANDN U28538 ( .A(n27881), .B(n27880), .Z(n27885) );
  NAND U28539 ( .A(n27883), .B(n27882), .Z(n27884) );
  AND U28540 ( .A(n27885), .B(n27884), .Z(n28020) );
  XNOR U28541 ( .A(n28019), .B(n28020), .Z(n28021) );
  XNOR U28542 ( .A(b[9]), .B(a[192]), .Z(n28041) );
  NANDN U28543 ( .A(n28041), .B(n36925), .Z(n27888) );
  NANDN U28544 ( .A(n27886), .B(n36926), .Z(n27887) );
  NAND U28545 ( .A(n27888), .B(n27887), .Z(n28005) );
  XNOR U28546 ( .A(b[15]), .B(a[186]), .Z(n28044) );
  OR U28547 ( .A(n28044), .B(n37665), .Z(n27891) );
  NAND U28548 ( .A(n27889), .B(n37604), .Z(n27890) );
  AND U28549 ( .A(n27891), .B(n27890), .Z(n28003) );
  XNOR U28550 ( .A(b[21]), .B(a[180]), .Z(n28047) );
  NANDN U28551 ( .A(n28047), .B(n38101), .Z(n27894) );
  NANDN U28552 ( .A(n27892), .B(n38102), .Z(n27893) );
  AND U28553 ( .A(n27894), .B(n27893), .Z(n28004) );
  XOR U28554 ( .A(n28005), .B(n28006), .Z(n27994) );
  XNOR U28555 ( .A(b[11]), .B(a[190]), .Z(n28050) );
  OR U28556 ( .A(n28050), .B(n37311), .Z(n27897) );
  NANDN U28557 ( .A(n27895), .B(n37218), .Z(n27896) );
  NAND U28558 ( .A(n27897), .B(n27896), .Z(n27992) );
  XOR U28559 ( .A(n1053), .B(a[188]), .Z(n28053) );
  NANDN U28560 ( .A(n28053), .B(n37424), .Z(n27900) );
  NANDN U28561 ( .A(n27898), .B(n37425), .Z(n27899) );
  AND U28562 ( .A(n27900), .B(n27899), .Z(n27991) );
  XNOR U28563 ( .A(n27992), .B(n27991), .Z(n27993) );
  XOR U28564 ( .A(n27994), .B(n27993), .Z(n28011) );
  NANDN U28565 ( .A(n1049), .B(a[200]), .Z(n27901) );
  XNOR U28566 ( .A(b[1]), .B(n27901), .Z(n27903) );
  NANDN U28567 ( .A(b[0]), .B(a[199]), .Z(n27902) );
  AND U28568 ( .A(n27903), .B(n27902), .Z(n27969) );
  NAND U28569 ( .A(n38490), .B(n27904), .Z(n27906) );
  XNOR U28570 ( .A(n1058), .B(a[172]), .Z(n28056) );
  NANDN U28571 ( .A(n1048), .B(n28056), .Z(n27905) );
  NAND U28572 ( .A(n27906), .B(n27905), .Z(n27967) );
  NANDN U28573 ( .A(n1059), .B(a[168]), .Z(n27968) );
  XNOR U28574 ( .A(n27967), .B(n27968), .Z(n27970) );
  XOR U28575 ( .A(n27969), .B(n27970), .Z(n28009) );
  NANDN U28576 ( .A(n27907), .B(n38205), .Z(n27909) );
  XNOR U28577 ( .A(b[23]), .B(a[178]), .Z(n28062) );
  OR U28578 ( .A(n28062), .B(n38268), .Z(n27908) );
  NAND U28579 ( .A(n27909), .B(n27908), .Z(n28032) );
  XNOR U28580 ( .A(b[7]), .B(a[194]), .Z(n28065) );
  NANDN U28581 ( .A(n28065), .B(n36701), .Z(n27912) );
  NANDN U28582 ( .A(n27910), .B(n36702), .Z(n27911) );
  NAND U28583 ( .A(n27912), .B(n27911), .Z(n28029) );
  XOR U28584 ( .A(b[25]), .B(a[176]), .Z(n28068) );
  NAND U28585 ( .A(n28068), .B(n38325), .Z(n27915) );
  NAND U28586 ( .A(n27913), .B(n38326), .Z(n27914) );
  AND U28587 ( .A(n27915), .B(n27914), .Z(n28030) );
  XNOR U28588 ( .A(n28029), .B(n28030), .Z(n28031) );
  XNOR U28589 ( .A(n28032), .B(n28031), .Z(n28010) );
  XOR U28590 ( .A(n28009), .B(n28010), .Z(n28012) );
  XNOR U28591 ( .A(n28011), .B(n28012), .Z(n28022) );
  XNOR U28592 ( .A(n28021), .B(n28022), .Z(n27957) );
  XNOR U28593 ( .A(n27958), .B(n27957), .Z(n27960) );
  XNOR U28594 ( .A(n27959), .B(n27960), .Z(n28077) );
  XOR U28595 ( .A(n28078), .B(n28077), .Z(n28080) );
  NANDN U28596 ( .A(n27917), .B(n27916), .Z(n27921) );
  NAND U28597 ( .A(n27919), .B(n27918), .Z(n27920) );
  NAND U28598 ( .A(n27921), .B(n27920), .Z(n28072) );
  NAND U28599 ( .A(n27923), .B(n27922), .Z(n27927) );
  NANDN U28600 ( .A(n27925), .B(n27924), .Z(n27926) );
  AND U28601 ( .A(n27927), .B(n27926), .Z(n28071) );
  XNOR U28602 ( .A(n28072), .B(n28071), .Z(n28073) );
  XOR U28603 ( .A(n28074), .B(n28073), .Z(n27953) );
  NANDN U28604 ( .A(n27929), .B(n27928), .Z(n27933) );
  NAND U28605 ( .A(n27931), .B(n27930), .Z(n27932) );
  NAND U28606 ( .A(n27933), .B(n27932), .Z(n27951) );
  NANDN U28607 ( .A(n27935), .B(n27934), .Z(n27939) );
  NANDN U28608 ( .A(n27937), .B(n27936), .Z(n27938) );
  NAND U28609 ( .A(n27939), .B(n27938), .Z(n27952) );
  XNOR U28610 ( .A(n27951), .B(n27952), .Z(n27954) );
  XOR U28611 ( .A(n27953), .B(n27954), .Z(n27945) );
  XOR U28612 ( .A(n27946), .B(n27945), .Z(n27947) );
  XNOR U28613 ( .A(n27948), .B(n27947), .Z(n28083) );
  XNOR U28614 ( .A(n28083), .B(sreg[424]), .Z(n28085) );
  NAND U28615 ( .A(n27940), .B(sreg[423]), .Z(n27944) );
  OR U28616 ( .A(n27942), .B(n27941), .Z(n27943) );
  AND U28617 ( .A(n27944), .B(n27943), .Z(n28084) );
  XOR U28618 ( .A(n28085), .B(n28084), .Z(c[424]) );
  NAND U28619 ( .A(n27946), .B(n27945), .Z(n27950) );
  NAND U28620 ( .A(n27948), .B(n27947), .Z(n27949) );
  NAND U28621 ( .A(n27950), .B(n27949), .Z(n28091) );
  NANDN U28622 ( .A(n27952), .B(n27951), .Z(n27956) );
  NAND U28623 ( .A(n27954), .B(n27953), .Z(n27955) );
  NAND U28624 ( .A(n27956), .B(n27955), .Z(n28088) );
  NAND U28625 ( .A(n27958), .B(n27957), .Z(n27962) );
  NANDN U28626 ( .A(n27960), .B(n27959), .Z(n27961) );
  NAND U28627 ( .A(n27962), .B(n27961), .Z(n28100) );
  XNOR U28628 ( .A(n28100), .B(n28101), .Z(n28102) );
  NANDN U28629 ( .A(n27968), .B(n27967), .Z(n27972) );
  NAND U28630 ( .A(n27970), .B(n27969), .Z(n27971) );
  NAND U28631 ( .A(n27972), .B(n27971), .Z(n28175) );
  XNOR U28632 ( .A(b[19]), .B(a[183]), .Z(n28142) );
  NANDN U28633 ( .A(n28142), .B(n37934), .Z(n27975) );
  NANDN U28634 ( .A(n27973), .B(n37935), .Z(n27974) );
  NAND U28635 ( .A(n27975), .B(n27974), .Z(n28187) );
  XOR U28636 ( .A(b[27]), .B(a[175]), .Z(n28145) );
  NAND U28637 ( .A(n38423), .B(n28145), .Z(n27978) );
  NAND U28638 ( .A(n27976), .B(n38424), .Z(n27977) );
  NAND U28639 ( .A(n27978), .B(n27977), .Z(n28184) );
  XNOR U28640 ( .A(b[5]), .B(a[197]), .Z(n28148) );
  NANDN U28641 ( .A(n28148), .B(n36587), .Z(n27981) );
  NANDN U28642 ( .A(n27979), .B(n36588), .Z(n27980) );
  AND U28643 ( .A(n27981), .B(n27980), .Z(n28185) );
  XNOR U28644 ( .A(n28184), .B(n28185), .Z(n28186) );
  XNOR U28645 ( .A(n28187), .B(n28186), .Z(n28172) );
  NAND U28646 ( .A(n27982), .B(n37762), .Z(n27984) );
  XOR U28647 ( .A(b[17]), .B(a[185]), .Z(n28151) );
  NAND U28648 ( .A(n28151), .B(n37764), .Z(n27983) );
  NAND U28649 ( .A(n27984), .B(n27983), .Z(n28126) );
  XNOR U28650 ( .A(b[31]), .B(a[171]), .Z(n28154) );
  NANDN U28651 ( .A(n28154), .B(n38552), .Z(n27987) );
  NANDN U28652 ( .A(n27985), .B(n38553), .Z(n27986) );
  AND U28653 ( .A(n27987), .B(n27986), .Z(n28124) );
  OR U28654 ( .A(n27988), .B(n36105), .Z(n27990) );
  XNOR U28655 ( .A(b[3]), .B(a[199]), .Z(n28157) );
  NANDN U28656 ( .A(n28157), .B(n36107), .Z(n27989) );
  AND U28657 ( .A(n27990), .B(n27989), .Z(n28125) );
  XOR U28658 ( .A(n28126), .B(n28127), .Z(n28173) );
  XOR U28659 ( .A(n28172), .B(n28173), .Z(n28174) );
  XNOR U28660 ( .A(n28175), .B(n28174), .Z(n28220) );
  NANDN U28661 ( .A(n27992), .B(n27991), .Z(n27996) );
  NAND U28662 ( .A(n27994), .B(n27993), .Z(n27995) );
  NAND U28663 ( .A(n27996), .B(n27995), .Z(n28163) );
  NANDN U28664 ( .A(n27998), .B(n27997), .Z(n28002) );
  NAND U28665 ( .A(n28000), .B(n27999), .Z(n28001) );
  NAND U28666 ( .A(n28002), .B(n28001), .Z(n28161) );
  OR U28667 ( .A(n28004), .B(n28003), .Z(n28008) );
  NANDN U28668 ( .A(n28006), .B(n28005), .Z(n28007) );
  NAND U28669 ( .A(n28008), .B(n28007), .Z(n28160) );
  XNOR U28670 ( .A(n28163), .B(n28162), .Z(n28221) );
  XNOR U28671 ( .A(n28220), .B(n28221), .Z(n28222) );
  NANDN U28672 ( .A(n28010), .B(n28009), .Z(n28014) );
  OR U28673 ( .A(n28012), .B(n28011), .Z(n28013) );
  AND U28674 ( .A(n28014), .B(n28013), .Z(n28223) );
  XOR U28675 ( .A(n28222), .B(n28223), .Z(n28108) );
  NANDN U28676 ( .A(n28020), .B(n28019), .Z(n28024) );
  NANDN U28677 ( .A(n28022), .B(n28021), .Z(n28023) );
  NAND U28678 ( .A(n28024), .B(n28023), .Z(n28229) );
  NANDN U28679 ( .A(n28030), .B(n28029), .Z(n28034) );
  NAND U28680 ( .A(n28032), .B(n28031), .Z(n28033) );
  NAND U28681 ( .A(n28034), .B(n28033), .Z(n28166) );
  NANDN U28682 ( .A(n28036), .B(n28035), .Z(n28040) );
  NAND U28683 ( .A(n28038), .B(n28037), .Z(n28039) );
  AND U28684 ( .A(n28040), .B(n28039), .Z(n28167) );
  XNOR U28685 ( .A(n28166), .B(n28167), .Z(n28168) );
  XOR U28686 ( .A(b[9]), .B(n31508), .Z(n28190) );
  NANDN U28687 ( .A(n28190), .B(n36925), .Z(n28043) );
  NANDN U28688 ( .A(n28041), .B(n36926), .Z(n28042) );
  NAND U28689 ( .A(n28043), .B(n28042), .Z(n28132) );
  XNOR U28690 ( .A(b[15]), .B(a[187]), .Z(n28193) );
  OR U28691 ( .A(n28193), .B(n37665), .Z(n28046) );
  NANDN U28692 ( .A(n28044), .B(n37604), .Z(n28045) );
  AND U28693 ( .A(n28046), .B(n28045), .Z(n28130) );
  XNOR U28694 ( .A(b[21]), .B(a[181]), .Z(n28196) );
  NANDN U28695 ( .A(n28196), .B(n38101), .Z(n28049) );
  NANDN U28696 ( .A(n28047), .B(n38102), .Z(n28048) );
  AND U28697 ( .A(n28049), .B(n28048), .Z(n28131) );
  XOR U28698 ( .A(n28132), .B(n28133), .Z(n28121) );
  XNOR U28699 ( .A(b[11]), .B(a[191]), .Z(n28199) );
  OR U28700 ( .A(n28199), .B(n37311), .Z(n28052) );
  NANDN U28701 ( .A(n28050), .B(n37218), .Z(n28051) );
  NAND U28702 ( .A(n28052), .B(n28051), .Z(n28119) );
  XOR U28703 ( .A(n1053), .B(a[189]), .Z(n28202) );
  NANDN U28704 ( .A(n28202), .B(n37424), .Z(n28055) );
  NANDN U28705 ( .A(n28053), .B(n37425), .Z(n28054) );
  NAND U28706 ( .A(n28055), .B(n28054), .Z(n28118) );
  XOR U28707 ( .A(n28121), .B(n28120), .Z(n28115) );
  NAND U28708 ( .A(n38490), .B(n28056), .Z(n28058) );
  XNOR U28709 ( .A(n1058), .B(a[173]), .Z(n28205) );
  NANDN U28710 ( .A(n1048), .B(n28205), .Z(n28057) );
  NAND U28711 ( .A(n28058), .B(n28057), .Z(n28136) );
  NANDN U28712 ( .A(n1059), .B(a[169]), .Z(n28137) );
  XNOR U28713 ( .A(n28136), .B(n28137), .Z(n28139) );
  NANDN U28714 ( .A(n1049), .B(a[201]), .Z(n28059) );
  XNOR U28715 ( .A(b[1]), .B(n28059), .Z(n28061) );
  NANDN U28716 ( .A(b[0]), .B(a[200]), .Z(n28060) );
  AND U28717 ( .A(n28061), .B(n28060), .Z(n28138) );
  XNOR U28718 ( .A(n28139), .B(n28138), .Z(n28113) );
  NANDN U28719 ( .A(n28062), .B(n38205), .Z(n28064) );
  XNOR U28720 ( .A(b[23]), .B(a[179]), .Z(n28211) );
  OR U28721 ( .A(n28211), .B(n38268), .Z(n28063) );
  NAND U28722 ( .A(n28064), .B(n28063), .Z(n28181) );
  XNOR U28723 ( .A(b[7]), .B(a[195]), .Z(n28214) );
  NANDN U28724 ( .A(n28214), .B(n36701), .Z(n28067) );
  NANDN U28725 ( .A(n28065), .B(n36702), .Z(n28066) );
  NAND U28726 ( .A(n28067), .B(n28066), .Z(n28178) );
  XOR U28727 ( .A(b[25]), .B(a[177]), .Z(n28217) );
  NAND U28728 ( .A(n28217), .B(n38325), .Z(n28070) );
  NAND U28729 ( .A(n28068), .B(n38326), .Z(n28069) );
  AND U28730 ( .A(n28070), .B(n28069), .Z(n28179) );
  XNOR U28731 ( .A(n28178), .B(n28179), .Z(n28180) );
  XOR U28732 ( .A(n28181), .B(n28180), .Z(n28112) );
  XOR U28733 ( .A(n28115), .B(n28114), .Z(n28169) );
  XNOR U28734 ( .A(n28168), .B(n28169), .Z(n28226) );
  XOR U28735 ( .A(n28227), .B(n28226), .Z(n28228) );
  XNOR U28736 ( .A(n28229), .B(n28228), .Z(n28106) );
  XNOR U28737 ( .A(n28107), .B(n28106), .Z(n28109) );
  XNOR U28738 ( .A(n28108), .B(n28109), .Z(n28103) );
  XOR U28739 ( .A(n28102), .B(n28103), .Z(n28097) );
  NANDN U28740 ( .A(n28072), .B(n28071), .Z(n28076) );
  NAND U28741 ( .A(n28074), .B(n28073), .Z(n28075) );
  NAND U28742 ( .A(n28076), .B(n28075), .Z(n28094) );
  NANDN U28743 ( .A(n28078), .B(n28077), .Z(n28082) );
  OR U28744 ( .A(n28080), .B(n28079), .Z(n28081) );
  NAND U28745 ( .A(n28082), .B(n28081), .Z(n28095) );
  XNOR U28746 ( .A(n28094), .B(n28095), .Z(n28096) );
  XNOR U28747 ( .A(n28097), .B(n28096), .Z(n28089) );
  XNOR U28748 ( .A(n28088), .B(n28089), .Z(n28090) );
  XNOR U28749 ( .A(n28091), .B(n28090), .Z(n28232) );
  XNOR U28750 ( .A(n28232), .B(sreg[425]), .Z(n28234) );
  NAND U28751 ( .A(n28083), .B(sreg[424]), .Z(n28087) );
  OR U28752 ( .A(n28085), .B(n28084), .Z(n28086) );
  AND U28753 ( .A(n28087), .B(n28086), .Z(n28233) );
  XOR U28754 ( .A(n28234), .B(n28233), .Z(c[425]) );
  NANDN U28755 ( .A(n28089), .B(n28088), .Z(n28093) );
  NAND U28756 ( .A(n28091), .B(n28090), .Z(n28092) );
  NAND U28757 ( .A(n28093), .B(n28092), .Z(n28240) );
  NANDN U28758 ( .A(n28095), .B(n28094), .Z(n28099) );
  NAND U28759 ( .A(n28097), .B(n28096), .Z(n28098) );
  NAND U28760 ( .A(n28099), .B(n28098), .Z(n28238) );
  NANDN U28761 ( .A(n28101), .B(n28100), .Z(n28105) );
  NANDN U28762 ( .A(n28103), .B(n28102), .Z(n28104) );
  NAND U28763 ( .A(n28105), .B(n28104), .Z(n28244) );
  OR U28764 ( .A(n28107), .B(n28106), .Z(n28111) );
  OR U28765 ( .A(n28109), .B(n28108), .Z(n28110) );
  AND U28766 ( .A(n28111), .B(n28110), .Z(n28243) );
  XNOR U28767 ( .A(n28244), .B(n28243), .Z(n28245) );
  NANDN U28768 ( .A(n28113), .B(n28112), .Z(n28117) );
  NANDN U28769 ( .A(n28115), .B(n28114), .Z(n28116) );
  NAND U28770 ( .A(n28117), .B(n28116), .Z(n28372) );
  OR U28771 ( .A(n28119), .B(n28118), .Z(n28123) );
  NAND U28772 ( .A(n28121), .B(n28120), .Z(n28122) );
  NAND U28773 ( .A(n28123), .B(n28122), .Z(n28311) );
  OR U28774 ( .A(n28125), .B(n28124), .Z(n28129) );
  NANDN U28775 ( .A(n28127), .B(n28126), .Z(n28128) );
  NAND U28776 ( .A(n28129), .B(n28128), .Z(n28310) );
  OR U28777 ( .A(n28131), .B(n28130), .Z(n28135) );
  NANDN U28778 ( .A(n28133), .B(n28132), .Z(n28134) );
  NAND U28779 ( .A(n28135), .B(n28134), .Z(n28309) );
  XOR U28780 ( .A(n28311), .B(n28312), .Z(n28369) );
  NANDN U28781 ( .A(n28137), .B(n28136), .Z(n28141) );
  NAND U28782 ( .A(n28139), .B(n28138), .Z(n28140) );
  NAND U28783 ( .A(n28141), .B(n28140), .Z(n28324) );
  XNOR U28784 ( .A(b[19]), .B(a[184]), .Z(n28291) );
  NANDN U28785 ( .A(n28291), .B(n37934), .Z(n28144) );
  NANDN U28786 ( .A(n28142), .B(n37935), .Z(n28143) );
  NAND U28787 ( .A(n28144), .B(n28143), .Z(n28336) );
  XOR U28788 ( .A(b[27]), .B(a[176]), .Z(n28294) );
  NAND U28789 ( .A(n38423), .B(n28294), .Z(n28147) );
  NAND U28790 ( .A(n28145), .B(n38424), .Z(n28146) );
  NAND U28791 ( .A(n28147), .B(n28146), .Z(n28333) );
  XOR U28792 ( .A(b[5]), .B(n32246), .Z(n28297) );
  NANDN U28793 ( .A(n28297), .B(n36587), .Z(n28150) );
  NANDN U28794 ( .A(n28148), .B(n36588), .Z(n28149) );
  AND U28795 ( .A(n28150), .B(n28149), .Z(n28334) );
  XNOR U28796 ( .A(n28333), .B(n28334), .Z(n28335) );
  XNOR U28797 ( .A(n28336), .B(n28335), .Z(n28321) );
  NAND U28798 ( .A(n28151), .B(n37762), .Z(n28153) );
  XOR U28799 ( .A(b[17]), .B(a[186]), .Z(n28300) );
  NAND U28800 ( .A(n28300), .B(n37764), .Z(n28152) );
  NAND U28801 ( .A(n28153), .B(n28152), .Z(n28275) );
  XNOR U28802 ( .A(b[31]), .B(a[172]), .Z(n28303) );
  NANDN U28803 ( .A(n28303), .B(n38552), .Z(n28156) );
  NANDN U28804 ( .A(n28154), .B(n38553), .Z(n28155) );
  AND U28805 ( .A(n28156), .B(n28155), .Z(n28273) );
  OR U28806 ( .A(n28157), .B(n36105), .Z(n28159) );
  XNOR U28807 ( .A(b[3]), .B(a[200]), .Z(n28306) );
  NANDN U28808 ( .A(n28306), .B(n36107), .Z(n28158) );
  AND U28809 ( .A(n28159), .B(n28158), .Z(n28274) );
  XOR U28810 ( .A(n28275), .B(n28276), .Z(n28322) );
  XOR U28811 ( .A(n28321), .B(n28322), .Z(n28323) );
  XNOR U28812 ( .A(n28324), .B(n28323), .Z(n28370) );
  XNOR U28813 ( .A(n28369), .B(n28370), .Z(n28371) );
  XNOR U28814 ( .A(n28372), .B(n28371), .Z(n28258) );
  OR U28815 ( .A(n28161), .B(n28160), .Z(n28165) );
  NAND U28816 ( .A(n28163), .B(n28162), .Z(n28164) );
  NAND U28817 ( .A(n28165), .B(n28164), .Z(n28256) );
  NANDN U28818 ( .A(n28167), .B(n28166), .Z(n28171) );
  NANDN U28819 ( .A(n28169), .B(n28168), .Z(n28170) );
  NAND U28820 ( .A(n28171), .B(n28170), .Z(n28377) );
  OR U28821 ( .A(n28173), .B(n28172), .Z(n28177) );
  NAND U28822 ( .A(n28175), .B(n28174), .Z(n28176) );
  NAND U28823 ( .A(n28177), .B(n28176), .Z(n28376) );
  NANDN U28824 ( .A(n28179), .B(n28178), .Z(n28183) );
  NAND U28825 ( .A(n28181), .B(n28180), .Z(n28182) );
  NAND U28826 ( .A(n28183), .B(n28182), .Z(n28315) );
  NANDN U28827 ( .A(n28185), .B(n28184), .Z(n28189) );
  NAND U28828 ( .A(n28187), .B(n28186), .Z(n28188) );
  AND U28829 ( .A(n28189), .B(n28188), .Z(n28316) );
  XNOR U28830 ( .A(n28315), .B(n28316), .Z(n28317) );
  XOR U28831 ( .A(b[9]), .B(n31644), .Z(n28339) );
  NANDN U28832 ( .A(n28339), .B(n36925), .Z(n28192) );
  NANDN U28833 ( .A(n28190), .B(n36926), .Z(n28191) );
  NAND U28834 ( .A(n28192), .B(n28191), .Z(n28281) );
  XNOR U28835 ( .A(b[15]), .B(a[188]), .Z(n28342) );
  OR U28836 ( .A(n28342), .B(n37665), .Z(n28195) );
  NANDN U28837 ( .A(n28193), .B(n37604), .Z(n28194) );
  AND U28838 ( .A(n28195), .B(n28194), .Z(n28279) );
  XNOR U28839 ( .A(b[21]), .B(a[182]), .Z(n28345) );
  NANDN U28840 ( .A(n28345), .B(n38101), .Z(n28198) );
  NANDN U28841 ( .A(n28196), .B(n38102), .Z(n28197) );
  AND U28842 ( .A(n28198), .B(n28197), .Z(n28280) );
  XOR U28843 ( .A(n28281), .B(n28282), .Z(n28270) );
  XNOR U28844 ( .A(b[11]), .B(a[192]), .Z(n28348) );
  OR U28845 ( .A(n28348), .B(n37311), .Z(n28201) );
  NANDN U28846 ( .A(n28199), .B(n37218), .Z(n28200) );
  NAND U28847 ( .A(n28201), .B(n28200), .Z(n28268) );
  XOR U28848 ( .A(n1053), .B(a[190]), .Z(n28351) );
  NANDN U28849 ( .A(n28351), .B(n37424), .Z(n28204) );
  NANDN U28850 ( .A(n28202), .B(n37425), .Z(n28203) );
  NAND U28851 ( .A(n28204), .B(n28203), .Z(n28267) );
  XOR U28852 ( .A(n28270), .B(n28269), .Z(n28264) );
  NAND U28853 ( .A(n38490), .B(n28205), .Z(n28207) );
  XNOR U28854 ( .A(n1058), .B(a[174]), .Z(n28357) );
  NANDN U28855 ( .A(n1048), .B(n28357), .Z(n28206) );
  NAND U28856 ( .A(n28207), .B(n28206), .Z(n28285) );
  NANDN U28857 ( .A(n1059), .B(a[170]), .Z(n28286) );
  XNOR U28858 ( .A(n28285), .B(n28286), .Z(n28288) );
  NANDN U28859 ( .A(n1049), .B(a[202]), .Z(n28208) );
  XNOR U28860 ( .A(b[1]), .B(n28208), .Z(n28210) );
  IV U28861 ( .A(a[201]), .Z(n32687) );
  NANDN U28862 ( .A(n32687), .B(n1049), .Z(n28209) );
  AND U28863 ( .A(n28210), .B(n28209), .Z(n28287) );
  XNOR U28864 ( .A(n28288), .B(n28287), .Z(n28262) );
  NANDN U28865 ( .A(n28211), .B(n38205), .Z(n28213) );
  XNOR U28866 ( .A(b[23]), .B(a[180]), .Z(n28360) );
  OR U28867 ( .A(n28360), .B(n38268), .Z(n28212) );
  NAND U28868 ( .A(n28213), .B(n28212), .Z(n28330) );
  XOR U28869 ( .A(b[7]), .B(a[196]), .Z(n28363) );
  NAND U28870 ( .A(n28363), .B(n36701), .Z(n28216) );
  NANDN U28871 ( .A(n28214), .B(n36702), .Z(n28215) );
  NAND U28872 ( .A(n28216), .B(n28215), .Z(n28327) );
  XOR U28873 ( .A(b[25]), .B(a[178]), .Z(n28366) );
  NAND U28874 ( .A(n28366), .B(n38325), .Z(n28219) );
  NAND U28875 ( .A(n28217), .B(n38326), .Z(n28218) );
  AND U28876 ( .A(n28219), .B(n28218), .Z(n28328) );
  XNOR U28877 ( .A(n28327), .B(n28328), .Z(n28329) );
  XOR U28878 ( .A(n28330), .B(n28329), .Z(n28261) );
  XOR U28879 ( .A(n28264), .B(n28263), .Z(n28318) );
  XNOR U28880 ( .A(n28317), .B(n28318), .Z(n28375) );
  XNOR U28881 ( .A(n28376), .B(n28375), .Z(n28378) );
  XNOR U28882 ( .A(n28377), .B(n28378), .Z(n28255) );
  XNOR U28883 ( .A(n28256), .B(n28255), .Z(n28257) );
  XOR U28884 ( .A(n28258), .B(n28257), .Z(n28252) );
  NANDN U28885 ( .A(n28221), .B(n28220), .Z(n28225) );
  NAND U28886 ( .A(n28223), .B(n28222), .Z(n28224) );
  NAND U28887 ( .A(n28225), .B(n28224), .Z(n28249) );
  NAND U28888 ( .A(n28227), .B(n28226), .Z(n28231) );
  NAND U28889 ( .A(n28229), .B(n28228), .Z(n28230) );
  NAND U28890 ( .A(n28231), .B(n28230), .Z(n28250) );
  XNOR U28891 ( .A(n28249), .B(n28250), .Z(n28251) );
  XOR U28892 ( .A(n28252), .B(n28251), .Z(n28246) );
  XOR U28893 ( .A(n28245), .B(n28246), .Z(n28237) );
  XOR U28894 ( .A(n28238), .B(n28237), .Z(n28239) );
  XNOR U28895 ( .A(n28240), .B(n28239), .Z(n28381) );
  XNOR U28896 ( .A(n28381), .B(sreg[426]), .Z(n28383) );
  NAND U28897 ( .A(n28232), .B(sreg[425]), .Z(n28236) );
  OR U28898 ( .A(n28234), .B(n28233), .Z(n28235) );
  AND U28899 ( .A(n28236), .B(n28235), .Z(n28382) );
  XOR U28900 ( .A(n28383), .B(n28382), .Z(c[426]) );
  NAND U28901 ( .A(n28238), .B(n28237), .Z(n28242) );
  NAND U28902 ( .A(n28240), .B(n28239), .Z(n28241) );
  NAND U28903 ( .A(n28242), .B(n28241), .Z(n28389) );
  NANDN U28904 ( .A(n28244), .B(n28243), .Z(n28248) );
  NAND U28905 ( .A(n28246), .B(n28245), .Z(n28247) );
  NAND U28906 ( .A(n28248), .B(n28247), .Z(n28387) );
  NANDN U28907 ( .A(n28250), .B(n28249), .Z(n28254) );
  NAND U28908 ( .A(n28252), .B(n28251), .Z(n28253) );
  NAND U28909 ( .A(n28254), .B(n28253), .Z(n28392) );
  NANDN U28910 ( .A(n28256), .B(n28255), .Z(n28260) );
  NANDN U28911 ( .A(n28258), .B(n28257), .Z(n28259) );
  NAND U28912 ( .A(n28260), .B(n28259), .Z(n28393) );
  XNOR U28913 ( .A(n28392), .B(n28393), .Z(n28394) );
  NANDN U28914 ( .A(n28262), .B(n28261), .Z(n28266) );
  NANDN U28915 ( .A(n28264), .B(n28263), .Z(n28265) );
  NAND U28916 ( .A(n28266), .B(n28265), .Z(n28521) );
  OR U28917 ( .A(n28268), .B(n28267), .Z(n28272) );
  NAND U28918 ( .A(n28270), .B(n28269), .Z(n28271) );
  NAND U28919 ( .A(n28272), .B(n28271), .Z(n28460) );
  OR U28920 ( .A(n28274), .B(n28273), .Z(n28278) );
  NANDN U28921 ( .A(n28276), .B(n28275), .Z(n28277) );
  NAND U28922 ( .A(n28278), .B(n28277), .Z(n28459) );
  OR U28923 ( .A(n28280), .B(n28279), .Z(n28284) );
  NANDN U28924 ( .A(n28282), .B(n28281), .Z(n28283) );
  NAND U28925 ( .A(n28284), .B(n28283), .Z(n28458) );
  XOR U28926 ( .A(n28460), .B(n28461), .Z(n28518) );
  NANDN U28927 ( .A(n28286), .B(n28285), .Z(n28290) );
  NAND U28928 ( .A(n28288), .B(n28287), .Z(n28289) );
  NAND U28929 ( .A(n28290), .B(n28289), .Z(n28473) );
  XNOR U28930 ( .A(b[19]), .B(a[185]), .Z(n28416) );
  NANDN U28931 ( .A(n28416), .B(n37934), .Z(n28293) );
  NANDN U28932 ( .A(n28291), .B(n37935), .Z(n28292) );
  NAND U28933 ( .A(n28293), .B(n28292), .Z(n28485) );
  XOR U28934 ( .A(b[27]), .B(a[177]), .Z(n28419) );
  NAND U28935 ( .A(n38423), .B(n28419), .Z(n28296) );
  NAND U28936 ( .A(n28294), .B(n38424), .Z(n28295) );
  NAND U28937 ( .A(n28296), .B(n28295), .Z(n28482) );
  XNOR U28938 ( .A(b[5]), .B(a[199]), .Z(n28422) );
  NANDN U28939 ( .A(n28422), .B(n36587), .Z(n28299) );
  NANDN U28940 ( .A(n28297), .B(n36588), .Z(n28298) );
  AND U28941 ( .A(n28299), .B(n28298), .Z(n28483) );
  XNOR U28942 ( .A(n28482), .B(n28483), .Z(n28484) );
  XNOR U28943 ( .A(n28485), .B(n28484), .Z(n28471) );
  NAND U28944 ( .A(n28300), .B(n37762), .Z(n28302) );
  XOR U28945 ( .A(b[17]), .B(a[187]), .Z(n28425) );
  NAND U28946 ( .A(n28425), .B(n37764), .Z(n28301) );
  NAND U28947 ( .A(n28302), .B(n28301), .Z(n28443) );
  XNOR U28948 ( .A(b[31]), .B(a[173]), .Z(n28428) );
  NANDN U28949 ( .A(n28428), .B(n38552), .Z(n28305) );
  NANDN U28950 ( .A(n28303), .B(n38553), .Z(n28304) );
  NAND U28951 ( .A(n28305), .B(n28304), .Z(n28440) );
  OR U28952 ( .A(n28306), .B(n36105), .Z(n28308) );
  XOR U28953 ( .A(b[3]), .B(n32687), .Z(n28431) );
  NANDN U28954 ( .A(n28431), .B(n36107), .Z(n28307) );
  AND U28955 ( .A(n28308), .B(n28307), .Z(n28441) );
  XNOR U28956 ( .A(n28440), .B(n28441), .Z(n28442) );
  XOR U28957 ( .A(n28443), .B(n28442), .Z(n28470) );
  XNOR U28958 ( .A(n28471), .B(n28470), .Z(n28472) );
  XNOR U28959 ( .A(n28473), .B(n28472), .Z(n28519) );
  XNOR U28960 ( .A(n28518), .B(n28519), .Z(n28520) );
  XNOR U28961 ( .A(n28521), .B(n28520), .Z(n28407) );
  OR U28962 ( .A(n28310), .B(n28309), .Z(n28314) );
  NANDN U28963 ( .A(n28312), .B(n28311), .Z(n28313) );
  NAND U28964 ( .A(n28314), .B(n28313), .Z(n28405) );
  NANDN U28965 ( .A(n28316), .B(n28315), .Z(n28320) );
  NANDN U28966 ( .A(n28318), .B(n28317), .Z(n28319) );
  NAND U28967 ( .A(n28320), .B(n28319), .Z(n28526) );
  OR U28968 ( .A(n28322), .B(n28321), .Z(n28326) );
  NAND U28969 ( .A(n28324), .B(n28323), .Z(n28325) );
  NAND U28970 ( .A(n28326), .B(n28325), .Z(n28525) );
  NANDN U28971 ( .A(n28328), .B(n28327), .Z(n28332) );
  NAND U28972 ( .A(n28330), .B(n28329), .Z(n28331) );
  NAND U28973 ( .A(n28332), .B(n28331), .Z(n28464) );
  NANDN U28974 ( .A(n28334), .B(n28333), .Z(n28338) );
  NAND U28975 ( .A(n28336), .B(n28335), .Z(n28337) );
  AND U28976 ( .A(n28338), .B(n28337), .Z(n28465) );
  XNOR U28977 ( .A(n28464), .B(n28465), .Z(n28466) );
  XOR U28978 ( .A(b[9]), .B(n31434), .Z(n28488) );
  NANDN U28979 ( .A(n28488), .B(n36925), .Z(n28341) );
  NANDN U28980 ( .A(n28339), .B(n36926), .Z(n28340) );
  NAND U28981 ( .A(n28341), .B(n28340), .Z(n28448) );
  XOR U28982 ( .A(b[15]), .B(n30936), .Z(n28491) );
  OR U28983 ( .A(n28491), .B(n37665), .Z(n28344) );
  NANDN U28984 ( .A(n28342), .B(n37604), .Z(n28343) );
  AND U28985 ( .A(n28344), .B(n28343), .Z(n28446) );
  XNOR U28986 ( .A(b[21]), .B(a[183]), .Z(n28494) );
  NANDN U28987 ( .A(n28494), .B(n38101), .Z(n28347) );
  NANDN U28988 ( .A(n28345), .B(n38102), .Z(n28346) );
  AND U28989 ( .A(n28347), .B(n28346), .Z(n28447) );
  XOR U28990 ( .A(n28448), .B(n28449), .Z(n28437) );
  XOR U28991 ( .A(b[11]), .B(n31508), .Z(n28497) );
  OR U28992 ( .A(n28497), .B(n37311), .Z(n28350) );
  NANDN U28993 ( .A(n28348), .B(n37218), .Z(n28349) );
  NAND U28994 ( .A(n28350), .B(n28349), .Z(n28435) );
  XOR U28995 ( .A(n1053), .B(a[191]), .Z(n28500) );
  NANDN U28996 ( .A(n28500), .B(n37424), .Z(n28353) );
  NANDN U28997 ( .A(n28351), .B(n37425), .Z(n28352) );
  AND U28998 ( .A(n28353), .B(n28352), .Z(n28434) );
  XNOR U28999 ( .A(n28435), .B(n28434), .Z(n28436) );
  XOR U29000 ( .A(n28437), .B(n28436), .Z(n28454) );
  NANDN U29001 ( .A(n1049), .B(a[203]), .Z(n28354) );
  XNOR U29002 ( .A(b[1]), .B(n28354), .Z(n28356) );
  NANDN U29003 ( .A(b[0]), .B(a[202]), .Z(n28355) );
  AND U29004 ( .A(n28356), .B(n28355), .Z(n28412) );
  NAND U29005 ( .A(n38490), .B(n28357), .Z(n28359) );
  XNOR U29006 ( .A(n1058), .B(a[175]), .Z(n28506) );
  NANDN U29007 ( .A(n1048), .B(n28506), .Z(n28358) );
  NAND U29008 ( .A(n28359), .B(n28358), .Z(n28410) );
  NANDN U29009 ( .A(n1059), .B(a[171]), .Z(n28411) );
  XNOR U29010 ( .A(n28410), .B(n28411), .Z(n28413) );
  XOR U29011 ( .A(n28412), .B(n28413), .Z(n28452) );
  NANDN U29012 ( .A(n28360), .B(n38205), .Z(n28362) );
  XNOR U29013 ( .A(b[23]), .B(a[181]), .Z(n28509) );
  OR U29014 ( .A(n28509), .B(n38268), .Z(n28361) );
  NAND U29015 ( .A(n28362), .B(n28361), .Z(n28479) );
  XOR U29016 ( .A(b[7]), .B(a[197]), .Z(n28512) );
  NAND U29017 ( .A(n28512), .B(n36701), .Z(n28365) );
  NAND U29018 ( .A(n28363), .B(n36702), .Z(n28364) );
  NAND U29019 ( .A(n28365), .B(n28364), .Z(n28476) );
  XOR U29020 ( .A(b[25]), .B(a[179]), .Z(n28515) );
  NAND U29021 ( .A(n28515), .B(n38325), .Z(n28368) );
  NAND U29022 ( .A(n28366), .B(n38326), .Z(n28367) );
  AND U29023 ( .A(n28368), .B(n28367), .Z(n28477) );
  XNOR U29024 ( .A(n28476), .B(n28477), .Z(n28478) );
  XNOR U29025 ( .A(n28479), .B(n28478), .Z(n28453) );
  XOR U29026 ( .A(n28452), .B(n28453), .Z(n28455) );
  XNOR U29027 ( .A(n28454), .B(n28455), .Z(n28467) );
  XNOR U29028 ( .A(n28466), .B(n28467), .Z(n28524) );
  XNOR U29029 ( .A(n28525), .B(n28524), .Z(n28527) );
  XNOR U29030 ( .A(n28526), .B(n28527), .Z(n28404) );
  XNOR U29031 ( .A(n28405), .B(n28404), .Z(n28406) );
  XOR U29032 ( .A(n28407), .B(n28406), .Z(n28401) );
  NANDN U29033 ( .A(n28370), .B(n28369), .Z(n28374) );
  NAND U29034 ( .A(n28372), .B(n28371), .Z(n28373) );
  NAND U29035 ( .A(n28374), .B(n28373), .Z(n28399) );
  NAND U29036 ( .A(n28376), .B(n28375), .Z(n28380) );
  NANDN U29037 ( .A(n28378), .B(n28377), .Z(n28379) );
  AND U29038 ( .A(n28380), .B(n28379), .Z(n28398) );
  XNOR U29039 ( .A(n28399), .B(n28398), .Z(n28400) );
  XOR U29040 ( .A(n28401), .B(n28400), .Z(n28395) );
  XOR U29041 ( .A(n28394), .B(n28395), .Z(n28386) );
  XOR U29042 ( .A(n28387), .B(n28386), .Z(n28388) );
  XNOR U29043 ( .A(n28389), .B(n28388), .Z(n28530) );
  XNOR U29044 ( .A(n28530), .B(sreg[427]), .Z(n28532) );
  NAND U29045 ( .A(n28381), .B(sreg[426]), .Z(n28385) );
  OR U29046 ( .A(n28383), .B(n28382), .Z(n28384) );
  AND U29047 ( .A(n28385), .B(n28384), .Z(n28531) );
  XOR U29048 ( .A(n28532), .B(n28531), .Z(c[427]) );
  NAND U29049 ( .A(n28387), .B(n28386), .Z(n28391) );
  NAND U29050 ( .A(n28389), .B(n28388), .Z(n28390) );
  NAND U29051 ( .A(n28391), .B(n28390), .Z(n28538) );
  NANDN U29052 ( .A(n28393), .B(n28392), .Z(n28397) );
  NAND U29053 ( .A(n28395), .B(n28394), .Z(n28396) );
  NAND U29054 ( .A(n28397), .B(n28396), .Z(n28536) );
  NANDN U29055 ( .A(n28399), .B(n28398), .Z(n28403) );
  NAND U29056 ( .A(n28401), .B(n28400), .Z(n28402) );
  NAND U29057 ( .A(n28403), .B(n28402), .Z(n28541) );
  NANDN U29058 ( .A(n28405), .B(n28404), .Z(n28409) );
  NANDN U29059 ( .A(n28407), .B(n28406), .Z(n28408) );
  NAND U29060 ( .A(n28409), .B(n28408), .Z(n28542) );
  XNOR U29061 ( .A(n28541), .B(n28542), .Z(n28543) );
  NANDN U29062 ( .A(n28411), .B(n28410), .Z(n28415) );
  NAND U29063 ( .A(n28413), .B(n28412), .Z(n28414) );
  NAND U29064 ( .A(n28415), .B(n28414), .Z(n28610) );
  XNOR U29065 ( .A(b[19]), .B(a[186]), .Z(n28553) );
  NANDN U29066 ( .A(n28553), .B(n37934), .Z(n28418) );
  NANDN U29067 ( .A(n28416), .B(n37935), .Z(n28417) );
  NAND U29068 ( .A(n28418), .B(n28417), .Z(n28620) );
  XOR U29069 ( .A(b[27]), .B(a[178]), .Z(n28556) );
  NAND U29070 ( .A(n38423), .B(n28556), .Z(n28421) );
  NAND U29071 ( .A(n28419), .B(n38424), .Z(n28420) );
  NAND U29072 ( .A(n28421), .B(n28420), .Z(n28617) );
  XNOR U29073 ( .A(b[5]), .B(a[200]), .Z(n28559) );
  NANDN U29074 ( .A(n28559), .B(n36587), .Z(n28424) );
  NANDN U29075 ( .A(n28422), .B(n36588), .Z(n28423) );
  AND U29076 ( .A(n28424), .B(n28423), .Z(n28618) );
  XNOR U29077 ( .A(n28617), .B(n28618), .Z(n28619) );
  XNOR U29078 ( .A(n28620), .B(n28619), .Z(n28608) );
  NAND U29079 ( .A(n28425), .B(n37762), .Z(n28427) );
  XOR U29080 ( .A(b[17]), .B(a[188]), .Z(n28562) );
  NAND U29081 ( .A(n28562), .B(n37764), .Z(n28426) );
  NAND U29082 ( .A(n28427), .B(n28426), .Z(n28580) );
  XNOR U29083 ( .A(b[31]), .B(a[174]), .Z(n28565) );
  NANDN U29084 ( .A(n28565), .B(n38552), .Z(n28430) );
  NANDN U29085 ( .A(n28428), .B(n38553), .Z(n28429) );
  NAND U29086 ( .A(n28430), .B(n28429), .Z(n28577) );
  OR U29087 ( .A(n28431), .B(n36105), .Z(n28433) );
  XNOR U29088 ( .A(b[3]), .B(a[202]), .Z(n28568) );
  NANDN U29089 ( .A(n28568), .B(n36107), .Z(n28432) );
  AND U29090 ( .A(n28433), .B(n28432), .Z(n28578) );
  XNOR U29091 ( .A(n28577), .B(n28578), .Z(n28579) );
  XOR U29092 ( .A(n28580), .B(n28579), .Z(n28607) );
  XNOR U29093 ( .A(n28608), .B(n28607), .Z(n28609) );
  XNOR U29094 ( .A(n28610), .B(n28609), .Z(n28653) );
  NANDN U29095 ( .A(n28435), .B(n28434), .Z(n28439) );
  NAND U29096 ( .A(n28437), .B(n28436), .Z(n28438) );
  NAND U29097 ( .A(n28439), .B(n28438), .Z(n28598) );
  NANDN U29098 ( .A(n28441), .B(n28440), .Z(n28445) );
  NAND U29099 ( .A(n28443), .B(n28442), .Z(n28444) );
  NAND U29100 ( .A(n28445), .B(n28444), .Z(n28596) );
  OR U29101 ( .A(n28447), .B(n28446), .Z(n28451) );
  NANDN U29102 ( .A(n28449), .B(n28448), .Z(n28450) );
  NAND U29103 ( .A(n28451), .B(n28450), .Z(n28595) );
  XNOR U29104 ( .A(n28598), .B(n28597), .Z(n28654) );
  XOR U29105 ( .A(n28653), .B(n28654), .Z(n28656) );
  NANDN U29106 ( .A(n28453), .B(n28452), .Z(n28457) );
  OR U29107 ( .A(n28455), .B(n28454), .Z(n28456) );
  NAND U29108 ( .A(n28457), .B(n28456), .Z(n28655) );
  XOR U29109 ( .A(n28656), .B(n28655), .Z(n28673) );
  OR U29110 ( .A(n28459), .B(n28458), .Z(n28463) );
  NANDN U29111 ( .A(n28461), .B(n28460), .Z(n28462) );
  NAND U29112 ( .A(n28463), .B(n28462), .Z(n28672) );
  NANDN U29113 ( .A(n28465), .B(n28464), .Z(n28469) );
  NANDN U29114 ( .A(n28467), .B(n28466), .Z(n28468) );
  NAND U29115 ( .A(n28469), .B(n28468), .Z(n28661) );
  NANDN U29116 ( .A(n28471), .B(n28470), .Z(n28475) );
  NAND U29117 ( .A(n28473), .B(n28472), .Z(n28474) );
  NAND U29118 ( .A(n28475), .B(n28474), .Z(n28660) );
  NANDN U29119 ( .A(n28477), .B(n28476), .Z(n28481) );
  NAND U29120 ( .A(n28479), .B(n28478), .Z(n28480) );
  NAND U29121 ( .A(n28481), .B(n28480), .Z(n28601) );
  NANDN U29122 ( .A(n28483), .B(n28482), .Z(n28487) );
  NAND U29123 ( .A(n28485), .B(n28484), .Z(n28486) );
  AND U29124 ( .A(n28487), .B(n28486), .Z(n28602) );
  XNOR U29125 ( .A(n28601), .B(n28602), .Z(n28603) );
  XNOR U29126 ( .A(n1052), .B(a[196]), .Z(n28629) );
  NAND U29127 ( .A(n36925), .B(n28629), .Z(n28490) );
  NANDN U29128 ( .A(n28488), .B(n36926), .Z(n28489) );
  NAND U29129 ( .A(n28490), .B(n28489), .Z(n28585) );
  XNOR U29130 ( .A(b[15]), .B(a[190]), .Z(n28626) );
  OR U29131 ( .A(n28626), .B(n37665), .Z(n28493) );
  NANDN U29132 ( .A(n28491), .B(n37604), .Z(n28492) );
  AND U29133 ( .A(n28493), .B(n28492), .Z(n28583) );
  XNOR U29134 ( .A(n1056), .B(a[184]), .Z(n28623) );
  NAND U29135 ( .A(n28623), .B(n38101), .Z(n28496) );
  NANDN U29136 ( .A(n28494), .B(n38102), .Z(n28495) );
  AND U29137 ( .A(n28496), .B(n28495), .Z(n28584) );
  XOR U29138 ( .A(n28585), .B(n28586), .Z(n28574) );
  XOR U29139 ( .A(b[11]), .B(n31644), .Z(n28632) );
  OR U29140 ( .A(n28632), .B(n37311), .Z(n28499) );
  NANDN U29141 ( .A(n28497), .B(n37218), .Z(n28498) );
  NAND U29142 ( .A(n28499), .B(n28498), .Z(n28572) );
  XOR U29143 ( .A(n1053), .B(a[192]), .Z(n28635) );
  NANDN U29144 ( .A(n28635), .B(n37424), .Z(n28502) );
  NANDN U29145 ( .A(n28500), .B(n37425), .Z(n28501) );
  AND U29146 ( .A(n28502), .B(n28501), .Z(n28571) );
  XNOR U29147 ( .A(n28572), .B(n28571), .Z(n28573) );
  XOR U29148 ( .A(n28574), .B(n28573), .Z(n28591) );
  NANDN U29149 ( .A(n1049), .B(a[204]), .Z(n28503) );
  XNOR U29150 ( .A(b[1]), .B(n28503), .Z(n28505) );
  NANDN U29151 ( .A(b[0]), .B(a[203]), .Z(n28504) );
  AND U29152 ( .A(n28505), .B(n28504), .Z(n28549) );
  NAND U29153 ( .A(n38490), .B(n28506), .Z(n28508) );
  XNOR U29154 ( .A(n1058), .B(a[176]), .Z(n28641) );
  NANDN U29155 ( .A(n1048), .B(n28641), .Z(n28507) );
  NAND U29156 ( .A(n28508), .B(n28507), .Z(n28547) );
  NANDN U29157 ( .A(n1059), .B(a[172]), .Z(n28548) );
  XNOR U29158 ( .A(n28547), .B(n28548), .Z(n28550) );
  XOR U29159 ( .A(n28549), .B(n28550), .Z(n28589) );
  NANDN U29160 ( .A(n28509), .B(n38205), .Z(n28511) );
  XNOR U29161 ( .A(b[23]), .B(a[182]), .Z(n28644) );
  OR U29162 ( .A(n28644), .B(n38268), .Z(n28510) );
  NAND U29163 ( .A(n28511), .B(n28510), .Z(n28614) );
  XNOR U29164 ( .A(b[7]), .B(a[198]), .Z(n28647) );
  NANDN U29165 ( .A(n28647), .B(n36701), .Z(n28514) );
  NAND U29166 ( .A(n28512), .B(n36702), .Z(n28513) );
  NAND U29167 ( .A(n28514), .B(n28513), .Z(n28611) );
  XOR U29168 ( .A(b[25]), .B(a[180]), .Z(n28650) );
  NAND U29169 ( .A(n28650), .B(n38325), .Z(n28517) );
  NAND U29170 ( .A(n28515), .B(n38326), .Z(n28516) );
  AND U29171 ( .A(n28517), .B(n28516), .Z(n28612) );
  XNOR U29172 ( .A(n28611), .B(n28612), .Z(n28613) );
  XNOR U29173 ( .A(n28614), .B(n28613), .Z(n28590) );
  XOR U29174 ( .A(n28589), .B(n28590), .Z(n28592) );
  XNOR U29175 ( .A(n28591), .B(n28592), .Z(n28604) );
  XNOR U29176 ( .A(n28603), .B(n28604), .Z(n28659) );
  XNOR U29177 ( .A(n28660), .B(n28659), .Z(n28662) );
  XNOR U29178 ( .A(n28661), .B(n28662), .Z(n28671) );
  XOR U29179 ( .A(n28672), .B(n28671), .Z(n28674) );
  NANDN U29180 ( .A(n28519), .B(n28518), .Z(n28523) );
  NAND U29181 ( .A(n28521), .B(n28520), .Z(n28522) );
  NAND U29182 ( .A(n28523), .B(n28522), .Z(n28666) );
  NAND U29183 ( .A(n28525), .B(n28524), .Z(n28529) );
  NANDN U29184 ( .A(n28527), .B(n28526), .Z(n28528) );
  AND U29185 ( .A(n28529), .B(n28528), .Z(n28665) );
  XNOR U29186 ( .A(n28666), .B(n28665), .Z(n28667) );
  XOR U29187 ( .A(n28668), .B(n28667), .Z(n28544) );
  XOR U29188 ( .A(n28543), .B(n28544), .Z(n28535) );
  XOR U29189 ( .A(n28536), .B(n28535), .Z(n28537) );
  XNOR U29190 ( .A(n28538), .B(n28537), .Z(n28677) );
  XNOR U29191 ( .A(n28677), .B(sreg[428]), .Z(n28679) );
  NAND U29192 ( .A(n28530), .B(sreg[427]), .Z(n28534) );
  OR U29193 ( .A(n28532), .B(n28531), .Z(n28533) );
  AND U29194 ( .A(n28534), .B(n28533), .Z(n28678) );
  XOR U29195 ( .A(n28679), .B(n28678), .Z(c[428]) );
  NAND U29196 ( .A(n28536), .B(n28535), .Z(n28540) );
  NAND U29197 ( .A(n28538), .B(n28537), .Z(n28539) );
  NAND U29198 ( .A(n28540), .B(n28539), .Z(n28685) );
  NANDN U29199 ( .A(n28542), .B(n28541), .Z(n28546) );
  NAND U29200 ( .A(n28544), .B(n28543), .Z(n28545) );
  NAND U29201 ( .A(n28546), .B(n28545), .Z(n28683) );
  NANDN U29202 ( .A(n28548), .B(n28547), .Z(n28552) );
  NAND U29203 ( .A(n28550), .B(n28549), .Z(n28551) );
  NAND U29204 ( .A(n28552), .B(n28551), .Z(n28767) );
  XNOR U29205 ( .A(b[19]), .B(a[187]), .Z(n28712) );
  NANDN U29206 ( .A(n28712), .B(n37934), .Z(n28555) );
  NANDN U29207 ( .A(n28553), .B(n37935), .Z(n28554) );
  NAND U29208 ( .A(n28555), .B(n28554), .Z(n28777) );
  XOR U29209 ( .A(b[27]), .B(a[179]), .Z(n28715) );
  NAND U29210 ( .A(n38423), .B(n28715), .Z(n28558) );
  NAND U29211 ( .A(n28556), .B(n38424), .Z(n28557) );
  NAND U29212 ( .A(n28558), .B(n28557), .Z(n28774) );
  XOR U29213 ( .A(b[5]), .B(n32687), .Z(n28718) );
  NANDN U29214 ( .A(n28718), .B(n36587), .Z(n28561) );
  NANDN U29215 ( .A(n28559), .B(n36588), .Z(n28560) );
  AND U29216 ( .A(n28561), .B(n28560), .Z(n28775) );
  XNOR U29217 ( .A(n28774), .B(n28775), .Z(n28776) );
  XNOR U29218 ( .A(n28777), .B(n28776), .Z(n28765) );
  NAND U29219 ( .A(n28562), .B(n37762), .Z(n28564) );
  XNOR U29220 ( .A(b[17]), .B(a[189]), .Z(n28721) );
  NANDN U29221 ( .A(n28721), .B(n37764), .Z(n28563) );
  NAND U29222 ( .A(n28564), .B(n28563), .Z(n28739) );
  XNOR U29223 ( .A(b[31]), .B(a[175]), .Z(n28724) );
  NANDN U29224 ( .A(n28724), .B(n38552), .Z(n28567) );
  NANDN U29225 ( .A(n28565), .B(n38553), .Z(n28566) );
  NAND U29226 ( .A(n28567), .B(n28566), .Z(n28736) );
  OR U29227 ( .A(n28568), .B(n36105), .Z(n28570) );
  XNOR U29228 ( .A(b[3]), .B(a[203]), .Z(n28727) );
  NANDN U29229 ( .A(n28727), .B(n36107), .Z(n28569) );
  AND U29230 ( .A(n28570), .B(n28569), .Z(n28737) );
  XNOR U29231 ( .A(n28736), .B(n28737), .Z(n28738) );
  XOR U29232 ( .A(n28739), .B(n28738), .Z(n28764) );
  XNOR U29233 ( .A(n28765), .B(n28764), .Z(n28766) );
  XNOR U29234 ( .A(n28767), .B(n28766), .Z(n28810) );
  NANDN U29235 ( .A(n28572), .B(n28571), .Z(n28576) );
  NAND U29236 ( .A(n28574), .B(n28573), .Z(n28575) );
  NAND U29237 ( .A(n28576), .B(n28575), .Z(n28755) );
  NANDN U29238 ( .A(n28578), .B(n28577), .Z(n28582) );
  NAND U29239 ( .A(n28580), .B(n28579), .Z(n28581) );
  NAND U29240 ( .A(n28582), .B(n28581), .Z(n28753) );
  OR U29241 ( .A(n28584), .B(n28583), .Z(n28588) );
  NANDN U29242 ( .A(n28586), .B(n28585), .Z(n28587) );
  NAND U29243 ( .A(n28588), .B(n28587), .Z(n28752) );
  XNOR U29244 ( .A(n28755), .B(n28754), .Z(n28811) );
  XOR U29245 ( .A(n28810), .B(n28811), .Z(n28813) );
  NANDN U29246 ( .A(n28590), .B(n28589), .Z(n28594) );
  OR U29247 ( .A(n28592), .B(n28591), .Z(n28593) );
  NAND U29248 ( .A(n28594), .B(n28593), .Z(n28812) );
  XOR U29249 ( .A(n28813), .B(n28812), .Z(n28702) );
  OR U29250 ( .A(n28596), .B(n28595), .Z(n28600) );
  NAND U29251 ( .A(n28598), .B(n28597), .Z(n28599) );
  NAND U29252 ( .A(n28600), .B(n28599), .Z(n28701) );
  NANDN U29253 ( .A(n28602), .B(n28601), .Z(n28606) );
  NANDN U29254 ( .A(n28604), .B(n28603), .Z(n28605) );
  NAND U29255 ( .A(n28606), .B(n28605), .Z(n28818) );
  NANDN U29256 ( .A(n28612), .B(n28611), .Z(n28616) );
  NAND U29257 ( .A(n28614), .B(n28613), .Z(n28615) );
  NAND U29258 ( .A(n28616), .B(n28615), .Z(n28758) );
  NANDN U29259 ( .A(n28618), .B(n28617), .Z(n28622) );
  NAND U29260 ( .A(n28620), .B(n28619), .Z(n28621) );
  AND U29261 ( .A(n28622), .B(n28621), .Z(n28759) );
  XNOR U29262 ( .A(n28758), .B(n28759), .Z(n28760) );
  XNOR U29263 ( .A(b[21]), .B(a[185]), .Z(n28786) );
  NANDN U29264 ( .A(n28786), .B(n38101), .Z(n28625) );
  NAND U29265 ( .A(n38102), .B(n28623), .Z(n28624) );
  NAND U29266 ( .A(n28625), .B(n28624), .Z(n28748) );
  XNOR U29267 ( .A(b[15]), .B(a[191]), .Z(n28783) );
  OR U29268 ( .A(n28783), .B(n37665), .Z(n28628) );
  NANDN U29269 ( .A(n28626), .B(n37604), .Z(n28627) );
  AND U29270 ( .A(n28628), .B(n28627), .Z(n28749) );
  XNOR U29271 ( .A(n28748), .B(n28749), .Z(n28751) );
  XNOR U29272 ( .A(b[9]), .B(a[197]), .Z(n28780) );
  NANDN U29273 ( .A(n28780), .B(n36925), .Z(n28631) );
  NAND U29274 ( .A(n36926), .B(n28629), .Z(n28630) );
  NAND U29275 ( .A(n28631), .B(n28630), .Z(n28750) );
  XNOR U29276 ( .A(n28751), .B(n28750), .Z(n28744) );
  XOR U29277 ( .A(b[11]), .B(n31434), .Z(n28789) );
  OR U29278 ( .A(n28789), .B(n37311), .Z(n28634) );
  NANDN U29279 ( .A(n28632), .B(n37218), .Z(n28633) );
  NAND U29280 ( .A(n28634), .B(n28633), .Z(n28743) );
  XOR U29281 ( .A(n1053), .B(a[193]), .Z(n28792) );
  NANDN U29282 ( .A(n28792), .B(n37424), .Z(n28637) );
  NANDN U29283 ( .A(n28635), .B(n37425), .Z(n28636) );
  NAND U29284 ( .A(n28637), .B(n28636), .Z(n28742) );
  XNOR U29285 ( .A(n28743), .B(n28742), .Z(n28745) );
  XNOR U29286 ( .A(n28744), .B(n28745), .Z(n28733) );
  NANDN U29287 ( .A(n1049), .B(a[205]), .Z(n28638) );
  XNOR U29288 ( .A(b[1]), .B(n28638), .Z(n28640) );
  IV U29289 ( .A(a[204]), .Z(n33130) );
  NANDN U29290 ( .A(n33130), .B(n1049), .Z(n28639) );
  AND U29291 ( .A(n28640), .B(n28639), .Z(n28708) );
  NAND U29292 ( .A(n38490), .B(n28641), .Z(n28643) );
  XNOR U29293 ( .A(n1058), .B(a[177]), .Z(n28798) );
  NANDN U29294 ( .A(n1048), .B(n28798), .Z(n28642) );
  NAND U29295 ( .A(n28643), .B(n28642), .Z(n28706) );
  NANDN U29296 ( .A(n1059), .B(a[173]), .Z(n28707) );
  XNOR U29297 ( .A(n28706), .B(n28707), .Z(n28709) );
  XNOR U29298 ( .A(n28708), .B(n28709), .Z(n28731) );
  NANDN U29299 ( .A(n28644), .B(n38205), .Z(n28646) );
  XNOR U29300 ( .A(b[23]), .B(a[183]), .Z(n28801) );
  OR U29301 ( .A(n28801), .B(n38268), .Z(n28645) );
  NAND U29302 ( .A(n28646), .B(n28645), .Z(n28771) );
  XOR U29303 ( .A(b[7]), .B(a[199]), .Z(n28804) );
  NAND U29304 ( .A(n28804), .B(n36701), .Z(n28649) );
  NANDN U29305 ( .A(n28647), .B(n36702), .Z(n28648) );
  NAND U29306 ( .A(n28649), .B(n28648), .Z(n28768) );
  XOR U29307 ( .A(b[25]), .B(a[181]), .Z(n28807) );
  NAND U29308 ( .A(n28807), .B(n38325), .Z(n28652) );
  NAND U29309 ( .A(n28650), .B(n38326), .Z(n28651) );
  AND U29310 ( .A(n28652), .B(n28651), .Z(n28769) );
  XNOR U29311 ( .A(n28768), .B(n28769), .Z(n28770) );
  XOR U29312 ( .A(n28771), .B(n28770), .Z(n28730) );
  XOR U29313 ( .A(n28733), .B(n28732), .Z(n28761) );
  XNOR U29314 ( .A(n28760), .B(n28761), .Z(n28816) );
  XNOR U29315 ( .A(n28817), .B(n28816), .Z(n28819) );
  XNOR U29316 ( .A(n28818), .B(n28819), .Z(n28700) );
  XOR U29317 ( .A(n28701), .B(n28700), .Z(n28703) );
  NANDN U29318 ( .A(n28654), .B(n28653), .Z(n28658) );
  OR U29319 ( .A(n28656), .B(n28655), .Z(n28657) );
  NAND U29320 ( .A(n28658), .B(n28657), .Z(n28694) );
  NAND U29321 ( .A(n28660), .B(n28659), .Z(n28664) );
  NANDN U29322 ( .A(n28662), .B(n28661), .Z(n28663) );
  NAND U29323 ( .A(n28664), .B(n28663), .Z(n28695) );
  XNOR U29324 ( .A(n28694), .B(n28695), .Z(n28696) );
  XOR U29325 ( .A(n28697), .B(n28696), .Z(n28690) );
  NANDN U29326 ( .A(n28666), .B(n28665), .Z(n28670) );
  NAND U29327 ( .A(n28668), .B(n28667), .Z(n28669) );
  NAND U29328 ( .A(n28670), .B(n28669), .Z(n28688) );
  NANDN U29329 ( .A(n28672), .B(n28671), .Z(n28676) );
  OR U29330 ( .A(n28674), .B(n28673), .Z(n28675) );
  NAND U29331 ( .A(n28676), .B(n28675), .Z(n28689) );
  XNOR U29332 ( .A(n28688), .B(n28689), .Z(n28691) );
  XOR U29333 ( .A(n28690), .B(n28691), .Z(n28682) );
  XOR U29334 ( .A(n28683), .B(n28682), .Z(n28684) );
  XNOR U29335 ( .A(n28685), .B(n28684), .Z(n28822) );
  XNOR U29336 ( .A(n28822), .B(sreg[429]), .Z(n28824) );
  NAND U29337 ( .A(n28677), .B(sreg[428]), .Z(n28681) );
  OR U29338 ( .A(n28679), .B(n28678), .Z(n28680) );
  AND U29339 ( .A(n28681), .B(n28680), .Z(n28823) );
  XOR U29340 ( .A(n28824), .B(n28823), .Z(c[429]) );
  NAND U29341 ( .A(n28683), .B(n28682), .Z(n28687) );
  NAND U29342 ( .A(n28685), .B(n28684), .Z(n28686) );
  NAND U29343 ( .A(n28687), .B(n28686), .Z(n28830) );
  NANDN U29344 ( .A(n28689), .B(n28688), .Z(n28693) );
  NAND U29345 ( .A(n28691), .B(n28690), .Z(n28692) );
  NAND U29346 ( .A(n28693), .B(n28692), .Z(n28828) );
  NANDN U29347 ( .A(n28695), .B(n28694), .Z(n28699) );
  NAND U29348 ( .A(n28697), .B(n28696), .Z(n28698) );
  NAND U29349 ( .A(n28699), .B(n28698), .Z(n28833) );
  NANDN U29350 ( .A(n28701), .B(n28700), .Z(n28705) );
  OR U29351 ( .A(n28703), .B(n28702), .Z(n28704) );
  NAND U29352 ( .A(n28705), .B(n28704), .Z(n28834) );
  XNOR U29353 ( .A(n28833), .B(n28834), .Z(n28835) );
  NANDN U29354 ( .A(n28707), .B(n28706), .Z(n28711) );
  NAND U29355 ( .A(n28709), .B(n28708), .Z(n28710) );
  NAND U29356 ( .A(n28711), .B(n28710), .Z(n28852) );
  XNOR U29357 ( .A(b[19]), .B(a[188]), .Z(n28901) );
  NANDN U29358 ( .A(n28901), .B(n37934), .Z(n28714) );
  NANDN U29359 ( .A(n28712), .B(n37935), .Z(n28713) );
  NAND U29360 ( .A(n28714), .B(n28713), .Z(n28862) );
  XOR U29361 ( .A(b[27]), .B(a[180]), .Z(n28904) );
  NAND U29362 ( .A(n38423), .B(n28904), .Z(n28717) );
  NAND U29363 ( .A(n28715), .B(n38424), .Z(n28716) );
  NAND U29364 ( .A(n28717), .B(n28716), .Z(n28859) );
  XNOR U29365 ( .A(b[5]), .B(a[202]), .Z(n28907) );
  NANDN U29366 ( .A(n28907), .B(n36587), .Z(n28720) );
  NANDN U29367 ( .A(n28718), .B(n36588), .Z(n28719) );
  AND U29368 ( .A(n28720), .B(n28719), .Z(n28860) );
  XNOR U29369 ( .A(n28859), .B(n28860), .Z(n28861) );
  XNOR U29370 ( .A(n28862), .B(n28861), .Z(n28850) );
  NANDN U29371 ( .A(n28721), .B(n37762), .Z(n28723) );
  XOR U29372 ( .A(b[17]), .B(a[190]), .Z(n28910) );
  NAND U29373 ( .A(n28910), .B(n37764), .Z(n28722) );
  NAND U29374 ( .A(n28723), .B(n28722), .Z(n28928) );
  XNOR U29375 ( .A(b[31]), .B(a[176]), .Z(n28913) );
  NANDN U29376 ( .A(n28913), .B(n38552), .Z(n28726) );
  NANDN U29377 ( .A(n28724), .B(n38553), .Z(n28725) );
  NAND U29378 ( .A(n28726), .B(n28725), .Z(n28925) );
  OR U29379 ( .A(n28727), .B(n36105), .Z(n28729) );
  XOR U29380 ( .A(b[3]), .B(n33130), .Z(n28916) );
  NANDN U29381 ( .A(n28916), .B(n36107), .Z(n28728) );
  AND U29382 ( .A(n28729), .B(n28728), .Z(n28926) );
  XNOR U29383 ( .A(n28925), .B(n28926), .Z(n28927) );
  XOR U29384 ( .A(n28928), .B(n28927), .Z(n28849) );
  XNOR U29385 ( .A(n28850), .B(n28849), .Z(n28851) );
  XNOR U29386 ( .A(n28852), .B(n28851), .Z(n28949) );
  NANDN U29387 ( .A(n28731), .B(n28730), .Z(n28735) );
  NANDN U29388 ( .A(n28733), .B(n28732), .Z(n28734) );
  NAND U29389 ( .A(n28735), .B(n28734), .Z(n28950) );
  XNOR U29390 ( .A(n28949), .B(n28950), .Z(n28951) );
  NANDN U29391 ( .A(n28737), .B(n28736), .Z(n28741) );
  NAND U29392 ( .A(n28739), .B(n28738), .Z(n28740) );
  NAND U29393 ( .A(n28741), .B(n28740), .Z(n28842) );
  OR U29394 ( .A(n28743), .B(n28742), .Z(n28747) );
  NANDN U29395 ( .A(n28745), .B(n28744), .Z(n28746) );
  NAND U29396 ( .A(n28747), .B(n28746), .Z(n28840) );
  XNOR U29397 ( .A(n28840), .B(n28839), .Z(n28841) );
  XOR U29398 ( .A(n28842), .B(n28841), .Z(n28952) );
  XOR U29399 ( .A(n28951), .B(n28952), .Z(n28962) );
  OR U29400 ( .A(n28753), .B(n28752), .Z(n28757) );
  NAND U29401 ( .A(n28755), .B(n28754), .Z(n28756) );
  NAND U29402 ( .A(n28757), .B(n28756), .Z(n28960) );
  NANDN U29403 ( .A(n28759), .B(n28758), .Z(n28763) );
  NANDN U29404 ( .A(n28761), .B(n28760), .Z(n28762) );
  NAND U29405 ( .A(n28763), .B(n28762), .Z(n28945) );
  NANDN U29406 ( .A(n28769), .B(n28768), .Z(n28773) );
  NAND U29407 ( .A(n28771), .B(n28770), .Z(n28772) );
  NAND U29408 ( .A(n28773), .B(n28772), .Z(n28843) );
  NANDN U29409 ( .A(n28775), .B(n28774), .Z(n28779) );
  NAND U29410 ( .A(n28777), .B(n28776), .Z(n28778) );
  AND U29411 ( .A(n28779), .B(n28778), .Z(n28844) );
  XNOR U29412 ( .A(n28843), .B(n28844), .Z(n28845) );
  XOR U29413 ( .A(b[9]), .B(n32246), .Z(n28865) );
  NANDN U29414 ( .A(n28865), .B(n36925), .Z(n28782) );
  NANDN U29415 ( .A(n28780), .B(n36926), .Z(n28781) );
  NAND U29416 ( .A(n28782), .B(n28781), .Z(n28939) );
  XNOR U29417 ( .A(b[15]), .B(a[192]), .Z(n28868) );
  OR U29418 ( .A(n28868), .B(n37665), .Z(n28785) );
  NANDN U29419 ( .A(n28783), .B(n37604), .Z(n28784) );
  AND U29420 ( .A(n28785), .B(n28784), .Z(n28937) );
  XNOR U29421 ( .A(b[21]), .B(a[186]), .Z(n28871) );
  NANDN U29422 ( .A(n28871), .B(n38101), .Z(n28788) );
  NANDN U29423 ( .A(n28786), .B(n38102), .Z(n28787) );
  AND U29424 ( .A(n28788), .B(n28787), .Z(n28938) );
  XOR U29425 ( .A(n28939), .B(n28940), .Z(n28934) );
  XNOR U29426 ( .A(b[11]), .B(a[196]), .Z(n28874) );
  OR U29427 ( .A(n28874), .B(n37311), .Z(n28791) );
  NANDN U29428 ( .A(n28789), .B(n37218), .Z(n28790) );
  NAND U29429 ( .A(n28791), .B(n28790), .Z(n28932) );
  XOR U29430 ( .A(n1053), .B(a[194]), .Z(n28877) );
  NANDN U29431 ( .A(n28877), .B(n37424), .Z(n28794) );
  NANDN U29432 ( .A(n28792), .B(n37425), .Z(n28793) );
  AND U29433 ( .A(n28794), .B(n28793), .Z(n28931) );
  XNOR U29434 ( .A(n28932), .B(n28931), .Z(n28933) );
  XOR U29435 ( .A(n28934), .B(n28933), .Z(n28921) );
  NANDN U29436 ( .A(n1049), .B(a[206]), .Z(n28795) );
  XNOR U29437 ( .A(b[1]), .B(n28795), .Z(n28797) );
  NANDN U29438 ( .A(b[0]), .B(a[205]), .Z(n28796) );
  AND U29439 ( .A(n28797), .B(n28796), .Z(n28897) );
  NAND U29440 ( .A(n38490), .B(n28798), .Z(n28800) );
  XNOR U29441 ( .A(n1058), .B(a[178]), .Z(n28883) );
  NANDN U29442 ( .A(n1048), .B(n28883), .Z(n28799) );
  NAND U29443 ( .A(n28800), .B(n28799), .Z(n28895) );
  NANDN U29444 ( .A(n1059), .B(a[174]), .Z(n28896) );
  XNOR U29445 ( .A(n28895), .B(n28896), .Z(n28898) );
  XOR U29446 ( .A(n28897), .B(n28898), .Z(n28919) );
  NANDN U29447 ( .A(n28801), .B(n38205), .Z(n28803) );
  XNOR U29448 ( .A(b[23]), .B(a[184]), .Z(n28886) );
  OR U29449 ( .A(n28886), .B(n38268), .Z(n28802) );
  NAND U29450 ( .A(n28803), .B(n28802), .Z(n28856) );
  XOR U29451 ( .A(b[7]), .B(a[200]), .Z(n28889) );
  NAND U29452 ( .A(n28889), .B(n36701), .Z(n28806) );
  NAND U29453 ( .A(n28804), .B(n36702), .Z(n28805) );
  NAND U29454 ( .A(n28806), .B(n28805), .Z(n28853) );
  XOR U29455 ( .A(b[25]), .B(a[182]), .Z(n28892) );
  NAND U29456 ( .A(n28892), .B(n38325), .Z(n28809) );
  NAND U29457 ( .A(n28807), .B(n38326), .Z(n28808) );
  AND U29458 ( .A(n28809), .B(n28808), .Z(n28854) );
  XNOR U29459 ( .A(n28853), .B(n28854), .Z(n28855) );
  XNOR U29460 ( .A(n28856), .B(n28855), .Z(n28920) );
  XOR U29461 ( .A(n28919), .B(n28920), .Z(n28922) );
  XNOR U29462 ( .A(n28921), .B(n28922), .Z(n28846) );
  XNOR U29463 ( .A(n28845), .B(n28846), .Z(n28943) );
  XNOR U29464 ( .A(n28944), .B(n28943), .Z(n28946) );
  XNOR U29465 ( .A(n28945), .B(n28946), .Z(n28959) );
  XOR U29466 ( .A(n28960), .B(n28959), .Z(n28961) );
  XNOR U29467 ( .A(n28962), .B(n28961), .Z(n28956) );
  NANDN U29468 ( .A(n28811), .B(n28810), .Z(n28815) );
  OR U29469 ( .A(n28813), .B(n28812), .Z(n28814) );
  NAND U29470 ( .A(n28815), .B(n28814), .Z(n28953) );
  NAND U29471 ( .A(n28817), .B(n28816), .Z(n28821) );
  NANDN U29472 ( .A(n28819), .B(n28818), .Z(n28820) );
  NAND U29473 ( .A(n28821), .B(n28820), .Z(n28954) );
  XNOR U29474 ( .A(n28953), .B(n28954), .Z(n28955) );
  XOR U29475 ( .A(n28956), .B(n28955), .Z(n28836) );
  XOR U29476 ( .A(n28835), .B(n28836), .Z(n28827) );
  XOR U29477 ( .A(n28828), .B(n28827), .Z(n28829) );
  XNOR U29478 ( .A(n28830), .B(n28829), .Z(n28965) );
  XNOR U29479 ( .A(n28965), .B(sreg[430]), .Z(n28967) );
  NAND U29480 ( .A(n28822), .B(sreg[429]), .Z(n28826) );
  OR U29481 ( .A(n28824), .B(n28823), .Z(n28825) );
  AND U29482 ( .A(n28826), .B(n28825), .Z(n28966) );
  XOR U29483 ( .A(n28967), .B(n28966), .Z(c[430]) );
  NAND U29484 ( .A(n28828), .B(n28827), .Z(n28832) );
  NAND U29485 ( .A(n28830), .B(n28829), .Z(n28831) );
  NAND U29486 ( .A(n28832), .B(n28831), .Z(n28973) );
  NANDN U29487 ( .A(n28834), .B(n28833), .Z(n28838) );
  NAND U29488 ( .A(n28836), .B(n28835), .Z(n28837) );
  NAND U29489 ( .A(n28838), .B(n28837), .Z(n28971) );
  NANDN U29490 ( .A(n28844), .B(n28843), .Z(n28848) );
  NANDN U29491 ( .A(n28846), .B(n28845), .Z(n28847) );
  NAND U29492 ( .A(n28848), .B(n28847), .Z(n28987) );
  NANDN U29493 ( .A(n28854), .B(n28853), .Z(n28858) );
  NAND U29494 ( .A(n28856), .B(n28855), .Z(n28857) );
  NAND U29495 ( .A(n28858), .B(n28857), .Z(n29044) );
  NANDN U29496 ( .A(n28860), .B(n28859), .Z(n28864) );
  NAND U29497 ( .A(n28862), .B(n28861), .Z(n28863) );
  AND U29498 ( .A(n28864), .B(n28863), .Z(n29045) );
  XNOR U29499 ( .A(n29044), .B(n29045), .Z(n29046) );
  XNOR U29500 ( .A(n1052), .B(a[199]), .Z(n29068) );
  NAND U29501 ( .A(n36925), .B(n29068), .Z(n28867) );
  NANDN U29502 ( .A(n28865), .B(n36926), .Z(n28866) );
  NAND U29503 ( .A(n28867), .B(n28866), .Z(n29010) );
  XOR U29504 ( .A(b[15]), .B(n31508), .Z(n29071) );
  OR U29505 ( .A(n29071), .B(n37665), .Z(n28870) );
  NANDN U29506 ( .A(n28868), .B(n37604), .Z(n28869) );
  AND U29507 ( .A(n28870), .B(n28869), .Z(n29008) );
  XNOR U29508 ( .A(n1056), .B(a[187]), .Z(n29074) );
  NAND U29509 ( .A(n29074), .B(n38101), .Z(n28873) );
  NANDN U29510 ( .A(n28871), .B(n38102), .Z(n28872) );
  AND U29511 ( .A(n28873), .B(n28872), .Z(n29009) );
  XOR U29512 ( .A(n29010), .B(n29011), .Z(n28999) );
  XNOR U29513 ( .A(b[11]), .B(a[197]), .Z(n29077) );
  OR U29514 ( .A(n29077), .B(n37311), .Z(n28876) );
  NANDN U29515 ( .A(n28874), .B(n37218), .Z(n28875) );
  NAND U29516 ( .A(n28876), .B(n28875), .Z(n28997) );
  XOR U29517 ( .A(n1053), .B(a[195]), .Z(n29080) );
  NANDN U29518 ( .A(n29080), .B(n37424), .Z(n28879) );
  NANDN U29519 ( .A(n28877), .B(n37425), .Z(n28878) );
  NAND U29520 ( .A(n28879), .B(n28878), .Z(n28996) );
  XOR U29521 ( .A(n28999), .B(n28998), .Z(n28993) );
  NANDN U29522 ( .A(n1049), .B(a[207]), .Z(n28880) );
  XNOR U29523 ( .A(b[1]), .B(n28880), .Z(n28882) );
  NANDN U29524 ( .A(b[0]), .B(a[206]), .Z(n28881) );
  AND U29525 ( .A(n28882), .B(n28881), .Z(n29016) );
  NAND U29526 ( .A(n38490), .B(n28883), .Z(n28885) );
  XNOR U29527 ( .A(n1058), .B(a[179]), .Z(n29086) );
  NANDN U29528 ( .A(n1048), .B(n29086), .Z(n28884) );
  NAND U29529 ( .A(n28885), .B(n28884), .Z(n29014) );
  NANDN U29530 ( .A(n1059), .B(a[175]), .Z(n29015) );
  XNOR U29531 ( .A(n29014), .B(n29015), .Z(n29017) );
  XNOR U29532 ( .A(n29016), .B(n29017), .Z(n28991) );
  NANDN U29533 ( .A(n28886), .B(n38205), .Z(n28888) );
  XNOR U29534 ( .A(b[23]), .B(a[185]), .Z(n29089) );
  OR U29535 ( .A(n29089), .B(n38268), .Z(n28887) );
  NAND U29536 ( .A(n28888), .B(n28887), .Z(n29059) );
  XNOR U29537 ( .A(b[7]), .B(a[201]), .Z(n29092) );
  NANDN U29538 ( .A(n29092), .B(n36701), .Z(n28891) );
  NAND U29539 ( .A(n28889), .B(n36702), .Z(n28890) );
  NAND U29540 ( .A(n28891), .B(n28890), .Z(n29056) );
  XOR U29541 ( .A(b[25]), .B(a[183]), .Z(n29095) );
  NAND U29542 ( .A(n29095), .B(n38325), .Z(n28894) );
  NAND U29543 ( .A(n28892), .B(n38326), .Z(n28893) );
  AND U29544 ( .A(n28894), .B(n28893), .Z(n29057) );
  XNOR U29545 ( .A(n29056), .B(n29057), .Z(n29058) );
  XOR U29546 ( .A(n29059), .B(n29058), .Z(n28990) );
  XOR U29547 ( .A(n28993), .B(n28992), .Z(n29047) );
  XNOR U29548 ( .A(n29046), .B(n29047), .Z(n28984) );
  XOR U29549 ( .A(n28985), .B(n28984), .Z(n28986) );
  XOR U29550 ( .A(n28987), .B(n28986), .Z(n29099) );
  XNOR U29551 ( .A(n29098), .B(n29099), .Z(n29101) );
  NANDN U29552 ( .A(n28896), .B(n28895), .Z(n28900) );
  NAND U29553 ( .A(n28898), .B(n28897), .Z(n28899) );
  NAND U29554 ( .A(n28900), .B(n28899), .Z(n29053) );
  XOR U29555 ( .A(b[19]), .B(n30936), .Z(n29020) );
  NANDN U29556 ( .A(n29020), .B(n37934), .Z(n28903) );
  NANDN U29557 ( .A(n28901), .B(n37935), .Z(n28902) );
  NAND U29558 ( .A(n28903), .B(n28902), .Z(n29065) );
  XOR U29559 ( .A(b[27]), .B(a[181]), .Z(n29023) );
  NAND U29560 ( .A(n38423), .B(n29023), .Z(n28906) );
  NAND U29561 ( .A(n28904), .B(n38424), .Z(n28905) );
  NAND U29562 ( .A(n28906), .B(n28905), .Z(n29062) );
  XNOR U29563 ( .A(b[5]), .B(a[203]), .Z(n29026) );
  NANDN U29564 ( .A(n29026), .B(n36587), .Z(n28909) );
  NANDN U29565 ( .A(n28907), .B(n36588), .Z(n28908) );
  AND U29566 ( .A(n28909), .B(n28908), .Z(n29063) );
  XNOR U29567 ( .A(n29062), .B(n29063), .Z(n29064) );
  XNOR U29568 ( .A(n29065), .B(n29064), .Z(n29050) );
  NAND U29569 ( .A(n28910), .B(n37762), .Z(n28912) );
  XOR U29570 ( .A(b[17]), .B(a[191]), .Z(n29029) );
  NAND U29571 ( .A(n29029), .B(n37764), .Z(n28911) );
  NAND U29572 ( .A(n28912), .B(n28911), .Z(n29004) );
  XNOR U29573 ( .A(b[31]), .B(a[177]), .Z(n29032) );
  NANDN U29574 ( .A(n29032), .B(n38552), .Z(n28915) );
  NANDN U29575 ( .A(n28913), .B(n38553), .Z(n28914) );
  AND U29576 ( .A(n28915), .B(n28914), .Z(n29002) );
  OR U29577 ( .A(n28916), .B(n36105), .Z(n28918) );
  XNOR U29578 ( .A(b[3]), .B(a[205]), .Z(n29035) );
  NANDN U29579 ( .A(n29035), .B(n36107), .Z(n28917) );
  AND U29580 ( .A(n28918), .B(n28917), .Z(n29003) );
  XOR U29581 ( .A(n29004), .B(n29005), .Z(n29051) );
  XOR U29582 ( .A(n29050), .B(n29051), .Z(n29052) );
  XNOR U29583 ( .A(n29053), .B(n29052), .Z(n28980) );
  NANDN U29584 ( .A(n28920), .B(n28919), .Z(n28924) );
  OR U29585 ( .A(n28922), .B(n28921), .Z(n28923) );
  NAND U29586 ( .A(n28924), .B(n28923), .Z(n28981) );
  XNOR U29587 ( .A(n28980), .B(n28981), .Z(n28982) );
  NANDN U29588 ( .A(n28926), .B(n28925), .Z(n28930) );
  NAND U29589 ( .A(n28928), .B(n28927), .Z(n28929) );
  NAND U29590 ( .A(n28930), .B(n28929), .Z(n29041) );
  NANDN U29591 ( .A(n28932), .B(n28931), .Z(n28936) );
  NAND U29592 ( .A(n28934), .B(n28933), .Z(n28935) );
  NAND U29593 ( .A(n28936), .B(n28935), .Z(n29038) );
  OR U29594 ( .A(n28938), .B(n28937), .Z(n28942) );
  NANDN U29595 ( .A(n28940), .B(n28939), .Z(n28941) );
  NAND U29596 ( .A(n28942), .B(n28941), .Z(n29039) );
  XNOR U29597 ( .A(n29038), .B(n29039), .Z(n29040) );
  XOR U29598 ( .A(n29041), .B(n29040), .Z(n28983) );
  XNOR U29599 ( .A(n28982), .B(n28983), .Z(n29100) );
  XOR U29600 ( .A(n29101), .B(n29100), .Z(n29105) );
  NAND U29601 ( .A(n28944), .B(n28943), .Z(n28948) );
  NANDN U29602 ( .A(n28946), .B(n28945), .Z(n28947) );
  NAND U29603 ( .A(n28948), .B(n28947), .Z(n29102) );
  XNOR U29604 ( .A(n29102), .B(n29103), .Z(n29104) );
  XNOR U29605 ( .A(n29105), .B(n29104), .Z(n28977) );
  NANDN U29606 ( .A(n28954), .B(n28953), .Z(n28958) );
  NAND U29607 ( .A(n28956), .B(n28955), .Z(n28957) );
  NAND U29608 ( .A(n28958), .B(n28957), .Z(n28974) );
  NANDN U29609 ( .A(n28960), .B(n28959), .Z(n28964) );
  OR U29610 ( .A(n28962), .B(n28961), .Z(n28963) );
  NAND U29611 ( .A(n28964), .B(n28963), .Z(n28975) );
  XNOR U29612 ( .A(n28974), .B(n28975), .Z(n28976) );
  XNOR U29613 ( .A(n28977), .B(n28976), .Z(n28970) );
  XOR U29614 ( .A(n28971), .B(n28970), .Z(n28972) );
  XNOR U29615 ( .A(n28973), .B(n28972), .Z(n29108) );
  XNOR U29616 ( .A(n29108), .B(sreg[431]), .Z(n29110) );
  NAND U29617 ( .A(n28965), .B(sreg[430]), .Z(n28969) );
  OR U29618 ( .A(n28967), .B(n28966), .Z(n28968) );
  AND U29619 ( .A(n28969), .B(n28968), .Z(n29109) );
  XOR U29620 ( .A(n29110), .B(n29109), .Z(c[431]) );
  NANDN U29621 ( .A(n28975), .B(n28974), .Z(n28979) );
  NANDN U29622 ( .A(n28977), .B(n28976), .Z(n28978) );
  NAND U29623 ( .A(n28979), .B(n28978), .Z(n29114) );
  NAND U29624 ( .A(n28985), .B(n28984), .Z(n28989) );
  NAND U29625 ( .A(n28987), .B(n28986), .Z(n28988) );
  NAND U29626 ( .A(n28989), .B(n28988), .Z(n29248) );
  XNOR U29627 ( .A(n29247), .B(n29248), .Z(n29249) );
  NANDN U29628 ( .A(n28991), .B(n28990), .Z(n28995) );
  NANDN U29629 ( .A(n28993), .B(n28992), .Z(n28994) );
  NAND U29630 ( .A(n28995), .B(n28994), .Z(n29234) );
  OR U29631 ( .A(n28997), .B(n28996), .Z(n29001) );
  NAND U29632 ( .A(n28999), .B(n28998), .Z(n29000) );
  NAND U29633 ( .A(n29001), .B(n29000), .Z(n29173) );
  OR U29634 ( .A(n29003), .B(n29002), .Z(n29007) );
  NANDN U29635 ( .A(n29005), .B(n29004), .Z(n29006) );
  NAND U29636 ( .A(n29007), .B(n29006), .Z(n29172) );
  OR U29637 ( .A(n29009), .B(n29008), .Z(n29013) );
  NANDN U29638 ( .A(n29011), .B(n29010), .Z(n29012) );
  NAND U29639 ( .A(n29013), .B(n29012), .Z(n29171) );
  XOR U29640 ( .A(n29173), .B(n29174), .Z(n29231) );
  NANDN U29641 ( .A(n29015), .B(n29014), .Z(n29019) );
  NAND U29642 ( .A(n29017), .B(n29016), .Z(n29018) );
  NAND U29643 ( .A(n29019), .B(n29018), .Z(n29186) );
  XNOR U29644 ( .A(b[19]), .B(a[190]), .Z(n29131) );
  NANDN U29645 ( .A(n29131), .B(n37934), .Z(n29022) );
  NANDN U29646 ( .A(n29020), .B(n37935), .Z(n29021) );
  NAND U29647 ( .A(n29022), .B(n29021), .Z(n29198) );
  XOR U29648 ( .A(b[27]), .B(a[182]), .Z(n29134) );
  NAND U29649 ( .A(n38423), .B(n29134), .Z(n29025) );
  NAND U29650 ( .A(n29023), .B(n38424), .Z(n29024) );
  NAND U29651 ( .A(n29025), .B(n29024), .Z(n29195) );
  XOR U29652 ( .A(b[5]), .B(n33130), .Z(n29137) );
  NANDN U29653 ( .A(n29137), .B(n36587), .Z(n29028) );
  NANDN U29654 ( .A(n29026), .B(n36588), .Z(n29027) );
  AND U29655 ( .A(n29028), .B(n29027), .Z(n29196) );
  XNOR U29656 ( .A(n29195), .B(n29196), .Z(n29197) );
  XNOR U29657 ( .A(n29198), .B(n29197), .Z(n29184) );
  NAND U29658 ( .A(n29029), .B(n37762), .Z(n29031) );
  XOR U29659 ( .A(b[17]), .B(a[192]), .Z(n29140) );
  NAND U29660 ( .A(n29140), .B(n37764), .Z(n29030) );
  NAND U29661 ( .A(n29031), .B(n29030), .Z(n29158) );
  XNOR U29662 ( .A(b[31]), .B(a[178]), .Z(n29143) );
  NANDN U29663 ( .A(n29143), .B(n38552), .Z(n29034) );
  NANDN U29664 ( .A(n29032), .B(n38553), .Z(n29033) );
  NAND U29665 ( .A(n29034), .B(n29033), .Z(n29155) );
  OR U29666 ( .A(n29035), .B(n36105), .Z(n29037) );
  XNOR U29667 ( .A(b[3]), .B(a[206]), .Z(n29146) );
  NANDN U29668 ( .A(n29146), .B(n36107), .Z(n29036) );
  AND U29669 ( .A(n29037), .B(n29036), .Z(n29156) );
  XNOR U29670 ( .A(n29155), .B(n29156), .Z(n29157) );
  XOR U29671 ( .A(n29158), .B(n29157), .Z(n29183) );
  XNOR U29672 ( .A(n29184), .B(n29183), .Z(n29185) );
  XNOR U29673 ( .A(n29186), .B(n29185), .Z(n29232) );
  XNOR U29674 ( .A(n29231), .B(n29232), .Z(n29233) );
  XNOR U29675 ( .A(n29234), .B(n29233), .Z(n29244) );
  NANDN U29676 ( .A(n29039), .B(n29038), .Z(n29043) );
  NANDN U29677 ( .A(n29041), .B(n29040), .Z(n29042) );
  NAND U29678 ( .A(n29043), .B(n29042), .Z(n29241) );
  NANDN U29679 ( .A(n29045), .B(n29044), .Z(n29049) );
  NANDN U29680 ( .A(n29047), .B(n29046), .Z(n29048) );
  NAND U29681 ( .A(n29049), .B(n29048), .Z(n29238) );
  OR U29682 ( .A(n29051), .B(n29050), .Z(n29055) );
  NAND U29683 ( .A(n29053), .B(n29052), .Z(n29054) );
  NAND U29684 ( .A(n29055), .B(n29054), .Z(n29236) );
  NANDN U29685 ( .A(n29057), .B(n29056), .Z(n29061) );
  NAND U29686 ( .A(n29059), .B(n29058), .Z(n29060) );
  NAND U29687 ( .A(n29061), .B(n29060), .Z(n29177) );
  NANDN U29688 ( .A(n29063), .B(n29062), .Z(n29067) );
  NAND U29689 ( .A(n29065), .B(n29064), .Z(n29066) );
  AND U29690 ( .A(n29067), .B(n29066), .Z(n29178) );
  XNOR U29691 ( .A(n29177), .B(n29178), .Z(n29179) );
  XOR U29692 ( .A(n1052), .B(a[200]), .Z(n29207) );
  NANDN U29693 ( .A(n29207), .B(n36925), .Z(n29070) );
  NAND U29694 ( .A(n36926), .B(n29068), .Z(n29069) );
  NAND U29695 ( .A(n29070), .B(n29069), .Z(n29163) );
  XNOR U29696 ( .A(n1054), .B(a[194]), .Z(n29204) );
  NANDN U29697 ( .A(n37665), .B(n29204), .Z(n29073) );
  NANDN U29698 ( .A(n29071), .B(n37604), .Z(n29072) );
  NAND U29699 ( .A(n29073), .B(n29072), .Z(n29161) );
  XOR U29700 ( .A(n1056), .B(a[188]), .Z(n29201) );
  NANDN U29701 ( .A(n29201), .B(n38101), .Z(n29076) );
  NAND U29702 ( .A(n38102), .B(n29074), .Z(n29075) );
  NAND U29703 ( .A(n29076), .B(n29075), .Z(n29162) );
  XNOR U29704 ( .A(n29161), .B(n29162), .Z(n29164) );
  XOR U29705 ( .A(n29163), .B(n29164), .Z(n29152) );
  XOR U29706 ( .A(b[11]), .B(n32246), .Z(n29210) );
  OR U29707 ( .A(n29210), .B(n37311), .Z(n29079) );
  NANDN U29708 ( .A(n29077), .B(n37218), .Z(n29078) );
  NAND U29709 ( .A(n29079), .B(n29078), .Z(n29150) );
  XOR U29710 ( .A(n1053), .B(a[196]), .Z(n29213) );
  NANDN U29711 ( .A(n29213), .B(n37424), .Z(n29082) );
  NANDN U29712 ( .A(n29080), .B(n37425), .Z(n29081) );
  AND U29713 ( .A(n29082), .B(n29081), .Z(n29149) );
  XNOR U29714 ( .A(n29150), .B(n29149), .Z(n29151) );
  XNOR U29715 ( .A(n29152), .B(n29151), .Z(n29168) );
  NANDN U29716 ( .A(n1049), .B(a[208]), .Z(n29083) );
  XNOR U29717 ( .A(b[1]), .B(n29083), .Z(n29085) );
  NANDN U29718 ( .A(b[0]), .B(a[207]), .Z(n29084) );
  AND U29719 ( .A(n29085), .B(n29084), .Z(n29127) );
  NAND U29720 ( .A(n38490), .B(n29086), .Z(n29088) );
  XNOR U29721 ( .A(n1058), .B(a[180]), .Z(n29219) );
  NANDN U29722 ( .A(n1048), .B(n29219), .Z(n29087) );
  NAND U29723 ( .A(n29088), .B(n29087), .Z(n29125) );
  NANDN U29724 ( .A(n1059), .B(a[176]), .Z(n29126) );
  XNOR U29725 ( .A(n29125), .B(n29126), .Z(n29128) );
  XNOR U29726 ( .A(n29127), .B(n29128), .Z(n29166) );
  NANDN U29727 ( .A(n29089), .B(n38205), .Z(n29091) );
  XNOR U29728 ( .A(b[23]), .B(a[186]), .Z(n29222) );
  OR U29729 ( .A(n29222), .B(n38268), .Z(n29090) );
  NAND U29730 ( .A(n29091), .B(n29090), .Z(n29192) );
  XOR U29731 ( .A(b[7]), .B(a[202]), .Z(n29225) );
  NAND U29732 ( .A(n29225), .B(n36701), .Z(n29094) );
  NANDN U29733 ( .A(n29092), .B(n36702), .Z(n29093) );
  NAND U29734 ( .A(n29094), .B(n29093), .Z(n29189) );
  XOR U29735 ( .A(b[25]), .B(a[184]), .Z(n29228) );
  NAND U29736 ( .A(n29228), .B(n38325), .Z(n29097) );
  NAND U29737 ( .A(n29095), .B(n38326), .Z(n29096) );
  AND U29738 ( .A(n29097), .B(n29096), .Z(n29190) );
  XNOR U29739 ( .A(n29189), .B(n29190), .Z(n29191) );
  XOR U29740 ( .A(n29192), .B(n29191), .Z(n29165) );
  XOR U29741 ( .A(n29168), .B(n29167), .Z(n29180) );
  XOR U29742 ( .A(n29179), .B(n29180), .Z(n29235) );
  XOR U29743 ( .A(n29236), .B(n29235), .Z(n29237) );
  XOR U29744 ( .A(n29238), .B(n29237), .Z(n29242) );
  XNOR U29745 ( .A(n29241), .B(n29242), .Z(n29243) );
  XOR U29746 ( .A(n29244), .B(n29243), .Z(n29250) );
  XOR U29747 ( .A(n29249), .B(n29250), .Z(n29121) );
  NANDN U29748 ( .A(n29103), .B(n29102), .Z(n29107) );
  NANDN U29749 ( .A(n29105), .B(n29104), .Z(n29106) );
  NAND U29750 ( .A(n29107), .B(n29106), .Z(n29120) );
  XNOR U29751 ( .A(n29119), .B(n29120), .Z(n29122) );
  XOR U29752 ( .A(n29121), .B(n29122), .Z(n29113) );
  XOR U29753 ( .A(n29114), .B(n29113), .Z(n29115) );
  XNOR U29754 ( .A(n29116), .B(n29115), .Z(n29253) );
  XNOR U29755 ( .A(n29253), .B(sreg[432]), .Z(n29255) );
  NAND U29756 ( .A(n29108), .B(sreg[431]), .Z(n29112) );
  OR U29757 ( .A(n29110), .B(n29109), .Z(n29111) );
  AND U29758 ( .A(n29112), .B(n29111), .Z(n29254) );
  XOR U29759 ( .A(n29255), .B(n29254), .Z(c[432]) );
  NAND U29760 ( .A(n29114), .B(n29113), .Z(n29118) );
  NAND U29761 ( .A(n29116), .B(n29115), .Z(n29117) );
  NAND U29762 ( .A(n29118), .B(n29117), .Z(n29261) );
  NANDN U29763 ( .A(n29120), .B(n29119), .Z(n29124) );
  NAND U29764 ( .A(n29122), .B(n29121), .Z(n29123) );
  NAND U29765 ( .A(n29124), .B(n29123), .Z(n29259) );
  NANDN U29766 ( .A(n29126), .B(n29125), .Z(n29130) );
  NAND U29767 ( .A(n29128), .B(n29127), .Z(n29129) );
  NAND U29768 ( .A(n29130), .B(n29129), .Z(n29339) );
  XNOR U29769 ( .A(b[19]), .B(a[191]), .Z(n29286) );
  NANDN U29770 ( .A(n29286), .B(n37934), .Z(n29133) );
  NANDN U29771 ( .A(n29131), .B(n37935), .Z(n29132) );
  NAND U29772 ( .A(n29133), .B(n29132), .Z(n29373) );
  XOR U29773 ( .A(b[27]), .B(a[183]), .Z(n29289) );
  NAND U29774 ( .A(n38423), .B(n29289), .Z(n29136) );
  NAND U29775 ( .A(n29134), .B(n38424), .Z(n29135) );
  NAND U29776 ( .A(n29136), .B(n29135), .Z(n29370) );
  XNOR U29777 ( .A(b[5]), .B(a[205]), .Z(n29292) );
  NANDN U29778 ( .A(n29292), .B(n36587), .Z(n29139) );
  NANDN U29779 ( .A(n29137), .B(n36588), .Z(n29138) );
  AND U29780 ( .A(n29139), .B(n29138), .Z(n29371) );
  XNOR U29781 ( .A(n29370), .B(n29371), .Z(n29372) );
  XNOR U29782 ( .A(n29373), .B(n29372), .Z(n29337) );
  NAND U29783 ( .A(n29140), .B(n37762), .Z(n29142) );
  XNOR U29784 ( .A(b[17]), .B(a[193]), .Z(n29295) );
  NANDN U29785 ( .A(n29295), .B(n37764), .Z(n29141) );
  NAND U29786 ( .A(n29142), .B(n29141), .Z(n29313) );
  XNOR U29787 ( .A(b[31]), .B(a[179]), .Z(n29298) );
  NANDN U29788 ( .A(n29298), .B(n38552), .Z(n29145) );
  NANDN U29789 ( .A(n29143), .B(n38553), .Z(n29144) );
  NAND U29790 ( .A(n29145), .B(n29144), .Z(n29310) );
  OR U29791 ( .A(n29146), .B(n36105), .Z(n29148) );
  XNOR U29792 ( .A(b[3]), .B(a[207]), .Z(n29301) );
  NANDN U29793 ( .A(n29301), .B(n36107), .Z(n29147) );
  AND U29794 ( .A(n29148), .B(n29147), .Z(n29311) );
  XNOR U29795 ( .A(n29310), .B(n29311), .Z(n29312) );
  XOR U29796 ( .A(n29313), .B(n29312), .Z(n29336) );
  XNOR U29797 ( .A(n29337), .B(n29336), .Z(n29338) );
  XNOR U29798 ( .A(n29339), .B(n29338), .Z(n29277) );
  NANDN U29799 ( .A(n29150), .B(n29149), .Z(n29154) );
  NAND U29800 ( .A(n29152), .B(n29151), .Z(n29153) );
  NAND U29801 ( .A(n29154), .B(n29153), .Z(n29328) );
  NANDN U29802 ( .A(n29156), .B(n29155), .Z(n29160) );
  NAND U29803 ( .A(n29158), .B(n29157), .Z(n29159) );
  NAND U29804 ( .A(n29160), .B(n29159), .Z(n29327) );
  XNOR U29805 ( .A(n29327), .B(n29326), .Z(n29329) );
  XOR U29806 ( .A(n29328), .B(n29329), .Z(n29276) );
  XOR U29807 ( .A(n29277), .B(n29276), .Z(n29278) );
  NANDN U29808 ( .A(n29166), .B(n29165), .Z(n29170) );
  NAND U29809 ( .A(n29168), .B(n29167), .Z(n29169) );
  NAND U29810 ( .A(n29170), .B(n29169), .Z(n29279) );
  XNOR U29811 ( .A(n29278), .B(n29279), .Z(n29390) );
  OR U29812 ( .A(n29172), .B(n29171), .Z(n29176) );
  NANDN U29813 ( .A(n29174), .B(n29173), .Z(n29175) );
  NAND U29814 ( .A(n29176), .B(n29175), .Z(n29389) );
  NANDN U29815 ( .A(n29178), .B(n29177), .Z(n29182) );
  NAND U29816 ( .A(n29180), .B(n29179), .Z(n29181) );
  NAND U29817 ( .A(n29182), .B(n29181), .Z(n29272) );
  NANDN U29818 ( .A(n29184), .B(n29183), .Z(n29188) );
  NAND U29819 ( .A(n29186), .B(n29185), .Z(n29187) );
  NAND U29820 ( .A(n29188), .B(n29187), .Z(n29271) );
  NANDN U29821 ( .A(n29190), .B(n29189), .Z(n29194) );
  NAND U29822 ( .A(n29192), .B(n29191), .Z(n29193) );
  NAND U29823 ( .A(n29194), .B(n29193), .Z(n29330) );
  NANDN U29824 ( .A(n29196), .B(n29195), .Z(n29200) );
  NAND U29825 ( .A(n29198), .B(n29197), .Z(n29199) );
  AND U29826 ( .A(n29200), .B(n29199), .Z(n29331) );
  XNOR U29827 ( .A(n29330), .B(n29331), .Z(n29332) );
  XOR U29828 ( .A(n1056), .B(a[189]), .Z(n29346) );
  NANDN U29829 ( .A(n29346), .B(n38101), .Z(n29203) );
  NANDN U29830 ( .A(n29201), .B(n38102), .Z(n29202) );
  NAND U29831 ( .A(n29203), .B(n29202), .Z(n29322) );
  XOR U29832 ( .A(b[15]), .B(n31434), .Z(n29343) );
  OR U29833 ( .A(n29343), .B(n37665), .Z(n29206) );
  NAND U29834 ( .A(n29204), .B(n37604), .Z(n29205) );
  AND U29835 ( .A(n29206), .B(n29205), .Z(n29323) );
  XNOR U29836 ( .A(n29322), .B(n29323), .Z(n29325) );
  XOR U29837 ( .A(n1052), .B(a[201]), .Z(n29340) );
  NANDN U29838 ( .A(n29340), .B(n36925), .Z(n29209) );
  NANDN U29839 ( .A(n29207), .B(n36926), .Z(n29208) );
  NAND U29840 ( .A(n29209), .B(n29208), .Z(n29324) );
  XNOR U29841 ( .A(n29325), .B(n29324), .Z(n29318) );
  XNOR U29842 ( .A(b[11]), .B(a[199]), .Z(n29349) );
  OR U29843 ( .A(n29349), .B(n37311), .Z(n29212) );
  NANDN U29844 ( .A(n29210), .B(n37218), .Z(n29211) );
  NAND U29845 ( .A(n29212), .B(n29211), .Z(n29317) );
  XOR U29846 ( .A(n1053), .B(a[197]), .Z(n29352) );
  NANDN U29847 ( .A(n29352), .B(n37424), .Z(n29215) );
  NANDN U29848 ( .A(n29213), .B(n37425), .Z(n29214) );
  NAND U29849 ( .A(n29215), .B(n29214), .Z(n29316) );
  XNOR U29850 ( .A(n29317), .B(n29316), .Z(n29319) );
  XNOR U29851 ( .A(n29318), .B(n29319), .Z(n29307) );
  NANDN U29852 ( .A(n1049), .B(a[209]), .Z(n29216) );
  XNOR U29853 ( .A(b[1]), .B(n29216), .Z(n29218) );
  NANDN U29854 ( .A(b[0]), .B(a[208]), .Z(n29217) );
  AND U29855 ( .A(n29218), .B(n29217), .Z(n29282) );
  NAND U29856 ( .A(n38490), .B(n29219), .Z(n29221) );
  XNOR U29857 ( .A(n1058), .B(a[181]), .Z(n29358) );
  NANDN U29858 ( .A(n1048), .B(n29358), .Z(n29220) );
  NAND U29859 ( .A(n29221), .B(n29220), .Z(n29280) );
  NANDN U29860 ( .A(n1059), .B(a[177]), .Z(n29281) );
  XNOR U29861 ( .A(n29280), .B(n29281), .Z(n29283) );
  XNOR U29862 ( .A(n29282), .B(n29283), .Z(n29305) );
  NANDN U29863 ( .A(n29222), .B(n38205), .Z(n29224) );
  XNOR U29864 ( .A(b[23]), .B(a[187]), .Z(n29361) );
  OR U29865 ( .A(n29361), .B(n38268), .Z(n29223) );
  NAND U29866 ( .A(n29224), .B(n29223), .Z(n29379) );
  XOR U29867 ( .A(b[7]), .B(a[203]), .Z(n29364) );
  NAND U29868 ( .A(n29364), .B(n36701), .Z(n29227) );
  NAND U29869 ( .A(n29225), .B(n36702), .Z(n29226) );
  NAND U29870 ( .A(n29227), .B(n29226), .Z(n29376) );
  XOR U29871 ( .A(b[25]), .B(a[185]), .Z(n29367) );
  NAND U29872 ( .A(n29367), .B(n38325), .Z(n29230) );
  NAND U29873 ( .A(n29228), .B(n38326), .Z(n29229) );
  AND U29874 ( .A(n29230), .B(n29229), .Z(n29377) );
  XNOR U29875 ( .A(n29376), .B(n29377), .Z(n29378) );
  XOR U29876 ( .A(n29379), .B(n29378), .Z(n29304) );
  XOR U29877 ( .A(n29307), .B(n29306), .Z(n29333) );
  XNOR U29878 ( .A(n29332), .B(n29333), .Z(n29270) );
  XNOR U29879 ( .A(n29271), .B(n29270), .Z(n29273) );
  XNOR U29880 ( .A(n29272), .B(n29273), .Z(n29388) );
  XOR U29881 ( .A(n29389), .B(n29388), .Z(n29391) );
  NAND U29882 ( .A(n29236), .B(n29235), .Z(n29240) );
  NAND U29883 ( .A(n29238), .B(n29237), .Z(n29239) );
  AND U29884 ( .A(n29240), .B(n29239), .Z(n29382) );
  XNOR U29885 ( .A(n29383), .B(n29382), .Z(n29384) );
  XOR U29886 ( .A(n29385), .B(n29384), .Z(n29266) );
  NANDN U29887 ( .A(n29242), .B(n29241), .Z(n29246) );
  NAND U29888 ( .A(n29244), .B(n29243), .Z(n29245) );
  NAND U29889 ( .A(n29246), .B(n29245), .Z(n29264) );
  NANDN U29890 ( .A(n29248), .B(n29247), .Z(n29252) );
  NAND U29891 ( .A(n29250), .B(n29249), .Z(n29251) );
  AND U29892 ( .A(n29252), .B(n29251), .Z(n29265) );
  XNOR U29893 ( .A(n29264), .B(n29265), .Z(n29267) );
  XOR U29894 ( .A(n29266), .B(n29267), .Z(n29258) );
  XOR U29895 ( .A(n29259), .B(n29258), .Z(n29260) );
  XNOR U29896 ( .A(n29261), .B(n29260), .Z(n29394) );
  XNOR U29897 ( .A(n29394), .B(sreg[433]), .Z(n29396) );
  NAND U29898 ( .A(n29253), .B(sreg[432]), .Z(n29257) );
  OR U29899 ( .A(n29255), .B(n29254), .Z(n29256) );
  AND U29900 ( .A(n29257), .B(n29256), .Z(n29395) );
  XOR U29901 ( .A(n29396), .B(n29395), .Z(c[433]) );
  NAND U29902 ( .A(n29259), .B(n29258), .Z(n29263) );
  NAND U29903 ( .A(n29261), .B(n29260), .Z(n29262) );
  NAND U29904 ( .A(n29263), .B(n29262), .Z(n29402) );
  NANDN U29905 ( .A(n29265), .B(n29264), .Z(n29269) );
  NAND U29906 ( .A(n29267), .B(n29266), .Z(n29268) );
  NAND U29907 ( .A(n29269), .B(n29268), .Z(n29399) );
  NAND U29908 ( .A(n29271), .B(n29270), .Z(n29275) );
  NANDN U29909 ( .A(n29273), .B(n29272), .Z(n29274) );
  NAND U29910 ( .A(n29275), .B(n29274), .Z(n29525) );
  XNOR U29911 ( .A(n29525), .B(n29526), .Z(n29527) );
  NANDN U29912 ( .A(n29281), .B(n29280), .Z(n29285) );
  NAND U29913 ( .A(n29283), .B(n29282), .Z(n29284) );
  NAND U29914 ( .A(n29285), .B(n29284), .Z(n29470) );
  XNOR U29915 ( .A(b[19]), .B(a[192]), .Z(n29417) );
  NANDN U29916 ( .A(n29417), .B(n37934), .Z(n29288) );
  NANDN U29917 ( .A(n29286), .B(n37935), .Z(n29287) );
  NAND U29918 ( .A(n29288), .B(n29287), .Z(n29480) );
  XOR U29919 ( .A(b[27]), .B(a[184]), .Z(n29420) );
  NAND U29920 ( .A(n38423), .B(n29420), .Z(n29291) );
  NAND U29921 ( .A(n29289), .B(n38424), .Z(n29290) );
  NAND U29922 ( .A(n29291), .B(n29290), .Z(n29477) );
  XNOR U29923 ( .A(b[5]), .B(a[206]), .Z(n29423) );
  NANDN U29924 ( .A(n29423), .B(n36587), .Z(n29294) );
  NANDN U29925 ( .A(n29292), .B(n36588), .Z(n29293) );
  AND U29926 ( .A(n29294), .B(n29293), .Z(n29478) );
  XNOR U29927 ( .A(n29477), .B(n29478), .Z(n29479) );
  XNOR U29928 ( .A(n29480), .B(n29479), .Z(n29468) );
  NANDN U29929 ( .A(n29295), .B(n37762), .Z(n29297) );
  XNOR U29930 ( .A(b[17]), .B(a[194]), .Z(n29426) );
  NANDN U29931 ( .A(n29426), .B(n37764), .Z(n29296) );
  NAND U29932 ( .A(n29297), .B(n29296), .Z(n29444) );
  XNOR U29933 ( .A(b[31]), .B(a[180]), .Z(n29429) );
  NANDN U29934 ( .A(n29429), .B(n38552), .Z(n29300) );
  NANDN U29935 ( .A(n29298), .B(n38553), .Z(n29299) );
  NAND U29936 ( .A(n29300), .B(n29299), .Z(n29441) );
  OR U29937 ( .A(n29301), .B(n36105), .Z(n29303) );
  XNOR U29938 ( .A(b[3]), .B(a[208]), .Z(n29432) );
  NANDN U29939 ( .A(n29432), .B(n36107), .Z(n29302) );
  AND U29940 ( .A(n29303), .B(n29302), .Z(n29442) );
  XNOR U29941 ( .A(n29441), .B(n29442), .Z(n29443) );
  XOR U29942 ( .A(n29444), .B(n29443), .Z(n29467) );
  XNOR U29943 ( .A(n29468), .B(n29467), .Z(n29469) );
  XNOR U29944 ( .A(n29470), .B(n29469), .Z(n29519) );
  NANDN U29945 ( .A(n29305), .B(n29304), .Z(n29309) );
  NANDN U29946 ( .A(n29307), .B(n29306), .Z(n29308) );
  NAND U29947 ( .A(n29309), .B(n29308), .Z(n29520) );
  XNOR U29948 ( .A(n29519), .B(n29520), .Z(n29521) );
  NANDN U29949 ( .A(n29311), .B(n29310), .Z(n29315) );
  NAND U29950 ( .A(n29313), .B(n29312), .Z(n29314) );
  NAND U29951 ( .A(n29315), .B(n29314), .Z(n29460) );
  OR U29952 ( .A(n29317), .B(n29316), .Z(n29321) );
  NANDN U29953 ( .A(n29319), .B(n29318), .Z(n29320) );
  NAND U29954 ( .A(n29321), .B(n29320), .Z(n29458) );
  XNOR U29955 ( .A(n29458), .B(n29457), .Z(n29459) );
  XOR U29956 ( .A(n29460), .B(n29459), .Z(n29522) );
  XOR U29957 ( .A(n29521), .B(n29522), .Z(n29533) );
  NANDN U29958 ( .A(n29331), .B(n29330), .Z(n29335) );
  NANDN U29959 ( .A(n29333), .B(n29332), .Z(n29334) );
  NAND U29960 ( .A(n29335), .B(n29334), .Z(n29516) );
  XNOR U29961 ( .A(b[9]), .B(a[202]), .Z(n29483) );
  NANDN U29962 ( .A(n29483), .B(n36925), .Z(n29342) );
  NANDN U29963 ( .A(n29340), .B(n36926), .Z(n29341) );
  NAND U29964 ( .A(n29342), .B(n29341), .Z(n29449) );
  XNOR U29965 ( .A(n1054), .B(a[196]), .Z(n29486) );
  NANDN U29966 ( .A(n37665), .B(n29486), .Z(n29345) );
  NANDN U29967 ( .A(n29343), .B(n37604), .Z(n29344) );
  NAND U29968 ( .A(n29345), .B(n29344), .Z(n29447) );
  XNOR U29969 ( .A(b[21]), .B(a[190]), .Z(n29489) );
  NANDN U29970 ( .A(n29489), .B(n38101), .Z(n29348) );
  NANDN U29971 ( .A(n29346), .B(n38102), .Z(n29347) );
  NAND U29972 ( .A(n29348), .B(n29347), .Z(n29448) );
  XNOR U29973 ( .A(n29447), .B(n29448), .Z(n29450) );
  XOR U29974 ( .A(n29449), .B(n29450), .Z(n29438) );
  XNOR U29975 ( .A(b[11]), .B(a[200]), .Z(n29492) );
  OR U29976 ( .A(n29492), .B(n37311), .Z(n29351) );
  NANDN U29977 ( .A(n29349), .B(n37218), .Z(n29350) );
  NAND U29978 ( .A(n29351), .B(n29350), .Z(n29436) );
  XOR U29979 ( .A(n1053), .B(a[198]), .Z(n29495) );
  NANDN U29980 ( .A(n29495), .B(n37424), .Z(n29354) );
  NANDN U29981 ( .A(n29352), .B(n37425), .Z(n29353) );
  AND U29982 ( .A(n29354), .B(n29353), .Z(n29435) );
  XNOR U29983 ( .A(n29436), .B(n29435), .Z(n29437) );
  XNOR U29984 ( .A(n29438), .B(n29437), .Z(n29454) );
  NANDN U29985 ( .A(n1049), .B(a[210]), .Z(n29355) );
  XNOR U29986 ( .A(b[1]), .B(n29355), .Z(n29357) );
  NANDN U29987 ( .A(b[0]), .B(a[209]), .Z(n29356) );
  AND U29988 ( .A(n29357), .B(n29356), .Z(n29413) );
  NAND U29989 ( .A(n38490), .B(n29358), .Z(n29360) );
  XNOR U29990 ( .A(n1058), .B(a[182]), .Z(n29501) );
  NANDN U29991 ( .A(n1048), .B(n29501), .Z(n29359) );
  NAND U29992 ( .A(n29360), .B(n29359), .Z(n29411) );
  NANDN U29993 ( .A(n1059), .B(a[178]), .Z(n29412) );
  XNOR U29994 ( .A(n29411), .B(n29412), .Z(n29414) );
  XNOR U29995 ( .A(n29413), .B(n29414), .Z(n29452) );
  NANDN U29996 ( .A(n29361), .B(n38205), .Z(n29363) );
  XNOR U29997 ( .A(b[23]), .B(a[188]), .Z(n29504) );
  OR U29998 ( .A(n29504), .B(n38268), .Z(n29362) );
  NAND U29999 ( .A(n29363), .B(n29362), .Z(n29474) );
  XNOR U30000 ( .A(b[7]), .B(a[204]), .Z(n29507) );
  NANDN U30001 ( .A(n29507), .B(n36701), .Z(n29366) );
  NAND U30002 ( .A(n29364), .B(n36702), .Z(n29365) );
  NAND U30003 ( .A(n29366), .B(n29365), .Z(n29471) );
  XOR U30004 ( .A(b[25]), .B(a[186]), .Z(n29510) );
  NAND U30005 ( .A(n29510), .B(n38325), .Z(n29369) );
  NAND U30006 ( .A(n29367), .B(n38326), .Z(n29368) );
  AND U30007 ( .A(n29369), .B(n29368), .Z(n29472) );
  XNOR U30008 ( .A(n29471), .B(n29472), .Z(n29473) );
  XOR U30009 ( .A(n29474), .B(n29473), .Z(n29451) );
  XOR U30010 ( .A(n29454), .B(n29453), .Z(n29464) );
  NANDN U30011 ( .A(n29371), .B(n29370), .Z(n29375) );
  NAND U30012 ( .A(n29373), .B(n29372), .Z(n29374) );
  NAND U30013 ( .A(n29375), .B(n29374), .Z(n29462) );
  NANDN U30014 ( .A(n29377), .B(n29376), .Z(n29381) );
  NAND U30015 ( .A(n29379), .B(n29378), .Z(n29380) );
  AND U30016 ( .A(n29381), .B(n29380), .Z(n29461) );
  XNOR U30017 ( .A(n29462), .B(n29461), .Z(n29463) );
  XNOR U30018 ( .A(n29464), .B(n29463), .Z(n29514) );
  XNOR U30019 ( .A(n29513), .B(n29514), .Z(n29515) );
  XNOR U30020 ( .A(n29516), .B(n29515), .Z(n29531) );
  XNOR U30021 ( .A(n29532), .B(n29531), .Z(n29534) );
  XNOR U30022 ( .A(n29533), .B(n29534), .Z(n29528) );
  XOR U30023 ( .A(n29527), .B(n29528), .Z(n29408) );
  NANDN U30024 ( .A(n29383), .B(n29382), .Z(n29387) );
  NAND U30025 ( .A(n29385), .B(n29384), .Z(n29386) );
  NAND U30026 ( .A(n29387), .B(n29386), .Z(n29405) );
  NANDN U30027 ( .A(n29389), .B(n29388), .Z(n29393) );
  OR U30028 ( .A(n29391), .B(n29390), .Z(n29392) );
  NAND U30029 ( .A(n29393), .B(n29392), .Z(n29406) );
  XNOR U30030 ( .A(n29405), .B(n29406), .Z(n29407) );
  XNOR U30031 ( .A(n29408), .B(n29407), .Z(n29400) );
  XNOR U30032 ( .A(n29399), .B(n29400), .Z(n29401) );
  XNOR U30033 ( .A(n29402), .B(n29401), .Z(n29537) );
  XNOR U30034 ( .A(n29537), .B(sreg[434]), .Z(n29539) );
  NAND U30035 ( .A(n29394), .B(sreg[433]), .Z(n29398) );
  OR U30036 ( .A(n29396), .B(n29395), .Z(n29397) );
  AND U30037 ( .A(n29398), .B(n29397), .Z(n29538) );
  XOR U30038 ( .A(n29539), .B(n29538), .Z(c[434]) );
  NANDN U30039 ( .A(n29400), .B(n29399), .Z(n29404) );
  NAND U30040 ( .A(n29402), .B(n29401), .Z(n29403) );
  NAND U30041 ( .A(n29404), .B(n29403), .Z(n29545) );
  NANDN U30042 ( .A(n29406), .B(n29405), .Z(n29410) );
  NAND U30043 ( .A(n29408), .B(n29407), .Z(n29409) );
  NAND U30044 ( .A(n29410), .B(n29409), .Z(n29543) );
  NANDN U30045 ( .A(n29412), .B(n29411), .Z(n29416) );
  NAND U30046 ( .A(n29414), .B(n29413), .Z(n29415) );
  NAND U30047 ( .A(n29416), .B(n29415), .Z(n29623) );
  XOR U30048 ( .A(b[19]), .B(n31508), .Z(n29568) );
  NANDN U30049 ( .A(n29568), .B(n37934), .Z(n29419) );
  NANDN U30050 ( .A(n29417), .B(n37935), .Z(n29418) );
  NAND U30051 ( .A(n29419), .B(n29418), .Z(n29633) );
  XOR U30052 ( .A(b[27]), .B(a[185]), .Z(n29571) );
  NAND U30053 ( .A(n38423), .B(n29571), .Z(n29422) );
  NAND U30054 ( .A(n29420), .B(n38424), .Z(n29421) );
  NAND U30055 ( .A(n29422), .B(n29421), .Z(n29630) );
  XNOR U30056 ( .A(b[5]), .B(a[207]), .Z(n29574) );
  NANDN U30057 ( .A(n29574), .B(n36587), .Z(n29425) );
  NANDN U30058 ( .A(n29423), .B(n36588), .Z(n29424) );
  AND U30059 ( .A(n29425), .B(n29424), .Z(n29631) );
  XNOR U30060 ( .A(n29630), .B(n29631), .Z(n29632) );
  XNOR U30061 ( .A(n29633), .B(n29632), .Z(n29621) );
  NANDN U30062 ( .A(n29426), .B(n37762), .Z(n29428) );
  XNOR U30063 ( .A(b[17]), .B(a[195]), .Z(n29577) );
  NANDN U30064 ( .A(n29577), .B(n37764), .Z(n29427) );
  NAND U30065 ( .A(n29428), .B(n29427), .Z(n29595) );
  XNOR U30066 ( .A(b[31]), .B(a[181]), .Z(n29580) );
  NANDN U30067 ( .A(n29580), .B(n38552), .Z(n29431) );
  NANDN U30068 ( .A(n29429), .B(n38553), .Z(n29430) );
  NAND U30069 ( .A(n29431), .B(n29430), .Z(n29592) );
  OR U30070 ( .A(n29432), .B(n36105), .Z(n29434) );
  XNOR U30071 ( .A(b[3]), .B(a[209]), .Z(n29583) );
  NANDN U30072 ( .A(n29583), .B(n36107), .Z(n29433) );
  AND U30073 ( .A(n29434), .B(n29433), .Z(n29593) );
  XNOR U30074 ( .A(n29592), .B(n29593), .Z(n29594) );
  XOR U30075 ( .A(n29595), .B(n29594), .Z(n29620) );
  XNOR U30076 ( .A(n29621), .B(n29620), .Z(n29622) );
  XNOR U30077 ( .A(n29623), .B(n29622), .Z(n29559) );
  NANDN U30078 ( .A(n29436), .B(n29435), .Z(n29440) );
  NAND U30079 ( .A(n29438), .B(n29437), .Z(n29439) );
  NAND U30080 ( .A(n29440), .B(n29439), .Z(n29612) );
  NANDN U30081 ( .A(n29442), .B(n29441), .Z(n29446) );
  NAND U30082 ( .A(n29444), .B(n29443), .Z(n29445) );
  NAND U30083 ( .A(n29446), .B(n29445), .Z(n29611) );
  XNOR U30084 ( .A(n29611), .B(n29610), .Z(n29613) );
  XOR U30085 ( .A(n29612), .B(n29613), .Z(n29558) );
  XOR U30086 ( .A(n29559), .B(n29558), .Z(n29560) );
  NANDN U30087 ( .A(n29452), .B(n29451), .Z(n29456) );
  NAND U30088 ( .A(n29454), .B(n29453), .Z(n29455) );
  AND U30089 ( .A(n29456), .B(n29455), .Z(n29561) );
  XNOR U30090 ( .A(n29560), .B(n29561), .Z(n29669) );
  NANDN U30091 ( .A(n29462), .B(n29461), .Z(n29466) );
  NANDN U30092 ( .A(n29464), .B(n29463), .Z(n29465) );
  NAND U30093 ( .A(n29466), .B(n29465), .Z(n29555) );
  NANDN U30094 ( .A(n29472), .B(n29471), .Z(n29476) );
  NAND U30095 ( .A(n29474), .B(n29473), .Z(n29475) );
  NAND U30096 ( .A(n29476), .B(n29475), .Z(n29614) );
  NANDN U30097 ( .A(n29478), .B(n29477), .Z(n29482) );
  NAND U30098 ( .A(n29480), .B(n29479), .Z(n29481) );
  AND U30099 ( .A(n29482), .B(n29481), .Z(n29615) );
  XNOR U30100 ( .A(n29614), .B(n29615), .Z(n29616) );
  XNOR U30101 ( .A(n1052), .B(a[203]), .Z(n29636) );
  NAND U30102 ( .A(n36925), .B(n29636), .Z(n29485) );
  NANDN U30103 ( .A(n29483), .B(n36926), .Z(n29484) );
  NAND U30104 ( .A(n29485), .B(n29484), .Z(n29600) );
  XNOR U30105 ( .A(b[15]), .B(a[197]), .Z(n29639) );
  OR U30106 ( .A(n29639), .B(n37665), .Z(n29488) );
  NAND U30107 ( .A(n29486), .B(n37604), .Z(n29487) );
  AND U30108 ( .A(n29488), .B(n29487), .Z(n29598) );
  XNOR U30109 ( .A(n1056), .B(a[191]), .Z(n29642) );
  NAND U30110 ( .A(n29642), .B(n38101), .Z(n29491) );
  NANDN U30111 ( .A(n29489), .B(n38102), .Z(n29490) );
  AND U30112 ( .A(n29491), .B(n29490), .Z(n29599) );
  XOR U30113 ( .A(n29600), .B(n29601), .Z(n29589) );
  XOR U30114 ( .A(b[11]), .B(n32687), .Z(n29645) );
  OR U30115 ( .A(n29645), .B(n37311), .Z(n29494) );
  NANDN U30116 ( .A(n29492), .B(n37218), .Z(n29493) );
  NAND U30117 ( .A(n29494), .B(n29493), .Z(n29587) );
  XOR U30118 ( .A(n1053), .B(a[199]), .Z(n29648) );
  NANDN U30119 ( .A(n29648), .B(n37424), .Z(n29497) );
  NANDN U30120 ( .A(n29495), .B(n37425), .Z(n29496) );
  AND U30121 ( .A(n29497), .B(n29496), .Z(n29586) );
  XNOR U30122 ( .A(n29587), .B(n29586), .Z(n29588) );
  XOR U30123 ( .A(n29589), .B(n29588), .Z(n29606) );
  NANDN U30124 ( .A(n1049), .B(a[211]), .Z(n29498) );
  XNOR U30125 ( .A(b[1]), .B(n29498), .Z(n29500) );
  NANDN U30126 ( .A(b[0]), .B(a[210]), .Z(n29499) );
  AND U30127 ( .A(n29500), .B(n29499), .Z(n29564) );
  NAND U30128 ( .A(n38490), .B(n29501), .Z(n29503) );
  XNOR U30129 ( .A(n1058), .B(a[183]), .Z(n29654) );
  NANDN U30130 ( .A(n1048), .B(n29654), .Z(n29502) );
  NAND U30131 ( .A(n29503), .B(n29502), .Z(n29562) );
  NANDN U30132 ( .A(n1059), .B(a[179]), .Z(n29563) );
  XNOR U30133 ( .A(n29562), .B(n29563), .Z(n29565) );
  XOR U30134 ( .A(n29564), .B(n29565), .Z(n29604) );
  NANDN U30135 ( .A(n29504), .B(n38205), .Z(n29506) );
  XOR U30136 ( .A(b[23]), .B(n30936), .Z(n29657) );
  OR U30137 ( .A(n29657), .B(n38268), .Z(n29505) );
  NAND U30138 ( .A(n29506), .B(n29505), .Z(n29627) );
  XOR U30139 ( .A(b[7]), .B(a[205]), .Z(n29660) );
  NAND U30140 ( .A(n29660), .B(n36701), .Z(n29509) );
  NANDN U30141 ( .A(n29507), .B(n36702), .Z(n29508) );
  NAND U30142 ( .A(n29509), .B(n29508), .Z(n29624) );
  XOR U30143 ( .A(b[25]), .B(a[187]), .Z(n29663) );
  NAND U30144 ( .A(n29663), .B(n38325), .Z(n29512) );
  NAND U30145 ( .A(n29510), .B(n38326), .Z(n29511) );
  AND U30146 ( .A(n29512), .B(n29511), .Z(n29625) );
  XNOR U30147 ( .A(n29624), .B(n29625), .Z(n29626) );
  XNOR U30148 ( .A(n29627), .B(n29626), .Z(n29605) );
  XOR U30149 ( .A(n29604), .B(n29605), .Z(n29607) );
  XNOR U30150 ( .A(n29606), .B(n29607), .Z(n29617) );
  XNOR U30151 ( .A(n29616), .B(n29617), .Z(n29552) );
  XNOR U30152 ( .A(n29553), .B(n29552), .Z(n29554) );
  XOR U30153 ( .A(n29555), .B(n29554), .Z(n29667) );
  XNOR U30154 ( .A(n29666), .B(n29667), .Z(n29668) );
  XNOR U30155 ( .A(n29669), .B(n29668), .Z(n29673) );
  NANDN U30156 ( .A(n29514), .B(n29513), .Z(n29518) );
  NAND U30157 ( .A(n29516), .B(n29515), .Z(n29517) );
  NAND U30158 ( .A(n29518), .B(n29517), .Z(n29670) );
  NANDN U30159 ( .A(n29520), .B(n29519), .Z(n29524) );
  NAND U30160 ( .A(n29522), .B(n29521), .Z(n29523) );
  NAND U30161 ( .A(n29524), .B(n29523), .Z(n29671) );
  XNOR U30162 ( .A(n29670), .B(n29671), .Z(n29672) );
  XNOR U30163 ( .A(n29673), .B(n29672), .Z(n29549) );
  NANDN U30164 ( .A(n29526), .B(n29525), .Z(n29530) );
  NANDN U30165 ( .A(n29528), .B(n29527), .Z(n29529) );
  NAND U30166 ( .A(n29530), .B(n29529), .Z(n29547) );
  OR U30167 ( .A(n29532), .B(n29531), .Z(n29536) );
  OR U30168 ( .A(n29534), .B(n29533), .Z(n29535) );
  AND U30169 ( .A(n29536), .B(n29535), .Z(n29546) );
  XNOR U30170 ( .A(n29547), .B(n29546), .Z(n29548) );
  XNOR U30171 ( .A(n29549), .B(n29548), .Z(n29542) );
  XOR U30172 ( .A(n29543), .B(n29542), .Z(n29544) );
  XNOR U30173 ( .A(n29545), .B(n29544), .Z(n29676) );
  XNOR U30174 ( .A(n29676), .B(sreg[435]), .Z(n29678) );
  NAND U30175 ( .A(n29537), .B(sreg[434]), .Z(n29541) );
  OR U30176 ( .A(n29539), .B(n29538), .Z(n29540) );
  AND U30177 ( .A(n29541), .B(n29540), .Z(n29677) );
  XOR U30178 ( .A(n29678), .B(n29677), .Z(c[435]) );
  NANDN U30179 ( .A(n29547), .B(n29546), .Z(n29551) );
  NANDN U30180 ( .A(n29549), .B(n29548), .Z(n29550) );
  NAND U30181 ( .A(n29551), .B(n29550), .Z(n29681) );
  NAND U30182 ( .A(n29553), .B(n29552), .Z(n29557) );
  OR U30183 ( .A(n29555), .B(n29554), .Z(n29556) );
  NAND U30184 ( .A(n29557), .B(n29556), .Z(n29693) );
  XNOR U30185 ( .A(n29693), .B(n29694), .Z(n29695) );
  NANDN U30186 ( .A(n29563), .B(n29562), .Z(n29567) );
  NAND U30187 ( .A(n29565), .B(n29564), .Z(n29566) );
  NAND U30188 ( .A(n29567), .B(n29566), .Z(n29766) );
  XOR U30189 ( .A(b[19]), .B(n31644), .Z(n29711) );
  NANDN U30190 ( .A(n29711), .B(n37934), .Z(n29570) );
  NANDN U30191 ( .A(n29568), .B(n37935), .Z(n29569) );
  NAND U30192 ( .A(n29570), .B(n29569), .Z(n29776) );
  XOR U30193 ( .A(b[27]), .B(a[186]), .Z(n29714) );
  NAND U30194 ( .A(n38423), .B(n29714), .Z(n29573) );
  NAND U30195 ( .A(n29571), .B(n38424), .Z(n29572) );
  NAND U30196 ( .A(n29573), .B(n29572), .Z(n29773) );
  XNOR U30197 ( .A(b[5]), .B(a[208]), .Z(n29717) );
  NANDN U30198 ( .A(n29717), .B(n36587), .Z(n29576) );
  NANDN U30199 ( .A(n29574), .B(n36588), .Z(n29575) );
  AND U30200 ( .A(n29576), .B(n29575), .Z(n29774) );
  XNOR U30201 ( .A(n29773), .B(n29774), .Z(n29775) );
  XNOR U30202 ( .A(n29776), .B(n29775), .Z(n29764) );
  NANDN U30203 ( .A(n29577), .B(n37762), .Z(n29579) );
  XOR U30204 ( .A(b[17]), .B(a[196]), .Z(n29720) );
  NAND U30205 ( .A(n29720), .B(n37764), .Z(n29578) );
  NAND U30206 ( .A(n29579), .B(n29578), .Z(n29738) );
  XNOR U30207 ( .A(b[31]), .B(a[182]), .Z(n29723) );
  NANDN U30208 ( .A(n29723), .B(n38552), .Z(n29582) );
  NANDN U30209 ( .A(n29580), .B(n38553), .Z(n29581) );
  NAND U30210 ( .A(n29582), .B(n29581), .Z(n29735) );
  OR U30211 ( .A(n29583), .B(n36105), .Z(n29585) );
  XNOR U30212 ( .A(b[3]), .B(a[210]), .Z(n29726) );
  NANDN U30213 ( .A(n29726), .B(n36107), .Z(n29584) );
  AND U30214 ( .A(n29585), .B(n29584), .Z(n29736) );
  XNOR U30215 ( .A(n29735), .B(n29736), .Z(n29737) );
  XOR U30216 ( .A(n29738), .B(n29737), .Z(n29763) );
  XNOR U30217 ( .A(n29764), .B(n29763), .Z(n29765) );
  XNOR U30218 ( .A(n29766), .B(n29765), .Z(n29809) );
  NANDN U30219 ( .A(n29587), .B(n29586), .Z(n29591) );
  NAND U30220 ( .A(n29589), .B(n29588), .Z(n29590) );
  NAND U30221 ( .A(n29591), .B(n29590), .Z(n29754) );
  NANDN U30222 ( .A(n29593), .B(n29592), .Z(n29597) );
  NAND U30223 ( .A(n29595), .B(n29594), .Z(n29596) );
  NAND U30224 ( .A(n29597), .B(n29596), .Z(n29752) );
  OR U30225 ( .A(n29599), .B(n29598), .Z(n29603) );
  NANDN U30226 ( .A(n29601), .B(n29600), .Z(n29602) );
  NAND U30227 ( .A(n29603), .B(n29602), .Z(n29751) );
  XNOR U30228 ( .A(n29754), .B(n29753), .Z(n29810) );
  XNOR U30229 ( .A(n29809), .B(n29810), .Z(n29811) );
  NANDN U30230 ( .A(n29605), .B(n29604), .Z(n29609) );
  OR U30231 ( .A(n29607), .B(n29606), .Z(n29608) );
  AND U30232 ( .A(n29609), .B(n29608), .Z(n29812) );
  XOR U30233 ( .A(n29811), .B(n29812), .Z(n29701) );
  NANDN U30234 ( .A(n29615), .B(n29614), .Z(n29619) );
  NANDN U30235 ( .A(n29617), .B(n29616), .Z(n29618) );
  NAND U30236 ( .A(n29619), .B(n29618), .Z(n29818) );
  NANDN U30237 ( .A(n29625), .B(n29624), .Z(n29629) );
  NAND U30238 ( .A(n29627), .B(n29626), .Z(n29628) );
  NAND U30239 ( .A(n29629), .B(n29628), .Z(n29757) );
  NANDN U30240 ( .A(n29631), .B(n29630), .Z(n29635) );
  NAND U30241 ( .A(n29633), .B(n29632), .Z(n29634) );
  AND U30242 ( .A(n29635), .B(n29634), .Z(n29758) );
  XNOR U30243 ( .A(n29757), .B(n29758), .Z(n29759) );
  XOR U30244 ( .A(b[9]), .B(n33130), .Z(n29779) );
  NANDN U30245 ( .A(n29779), .B(n36925), .Z(n29638) );
  NAND U30246 ( .A(n36926), .B(n29636), .Z(n29637) );
  NAND U30247 ( .A(n29638), .B(n29637), .Z(n29743) );
  XNOR U30248 ( .A(n1054), .B(a[198]), .Z(n29782) );
  NANDN U30249 ( .A(n37665), .B(n29782), .Z(n29641) );
  NANDN U30250 ( .A(n29639), .B(n37604), .Z(n29640) );
  NAND U30251 ( .A(n29641), .B(n29640), .Z(n29741) );
  XNOR U30252 ( .A(b[21]), .B(a[192]), .Z(n29785) );
  NANDN U30253 ( .A(n29785), .B(n38101), .Z(n29644) );
  NAND U30254 ( .A(n38102), .B(n29642), .Z(n29643) );
  NAND U30255 ( .A(n29644), .B(n29643), .Z(n29742) );
  XNOR U30256 ( .A(n29741), .B(n29742), .Z(n29744) );
  XOR U30257 ( .A(n29743), .B(n29744), .Z(n29732) );
  XNOR U30258 ( .A(b[11]), .B(a[202]), .Z(n29788) );
  OR U30259 ( .A(n29788), .B(n37311), .Z(n29647) );
  NANDN U30260 ( .A(n29645), .B(n37218), .Z(n29646) );
  NAND U30261 ( .A(n29647), .B(n29646), .Z(n29730) );
  XOR U30262 ( .A(n1053), .B(a[200]), .Z(n29791) );
  NANDN U30263 ( .A(n29791), .B(n37424), .Z(n29650) );
  NANDN U30264 ( .A(n29648), .B(n37425), .Z(n29649) );
  AND U30265 ( .A(n29650), .B(n29649), .Z(n29729) );
  XNOR U30266 ( .A(n29730), .B(n29729), .Z(n29731) );
  XNOR U30267 ( .A(n29732), .B(n29731), .Z(n29748) );
  NANDN U30268 ( .A(n1049), .B(a[212]), .Z(n29651) );
  XNOR U30269 ( .A(b[1]), .B(n29651), .Z(n29653) );
  NANDN U30270 ( .A(b[0]), .B(a[211]), .Z(n29652) );
  AND U30271 ( .A(n29653), .B(n29652), .Z(n29707) );
  NAND U30272 ( .A(n38490), .B(n29654), .Z(n29656) );
  XNOR U30273 ( .A(n1058), .B(a[184]), .Z(n29797) );
  NANDN U30274 ( .A(n1048), .B(n29797), .Z(n29655) );
  NAND U30275 ( .A(n29656), .B(n29655), .Z(n29705) );
  NANDN U30276 ( .A(n1059), .B(a[180]), .Z(n29706) );
  XNOR U30277 ( .A(n29705), .B(n29706), .Z(n29708) );
  XNOR U30278 ( .A(n29707), .B(n29708), .Z(n29746) );
  NANDN U30279 ( .A(n29657), .B(n38205), .Z(n29659) );
  XNOR U30280 ( .A(b[23]), .B(a[190]), .Z(n29800) );
  OR U30281 ( .A(n29800), .B(n38268), .Z(n29658) );
  NAND U30282 ( .A(n29659), .B(n29658), .Z(n29770) );
  XOR U30283 ( .A(b[7]), .B(a[206]), .Z(n29803) );
  NAND U30284 ( .A(n29803), .B(n36701), .Z(n29662) );
  NAND U30285 ( .A(n29660), .B(n36702), .Z(n29661) );
  NAND U30286 ( .A(n29662), .B(n29661), .Z(n29767) );
  XOR U30287 ( .A(b[25]), .B(a[188]), .Z(n29806) );
  NAND U30288 ( .A(n29806), .B(n38325), .Z(n29665) );
  NAND U30289 ( .A(n29663), .B(n38326), .Z(n29664) );
  AND U30290 ( .A(n29665), .B(n29664), .Z(n29768) );
  XNOR U30291 ( .A(n29767), .B(n29768), .Z(n29769) );
  XOR U30292 ( .A(n29770), .B(n29769), .Z(n29745) );
  XOR U30293 ( .A(n29748), .B(n29747), .Z(n29760) );
  XOR U30294 ( .A(n29759), .B(n29760), .Z(n29815) );
  XOR U30295 ( .A(n29816), .B(n29815), .Z(n29817) );
  XNOR U30296 ( .A(n29818), .B(n29817), .Z(n29699) );
  XNOR U30297 ( .A(n29700), .B(n29699), .Z(n29702) );
  XNOR U30298 ( .A(n29701), .B(n29702), .Z(n29696) );
  XOR U30299 ( .A(n29695), .B(n29696), .Z(n29690) );
  NANDN U30300 ( .A(n29671), .B(n29670), .Z(n29675) );
  NANDN U30301 ( .A(n29673), .B(n29672), .Z(n29674) );
  NAND U30302 ( .A(n29675), .B(n29674), .Z(n29688) );
  XNOR U30303 ( .A(n29687), .B(n29688), .Z(n29689) );
  XNOR U30304 ( .A(n29690), .B(n29689), .Z(n29682) );
  XNOR U30305 ( .A(n29681), .B(n29682), .Z(n29683) );
  XNOR U30306 ( .A(n29684), .B(n29683), .Z(n29821) );
  XNOR U30307 ( .A(n29821), .B(sreg[436]), .Z(n29823) );
  NAND U30308 ( .A(n29676), .B(sreg[435]), .Z(n29680) );
  OR U30309 ( .A(n29678), .B(n29677), .Z(n29679) );
  AND U30310 ( .A(n29680), .B(n29679), .Z(n29822) );
  XOR U30311 ( .A(n29823), .B(n29822), .Z(c[436]) );
  NANDN U30312 ( .A(n29682), .B(n29681), .Z(n29686) );
  NAND U30313 ( .A(n29684), .B(n29683), .Z(n29685) );
  NAND U30314 ( .A(n29686), .B(n29685), .Z(n29829) );
  NANDN U30315 ( .A(n29688), .B(n29687), .Z(n29692) );
  NAND U30316 ( .A(n29690), .B(n29689), .Z(n29691) );
  NAND U30317 ( .A(n29692), .B(n29691), .Z(n29827) );
  NANDN U30318 ( .A(n29694), .B(n29693), .Z(n29698) );
  NANDN U30319 ( .A(n29696), .B(n29695), .Z(n29697) );
  NAND U30320 ( .A(n29698), .B(n29697), .Z(n29833) );
  OR U30321 ( .A(n29700), .B(n29699), .Z(n29704) );
  OR U30322 ( .A(n29702), .B(n29701), .Z(n29703) );
  AND U30323 ( .A(n29704), .B(n29703), .Z(n29832) );
  XNOR U30324 ( .A(n29833), .B(n29832), .Z(n29834) );
  NANDN U30325 ( .A(n29706), .B(n29705), .Z(n29710) );
  NAND U30326 ( .A(n29708), .B(n29707), .Z(n29709) );
  NAND U30327 ( .A(n29710), .B(n29709), .Z(n29909) );
  XOR U30328 ( .A(b[19]), .B(n31434), .Z(n29854) );
  NANDN U30329 ( .A(n29854), .B(n37934), .Z(n29713) );
  NANDN U30330 ( .A(n29711), .B(n37935), .Z(n29712) );
  NAND U30331 ( .A(n29713), .B(n29712), .Z(n29919) );
  XOR U30332 ( .A(b[27]), .B(a[187]), .Z(n29857) );
  NAND U30333 ( .A(n38423), .B(n29857), .Z(n29716) );
  NAND U30334 ( .A(n29714), .B(n38424), .Z(n29715) );
  NAND U30335 ( .A(n29716), .B(n29715), .Z(n29916) );
  XNOR U30336 ( .A(b[5]), .B(a[209]), .Z(n29860) );
  NANDN U30337 ( .A(n29860), .B(n36587), .Z(n29719) );
  NANDN U30338 ( .A(n29717), .B(n36588), .Z(n29718) );
  AND U30339 ( .A(n29719), .B(n29718), .Z(n29917) );
  XNOR U30340 ( .A(n29916), .B(n29917), .Z(n29918) );
  XNOR U30341 ( .A(n29919), .B(n29918), .Z(n29907) );
  NAND U30342 ( .A(n29720), .B(n37762), .Z(n29722) );
  XOR U30343 ( .A(b[17]), .B(a[197]), .Z(n29863) );
  NAND U30344 ( .A(n29863), .B(n37764), .Z(n29721) );
  NAND U30345 ( .A(n29722), .B(n29721), .Z(n29881) );
  XNOR U30346 ( .A(b[31]), .B(a[183]), .Z(n29866) );
  NANDN U30347 ( .A(n29866), .B(n38552), .Z(n29725) );
  NANDN U30348 ( .A(n29723), .B(n38553), .Z(n29724) );
  NAND U30349 ( .A(n29725), .B(n29724), .Z(n29878) );
  OR U30350 ( .A(n29726), .B(n36105), .Z(n29728) );
  XNOR U30351 ( .A(b[3]), .B(a[211]), .Z(n29869) );
  NANDN U30352 ( .A(n29869), .B(n36107), .Z(n29727) );
  AND U30353 ( .A(n29728), .B(n29727), .Z(n29879) );
  XNOR U30354 ( .A(n29878), .B(n29879), .Z(n29880) );
  XOR U30355 ( .A(n29881), .B(n29880), .Z(n29906) );
  XNOR U30356 ( .A(n29907), .B(n29906), .Z(n29908) );
  XNOR U30357 ( .A(n29909), .B(n29908), .Z(n29845) );
  NANDN U30358 ( .A(n29730), .B(n29729), .Z(n29734) );
  NAND U30359 ( .A(n29732), .B(n29731), .Z(n29733) );
  NAND U30360 ( .A(n29734), .B(n29733), .Z(n29898) );
  NANDN U30361 ( .A(n29736), .B(n29735), .Z(n29740) );
  NAND U30362 ( .A(n29738), .B(n29737), .Z(n29739) );
  NAND U30363 ( .A(n29740), .B(n29739), .Z(n29897) );
  XNOR U30364 ( .A(n29897), .B(n29896), .Z(n29899) );
  XOR U30365 ( .A(n29898), .B(n29899), .Z(n29844) );
  XOR U30366 ( .A(n29845), .B(n29844), .Z(n29846) );
  NANDN U30367 ( .A(n29746), .B(n29745), .Z(n29750) );
  NAND U30368 ( .A(n29748), .B(n29747), .Z(n29749) );
  NAND U30369 ( .A(n29750), .B(n29749), .Z(n29847) );
  XNOR U30370 ( .A(n29846), .B(n29847), .Z(n29960) );
  OR U30371 ( .A(n29752), .B(n29751), .Z(n29756) );
  NAND U30372 ( .A(n29754), .B(n29753), .Z(n29755) );
  NAND U30373 ( .A(n29756), .B(n29755), .Z(n29959) );
  NANDN U30374 ( .A(n29758), .B(n29757), .Z(n29762) );
  NAND U30375 ( .A(n29760), .B(n29759), .Z(n29761) );
  NAND U30376 ( .A(n29762), .B(n29761), .Z(n29840) );
  NANDN U30377 ( .A(n29768), .B(n29767), .Z(n29772) );
  NAND U30378 ( .A(n29770), .B(n29769), .Z(n29771) );
  NAND U30379 ( .A(n29772), .B(n29771), .Z(n29900) );
  NANDN U30380 ( .A(n29774), .B(n29773), .Z(n29778) );
  NAND U30381 ( .A(n29776), .B(n29775), .Z(n29777) );
  AND U30382 ( .A(n29778), .B(n29777), .Z(n29901) );
  XNOR U30383 ( .A(n29900), .B(n29901), .Z(n29902) );
  XNOR U30384 ( .A(n1052), .B(a[205]), .Z(n29922) );
  NAND U30385 ( .A(n36925), .B(n29922), .Z(n29781) );
  NANDN U30386 ( .A(n29779), .B(n36926), .Z(n29780) );
  NAND U30387 ( .A(n29781), .B(n29780), .Z(n29886) );
  XNOR U30388 ( .A(b[15]), .B(a[199]), .Z(n29925) );
  OR U30389 ( .A(n29925), .B(n37665), .Z(n29784) );
  NAND U30390 ( .A(n29782), .B(n37604), .Z(n29783) );
  AND U30391 ( .A(n29784), .B(n29783), .Z(n29884) );
  XOR U30392 ( .A(n1056), .B(n31508), .Z(n29928) );
  NAND U30393 ( .A(n29928), .B(n38101), .Z(n29787) );
  NANDN U30394 ( .A(n29785), .B(n38102), .Z(n29786) );
  AND U30395 ( .A(n29787), .B(n29786), .Z(n29885) );
  XOR U30396 ( .A(n29886), .B(n29887), .Z(n29875) );
  XNOR U30397 ( .A(b[11]), .B(a[203]), .Z(n29931) );
  OR U30398 ( .A(n29931), .B(n37311), .Z(n29790) );
  NANDN U30399 ( .A(n29788), .B(n37218), .Z(n29789) );
  NAND U30400 ( .A(n29790), .B(n29789), .Z(n29873) );
  XOR U30401 ( .A(n1053), .B(a[201]), .Z(n29934) );
  NANDN U30402 ( .A(n29934), .B(n37424), .Z(n29793) );
  NANDN U30403 ( .A(n29791), .B(n37425), .Z(n29792) );
  AND U30404 ( .A(n29793), .B(n29792), .Z(n29872) );
  XNOR U30405 ( .A(n29873), .B(n29872), .Z(n29874) );
  XOR U30406 ( .A(n29875), .B(n29874), .Z(n29892) );
  NANDN U30407 ( .A(n1049), .B(a[213]), .Z(n29794) );
  XNOR U30408 ( .A(b[1]), .B(n29794), .Z(n29796) );
  NANDN U30409 ( .A(b[0]), .B(a[212]), .Z(n29795) );
  AND U30410 ( .A(n29796), .B(n29795), .Z(n29850) );
  NAND U30411 ( .A(n38490), .B(n29797), .Z(n29799) );
  XNOR U30412 ( .A(n1058), .B(a[185]), .Z(n29940) );
  NANDN U30413 ( .A(n1048), .B(n29940), .Z(n29798) );
  NAND U30414 ( .A(n29799), .B(n29798), .Z(n29848) );
  NANDN U30415 ( .A(n1059), .B(a[181]), .Z(n29849) );
  XNOR U30416 ( .A(n29848), .B(n29849), .Z(n29851) );
  XOR U30417 ( .A(n29850), .B(n29851), .Z(n29890) );
  NANDN U30418 ( .A(n29800), .B(n38205), .Z(n29802) );
  XNOR U30419 ( .A(b[23]), .B(a[191]), .Z(n29943) );
  OR U30420 ( .A(n29943), .B(n38268), .Z(n29801) );
  NAND U30421 ( .A(n29802), .B(n29801), .Z(n29913) );
  XOR U30422 ( .A(b[7]), .B(a[207]), .Z(n29946) );
  NAND U30423 ( .A(n29946), .B(n36701), .Z(n29805) );
  NAND U30424 ( .A(n29803), .B(n36702), .Z(n29804) );
  NAND U30425 ( .A(n29805), .B(n29804), .Z(n29910) );
  XNOR U30426 ( .A(b[25]), .B(a[189]), .Z(n29949) );
  NANDN U30427 ( .A(n29949), .B(n38325), .Z(n29808) );
  NAND U30428 ( .A(n29806), .B(n38326), .Z(n29807) );
  AND U30429 ( .A(n29808), .B(n29807), .Z(n29911) );
  XNOR U30430 ( .A(n29910), .B(n29911), .Z(n29912) );
  XNOR U30431 ( .A(n29913), .B(n29912), .Z(n29891) );
  XOR U30432 ( .A(n29890), .B(n29891), .Z(n29893) );
  XNOR U30433 ( .A(n29892), .B(n29893), .Z(n29903) );
  XNOR U30434 ( .A(n29902), .B(n29903), .Z(n29838) );
  XNOR U30435 ( .A(n29839), .B(n29838), .Z(n29841) );
  XNOR U30436 ( .A(n29840), .B(n29841), .Z(n29958) );
  XOR U30437 ( .A(n29959), .B(n29958), .Z(n29961) );
  NANDN U30438 ( .A(n29810), .B(n29809), .Z(n29814) );
  NAND U30439 ( .A(n29812), .B(n29811), .Z(n29813) );
  NAND U30440 ( .A(n29814), .B(n29813), .Z(n29952) );
  NAND U30441 ( .A(n29816), .B(n29815), .Z(n29820) );
  NAND U30442 ( .A(n29818), .B(n29817), .Z(n29819) );
  NAND U30443 ( .A(n29820), .B(n29819), .Z(n29953) );
  XNOR U30444 ( .A(n29952), .B(n29953), .Z(n29954) );
  XOR U30445 ( .A(n29955), .B(n29954), .Z(n29835) );
  XOR U30446 ( .A(n29834), .B(n29835), .Z(n29826) );
  XOR U30447 ( .A(n29827), .B(n29826), .Z(n29828) );
  XNOR U30448 ( .A(n29829), .B(n29828), .Z(n29964) );
  XNOR U30449 ( .A(n29964), .B(sreg[437]), .Z(n29966) );
  NAND U30450 ( .A(n29821), .B(sreg[436]), .Z(n29825) );
  OR U30451 ( .A(n29823), .B(n29822), .Z(n29824) );
  AND U30452 ( .A(n29825), .B(n29824), .Z(n29965) );
  XOR U30453 ( .A(n29966), .B(n29965), .Z(c[437]) );
  NAND U30454 ( .A(n29827), .B(n29826), .Z(n29831) );
  NAND U30455 ( .A(n29829), .B(n29828), .Z(n29830) );
  NAND U30456 ( .A(n29831), .B(n29830), .Z(n29972) );
  NANDN U30457 ( .A(n29833), .B(n29832), .Z(n29837) );
  NAND U30458 ( .A(n29835), .B(n29834), .Z(n29836) );
  NAND U30459 ( .A(n29837), .B(n29836), .Z(n29969) );
  NAND U30460 ( .A(n29839), .B(n29838), .Z(n29843) );
  NANDN U30461 ( .A(n29841), .B(n29840), .Z(n29842) );
  NAND U30462 ( .A(n29843), .B(n29842), .Z(n30097) );
  XNOR U30463 ( .A(n30097), .B(n30098), .Z(n30099) );
  NANDN U30464 ( .A(n29849), .B(n29848), .Z(n29853) );
  NAND U30465 ( .A(n29851), .B(n29850), .Z(n29852) );
  NAND U30466 ( .A(n29853), .B(n29852), .Z(n30042) );
  XNOR U30467 ( .A(b[19]), .B(a[196]), .Z(n29987) );
  NANDN U30468 ( .A(n29987), .B(n37934), .Z(n29856) );
  NANDN U30469 ( .A(n29854), .B(n37935), .Z(n29855) );
  NAND U30470 ( .A(n29856), .B(n29855), .Z(n30052) );
  XOR U30471 ( .A(b[27]), .B(a[188]), .Z(n29990) );
  NAND U30472 ( .A(n38423), .B(n29990), .Z(n29859) );
  NAND U30473 ( .A(n29857), .B(n38424), .Z(n29858) );
  NAND U30474 ( .A(n29859), .B(n29858), .Z(n30049) );
  XNOR U30475 ( .A(b[5]), .B(a[210]), .Z(n29993) );
  NANDN U30476 ( .A(n29993), .B(n36587), .Z(n29862) );
  NANDN U30477 ( .A(n29860), .B(n36588), .Z(n29861) );
  AND U30478 ( .A(n29862), .B(n29861), .Z(n30050) );
  XNOR U30479 ( .A(n30049), .B(n30050), .Z(n30051) );
  XNOR U30480 ( .A(n30052), .B(n30051), .Z(n30040) );
  NAND U30481 ( .A(n29863), .B(n37762), .Z(n29865) );
  XNOR U30482 ( .A(b[17]), .B(a[198]), .Z(n29996) );
  NANDN U30483 ( .A(n29996), .B(n37764), .Z(n29864) );
  NAND U30484 ( .A(n29865), .B(n29864), .Z(n30014) );
  XNOR U30485 ( .A(b[31]), .B(a[184]), .Z(n29999) );
  NANDN U30486 ( .A(n29999), .B(n38552), .Z(n29868) );
  NANDN U30487 ( .A(n29866), .B(n38553), .Z(n29867) );
  NAND U30488 ( .A(n29868), .B(n29867), .Z(n30011) );
  OR U30489 ( .A(n29869), .B(n36105), .Z(n29871) );
  XNOR U30490 ( .A(b[3]), .B(a[212]), .Z(n30002) );
  NANDN U30491 ( .A(n30002), .B(n36107), .Z(n29870) );
  AND U30492 ( .A(n29871), .B(n29870), .Z(n30012) );
  XNOR U30493 ( .A(n30011), .B(n30012), .Z(n30013) );
  XOR U30494 ( .A(n30014), .B(n30013), .Z(n30039) );
  XNOR U30495 ( .A(n30040), .B(n30039), .Z(n30041) );
  XNOR U30496 ( .A(n30042), .B(n30041), .Z(n30085) );
  NANDN U30497 ( .A(n29873), .B(n29872), .Z(n29877) );
  NAND U30498 ( .A(n29875), .B(n29874), .Z(n29876) );
  NAND U30499 ( .A(n29877), .B(n29876), .Z(n30030) );
  NANDN U30500 ( .A(n29879), .B(n29878), .Z(n29883) );
  NAND U30501 ( .A(n29881), .B(n29880), .Z(n29882) );
  NAND U30502 ( .A(n29883), .B(n29882), .Z(n30028) );
  OR U30503 ( .A(n29885), .B(n29884), .Z(n29889) );
  NANDN U30504 ( .A(n29887), .B(n29886), .Z(n29888) );
  NAND U30505 ( .A(n29889), .B(n29888), .Z(n30027) );
  XNOR U30506 ( .A(n30030), .B(n30029), .Z(n30086) );
  XNOR U30507 ( .A(n30085), .B(n30086), .Z(n30087) );
  NANDN U30508 ( .A(n29891), .B(n29890), .Z(n29895) );
  OR U30509 ( .A(n29893), .B(n29892), .Z(n29894) );
  AND U30510 ( .A(n29895), .B(n29894), .Z(n30088) );
  XOR U30511 ( .A(n30087), .B(n30088), .Z(n30105) );
  NANDN U30512 ( .A(n29901), .B(n29900), .Z(n29905) );
  NANDN U30513 ( .A(n29903), .B(n29902), .Z(n29904) );
  NAND U30514 ( .A(n29905), .B(n29904), .Z(n30094) );
  NANDN U30515 ( .A(n29911), .B(n29910), .Z(n29915) );
  NAND U30516 ( .A(n29913), .B(n29912), .Z(n29914) );
  NAND U30517 ( .A(n29915), .B(n29914), .Z(n30033) );
  NANDN U30518 ( .A(n29917), .B(n29916), .Z(n29921) );
  NAND U30519 ( .A(n29919), .B(n29918), .Z(n29920) );
  AND U30520 ( .A(n29921), .B(n29920), .Z(n30034) );
  XNOR U30521 ( .A(n30033), .B(n30034), .Z(n30035) );
  XOR U30522 ( .A(n1052), .B(a[206]), .Z(n30061) );
  NANDN U30523 ( .A(n30061), .B(n36925), .Z(n29924) );
  NAND U30524 ( .A(n36926), .B(n29922), .Z(n29923) );
  NAND U30525 ( .A(n29924), .B(n29923), .Z(n30019) );
  XNOR U30526 ( .A(n1054), .B(a[200]), .Z(n30058) );
  NANDN U30527 ( .A(n37665), .B(n30058), .Z(n29927) );
  NANDN U30528 ( .A(n29925), .B(n37604), .Z(n29926) );
  NAND U30529 ( .A(n29927), .B(n29926), .Z(n30017) );
  XOR U30530 ( .A(n1056), .B(a[194]), .Z(n30055) );
  NANDN U30531 ( .A(n30055), .B(n38101), .Z(n29930) );
  NAND U30532 ( .A(n38102), .B(n29928), .Z(n29929) );
  NAND U30533 ( .A(n29930), .B(n29929), .Z(n30018) );
  XNOR U30534 ( .A(n30017), .B(n30018), .Z(n30020) );
  XOR U30535 ( .A(n30019), .B(n30020), .Z(n30008) );
  XOR U30536 ( .A(b[11]), .B(n33130), .Z(n30064) );
  OR U30537 ( .A(n30064), .B(n37311), .Z(n29933) );
  NANDN U30538 ( .A(n29931), .B(n37218), .Z(n29932) );
  NAND U30539 ( .A(n29933), .B(n29932), .Z(n30006) );
  XOR U30540 ( .A(n1053), .B(a[202]), .Z(n30067) );
  NANDN U30541 ( .A(n30067), .B(n37424), .Z(n29936) );
  NANDN U30542 ( .A(n29934), .B(n37425), .Z(n29935) );
  AND U30543 ( .A(n29936), .B(n29935), .Z(n30005) );
  XNOR U30544 ( .A(n30006), .B(n30005), .Z(n30007) );
  XNOR U30545 ( .A(n30008), .B(n30007), .Z(n30024) );
  NANDN U30546 ( .A(n1049), .B(a[214]), .Z(n29937) );
  XNOR U30547 ( .A(b[1]), .B(n29937), .Z(n29939) );
  NANDN U30548 ( .A(b[0]), .B(a[213]), .Z(n29938) );
  AND U30549 ( .A(n29939), .B(n29938), .Z(n29983) );
  NAND U30550 ( .A(n38490), .B(n29940), .Z(n29942) );
  XNOR U30551 ( .A(n1058), .B(a[186]), .Z(n30073) );
  NANDN U30552 ( .A(n1048), .B(n30073), .Z(n29941) );
  NAND U30553 ( .A(n29942), .B(n29941), .Z(n29981) );
  NANDN U30554 ( .A(n1059), .B(a[182]), .Z(n29982) );
  XNOR U30555 ( .A(n29981), .B(n29982), .Z(n29984) );
  XNOR U30556 ( .A(n29983), .B(n29984), .Z(n30022) );
  NANDN U30557 ( .A(n29943), .B(n38205), .Z(n29945) );
  XNOR U30558 ( .A(b[23]), .B(a[192]), .Z(n30076) );
  OR U30559 ( .A(n30076), .B(n38268), .Z(n29944) );
  NAND U30560 ( .A(n29945), .B(n29944), .Z(n30046) );
  XOR U30561 ( .A(b[7]), .B(a[208]), .Z(n30079) );
  NAND U30562 ( .A(n30079), .B(n36701), .Z(n29948) );
  NAND U30563 ( .A(n29946), .B(n36702), .Z(n29947) );
  NAND U30564 ( .A(n29948), .B(n29947), .Z(n30043) );
  XOR U30565 ( .A(b[25]), .B(a[190]), .Z(n30082) );
  NAND U30566 ( .A(n30082), .B(n38325), .Z(n29951) );
  NANDN U30567 ( .A(n29949), .B(n38326), .Z(n29950) );
  AND U30568 ( .A(n29951), .B(n29950), .Z(n30044) );
  XNOR U30569 ( .A(n30043), .B(n30044), .Z(n30045) );
  XOR U30570 ( .A(n30046), .B(n30045), .Z(n30021) );
  XOR U30571 ( .A(n30024), .B(n30023), .Z(n30036) );
  XOR U30572 ( .A(n30035), .B(n30036), .Z(n30091) );
  XOR U30573 ( .A(n30092), .B(n30091), .Z(n30093) );
  XNOR U30574 ( .A(n30094), .B(n30093), .Z(n30103) );
  XNOR U30575 ( .A(n30104), .B(n30103), .Z(n30106) );
  XNOR U30576 ( .A(n30105), .B(n30106), .Z(n30100) );
  XOR U30577 ( .A(n30099), .B(n30100), .Z(n29978) );
  NANDN U30578 ( .A(n29953), .B(n29952), .Z(n29957) );
  NAND U30579 ( .A(n29955), .B(n29954), .Z(n29956) );
  NAND U30580 ( .A(n29957), .B(n29956), .Z(n29975) );
  NANDN U30581 ( .A(n29959), .B(n29958), .Z(n29963) );
  OR U30582 ( .A(n29961), .B(n29960), .Z(n29962) );
  NAND U30583 ( .A(n29963), .B(n29962), .Z(n29976) );
  XNOR U30584 ( .A(n29975), .B(n29976), .Z(n29977) );
  XNOR U30585 ( .A(n29978), .B(n29977), .Z(n29970) );
  XNOR U30586 ( .A(n29969), .B(n29970), .Z(n29971) );
  XNOR U30587 ( .A(n29972), .B(n29971), .Z(n30109) );
  XNOR U30588 ( .A(n30109), .B(sreg[438]), .Z(n30111) );
  NAND U30589 ( .A(n29964), .B(sreg[437]), .Z(n29968) );
  OR U30590 ( .A(n29966), .B(n29965), .Z(n29967) );
  AND U30591 ( .A(n29968), .B(n29967), .Z(n30110) );
  XOR U30592 ( .A(n30111), .B(n30110), .Z(c[438]) );
  NANDN U30593 ( .A(n29970), .B(n29969), .Z(n29974) );
  NAND U30594 ( .A(n29972), .B(n29971), .Z(n29973) );
  NAND U30595 ( .A(n29974), .B(n29973), .Z(n30117) );
  NANDN U30596 ( .A(n29976), .B(n29975), .Z(n29980) );
  NAND U30597 ( .A(n29978), .B(n29977), .Z(n29979) );
  NAND U30598 ( .A(n29980), .B(n29979), .Z(n30115) );
  NANDN U30599 ( .A(n29982), .B(n29981), .Z(n29986) );
  NAND U30600 ( .A(n29984), .B(n29983), .Z(n29985) );
  NAND U30601 ( .A(n29986), .B(n29985), .Z(n30195) );
  XNOR U30602 ( .A(b[19]), .B(a[197]), .Z(n30142) );
  NANDN U30603 ( .A(n30142), .B(n37934), .Z(n29989) );
  NANDN U30604 ( .A(n29987), .B(n37935), .Z(n29988) );
  NAND U30605 ( .A(n29989), .B(n29988), .Z(n30205) );
  XNOR U30606 ( .A(b[27]), .B(a[189]), .Z(n30145) );
  NANDN U30607 ( .A(n30145), .B(n38423), .Z(n29992) );
  NAND U30608 ( .A(n29990), .B(n38424), .Z(n29991) );
  NAND U30609 ( .A(n29992), .B(n29991), .Z(n30202) );
  XNOR U30610 ( .A(b[5]), .B(a[211]), .Z(n30148) );
  NANDN U30611 ( .A(n30148), .B(n36587), .Z(n29995) );
  NANDN U30612 ( .A(n29993), .B(n36588), .Z(n29994) );
  AND U30613 ( .A(n29995), .B(n29994), .Z(n30203) );
  XNOR U30614 ( .A(n30202), .B(n30203), .Z(n30204) );
  XNOR U30615 ( .A(n30205), .B(n30204), .Z(n30193) );
  NANDN U30616 ( .A(n29996), .B(n37762), .Z(n29998) );
  XOR U30617 ( .A(b[17]), .B(a[199]), .Z(n30151) );
  NAND U30618 ( .A(n30151), .B(n37764), .Z(n29997) );
  NAND U30619 ( .A(n29998), .B(n29997), .Z(n30169) );
  XNOR U30620 ( .A(b[31]), .B(a[185]), .Z(n30154) );
  NANDN U30621 ( .A(n30154), .B(n38552), .Z(n30001) );
  NANDN U30622 ( .A(n29999), .B(n38553), .Z(n30000) );
  NAND U30623 ( .A(n30001), .B(n30000), .Z(n30166) );
  OR U30624 ( .A(n30002), .B(n36105), .Z(n30004) );
  XNOR U30625 ( .A(b[3]), .B(a[213]), .Z(n30157) );
  NANDN U30626 ( .A(n30157), .B(n36107), .Z(n30003) );
  AND U30627 ( .A(n30004), .B(n30003), .Z(n30167) );
  XNOR U30628 ( .A(n30166), .B(n30167), .Z(n30168) );
  XOR U30629 ( .A(n30169), .B(n30168), .Z(n30192) );
  XNOR U30630 ( .A(n30193), .B(n30192), .Z(n30194) );
  XNOR U30631 ( .A(n30195), .B(n30194), .Z(n30133) );
  NANDN U30632 ( .A(n30006), .B(n30005), .Z(n30010) );
  NAND U30633 ( .A(n30008), .B(n30007), .Z(n30009) );
  NAND U30634 ( .A(n30010), .B(n30009), .Z(n30184) );
  NANDN U30635 ( .A(n30012), .B(n30011), .Z(n30016) );
  NAND U30636 ( .A(n30014), .B(n30013), .Z(n30015) );
  NAND U30637 ( .A(n30016), .B(n30015), .Z(n30183) );
  XNOR U30638 ( .A(n30183), .B(n30182), .Z(n30185) );
  XOR U30639 ( .A(n30184), .B(n30185), .Z(n30132) );
  XOR U30640 ( .A(n30133), .B(n30132), .Z(n30134) );
  NANDN U30641 ( .A(n30022), .B(n30021), .Z(n30026) );
  NAND U30642 ( .A(n30024), .B(n30023), .Z(n30025) );
  NAND U30643 ( .A(n30026), .B(n30025), .Z(n30135) );
  XNOR U30644 ( .A(n30134), .B(n30135), .Z(n30246) );
  OR U30645 ( .A(n30028), .B(n30027), .Z(n30032) );
  NAND U30646 ( .A(n30030), .B(n30029), .Z(n30031) );
  NAND U30647 ( .A(n30032), .B(n30031), .Z(n30245) );
  NANDN U30648 ( .A(n30034), .B(n30033), .Z(n30038) );
  NAND U30649 ( .A(n30036), .B(n30035), .Z(n30037) );
  NAND U30650 ( .A(n30038), .B(n30037), .Z(n30128) );
  NANDN U30651 ( .A(n30044), .B(n30043), .Z(n30048) );
  NAND U30652 ( .A(n30046), .B(n30045), .Z(n30047) );
  NAND U30653 ( .A(n30048), .B(n30047), .Z(n30186) );
  NANDN U30654 ( .A(n30050), .B(n30049), .Z(n30054) );
  NAND U30655 ( .A(n30052), .B(n30051), .Z(n30053) );
  AND U30656 ( .A(n30054), .B(n30053), .Z(n30187) );
  XNOR U30657 ( .A(n30186), .B(n30187), .Z(n30188) );
  XOR U30658 ( .A(n1056), .B(a[195]), .Z(n30208) );
  NANDN U30659 ( .A(n30208), .B(n38101), .Z(n30057) );
  NANDN U30660 ( .A(n30055), .B(n38102), .Z(n30056) );
  NAND U30661 ( .A(n30057), .B(n30056), .Z(n30178) );
  XOR U30662 ( .A(b[15]), .B(n32687), .Z(n30211) );
  OR U30663 ( .A(n30211), .B(n37665), .Z(n30060) );
  NAND U30664 ( .A(n30058), .B(n37604), .Z(n30059) );
  AND U30665 ( .A(n30060), .B(n30059), .Z(n30179) );
  XNOR U30666 ( .A(n30178), .B(n30179), .Z(n30181) );
  XOR U30667 ( .A(n1052), .B(a[207]), .Z(n30214) );
  NANDN U30668 ( .A(n30214), .B(n36925), .Z(n30063) );
  NANDN U30669 ( .A(n30061), .B(n36926), .Z(n30062) );
  NAND U30670 ( .A(n30063), .B(n30062), .Z(n30180) );
  XNOR U30671 ( .A(n30181), .B(n30180), .Z(n30174) );
  XNOR U30672 ( .A(b[11]), .B(a[205]), .Z(n30217) );
  OR U30673 ( .A(n30217), .B(n37311), .Z(n30066) );
  NANDN U30674 ( .A(n30064), .B(n37218), .Z(n30065) );
  NAND U30675 ( .A(n30066), .B(n30065), .Z(n30173) );
  XOR U30676 ( .A(n1053), .B(a[203]), .Z(n30220) );
  NANDN U30677 ( .A(n30220), .B(n37424), .Z(n30069) );
  NANDN U30678 ( .A(n30067), .B(n37425), .Z(n30068) );
  NAND U30679 ( .A(n30069), .B(n30068), .Z(n30172) );
  XNOR U30680 ( .A(n30173), .B(n30172), .Z(n30175) );
  XNOR U30681 ( .A(n30174), .B(n30175), .Z(n30163) );
  NANDN U30682 ( .A(n1049), .B(a[215]), .Z(n30070) );
  XNOR U30683 ( .A(b[1]), .B(n30070), .Z(n30072) );
  NANDN U30684 ( .A(b[0]), .B(a[214]), .Z(n30071) );
  AND U30685 ( .A(n30072), .B(n30071), .Z(n30138) );
  NAND U30686 ( .A(n38490), .B(n30073), .Z(n30075) );
  XNOR U30687 ( .A(n1058), .B(a[187]), .Z(n30223) );
  NANDN U30688 ( .A(n1048), .B(n30223), .Z(n30074) );
  NAND U30689 ( .A(n30075), .B(n30074), .Z(n30136) );
  NANDN U30690 ( .A(n1059), .B(a[183]), .Z(n30137) );
  XNOR U30691 ( .A(n30136), .B(n30137), .Z(n30139) );
  XNOR U30692 ( .A(n30138), .B(n30139), .Z(n30161) );
  NANDN U30693 ( .A(n30076), .B(n38205), .Z(n30078) );
  XOR U30694 ( .A(b[23]), .B(n31508), .Z(n30229) );
  OR U30695 ( .A(n30229), .B(n38268), .Z(n30077) );
  NAND U30696 ( .A(n30078), .B(n30077), .Z(n30199) );
  XOR U30697 ( .A(b[7]), .B(a[209]), .Z(n30232) );
  NAND U30698 ( .A(n30232), .B(n36701), .Z(n30081) );
  NAND U30699 ( .A(n30079), .B(n36702), .Z(n30080) );
  NAND U30700 ( .A(n30081), .B(n30080), .Z(n30196) );
  XOR U30701 ( .A(b[25]), .B(a[191]), .Z(n30235) );
  NAND U30702 ( .A(n30235), .B(n38325), .Z(n30084) );
  NAND U30703 ( .A(n30082), .B(n38326), .Z(n30083) );
  AND U30704 ( .A(n30084), .B(n30083), .Z(n30197) );
  XNOR U30705 ( .A(n30196), .B(n30197), .Z(n30198) );
  XOR U30706 ( .A(n30199), .B(n30198), .Z(n30160) );
  XOR U30707 ( .A(n30163), .B(n30162), .Z(n30189) );
  XNOR U30708 ( .A(n30188), .B(n30189), .Z(n30126) );
  XNOR U30709 ( .A(n30127), .B(n30126), .Z(n30129) );
  XNOR U30710 ( .A(n30128), .B(n30129), .Z(n30244) );
  XOR U30711 ( .A(n30245), .B(n30244), .Z(n30247) );
  NANDN U30712 ( .A(n30086), .B(n30085), .Z(n30090) );
  NAND U30713 ( .A(n30088), .B(n30087), .Z(n30089) );
  NAND U30714 ( .A(n30090), .B(n30089), .Z(n30238) );
  NAND U30715 ( .A(n30092), .B(n30091), .Z(n30096) );
  NAND U30716 ( .A(n30094), .B(n30093), .Z(n30095) );
  NAND U30717 ( .A(n30096), .B(n30095), .Z(n30239) );
  XNOR U30718 ( .A(n30238), .B(n30239), .Z(n30240) );
  XOR U30719 ( .A(n30241), .B(n30240), .Z(n30122) );
  NANDN U30720 ( .A(n30098), .B(n30097), .Z(n30102) );
  NANDN U30721 ( .A(n30100), .B(n30099), .Z(n30101) );
  NAND U30722 ( .A(n30102), .B(n30101), .Z(n30121) );
  OR U30723 ( .A(n30104), .B(n30103), .Z(n30108) );
  OR U30724 ( .A(n30106), .B(n30105), .Z(n30107) );
  AND U30725 ( .A(n30108), .B(n30107), .Z(n30120) );
  XNOR U30726 ( .A(n30121), .B(n30120), .Z(n30123) );
  XOR U30727 ( .A(n30122), .B(n30123), .Z(n30114) );
  XOR U30728 ( .A(n30115), .B(n30114), .Z(n30116) );
  XNOR U30729 ( .A(n30117), .B(n30116), .Z(n30250) );
  XNOR U30730 ( .A(n30250), .B(sreg[439]), .Z(n30252) );
  NAND U30731 ( .A(n30109), .B(sreg[438]), .Z(n30113) );
  OR U30732 ( .A(n30111), .B(n30110), .Z(n30112) );
  AND U30733 ( .A(n30113), .B(n30112), .Z(n30251) );
  XOR U30734 ( .A(n30252), .B(n30251), .Z(c[439]) );
  NAND U30735 ( .A(n30115), .B(n30114), .Z(n30119) );
  NAND U30736 ( .A(n30117), .B(n30116), .Z(n30118) );
  NAND U30737 ( .A(n30119), .B(n30118), .Z(n30258) );
  NANDN U30738 ( .A(n30121), .B(n30120), .Z(n30125) );
  NAND U30739 ( .A(n30123), .B(n30122), .Z(n30124) );
  NAND U30740 ( .A(n30125), .B(n30124), .Z(n30255) );
  NAND U30741 ( .A(n30127), .B(n30126), .Z(n30131) );
  NANDN U30742 ( .A(n30129), .B(n30128), .Z(n30130) );
  NAND U30743 ( .A(n30131), .B(n30130), .Z(n30381) );
  XNOR U30744 ( .A(n30381), .B(n30382), .Z(n30383) );
  NANDN U30745 ( .A(n30137), .B(n30136), .Z(n30141) );
  NAND U30746 ( .A(n30139), .B(n30138), .Z(n30140) );
  NAND U30747 ( .A(n30141), .B(n30140), .Z(n30280) );
  XOR U30748 ( .A(b[19]), .B(n32246), .Z(n30329) );
  NANDN U30749 ( .A(n30329), .B(n37934), .Z(n30144) );
  NANDN U30750 ( .A(n30142), .B(n37935), .Z(n30143) );
  NAND U30751 ( .A(n30144), .B(n30143), .Z(n30290) );
  XOR U30752 ( .A(b[27]), .B(a[190]), .Z(n30332) );
  NAND U30753 ( .A(n38423), .B(n30332), .Z(n30147) );
  NANDN U30754 ( .A(n30145), .B(n38424), .Z(n30146) );
  NAND U30755 ( .A(n30147), .B(n30146), .Z(n30287) );
  XNOR U30756 ( .A(b[5]), .B(a[212]), .Z(n30335) );
  NANDN U30757 ( .A(n30335), .B(n36587), .Z(n30150) );
  NANDN U30758 ( .A(n30148), .B(n36588), .Z(n30149) );
  AND U30759 ( .A(n30150), .B(n30149), .Z(n30288) );
  XNOR U30760 ( .A(n30287), .B(n30288), .Z(n30289) );
  XNOR U30761 ( .A(n30290), .B(n30289), .Z(n30278) );
  NAND U30762 ( .A(n30151), .B(n37762), .Z(n30153) );
  XOR U30763 ( .A(b[17]), .B(a[200]), .Z(n30338) );
  NAND U30764 ( .A(n30338), .B(n37764), .Z(n30152) );
  NAND U30765 ( .A(n30153), .B(n30152), .Z(n30356) );
  XNOR U30766 ( .A(b[31]), .B(a[186]), .Z(n30341) );
  NANDN U30767 ( .A(n30341), .B(n38552), .Z(n30156) );
  NANDN U30768 ( .A(n30154), .B(n38553), .Z(n30155) );
  NAND U30769 ( .A(n30156), .B(n30155), .Z(n30353) );
  OR U30770 ( .A(n30157), .B(n36105), .Z(n30159) );
  XNOR U30771 ( .A(b[3]), .B(a[214]), .Z(n30344) );
  NANDN U30772 ( .A(n30344), .B(n36107), .Z(n30158) );
  AND U30773 ( .A(n30159), .B(n30158), .Z(n30354) );
  XNOR U30774 ( .A(n30353), .B(n30354), .Z(n30355) );
  XOR U30775 ( .A(n30356), .B(n30355), .Z(n30277) );
  XNOR U30776 ( .A(n30278), .B(n30277), .Z(n30279) );
  XNOR U30777 ( .A(n30280), .B(n30279), .Z(n30375) );
  NANDN U30778 ( .A(n30161), .B(n30160), .Z(n30165) );
  NANDN U30779 ( .A(n30163), .B(n30162), .Z(n30164) );
  NAND U30780 ( .A(n30165), .B(n30164), .Z(n30376) );
  XNOR U30781 ( .A(n30375), .B(n30376), .Z(n30377) );
  NANDN U30782 ( .A(n30167), .B(n30166), .Z(n30171) );
  NAND U30783 ( .A(n30169), .B(n30168), .Z(n30170) );
  NAND U30784 ( .A(n30171), .B(n30170), .Z(n30270) );
  OR U30785 ( .A(n30173), .B(n30172), .Z(n30177) );
  NANDN U30786 ( .A(n30175), .B(n30174), .Z(n30176) );
  NAND U30787 ( .A(n30177), .B(n30176), .Z(n30268) );
  XNOR U30788 ( .A(n30268), .B(n30267), .Z(n30269) );
  XOR U30789 ( .A(n30270), .B(n30269), .Z(n30378) );
  XOR U30790 ( .A(n30377), .B(n30378), .Z(n30389) );
  NANDN U30791 ( .A(n30187), .B(n30186), .Z(n30191) );
  NANDN U30792 ( .A(n30189), .B(n30188), .Z(n30190) );
  NAND U30793 ( .A(n30191), .B(n30190), .Z(n30372) );
  NANDN U30794 ( .A(n30197), .B(n30196), .Z(n30201) );
  NAND U30795 ( .A(n30199), .B(n30198), .Z(n30200) );
  NAND U30796 ( .A(n30201), .B(n30200), .Z(n30271) );
  NANDN U30797 ( .A(n30203), .B(n30202), .Z(n30207) );
  NAND U30798 ( .A(n30205), .B(n30204), .Z(n30206) );
  AND U30799 ( .A(n30207), .B(n30206), .Z(n30272) );
  XNOR U30800 ( .A(n30271), .B(n30272), .Z(n30273) );
  XNOR U30801 ( .A(b[21]), .B(a[196]), .Z(n30299) );
  NANDN U30802 ( .A(n30299), .B(n38101), .Z(n30210) );
  NANDN U30803 ( .A(n30208), .B(n38102), .Z(n30209) );
  NAND U30804 ( .A(n30210), .B(n30209), .Z(n30365) );
  XNOR U30805 ( .A(b[15]), .B(a[202]), .Z(n30296) );
  OR U30806 ( .A(n30296), .B(n37665), .Z(n30213) );
  NANDN U30807 ( .A(n30211), .B(n37604), .Z(n30212) );
  AND U30808 ( .A(n30213), .B(n30212), .Z(n30366) );
  XNOR U30809 ( .A(n30365), .B(n30366), .Z(n30368) );
  XNOR U30810 ( .A(b[9]), .B(a[208]), .Z(n30293) );
  NANDN U30811 ( .A(n30293), .B(n36925), .Z(n30216) );
  NANDN U30812 ( .A(n30214), .B(n36926), .Z(n30215) );
  NAND U30813 ( .A(n30216), .B(n30215), .Z(n30367) );
  XNOR U30814 ( .A(n30368), .B(n30367), .Z(n30361) );
  XNOR U30815 ( .A(b[11]), .B(a[206]), .Z(n30302) );
  OR U30816 ( .A(n30302), .B(n37311), .Z(n30219) );
  NANDN U30817 ( .A(n30217), .B(n37218), .Z(n30218) );
  NAND U30818 ( .A(n30219), .B(n30218), .Z(n30360) );
  XOR U30819 ( .A(n1053), .B(a[204]), .Z(n30305) );
  NANDN U30820 ( .A(n30305), .B(n37424), .Z(n30222) );
  NANDN U30821 ( .A(n30220), .B(n37425), .Z(n30221) );
  NAND U30822 ( .A(n30222), .B(n30221), .Z(n30359) );
  XNOR U30823 ( .A(n30360), .B(n30359), .Z(n30362) );
  XNOR U30824 ( .A(n30361), .B(n30362), .Z(n30350) );
  NAND U30825 ( .A(n38490), .B(n30223), .Z(n30225) );
  XNOR U30826 ( .A(n1058), .B(a[188]), .Z(n30311) );
  NANDN U30827 ( .A(n1048), .B(n30311), .Z(n30224) );
  NAND U30828 ( .A(n30225), .B(n30224), .Z(n30323) );
  NANDN U30829 ( .A(n1059), .B(a[184]), .Z(n30324) );
  XNOR U30830 ( .A(n30323), .B(n30324), .Z(n30326) );
  NANDN U30831 ( .A(n1049), .B(a[216]), .Z(n30226) );
  XNOR U30832 ( .A(b[1]), .B(n30226), .Z(n30228) );
  IV U30833 ( .A(a[215]), .Z(n34725) );
  NANDN U30834 ( .A(n34725), .B(n1049), .Z(n30227) );
  AND U30835 ( .A(n30228), .B(n30227), .Z(n30325) );
  XNOR U30836 ( .A(n30326), .B(n30325), .Z(n30348) );
  NANDN U30837 ( .A(n30229), .B(n38205), .Z(n30231) );
  XOR U30838 ( .A(b[23]), .B(n31644), .Z(n30314) );
  OR U30839 ( .A(n30314), .B(n38268), .Z(n30230) );
  NAND U30840 ( .A(n30231), .B(n30230), .Z(n30284) );
  XOR U30841 ( .A(b[7]), .B(a[210]), .Z(n30317) );
  NAND U30842 ( .A(n30317), .B(n36701), .Z(n30234) );
  NAND U30843 ( .A(n30232), .B(n36702), .Z(n30233) );
  NAND U30844 ( .A(n30234), .B(n30233), .Z(n30281) );
  XOR U30845 ( .A(b[25]), .B(a[192]), .Z(n30320) );
  NAND U30846 ( .A(n30320), .B(n38325), .Z(n30237) );
  NAND U30847 ( .A(n30235), .B(n38326), .Z(n30236) );
  AND U30848 ( .A(n30237), .B(n30236), .Z(n30282) );
  XNOR U30849 ( .A(n30281), .B(n30282), .Z(n30283) );
  XOR U30850 ( .A(n30284), .B(n30283), .Z(n30347) );
  XOR U30851 ( .A(n30350), .B(n30349), .Z(n30274) );
  XNOR U30852 ( .A(n30273), .B(n30274), .Z(n30369) );
  XOR U30853 ( .A(n30370), .B(n30369), .Z(n30371) );
  XNOR U30854 ( .A(n30372), .B(n30371), .Z(n30387) );
  XNOR U30855 ( .A(n30388), .B(n30387), .Z(n30390) );
  XNOR U30856 ( .A(n30389), .B(n30390), .Z(n30384) );
  XOR U30857 ( .A(n30383), .B(n30384), .Z(n30264) );
  NANDN U30858 ( .A(n30239), .B(n30238), .Z(n30243) );
  NAND U30859 ( .A(n30241), .B(n30240), .Z(n30242) );
  NAND U30860 ( .A(n30243), .B(n30242), .Z(n30261) );
  NANDN U30861 ( .A(n30245), .B(n30244), .Z(n30249) );
  OR U30862 ( .A(n30247), .B(n30246), .Z(n30248) );
  NAND U30863 ( .A(n30249), .B(n30248), .Z(n30262) );
  XNOR U30864 ( .A(n30261), .B(n30262), .Z(n30263) );
  XNOR U30865 ( .A(n30264), .B(n30263), .Z(n30256) );
  XNOR U30866 ( .A(n30255), .B(n30256), .Z(n30257) );
  XNOR U30867 ( .A(n30258), .B(n30257), .Z(n30393) );
  XNOR U30868 ( .A(n30393), .B(sreg[440]), .Z(n30395) );
  NAND U30869 ( .A(n30250), .B(sreg[439]), .Z(n30254) );
  OR U30870 ( .A(n30252), .B(n30251), .Z(n30253) );
  AND U30871 ( .A(n30254), .B(n30253), .Z(n30394) );
  XOR U30872 ( .A(n30395), .B(n30394), .Z(c[440]) );
  NANDN U30873 ( .A(n30256), .B(n30255), .Z(n30260) );
  NAND U30874 ( .A(n30258), .B(n30257), .Z(n30259) );
  NAND U30875 ( .A(n30260), .B(n30259), .Z(n30401) );
  NANDN U30876 ( .A(n30262), .B(n30261), .Z(n30266) );
  NAND U30877 ( .A(n30264), .B(n30263), .Z(n30265) );
  NAND U30878 ( .A(n30266), .B(n30265), .Z(n30399) );
  NANDN U30879 ( .A(n30272), .B(n30271), .Z(n30276) );
  NANDN U30880 ( .A(n30274), .B(n30273), .Z(n30275) );
  NAND U30881 ( .A(n30276), .B(n30275), .Z(n30515) );
  NANDN U30882 ( .A(n30282), .B(n30281), .Z(n30286) );
  NAND U30883 ( .A(n30284), .B(n30283), .Z(n30285) );
  NAND U30884 ( .A(n30286), .B(n30285), .Z(n30460) );
  NANDN U30885 ( .A(n30288), .B(n30287), .Z(n30292) );
  NAND U30886 ( .A(n30290), .B(n30289), .Z(n30291) );
  AND U30887 ( .A(n30292), .B(n30291), .Z(n30461) );
  XNOR U30888 ( .A(n30460), .B(n30461), .Z(n30462) );
  XNOR U30889 ( .A(b[9]), .B(a[209]), .Z(n30482) );
  NANDN U30890 ( .A(n30482), .B(n36925), .Z(n30295) );
  NANDN U30891 ( .A(n30293), .B(n36926), .Z(n30294) );
  NAND U30892 ( .A(n30295), .B(n30294), .Z(n30446) );
  XNOR U30893 ( .A(b[15]), .B(a[203]), .Z(n30485) );
  OR U30894 ( .A(n30485), .B(n37665), .Z(n30298) );
  NANDN U30895 ( .A(n30296), .B(n37604), .Z(n30297) );
  AND U30896 ( .A(n30298), .B(n30297), .Z(n30444) );
  XNOR U30897 ( .A(b[21]), .B(a[197]), .Z(n30488) );
  NANDN U30898 ( .A(n30488), .B(n38101), .Z(n30301) );
  NANDN U30899 ( .A(n30299), .B(n38102), .Z(n30300) );
  AND U30900 ( .A(n30301), .B(n30300), .Z(n30445) );
  XOR U30901 ( .A(n30446), .B(n30447), .Z(n30435) );
  XNOR U30902 ( .A(b[11]), .B(a[207]), .Z(n30491) );
  OR U30903 ( .A(n30491), .B(n37311), .Z(n30304) );
  NANDN U30904 ( .A(n30302), .B(n37218), .Z(n30303) );
  NAND U30905 ( .A(n30304), .B(n30303), .Z(n30433) );
  XOR U30906 ( .A(n1053), .B(a[205]), .Z(n30494) );
  NANDN U30907 ( .A(n30494), .B(n37424), .Z(n30307) );
  NANDN U30908 ( .A(n30305), .B(n37425), .Z(n30306) );
  AND U30909 ( .A(n30307), .B(n30306), .Z(n30432) );
  XNOR U30910 ( .A(n30433), .B(n30432), .Z(n30434) );
  XOR U30911 ( .A(n30435), .B(n30434), .Z(n30452) );
  ANDN U30912 ( .B(a[217]), .A(n1049), .Z(n30308) );
  XOR U30913 ( .A(b[1]), .B(n30308), .Z(n30310) );
  NANDN U30914 ( .A(b[0]), .B(a[216]), .Z(n30309) );
  NAND U30915 ( .A(n30310), .B(n30309), .Z(n30411) );
  NAND U30916 ( .A(n38490), .B(n30311), .Z(n30313) );
  XOR U30917 ( .A(n1058), .B(n30936), .Z(n30500) );
  NANDN U30918 ( .A(n1048), .B(n30500), .Z(n30312) );
  NAND U30919 ( .A(n30313), .B(n30312), .Z(n30408) );
  NANDN U30920 ( .A(n1059), .B(a[185]), .Z(n30409) );
  XNOR U30921 ( .A(n30408), .B(n30409), .Z(n30410) );
  XNOR U30922 ( .A(n30411), .B(n30410), .Z(n30450) );
  NANDN U30923 ( .A(n30314), .B(n38205), .Z(n30316) );
  XOR U30924 ( .A(b[23]), .B(n31434), .Z(n30503) );
  OR U30925 ( .A(n30503), .B(n38268), .Z(n30315) );
  NAND U30926 ( .A(n30316), .B(n30315), .Z(n30473) );
  XOR U30927 ( .A(b[7]), .B(a[211]), .Z(n30506) );
  NAND U30928 ( .A(n30506), .B(n36701), .Z(n30319) );
  NAND U30929 ( .A(n30317), .B(n36702), .Z(n30318) );
  NAND U30930 ( .A(n30319), .B(n30318), .Z(n30470) );
  XNOR U30931 ( .A(b[25]), .B(a[193]), .Z(n30509) );
  NANDN U30932 ( .A(n30509), .B(n38325), .Z(n30322) );
  NAND U30933 ( .A(n30320), .B(n38326), .Z(n30321) );
  AND U30934 ( .A(n30322), .B(n30321), .Z(n30471) );
  XNOR U30935 ( .A(n30470), .B(n30471), .Z(n30472) );
  XNOR U30936 ( .A(n30473), .B(n30472), .Z(n30451) );
  XOR U30937 ( .A(n30450), .B(n30451), .Z(n30453) );
  XNOR U30938 ( .A(n30452), .B(n30453), .Z(n30463) );
  XOR U30939 ( .A(n30462), .B(n30463), .Z(n30513) );
  XNOR U30940 ( .A(n30512), .B(n30513), .Z(n30514) );
  XOR U30941 ( .A(n30515), .B(n30514), .Z(n30523) );
  XNOR U30942 ( .A(n30522), .B(n30523), .Z(n30525) );
  NANDN U30943 ( .A(n30324), .B(n30323), .Z(n30328) );
  NAND U30944 ( .A(n30326), .B(n30325), .Z(n30327) );
  NAND U30945 ( .A(n30328), .B(n30327), .Z(n30469) );
  XNOR U30946 ( .A(b[19]), .B(a[199]), .Z(n30414) );
  NANDN U30947 ( .A(n30414), .B(n37934), .Z(n30331) );
  NANDN U30948 ( .A(n30329), .B(n37935), .Z(n30330) );
  NAND U30949 ( .A(n30331), .B(n30330), .Z(n30479) );
  XOR U30950 ( .A(b[27]), .B(a[191]), .Z(n30417) );
  NAND U30951 ( .A(n38423), .B(n30417), .Z(n30334) );
  NAND U30952 ( .A(n30332), .B(n38424), .Z(n30333) );
  NAND U30953 ( .A(n30334), .B(n30333), .Z(n30476) );
  XNOR U30954 ( .A(b[5]), .B(a[213]), .Z(n30420) );
  NANDN U30955 ( .A(n30420), .B(n36587), .Z(n30337) );
  NANDN U30956 ( .A(n30335), .B(n36588), .Z(n30336) );
  AND U30957 ( .A(n30337), .B(n30336), .Z(n30477) );
  XNOR U30958 ( .A(n30476), .B(n30477), .Z(n30478) );
  XNOR U30959 ( .A(n30479), .B(n30478), .Z(n30467) );
  NAND U30960 ( .A(n30338), .B(n37762), .Z(n30340) );
  XNOR U30961 ( .A(b[17]), .B(a[201]), .Z(n30423) );
  NANDN U30962 ( .A(n30423), .B(n37764), .Z(n30339) );
  NAND U30963 ( .A(n30340), .B(n30339), .Z(n30441) );
  XNOR U30964 ( .A(b[31]), .B(a[187]), .Z(n30426) );
  NANDN U30965 ( .A(n30426), .B(n38552), .Z(n30343) );
  NANDN U30966 ( .A(n30341), .B(n38553), .Z(n30342) );
  NAND U30967 ( .A(n30343), .B(n30342), .Z(n30438) );
  OR U30968 ( .A(n30344), .B(n36105), .Z(n30346) );
  XOR U30969 ( .A(b[3]), .B(n34725), .Z(n30429) );
  NANDN U30970 ( .A(n30429), .B(n36107), .Z(n30345) );
  AND U30971 ( .A(n30346), .B(n30345), .Z(n30439) );
  XNOR U30972 ( .A(n30438), .B(n30439), .Z(n30440) );
  XOR U30973 ( .A(n30441), .B(n30440), .Z(n30466) );
  XNOR U30974 ( .A(n30467), .B(n30466), .Z(n30468) );
  XNOR U30975 ( .A(n30469), .B(n30468), .Z(n30518) );
  NANDN U30976 ( .A(n30348), .B(n30347), .Z(n30352) );
  NANDN U30977 ( .A(n30350), .B(n30349), .Z(n30351) );
  NAND U30978 ( .A(n30352), .B(n30351), .Z(n30519) );
  XNOR U30979 ( .A(n30518), .B(n30519), .Z(n30520) );
  NANDN U30980 ( .A(n30354), .B(n30353), .Z(n30358) );
  NAND U30981 ( .A(n30356), .B(n30355), .Z(n30357) );
  NAND U30982 ( .A(n30358), .B(n30357), .Z(n30459) );
  OR U30983 ( .A(n30360), .B(n30359), .Z(n30364) );
  NANDN U30984 ( .A(n30362), .B(n30361), .Z(n30363) );
  NAND U30985 ( .A(n30364), .B(n30363), .Z(n30457) );
  XNOR U30986 ( .A(n30457), .B(n30456), .Z(n30458) );
  XOR U30987 ( .A(n30459), .B(n30458), .Z(n30521) );
  XOR U30988 ( .A(n30520), .B(n30521), .Z(n30524) );
  XOR U30989 ( .A(n30525), .B(n30524), .Z(n30529) );
  NAND U30990 ( .A(n30370), .B(n30369), .Z(n30374) );
  NAND U30991 ( .A(n30372), .B(n30371), .Z(n30373) );
  NAND U30992 ( .A(n30374), .B(n30373), .Z(n30526) );
  NANDN U30993 ( .A(n30376), .B(n30375), .Z(n30380) );
  NAND U30994 ( .A(n30378), .B(n30377), .Z(n30379) );
  NAND U30995 ( .A(n30380), .B(n30379), .Z(n30527) );
  XNOR U30996 ( .A(n30526), .B(n30527), .Z(n30528) );
  XNOR U30997 ( .A(n30529), .B(n30528), .Z(n30405) );
  NANDN U30998 ( .A(n30382), .B(n30381), .Z(n30386) );
  NANDN U30999 ( .A(n30384), .B(n30383), .Z(n30385) );
  NAND U31000 ( .A(n30386), .B(n30385), .Z(n30403) );
  OR U31001 ( .A(n30388), .B(n30387), .Z(n30392) );
  OR U31002 ( .A(n30390), .B(n30389), .Z(n30391) );
  AND U31003 ( .A(n30392), .B(n30391), .Z(n30402) );
  XNOR U31004 ( .A(n30403), .B(n30402), .Z(n30404) );
  XNOR U31005 ( .A(n30405), .B(n30404), .Z(n30398) );
  XOR U31006 ( .A(n30399), .B(n30398), .Z(n30400) );
  XNOR U31007 ( .A(n30401), .B(n30400), .Z(n30532) );
  XNOR U31008 ( .A(n30532), .B(sreg[441]), .Z(n30534) );
  NAND U31009 ( .A(n30393), .B(sreg[440]), .Z(n30397) );
  OR U31010 ( .A(n30395), .B(n30394), .Z(n30396) );
  AND U31011 ( .A(n30397), .B(n30396), .Z(n30533) );
  XOR U31012 ( .A(n30534), .B(n30533), .Z(c[441]) );
  NANDN U31013 ( .A(n30403), .B(n30402), .Z(n30407) );
  NANDN U31014 ( .A(n30405), .B(n30404), .Z(n30406) );
  NAND U31015 ( .A(n30407), .B(n30406), .Z(n30538) );
  NANDN U31016 ( .A(n30409), .B(n30408), .Z(n30413) );
  NANDN U31017 ( .A(n30411), .B(n30410), .Z(n30412) );
  NAND U31018 ( .A(n30413), .B(n30412), .Z(n30620) );
  XNOR U31019 ( .A(b[19]), .B(a[200]), .Z(n30563) );
  NANDN U31020 ( .A(n30563), .B(n37934), .Z(n30416) );
  NANDN U31021 ( .A(n30414), .B(n37935), .Z(n30415) );
  NAND U31022 ( .A(n30416), .B(n30415), .Z(n30630) );
  XOR U31023 ( .A(b[27]), .B(a[192]), .Z(n30566) );
  NAND U31024 ( .A(n38423), .B(n30566), .Z(n30419) );
  NAND U31025 ( .A(n30417), .B(n38424), .Z(n30418) );
  NAND U31026 ( .A(n30419), .B(n30418), .Z(n30627) );
  XNOR U31027 ( .A(b[5]), .B(a[214]), .Z(n30569) );
  NANDN U31028 ( .A(n30569), .B(n36587), .Z(n30422) );
  NANDN U31029 ( .A(n30420), .B(n36588), .Z(n30421) );
  AND U31030 ( .A(n30422), .B(n30421), .Z(n30628) );
  XNOR U31031 ( .A(n30627), .B(n30628), .Z(n30629) );
  XNOR U31032 ( .A(n30630), .B(n30629), .Z(n30618) );
  NANDN U31033 ( .A(n30423), .B(n37762), .Z(n30425) );
  XOR U31034 ( .A(b[17]), .B(a[202]), .Z(n30572) );
  NAND U31035 ( .A(n30572), .B(n37764), .Z(n30424) );
  NAND U31036 ( .A(n30425), .B(n30424), .Z(n30590) );
  XNOR U31037 ( .A(b[31]), .B(a[188]), .Z(n30575) );
  NANDN U31038 ( .A(n30575), .B(n38552), .Z(n30428) );
  NANDN U31039 ( .A(n30426), .B(n38553), .Z(n30427) );
  NAND U31040 ( .A(n30428), .B(n30427), .Z(n30587) );
  OR U31041 ( .A(n30429), .B(n36105), .Z(n30431) );
  XNOR U31042 ( .A(b[3]), .B(a[216]), .Z(n30578) );
  NANDN U31043 ( .A(n30578), .B(n36107), .Z(n30430) );
  AND U31044 ( .A(n30431), .B(n30430), .Z(n30588) );
  XNOR U31045 ( .A(n30587), .B(n30588), .Z(n30589) );
  XOR U31046 ( .A(n30590), .B(n30589), .Z(n30617) );
  XNOR U31047 ( .A(n30618), .B(n30617), .Z(n30619) );
  XNOR U31048 ( .A(n30620), .B(n30619), .Z(n30663) );
  NANDN U31049 ( .A(n30433), .B(n30432), .Z(n30437) );
  NAND U31050 ( .A(n30435), .B(n30434), .Z(n30436) );
  NAND U31051 ( .A(n30437), .B(n30436), .Z(n30608) );
  NANDN U31052 ( .A(n30439), .B(n30438), .Z(n30443) );
  NAND U31053 ( .A(n30441), .B(n30440), .Z(n30442) );
  NAND U31054 ( .A(n30443), .B(n30442), .Z(n30606) );
  OR U31055 ( .A(n30445), .B(n30444), .Z(n30449) );
  NANDN U31056 ( .A(n30447), .B(n30446), .Z(n30448) );
  NAND U31057 ( .A(n30449), .B(n30448), .Z(n30605) );
  XNOR U31058 ( .A(n30608), .B(n30607), .Z(n30664) );
  XNOR U31059 ( .A(n30663), .B(n30664), .Z(n30665) );
  NANDN U31060 ( .A(n30451), .B(n30450), .Z(n30455) );
  OR U31061 ( .A(n30453), .B(n30452), .Z(n30454) );
  AND U31062 ( .A(n30455), .B(n30454), .Z(n30666) );
  XNOR U31063 ( .A(n30665), .B(n30666), .Z(n30550) );
  NANDN U31064 ( .A(n30461), .B(n30460), .Z(n30465) );
  NANDN U31065 ( .A(n30463), .B(n30462), .Z(n30464) );
  NAND U31066 ( .A(n30465), .B(n30464), .Z(n30672) );
  NANDN U31067 ( .A(n30471), .B(n30470), .Z(n30475) );
  NAND U31068 ( .A(n30473), .B(n30472), .Z(n30474) );
  NAND U31069 ( .A(n30475), .B(n30474), .Z(n30611) );
  NANDN U31070 ( .A(n30477), .B(n30476), .Z(n30481) );
  NAND U31071 ( .A(n30479), .B(n30478), .Z(n30480) );
  AND U31072 ( .A(n30481), .B(n30480), .Z(n30612) );
  XNOR U31073 ( .A(n30611), .B(n30612), .Z(n30613) );
  XNOR U31074 ( .A(n1052), .B(a[210]), .Z(n30633) );
  NAND U31075 ( .A(n36925), .B(n30633), .Z(n30484) );
  NANDN U31076 ( .A(n30482), .B(n36926), .Z(n30483) );
  NAND U31077 ( .A(n30484), .B(n30483), .Z(n30595) );
  XOR U31078 ( .A(b[15]), .B(n33130), .Z(n30636) );
  OR U31079 ( .A(n30636), .B(n37665), .Z(n30487) );
  NANDN U31080 ( .A(n30485), .B(n37604), .Z(n30486) );
  AND U31081 ( .A(n30487), .B(n30486), .Z(n30593) );
  XOR U31082 ( .A(n1056), .B(n32246), .Z(n30639) );
  NAND U31083 ( .A(n30639), .B(n38101), .Z(n30490) );
  NANDN U31084 ( .A(n30488), .B(n38102), .Z(n30489) );
  AND U31085 ( .A(n30490), .B(n30489), .Z(n30594) );
  XOR U31086 ( .A(n30595), .B(n30596), .Z(n30584) );
  XNOR U31087 ( .A(b[11]), .B(a[208]), .Z(n30642) );
  OR U31088 ( .A(n30642), .B(n37311), .Z(n30493) );
  NANDN U31089 ( .A(n30491), .B(n37218), .Z(n30492) );
  NAND U31090 ( .A(n30493), .B(n30492), .Z(n30582) );
  XOR U31091 ( .A(n1053), .B(a[206]), .Z(n30645) );
  NANDN U31092 ( .A(n30645), .B(n37424), .Z(n30496) );
  NANDN U31093 ( .A(n30494), .B(n37425), .Z(n30495) );
  AND U31094 ( .A(n30496), .B(n30495), .Z(n30581) );
  XNOR U31095 ( .A(n30582), .B(n30581), .Z(n30583) );
  XOR U31096 ( .A(n30584), .B(n30583), .Z(n30601) );
  NANDN U31097 ( .A(n1049), .B(a[218]), .Z(n30497) );
  XNOR U31098 ( .A(b[1]), .B(n30497), .Z(n30499) );
  IV U31099 ( .A(a[217]), .Z(n34670) );
  NANDN U31100 ( .A(n34670), .B(n1049), .Z(n30498) );
  AND U31101 ( .A(n30499), .B(n30498), .Z(n30559) );
  NAND U31102 ( .A(n38490), .B(n30500), .Z(n30502) );
  XNOR U31103 ( .A(n1058), .B(a[190]), .Z(n30651) );
  NANDN U31104 ( .A(n1048), .B(n30651), .Z(n30501) );
  NAND U31105 ( .A(n30502), .B(n30501), .Z(n30557) );
  NANDN U31106 ( .A(n1059), .B(a[186]), .Z(n30558) );
  XNOR U31107 ( .A(n30557), .B(n30558), .Z(n30560) );
  XOR U31108 ( .A(n30559), .B(n30560), .Z(n30599) );
  NANDN U31109 ( .A(n30503), .B(n38205), .Z(n30505) );
  XNOR U31110 ( .A(b[23]), .B(a[196]), .Z(n30654) );
  OR U31111 ( .A(n30654), .B(n38268), .Z(n30504) );
  NAND U31112 ( .A(n30505), .B(n30504), .Z(n30624) );
  XOR U31113 ( .A(b[7]), .B(a[212]), .Z(n30657) );
  NAND U31114 ( .A(n30657), .B(n36701), .Z(n30508) );
  NAND U31115 ( .A(n30506), .B(n36702), .Z(n30507) );
  NAND U31116 ( .A(n30508), .B(n30507), .Z(n30621) );
  XNOR U31117 ( .A(b[25]), .B(a[194]), .Z(n30660) );
  NANDN U31118 ( .A(n30660), .B(n38325), .Z(n30511) );
  NANDN U31119 ( .A(n30509), .B(n38326), .Z(n30510) );
  AND U31120 ( .A(n30511), .B(n30510), .Z(n30622) );
  XNOR U31121 ( .A(n30621), .B(n30622), .Z(n30623) );
  XNOR U31122 ( .A(n30624), .B(n30623), .Z(n30600) );
  XOR U31123 ( .A(n30599), .B(n30600), .Z(n30602) );
  XNOR U31124 ( .A(n30601), .B(n30602), .Z(n30614) );
  XOR U31125 ( .A(n30613), .B(n30614), .Z(n30670) );
  XNOR U31126 ( .A(n30669), .B(n30670), .Z(n30671) );
  XOR U31127 ( .A(n30672), .B(n30671), .Z(n30548) );
  XNOR U31128 ( .A(n30547), .B(n30548), .Z(n30549) );
  XNOR U31129 ( .A(n30550), .B(n30549), .Z(n30554) );
  NANDN U31130 ( .A(n30513), .B(n30512), .Z(n30517) );
  NAND U31131 ( .A(n30515), .B(n30514), .Z(n30516) );
  NAND U31132 ( .A(n30517), .B(n30516), .Z(n30551) );
  XNOR U31133 ( .A(n30551), .B(n30552), .Z(n30553) );
  XNOR U31134 ( .A(n30554), .B(n30553), .Z(n30544) );
  NANDN U31135 ( .A(n30527), .B(n30526), .Z(n30531) );
  NANDN U31136 ( .A(n30529), .B(n30528), .Z(n30530) );
  NAND U31137 ( .A(n30531), .B(n30530), .Z(n30542) );
  XNOR U31138 ( .A(n30541), .B(n30542), .Z(n30543) );
  XNOR U31139 ( .A(n30544), .B(n30543), .Z(n30537) );
  XOR U31140 ( .A(n30538), .B(n30537), .Z(n30539) );
  XNOR U31141 ( .A(n30540), .B(n30539), .Z(n30675) );
  XNOR U31142 ( .A(n30675), .B(sreg[442]), .Z(n30677) );
  NAND U31143 ( .A(n30532), .B(sreg[441]), .Z(n30536) );
  OR U31144 ( .A(n30534), .B(n30533), .Z(n30535) );
  AND U31145 ( .A(n30536), .B(n30535), .Z(n30676) );
  XOR U31146 ( .A(n30677), .B(n30676), .Z(c[442]) );
  NANDN U31147 ( .A(n30542), .B(n30541), .Z(n30546) );
  NANDN U31148 ( .A(n30544), .B(n30543), .Z(n30545) );
  NAND U31149 ( .A(n30546), .B(n30545), .Z(n30681) );
  NANDN U31150 ( .A(n30552), .B(n30551), .Z(n30556) );
  NANDN U31151 ( .A(n30554), .B(n30553), .Z(n30555) );
  NAND U31152 ( .A(n30556), .B(n30555), .Z(n30687) );
  XNOR U31153 ( .A(n30686), .B(n30687), .Z(n30688) );
  NANDN U31154 ( .A(n30558), .B(n30557), .Z(n30562) );
  NAND U31155 ( .A(n30560), .B(n30559), .Z(n30561) );
  NAND U31156 ( .A(n30562), .B(n30561), .Z(n30765) );
  XOR U31157 ( .A(b[19]), .B(n32687), .Z(n30710) );
  NANDN U31158 ( .A(n30710), .B(n37934), .Z(n30565) );
  NANDN U31159 ( .A(n30563), .B(n37935), .Z(n30564) );
  NAND U31160 ( .A(n30565), .B(n30564), .Z(n30775) );
  XNOR U31161 ( .A(b[27]), .B(a[193]), .Z(n30713) );
  NANDN U31162 ( .A(n30713), .B(n38423), .Z(n30568) );
  NAND U31163 ( .A(n30566), .B(n38424), .Z(n30567) );
  NAND U31164 ( .A(n30568), .B(n30567), .Z(n30772) );
  XOR U31165 ( .A(b[5]), .B(n34725), .Z(n30716) );
  NANDN U31166 ( .A(n30716), .B(n36587), .Z(n30571) );
  NANDN U31167 ( .A(n30569), .B(n36588), .Z(n30570) );
  AND U31168 ( .A(n30571), .B(n30570), .Z(n30773) );
  XNOR U31169 ( .A(n30772), .B(n30773), .Z(n30774) );
  XNOR U31170 ( .A(n30775), .B(n30774), .Z(n30763) );
  NAND U31171 ( .A(n30572), .B(n37762), .Z(n30574) );
  XOR U31172 ( .A(b[17]), .B(a[203]), .Z(n30719) );
  NAND U31173 ( .A(n30719), .B(n37764), .Z(n30573) );
  NAND U31174 ( .A(n30574), .B(n30573), .Z(n30737) );
  XOR U31175 ( .A(b[31]), .B(n30936), .Z(n30722) );
  NANDN U31176 ( .A(n30722), .B(n38552), .Z(n30577) );
  NANDN U31177 ( .A(n30575), .B(n38553), .Z(n30576) );
  NAND U31178 ( .A(n30577), .B(n30576), .Z(n30734) );
  OR U31179 ( .A(n30578), .B(n36105), .Z(n30580) );
  XOR U31180 ( .A(b[3]), .B(n34670), .Z(n30725) );
  NANDN U31181 ( .A(n30725), .B(n36107), .Z(n30579) );
  AND U31182 ( .A(n30580), .B(n30579), .Z(n30735) );
  XNOR U31183 ( .A(n30734), .B(n30735), .Z(n30736) );
  XOR U31184 ( .A(n30737), .B(n30736), .Z(n30762) );
  XNOR U31185 ( .A(n30763), .B(n30762), .Z(n30764) );
  XNOR U31186 ( .A(n30765), .B(n30764), .Z(n30808) );
  NANDN U31187 ( .A(n30582), .B(n30581), .Z(n30586) );
  NAND U31188 ( .A(n30584), .B(n30583), .Z(n30585) );
  NAND U31189 ( .A(n30586), .B(n30585), .Z(n30753) );
  NANDN U31190 ( .A(n30588), .B(n30587), .Z(n30592) );
  NAND U31191 ( .A(n30590), .B(n30589), .Z(n30591) );
  NAND U31192 ( .A(n30592), .B(n30591), .Z(n30751) );
  OR U31193 ( .A(n30594), .B(n30593), .Z(n30598) );
  NANDN U31194 ( .A(n30596), .B(n30595), .Z(n30597) );
  NAND U31195 ( .A(n30598), .B(n30597), .Z(n30750) );
  XNOR U31196 ( .A(n30753), .B(n30752), .Z(n30809) );
  XOR U31197 ( .A(n30808), .B(n30809), .Z(n30811) );
  NANDN U31198 ( .A(n30600), .B(n30599), .Z(n30604) );
  OR U31199 ( .A(n30602), .B(n30601), .Z(n30603) );
  NAND U31200 ( .A(n30604), .B(n30603), .Z(n30810) );
  XOR U31201 ( .A(n30811), .B(n30810), .Z(n30700) );
  OR U31202 ( .A(n30606), .B(n30605), .Z(n30610) );
  NAND U31203 ( .A(n30608), .B(n30607), .Z(n30609) );
  NAND U31204 ( .A(n30610), .B(n30609), .Z(n30699) );
  NANDN U31205 ( .A(n30612), .B(n30611), .Z(n30616) );
  NANDN U31206 ( .A(n30614), .B(n30613), .Z(n30615) );
  NAND U31207 ( .A(n30616), .B(n30615), .Z(n30816) );
  NANDN U31208 ( .A(n30622), .B(n30621), .Z(n30626) );
  NAND U31209 ( .A(n30624), .B(n30623), .Z(n30625) );
  NAND U31210 ( .A(n30626), .B(n30625), .Z(n30756) );
  NANDN U31211 ( .A(n30628), .B(n30627), .Z(n30632) );
  NAND U31212 ( .A(n30630), .B(n30629), .Z(n30631) );
  AND U31213 ( .A(n30632), .B(n30631), .Z(n30757) );
  XNOR U31214 ( .A(n30756), .B(n30757), .Z(n30758) );
  XNOR U31215 ( .A(b[9]), .B(a[211]), .Z(n30778) );
  NANDN U31216 ( .A(n30778), .B(n36925), .Z(n30635) );
  NAND U31217 ( .A(n36926), .B(n30633), .Z(n30634) );
  NAND U31218 ( .A(n30635), .B(n30634), .Z(n30742) );
  XNOR U31219 ( .A(n1054), .B(a[205]), .Z(n30781) );
  NANDN U31220 ( .A(n37665), .B(n30781), .Z(n30638) );
  NANDN U31221 ( .A(n30636), .B(n37604), .Z(n30637) );
  NAND U31222 ( .A(n30638), .B(n30637), .Z(n30740) );
  XNOR U31223 ( .A(b[21]), .B(a[199]), .Z(n30784) );
  NANDN U31224 ( .A(n30784), .B(n38101), .Z(n30641) );
  NAND U31225 ( .A(n38102), .B(n30639), .Z(n30640) );
  NAND U31226 ( .A(n30641), .B(n30640), .Z(n30741) );
  XNOR U31227 ( .A(n30740), .B(n30741), .Z(n30743) );
  XOR U31228 ( .A(n30742), .B(n30743), .Z(n30731) );
  XNOR U31229 ( .A(b[11]), .B(a[209]), .Z(n30787) );
  OR U31230 ( .A(n30787), .B(n37311), .Z(n30644) );
  NANDN U31231 ( .A(n30642), .B(n37218), .Z(n30643) );
  NAND U31232 ( .A(n30644), .B(n30643), .Z(n30729) );
  XOR U31233 ( .A(n1053), .B(a[207]), .Z(n30790) );
  NANDN U31234 ( .A(n30790), .B(n37424), .Z(n30647) );
  NANDN U31235 ( .A(n30645), .B(n37425), .Z(n30646) );
  AND U31236 ( .A(n30647), .B(n30646), .Z(n30728) );
  XNOR U31237 ( .A(n30729), .B(n30728), .Z(n30730) );
  XNOR U31238 ( .A(n30731), .B(n30730), .Z(n30747) );
  NANDN U31239 ( .A(n1049), .B(a[219]), .Z(n30648) );
  XNOR U31240 ( .A(b[1]), .B(n30648), .Z(n30650) );
  NANDN U31241 ( .A(b[0]), .B(a[218]), .Z(n30649) );
  AND U31242 ( .A(n30650), .B(n30649), .Z(n30706) );
  NAND U31243 ( .A(n38490), .B(n30651), .Z(n30653) );
  XNOR U31244 ( .A(n1058), .B(a[191]), .Z(n30796) );
  NANDN U31245 ( .A(n1048), .B(n30796), .Z(n30652) );
  NAND U31246 ( .A(n30653), .B(n30652), .Z(n30704) );
  NANDN U31247 ( .A(n1059), .B(a[187]), .Z(n30705) );
  XNOR U31248 ( .A(n30704), .B(n30705), .Z(n30707) );
  XNOR U31249 ( .A(n30706), .B(n30707), .Z(n30745) );
  NANDN U31250 ( .A(n30654), .B(n38205), .Z(n30656) );
  XNOR U31251 ( .A(b[23]), .B(a[197]), .Z(n30799) );
  OR U31252 ( .A(n30799), .B(n38268), .Z(n30655) );
  NAND U31253 ( .A(n30656), .B(n30655), .Z(n30769) );
  XOR U31254 ( .A(b[7]), .B(a[213]), .Z(n30802) );
  NAND U31255 ( .A(n30802), .B(n36701), .Z(n30659) );
  NAND U31256 ( .A(n30657), .B(n36702), .Z(n30658) );
  NAND U31257 ( .A(n30659), .B(n30658), .Z(n30766) );
  XNOR U31258 ( .A(b[25]), .B(a[195]), .Z(n30805) );
  NANDN U31259 ( .A(n30805), .B(n38325), .Z(n30662) );
  NANDN U31260 ( .A(n30660), .B(n38326), .Z(n30661) );
  AND U31261 ( .A(n30662), .B(n30661), .Z(n30767) );
  XNOR U31262 ( .A(n30766), .B(n30767), .Z(n30768) );
  XOR U31263 ( .A(n30769), .B(n30768), .Z(n30744) );
  XOR U31264 ( .A(n30747), .B(n30746), .Z(n30759) );
  XOR U31265 ( .A(n30758), .B(n30759), .Z(n30814) );
  XNOR U31266 ( .A(n30815), .B(n30814), .Z(n30817) );
  XNOR U31267 ( .A(n30816), .B(n30817), .Z(n30698) );
  XOR U31268 ( .A(n30699), .B(n30698), .Z(n30701) );
  NANDN U31269 ( .A(n30664), .B(n30663), .Z(n30668) );
  NAND U31270 ( .A(n30666), .B(n30665), .Z(n30667) );
  NAND U31271 ( .A(n30668), .B(n30667), .Z(n30692) );
  NANDN U31272 ( .A(n30670), .B(n30669), .Z(n30674) );
  NAND U31273 ( .A(n30672), .B(n30671), .Z(n30673) );
  NAND U31274 ( .A(n30674), .B(n30673), .Z(n30693) );
  XNOR U31275 ( .A(n30692), .B(n30693), .Z(n30694) );
  XOR U31276 ( .A(n30695), .B(n30694), .Z(n30689) );
  XOR U31277 ( .A(n30688), .B(n30689), .Z(n30680) );
  XOR U31278 ( .A(n30681), .B(n30680), .Z(n30682) );
  XNOR U31279 ( .A(n30683), .B(n30682), .Z(n30820) );
  XNOR U31280 ( .A(n30820), .B(sreg[443]), .Z(n30822) );
  NAND U31281 ( .A(n30675), .B(sreg[442]), .Z(n30679) );
  OR U31282 ( .A(n30677), .B(n30676), .Z(n30678) );
  AND U31283 ( .A(n30679), .B(n30678), .Z(n30821) );
  XOR U31284 ( .A(n30822), .B(n30821), .Z(c[443]) );
  NAND U31285 ( .A(n30681), .B(n30680), .Z(n30685) );
  NAND U31286 ( .A(n30683), .B(n30682), .Z(n30684) );
  NAND U31287 ( .A(n30685), .B(n30684), .Z(n30828) );
  NANDN U31288 ( .A(n30687), .B(n30686), .Z(n30691) );
  NAND U31289 ( .A(n30689), .B(n30688), .Z(n30690) );
  NAND U31290 ( .A(n30691), .B(n30690), .Z(n30826) );
  NANDN U31291 ( .A(n30693), .B(n30692), .Z(n30697) );
  NAND U31292 ( .A(n30695), .B(n30694), .Z(n30696) );
  NAND U31293 ( .A(n30697), .B(n30696), .Z(n30831) );
  NANDN U31294 ( .A(n30699), .B(n30698), .Z(n30703) );
  OR U31295 ( .A(n30701), .B(n30700), .Z(n30702) );
  NAND U31296 ( .A(n30703), .B(n30702), .Z(n30832) );
  XNOR U31297 ( .A(n30831), .B(n30832), .Z(n30833) );
  NANDN U31298 ( .A(n30705), .B(n30704), .Z(n30709) );
  NAND U31299 ( .A(n30707), .B(n30706), .Z(n30708) );
  NAND U31300 ( .A(n30709), .B(n30708), .Z(n30908) );
  XNOR U31301 ( .A(b[19]), .B(a[202]), .Z(n30853) );
  NANDN U31302 ( .A(n30853), .B(n37934), .Z(n30712) );
  NANDN U31303 ( .A(n30710), .B(n37935), .Z(n30711) );
  NAND U31304 ( .A(n30712), .B(n30711), .Z(n30918) );
  XNOR U31305 ( .A(b[27]), .B(a[194]), .Z(n30856) );
  NANDN U31306 ( .A(n30856), .B(n38423), .Z(n30715) );
  NANDN U31307 ( .A(n30713), .B(n38424), .Z(n30714) );
  NAND U31308 ( .A(n30715), .B(n30714), .Z(n30915) );
  XNOR U31309 ( .A(b[5]), .B(a[216]), .Z(n30859) );
  NANDN U31310 ( .A(n30859), .B(n36587), .Z(n30718) );
  NANDN U31311 ( .A(n30716), .B(n36588), .Z(n30717) );
  AND U31312 ( .A(n30718), .B(n30717), .Z(n30916) );
  XNOR U31313 ( .A(n30915), .B(n30916), .Z(n30917) );
  XNOR U31314 ( .A(n30918), .B(n30917), .Z(n30906) );
  NAND U31315 ( .A(n30719), .B(n37762), .Z(n30721) );
  XNOR U31316 ( .A(b[17]), .B(a[204]), .Z(n30862) );
  NANDN U31317 ( .A(n30862), .B(n37764), .Z(n30720) );
  NAND U31318 ( .A(n30721), .B(n30720), .Z(n30880) );
  XNOR U31319 ( .A(b[31]), .B(a[190]), .Z(n30865) );
  NANDN U31320 ( .A(n30865), .B(n38552), .Z(n30724) );
  NANDN U31321 ( .A(n30722), .B(n38553), .Z(n30723) );
  NAND U31322 ( .A(n30724), .B(n30723), .Z(n30877) );
  OR U31323 ( .A(n30725), .B(n36105), .Z(n30727) );
  XNOR U31324 ( .A(b[3]), .B(a[218]), .Z(n30868) );
  NANDN U31325 ( .A(n30868), .B(n36107), .Z(n30726) );
  AND U31326 ( .A(n30727), .B(n30726), .Z(n30878) );
  XNOR U31327 ( .A(n30877), .B(n30878), .Z(n30879) );
  XOR U31328 ( .A(n30880), .B(n30879), .Z(n30905) );
  XNOR U31329 ( .A(n30906), .B(n30905), .Z(n30907) );
  XNOR U31330 ( .A(n30908), .B(n30907), .Z(n30844) );
  NANDN U31331 ( .A(n30729), .B(n30728), .Z(n30733) );
  NAND U31332 ( .A(n30731), .B(n30730), .Z(n30732) );
  NAND U31333 ( .A(n30733), .B(n30732), .Z(n30897) );
  NANDN U31334 ( .A(n30735), .B(n30734), .Z(n30739) );
  NAND U31335 ( .A(n30737), .B(n30736), .Z(n30738) );
  NAND U31336 ( .A(n30739), .B(n30738), .Z(n30896) );
  XNOR U31337 ( .A(n30896), .B(n30895), .Z(n30898) );
  XOR U31338 ( .A(n30897), .B(n30898), .Z(n30843) );
  XOR U31339 ( .A(n30844), .B(n30843), .Z(n30845) );
  NANDN U31340 ( .A(n30745), .B(n30744), .Z(n30749) );
  NAND U31341 ( .A(n30747), .B(n30746), .Z(n30748) );
  NAND U31342 ( .A(n30749), .B(n30748), .Z(n30846) );
  XNOR U31343 ( .A(n30845), .B(n30846), .Z(n30960) );
  OR U31344 ( .A(n30751), .B(n30750), .Z(n30755) );
  NAND U31345 ( .A(n30753), .B(n30752), .Z(n30754) );
  NAND U31346 ( .A(n30755), .B(n30754), .Z(n30959) );
  NANDN U31347 ( .A(n30757), .B(n30756), .Z(n30761) );
  NAND U31348 ( .A(n30759), .B(n30758), .Z(n30760) );
  NAND U31349 ( .A(n30761), .B(n30760), .Z(n30839) );
  NANDN U31350 ( .A(n30767), .B(n30766), .Z(n30771) );
  NAND U31351 ( .A(n30769), .B(n30768), .Z(n30770) );
  NAND U31352 ( .A(n30771), .B(n30770), .Z(n30899) );
  NANDN U31353 ( .A(n30773), .B(n30772), .Z(n30777) );
  NAND U31354 ( .A(n30775), .B(n30774), .Z(n30776) );
  AND U31355 ( .A(n30777), .B(n30776), .Z(n30900) );
  XNOR U31356 ( .A(n30899), .B(n30900), .Z(n30901) );
  XNOR U31357 ( .A(b[9]), .B(a[212]), .Z(n30921) );
  NANDN U31358 ( .A(n30921), .B(n36925), .Z(n30780) );
  NANDN U31359 ( .A(n30778), .B(n36926), .Z(n30779) );
  NAND U31360 ( .A(n30780), .B(n30779), .Z(n30885) );
  XNOR U31361 ( .A(b[15]), .B(a[206]), .Z(n30924) );
  OR U31362 ( .A(n30924), .B(n37665), .Z(n30783) );
  NAND U31363 ( .A(n30781), .B(n37604), .Z(n30782) );
  AND U31364 ( .A(n30783), .B(n30782), .Z(n30883) );
  XNOR U31365 ( .A(b[21]), .B(a[200]), .Z(n30927) );
  NANDN U31366 ( .A(n30927), .B(n38101), .Z(n30786) );
  NANDN U31367 ( .A(n30784), .B(n38102), .Z(n30785) );
  AND U31368 ( .A(n30786), .B(n30785), .Z(n30884) );
  XOR U31369 ( .A(n30885), .B(n30886), .Z(n30874) );
  XNOR U31370 ( .A(b[11]), .B(a[210]), .Z(n30930) );
  OR U31371 ( .A(n30930), .B(n37311), .Z(n30789) );
  NANDN U31372 ( .A(n30787), .B(n37218), .Z(n30788) );
  NAND U31373 ( .A(n30789), .B(n30788), .Z(n30872) );
  XOR U31374 ( .A(n1053), .B(a[208]), .Z(n30933) );
  NANDN U31375 ( .A(n30933), .B(n37424), .Z(n30792) );
  NANDN U31376 ( .A(n30790), .B(n37425), .Z(n30791) );
  AND U31377 ( .A(n30792), .B(n30791), .Z(n30871) );
  XNOR U31378 ( .A(n30872), .B(n30871), .Z(n30873) );
  XOR U31379 ( .A(n30874), .B(n30873), .Z(n30891) );
  NANDN U31380 ( .A(n1049), .B(a[220]), .Z(n30793) );
  XNOR U31381 ( .A(b[1]), .B(n30793), .Z(n30795) );
  NANDN U31382 ( .A(b[0]), .B(a[219]), .Z(n30794) );
  AND U31383 ( .A(n30795), .B(n30794), .Z(n30849) );
  NAND U31384 ( .A(n38490), .B(n30796), .Z(n30798) );
  XNOR U31385 ( .A(b[29]), .B(a[192]), .Z(n30937) );
  OR U31386 ( .A(n30937), .B(n1048), .Z(n30797) );
  NAND U31387 ( .A(n30798), .B(n30797), .Z(n30847) );
  NANDN U31388 ( .A(n1059), .B(a[188]), .Z(n30848) );
  XNOR U31389 ( .A(n30847), .B(n30848), .Z(n30850) );
  XOR U31390 ( .A(n30849), .B(n30850), .Z(n30889) );
  NANDN U31391 ( .A(n30799), .B(n38205), .Z(n30801) );
  XOR U31392 ( .A(b[23]), .B(n32246), .Z(n30943) );
  OR U31393 ( .A(n30943), .B(n38268), .Z(n30800) );
  NAND U31394 ( .A(n30801), .B(n30800), .Z(n30912) );
  XOR U31395 ( .A(b[7]), .B(a[214]), .Z(n30946) );
  NAND U31396 ( .A(n30946), .B(n36701), .Z(n30804) );
  NAND U31397 ( .A(n30802), .B(n36702), .Z(n30803) );
  NAND U31398 ( .A(n30804), .B(n30803), .Z(n30909) );
  XOR U31399 ( .A(b[25]), .B(a[196]), .Z(n30949) );
  NAND U31400 ( .A(n30949), .B(n38325), .Z(n30807) );
  NANDN U31401 ( .A(n30805), .B(n38326), .Z(n30806) );
  AND U31402 ( .A(n30807), .B(n30806), .Z(n30910) );
  XNOR U31403 ( .A(n30909), .B(n30910), .Z(n30911) );
  XNOR U31404 ( .A(n30912), .B(n30911), .Z(n30890) );
  XOR U31405 ( .A(n30889), .B(n30890), .Z(n30892) );
  XNOR U31406 ( .A(n30891), .B(n30892), .Z(n30902) );
  XNOR U31407 ( .A(n30901), .B(n30902), .Z(n30837) );
  XNOR U31408 ( .A(n30838), .B(n30837), .Z(n30840) );
  XNOR U31409 ( .A(n30839), .B(n30840), .Z(n30958) );
  XOR U31410 ( .A(n30959), .B(n30958), .Z(n30961) );
  NANDN U31411 ( .A(n30809), .B(n30808), .Z(n30813) );
  OR U31412 ( .A(n30811), .B(n30810), .Z(n30812) );
  NAND U31413 ( .A(n30813), .B(n30812), .Z(n30952) );
  NAND U31414 ( .A(n30815), .B(n30814), .Z(n30819) );
  NANDN U31415 ( .A(n30817), .B(n30816), .Z(n30818) );
  NAND U31416 ( .A(n30819), .B(n30818), .Z(n30953) );
  XNOR U31417 ( .A(n30952), .B(n30953), .Z(n30954) );
  XOR U31418 ( .A(n30955), .B(n30954), .Z(n30834) );
  XOR U31419 ( .A(n30833), .B(n30834), .Z(n30825) );
  XOR U31420 ( .A(n30826), .B(n30825), .Z(n30827) );
  XNOR U31421 ( .A(n30828), .B(n30827), .Z(n30964) );
  XNOR U31422 ( .A(n30964), .B(sreg[444]), .Z(n30966) );
  NAND U31423 ( .A(n30820), .B(sreg[443]), .Z(n30824) );
  OR U31424 ( .A(n30822), .B(n30821), .Z(n30823) );
  AND U31425 ( .A(n30824), .B(n30823), .Z(n30965) );
  XOR U31426 ( .A(n30966), .B(n30965), .Z(c[444]) );
  NAND U31427 ( .A(n30826), .B(n30825), .Z(n30830) );
  NAND U31428 ( .A(n30828), .B(n30827), .Z(n30829) );
  NAND U31429 ( .A(n30830), .B(n30829), .Z(n30972) );
  NANDN U31430 ( .A(n30832), .B(n30831), .Z(n30836) );
  NAND U31431 ( .A(n30834), .B(n30833), .Z(n30835) );
  NAND U31432 ( .A(n30836), .B(n30835), .Z(n30969) );
  NAND U31433 ( .A(n30838), .B(n30837), .Z(n30842) );
  NANDN U31434 ( .A(n30840), .B(n30839), .Z(n30841) );
  NAND U31435 ( .A(n30842), .B(n30841), .Z(n31101) );
  XNOR U31436 ( .A(n31101), .B(n31102), .Z(n31103) );
  NANDN U31437 ( .A(n30848), .B(n30847), .Z(n30852) );
  NAND U31438 ( .A(n30850), .B(n30849), .Z(n30851) );
  NAND U31439 ( .A(n30852), .B(n30851), .Z(n31044) );
  XNOR U31440 ( .A(b[19]), .B(a[203]), .Z(n31011) );
  NANDN U31441 ( .A(n31011), .B(n37934), .Z(n30855) );
  NANDN U31442 ( .A(n30853), .B(n37935), .Z(n30854) );
  NAND U31443 ( .A(n30855), .B(n30854), .Z(n31056) );
  XNOR U31444 ( .A(b[27]), .B(a[195]), .Z(n31014) );
  NANDN U31445 ( .A(n31014), .B(n38423), .Z(n30858) );
  NANDN U31446 ( .A(n30856), .B(n38424), .Z(n30857) );
  NAND U31447 ( .A(n30858), .B(n30857), .Z(n31053) );
  XOR U31448 ( .A(b[5]), .B(n34670), .Z(n31017) );
  NANDN U31449 ( .A(n31017), .B(n36587), .Z(n30861) );
  NANDN U31450 ( .A(n30859), .B(n36588), .Z(n30860) );
  AND U31451 ( .A(n30861), .B(n30860), .Z(n31054) );
  XNOR U31452 ( .A(n31053), .B(n31054), .Z(n31055) );
  XNOR U31453 ( .A(n31056), .B(n31055), .Z(n31041) );
  NANDN U31454 ( .A(n30862), .B(n37762), .Z(n30864) );
  XOR U31455 ( .A(b[17]), .B(a[205]), .Z(n31020) );
  NAND U31456 ( .A(n31020), .B(n37764), .Z(n30863) );
  NAND U31457 ( .A(n30864), .B(n30863), .Z(n30995) );
  XNOR U31458 ( .A(b[31]), .B(a[191]), .Z(n31023) );
  NANDN U31459 ( .A(n31023), .B(n38552), .Z(n30867) );
  NANDN U31460 ( .A(n30865), .B(n38553), .Z(n30866) );
  AND U31461 ( .A(n30867), .B(n30866), .Z(n30993) );
  OR U31462 ( .A(n30868), .B(n36105), .Z(n30870) );
  XNOR U31463 ( .A(b[3]), .B(a[219]), .Z(n31026) );
  NANDN U31464 ( .A(n31026), .B(n36107), .Z(n30869) );
  AND U31465 ( .A(n30870), .B(n30869), .Z(n30994) );
  XOR U31466 ( .A(n30995), .B(n30996), .Z(n31042) );
  XOR U31467 ( .A(n31041), .B(n31042), .Z(n31043) );
  XNOR U31468 ( .A(n31044), .B(n31043), .Z(n31089) );
  NANDN U31469 ( .A(n30872), .B(n30871), .Z(n30876) );
  NAND U31470 ( .A(n30874), .B(n30873), .Z(n30875) );
  NAND U31471 ( .A(n30876), .B(n30875), .Z(n31032) );
  NANDN U31472 ( .A(n30878), .B(n30877), .Z(n30882) );
  NAND U31473 ( .A(n30880), .B(n30879), .Z(n30881) );
  NAND U31474 ( .A(n30882), .B(n30881), .Z(n31030) );
  OR U31475 ( .A(n30884), .B(n30883), .Z(n30888) );
  NANDN U31476 ( .A(n30886), .B(n30885), .Z(n30887) );
  NAND U31477 ( .A(n30888), .B(n30887), .Z(n31029) );
  XNOR U31478 ( .A(n31032), .B(n31031), .Z(n31090) );
  XNOR U31479 ( .A(n31089), .B(n31090), .Z(n31091) );
  NANDN U31480 ( .A(n30890), .B(n30889), .Z(n30894) );
  OR U31481 ( .A(n30892), .B(n30891), .Z(n30893) );
  AND U31482 ( .A(n30894), .B(n30893), .Z(n31092) );
  XOR U31483 ( .A(n31091), .B(n31092), .Z(n31109) );
  NANDN U31484 ( .A(n30900), .B(n30899), .Z(n30904) );
  NANDN U31485 ( .A(n30902), .B(n30901), .Z(n30903) );
  NAND U31486 ( .A(n30904), .B(n30903), .Z(n31098) );
  NANDN U31487 ( .A(n30910), .B(n30909), .Z(n30914) );
  NAND U31488 ( .A(n30912), .B(n30911), .Z(n30913) );
  NAND U31489 ( .A(n30914), .B(n30913), .Z(n31035) );
  NANDN U31490 ( .A(n30916), .B(n30915), .Z(n30920) );
  NAND U31491 ( .A(n30918), .B(n30917), .Z(n30919) );
  AND U31492 ( .A(n30920), .B(n30919), .Z(n31036) );
  XNOR U31493 ( .A(n31035), .B(n31036), .Z(n31037) );
  XNOR U31494 ( .A(n1052), .B(a[213]), .Z(n31065) );
  NAND U31495 ( .A(n36925), .B(n31065), .Z(n30923) );
  NANDN U31496 ( .A(n30921), .B(n36926), .Z(n30922) );
  NAND U31497 ( .A(n30923), .B(n30922), .Z(n31001) );
  XNOR U31498 ( .A(b[15]), .B(a[207]), .Z(n31062) );
  OR U31499 ( .A(n31062), .B(n37665), .Z(n30926) );
  NANDN U31500 ( .A(n30924), .B(n37604), .Z(n30925) );
  AND U31501 ( .A(n30926), .B(n30925), .Z(n30999) );
  XOR U31502 ( .A(n1056), .B(n32687), .Z(n31059) );
  NAND U31503 ( .A(n31059), .B(n38101), .Z(n30929) );
  NANDN U31504 ( .A(n30927), .B(n38102), .Z(n30928) );
  AND U31505 ( .A(n30929), .B(n30928), .Z(n31000) );
  XOR U31506 ( .A(n31001), .B(n31002), .Z(n30990) );
  XNOR U31507 ( .A(b[11]), .B(a[211]), .Z(n31068) );
  OR U31508 ( .A(n31068), .B(n37311), .Z(n30932) );
  NANDN U31509 ( .A(n30930), .B(n37218), .Z(n30931) );
  NAND U31510 ( .A(n30932), .B(n30931), .Z(n30988) );
  XOR U31511 ( .A(n1053), .B(a[209]), .Z(n31071) );
  NANDN U31512 ( .A(n31071), .B(n37424), .Z(n30935) );
  NANDN U31513 ( .A(n30933), .B(n37425), .Z(n30934) );
  NAND U31514 ( .A(n30935), .B(n30934), .Z(n30987) );
  XOR U31515 ( .A(n30990), .B(n30989), .Z(n30984) );
  ANDN U31516 ( .B(b[31]), .A(n30936), .Z(n31005) );
  NANDN U31517 ( .A(n30937), .B(n38490), .Z(n30939) );
  XNOR U31518 ( .A(n1058), .B(a[193]), .Z(n31077) );
  NANDN U31519 ( .A(n1048), .B(n31077), .Z(n30938) );
  NAND U31520 ( .A(n30939), .B(n30938), .Z(n31006) );
  XOR U31521 ( .A(n31005), .B(n31006), .Z(n31007) );
  NANDN U31522 ( .A(n1049), .B(a[221]), .Z(n30940) );
  XNOR U31523 ( .A(b[1]), .B(n30940), .Z(n30942) );
  NANDN U31524 ( .A(b[0]), .B(a[220]), .Z(n30941) );
  AND U31525 ( .A(n30942), .B(n30941), .Z(n31008) );
  XNOR U31526 ( .A(n31007), .B(n31008), .Z(n30981) );
  NANDN U31527 ( .A(n30943), .B(n38205), .Z(n30945) );
  XNOR U31528 ( .A(b[23]), .B(a[199]), .Z(n31080) );
  OR U31529 ( .A(n31080), .B(n38268), .Z(n30944) );
  NAND U31530 ( .A(n30945), .B(n30944), .Z(n31050) );
  XNOR U31531 ( .A(b[7]), .B(a[215]), .Z(n31083) );
  NANDN U31532 ( .A(n31083), .B(n36701), .Z(n30948) );
  NAND U31533 ( .A(n30946), .B(n36702), .Z(n30947) );
  NAND U31534 ( .A(n30948), .B(n30947), .Z(n31047) );
  XOR U31535 ( .A(b[25]), .B(a[197]), .Z(n31086) );
  NAND U31536 ( .A(n31086), .B(n38325), .Z(n30951) );
  NAND U31537 ( .A(n30949), .B(n38326), .Z(n30950) );
  AND U31538 ( .A(n30951), .B(n30950), .Z(n31048) );
  XNOR U31539 ( .A(n31047), .B(n31048), .Z(n31049) );
  XNOR U31540 ( .A(n31050), .B(n31049), .Z(n30982) );
  XOR U31541 ( .A(n30984), .B(n30983), .Z(n31038) );
  XNOR U31542 ( .A(n31037), .B(n31038), .Z(n31095) );
  XOR U31543 ( .A(n31096), .B(n31095), .Z(n31097) );
  XNOR U31544 ( .A(n31098), .B(n31097), .Z(n31107) );
  XNOR U31545 ( .A(n31108), .B(n31107), .Z(n31110) );
  XNOR U31546 ( .A(n31109), .B(n31110), .Z(n31104) );
  XOR U31547 ( .A(n31103), .B(n31104), .Z(n30978) );
  NANDN U31548 ( .A(n30953), .B(n30952), .Z(n30957) );
  NAND U31549 ( .A(n30955), .B(n30954), .Z(n30956) );
  NAND U31550 ( .A(n30957), .B(n30956), .Z(n30975) );
  NANDN U31551 ( .A(n30959), .B(n30958), .Z(n30963) );
  OR U31552 ( .A(n30961), .B(n30960), .Z(n30962) );
  NAND U31553 ( .A(n30963), .B(n30962), .Z(n30976) );
  XNOR U31554 ( .A(n30975), .B(n30976), .Z(n30977) );
  XNOR U31555 ( .A(n30978), .B(n30977), .Z(n30970) );
  XNOR U31556 ( .A(n30969), .B(n30970), .Z(n30971) );
  XNOR U31557 ( .A(n30972), .B(n30971), .Z(n31113) );
  XNOR U31558 ( .A(n31113), .B(sreg[445]), .Z(n31115) );
  NAND U31559 ( .A(n30964), .B(sreg[444]), .Z(n30968) );
  OR U31560 ( .A(n30966), .B(n30965), .Z(n30967) );
  AND U31561 ( .A(n30968), .B(n30967), .Z(n31114) );
  XOR U31562 ( .A(n31115), .B(n31114), .Z(c[445]) );
  NANDN U31563 ( .A(n30970), .B(n30969), .Z(n30974) );
  NAND U31564 ( .A(n30972), .B(n30971), .Z(n30973) );
  NAND U31565 ( .A(n30974), .B(n30973), .Z(n31121) );
  NANDN U31566 ( .A(n30976), .B(n30975), .Z(n30980) );
  NAND U31567 ( .A(n30978), .B(n30977), .Z(n30979) );
  NAND U31568 ( .A(n30980), .B(n30979), .Z(n31119) );
  OR U31569 ( .A(n30982), .B(n30981), .Z(n30986) );
  NANDN U31570 ( .A(n30984), .B(n30983), .Z(n30985) );
  NAND U31571 ( .A(n30986), .B(n30985), .Z(n31249) );
  OR U31572 ( .A(n30988), .B(n30987), .Z(n30992) );
  NAND U31573 ( .A(n30990), .B(n30989), .Z(n30991) );
  NAND U31574 ( .A(n30992), .B(n30991), .Z(n31188) );
  OR U31575 ( .A(n30994), .B(n30993), .Z(n30998) );
  NANDN U31576 ( .A(n30996), .B(n30995), .Z(n30997) );
  NAND U31577 ( .A(n30998), .B(n30997), .Z(n31187) );
  OR U31578 ( .A(n31000), .B(n30999), .Z(n31004) );
  NANDN U31579 ( .A(n31002), .B(n31001), .Z(n31003) );
  NAND U31580 ( .A(n31004), .B(n31003), .Z(n31186) );
  XOR U31581 ( .A(n31188), .B(n31189), .Z(n31247) );
  OR U31582 ( .A(n31006), .B(n31005), .Z(n31010) );
  NANDN U31583 ( .A(n31008), .B(n31007), .Z(n31009) );
  NAND U31584 ( .A(n31010), .B(n31009), .Z(n31200) );
  XOR U31585 ( .A(b[19]), .B(n33130), .Z(n31146) );
  NANDN U31586 ( .A(n31146), .B(n37934), .Z(n31013) );
  NANDN U31587 ( .A(n31011), .B(n37935), .Z(n31012) );
  NAND U31588 ( .A(n31013), .B(n31012), .Z(n31213) );
  XOR U31589 ( .A(b[27]), .B(a[196]), .Z(n31149) );
  NAND U31590 ( .A(n38423), .B(n31149), .Z(n31016) );
  NANDN U31591 ( .A(n31014), .B(n38424), .Z(n31015) );
  NAND U31592 ( .A(n31016), .B(n31015), .Z(n31210) );
  XNOR U31593 ( .A(b[5]), .B(a[218]), .Z(n31152) );
  NANDN U31594 ( .A(n31152), .B(n36587), .Z(n31019) );
  NANDN U31595 ( .A(n31017), .B(n36588), .Z(n31018) );
  AND U31596 ( .A(n31019), .B(n31018), .Z(n31211) );
  XNOR U31597 ( .A(n31210), .B(n31211), .Z(n31212) );
  XNOR U31598 ( .A(n31213), .B(n31212), .Z(n31199) );
  NAND U31599 ( .A(n31020), .B(n37762), .Z(n31022) );
  XOR U31600 ( .A(b[17]), .B(a[206]), .Z(n31155) );
  NAND U31601 ( .A(n31155), .B(n37764), .Z(n31021) );
  NAND U31602 ( .A(n31022), .B(n31021), .Z(n31173) );
  XNOR U31603 ( .A(b[31]), .B(a[192]), .Z(n31158) );
  NANDN U31604 ( .A(n31158), .B(n38552), .Z(n31025) );
  NANDN U31605 ( .A(n31023), .B(n38553), .Z(n31024) );
  NAND U31606 ( .A(n31025), .B(n31024), .Z(n31170) );
  OR U31607 ( .A(n31026), .B(n36105), .Z(n31028) );
  XNOR U31608 ( .A(b[3]), .B(a[220]), .Z(n31161) );
  NANDN U31609 ( .A(n31161), .B(n36107), .Z(n31027) );
  AND U31610 ( .A(n31028), .B(n31027), .Z(n31171) );
  XNOR U31611 ( .A(n31170), .B(n31171), .Z(n31172) );
  XOR U31612 ( .A(n31173), .B(n31172), .Z(n31198) );
  XOR U31613 ( .A(n31199), .B(n31198), .Z(n31201) );
  XOR U31614 ( .A(n31200), .B(n31201), .Z(n31246) );
  XOR U31615 ( .A(n31247), .B(n31246), .Z(n31248) );
  XNOR U31616 ( .A(n31249), .B(n31248), .Z(n31137) );
  OR U31617 ( .A(n31030), .B(n31029), .Z(n31034) );
  NAND U31618 ( .A(n31032), .B(n31031), .Z(n31033) );
  NAND U31619 ( .A(n31034), .B(n31033), .Z(n31135) );
  NANDN U31620 ( .A(n31036), .B(n31035), .Z(n31040) );
  NANDN U31621 ( .A(n31038), .B(n31037), .Z(n31039) );
  NAND U31622 ( .A(n31040), .B(n31039), .Z(n31254) );
  OR U31623 ( .A(n31042), .B(n31041), .Z(n31046) );
  NAND U31624 ( .A(n31044), .B(n31043), .Z(n31045) );
  NAND U31625 ( .A(n31046), .B(n31045), .Z(n31253) );
  NANDN U31626 ( .A(n31048), .B(n31047), .Z(n31052) );
  NAND U31627 ( .A(n31050), .B(n31049), .Z(n31051) );
  NAND U31628 ( .A(n31052), .B(n31051), .Z(n31192) );
  NANDN U31629 ( .A(n31054), .B(n31053), .Z(n31058) );
  NAND U31630 ( .A(n31056), .B(n31055), .Z(n31057) );
  AND U31631 ( .A(n31058), .B(n31057), .Z(n31193) );
  XNOR U31632 ( .A(n31192), .B(n31193), .Z(n31194) );
  XNOR U31633 ( .A(b[21]), .B(a[202]), .Z(n31222) );
  NANDN U31634 ( .A(n31222), .B(n38101), .Z(n31061) );
  NAND U31635 ( .A(n38102), .B(n31059), .Z(n31060) );
  NAND U31636 ( .A(n31061), .B(n31060), .Z(n31182) );
  XNOR U31637 ( .A(b[15]), .B(a[208]), .Z(n31219) );
  OR U31638 ( .A(n31219), .B(n37665), .Z(n31064) );
  NANDN U31639 ( .A(n31062), .B(n37604), .Z(n31063) );
  AND U31640 ( .A(n31064), .B(n31063), .Z(n31183) );
  XNOR U31641 ( .A(n31182), .B(n31183), .Z(n31185) );
  XNOR U31642 ( .A(b[9]), .B(a[214]), .Z(n31216) );
  NANDN U31643 ( .A(n31216), .B(n36925), .Z(n31067) );
  NAND U31644 ( .A(n36926), .B(n31065), .Z(n31066) );
  NAND U31645 ( .A(n31067), .B(n31066), .Z(n31184) );
  XNOR U31646 ( .A(n31185), .B(n31184), .Z(n31178) );
  XNOR U31647 ( .A(b[11]), .B(a[212]), .Z(n31225) );
  OR U31648 ( .A(n31225), .B(n37311), .Z(n31070) );
  NANDN U31649 ( .A(n31068), .B(n37218), .Z(n31069) );
  NAND U31650 ( .A(n31070), .B(n31069), .Z(n31177) );
  XOR U31651 ( .A(n1053), .B(a[210]), .Z(n31228) );
  NANDN U31652 ( .A(n31228), .B(n37424), .Z(n31073) );
  NANDN U31653 ( .A(n31071), .B(n37425), .Z(n31072) );
  NAND U31654 ( .A(n31073), .B(n31072), .Z(n31176) );
  XNOR U31655 ( .A(n31177), .B(n31176), .Z(n31179) );
  XNOR U31656 ( .A(n31178), .B(n31179), .Z(n31167) );
  NANDN U31657 ( .A(n1049), .B(a[222]), .Z(n31074) );
  XNOR U31658 ( .A(b[1]), .B(n31074), .Z(n31076) );
  NANDN U31659 ( .A(b[0]), .B(a[221]), .Z(n31075) );
  AND U31660 ( .A(n31076), .B(n31075), .Z(n31142) );
  NAND U31661 ( .A(n31077), .B(n38490), .Z(n31079) );
  XOR U31662 ( .A(n1058), .B(n31644), .Z(n31231) );
  NANDN U31663 ( .A(n1048), .B(n31231), .Z(n31078) );
  NAND U31664 ( .A(n31079), .B(n31078), .Z(n31140) );
  NANDN U31665 ( .A(n1059), .B(a[190]), .Z(n31141) );
  XNOR U31666 ( .A(n31140), .B(n31141), .Z(n31143) );
  XNOR U31667 ( .A(n31142), .B(n31143), .Z(n31165) );
  NANDN U31668 ( .A(n31080), .B(n38205), .Z(n31082) );
  XNOR U31669 ( .A(b[23]), .B(a[200]), .Z(n31237) );
  OR U31670 ( .A(n31237), .B(n38268), .Z(n31081) );
  NAND U31671 ( .A(n31082), .B(n31081), .Z(n31207) );
  XOR U31672 ( .A(b[7]), .B(a[216]), .Z(n31240) );
  NAND U31673 ( .A(n31240), .B(n36701), .Z(n31085) );
  NANDN U31674 ( .A(n31083), .B(n36702), .Z(n31084) );
  NAND U31675 ( .A(n31085), .B(n31084), .Z(n31204) );
  XNOR U31676 ( .A(b[25]), .B(a[198]), .Z(n31243) );
  NANDN U31677 ( .A(n31243), .B(n38325), .Z(n31088) );
  NAND U31678 ( .A(n31086), .B(n38326), .Z(n31087) );
  AND U31679 ( .A(n31088), .B(n31087), .Z(n31205) );
  XNOR U31680 ( .A(n31204), .B(n31205), .Z(n31206) );
  XOR U31681 ( .A(n31207), .B(n31206), .Z(n31164) );
  XOR U31682 ( .A(n31167), .B(n31166), .Z(n31195) );
  XNOR U31683 ( .A(n31194), .B(n31195), .Z(n31252) );
  XNOR U31684 ( .A(n31253), .B(n31252), .Z(n31255) );
  XNOR U31685 ( .A(n31254), .B(n31255), .Z(n31134) );
  XNOR U31686 ( .A(n31135), .B(n31134), .Z(n31136) );
  XOR U31687 ( .A(n31137), .B(n31136), .Z(n31131) );
  NANDN U31688 ( .A(n31090), .B(n31089), .Z(n31094) );
  NAND U31689 ( .A(n31092), .B(n31091), .Z(n31093) );
  NAND U31690 ( .A(n31094), .B(n31093), .Z(n31128) );
  NAND U31691 ( .A(n31096), .B(n31095), .Z(n31100) );
  NAND U31692 ( .A(n31098), .B(n31097), .Z(n31099) );
  NAND U31693 ( .A(n31100), .B(n31099), .Z(n31129) );
  XNOR U31694 ( .A(n31128), .B(n31129), .Z(n31130) );
  XNOR U31695 ( .A(n31131), .B(n31130), .Z(n31125) );
  NANDN U31696 ( .A(n31102), .B(n31101), .Z(n31106) );
  NANDN U31697 ( .A(n31104), .B(n31103), .Z(n31105) );
  NAND U31698 ( .A(n31106), .B(n31105), .Z(n31123) );
  OR U31699 ( .A(n31108), .B(n31107), .Z(n31112) );
  OR U31700 ( .A(n31110), .B(n31109), .Z(n31111) );
  AND U31701 ( .A(n31112), .B(n31111), .Z(n31122) );
  XNOR U31702 ( .A(n31123), .B(n31122), .Z(n31124) );
  XNOR U31703 ( .A(n31125), .B(n31124), .Z(n31118) );
  XOR U31704 ( .A(n31119), .B(n31118), .Z(n31120) );
  XNOR U31705 ( .A(n31121), .B(n31120), .Z(n31258) );
  XNOR U31706 ( .A(n31258), .B(sreg[446]), .Z(n31260) );
  NAND U31707 ( .A(n31113), .B(sreg[445]), .Z(n31117) );
  OR U31708 ( .A(n31115), .B(n31114), .Z(n31116) );
  AND U31709 ( .A(n31117), .B(n31116), .Z(n31259) );
  XOR U31710 ( .A(n31260), .B(n31259), .Z(c[446]) );
  NANDN U31711 ( .A(n31123), .B(n31122), .Z(n31127) );
  NANDN U31712 ( .A(n31125), .B(n31124), .Z(n31126) );
  NAND U31713 ( .A(n31127), .B(n31126), .Z(n31264) );
  NANDN U31714 ( .A(n31129), .B(n31128), .Z(n31133) );
  NAND U31715 ( .A(n31131), .B(n31130), .Z(n31132) );
  NAND U31716 ( .A(n31133), .B(n31132), .Z(n31269) );
  NANDN U31717 ( .A(n31135), .B(n31134), .Z(n31139) );
  NANDN U31718 ( .A(n31137), .B(n31136), .Z(n31138) );
  NAND U31719 ( .A(n31139), .B(n31138), .Z(n31270) );
  XNOR U31720 ( .A(n31269), .B(n31270), .Z(n31271) );
  NANDN U31721 ( .A(n31141), .B(n31140), .Z(n31145) );
  NAND U31722 ( .A(n31143), .B(n31142), .Z(n31144) );
  NAND U31723 ( .A(n31145), .B(n31144), .Z(n31336) );
  XNOR U31724 ( .A(b[19]), .B(a[205]), .Z(n31281) );
  NANDN U31725 ( .A(n31281), .B(n37934), .Z(n31148) );
  NANDN U31726 ( .A(n31146), .B(n37935), .Z(n31147) );
  NAND U31727 ( .A(n31148), .B(n31147), .Z(n31346) );
  XOR U31728 ( .A(b[27]), .B(a[197]), .Z(n31284) );
  NAND U31729 ( .A(n38423), .B(n31284), .Z(n31151) );
  NAND U31730 ( .A(n31149), .B(n38424), .Z(n31150) );
  NAND U31731 ( .A(n31151), .B(n31150), .Z(n31343) );
  XNOR U31732 ( .A(b[5]), .B(a[219]), .Z(n31287) );
  NANDN U31733 ( .A(n31287), .B(n36587), .Z(n31154) );
  NANDN U31734 ( .A(n31152), .B(n36588), .Z(n31153) );
  AND U31735 ( .A(n31154), .B(n31153), .Z(n31344) );
  XNOR U31736 ( .A(n31343), .B(n31344), .Z(n31345) );
  XNOR U31737 ( .A(n31346), .B(n31345), .Z(n31334) );
  NAND U31738 ( .A(n31155), .B(n37762), .Z(n31157) );
  XOR U31739 ( .A(b[17]), .B(a[207]), .Z(n31290) );
  NAND U31740 ( .A(n31290), .B(n37764), .Z(n31156) );
  NAND U31741 ( .A(n31157), .B(n31156), .Z(n31308) );
  XOR U31742 ( .A(b[31]), .B(n31508), .Z(n31293) );
  NANDN U31743 ( .A(n31293), .B(n38552), .Z(n31160) );
  NANDN U31744 ( .A(n31158), .B(n38553), .Z(n31159) );
  NAND U31745 ( .A(n31160), .B(n31159), .Z(n31305) );
  OR U31746 ( .A(n31161), .B(n36105), .Z(n31163) );
  XNOR U31747 ( .A(b[3]), .B(a[221]), .Z(n31296) );
  NANDN U31748 ( .A(n31296), .B(n36107), .Z(n31162) );
  AND U31749 ( .A(n31163), .B(n31162), .Z(n31306) );
  XNOR U31750 ( .A(n31305), .B(n31306), .Z(n31307) );
  XOR U31751 ( .A(n31308), .B(n31307), .Z(n31333) );
  XNOR U31752 ( .A(n31334), .B(n31333), .Z(n31335) );
  XNOR U31753 ( .A(n31336), .B(n31335), .Z(n31385) );
  NANDN U31754 ( .A(n31165), .B(n31164), .Z(n31169) );
  NANDN U31755 ( .A(n31167), .B(n31166), .Z(n31168) );
  NAND U31756 ( .A(n31169), .B(n31168), .Z(n31386) );
  XNOR U31757 ( .A(n31385), .B(n31386), .Z(n31387) );
  NANDN U31758 ( .A(n31171), .B(n31170), .Z(n31175) );
  NAND U31759 ( .A(n31173), .B(n31172), .Z(n31174) );
  NAND U31760 ( .A(n31175), .B(n31174), .Z(n31326) );
  OR U31761 ( .A(n31177), .B(n31176), .Z(n31181) );
  NANDN U31762 ( .A(n31179), .B(n31178), .Z(n31180) );
  NAND U31763 ( .A(n31181), .B(n31180), .Z(n31324) );
  XNOR U31764 ( .A(n31324), .B(n31323), .Z(n31325) );
  XOR U31765 ( .A(n31326), .B(n31325), .Z(n31388) );
  XOR U31766 ( .A(n31387), .B(n31388), .Z(n31398) );
  OR U31767 ( .A(n31187), .B(n31186), .Z(n31191) );
  NANDN U31768 ( .A(n31189), .B(n31188), .Z(n31190) );
  NAND U31769 ( .A(n31191), .B(n31190), .Z(n31396) );
  NANDN U31770 ( .A(n31193), .B(n31192), .Z(n31197) );
  NANDN U31771 ( .A(n31195), .B(n31194), .Z(n31196) );
  NAND U31772 ( .A(n31197), .B(n31196), .Z(n31381) );
  NANDN U31773 ( .A(n31199), .B(n31198), .Z(n31203) );
  OR U31774 ( .A(n31201), .B(n31200), .Z(n31202) );
  NAND U31775 ( .A(n31203), .B(n31202), .Z(n31380) );
  NANDN U31776 ( .A(n31205), .B(n31204), .Z(n31209) );
  NAND U31777 ( .A(n31207), .B(n31206), .Z(n31208) );
  NAND U31778 ( .A(n31209), .B(n31208), .Z(n31327) );
  NANDN U31779 ( .A(n31211), .B(n31210), .Z(n31215) );
  NAND U31780 ( .A(n31213), .B(n31212), .Z(n31214) );
  AND U31781 ( .A(n31215), .B(n31214), .Z(n31328) );
  XNOR U31782 ( .A(n31327), .B(n31328), .Z(n31329) );
  XOR U31783 ( .A(b[9]), .B(n34725), .Z(n31349) );
  NANDN U31784 ( .A(n31349), .B(n36925), .Z(n31218) );
  NANDN U31785 ( .A(n31216), .B(n36926), .Z(n31217) );
  NAND U31786 ( .A(n31218), .B(n31217), .Z(n31313) );
  XNOR U31787 ( .A(b[15]), .B(a[209]), .Z(n31352) );
  OR U31788 ( .A(n31352), .B(n37665), .Z(n31221) );
  NANDN U31789 ( .A(n31219), .B(n37604), .Z(n31220) );
  AND U31790 ( .A(n31221), .B(n31220), .Z(n31311) );
  XNOR U31791 ( .A(b[21]), .B(a[203]), .Z(n31355) );
  NANDN U31792 ( .A(n31355), .B(n38101), .Z(n31224) );
  NANDN U31793 ( .A(n31222), .B(n38102), .Z(n31223) );
  AND U31794 ( .A(n31224), .B(n31223), .Z(n31312) );
  XOR U31795 ( .A(n31313), .B(n31314), .Z(n31302) );
  XNOR U31796 ( .A(b[11]), .B(a[213]), .Z(n31358) );
  OR U31797 ( .A(n31358), .B(n37311), .Z(n31227) );
  NANDN U31798 ( .A(n31225), .B(n37218), .Z(n31226) );
  NAND U31799 ( .A(n31227), .B(n31226), .Z(n31300) );
  XOR U31800 ( .A(n1053), .B(a[211]), .Z(n31361) );
  NANDN U31801 ( .A(n31361), .B(n37424), .Z(n31230) );
  NANDN U31802 ( .A(n31228), .B(n37425), .Z(n31229) );
  AND U31803 ( .A(n31230), .B(n31229), .Z(n31299) );
  XNOR U31804 ( .A(n31300), .B(n31299), .Z(n31301) );
  XOR U31805 ( .A(n31302), .B(n31301), .Z(n31319) );
  NAND U31806 ( .A(n38490), .B(n31231), .Z(n31233) );
  XOR U31807 ( .A(n1058), .B(n31434), .Z(n31367) );
  NANDN U31808 ( .A(n1048), .B(n31367), .Z(n31232) );
  NAND U31809 ( .A(n31233), .B(n31232), .Z(n31275) );
  NANDN U31810 ( .A(n1059), .B(a[191]), .Z(n31276) );
  XNOR U31811 ( .A(n31275), .B(n31276), .Z(n31278) );
  NANDN U31812 ( .A(n1049), .B(a[223]), .Z(n31234) );
  XNOR U31813 ( .A(b[1]), .B(n31234), .Z(n31236) );
  IV U31814 ( .A(a[222]), .Z(n35381) );
  NANDN U31815 ( .A(n35381), .B(n1049), .Z(n31235) );
  AND U31816 ( .A(n31236), .B(n31235), .Z(n31277) );
  XOR U31817 ( .A(n31278), .B(n31277), .Z(n31317) );
  NANDN U31818 ( .A(n31237), .B(n38205), .Z(n31239) );
  XOR U31819 ( .A(b[23]), .B(n32687), .Z(n31370) );
  OR U31820 ( .A(n31370), .B(n38268), .Z(n31238) );
  NAND U31821 ( .A(n31239), .B(n31238), .Z(n31340) );
  XNOR U31822 ( .A(b[7]), .B(a[217]), .Z(n31373) );
  NANDN U31823 ( .A(n31373), .B(n36701), .Z(n31242) );
  NAND U31824 ( .A(n31240), .B(n36702), .Z(n31241) );
  NAND U31825 ( .A(n31242), .B(n31241), .Z(n31337) );
  XOR U31826 ( .A(b[25]), .B(a[199]), .Z(n31376) );
  NAND U31827 ( .A(n31376), .B(n38325), .Z(n31245) );
  NANDN U31828 ( .A(n31243), .B(n38326), .Z(n31244) );
  AND U31829 ( .A(n31245), .B(n31244), .Z(n31338) );
  XNOR U31830 ( .A(n31337), .B(n31338), .Z(n31339) );
  XNOR U31831 ( .A(n31340), .B(n31339), .Z(n31318) );
  XOR U31832 ( .A(n31317), .B(n31318), .Z(n31320) );
  XNOR U31833 ( .A(n31319), .B(n31320), .Z(n31330) );
  XNOR U31834 ( .A(n31329), .B(n31330), .Z(n31379) );
  XNOR U31835 ( .A(n31380), .B(n31379), .Z(n31382) );
  XNOR U31836 ( .A(n31381), .B(n31382), .Z(n31395) );
  XOR U31837 ( .A(n31396), .B(n31395), .Z(n31397) );
  XNOR U31838 ( .A(n31398), .B(n31397), .Z(n31392) );
  NAND U31839 ( .A(n31247), .B(n31246), .Z(n31251) );
  NAND U31840 ( .A(n31249), .B(n31248), .Z(n31250) );
  NAND U31841 ( .A(n31251), .B(n31250), .Z(n31390) );
  NAND U31842 ( .A(n31253), .B(n31252), .Z(n31257) );
  NANDN U31843 ( .A(n31255), .B(n31254), .Z(n31256) );
  AND U31844 ( .A(n31257), .B(n31256), .Z(n31389) );
  XNOR U31845 ( .A(n31390), .B(n31389), .Z(n31391) );
  XOR U31846 ( .A(n31392), .B(n31391), .Z(n31272) );
  XOR U31847 ( .A(n31271), .B(n31272), .Z(n31263) );
  XOR U31848 ( .A(n31264), .B(n31263), .Z(n31265) );
  XNOR U31849 ( .A(n31266), .B(n31265), .Z(n31401) );
  XNOR U31850 ( .A(n31401), .B(sreg[447]), .Z(n31403) );
  NAND U31851 ( .A(n31258), .B(sreg[446]), .Z(n31262) );
  OR U31852 ( .A(n31260), .B(n31259), .Z(n31261) );
  AND U31853 ( .A(n31262), .B(n31261), .Z(n31402) );
  XOR U31854 ( .A(n31403), .B(n31402), .Z(c[447]) );
  NAND U31855 ( .A(n31264), .B(n31263), .Z(n31268) );
  NAND U31856 ( .A(n31266), .B(n31265), .Z(n31267) );
  NAND U31857 ( .A(n31268), .B(n31267), .Z(n31409) );
  NANDN U31858 ( .A(n31270), .B(n31269), .Z(n31274) );
  NAND U31859 ( .A(n31272), .B(n31271), .Z(n31273) );
  NAND U31860 ( .A(n31274), .B(n31273), .Z(n31407) );
  NANDN U31861 ( .A(n31276), .B(n31275), .Z(n31280) );
  NAND U31862 ( .A(n31278), .B(n31277), .Z(n31279) );
  NAND U31863 ( .A(n31280), .B(n31279), .Z(n31480) );
  XNOR U31864 ( .A(b[19]), .B(a[206]), .Z(n31422) );
  NANDN U31865 ( .A(n31422), .B(n37934), .Z(n31283) );
  NANDN U31866 ( .A(n31281), .B(n37935), .Z(n31282) );
  NAND U31867 ( .A(n31283), .B(n31282), .Z(n31490) );
  XNOR U31868 ( .A(b[27]), .B(a[198]), .Z(n31425) );
  NANDN U31869 ( .A(n31425), .B(n38423), .Z(n31286) );
  NAND U31870 ( .A(n31284), .B(n38424), .Z(n31285) );
  NAND U31871 ( .A(n31286), .B(n31285), .Z(n31487) );
  XNOR U31872 ( .A(b[5]), .B(a[220]), .Z(n31428) );
  NANDN U31873 ( .A(n31428), .B(n36587), .Z(n31289) );
  NANDN U31874 ( .A(n31287), .B(n36588), .Z(n31288) );
  AND U31875 ( .A(n31289), .B(n31288), .Z(n31488) );
  XNOR U31876 ( .A(n31487), .B(n31488), .Z(n31489) );
  XNOR U31877 ( .A(n31490), .B(n31489), .Z(n31478) );
  NAND U31878 ( .A(n31290), .B(n37762), .Z(n31292) );
  XOR U31879 ( .A(b[17]), .B(a[208]), .Z(n31431) );
  NAND U31880 ( .A(n31431), .B(n37764), .Z(n31291) );
  NAND U31881 ( .A(n31292), .B(n31291), .Z(n31450) );
  XOR U31882 ( .A(b[31]), .B(n31644), .Z(n31435) );
  NANDN U31883 ( .A(n31435), .B(n38552), .Z(n31295) );
  NANDN U31884 ( .A(n31293), .B(n38553), .Z(n31294) );
  NAND U31885 ( .A(n31295), .B(n31294), .Z(n31447) );
  OR U31886 ( .A(n31296), .B(n36105), .Z(n31298) );
  XOR U31887 ( .A(b[3]), .B(n35381), .Z(n31438) );
  NANDN U31888 ( .A(n31438), .B(n36107), .Z(n31297) );
  AND U31889 ( .A(n31298), .B(n31297), .Z(n31448) );
  XNOR U31890 ( .A(n31447), .B(n31448), .Z(n31449) );
  XOR U31891 ( .A(n31450), .B(n31449), .Z(n31477) );
  XNOR U31892 ( .A(n31478), .B(n31477), .Z(n31479) );
  XNOR U31893 ( .A(n31480), .B(n31479), .Z(n31524) );
  NANDN U31894 ( .A(n31300), .B(n31299), .Z(n31304) );
  NAND U31895 ( .A(n31302), .B(n31301), .Z(n31303) );
  NAND U31896 ( .A(n31304), .B(n31303), .Z(n31468) );
  NANDN U31897 ( .A(n31306), .B(n31305), .Z(n31310) );
  NAND U31898 ( .A(n31308), .B(n31307), .Z(n31309) );
  NAND U31899 ( .A(n31310), .B(n31309), .Z(n31466) );
  OR U31900 ( .A(n31312), .B(n31311), .Z(n31316) );
  NANDN U31901 ( .A(n31314), .B(n31313), .Z(n31315) );
  NAND U31902 ( .A(n31316), .B(n31315), .Z(n31465) );
  XNOR U31903 ( .A(n31468), .B(n31467), .Z(n31525) );
  XNOR U31904 ( .A(n31524), .B(n31525), .Z(n31526) );
  NANDN U31905 ( .A(n31318), .B(n31317), .Z(n31322) );
  OR U31906 ( .A(n31320), .B(n31319), .Z(n31321) );
  AND U31907 ( .A(n31322), .B(n31321), .Z(n31527) );
  XNOR U31908 ( .A(n31526), .B(n31527), .Z(n31539) );
  NANDN U31909 ( .A(n31328), .B(n31327), .Z(n31332) );
  NANDN U31910 ( .A(n31330), .B(n31329), .Z(n31331) );
  NAND U31911 ( .A(n31332), .B(n31331), .Z(n31533) );
  NANDN U31912 ( .A(n31338), .B(n31337), .Z(n31342) );
  NAND U31913 ( .A(n31340), .B(n31339), .Z(n31341) );
  NAND U31914 ( .A(n31342), .B(n31341), .Z(n31471) );
  NANDN U31915 ( .A(n31344), .B(n31343), .Z(n31348) );
  NAND U31916 ( .A(n31346), .B(n31345), .Z(n31347) );
  AND U31917 ( .A(n31348), .B(n31347), .Z(n31472) );
  XNOR U31918 ( .A(n31471), .B(n31472), .Z(n31473) );
  XNOR U31919 ( .A(b[9]), .B(a[216]), .Z(n31493) );
  NANDN U31920 ( .A(n31493), .B(n36925), .Z(n31351) );
  NANDN U31921 ( .A(n31349), .B(n36926), .Z(n31350) );
  NAND U31922 ( .A(n31351), .B(n31350), .Z(n31455) );
  XNOR U31923 ( .A(b[15]), .B(a[210]), .Z(n31496) );
  OR U31924 ( .A(n31496), .B(n37665), .Z(n31354) );
  NANDN U31925 ( .A(n31352), .B(n37604), .Z(n31353) );
  AND U31926 ( .A(n31354), .B(n31353), .Z(n31453) );
  XOR U31927 ( .A(b[21]), .B(n33130), .Z(n31499) );
  NANDN U31928 ( .A(n31499), .B(n38101), .Z(n31357) );
  NANDN U31929 ( .A(n31355), .B(n38102), .Z(n31356) );
  AND U31930 ( .A(n31357), .B(n31356), .Z(n31454) );
  XOR U31931 ( .A(n31455), .B(n31456), .Z(n31444) );
  XNOR U31932 ( .A(b[11]), .B(a[214]), .Z(n31502) );
  OR U31933 ( .A(n31502), .B(n37311), .Z(n31360) );
  NANDN U31934 ( .A(n31358), .B(n37218), .Z(n31359) );
  NAND U31935 ( .A(n31360), .B(n31359), .Z(n31442) );
  XOR U31936 ( .A(n1053), .B(a[212]), .Z(n31505) );
  NANDN U31937 ( .A(n31505), .B(n37424), .Z(n31363) );
  NANDN U31938 ( .A(n31361), .B(n37425), .Z(n31362) );
  AND U31939 ( .A(n31363), .B(n31362), .Z(n31441) );
  XNOR U31940 ( .A(n31442), .B(n31441), .Z(n31443) );
  XOR U31941 ( .A(n31444), .B(n31443), .Z(n31461) );
  NANDN U31942 ( .A(n1049), .B(a[224]), .Z(n31364) );
  XNOR U31943 ( .A(b[1]), .B(n31364), .Z(n31366) );
  NANDN U31944 ( .A(b[0]), .B(a[223]), .Z(n31365) );
  AND U31945 ( .A(n31366), .B(n31365), .Z(n31418) );
  NAND U31946 ( .A(n38490), .B(n31367), .Z(n31369) );
  XNOR U31947 ( .A(b[29]), .B(a[196]), .Z(n31509) );
  OR U31948 ( .A(n31509), .B(n1048), .Z(n31368) );
  NAND U31949 ( .A(n31369), .B(n31368), .Z(n31416) );
  NANDN U31950 ( .A(n1059), .B(a[192]), .Z(n31417) );
  XNOR U31951 ( .A(n31416), .B(n31417), .Z(n31419) );
  XOR U31952 ( .A(n31418), .B(n31419), .Z(n31459) );
  NANDN U31953 ( .A(n31370), .B(n38205), .Z(n31372) );
  XNOR U31954 ( .A(b[23]), .B(a[202]), .Z(n31515) );
  OR U31955 ( .A(n31515), .B(n38268), .Z(n31371) );
  NAND U31956 ( .A(n31372), .B(n31371), .Z(n31484) );
  XOR U31957 ( .A(b[7]), .B(a[218]), .Z(n31518) );
  NAND U31958 ( .A(n31518), .B(n36701), .Z(n31375) );
  NANDN U31959 ( .A(n31373), .B(n36702), .Z(n31374) );
  NAND U31960 ( .A(n31375), .B(n31374), .Z(n31481) );
  XOR U31961 ( .A(b[25]), .B(a[200]), .Z(n31521) );
  NAND U31962 ( .A(n31521), .B(n38325), .Z(n31378) );
  NAND U31963 ( .A(n31376), .B(n38326), .Z(n31377) );
  AND U31964 ( .A(n31378), .B(n31377), .Z(n31482) );
  XNOR U31965 ( .A(n31481), .B(n31482), .Z(n31483) );
  XNOR U31966 ( .A(n31484), .B(n31483), .Z(n31460) );
  XOR U31967 ( .A(n31459), .B(n31460), .Z(n31462) );
  XNOR U31968 ( .A(n31461), .B(n31462), .Z(n31474) );
  XOR U31969 ( .A(n31473), .B(n31474), .Z(n31531) );
  XNOR U31970 ( .A(n31530), .B(n31531), .Z(n31532) );
  XOR U31971 ( .A(n31533), .B(n31532), .Z(n31537) );
  XNOR U31972 ( .A(n31536), .B(n31537), .Z(n31538) );
  XNOR U31973 ( .A(n31539), .B(n31538), .Z(n31543) );
  NAND U31974 ( .A(n31380), .B(n31379), .Z(n31384) );
  NANDN U31975 ( .A(n31382), .B(n31381), .Z(n31383) );
  NAND U31976 ( .A(n31384), .B(n31383), .Z(n31540) );
  XNOR U31977 ( .A(n31540), .B(n31541), .Z(n31542) );
  XNOR U31978 ( .A(n31543), .B(n31542), .Z(n31413) );
  NANDN U31979 ( .A(n31390), .B(n31389), .Z(n31394) );
  NAND U31980 ( .A(n31392), .B(n31391), .Z(n31393) );
  NAND U31981 ( .A(n31394), .B(n31393), .Z(n31410) );
  NANDN U31982 ( .A(n31396), .B(n31395), .Z(n31400) );
  OR U31983 ( .A(n31398), .B(n31397), .Z(n31399) );
  NAND U31984 ( .A(n31400), .B(n31399), .Z(n31411) );
  XNOR U31985 ( .A(n31410), .B(n31411), .Z(n31412) );
  XNOR U31986 ( .A(n31413), .B(n31412), .Z(n31406) );
  XOR U31987 ( .A(n31407), .B(n31406), .Z(n31408) );
  XNOR U31988 ( .A(n31409), .B(n31408), .Z(n31546) );
  XNOR U31989 ( .A(n31546), .B(sreg[448]), .Z(n31548) );
  NAND U31990 ( .A(n31401), .B(sreg[447]), .Z(n31405) );
  OR U31991 ( .A(n31403), .B(n31402), .Z(n31404) );
  AND U31992 ( .A(n31405), .B(n31404), .Z(n31547) );
  XOR U31993 ( .A(n31548), .B(n31547), .Z(c[448]) );
  NANDN U31994 ( .A(n31411), .B(n31410), .Z(n31415) );
  NANDN U31995 ( .A(n31413), .B(n31412), .Z(n31414) );
  NAND U31996 ( .A(n31415), .B(n31414), .Z(n31552) );
  NANDN U31997 ( .A(n31417), .B(n31416), .Z(n31421) );
  NAND U31998 ( .A(n31419), .B(n31418), .Z(n31420) );
  NAND U31999 ( .A(n31421), .B(n31420), .Z(n31626) );
  XNOR U32000 ( .A(b[19]), .B(a[207]), .Z(n31593) );
  NANDN U32001 ( .A(n31593), .B(n37934), .Z(n31424) );
  NANDN U32002 ( .A(n31422), .B(n37935), .Z(n31423) );
  NAND U32003 ( .A(n31424), .B(n31423), .Z(n31663) );
  XOR U32004 ( .A(b[27]), .B(a[199]), .Z(n31596) );
  NAND U32005 ( .A(n38423), .B(n31596), .Z(n31427) );
  NANDN U32006 ( .A(n31425), .B(n38424), .Z(n31426) );
  NAND U32007 ( .A(n31427), .B(n31426), .Z(n31660) );
  XNOR U32008 ( .A(b[5]), .B(a[221]), .Z(n31599) );
  NANDN U32009 ( .A(n31599), .B(n36587), .Z(n31430) );
  NANDN U32010 ( .A(n31428), .B(n36588), .Z(n31429) );
  AND U32011 ( .A(n31430), .B(n31429), .Z(n31661) );
  XNOR U32012 ( .A(n31660), .B(n31661), .Z(n31662) );
  XNOR U32013 ( .A(n31663), .B(n31662), .Z(n31623) );
  NAND U32014 ( .A(n31431), .B(n37762), .Z(n31433) );
  XOR U32015 ( .A(b[17]), .B(a[209]), .Z(n31602) );
  NAND U32016 ( .A(n31602), .B(n37764), .Z(n31432) );
  NAND U32017 ( .A(n31433), .B(n31432), .Z(n31577) );
  XOR U32018 ( .A(b[31]), .B(n31434), .Z(n31605) );
  NANDN U32019 ( .A(n31605), .B(n38552), .Z(n31437) );
  NANDN U32020 ( .A(n31435), .B(n38553), .Z(n31436) );
  AND U32021 ( .A(n31437), .B(n31436), .Z(n31575) );
  OR U32022 ( .A(n31438), .B(n36105), .Z(n31440) );
  XNOR U32023 ( .A(b[3]), .B(a[223]), .Z(n31608) );
  NANDN U32024 ( .A(n31608), .B(n36107), .Z(n31439) );
  AND U32025 ( .A(n31440), .B(n31439), .Z(n31576) );
  XOR U32026 ( .A(n31577), .B(n31578), .Z(n31624) );
  XOR U32027 ( .A(n31623), .B(n31624), .Z(n31625) );
  XNOR U32028 ( .A(n31626), .B(n31625), .Z(n31672) );
  NANDN U32029 ( .A(n31442), .B(n31441), .Z(n31446) );
  NAND U32030 ( .A(n31444), .B(n31443), .Z(n31445) );
  NAND U32031 ( .A(n31446), .B(n31445), .Z(n31614) );
  NANDN U32032 ( .A(n31448), .B(n31447), .Z(n31452) );
  NAND U32033 ( .A(n31450), .B(n31449), .Z(n31451) );
  NAND U32034 ( .A(n31452), .B(n31451), .Z(n31612) );
  OR U32035 ( .A(n31454), .B(n31453), .Z(n31458) );
  NANDN U32036 ( .A(n31456), .B(n31455), .Z(n31457) );
  NAND U32037 ( .A(n31458), .B(n31457), .Z(n31611) );
  XNOR U32038 ( .A(n31614), .B(n31613), .Z(n31673) );
  XOR U32039 ( .A(n31672), .B(n31673), .Z(n31675) );
  NANDN U32040 ( .A(n31460), .B(n31459), .Z(n31464) );
  OR U32041 ( .A(n31462), .B(n31461), .Z(n31463) );
  NAND U32042 ( .A(n31464), .B(n31463), .Z(n31674) );
  XOR U32043 ( .A(n31675), .B(n31674), .Z(n31692) );
  OR U32044 ( .A(n31466), .B(n31465), .Z(n31470) );
  NAND U32045 ( .A(n31468), .B(n31467), .Z(n31469) );
  NAND U32046 ( .A(n31470), .B(n31469), .Z(n31691) );
  NANDN U32047 ( .A(n31472), .B(n31471), .Z(n31476) );
  NANDN U32048 ( .A(n31474), .B(n31473), .Z(n31475) );
  NAND U32049 ( .A(n31476), .B(n31475), .Z(n31680) );
  NANDN U32050 ( .A(n31482), .B(n31481), .Z(n31486) );
  NAND U32051 ( .A(n31484), .B(n31483), .Z(n31485) );
  NAND U32052 ( .A(n31486), .B(n31485), .Z(n31617) );
  NANDN U32053 ( .A(n31488), .B(n31487), .Z(n31492) );
  NAND U32054 ( .A(n31490), .B(n31489), .Z(n31491) );
  AND U32055 ( .A(n31492), .B(n31491), .Z(n31618) );
  XNOR U32056 ( .A(n31617), .B(n31618), .Z(n31619) );
  XOR U32057 ( .A(b[9]), .B(n34670), .Z(n31629) );
  NANDN U32058 ( .A(n31629), .B(n36925), .Z(n31495) );
  NANDN U32059 ( .A(n31493), .B(n36926), .Z(n31494) );
  NAND U32060 ( .A(n31495), .B(n31494), .Z(n31583) );
  XNOR U32061 ( .A(b[15]), .B(a[211]), .Z(n31632) );
  OR U32062 ( .A(n31632), .B(n37665), .Z(n31498) );
  NANDN U32063 ( .A(n31496), .B(n37604), .Z(n31497) );
  AND U32064 ( .A(n31498), .B(n31497), .Z(n31581) );
  XNOR U32065 ( .A(b[21]), .B(a[205]), .Z(n31635) );
  NANDN U32066 ( .A(n31635), .B(n38101), .Z(n31501) );
  NANDN U32067 ( .A(n31499), .B(n38102), .Z(n31500) );
  AND U32068 ( .A(n31501), .B(n31500), .Z(n31582) );
  XOR U32069 ( .A(n31583), .B(n31584), .Z(n31572) );
  XOR U32070 ( .A(b[11]), .B(n34725), .Z(n31638) );
  OR U32071 ( .A(n31638), .B(n37311), .Z(n31504) );
  NANDN U32072 ( .A(n31502), .B(n37218), .Z(n31503) );
  NAND U32073 ( .A(n31504), .B(n31503), .Z(n31570) );
  XOR U32074 ( .A(n1053), .B(a[213]), .Z(n31641) );
  NANDN U32075 ( .A(n31641), .B(n37424), .Z(n31507) );
  NANDN U32076 ( .A(n31505), .B(n37425), .Z(n31506) );
  NAND U32077 ( .A(n31507), .B(n31506), .Z(n31569) );
  XOR U32078 ( .A(n31572), .B(n31571), .Z(n31566) );
  ANDN U32079 ( .B(b[31]), .A(n31508), .Z(n31587) );
  NANDN U32080 ( .A(n31509), .B(n38490), .Z(n31511) );
  XNOR U32081 ( .A(b[29]), .B(a[197]), .Z(n31645) );
  OR U32082 ( .A(n31645), .B(n1048), .Z(n31510) );
  NAND U32083 ( .A(n31511), .B(n31510), .Z(n31588) );
  XOR U32084 ( .A(n31587), .B(n31588), .Z(n31589) );
  NANDN U32085 ( .A(n1049), .B(a[225]), .Z(n31512) );
  XNOR U32086 ( .A(b[1]), .B(n31512), .Z(n31514) );
  NANDN U32087 ( .A(b[0]), .B(a[224]), .Z(n31513) );
  AND U32088 ( .A(n31514), .B(n31513), .Z(n31590) );
  XNOR U32089 ( .A(n31589), .B(n31590), .Z(n31563) );
  NANDN U32090 ( .A(n31515), .B(n38205), .Z(n31517) );
  XNOR U32091 ( .A(b[23]), .B(a[203]), .Z(n31651) );
  OR U32092 ( .A(n31651), .B(n38268), .Z(n31516) );
  NAND U32093 ( .A(n31517), .B(n31516), .Z(n31669) );
  XOR U32094 ( .A(b[7]), .B(a[219]), .Z(n31654) );
  NAND U32095 ( .A(n31654), .B(n36701), .Z(n31520) );
  NAND U32096 ( .A(n31518), .B(n36702), .Z(n31519) );
  NAND U32097 ( .A(n31520), .B(n31519), .Z(n31666) );
  XNOR U32098 ( .A(b[25]), .B(a[201]), .Z(n31657) );
  NANDN U32099 ( .A(n31657), .B(n38325), .Z(n31523) );
  NAND U32100 ( .A(n31521), .B(n38326), .Z(n31522) );
  AND U32101 ( .A(n31523), .B(n31522), .Z(n31667) );
  XNOR U32102 ( .A(n31666), .B(n31667), .Z(n31668) );
  XNOR U32103 ( .A(n31669), .B(n31668), .Z(n31564) );
  XOR U32104 ( .A(n31566), .B(n31565), .Z(n31620) );
  XNOR U32105 ( .A(n31619), .B(n31620), .Z(n31678) );
  XNOR U32106 ( .A(n31679), .B(n31678), .Z(n31681) );
  XNOR U32107 ( .A(n31680), .B(n31681), .Z(n31690) );
  XOR U32108 ( .A(n31691), .B(n31690), .Z(n31693) );
  NANDN U32109 ( .A(n31525), .B(n31524), .Z(n31529) );
  NAND U32110 ( .A(n31527), .B(n31526), .Z(n31528) );
  NAND U32111 ( .A(n31529), .B(n31528), .Z(n31684) );
  NANDN U32112 ( .A(n31531), .B(n31530), .Z(n31535) );
  NAND U32113 ( .A(n31533), .B(n31532), .Z(n31534) );
  NAND U32114 ( .A(n31535), .B(n31534), .Z(n31685) );
  XNOR U32115 ( .A(n31684), .B(n31685), .Z(n31686) );
  XOR U32116 ( .A(n31687), .B(n31686), .Z(n31559) );
  NANDN U32117 ( .A(n31541), .B(n31540), .Z(n31545) );
  NANDN U32118 ( .A(n31543), .B(n31542), .Z(n31544) );
  NAND U32119 ( .A(n31545), .B(n31544), .Z(n31558) );
  XNOR U32120 ( .A(n31557), .B(n31558), .Z(n31560) );
  XOR U32121 ( .A(n31559), .B(n31560), .Z(n31551) );
  XOR U32122 ( .A(n31552), .B(n31551), .Z(n31553) );
  XNOR U32123 ( .A(n31554), .B(n31553), .Z(n31696) );
  XNOR U32124 ( .A(n31696), .B(sreg[449]), .Z(n31698) );
  NAND U32125 ( .A(n31546), .B(sreg[448]), .Z(n31550) );
  OR U32126 ( .A(n31548), .B(n31547), .Z(n31549) );
  AND U32127 ( .A(n31550), .B(n31549), .Z(n31697) );
  XOR U32128 ( .A(n31698), .B(n31697), .Z(c[449]) );
  NAND U32129 ( .A(n31552), .B(n31551), .Z(n31556) );
  NAND U32130 ( .A(n31554), .B(n31553), .Z(n31555) );
  NAND U32131 ( .A(n31556), .B(n31555), .Z(n31704) );
  NANDN U32132 ( .A(n31558), .B(n31557), .Z(n31562) );
  NAND U32133 ( .A(n31560), .B(n31559), .Z(n31561) );
  NAND U32134 ( .A(n31562), .B(n31561), .Z(n31702) );
  OR U32135 ( .A(n31564), .B(n31563), .Z(n31568) );
  NANDN U32136 ( .A(n31566), .B(n31565), .Z(n31567) );
  NAND U32137 ( .A(n31568), .B(n31567), .Z(n31822) );
  OR U32138 ( .A(n31570), .B(n31569), .Z(n31574) );
  NAND U32139 ( .A(n31572), .B(n31571), .Z(n31573) );
  NAND U32140 ( .A(n31574), .B(n31573), .Z(n31761) );
  OR U32141 ( .A(n31576), .B(n31575), .Z(n31580) );
  NANDN U32142 ( .A(n31578), .B(n31577), .Z(n31579) );
  NAND U32143 ( .A(n31580), .B(n31579), .Z(n31760) );
  OR U32144 ( .A(n31582), .B(n31581), .Z(n31586) );
  NANDN U32145 ( .A(n31584), .B(n31583), .Z(n31585) );
  NAND U32146 ( .A(n31586), .B(n31585), .Z(n31759) );
  XOR U32147 ( .A(n31761), .B(n31762), .Z(n31820) );
  OR U32148 ( .A(n31588), .B(n31587), .Z(n31592) );
  NANDN U32149 ( .A(n31590), .B(n31589), .Z(n31591) );
  NAND U32150 ( .A(n31592), .B(n31591), .Z(n31774) );
  XNOR U32151 ( .A(b[19]), .B(a[208]), .Z(n31741) );
  NANDN U32152 ( .A(n31741), .B(n37934), .Z(n31595) );
  NANDN U32153 ( .A(n31593), .B(n37935), .Z(n31594) );
  NAND U32154 ( .A(n31595), .B(n31594), .Z(n31786) );
  XOR U32155 ( .A(b[27]), .B(a[200]), .Z(n31744) );
  NAND U32156 ( .A(n38423), .B(n31744), .Z(n31598) );
  NAND U32157 ( .A(n31596), .B(n38424), .Z(n31597) );
  NAND U32158 ( .A(n31598), .B(n31597), .Z(n31783) );
  XOR U32159 ( .A(b[5]), .B(n35381), .Z(n31747) );
  NANDN U32160 ( .A(n31747), .B(n36587), .Z(n31601) );
  NANDN U32161 ( .A(n31599), .B(n36588), .Z(n31600) );
  AND U32162 ( .A(n31601), .B(n31600), .Z(n31784) );
  XNOR U32163 ( .A(n31783), .B(n31784), .Z(n31785) );
  XNOR U32164 ( .A(n31786), .B(n31785), .Z(n31771) );
  NAND U32165 ( .A(n31602), .B(n37762), .Z(n31604) );
  XOR U32166 ( .A(b[17]), .B(a[210]), .Z(n31750) );
  NAND U32167 ( .A(n31750), .B(n37764), .Z(n31603) );
  NAND U32168 ( .A(n31604), .B(n31603), .Z(n31725) );
  XNOR U32169 ( .A(b[31]), .B(a[196]), .Z(n31753) );
  NANDN U32170 ( .A(n31753), .B(n38552), .Z(n31607) );
  NANDN U32171 ( .A(n31605), .B(n38553), .Z(n31606) );
  AND U32172 ( .A(n31607), .B(n31606), .Z(n31723) );
  OR U32173 ( .A(n31608), .B(n36105), .Z(n31610) );
  XNOR U32174 ( .A(b[3]), .B(a[224]), .Z(n31756) );
  NANDN U32175 ( .A(n31756), .B(n36107), .Z(n31609) );
  AND U32176 ( .A(n31610), .B(n31609), .Z(n31724) );
  XOR U32177 ( .A(n31725), .B(n31726), .Z(n31772) );
  XOR U32178 ( .A(n31771), .B(n31772), .Z(n31773) );
  XNOR U32179 ( .A(n31774), .B(n31773), .Z(n31819) );
  XOR U32180 ( .A(n31820), .B(n31819), .Z(n31821) );
  XNOR U32181 ( .A(n31822), .B(n31821), .Z(n31838) );
  OR U32182 ( .A(n31612), .B(n31611), .Z(n31616) );
  NAND U32183 ( .A(n31614), .B(n31613), .Z(n31615) );
  NAND U32184 ( .A(n31616), .B(n31615), .Z(n31836) );
  NANDN U32185 ( .A(n31618), .B(n31617), .Z(n31622) );
  NANDN U32186 ( .A(n31620), .B(n31619), .Z(n31621) );
  NAND U32187 ( .A(n31622), .B(n31621), .Z(n31826) );
  OR U32188 ( .A(n31624), .B(n31623), .Z(n31628) );
  NAND U32189 ( .A(n31626), .B(n31625), .Z(n31627) );
  NAND U32190 ( .A(n31628), .B(n31627), .Z(n31823) );
  XNOR U32191 ( .A(n1052), .B(a[218]), .Z(n31789) );
  NAND U32192 ( .A(n36925), .B(n31789), .Z(n31631) );
  NANDN U32193 ( .A(n31629), .B(n36926), .Z(n31630) );
  NAND U32194 ( .A(n31631), .B(n31630), .Z(n31731) );
  XNOR U32195 ( .A(b[15]), .B(a[212]), .Z(n31792) );
  OR U32196 ( .A(n31792), .B(n37665), .Z(n31634) );
  NANDN U32197 ( .A(n31632), .B(n37604), .Z(n31633) );
  AND U32198 ( .A(n31634), .B(n31633), .Z(n31729) );
  XNOR U32199 ( .A(n1056), .B(a[206]), .Z(n31795) );
  NAND U32200 ( .A(n31795), .B(n38101), .Z(n31637) );
  NANDN U32201 ( .A(n31635), .B(n38102), .Z(n31636) );
  AND U32202 ( .A(n31637), .B(n31636), .Z(n31730) );
  XOR U32203 ( .A(n31731), .B(n31732), .Z(n31720) );
  XNOR U32204 ( .A(b[11]), .B(a[216]), .Z(n31798) );
  OR U32205 ( .A(n31798), .B(n37311), .Z(n31640) );
  NANDN U32206 ( .A(n31638), .B(n37218), .Z(n31639) );
  NAND U32207 ( .A(n31640), .B(n31639), .Z(n31718) );
  XOR U32208 ( .A(n1053), .B(a[214]), .Z(n31801) );
  NANDN U32209 ( .A(n31801), .B(n37424), .Z(n31643) );
  NANDN U32210 ( .A(n31641), .B(n37425), .Z(n31642) );
  NAND U32211 ( .A(n31643), .B(n31642), .Z(n31717) );
  XOR U32212 ( .A(n31720), .B(n31719), .Z(n31714) );
  ANDN U32213 ( .B(b[31]), .A(n31644), .Z(n31735) );
  NANDN U32214 ( .A(n31645), .B(n38490), .Z(n31647) );
  XNOR U32215 ( .A(n1058), .B(a[198]), .Z(n31807) );
  NANDN U32216 ( .A(n1048), .B(n31807), .Z(n31646) );
  NAND U32217 ( .A(n31647), .B(n31646), .Z(n31736) );
  XOR U32218 ( .A(n31735), .B(n31736), .Z(n31737) );
  NANDN U32219 ( .A(n1049), .B(a[226]), .Z(n31648) );
  XNOR U32220 ( .A(b[1]), .B(n31648), .Z(n31650) );
  IV U32221 ( .A(a[225]), .Z(n36167) );
  NANDN U32222 ( .A(n36167), .B(n1049), .Z(n31649) );
  AND U32223 ( .A(n31650), .B(n31649), .Z(n31738) );
  XNOR U32224 ( .A(n31737), .B(n31738), .Z(n31711) );
  NANDN U32225 ( .A(n31651), .B(n38205), .Z(n31653) );
  XOR U32226 ( .A(b[23]), .B(n33130), .Z(n31810) );
  OR U32227 ( .A(n31810), .B(n38268), .Z(n31652) );
  NAND U32228 ( .A(n31653), .B(n31652), .Z(n31780) );
  XOR U32229 ( .A(b[7]), .B(a[220]), .Z(n31813) );
  NAND U32230 ( .A(n31813), .B(n36701), .Z(n31656) );
  NAND U32231 ( .A(n31654), .B(n36702), .Z(n31655) );
  NAND U32232 ( .A(n31656), .B(n31655), .Z(n31777) );
  XOR U32233 ( .A(b[25]), .B(a[202]), .Z(n31816) );
  NAND U32234 ( .A(n31816), .B(n38325), .Z(n31659) );
  NANDN U32235 ( .A(n31657), .B(n38326), .Z(n31658) );
  AND U32236 ( .A(n31659), .B(n31658), .Z(n31778) );
  XNOR U32237 ( .A(n31777), .B(n31778), .Z(n31779) );
  XNOR U32238 ( .A(n31780), .B(n31779), .Z(n31712) );
  XNOR U32239 ( .A(n31714), .B(n31713), .Z(n31768) );
  NANDN U32240 ( .A(n31661), .B(n31660), .Z(n31665) );
  NAND U32241 ( .A(n31663), .B(n31662), .Z(n31664) );
  NAND U32242 ( .A(n31665), .B(n31664), .Z(n31766) );
  NANDN U32243 ( .A(n31667), .B(n31666), .Z(n31671) );
  NAND U32244 ( .A(n31669), .B(n31668), .Z(n31670) );
  AND U32245 ( .A(n31671), .B(n31670), .Z(n31765) );
  XNOR U32246 ( .A(n31766), .B(n31765), .Z(n31767) );
  XNOR U32247 ( .A(n31768), .B(n31767), .Z(n31824) );
  XNOR U32248 ( .A(n31823), .B(n31824), .Z(n31825) );
  XOR U32249 ( .A(n31826), .B(n31825), .Z(n31835) );
  XNOR U32250 ( .A(n31836), .B(n31835), .Z(n31837) );
  XOR U32251 ( .A(n31838), .B(n31837), .Z(n31832) );
  NANDN U32252 ( .A(n31673), .B(n31672), .Z(n31677) );
  OR U32253 ( .A(n31675), .B(n31674), .Z(n31676) );
  NAND U32254 ( .A(n31677), .B(n31676), .Z(n31829) );
  NAND U32255 ( .A(n31679), .B(n31678), .Z(n31683) );
  NANDN U32256 ( .A(n31681), .B(n31680), .Z(n31682) );
  NAND U32257 ( .A(n31683), .B(n31682), .Z(n31830) );
  XNOR U32258 ( .A(n31829), .B(n31830), .Z(n31831) );
  XNOR U32259 ( .A(n31832), .B(n31831), .Z(n31708) );
  NANDN U32260 ( .A(n31685), .B(n31684), .Z(n31689) );
  NAND U32261 ( .A(n31687), .B(n31686), .Z(n31688) );
  NAND U32262 ( .A(n31689), .B(n31688), .Z(n31705) );
  NANDN U32263 ( .A(n31691), .B(n31690), .Z(n31695) );
  OR U32264 ( .A(n31693), .B(n31692), .Z(n31694) );
  NAND U32265 ( .A(n31695), .B(n31694), .Z(n31706) );
  XNOR U32266 ( .A(n31705), .B(n31706), .Z(n31707) );
  XNOR U32267 ( .A(n31708), .B(n31707), .Z(n31701) );
  XOR U32268 ( .A(n31702), .B(n31701), .Z(n31703) );
  XNOR U32269 ( .A(n31704), .B(n31703), .Z(n31841) );
  XNOR U32270 ( .A(n31841), .B(sreg[450]), .Z(n31843) );
  NAND U32271 ( .A(n31696), .B(sreg[449]), .Z(n31700) );
  OR U32272 ( .A(n31698), .B(n31697), .Z(n31699) );
  AND U32273 ( .A(n31700), .B(n31699), .Z(n31842) );
  XOR U32274 ( .A(n31843), .B(n31842), .Z(c[450]) );
  NANDN U32275 ( .A(n31706), .B(n31705), .Z(n31710) );
  NANDN U32276 ( .A(n31708), .B(n31707), .Z(n31709) );
  NAND U32277 ( .A(n31710), .B(n31709), .Z(n31847) );
  OR U32278 ( .A(n31712), .B(n31711), .Z(n31716) );
  NANDN U32279 ( .A(n31714), .B(n31713), .Z(n31715) );
  NAND U32280 ( .A(n31716), .B(n31715), .Z(n31977) );
  OR U32281 ( .A(n31718), .B(n31717), .Z(n31722) );
  NAND U32282 ( .A(n31720), .B(n31719), .Z(n31721) );
  NAND U32283 ( .A(n31722), .B(n31721), .Z(n31916) );
  OR U32284 ( .A(n31724), .B(n31723), .Z(n31728) );
  NANDN U32285 ( .A(n31726), .B(n31725), .Z(n31727) );
  NAND U32286 ( .A(n31728), .B(n31727), .Z(n31915) );
  OR U32287 ( .A(n31730), .B(n31729), .Z(n31734) );
  NANDN U32288 ( .A(n31732), .B(n31731), .Z(n31733) );
  NAND U32289 ( .A(n31734), .B(n31733), .Z(n31914) );
  XOR U32290 ( .A(n31916), .B(n31917), .Z(n31975) );
  OR U32291 ( .A(n31736), .B(n31735), .Z(n31740) );
  NANDN U32292 ( .A(n31738), .B(n31737), .Z(n31739) );
  NAND U32293 ( .A(n31740), .B(n31739), .Z(n31928) );
  XNOR U32294 ( .A(b[19]), .B(a[209]), .Z(n31874) );
  NANDN U32295 ( .A(n31874), .B(n37934), .Z(n31743) );
  NANDN U32296 ( .A(n31741), .B(n37935), .Z(n31742) );
  NAND U32297 ( .A(n31743), .B(n31742), .Z(n31941) );
  XNOR U32298 ( .A(b[27]), .B(a[201]), .Z(n31877) );
  NANDN U32299 ( .A(n31877), .B(n38423), .Z(n31746) );
  NAND U32300 ( .A(n31744), .B(n38424), .Z(n31745) );
  NAND U32301 ( .A(n31746), .B(n31745), .Z(n31938) );
  XNOR U32302 ( .A(b[5]), .B(a[223]), .Z(n31880) );
  NANDN U32303 ( .A(n31880), .B(n36587), .Z(n31749) );
  NANDN U32304 ( .A(n31747), .B(n36588), .Z(n31748) );
  AND U32305 ( .A(n31749), .B(n31748), .Z(n31939) );
  XNOR U32306 ( .A(n31938), .B(n31939), .Z(n31940) );
  XNOR U32307 ( .A(n31941), .B(n31940), .Z(n31927) );
  NAND U32308 ( .A(n31750), .B(n37762), .Z(n31752) );
  XOR U32309 ( .A(b[17]), .B(a[211]), .Z(n31883) );
  NAND U32310 ( .A(n31883), .B(n37764), .Z(n31751) );
  NAND U32311 ( .A(n31752), .B(n31751), .Z(n31901) );
  XNOR U32312 ( .A(b[31]), .B(a[197]), .Z(n31886) );
  NANDN U32313 ( .A(n31886), .B(n38552), .Z(n31755) );
  NANDN U32314 ( .A(n31753), .B(n38553), .Z(n31754) );
  NAND U32315 ( .A(n31755), .B(n31754), .Z(n31898) );
  OR U32316 ( .A(n31756), .B(n36105), .Z(n31758) );
  XOR U32317 ( .A(b[3]), .B(n36167), .Z(n31889) );
  NANDN U32318 ( .A(n31889), .B(n36107), .Z(n31757) );
  AND U32319 ( .A(n31758), .B(n31757), .Z(n31899) );
  XNOR U32320 ( .A(n31898), .B(n31899), .Z(n31900) );
  XOR U32321 ( .A(n31901), .B(n31900), .Z(n31926) );
  XOR U32322 ( .A(n31927), .B(n31926), .Z(n31929) );
  XOR U32323 ( .A(n31928), .B(n31929), .Z(n31974) );
  XOR U32324 ( .A(n31975), .B(n31974), .Z(n31976) );
  XNOR U32325 ( .A(n31977), .B(n31976), .Z(n31865) );
  OR U32326 ( .A(n31760), .B(n31759), .Z(n31764) );
  NANDN U32327 ( .A(n31762), .B(n31761), .Z(n31763) );
  NAND U32328 ( .A(n31764), .B(n31763), .Z(n31863) );
  NANDN U32329 ( .A(n31766), .B(n31765), .Z(n31770) );
  NANDN U32330 ( .A(n31768), .B(n31767), .Z(n31769) );
  NAND U32331 ( .A(n31770), .B(n31769), .Z(n31983) );
  OR U32332 ( .A(n31772), .B(n31771), .Z(n31776) );
  NANDN U32333 ( .A(n31774), .B(n31773), .Z(n31775) );
  NAND U32334 ( .A(n31776), .B(n31775), .Z(n31981) );
  NANDN U32335 ( .A(n31778), .B(n31777), .Z(n31782) );
  NAND U32336 ( .A(n31780), .B(n31779), .Z(n31781) );
  NAND U32337 ( .A(n31782), .B(n31781), .Z(n31920) );
  NANDN U32338 ( .A(n31784), .B(n31783), .Z(n31788) );
  NAND U32339 ( .A(n31786), .B(n31785), .Z(n31787) );
  AND U32340 ( .A(n31788), .B(n31787), .Z(n31921) );
  XNOR U32341 ( .A(n31920), .B(n31921), .Z(n31922) );
  XOR U32342 ( .A(n1052), .B(a[219]), .Z(n31944) );
  NANDN U32343 ( .A(n31944), .B(n36925), .Z(n31791) );
  NAND U32344 ( .A(n36926), .B(n31789), .Z(n31790) );
  NAND U32345 ( .A(n31791), .B(n31790), .Z(n31906) );
  XNOR U32346 ( .A(b[15]), .B(a[213]), .Z(n31947) );
  OR U32347 ( .A(n31947), .B(n37665), .Z(n31794) );
  NANDN U32348 ( .A(n31792), .B(n37604), .Z(n31793) );
  NAND U32349 ( .A(n31794), .B(n31793), .Z(n31904) );
  XOR U32350 ( .A(n1056), .B(a[207]), .Z(n31950) );
  NANDN U32351 ( .A(n31950), .B(n38101), .Z(n31797) );
  NAND U32352 ( .A(n38102), .B(n31795), .Z(n31796) );
  NAND U32353 ( .A(n31797), .B(n31796), .Z(n31905) );
  XNOR U32354 ( .A(n31904), .B(n31905), .Z(n31907) );
  XOR U32355 ( .A(n31906), .B(n31907), .Z(n31895) );
  XOR U32356 ( .A(b[11]), .B(n34670), .Z(n31953) );
  OR U32357 ( .A(n31953), .B(n37311), .Z(n31800) );
  NANDN U32358 ( .A(n31798), .B(n37218), .Z(n31799) );
  NAND U32359 ( .A(n31800), .B(n31799), .Z(n31893) );
  XOR U32360 ( .A(n1053), .B(a[215]), .Z(n31956) );
  NANDN U32361 ( .A(n31956), .B(n37424), .Z(n31803) );
  NANDN U32362 ( .A(n31801), .B(n37425), .Z(n31802) );
  AND U32363 ( .A(n31803), .B(n31802), .Z(n31892) );
  XNOR U32364 ( .A(n31893), .B(n31892), .Z(n31894) );
  XNOR U32365 ( .A(n31895), .B(n31894), .Z(n31911) );
  NANDN U32366 ( .A(n1049), .B(a[227]), .Z(n31804) );
  XNOR U32367 ( .A(b[1]), .B(n31804), .Z(n31806) );
  IV U32368 ( .A(a[226]), .Z(n36280) );
  NANDN U32369 ( .A(n36280), .B(n1049), .Z(n31805) );
  AND U32370 ( .A(n31806), .B(n31805), .Z(n31870) );
  NAND U32371 ( .A(n31807), .B(n38490), .Z(n31809) );
  XNOR U32372 ( .A(n1058), .B(a[199]), .Z(n31962) );
  NANDN U32373 ( .A(n1048), .B(n31962), .Z(n31808) );
  NAND U32374 ( .A(n31809), .B(n31808), .Z(n31868) );
  NANDN U32375 ( .A(n1059), .B(a[195]), .Z(n31869) );
  XNOR U32376 ( .A(n31868), .B(n31869), .Z(n31871) );
  XNOR U32377 ( .A(n31870), .B(n31871), .Z(n31909) );
  NANDN U32378 ( .A(n31810), .B(n38205), .Z(n31812) );
  XNOR U32379 ( .A(b[23]), .B(a[205]), .Z(n31965) );
  OR U32380 ( .A(n31965), .B(n38268), .Z(n31811) );
  NAND U32381 ( .A(n31812), .B(n31811), .Z(n31935) );
  XOR U32382 ( .A(b[7]), .B(a[221]), .Z(n31968) );
  NAND U32383 ( .A(n31968), .B(n36701), .Z(n31815) );
  NAND U32384 ( .A(n31813), .B(n36702), .Z(n31814) );
  NAND U32385 ( .A(n31815), .B(n31814), .Z(n31932) );
  XOR U32386 ( .A(b[25]), .B(a[203]), .Z(n31971) );
  NAND U32387 ( .A(n31971), .B(n38325), .Z(n31818) );
  NAND U32388 ( .A(n31816), .B(n38326), .Z(n31817) );
  AND U32389 ( .A(n31818), .B(n31817), .Z(n31933) );
  XNOR U32390 ( .A(n31932), .B(n31933), .Z(n31934) );
  XOR U32391 ( .A(n31935), .B(n31934), .Z(n31908) );
  XOR U32392 ( .A(n31911), .B(n31910), .Z(n31923) );
  XOR U32393 ( .A(n31922), .B(n31923), .Z(n31980) );
  XOR U32394 ( .A(n31981), .B(n31980), .Z(n31982) );
  XNOR U32395 ( .A(n31983), .B(n31982), .Z(n31862) );
  XNOR U32396 ( .A(n31863), .B(n31862), .Z(n31864) );
  XOR U32397 ( .A(n31865), .B(n31864), .Z(n31859) );
  NANDN U32398 ( .A(n31824), .B(n31823), .Z(n31828) );
  NAND U32399 ( .A(n31826), .B(n31825), .Z(n31827) );
  AND U32400 ( .A(n31828), .B(n31827), .Z(n31856) );
  XNOR U32401 ( .A(n31857), .B(n31856), .Z(n31858) );
  XNOR U32402 ( .A(n31859), .B(n31858), .Z(n31853) );
  NANDN U32403 ( .A(n31830), .B(n31829), .Z(n31834) );
  NAND U32404 ( .A(n31832), .B(n31831), .Z(n31833) );
  NAND U32405 ( .A(n31834), .B(n31833), .Z(n31850) );
  NANDN U32406 ( .A(n31836), .B(n31835), .Z(n31840) );
  NANDN U32407 ( .A(n31838), .B(n31837), .Z(n31839) );
  NAND U32408 ( .A(n31840), .B(n31839), .Z(n31851) );
  XNOR U32409 ( .A(n31850), .B(n31851), .Z(n31852) );
  XNOR U32410 ( .A(n31853), .B(n31852), .Z(n31846) );
  XOR U32411 ( .A(n31847), .B(n31846), .Z(n31848) );
  XNOR U32412 ( .A(n31849), .B(n31848), .Z(n31986) );
  XNOR U32413 ( .A(n31986), .B(sreg[451]), .Z(n31988) );
  NAND U32414 ( .A(n31841), .B(sreg[450]), .Z(n31845) );
  OR U32415 ( .A(n31843), .B(n31842), .Z(n31844) );
  AND U32416 ( .A(n31845), .B(n31844), .Z(n31987) );
  XOR U32417 ( .A(n31988), .B(n31987), .Z(c[451]) );
  NANDN U32418 ( .A(n31851), .B(n31850), .Z(n31855) );
  NANDN U32419 ( .A(n31853), .B(n31852), .Z(n31854) );
  NAND U32420 ( .A(n31855), .B(n31854), .Z(n31992) );
  NANDN U32421 ( .A(n31857), .B(n31856), .Z(n31861) );
  NAND U32422 ( .A(n31859), .B(n31858), .Z(n31860) );
  NAND U32423 ( .A(n31861), .B(n31860), .Z(n31997) );
  NANDN U32424 ( .A(n31863), .B(n31862), .Z(n31867) );
  NANDN U32425 ( .A(n31865), .B(n31864), .Z(n31866) );
  NAND U32426 ( .A(n31867), .B(n31866), .Z(n31998) );
  XNOR U32427 ( .A(n31997), .B(n31998), .Z(n31999) );
  NANDN U32428 ( .A(n31869), .B(n31868), .Z(n31873) );
  NAND U32429 ( .A(n31871), .B(n31870), .Z(n31872) );
  NAND U32430 ( .A(n31873), .B(n31872), .Z(n32072) );
  XNOR U32431 ( .A(b[19]), .B(a[210]), .Z(n32019) );
  NANDN U32432 ( .A(n32019), .B(n37934), .Z(n31876) );
  NANDN U32433 ( .A(n31874), .B(n37935), .Z(n31875) );
  NAND U32434 ( .A(n31876), .B(n31875), .Z(n32082) );
  XOR U32435 ( .A(b[27]), .B(a[202]), .Z(n32022) );
  NAND U32436 ( .A(n38423), .B(n32022), .Z(n31879) );
  NANDN U32437 ( .A(n31877), .B(n38424), .Z(n31878) );
  NAND U32438 ( .A(n31879), .B(n31878), .Z(n32079) );
  XNOR U32439 ( .A(b[5]), .B(a[224]), .Z(n32025) );
  NANDN U32440 ( .A(n32025), .B(n36587), .Z(n31882) );
  NANDN U32441 ( .A(n31880), .B(n36588), .Z(n31881) );
  AND U32442 ( .A(n31882), .B(n31881), .Z(n32080) );
  XNOR U32443 ( .A(n32079), .B(n32080), .Z(n32081) );
  XNOR U32444 ( .A(n32082), .B(n32081), .Z(n32070) );
  NAND U32445 ( .A(n31883), .B(n37762), .Z(n31885) );
  XOR U32446 ( .A(b[17]), .B(a[212]), .Z(n32028) );
  NAND U32447 ( .A(n32028), .B(n37764), .Z(n31884) );
  NAND U32448 ( .A(n31885), .B(n31884), .Z(n32046) );
  XOR U32449 ( .A(b[31]), .B(n32246), .Z(n32031) );
  NANDN U32450 ( .A(n32031), .B(n38552), .Z(n31888) );
  NANDN U32451 ( .A(n31886), .B(n38553), .Z(n31887) );
  NAND U32452 ( .A(n31888), .B(n31887), .Z(n32043) );
  OR U32453 ( .A(n31889), .B(n36105), .Z(n31891) );
  XOR U32454 ( .A(b[3]), .B(n36280), .Z(n32034) );
  NANDN U32455 ( .A(n32034), .B(n36107), .Z(n31890) );
  AND U32456 ( .A(n31891), .B(n31890), .Z(n32044) );
  XNOR U32457 ( .A(n32043), .B(n32044), .Z(n32045) );
  XOR U32458 ( .A(n32046), .B(n32045), .Z(n32069) );
  XNOR U32459 ( .A(n32070), .B(n32069), .Z(n32071) );
  XNOR U32460 ( .A(n32072), .B(n32071), .Z(n32010) );
  NANDN U32461 ( .A(n31893), .B(n31892), .Z(n31897) );
  NAND U32462 ( .A(n31895), .B(n31894), .Z(n31896) );
  NAND U32463 ( .A(n31897), .B(n31896), .Z(n32061) );
  NANDN U32464 ( .A(n31899), .B(n31898), .Z(n31903) );
  NAND U32465 ( .A(n31901), .B(n31900), .Z(n31902) );
  NAND U32466 ( .A(n31903), .B(n31902), .Z(n32060) );
  XNOR U32467 ( .A(n32060), .B(n32059), .Z(n32062) );
  XOR U32468 ( .A(n32061), .B(n32062), .Z(n32009) );
  XOR U32469 ( .A(n32010), .B(n32009), .Z(n32011) );
  NANDN U32470 ( .A(n31909), .B(n31908), .Z(n31913) );
  NAND U32471 ( .A(n31911), .B(n31910), .Z(n31912) );
  NAND U32472 ( .A(n31913), .B(n31912), .Z(n32012) );
  XNOR U32473 ( .A(n32011), .B(n32012), .Z(n32123) );
  OR U32474 ( .A(n31915), .B(n31914), .Z(n31919) );
  NANDN U32475 ( .A(n31917), .B(n31916), .Z(n31918) );
  NAND U32476 ( .A(n31919), .B(n31918), .Z(n32122) );
  NANDN U32477 ( .A(n31921), .B(n31920), .Z(n31925) );
  NAND U32478 ( .A(n31923), .B(n31922), .Z(n31924) );
  NAND U32479 ( .A(n31925), .B(n31924), .Z(n32005) );
  NANDN U32480 ( .A(n31927), .B(n31926), .Z(n31931) );
  OR U32481 ( .A(n31929), .B(n31928), .Z(n31930) );
  NAND U32482 ( .A(n31931), .B(n31930), .Z(n32004) );
  NANDN U32483 ( .A(n31933), .B(n31932), .Z(n31937) );
  NAND U32484 ( .A(n31935), .B(n31934), .Z(n31936) );
  NAND U32485 ( .A(n31937), .B(n31936), .Z(n32063) );
  NANDN U32486 ( .A(n31939), .B(n31938), .Z(n31943) );
  NAND U32487 ( .A(n31941), .B(n31940), .Z(n31942) );
  AND U32488 ( .A(n31943), .B(n31942), .Z(n32064) );
  XNOR U32489 ( .A(n32063), .B(n32064), .Z(n32065) );
  XNOR U32490 ( .A(b[9]), .B(a[220]), .Z(n32085) );
  NANDN U32491 ( .A(n32085), .B(n36925), .Z(n31946) );
  NANDN U32492 ( .A(n31944), .B(n36926), .Z(n31945) );
  NAND U32493 ( .A(n31946), .B(n31945), .Z(n32051) );
  XNOR U32494 ( .A(n1054), .B(a[214]), .Z(n32088) );
  NANDN U32495 ( .A(n37665), .B(n32088), .Z(n31949) );
  NANDN U32496 ( .A(n31947), .B(n37604), .Z(n31948) );
  NAND U32497 ( .A(n31949), .B(n31948), .Z(n32049) );
  XNOR U32498 ( .A(b[21]), .B(a[208]), .Z(n32091) );
  NANDN U32499 ( .A(n32091), .B(n38101), .Z(n31952) );
  NANDN U32500 ( .A(n31950), .B(n38102), .Z(n31951) );
  NAND U32501 ( .A(n31952), .B(n31951), .Z(n32050) );
  XNOR U32502 ( .A(n32049), .B(n32050), .Z(n32052) );
  XOR U32503 ( .A(n32051), .B(n32052), .Z(n32040) );
  XNOR U32504 ( .A(b[11]), .B(a[218]), .Z(n32094) );
  OR U32505 ( .A(n32094), .B(n37311), .Z(n31955) );
  NANDN U32506 ( .A(n31953), .B(n37218), .Z(n31954) );
  NAND U32507 ( .A(n31955), .B(n31954), .Z(n32038) );
  XOR U32508 ( .A(n1053), .B(a[216]), .Z(n32097) );
  NANDN U32509 ( .A(n32097), .B(n37424), .Z(n31958) );
  NANDN U32510 ( .A(n31956), .B(n37425), .Z(n31957) );
  AND U32511 ( .A(n31958), .B(n31957), .Z(n32037) );
  XNOR U32512 ( .A(n32038), .B(n32037), .Z(n32039) );
  XNOR U32513 ( .A(n32040), .B(n32039), .Z(n32056) );
  NANDN U32514 ( .A(n1049), .B(a[228]), .Z(n31959) );
  XNOR U32515 ( .A(b[1]), .B(n31959), .Z(n31961) );
  NANDN U32516 ( .A(b[0]), .B(a[227]), .Z(n31960) );
  AND U32517 ( .A(n31961), .B(n31960), .Z(n32015) );
  NAND U32518 ( .A(n38490), .B(n31962), .Z(n31964) );
  XNOR U32519 ( .A(n1058), .B(a[200]), .Z(n32100) );
  NANDN U32520 ( .A(n1048), .B(n32100), .Z(n31963) );
  NAND U32521 ( .A(n31964), .B(n31963), .Z(n32013) );
  NANDN U32522 ( .A(n1059), .B(a[196]), .Z(n32014) );
  XNOR U32523 ( .A(n32013), .B(n32014), .Z(n32016) );
  XNOR U32524 ( .A(n32015), .B(n32016), .Z(n32054) );
  NANDN U32525 ( .A(n31965), .B(n38205), .Z(n31967) );
  XNOR U32526 ( .A(b[23]), .B(a[206]), .Z(n32106) );
  OR U32527 ( .A(n32106), .B(n38268), .Z(n31966) );
  NAND U32528 ( .A(n31967), .B(n31966), .Z(n32076) );
  XNOR U32529 ( .A(b[7]), .B(a[222]), .Z(n32109) );
  NANDN U32530 ( .A(n32109), .B(n36701), .Z(n31970) );
  NAND U32531 ( .A(n31968), .B(n36702), .Z(n31969) );
  NAND U32532 ( .A(n31970), .B(n31969), .Z(n32073) );
  XNOR U32533 ( .A(b[25]), .B(a[204]), .Z(n32112) );
  NANDN U32534 ( .A(n32112), .B(n38325), .Z(n31973) );
  NAND U32535 ( .A(n31971), .B(n38326), .Z(n31972) );
  AND U32536 ( .A(n31973), .B(n31972), .Z(n32074) );
  XNOR U32537 ( .A(n32073), .B(n32074), .Z(n32075) );
  XOR U32538 ( .A(n32076), .B(n32075), .Z(n32053) );
  XOR U32539 ( .A(n32056), .B(n32055), .Z(n32066) );
  XOR U32540 ( .A(n32065), .B(n32066), .Z(n32003) );
  XNOR U32541 ( .A(n32004), .B(n32003), .Z(n32006) );
  XNOR U32542 ( .A(n32005), .B(n32006), .Z(n32121) );
  XOR U32543 ( .A(n32122), .B(n32121), .Z(n32124) );
  NAND U32544 ( .A(n31975), .B(n31974), .Z(n31979) );
  NAND U32545 ( .A(n31977), .B(n31976), .Z(n31978) );
  NAND U32546 ( .A(n31979), .B(n31978), .Z(n32116) );
  NAND U32547 ( .A(n31981), .B(n31980), .Z(n31985) );
  NANDN U32548 ( .A(n31983), .B(n31982), .Z(n31984) );
  AND U32549 ( .A(n31985), .B(n31984), .Z(n32115) );
  XNOR U32550 ( .A(n32116), .B(n32115), .Z(n32117) );
  XOR U32551 ( .A(n32118), .B(n32117), .Z(n32000) );
  XOR U32552 ( .A(n31999), .B(n32000), .Z(n31991) );
  XOR U32553 ( .A(n31992), .B(n31991), .Z(n31993) );
  XNOR U32554 ( .A(n31994), .B(n31993), .Z(n32127) );
  XNOR U32555 ( .A(n32127), .B(sreg[452]), .Z(n32129) );
  NAND U32556 ( .A(n31986), .B(sreg[451]), .Z(n31990) );
  OR U32557 ( .A(n31988), .B(n31987), .Z(n31989) );
  AND U32558 ( .A(n31990), .B(n31989), .Z(n32128) );
  XOR U32559 ( .A(n32129), .B(n32128), .Z(c[452]) );
  NAND U32560 ( .A(n31992), .B(n31991), .Z(n31996) );
  NAND U32561 ( .A(n31994), .B(n31993), .Z(n31995) );
  NAND U32562 ( .A(n31996), .B(n31995), .Z(n32135) );
  NANDN U32563 ( .A(n31998), .B(n31997), .Z(n32002) );
  NAND U32564 ( .A(n32000), .B(n31999), .Z(n32001) );
  NAND U32565 ( .A(n32002), .B(n32001), .Z(n32132) );
  NAND U32566 ( .A(n32004), .B(n32003), .Z(n32008) );
  NANDN U32567 ( .A(n32006), .B(n32005), .Z(n32007) );
  NAND U32568 ( .A(n32008), .B(n32007), .Z(n32259) );
  XNOR U32569 ( .A(n32259), .B(n32260), .Z(n32261) );
  NANDN U32570 ( .A(n32014), .B(n32013), .Z(n32018) );
  NAND U32571 ( .A(n32016), .B(n32015), .Z(n32017) );
  NAND U32572 ( .A(n32018), .B(n32017), .Z(n32215) );
  XNOR U32573 ( .A(b[19]), .B(a[211]), .Z(n32160) );
  NANDN U32574 ( .A(n32160), .B(n37934), .Z(n32021) );
  NANDN U32575 ( .A(n32019), .B(n37935), .Z(n32020) );
  NAND U32576 ( .A(n32021), .B(n32020), .Z(n32225) );
  XOR U32577 ( .A(b[27]), .B(a[203]), .Z(n32163) );
  NAND U32578 ( .A(n38423), .B(n32163), .Z(n32024) );
  NAND U32579 ( .A(n32022), .B(n38424), .Z(n32023) );
  NAND U32580 ( .A(n32024), .B(n32023), .Z(n32222) );
  XOR U32581 ( .A(b[5]), .B(n36167), .Z(n32166) );
  NANDN U32582 ( .A(n32166), .B(n36587), .Z(n32027) );
  NANDN U32583 ( .A(n32025), .B(n36588), .Z(n32026) );
  AND U32584 ( .A(n32027), .B(n32026), .Z(n32223) );
  XNOR U32585 ( .A(n32222), .B(n32223), .Z(n32224) );
  XNOR U32586 ( .A(n32225), .B(n32224), .Z(n32213) );
  NAND U32587 ( .A(n32028), .B(n37762), .Z(n32030) );
  XOR U32588 ( .A(b[17]), .B(a[213]), .Z(n32169) );
  NAND U32589 ( .A(n32169), .B(n37764), .Z(n32029) );
  NAND U32590 ( .A(n32030), .B(n32029), .Z(n32187) );
  XNOR U32591 ( .A(b[31]), .B(a[199]), .Z(n32172) );
  NANDN U32592 ( .A(n32172), .B(n38552), .Z(n32033) );
  NANDN U32593 ( .A(n32031), .B(n38553), .Z(n32032) );
  NAND U32594 ( .A(n32033), .B(n32032), .Z(n32184) );
  OR U32595 ( .A(n32034), .B(n36105), .Z(n32036) );
  XNOR U32596 ( .A(b[3]), .B(a[227]), .Z(n32175) );
  NANDN U32597 ( .A(n32175), .B(n36107), .Z(n32035) );
  AND U32598 ( .A(n32036), .B(n32035), .Z(n32185) );
  XNOR U32599 ( .A(n32184), .B(n32185), .Z(n32186) );
  XOR U32600 ( .A(n32187), .B(n32186), .Z(n32212) );
  XNOR U32601 ( .A(n32213), .B(n32212), .Z(n32214) );
  XNOR U32602 ( .A(n32215), .B(n32214), .Z(n32151) );
  NANDN U32603 ( .A(n32038), .B(n32037), .Z(n32042) );
  NAND U32604 ( .A(n32040), .B(n32039), .Z(n32041) );
  NAND U32605 ( .A(n32042), .B(n32041), .Z(n32204) );
  NANDN U32606 ( .A(n32044), .B(n32043), .Z(n32048) );
  NAND U32607 ( .A(n32046), .B(n32045), .Z(n32047) );
  NAND U32608 ( .A(n32048), .B(n32047), .Z(n32203) );
  XNOR U32609 ( .A(n32203), .B(n32202), .Z(n32205) );
  XOR U32610 ( .A(n32204), .B(n32205), .Z(n32150) );
  XOR U32611 ( .A(n32151), .B(n32150), .Z(n32152) );
  NANDN U32612 ( .A(n32054), .B(n32053), .Z(n32058) );
  NAND U32613 ( .A(n32056), .B(n32055), .Z(n32057) );
  AND U32614 ( .A(n32058), .B(n32057), .Z(n32153) );
  XOR U32615 ( .A(n32152), .B(n32153), .Z(n32267) );
  NANDN U32616 ( .A(n32064), .B(n32063), .Z(n32068) );
  NAND U32617 ( .A(n32066), .B(n32065), .Z(n32067) );
  NAND U32618 ( .A(n32068), .B(n32067), .Z(n32147) );
  NANDN U32619 ( .A(n32074), .B(n32073), .Z(n32078) );
  NAND U32620 ( .A(n32076), .B(n32075), .Z(n32077) );
  NAND U32621 ( .A(n32078), .B(n32077), .Z(n32206) );
  NANDN U32622 ( .A(n32080), .B(n32079), .Z(n32084) );
  NAND U32623 ( .A(n32082), .B(n32081), .Z(n32083) );
  AND U32624 ( .A(n32084), .B(n32083), .Z(n32207) );
  XNOR U32625 ( .A(n32206), .B(n32207), .Z(n32208) );
  XNOR U32626 ( .A(b[9]), .B(a[221]), .Z(n32228) );
  NANDN U32627 ( .A(n32228), .B(n36925), .Z(n32087) );
  NANDN U32628 ( .A(n32085), .B(n36926), .Z(n32086) );
  NAND U32629 ( .A(n32087), .B(n32086), .Z(n32192) );
  XOR U32630 ( .A(b[15]), .B(n34725), .Z(n32231) );
  OR U32631 ( .A(n32231), .B(n37665), .Z(n32090) );
  NAND U32632 ( .A(n32088), .B(n37604), .Z(n32089) );
  AND U32633 ( .A(n32090), .B(n32089), .Z(n32190) );
  XNOR U32634 ( .A(b[21]), .B(a[209]), .Z(n32234) );
  NANDN U32635 ( .A(n32234), .B(n38101), .Z(n32093) );
  NANDN U32636 ( .A(n32091), .B(n38102), .Z(n32092) );
  AND U32637 ( .A(n32093), .B(n32092), .Z(n32191) );
  XOR U32638 ( .A(n32192), .B(n32193), .Z(n32181) );
  XNOR U32639 ( .A(b[11]), .B(a[219]), .Z(n32237) );
  OR U32640 ( .A(n32237), .B(n37311), .Z(n32096) );
  NANDN U32641 ( .A(n32094), .B(n37218), .Z(n32095) );
  NAND U32642 ( .A(n32096), .B(n32095), .Z(n32179) );
  XOR U32643 ( .A(n1053), .B(a[217]), .Z(n32240) );
  NANDN U32644 ( .A(n32240), .B(n37424), .Z(n32099) );
  NANDN U32645 ( .A(n32097), .B(n37425), .Z(n32098) );
  AND U32646 ( .A(n32099), .B(n32098), .Z(n32178) );
  XNOR U32647 ( .A(n32179), .B(n32178), .Z(n32180) );
  XOR U32648 ( .A(n32181), .B(n32180), .Z(n32198) );
  NAND U32649 ( .A(n38490), .B(n32100), .Z(n32102) );
  XOR U32650 ( .A(b[29]), .B(n32687), .Z(n32247) );
  OR U32651 ( .A(n32247), .B(n1048), .Z(n32101) );
  NAND U32652 ( .A(n32102), .B(n32101), .Z(n32154) );
  NANDN U32653 ( .A(n1059), .B(a[197]), .Z(n32155) );
  XNOR U32654 ( .A(n32154), .B(n32155), .Z(n32157) );
  NANDN U32655 ( .A(n1049), .B(a[229]), .Z(n32103) );
  XNOR U32656 ( .A(b[1]), .B(n32103), .Z(n32105) );
  IV U32657 ( .A(a[228]), .Z(n36592) );
  NANDN U32658 ( .A(n36592), .B(n1049), .Z(n32104) );
  AND U32659 ( .A(n32105), .B(n32104), .Z(n32156) );
  XOR U32660 ( .A(n32157), .B(n32156), .Z(n32196) );
  NANDN U32661 ( .A(n32106), .B(n38205), .Z(n32108) );
  XNOR U32662 ( .A(b[23]), .B(a[207]), .Z(n32250) );
  OR U32663 ( .A(n32250), .B(n38268), .Z(n32107) );
  NAND U32664 ( .A(n32108), .B(n32107), .Z(n32219) );
  XOR U32665 ( .A(b[7]), .B(a[223]), .Z(n32253) );
  NAND U32666 ( .A(n32253), .B(n36701), .Z(n32111) );
  NANDN U32667 ( .A(n32109), .B(n36702), .Z(n32110) );
  NAND U32668 ( .A(n32111), .B(n32110), .Z(n32216) );
  XOR U32669 ( .A(b[25]), .B(a[205]), .Z(n32256) );
  NAND U32670 ( .A(n32256), .B(n38325), .Z(n32114) );
  NANDN U32671 ( .A(n32112), .B(n38326), .Z(n32113) );
  AND U32672 ( .A(n32114), .B(n32113), .Z(n32217) );
  XNOR U32673 ( .A(n32216), .B(n32217), .Z(n32218) );
  XNOR U32674 ( .A(n32219), .B(n32218), .Z(n32197) );
  XOR U32675 ( .A(n32196), .B(n32197), .Z(n32199) );
  XNOR U32676 ( .A(n32198), .B(n32199), .Z(n32209) );
  XOR U32677 ( .A(n32208), .B(n32209), .Z(n32145) );
  XNOR U32678 ( .A(n32144), .B(n32145), .Z(n32146) );
  XNOR U32679 ( .A(n32147), .B(n32146), .Z(n32265) );
  XNOR U32680 ( .A(n32266), .B(n32265), .Z(n32268) );
  XNOR U32681 ( .A(n32267), .B(n32268), .Z(n32262) );
  XOR U32682 ( .A(n32261), .B(n32262), .Z(n32141) );
  NANDN U32683 ( .A(n32116), .B(n32115), .Z(n32120) );
  NAND U32684 ( .A(n32118), .B(n32117), .Z(n32119) );
  NAND U32685 ( .A(n32120), .B(n32119), .Z(n32138) );
  NANDN U32686 ( .A(n32122), .B(n32121), .Z(n32126) );
  OR U32687 ( .A(n32124), .B(n32123), .Z(n32125) );
  NAND U32688 ( .A(n32126), .B(n32125), .Z(n32139) );
  XNOR U32689 ( .A(n32138), .B(n32139), .Z(n32140) );
  XNOR U32690 ( .A(n32141), .B(n32140), .Z(n32133) );
  XNOR U32691 ( .A(n32132), .B(n32133), .Z(n32134) );
  XNOR U32692 ( .A(n32135), .B(n32134), .Z(n32271) );
  XNOR U32693 ( .A(n32271), .B(sreg[453]), .Z(n32273) );
  NAND U32694 ( .A(n32127), .B(sreg[452]), .Z(n32131) );
  OR U32695 ( .A(n32129), .B(n32128), .Z(n32130) );
  AND U32696 ( .A(n32131), .B(n32130), .Z(n32272) );
  XOR U32697 ( .A(n32273), .B(n32272), .Z(c[453]) );
  NANDN U32698 ( .A(n32133), .B(n32132), .Z(n32137) );
  NAND U32699 ( .A(n32135), .B(n32134), .Z(n32136) );
  NAND U32700 ( .A(n32137), .B(n32136), .Z(n32279) );
  NANDN U32701 ( .A(n32139), .B(n32138), .Z(n32143) );
  NAND U32702 ( .A(n32141), .B(n32140), .Z(n32142) );
  NAND U32703 ( .A(n32143), .B(n32142), .Z(n32276) );
  NANDN U32704 ( .A(n32145), .B(n32144), .Z(n32149) );
  NAND U32705 ( .A(n32147), .B(n32146), .Z(n32148) );
  NAND U32706 ( .A(n32149), .B(n32148), .Z(n32408) );
  XNOR U32707 ( .A(n32408), .B(n32409), .Z(n32410) );
  NANDN U32708 ( .A(n32155), .B(n32154), .Z(n32159) );
  NAND U32709 ( .A(n32157), .B(n32156), .Z(n32158) );
  NAND U32710 ( .A(n32159), .B(n32158), .Z(n32351) );
  XNOR U32711 ( .A(b[19]), .B(a[212]), .Z(n32318) );
  NANDN U32712 ( .A(n32318), .B(n37934), .Z(n32162) );
  NANDN U32713 ( .A(n32160), .B(n37935), .Z(n32161) );
  NAND U32714 ( .A(n32162), .B(n32161), .Z(n32363) );
  XNOR U32715 ( .A(b[27]), .B(a[204]), .Z(n32321) );
  NANDN U32716 ( .A(n32321), .B(n38423), .Z(n32165) );
  NAND U32717 ( .A(n32163), .B(n38424), .Z(n32164) );
  NAND U32718 ( .A(n32165), .B(n32164), .Z(n32360) );
  XOR U32719 ( .A(b[5]), .B(n36280), .Z(n32324) );
  NANDN U32720 ( .A(n32324), .B(n36587), .Z(n32168) );
  NANDN U32721 ( .A(n32166), .B(n36588), .Z(n32167) );
  AND U32722 ( .A(n32168), .B(n32167), .Z(n32361) );
  XNOR U32723 ( .A(n32360), .B(n32361), .Z(n32362) );
  XNOR U32724 ( .A(n32363), .B(n32362), .Z(n32348) );
  NAND U32725 ( .A(n32169), .B(n37762), .Z(n32171) );
  XOR U32726 ( .A(b[17]), .B(a[214]), .Z(n32327) );
  NAND U32727 ( .A(n32327), .B(n37764), .Z(n32170) );
  NAND U32728 ( .A(n32171), .B(n32170), .Z(n32302) );
  XNOR U32729 ( .A(b[31]), .B(a[200]), .Z(n32330) );
  NANDN U32730 ( .A(n32330), .B(n38552), .Z(n32174) );
  NANDN U32731 ( .A(n32172), .B(n38553), .Z(n32173) );
  AND U32732 ( .A(n32174), .B(n32173), .Z(n32300) );
  OR U32733 ( .A(n32175), .B(n36105), .Z(n32177) );
  XOR U32734 ( .A(b[3]), .B(n36592), .Z(n32333) );
  NANDN U32735 ( .A(n32333), .B(n36107), .Z(n32176) );
  AND U32736 ( .A(n32177), .B(n32176), .Z(n32301) );
  XOR U32737 ( .A(n32302), .B(n32303), .Z(n32349) );
  XOR U32738 ( .A(n32348), .B(n32349), .Z(n32350) );
  XNOR U32739 ( .A(n32351), .B(n32350), .Z(n32396) );
  NANDN U32740 ( .A(n32179), .B(n32178), .Z(n32183) );
  NAND U32741 ( .A(n32181), .B(n32180), .Z(n32182) );
  NAND U32742 ( .A(n32183), .B(n32182), .Z(n32339) );
  NANDN U32743 ( .A(n32185), .B(n32184), .Z(n32189) );
  NAND U32744 ( .A(n32187), .B(n32186), .Z(n32188) );
  NAND U32745 ( .A(n32189), .B(n32188), .Z(n32337) );
  OR U32746 ( .A(n32191), .B(n32190), .Z(n32195) );
  NANDN U32747 ( .A(n32193), .B(n32192), .Z(n32194) );
  NAND U32748 ( .A(n32195), .B(n32194), .Z(n32336) );
  XNOR U32749 ( .A(n32339), .B(n32338), .Z(n32397) );
  XNOR U32750 ( .A(n32396), .B(n32397), .Z(n32398) );
  NANDN U32751 ( .A(n32197), .B(n32196), .Z(n32201) );
  OR U32752 ( .A(n32199), .B(n32198), .Z(n32200) );
  AND U32753 ( .A(n32201), .B(n32200), .Z(n32399) );
  XOR U32754 ( .A(n32398), .B(n32399), .Z(n32416) );
  NANDN U32755 ( .A(n32207), .B(n32206), .Z(n32211) );
  NANDN U32756 ( .A(n32209), .B(n32208), .Z(n32210) );
  NAND U32757 ( .A(n32211), .B(n32210), .Z(n32405) );
  NANDN U32758 ( .A(n32217), .B(n32216), .Z(n32221) );
  NAND U32759 ( .A(n32219), .B(n32218), .Z(n32220) );
  NAND U32760 ( .A(n32221), .B(n32220), .Z(n32342) );
  NANDN U32761 ( .A(n32223), .B(n32222), .Z(n32227) );
  NAND U32762 ( .A(n32225), .B(n32224), .Z(n32226) );
  AND U32763 ( .A(n32227), .B(n32226), .Z(n32343) );
  XNOR U32764 ( .A(n32342), .B(n32343), .Z(n32344) );
  XOR U32765 ( .A(b[9]), .B(n35381), .Z(n32366) );
  NANDN U32766 ( .A(n32366), .B(n36925), .Z(n32230) );
  NANDN U32767 ( .A(n32228), .B(n36926), .Z(n32229) );
  NAND U32768 ( .A(n32230), .B(n32229), .Z(n32308) );
  XNOR U32769 ( .A(b[15]), .B(a[216]), .Z(n32369) );
  OR U32770 ( .A(n32369), .B(n37665), .Z(n32233) );
  NANDN U32771 ( .A(n32231), .B(n37604), .Z(n32232) );
  AND U32772 ( .A(n32233), .B(n32232), .Z(n32306) );
  XNOR U32773 ( .A(b[21]), .B(a[210]), .Z(n32372) );
  NANDN U32774 ( .A(n32372), .B(n38101), .Z(n32236) );
  NANDN U32775 ( .A(n32234), .B(n38102), .Z(n32235) );
  AND U32776 ( .A(n32236), .B(n32235), .Z(n32307) );
  XOR U32777 ( .A(n32308), .B(n32309), .Z(n32297) );
  XNOR U32778 ( .A(b[11]), .B(a[220]), .Z(n32375) );
  OR U32779 ( .A(n32375), .B(n37311), .Z(n32239) );
  NANDN U32780 ( .A(n32237), .B(n37218), .Z(n32238) );
  NAND U32781 ( .A(n32239), .B(n32238), .Z(n32295) );
  XOR U32782 ( .A(n1053), .B(a[218]), .Z(n32378) );
  NANDN U32783 ( .A(n32378), .B(n37424), .Z(n32242) );
  NANDN U32784 ( .A(n32240), .B(n37425), .Z(n32241) );
  NAND U32785 ( .A(n32242), .B(n32241), .Z(n32294) );
  XOR U32786 ( .A(n32297), .B(n32296), .Z(n32291) );
  NANDN U32787 ( .A(n1049), .B(a[230]), .Z(n32243) );
  XNOR U32788 ( .A(b[1]), .B(n32243), .Z(n32245) );
  NANDN U32789 ( .A(b[0]), .B(a[229]), .Z(n32244) );
  AND U32790 ( .A(n32245), .B(n32244), .Z(n32315) );
  ANDN U32791 ( .B(b[31]), .A(n32246), .Z(n32312) );
  NANDN U32792 ( .A(n32247), .B(n38490), .Z(n32249) );
  XNOR U32793 ( .A(n1058), .B(a[202]), .Z(n32384) );
  NANDN U32794 ( .A(n1048), .B(n32384), .Z(n32248) );
  NAND U32795 ( .A(n32249), .B(n32248), .Z(n32313) );
  XOR U32796 ( .A(n32312), .B(n32313), .Z(n32314) );
  XNOR U32797 ( .A(n32315), .B(n32314), .Z(n32288) );
  NANDN U32798 ( .A(n32250), .B(n38205), .Z(n32252) );
  XNOR U32799 ( .A(b[23]), .B(a[208]), .Z(n32387) );
  OR U32800 ( .A(n32387), .B(n38268), .Z(n32251) );
  NAND U32801 ( .A(n32252), .B(n32251), .Z(n32357) );
  XOR U32802 ( .A(b[7]), .B(a[224]), .Z(n32390) );
  NAND U32803 ( .A(n32390), .B(n36701), .Z(n32255) );
  NAND U32804 ( .A(n32253), .B(n36702), .Z(n32254) );
  NAND U32805 ( .A(n32255), .B(n32254), .Z(n32354) );
  XOR U32806 ( .A(b[25]), .B(a[206]), .Z(n32393) );
  NAND U32807 ( .A(n32393), .B(n38325), .Z(n32258) );
  NAND U32808 ( .A(n32256), .B(n38326), .Z(n32257) );
  AND U32809 ( .A(n32258), .B(n32257), .Z(n32355) );
  XNOR U32810 ( .A(n32354), .B(n32355), .Z(n32356) );
  XNOR U32811 ( .A(n32357), .B(n32356), .Z(n32289) );
  XOR U32812 ( .A(n32291), .B(n32290), .Z(n32345) );
  XNOR U32813 ( .A(n32344), .B(n32345), .Z(n32402) );
  XOR U32814 ( .A(n32403), .B(n32402), .Z(n32404) );
  XNOR U32815 ( .A(n32405), .B(n32404), .Z(n32414) );
  XNOR U32816 ( .A(n32415), .B(n32414), .Z(n32417) );
  XNOR U32817 ( .A(n32416), .B(n32417), .Z(n32411) );
  XOR U32818 ( .A(n32410), .B(n32411), .Z(n32285) );
  NANDN U32819 ( .A(n32260), .B(n32259), .Z(n32264) );
  NANDN U32820 ( .A(n32262), .B(n32261), .Z(n32263) );
  NAND U32821 ( .A(n32264), .B(n32263), .Z(n32283) );
  OR U32822 ( .A(n32266), .B(n32265), .Z(n32270) );
  OR U32823 ( .A(n32268), .B(n32267), .Z(n32269) );
  AND U32824 ( .A(n32270), .B(n32269), .Z(n32282) );
  XNOR U32825 ( .A(n32283), .B(n32282), .Z(n32284) );
  XNOR U32826 ( .A(n32285), .B(n32284), .Z(n32277) );
  XNOR U32827 ( .A(n32276), .B(n32277), .Z(n32278) );
  XNOR U32828 ( .A(n32279), .B(n32278), .Z(n32420) );
  XNOR U32829 ( .A(n32420), .B(sreg[454]), .Z(n32422) );
  NAND U32830 ( .A(n32271), .B(sreg[453]), .Z(n32275) );
  OR U32831 ( .A(n32273), .B(n32272), .Z(n32274) );
  AND U32832 ( .A(n32275), .B(n32274), .Z(n32421) );
  XOR U32833 ( .A(n32422), .B(n32421), .Z(c[454]) );
  NANDN U32834 ( .A(n32277), .B(n32276), .Z(n32281) );
  NAND U32835 ( .A(n32279), .B(n32278), .Z(n32280) );
  NAND U32836 ( .A(n32281), .B(n32280), .Z(n32428) );
  NANDN U32837 ( .A(n32283), .B(n32282), .Z(n32287) );
  NAND U32838 ( .A(n32285), .B(n32284), .Z(n32286) );
  NAND U32839 ( .A(n32287), .B(n32286), .Z(n32426) );
  OR U32840 ( .A(n32289), .B(n32288), .Z(n32293) );
  NANDN U32841 ( .A(n32291), .B(n32290), .Z(n32292) );
  NAND U32842 ( .A(n32293), .B(n32292), .Z(n32546) );
  OR U32843 ( .A(n32295), .B(n32294), .Z(n32299) );
  NAND U32844 ( .A(n32297), .B(n32296), .Z(n32298) );
  NAND U32845 ( .A(n32299), .B(n32298), .Z(n32485) );
  OR U32846 ( .A(n32301), .B(n32300), .Z(n32305) );
  NANDN U32847 ( .A(n32303), .B(n32302), .Z(n32304) );
  NAND U32848 ( .A(n32305), .B(n32304), .Z(n32484) );
  OR U32849 ( .A(n32307), .B(n32306), .Z(n32311) );
  NANDN U32850 ( .A(n32309), .B(n32308), .Z(n32310) );
  NAND U32851 ( .A(n32311), .B(n32310), .Z(n32483) );
  XOR U32852 ( .A(n32485), .B(n32486), .Z(n32544) );
  OR U32853 ( .A(n32313), .B(n32312), .Z(n32317) );
  NANDN U32854 ( .A(n32315), .B(n32314), .Z(n32316) );
  NAND U32855 ( .A(n32317), .B(n32316), .Z(n32497) );
  XNOR U32856 ( .A(b[19]), .B(a[213]), .Z(n32441) );
  NANDN U32857 ( .A(n32441), .B(n37934), .Z(n32320) );
  NANDN U32858 ( .A(n32318), .B(n37935), .Z(n32319) );
  NAND U32859 ( .A(n32320), .B(n32319), .Z(n32510) );
  XOR U32860 ( .A(b[27]), .B(a[205]), .Z(n32444) );
  NAND U32861 ( .A(n38423), .B(n32444), .Z(n32323) );
  NANDN U32862 ( .A(n32321), .B(n38424), .Z(n32322) );
  NAND U32863 ( .A(n32323), .B(n32322), .Z(n32507) );
  XNOR U32864 ( .A(b[5]), .B(a[227]), .Z(n32447) );
  NANDN U32865 ( .A(n32447), .B(n36587), .Z(n32326) );
  NANDN U32866 ( .A(n32324), .B(n36588), .Z(n32325) );
  AND U32867 ( .A(n32326), .B(n32325), .Z(n32508) );
  XNOR U32868 ( .A(n32507), .B(n32508), .Z(n32509) );
  XNOR U32869 ( .A(n32510), .B(n32509), .Z(n32496) );
  NAND U32870 ( .A(n32327), .B(n37762), .Z(n32329) );
  XNOR U32871 ( .A(b[17]), .B(a[215]), .Z(n32450) );
  NANDN U32872 ( .A(n32450), .B(n37764), .Z(n32328) );
  NAND U32873 ( .A(n32329), .B(n32328), .Z(n32468) );
  XOR U32874 ( .A(b[31]), .B(n32687), .Z(n32453) );
  NANDN U32875 ( .A(n32453), .B(n38552), .Z(n32332) );
  NANDN U32876 ( .A(n32330), .B(n38553), .Z(n32331) );
  NAND U32877 ( .A(n32332), .B(n32331), .Z(n32465) );
  OR U32878 ( .A(n32333), .B(n36105), .Z(n32335) );
  XNOR U32879 ( .A(b[3]), .B(a[229]), .Z(n32456) );
  NANDN U32880 ( .A(n32456), .B(n36107), .Z(n32334) );
  AND U32881 ( .A(n32335), .B(n32334), .Z(n32466) );
  XNOR U32882 ( .A(n32465), .B(n32466), .Z(n32467) );
  XOR U32883 ( .A(n32468), .B(n32467), .Z(n32495) );
  XOR U32884 ( .A(n32496), .B(n32495), .Z(n32498) );
  XOR U32885 ( .A(n32497), .B(n32498), .Z(n32543) );
  XOR U32886 ( .A(n32544), .B(n32543), .Z(n32545) );
  XNOR U32887 ( .A(n32546), .B(n32545), .Z(n32564) );
  OR U32888 ( .A(n32337), .B(n32336), .Z(n32341) );
  NAND U32889 ( .A(n32339), .B(n32338), .Z(n32340) );
  NAND U32890 ( .A(n32341), .B(n32340), .Z(n32562) );
  NANDN U32891 ( .A(n32343), .B(n32342), .Z(n32347) );
  NANDN U32892 ( .A(n32345), .B(n32344), .Z(n32346) );
  NAND U32893 ( .A(n32347), .B(n32346), .Z(n32551) );
  OR U32894 ( .A(n32349), .B(n32348), .Z(n32353) );
  NAND U32895 ( .A(n32351), .B(n32350), .Z(n32352) );
  NAND U32896 ( .A(n32353), .B(n32352), .Z(n32550) );
  NANDN U32897 ( .A(n32355), .B(n32354), .Z(n32359) );
  NAND U32898 ( .A(n32357), .B(n32356), .Z(n32358) );
  NAND U32899 ( .A(n32359), .B(n32358), .Z(n32489) );
  NANDN U32900 ( .A(n32361), .B(n32360), .Z(n32365) );
  NAND U32901 ( .A(n32363), .B(n32362), .Z(n32364) );
  AND U32902 ( .A(n32365), .B(n32364), .Z(n32490) );
  XNOR U32903 ( .A(n32489), .B(n32490), .Z(n32491) );
  XNOR U32904 ( .A(b[9]), .B(a[223]), .Z(n32513) );
  NANDN U32905 ( .A(n32513), .B(n36925), .Z(n32368) );
  NANDN U32906 ( .A(n32366), .B(n36926), .Z(n32367) );
  NAND U32907 ( .A(n32368), .B(n32367), .Z(n32473) );
  XOR U32908 ( .A(b[15]), .B(n34670), .Z(n32516) );
  OR U32909 ( .A(n32516), .B(n37665), .Z(n32371) );
  NANDN U32910 ( .A(n32369), .B(n37604), .Z(n32370) );
  AND U32911 ( .A(n32371), .B(n32370), .Z(n32471) );
  XNOR U32912 ( .A(b[21]), .B(a[211]), .Z(n32519) );
  NANDN U32913 ( .A(n32519), .B(n38101), .Z(n32374) );
  NANDN U32914 ( .A(n32372), .B(n38102), .Z(n32373) );
  AND U32915 ( .A(n32374), .B(n32373), .Z(n32472) );
  XOR U32916 ( .A(n32473), .B(n32474), .Z(n32462) );
  XNOR U32917 ( .A(b[11]), .B(a[221]), .Z(n32522) );
  OR U32918 ( .A(n32522), .B(n37311), .Z(n32377) );
  NANDN U32919 ( .A(n32375), .B(n37218), .Z(n32376) );
  NAND U32920 ( .A(n32377), .B(n32376), .Z(n32460) );
  XOR U32921 ( .A(n1053), .B(a[219]), .Z(n32525) );
  NANDN U32922 ( .A(n32525), .B(n37424), .Z(n32380) );
  NANDN U32923 ( .A(n32378), .B(n37425), .Z(n32379) );
  AND U32924 ( .A(n32380), .B(n32379), .Z(n32459) );
  XNOR U32925 ( .A(n32460), .B(n32459), .Z(n32461) );
  XOR U32926 ( .A(n32462), .B(n32461), .Z(n32479) );
  NANDN U32927 ( .A(n1049), .B(a[231]), .Z(n32381) );
  XNOR U32928 ( .A(b[1]), .B(n32381), .Z(n32383) );
  IV U32929 ( .A(a[230]), .Z(n36333) );
  NANDN U32930 ( .A(n36333), .B(n1049), .Z(n32382) );
  AND U32931 ( .A(n32383), .B(n32382), .Z(n32437) );
  NAND U32932 ( .A(n32384), .B(n38490), .Z(n32386) );
  XNOR U32933 ( .A(n1058), .B(a[203]), .Z(n32528) );
  NANDN U32934 ( .A(n1048), .B(n32528), .Z(n32385) );
  NAND U32935 ( .A(n32386), .B(n32385), .Z(n32435) );
  NANDN U32936 ( .A(n1059), .B(a[199]), .Z(n32436) );
  XNOR U32937 ( .A(n32435), .B(n32436), .Z(n32438) );
  XOR U32938 ( .A(n32437), .B(n32438), .Z(n32477) );
  NANDN U32939 ( .A(n32387), .B(n38205), .Z(n32389) );
  XNOR U32940 ( .A(b[23]), .B(a[209]), .Z(n32534) );
  OR U32941 ( .A(n32534), .B(n38268), .Z(n32388) );
  NAND U32942 ( .A(n32389), .B(n32388), .Z(n32504) );
  XNOR U32943 ( .A(b[7]), .B(a[225]), .Z(n32537) );
  NANDN U32944 ( .A(n32537), .B(n36701), .Z(n32392) );
  NAND U32945 ( .A(n32390), .B(n36702), .Z(n32391) );
  NAND U32946 ( .A(n32392), .B(n32391), .Z(n32501) );
  XOR U32947 ( .A(b[25]), .B(a[207]), .Z(n32540) );
  NAND U32948 ( .A(n32540), .B(n38325), .Z(n32395) );
  NAND U32949 ( .A(n32393), .B(n38326), .Z(n32394) );
  AND U32950 ( .A(n32395), .B(n32394), .Z(n32502) );
  XNOR U32951 ( .A(n32501), .B(n32502), .Z(n32503) );
  XNOR U32952 ( .A(n32504), .B(n32503), .Z(n32478) );
  XOR U32953 ( .A(n32477), .B(n32478), .Z(n32480) );
  XNOR U32954 ( .A(n32479), .B(n32480), .Z(n32492) );
  XNOR U32955 ( .A(n32491), .B(n32492), .Z(n32549) );
  XNOR U32956 ( .A(n32550), .B(n32549), .Z(n32552) );
  XNOR U32957 ( .A(n32551), .B(n32552), .Z(n32561) );
  XNOR U32958 ( .A(n32562), .B(n32561), .Z(n32563) );
  XOR U32959 ( .A(n32564), .B(n32563), .Z(n32558) );
  NANDN U32960 ( .A(n32397), .B(n32396), .Z(n32401) );
  NAND U32961 ( .A(n32399), .B(n32398), .Z(n32400) );
  NAND U32962 ( .A(n32401), .B(n32400), .Z(n32555) );
  NAND U32963 ( .A(n32403), .B(n32402), .Z(n32407) );
  NAND U32964 ( .A(n32405), .B(n32404), .Z(n32406) );
  NAND U32965 ( .A(n32407), .B(n32406), .Z(n32556) );
  XNOR U32966 ( .A(n32555), .B(n32556), .Z(n32557) );
  XNOR U32967 ( .A(n32558), .B(n32557), .Z(n32432) );
  NANDN U32968 ( .A(n32409), .B(n32408), .Z(n32413) );
  NANDN U32969 ( .A(n32411), .B(n32410), .Z(n32412) );
  NAND U32970 ( .A(n32413), .B(n32412), .Z(n32430) );
  OR U32971 ( .A(n32415), .B(n32414), .Z(n32419) );
  OR U32972 ( .A(n32417), .B(n32416), .Z(n32418) );
  AND U32973 ( .A(n32419), .B(n32418), .Z(n32429) );
  XNOR U32974 ( .A(n32430), .B(n32429), .Z(n32431) );
  XNOR U32975 ( .A(n32432), .B(n32431), .Z(n32425) );
  XOR U32976 ( .A(n32426), .B(n32425), .Z(n32427) );
  XNOR U32977 ( .A(n32428), .B(n32427), .Z(n32567) );
  XNOR U32978 ( .A(n32567), .B(sreg[455]), .Z(n32569) );
  NAND U32979 ( .A(n32420), .B(sreg[454]), .Z(n32424) );
  OR U32980 ( .A(n32422), .B(n32421), .Z(n32423) );
  AND U32981 ( .A(n32424), .B(n32423), .Z(n32568) );
  XOR U32982 ( .A(n32569), .B(n32568), .Z(c[455]) );
  NANDN U32983 ( .A(n32430), .B(n32429), .Z(n32434) );
  NANDN U32984 ( .A(n32432), .B(n32431), .Z(n32433) );
  NAND U32985 ( .A(n32434), .B(n32433), .Z(n32573) );
  NANDN U32986 ( .A(n32436), .B(n32435), .Z(n32440) );
  NAND U32987 ( .A(n32438), .B(n32437), .Z(n32439) );
  NAND U32988 ( .A(n32440), .B(n32439), .Z(n32659) );
  XNOR U32989 ( .A(b[19]), .B(a[214]), .Z(n32602) );
  NANDN U32990 ( .A(n32602), .B(n37934), .Z(n32443) );
  NANDN U32991 ( .A(n32441), .B(n37935), .Z(n32442) );
  NAND U32992 ( .A(n32443), .B(n32442), .Z(n32669) );
  XOR U32993 ( .A(b[27]), .B(a[206]), .Z(n32605) );
  NAND U32994 ( .A(n38423), .B(n32605), .Z(n32446) );
  NAND U32995 ( .A(n32444), .B(n38424), .Z(n32445) );
  NAND U32996 ( .A(n32446), .B(n32445), .Z(n32666) );
  XOR U32997 ( .A(b[5]), .B(n36592), .Z(n32608) );
  NANDN U32998 ( .A(n32608), .B(n36587), .Z(n32449) );
  NANDN U32999 ( .A(n32447), .B(n36588), .Z(n32448) );
  AND U33000 ( .A(n32449), .B(n32448), .Z(n32667) );
  XNOR U33001 ( .A(n32666), .B(n32667), .Z(n32668) );
  XNOR U33002 ( .A(n32669), .B(n32668), .Z(n32657) );
  NANDN U33003 ( .A(n32450), .B(n37762), .Z(n32452) );
  XOR U33004 ( .A(b[17]), .B(a[216]), .Z(n32611) );
  NAND U33005 ( .A(n32611), .B(n37764), .Z(n32451) );
  NAND U33006 ( .A(n32452), .B(n32451), .Z(n32629) );
  XNOR U33007 ( .A(b[31]), .B(a[202]), .Z(n32614) );
  NANDN U33008 ( .A(n32614), .B(n38552), .Z(n32455) );
  NANDN U33009 ( .A(n32453), .B(n38553), .Z(n32454) );
  NAND U33010 ( .A(n32455), .B(n32454), .Z(n32626) );
  OR U33011 ( .A(n32456), .B(n36105), .Z(n32458) );
  XOR U33012 ( .A(a[230]), .B(n1050), .Z(n32617) );
  NANDN U33013 ( .A(n32617), .B(n36107), .Z(n32457) );
  AND U33014 ( .A(n32458), .B(n32457), .Z(n32627) );
  XNOR U33015 ( .A(n32626), .B(n32627), .Z(n32628) );
  XOR U33016 ( .A(n32629), .B(n32628), .Z(n32656) );
  XNOR U33017 ( .A(n32657), .B(n32656), .Z(n32658) );
  XNOR U33018 ( .A(n32659), .B(n32658), .Z(n32703) );
  NANDN U33019 ( .A(n32460), .B(n32459), .Z(n32464) );
  NAND U33020 ( .A(n32462), .B(n32461), .Z(n32463) );
  NAND U33021 ( .A(n32464), .B(n32463), .Z(n32647) );
  NANDN U33022 ( .A(n32466), .B(n32465), .Z(n32470) );
  NAND U33023 ( .A(n32468), .B(n32467), .Z(n32469) );
  NAND U33024 ( .A(n32470), .B(n32469), .Z(n32645) );
  OR U33025 ( .A(n32472), .B(n32471), .Z(n32476) );
  NANDN U33026 ( .A(n32474), .B(n32473), .Z(n32475) );
  NAND U33027 ( .A(n32476), .B(n32475), .Z(n32644) );
  XNOR U33028 ( .A(n32647), .B(n32646), .Z(n32704) );
  XOR U33029 ( .A(n32703), .B(n32704), .Z(n32706) );
  NANDN U33030 ( .A(n32478), .B(n32477), .Z(n32482) );
  OR U33031 ( .A(n32480), .B(n32479), .Z(n32481) );
  NAND U33032 ( .A(n32482), .B(n32481), .Z(n32705) );
  XOR U33033 ( .A(n32706), .B(n32705), .Z(n32592) );
  OR U33034 ( .A(n32484), .B(n32483), .Z(n32488) );
  NANDN U33035 ( .A(n32486), .B(n32485), .Z(n32487) );
  NAND U33036 ( .A(n32488), .B(n32487), .Z(n32591) );
  NANDN U33037 ( .A(n32490), .B(n32489), .Z(n32494) );
  NANDN U33038 ( .A(n32492), .B(n32491), .Z(n32493) );
  NAND U33039 ( .A(n32494), .B(n32493), .Z(n32711) );
  NANDN U33040 ( .A(n32496), .B(n32495), .Z(n32500) );
  OR U33041 ( .A(n32498), .B(n32497), .Z(n32499) );
  NAND U33042 ( .A(n32500), .B(n32499), .Z(n32710) );
  NANDN U33043 ( .A(n32502), .B(n32501), .Z(n32506) );
  NAND U33044 ( .A(n32504), .B(n32503), .Z(n32505) );
  NAND U33045 ( .A(n32506), .B(n32505), .Z(n32650) );
  NANDN U33046 ( .A(n32508), .B(n32507), .Z(n32512) );
  NAND U33047 ( .A(n32510), .B(n32509), .Z(n32511) );
  AND U33048 ( .A(n32512), .B(n32511), .Z(n32651) );
  XNOR U33049 ( .A(n32650), .B(n32651), .Z(n32652) );
  XNOR U33050 ( .A(n1052), .B(a[224]), .Z(n32678) );
  NAND U33051 ( .A(n36925), .B(n32678), .Z(n32515) );
  NANDN U33052 ( .A(n32513), .B(n36926), .Z(n32514) );
  NAND U33053 ( .A(n32515), .B(n32514), .Z(n32634) );
  XNOR U33054 ( .A(b[15]), .B(a[218]), .Z(n32675) );
  OR U33055 ( .A(n32675), .B(n37665), .Z(n32518) );
  NANDN U33056 ( .A(n32516), .B(n37604), .Z(n32517) );
  AND U33057 ( .A(n32518), .B(n32517), .Z(n32632) );
  XNOR U33058 ( .A(n1056), .B(a[212]), .Z(n32672) );
  NAND U33059 ( .A(n32672), .B(n38101), .Z(n32521) );
  NANDN U33060 ( .A(n32519), .B(n38102), .Z(n32520) );
  AND U33061 ( .A(n32521), .B(n32520), .Z(n32633) );
  XOR U33062 ( .A(n32634), .B(n32635), .Z(n32623) );
  XOR U33063 ( .A(b[11]), .B(n35381), .Z(n32681) );
  OR U33064 ( .A(n32681), .B(n37311), .Z(n32524) );
  NANDN U33065 ( .A(n32522), .B(n37218), .Z(n32523) );
  NAND U33066 ( .A(n32524), .B(n32523), .Z(n32621) );
  XOR U33067 ( .A(n1053), .B(a[220]), .Z(n32684) );
  NANDN U33068 ( .A(n32684), .B(n37424), .Z(n32527) );
  NANDN U33069 ( .A(n32525), .B(n37425), .Z(n32526) );
  AND U33070 ( .A(n32527), .B(n32526), .Z(n32620) );
  XNOR U33071 ( .A(n32621), .B(n32620), .Z(n32622) );
  XOR U33072 ( .A(n32623), .B(n32622), .Z(n32640) );
  NAND U33073 ( .A(n38490), .B(n32528), .Z(n32530) );
  XOR U33074 ( .A(b[29]), .B(n33130), .Z(n32688) );
  OR U33075 ( .A(n32688), .B(n1048), .Z(n32529) );
  NAND U33076 ( .A(n32530), .B(n32529), .Z(n32596) );
  NANDN U33077 ( .A(n1059), .B(a[200]), .Z(n32597) );
  XNOR U33078 ( .A(n32596), .B(n32597), .Z(n32599) );
  NANDN U33079 ( .A(n1049), .B(a[232]), .Z(n32531) );
  XNOR U33080 ( .A(b[1]), .B(n32531), .Z(n32533) );
  IV U33081 ( .A(a[231]), .Z(n36934) );
  NANDN U33082 ( .A(n36934), .B(n1049), .Z(n32532) );
  AND U33083 ( .A(n32533), .B(n32532), .Z(n32598) );
  XOR U33084 ( .A(n32599), .B(n32598), .Z(n32638) );
  NANDN U33085 ( .A(n32534), .B(n38205), .Z(n32536) );
  XNOR U33086 ( .A(b[23]), .B(a[210]), .Z(n32694) );
  OR U33087 ( .A(n32694), .B(n38268), .Z(n32535) );
  NAND U33088 ( .A(n32536), .B(n32535), .Z(n32663) );
  XNOR U33089 ( .A(b[7]), .B(a[226]), .Z(n32697) );
  NANDN U33090 ( .A(n32697), .B(n36701), .Z(n32539) );
  NANDN U33091 ( .A(n32537), .B(n36702), .Z(n32538) );
  NAND U33092 ( .A(n32539), .B(n32538), .Z(n32660) );
  XOR U33093 ( .A(b[25]), .B(a[208]), .Z(n32700) );
  NAND U33094 ( .A(n32700), .B(n38325), .Z(n32542) );
  NAND U33095 ( .A(n32540), .B(n38326), .Z(n32541) );
  AND U33096 ( .A(n32542), .B(n32541), .Z(n32661) );
  XNOR U33097 ( .A(n32660), .B(n32661), .Z(n32662) );
  XNOR U33098 ( .A(n32663), .B(n32662), .Z(n32639) );
  XOR U33099 ( .A(n32638), .B(n32639), .Z(n32641) );
  XNOR U33100 ( .A(n32640), .B(n32641), .Z(n32653) );
  XNOR U33101 ( .A(n32652), .B(n32653), .Z(n32709) );
  XNOR U33102 ( .A(n32710), .B(n32709), .Z(n32712) );
  XNOR U33103 ( .A(n32711), .B(n32712), .Z(n32590) );
  XOR U33104 ( .A(n32591), .B(n32590), .Z(n32593) );
  NAND U33105 ( .A(n32544), .B(n32543), .Z(n32548) );
  NAND U33106 ( .A(n32546), .B(n32545), .Z(n32547) );
  NAND U33107 ( .A(n32548), .B(n32547), .Z(n32585) );
  NAND U33108 ( .A(n32550), .B(n32549), .Z(n32554) );
  NANDN U33109 ( .A(n32552), .B(n32551), .Z(n32553) );
  AND U33110 ( .A(n32554), .B(n32553), .Z(n32584) );
  XNOR U33111 ( .A(n32585), .B(n32584), .Z(n32586) );
  XOR U33112 ( .A(n32587), .B(n32586), .Z(n32580) );
  NANDN U33113 ( .A(n32556), .B(n32555), .Z(n32560) );
  NAND U33114 ( .A(n32558), .B(n32557), .Z(n32559) );
  NAND U33115 ( .A(n32560), .B(n32559), .Z(n32578) );
  NANDN U33116 ( .A(n32562), .B(n32561), .Z(n32566) );
  NANDN U33117 ( .A(n32564), .B(n32563), .Z(n32565) );
  NAND U33118 ( .A(n32566), .B(n32565), .Z(n32579) );
  XNOR U33119 ( .A(n32578), .B(n32579), .Z(n32581) );
  XOR U33120 ( .A(n32580), .B(n32581), .Z(n32572) );
  XOR U33121 ( .A(n32573), .B(n32572), .Z(n32574) );
  XNOR U33122 ( .A(n32575), .B(n32574), .Z(n32715) );
  XNOR U33123 ( .A(n32715), .B(sreg[456]), .Z(n32717) );
  NAND U33124 ( .A(n32567), .B(sreg[455]), .Z(n32571) );
  OR U33125 ( .A(n32569), .B(n32568), .Z(n32570) );
  AND U33126 ( .A(n32571), .B(n32570), .Z(n32716) );
  XOR U33127 ( .A(n32717), .B(n32716), .Z(c[456]) );
  NAND U33128 ( .A(n32573), .B(n32572), .Z(n32577) );
  NAND U33129 ( .A(n32575), .B(n32574), .Z(n32576) );
  NAND U33130 ( .A(n32577), .B(n32576), .Z(n32723) );
  NANDN U33131 ( .A(n32579), .B(n32578), .Z(n32583) );
  NAND U33132 ( .A(n32581), .B(n32580), .Z(n32582) );
  NAND U33133 ( .A(n32583), .B(n32582), .Z(n32721) );
  NANDN U33134 ( .A(n32585), .B(n32584), .Z(n32589) );
  NAND U33135 ( .A(n32587), .B(n32586), .Z(n32588) );
  NAND U33136 ( .A(n32589), .B(n32588), .Z(n32726) );
  NANDN U33137 ( .A(n32591), .B(n32590), .Z(n32595) );
  OR U33138 ( .A(n32593), .B(n32592), .Z(n32594) );
  NAND U33139 ( .A(n32595), .B(n32594), .Z(n32727) );
  XNOR U33140 ( .A(n32726), .B(n32727), .Z(n32728) );
  NANDN U33141 ( .A(n32597), .B(n32596), .Z(n32601) );
  NAND U33142 ( .A(n32599), .B(n32598), .Z(n32600) );
  NAND U33143 ( .A(n32601), .B(n32600), .Z(n32793) );
  XOR U33144 ( .A(b[19]), .B(n34725), .Z(n32738) );
  NANDN U33145 ( .A(n32738), .B(n37934), .Z(n32604) );
  NANDN U33146 ( .A(n32602), .B(n37935), .Z(n32603) );
  NAND U33147 ( .A(n32604), .B(n32603), .Z(n32803) );
  XOR U33148 ( .A(b[27]), .B(a[207]), .Z(n32741) );
  NAND U33149 ( .A(n38423), .B(n32741), .Z(n32607) );
  NAND U33150 ( .A(n32605), .B(n38424), .Z(n32606) );
  NAND U33151 ( .A(n32607), .B(n32606), .Z(n32800) );
  XNOR U33152 ( .A(b[5]), .B(a[229]), .Z(n32744) );
  NANDN U33153 ( .A(n32744), .B(n36587), .Z(n32610) );
  NANDN U33154 ( .A(n32608), .B(n36588), .Z(n32609) );
  AND U33155 ( .A(n32610), .B(n32609), .Z(n32801) );
  XNOR U33156 ( .A(n32800), .B(n32801), .Z(n32802) );
  XNOR U33157 ( .A(n32803), .B(n32802), .Z(n32791) );
  NAND U33158 ( .A(n32611), .B(n37762), .Z(n32613) );
  XNOR U33159 ( .A(b[17]), .B(a[217]), .Z(n32747) );
  NANDN U33160 ( .A(n32747), .B(n37764), .Z(n32612) );
  NAND U33161 ( .A(n32613), .B(n32612), .Z(n32765) );
  XNOR U33162 ( .A(b[31]), .B(a[203]), .Z(n32750) );
  NANDN U33163 ( .A(n32750), .B(n38552), .Z(n32616) );
  NANDN U33164 ( .A(n32614), .B(n38553), .Z(n32615) );
  NAND U33165 ( .A(n32616), .B(n32615), .Z(n32762) );
  OR U33166 ( .A(n32617), .B(n36105), .Z(n32619) );
  XOR U33167 ( .A(a[231]), .B(n1050), .Z(n32753) );
  NANDN U33168 ( .A(n32753), .B(n36107), .Z(n32618) );
  AND U33169 ( .A(n32619), .B(n32618), .Z(n32763) );
  XNOR U33170 ( .A(n32762), .B(n32763), .Z(n32764) );
  XOR U33171 ( .A(n32765), .B(n32764), .Z(n32790) );
  XNOR U33172 ( .A(n32791), .B(n32790), .Z(n32792) );
  XNOR U33173 ( .A(n32793), .B(n32792), .Z(n32836) );
  NANDN U33174 ( .A(n32621), .B(n32620), .Z(n32625) );
  NAND U33175 ( .A(n32623), .B(n32622), .Z(n32624) );
  NAND U33176 ( .A(n32625), .B(n32624), .Z(n32781) );
  NANDN U33177 ( .A(n32627), .B(n32626), .Z(n32631) );
  NAND U33178 ( .A(n32629), .B(n32628), .Z(n32630) );
  NAND U33179 ( .A(n32631), .B(n32630), .Z(n32779) );
  OR U33180 ( .A(n32633), .B(n32632), .Z(n32637) );
  NANDN U33181 ( .A(n32635), .B(n32634), .Z(n32636) );
  NAND U33182 ( .A(n32637), .B(n32636), .Z(n32778) );
  XNOR U33183 ( .A(n32781), .B(n32780), .Z(n32837) );
  XOR U33184 ( .A(n32836), .B(n32837), .Z(n32839) );
  NANDN U33185 ( .A(n32639), .B(n32638), .Z(n32643) );
  OR U33186 ( .A(n32641), .B(n32640), .Z(n32642) );
  NAND U33187 ( .A(n32643), .B(n32642), .Z(n32838) );
  XOR U33188 ( .A(n32839), .B(n32838), .Z(n32856) );
  OR U33189 ( .A(n32645), .B(n32644), .Z(n32649) );
  NAND U33190 ( .A(n32647), .B(n32646), .Z(n32648) );
  NAND U33191 ( .A(n32649), .B(n32648), .Z(n32855) );
  NANDN U33192 ( .A(n32651), .B(n32650), .Z(n32655) );
  NANDN U33193 ( .A(n32653), .B(n32652), .Z(n32654) );
  NAND U33194 ( .A(n32655), .B(n32654), .Z(n32844) );
  NANDN U33195 ( .A(n32661), .B(n32660), .Z(n32665) );
  NAND U33196 ( .A(n32663), .B(n32662), .Z(n32664) );
  NAND U33197 ( .A(n32665), .B(n32664), .Z(n32784) );
  NANDN U33198 ( .A(n32667), .B(n32666), .Z(n32671) );
  NAND U33199 ( .A(n32669), .B(n32668), .Z(n32670) );
  AND U33200 ( .A(n32671), .B(n32670), .Z(n32785) );
  XNOR U33201 ( .A(n32784), .B(n32785), .Z(n32786) );
  XNOR U33202 ( .A(b[21]), .B(a[213]), .Z(n32812) );
  NANDN U33203 ( .A(n32812), .B(n38101), .Z(n32674) );
  NAND U33204 ( .A(n38102), .B(n32672), .Z(n32673) );
  NAND U33205 ( .A(n32674), .B(n32673), .Z(n32774) );
  XNOR U33206 ( .A(b[15]), .B(a[219]), .Z(n32809) );
  OR U33207 ( .A(n32809), .B(n37665), .Z(n32677) );
  NANDN U33208 ( .A(n32675), .B(n37604), .Z(n32676) );
  AND U33209 ( .A(n32677), .B(n32676), .Z(n32775) );
  XNOR U33210 ( .A(n32774), .B(n32775), .Z(n32777) );
  XOR U33211 ( .A(b[9]), .B(n36167), .Z(n32806) );
  NANDN U33212 ( .A(n32806), .B(n36925), .Z(n32680) );
  NAND U33213 ( .A(n36926), .B(n32678), .Z(n32679) );
  NAND U33214 ( .A(n32680), .B(n32679), .Z(n32776) );
  XNOR U33215 ( .A(n32777), .B(n32776), .Z(n32770) );
  XNOR U33216 ( .A(b[11]), .B(a[223]), .Z(n32815) );
  OR U33217 ( .A(n32815), .B(n37311), .Z(n32683) );
  NANDN U33218 ( .A(n32681), .B(n37218), .Z(n32682) );
  NAND U33219 ( .A(n32683), .B(n32682), .Z(n32769) );
  XOR U33220 ( .A(n1053), .B(a[221]), .Z(n32818) );
  NANDN U33221 ( .A(n32818), .B(n37424), .Z(n32686) );
  NANDN U33222 ( .A(n32684), .B(n37425), .Z(n32685) );
  NAND U33223 ( .A(n32686), .B(n32685), .Z(n32768) );
  XNOR U33224 ( .A(n32769), .B(n32768), .Z(n32771) );
  XNOR U33225 ( .A(n32770), .B(n32771), .Z(n32759) );
  ANDN U33226 ( .B(b[31]), .A(n32687), .Z(n32732) );
  NANDN U33227 ( .A(n32688), .B(n38490), .Z(n32690) );
  XNOR U33228 ( .A(n1058), .B(a[205]), .Z(n32824) );
  NANDN U33229 ( .A(n1048), .B(n32824), .Z(n32689) );
  NAND U33230 ( .A(n32690), .B(n32689), .Z(n32733) );
  XOR U33231 ( .A(n32732), .B(n32733), .Z(n32734) );
  NANDN U33232 ( .A(n1049), .B(a[233]), .Z(n32691) );
  XNOR U33233 ( .A(b[1]), .B(n32691), .Z(n32693) );
  IV U33234 ( .A(a[232]), .Z(n37079) );
  NANDN U33235 ( .A(n37079), .B(n1049), .Z(n32692) );
  AND U33236 ( .A(n32693), .B(n32692), .Z(n32735) );
  XNOR U33237 ( .A(n32734), .B(n32735), .Z(n32756) );
  NANDN U33238 ( .A(n32694), .B(n38205), .Z(n32696) );
  XNOR U33239 ( .A(b[23]), .B(a[211]), .Z(n32827) );
  OR U33240 ( .A(n32827), .B(n38268), .Z(n32695) );
  NAND U33241 ( .A(n32696), .B(n32695), .Z(n32797) );
  XOR U33242 ( .A(b[7]), .B(a[227]), .Z(n32830) );
  NAND U33243 ( .A(n32830), .B(n36701), .Z(n32699) );
  NANDN U33244 ( .A(n32697), .B(n36702), .Z(n32698) );
  NAND U33245 ( .A(n32699), .B(n32698), .Z(n32794) );
  XOR U33246 ( .A(b[25]), .B(a[209]), .Z(n32833) );
  NAND U33247 ( .A(n32833), .B(n38325), .Z(n32702) );
  NAND U33248 ( .A(n32700), .B(n38326), .Z(n32701) );
  AND U33249 ( .A(n32702), .B(n32701), .Z(n32795) );
  XNOR U33250 ( .A(n32794), .B(n32795), .Z(n32796) );
  XNOR U33251 ( .A(n32797), .B(n32796), .Z(n32757) );
  XOR U33252 ( .A(n32759), .B(n32758), .Z(n32787) );
  XNOR U33253 ( .A(n32786), .B(n32787), .Z(n32842) );
  XNOR U33254 ( .A(n32843), .B(n32842), .Z(n32845) );
  XNOR U33255 ( .A(n32844), .B(n32845), .Z(n32854) );
  XOR U33256 ( .A(n32855), .B(n32854), .Z(n32857) );
  NANDN U33257 ( .A(n32704), .B(n32703), .Z(n32708) );
  OR U33258 ( .A(n32706), .B(n32705), .Z(n32707) );
  NAND U33259 ( .A(n32708), .B(n32707), .Z(n32848) );
  NAND U33260 ( .A(n32710), .B(n32709), .Z(n32714) );
  NANDN U33261 ( .A(n32712), .B(n32711), .Z(n32713) );
  NAND U33262 ( .A(n32714), .B(n32713), .Z(n32849) );
  XNOR U33263 ( .A(n32848), .B(n32849), .Z(n32850) );
  XOR U33264 ( .A(n32851), .B(n32850), .Z(n32729) );
  XOR U33265 ( .A(n32728), .B(n32729), .Z(n32720) );
  XOR U33266 ( .A(n32721), .B(n32720), .Z(n32722) );
  XNOR U33267 ( .A(n32723), .B(n32722), .Z(n32860) );
  XNOR U33268 ( .A(n32860), .B(sreg[457]), .Z(n32862) );
  NAND U33269 ( .A(n32715), .B(sreg[456]), .Z(n32719) );
  OR U33270 ( .A(n32717), .B(n32716), .Z(n32718) );
  AND U33271 ( .A(n32719), .B(n32718), .Z(n32861) );
  XOR U33272 ( .A(n32862), .B(n32861), .Z(c[457]) );
  NAND U33273 ( .A(n32721), .B(n32720), .Z(n32725) );
  NAND U33274 ( .A(n32723), .B(n32722), .Z(n32724) );
  NAND U33275 ( .A(n32725), .B(n32724), .Z(n32868) );
  NANDN U33276 ( .A(n32727), .B(n32726), .Z(n32731) );
  NAND U33277 ( .A(n32729), .B(n32728), .Z(n32730) );
  NAND U33278 ( .A(n32731), .B(n32730), .Z(n32866) );
  OR U33279 ( .A(n32733), .B(n32732), .Z(n32737) );
  NANDN U33280 ( .A(n32735), .B(n32734), .Z(n32736) );
  NAND U33281 ( .A(n32737), .B(n32736), .Z(n32938) );
  XNOR U33282 ( .A(b[19]), .B(a[216]), .Z(n32907) );
  NANDN U33283 ( .A(n32907), .B(n37934), .Z(n32740) );
  NANDN U33284 ( .A(n32738), .B(n37935), .Z(n32739) );
  NAND U33285 ( .A(n32740), .B(n32739), .Z(n32950) );
  XOR U33286 ( .A(b[27]), .B(a[208]), .Z(n32910) );
  NAND U33287 ( .A(n38423), .B(n32910), .Z(n32743) );
  NAND U33288 ( .A(n32741), .B(n38424), .Z(n32742) );
  NAND U33289 ( .A(n32743), .B(n32742), .Z(n32947) );
  XOR U33290 ( .A(b[5]), .B(n36333), .Z(n32913) );
  NANDN U33291 ( .A(n32913), .B(n36587), .Z(n32746) );
  NANDN U33292 ( .A(n32744), .B(n36588), .Z(n32745) );
  AND U33293 ( .A(n32746), .B(n32745), .Z(n32948) );
  XNOR U33294 ( .A(n32947), .B(n32948), .Z(n32949) );
  XNOR U33295 ( .A(n32950), .B(n32949), .Z(n32935) );
  NANDN U33296 ( .A(n32747), .B(n37762), .Z(n32749) );
  XOR U33297 ( .A(b[17]), .B(a[218]), .Z(n32916) );
  NAND U33298 ( .A(n32916), .B(n37764), .Z(n32748) );
  NAND U33299 ( .A(n32749), .B(n32748), .Z(n32891) );
  XOR U33300 ( .A(b[31]), .B(n33130), .Z(n32919) );
  NANDN U33301 ( .A(n32919), .B(n38552), .Z(n32752) );
  NANDN U33302 ( .A(n32750), .B(n38553), .Z(n32751) );
  AND U33303 ( .A(n32752), .B(n32751), .Z(n32889) );
  OR U33304 ( .A(n32753), .B(n36105), .Z(n32755) );
  XOR U33305 ( .A(a[232]), .B(n1050), .Z(n32922) );
  NANDN U33306 ( .A(n32922), .B(n36107), .Z(n32754) );
  AND U33307 ( .A(n32755), .B(n32754), .Z(n32890) );
  XOR U33308 ( .A(n32891), .B(n32892), .Z(n32936) );
  XOR U33309 ( .A(n32935), .B(n32936), .Z(n32937) );
  XOR U33310 ( .A(n32938), .B(n32937), .Z(n32989) );
  OR U33311 ( .A(n32757), .B(n32756), .Z(n32761) );
  NANDN U33312 ( .A(n32759), .B(n32758), .Z(n32760) );
  NAND U33313 ( .A(n32761), .B(n32760), .Z(n32990) );
  XNOR U33314 ( .A(n32989), .B(n32990), .Z(n32991) );
  NANDN U33315 ( .A(n32763), .B(n32762), .Z(n32767) );
  NAND U33316 ( .A(n32765), .B(n32764), .Z(n32766) );
  NAND U33317 ( .A(n32767), .B(n32766), .Z(n32928) );
  OR U33318 ( .A(n32769), .B(n32768), .Z(n32773) );
  NANDN U33319 ( .A(n32771), .B(n32770), .Z(n32772) );
  NAND U33320 ( .A(n32773), .B(n32772), .Z(n32926) );
  XNOR U33321 ( .A(n32926), .B(n32925), .Z(n32927) );
  XOR U33322 ( .A(n32928), .B(n32927), .Z(n32992) );
  XOR U33323 ( .A(n32991), .B(n32992), .Z(n33004) );
  OR U33324 ( .A(n32779), .B(n32778), .Z(n32783) );
  NAND U33325 ( .A(n32781), .B(n32780), .Z(n32782) );
  NAND U33326 ( .A(n32783), .B(n32782), .Z(n33002) );
  NANDN U33327 ( .A(n32785), .B(n32784), .Z(n32789) );
  NANDN U33328 ( .A(n32787), .B(n32786), .Z(n32788) );
  NAND U33329 ( .A(n32789), .B(n32788), .Z(n32985) );
  NANDN U33330 ( .A(n32795), .B(n32794), .Z(n32799) );
  NAND U33331 ( .A(n32797), .B(n32796), .Z(n32798) );
  NAND U33332 ( .A(n32799), .B(n32798), .Z(n32929) );
  NANDN U33333 ( .A(n32801), .B(n32800), .Z(n32805) );
  NAND U33334 ( .A(n32803), .B(n32802), .Z(n32804) );
  AND U33335 ( .A(n32805), .B(n32804), .Z(n32930) );
  XNOR U33336 ( .A(n32929), .B(n32930), .Z(n32931) );
  XOR U33337 ( .A(b[9]), .B(n36280), .Z(n32953) );
  NANDN U33338 ( .A(n32953), .B(n36925), .Z(n32808) );
  NANDN U33339 ( .A(n32806), .B(n36926), .Z(n32807) );
  NAND U33340 ( .A(n32808), .B(n32807), .Z(n32897) );
  XNOR U33341 ( .A(b[15]), .B(a[220]), .Z(n32956) );
  OR U33342 ( .A(n32956), .B(n37665), .Z(n32811) );
  NANDN U33343 ( .A(n32809), .B(n37604), .Z(n32810) );
  AND U33344 ( .A(n32811), .B(n32810), .Z(n32895) );
  XNOR U33345 ( .A(b[21]), .B(a[214]), .Z(n32959) );
  NANDN U33346 ( .A(n32959), .B(n38101), .Z(n32814) );
  NANDN U33347 ( .A(n32812), .B(n38102), .Z(n32813) );
  AND U33348 ( .A(n32814), .B(n32813), .Z(n32896) );
  XOR U33349 ( .A(n32897), .B(n32898), .Z(n32886) );
  XNOR U33350 ( .A(b[11]), .B(a[224]), .Z(n32962) );
  OR U33351 ( .A(n32962), .B(n37311), .Z(n32817) );
  NANDN U33352 ( .A(n32815), .B(n37218), .Z(n32816) );
  NAND U33353 ( .A(n32817), .B(n32816), .Z(n32884) );
  XOR U33354 ( .A(n1053), .B(a[222]), .Z(n32965) );
  NANDN U33355 ( .A(n32965), .B(n37424), .Z(n32820) );
  NANDN U33356 ( .A(n32818), .B(n37425), .Z(n32819) );
  NAND U33357 ( .A(n32820), .B(n32819), .Z(n32883) );
  XOR U33358 ( .A(n32886), .B(n32885), .Z(n32880) );
  NANDN U33359 ( .A(n1049), .B(a[234]), .Z(n32821) );
  XNOR U33360 ( .A(b[1]), .B(n32821), .Z(n32823) );
  IV U33361 ( .A(a[233]), .Z(n37184) );
  NANDN U33362 ( .A(n37184), .B(n1049), .Z(n32822) );
  AND U33363 ( .A(n32823), .B(n32822), .Z(n32903) );
  NAND U33364 ( .A(n32824), .B(n38490), .Z(n32826) );
  XNOR U33365 ( .A(n1058), .B(a[206]), .Z(n32971) );
  NANDN U33366 ( .A(n1048), .B(n32971), .Z(n32825) );
  NAND U33367 ( .A(n32826), .B(n32825), .Z(n32901) );
  NANDN U33368 ( .A(n1059), .B(a[202]), .Z(n32902) );
  XNOR U33369 ( .A(n32901), .B(n32902), .Z(n32904) );
  XNOR U33370 ( .A(n32903), .B(n32904), .Z(n32878) );
  NANDN U33371 ( .A(n32827), .B(n38205), .Z(n32829) );
  XNOR U33372 ( .A(b[23]), .B(a[212]), .Z(n32974) );
  OR U33373 ( .A(n32974), .B(n38268), .Z(n32828) );
  NAND U33374 ( .A(n32829), .B(n32828), .Z(n32944) );
  XNOR U33375 ( .A(b[7]), .B(a[228]), .Z(n32977) );
  NANDN U33376 ( .A(n32977), .B(n36701), .Z(n32832) );
  NAND U33377 ( .A(n32830), .B(n36702), .Z(n32831) );
  NAND U33378 ( .A(n32832), .B(n32831), .Z(n32941) );
  XOR U33379 ( .A(b[25]), .B(a[210]), .Z(n32980) );
  NAND U33380 ( .A(n32980), .B(n38325), .Z(n32835) );
  NAND U33381 ( .A(n32833), .B(n38326), .Z(n32834) );
  AND U33382 ( .A(n32835), .B(n32834), .Z(n32942) );
  XNOR U33383 ( .A(n32941), .B(n32942), .Z(n32943) );
  XOR U33384 ( .A(n32944), .B(n32943), .Z(n32877) );
  XOR U33385 ( .A(n32880), .B(n32879), .Z(n32932) );
  XNOR U33386 ( .A(n32931), .B(n32932), .Z(n32983) );
  XNOR U33387 ( .A(n32984), .B(n32983), .Z(n32986) );
  XNOR U33388 ( .A(n32985), .B(n32986), .Z(n33001) );
  XOR U33389 ( .A(n33002), .B(n33001), .Z(n33003) );
  XNOR U33390 ( .A(n33004), .B(n33003), .Z(n32998) );
  NANDN U33391 ( .A(n32837), .B(n32836), .Z(n32841) );
  OR U33392 ( .A(n32839), .B(n32838), .Z(n32840) );
  NAND U33393 ( .A(n32841), .B(n32840), .Z(n32995) );
  NAND U33394 ( .A(n32843), .B(n32842), .Z(n32847) );
  NANDN U33395 ( .A(n32845), .B(n32844), .Z(n32846) );
  NAND U33396 ( .A(n32847), .B(n32846), .Z(n32996) );
  XNOR U33397 ( .A(n32995), .B(n32996), .Z(n32997) );
  XOR U33398 ( .A(n32998), .B(n32997), .Z(n32873) );
  NANDN U33399 ( .A(n32849), .B(n32848), .Z(n32853) );
  NAND U33400 ( .A(n32851), .B(n32850), .Z(n32852) );
  NAND U33401 ( .A(n32853), .B(n32852), .Z(n32871) );
  NANDN U33402 ( .A(n32855), .B(n32854), .Z(n32859) );
  OR U33403 ( .A(n32857), .B(n32856), .Z(n32858) );
  NAND U33404 ( .A(n32859), .B(n32858), .Z(n32872) );
  XNOR U33405 ( .A(n32871), .B(n32872), .Z(n32874) );
  XOR U33406 ( .A(n32873), .B(n32874), .Z(n32865) );
  XOR U33407 ( .A(n32866), .B(n32865), .Z(n32867) );
  XNOR U33408 ( .A(n32868), .B(n32867), .Z(n33007) );
  XNOR U33409 ( .A(n33007), .B(sreg[458]), .Z(n33009) );
  NAND U33410 ( .A(n32860), .B(sreg[457]), .Z(n32864) );
  OR U33411 ( .A(n32862), .B(n32861), .Z(n32863) );
  AND U33412 ( .A(n32864), .B(n32863), .Z(n33008) );
  XOR U33413 ( .A(n33009), .B(n33008), .Z(c[458]) );
  NAND U33414 ( .A(n32866), .B(n32865), .Z(n32870) );
  NAND U33415 ( .A(n32868), .B(n32867), .Z(n32869) );
  NAND U33416 ( .A(n32870), .B(n32869), .Z(n33015) );
  NANDN U33417 ( .A(n32872), .B(n32871), .Z(n32876) );
  NAND U33418 ( .A(n32874), .B(n32873), .Z(n32875) );
  NAND U33419 ( .A(n32876), .B(n32875), .Z(n33013) );
  NANDN U33420 ( .A(n32878), .B(n32877), .Z(n32882) );
  NANDN U33421 ( .A(n32880), .B(n32879), .Z(n32881) );
  NAND U33422 ( .A(n32882), .B(n32881), .Z(n33146) );
  OR U33423 ( .A(n32884), .B(n32883), .Z(n32888) );
  NAND U33424 ( .A(n32886), .B(n32885), .Z(n32887) );
  NAND U33425 ( .A(n32888), .B(n32887), .Z(n33084) );
  OR U33426 ( .A(n32890), .B(n32889), .Z(n32894) );
  NANDN U33427 ( .A(n32892), .B(n32891), .Z(n32893) );
  NAND U33428 ( .A(n32894), .B(n32893), .Z(n33083) );
  OR U33429 ( .A(n32896), .B(n32895), .Z(n32900) );
  NANDN U33430 ( .A(n32898), .B(n32897), .Z(n32899) );
  NAND U33431 ( .A(n32900), .B(n32899), .Z(n33082) );
  XOR U33432 ( .A(n33084), .B(n33085), .Z(n33143) );
  NANDN U33433 ( .A(n32902), .B(n32901), .Z(n32906) );
  NAND U33434 ( .A(n32904), .B(n32903), .Z(n32905) );
  NAND U33435 ( .A(n32906), .B(n32905), .Z(n33097) );
  XOR U33436 ( .A(b[19]), .B(n34670), .Z(n33040) );
  NANDN U33437 ( .A(n33040), .B(n37934), .Z(n32909) );
  NANDN U33438 ( .A(n32907), .B(n37935), .Z(n32908) );
  NAND U33439 ( .A(n32909), .B(n32908), .Z(n33109) );
  XOR U33440 ( .A(b[27]), .B(a[209]), .Z(n33043) );
  NAND U33441 ( .A(n38423), .B(n33043), .Z(n32912) );
  NAND U33442 ( .A(n32910), .B(n38424), .Z(n32911) );
  NAND U33443 ( .A(n32912), .B(n32911), .Z(n33106) );
  XOR U33444 ( .A(b[5]), .B(n36934), .Z(n33046) );
  NANDN U33445 ( .A(n33046), .B(n36587), .Z(n32915) );
  NANDN U33446 ( .A(n32913), .B(n36588), .Z(n32914) );
  AND U33447 ( .A(n32915), .B(n32914), .Z(n33107) );
  XNOR U33448 ( .A(n33106), .B(n33107), .Z(n33108) );
  XNOR U33449 ( .A(n33109), .B(n33108), .Z(n33095) );
  NAND U33450 ( .A(n32916), .B(n37762), .Z(n32918) );
  XOR U33451 ( .A(b[17]), .B(a[219]), .Z(n33049) );
  NAND U33452 ( .A(n33049), .B(n37764), .Z(n32917) );
  NAND U33453 ( .A(n32918), .B(n32917), .Z(n33067) );
  XNOR U33454 ( .A(b[31]), .B(a[205]), .Z(n33052) );
  NANDN U33455 ( .A(n33052), .B(n38552), .Z(n32921) );
  NANDN U33456 ( .A(n32919), .B(n38553), .Z(n32920) );
  NAND U33457 ( .A(n32921), .B(n32920), .Z(n33064) );
  OR U33458 ( .A(n32922), .B(n36105), .Z(n32924) );
  XOR U33459 ( .A(a[233]), .B(n1050), .Z(n33055) );
  NANDN U33460 ( .A(n33055), .B(n36107), .Z(n32923) );
  AND U33461 ( .A(n32924), .B(n32923), .Z(n33065) );
  XNOR U33462 ( .A(n33064), .B(n33065), .Z(n33066) );
  XOR U33463 ( .A(n33067), .B(n33066), .Z(n33094) );
  XNOR U33464 ( .A(n33095), .B(n33094), .Z(n33096) );
  XNOR U33465 ( .A(n33097), .B(n33096), .Z(n33144) );
  XNOR U33466 ( .A(n33143), .B(n33144), .Z(n33145) );
  XNOR U33467 ( .A(n33146), .B(n33145), .Z(n33024) );
  NANDN U33468 ( .A(n32930), .B(n32929), .Z(n32934) );
  NANDN U33469 ( .A(n32932), .B(n32931), .Z(n32933) );
  NAND U33470 ( .A(n32934), .B(n32933), .Z(n33149) );
  OR U33471 ( .A(n32936), .B(n32935), .Z(n32940) );
  NANDN U33472 ( .A(n32938), .B(n32937), .Z(n32939) );
  NAND U33473 ( .A(n32940), .B(n32939), .Z(n33148) );
  NANDN U33474 ( .A(n32942), .B(n32941), .Z(n32946) );
  NAND U33475 ( .A(n32944), .B(n32943), .Z(n32945) );
  NAND U33476 ( .A(n32946), .B(n32945), .Z(n33088) );
  NANDN U33477 ( .A(n32948), .B(n32947), .Z(n32952) );
  NAND U33478 ( .A(n32950), .B(n32949), .Z(n32951) );
  AND U33479 ( .A(n32952), .B(n32951), .Z(n33089) );
  XNOR U33480 ( .A(n33088), .B(n33089), .Z(n33090) );
  XNOR U33481 ( .A(b[9]), .B(a[227]), .Z(n33112) );
  NANDN U33482 ( .A(n33112), .B(n36925), .Z(n32955) );
  NANDN U33483 ( .A(n32953), .B(n36926), .Z(n32954) );
  NAND U33484 ( .A(n32955), .B(n32954), .Z(n33072) );
  XNOR U33485 ( .A(b[15]), .B(a[221]), .Z(n33115) );
  OR U33486 ( .A(n33115), .B(n37665), .Z(n32958) );
  NANDN U33487 ( .A(n32956), .B(n37604), .Z(n32957) );
  AND U33488 ( .A(n32958), .B(n32957), .Z(n33070) );
  XOR U33489 ( .A(b[21]), .B(n34725), .Z(n33118) );
  NANDN U33490 ( .A(n33118), .B(n38101), .Z(n32961) );
  NANDN U33491 ( .A(n32959), .B(n38102), .Z(n32960) );
  AND U33492 ( .A(n32961), .B(n32960), .Z(n33071) );
  XOR U33493 ( .A(n33072), .B(n33073), .Z(n33061) );
  XOR U33494 ( .A(b[11]), .B(n36167), .Z(n33121) );
  OR U33495 ( .A(n33121), .B(n37311), .Z(n32964) );
  NANDN U33496 ( .A(n32962), .B(n37218), .Z(n32963) );
  NAND U33497 ( .A(n32964), .B(n32963), .Z(n33059) );
  XOR U33498 ( .A(n1053), .B(a[223]), .Z(n33124) );
  NANDN U33499 ( .A(n33124), .B(n37424), .Z(n32967) );
  NANDN U33500 ( .A(n32965), .B(n37425), .Z(n32966) );
  AND U33501 ( .A(n32967), .B(n32966), .Z(n33058) );
  XNOR U33502 ( .A(n33059), .B(n33058), .Z(n33060) );
  XOR U33503 ( .A(n33061), .B(n33060), .Z(n33078) );
  NANDN U33504 ( .A(n1049), .B(a[235]), .Z(n32968) );
  XNOR U33505 ( .A(b[1]), .B(n32968), .Z(n32970) );
  IV U33506 ( .A(a[234]), .Z(n37080) );
  NANDN U33507 ( .A(n37080), .B(n1049), .Z(n32969) );
  AND U33508 ( .A(n32970), .B(n32969), .Z(n33036) );
  NAND U33509 ( .A(n38490), .B(n32971), .Z(n32973) );
  XNOR U33510 ( .A(b[29]), .B(a[207]), .Z(n33131) );
  OR U33511 ( .A(n33131), .B(n1048), .Z(n32972) );
  NAND U33512 ( .A(n32973), .B(n32972), .Z(n33034) );
  NANDN U33513 ( .A(n1059), .B(a[203]), .Z(n33035) );
  XNOR U33514 ( .A(n33034), .B(n33035), .Z(n33037) );
  XOR U33515 ( .A(n33036), .B(n33037), .Z(n33076) );
  NANDN U33516 ( .A(n32974), .B(n38205), .Z(n32976) );
  XNOR U33517 ( .A(b[23]), .B(a[213]), .Z(n33134) );
  OR U33518 ( .A(n33134), .B(n38268), .Z(n32975) );
  NAND U33519 ( .A(n32976), .B(n32975), .Z(n33103) );
  XOR U33520 ( .A(b[7]), .B(a[229]), .Z(n33137) );
  NAND U33521 ( .A(n33137), .B(n36701), .Z(n32979) );
  NANDN U33522 ( .A(n32977), .B(n36702), .Z(n32978) );
  NAND U33523 ( .A(n32979), .B(n32978), .Z(n33100) );
  XOR U33524 ( .A(b[25]), .B(a[211]), .Z(n33140) );
  NAND U33525 ( .A(n33140), .B(n38325), .Z(n32982) );
  NAND U33526 ( .A(n32980), .B(n38326), .Z(n32981) );
  AND U33527 ( .A(n32982), .B(n32981), .Z(n33101) );
  XNOR U33528 ( .A(n33100), .B(n33101), .Z(n33102) );
  XNOR U33529 ( .A(n33103), .B(n33102), .Z(n33077) );
  XOR U33530 ( .A(n33076), .B(n33077), .Z(n33079) );
  XNOR U33531 ( .A(n33078), .B(n33079), .Z(n33091) );
  XNOR U33532 ( .A(n33090), .B(n33091), .Z(n33147) );
  XNOR U33533 ( .A(n33148), .B(n33147), .Z(n33150) );
  XNOR U33534 ( .A(n33149), .B(n33150), .Z(n33023) );
  XOR U33535 ( .A(n33022), .B(n33023), .Z(n33025) );
  XNOR U33536 ( .A(n33024), .B(n33025), .Z(n33031) );
  NAND U33537 ( .A(n32984), .B(n32983), .Z(n32988) );
  NANDN U33538 ( .A(n32986), .B(n32985), .Z(n32987) );
  NAND U33539 ( .A(n32988), .B(n32987), .Z(n33028) );
  NANDN U33540 ( .A(n32990), .B(n32989), .Z(n32994) );
  NAND U33541 ( .A(n32992), .B(n32991), .Z(n32993) );
  NAND U33542 ( .A(n32994), .B(n32993), .Z(n33029) );
  XNOR U33543 ( .A(n33028), .B(n33029), .Z(n33030) );
  XNOR U33544 ( .A(n33031), .B(n33030), .Z(n33019) );
  NANDN U33545 ( .A(n32996), .B(n32995), .Z(n33000) );
  NAND U33546 ( .A(n32998), .B(n32997), .Z(n32999) );
  NAND U33547 ( .A(n33000), .B(n32999), .Z(n33016) );
  NANDN U33548 ( .A(n33002), .B(n33001), .Z(n33006) );
  OR U33549 ( .A(n33004), .B(n33003), .Z(n33005) );
  NAND U33550 ( .A(n33006), .B(n33005), .Z(n33017) );
  XNOR U33551 ( .A(n33016), .B(n33017), .Z(n33018) );
  XNOR U33552 ( .A(n33019), .B(n33018), .Z(n33012) );
  XOR U33553 ( .A(n33013), .B(n33012), .Z(n33014) );
  XNOR U33554 ( .A(n33015), .B(n33014), .Z(n33153) );
  XNOR U33555 ( .A(n33153), .B(sreg[459]), .Z(n33155) );
  NAND U33556 ( .A(n33007), .B(sreg[458]), .Z(n33011) );
  OR U33557 ( .A(n33009), .B(n33008), .Z(n33010) );
  AND U33558 ( .A(n33011), .B(n33010), .Z(n33154) );
  XOR U33559 ( .A(n33155), .B(n33154), .Z(c[459]) );
  NANDN U33560 ( .A(n33017), .B(n33016), .Z(n33021) );
  NANDN U33561 ( .A(n33019), .B(n33018), .Z(n33020) );
  NAND U33562 ( .A(n33021), .B(n33020), .Z(n33159) );
  NANDN U33563 ( .A(n33023), .B(n33022), .Z(n33027) );
  NANDN U33564 ( .A(n33025), .B(n33024), .Z(n33026) );
  NAND U33565 ( .A(n33027), .B(n33026), .Z(n33164) );
  NANDN U33566 ( .A(n33029), .B(n33028), .Z(n33033) );
  NANDN U33567 ( .A(n33031), .B(n33030), .Z(n33032) );
  NAND U33568 ( .A(n33033), .B(n33032), .Z(n33165) );
  XNOR U33569 ( .A(n33164), .B(n33165), .Z(n33166) );
  NANDN U33570 ( .A(n33035), .B(n33034), .Z(n33039) );
  NAND U33571 ( .A(n33037), .B(n33036), .Z(n33038) );
  NAND U33572 ( .A(n33039), .B(n33038), .Z(n33233) );
  XNOR U33573 ( .A(b[19]), .B(a[218]), .Z(n33200) );
  NANDN U33574 ( .A(n33200), .B(n37934), .Z(n33042) );
  NANDN U33575 ( .A(n33040), .B(n37935), .Z(n33041) );
  NAND U33576 ( .A(n33042), .B(n33041), .Z(n33245) );
  XOR U33577 ( .A(b[27]), .B(a[210]), .Z(n33203) );
  NAND U33578 ( .A(n38423), .B(n33203), .Z(n33045) );
  NAND U33579 ( .A(n33043), .B(n38424), .Z(n33044) );
  NAND U33580 ( .A(n33045), .B(n33044), .Z(n33242) );
  XOR U33581 ( .A(a[232]), .B(n1051), .Z(n33206) );
  NANDN U33582 ( .A(n33206), .B(n36587), .Z(n33048) );
  NANDN U33583 ( .A(n33046), .B(n36588), .Z(n33047) );
  AND U33584 ( .A(n33048), .B(n33047), .Z(n33243) );
  XNOR U33585 ( .A(n33242), .B(n33243), .Z(n33244) );
  XNOR U33586 ( .A(n33245), .B(n33244), .Z(n33230) );
  NAND U33587 ( .A(n33049), .B(n37762), .Z(n33051) );
  XOR U33588 ( .A(b[17]), .B(a[220]), .Z(n33209) );
  NAND U33589 ( .A(n33209), .B(n37764), .Z(n33050) );
  NAND U33590 ( .A(n33051), .B(n33050), .Z(n33184) );
  XNOR U33591 ( .A(b[31]), .B(a[206]), .Z(n33212) );
  NANDN U33592 ( .A(n33212), .B(n38552), .Z(n33054) );
  NANDN U33593 ( .A(n33052), .B(n38553), .Z(n33053) );
  AND U33594 ( .A(n33054), .B(n33053), .Z(n33182) );
  OR U33595 ( .A(n33055), .B(n36105), .Z(n33057) );
  XOR U33596 ( .A(a[234]), .B(n1050), .Z(n33215) );
  NANDN U33597 ( .A(n33215), .B(n36107), .Z(n33056) );
  AND U33598 ( .A(n33057), .B(n33056), .Z(n33183) );
  XOR U33599 ( .A(n33184), .B(n33185), .Z(n33231) );
  XOR U33600 ( .A(n33230), .B(n33231), .Z(n33232) );
  XNOR U33601 ( .A(n33233), .B(n33232), .Z(n33278) );
  NANDN U33602 ( .A(n33059), .B(n33058), .Z(n33063) );
  NAND U33603 ( .A(n33061), .B(n33060), .Z(n33062) );
  NAND U33604 ( .A(n33063), .B(n33062), .Z(n33221) );
  NANDN U33605 ( .A(n33065), .B(n33064), .Z(n33069) );
  NAND U33606 ( .A(n33067), .B(n33066), .Z(n33068) );
  NAND U33607 ( .A(n33069), .B(n33068), .Z(n33219) );
  OR U33608 ( .A(n33071), .B(n33070), .Z(n33075) );
  NANDN U33609 ( .A(n33073), .B(n33072), .Z(n33074) );
  NAND U33610 ( .A(n33075), .B(n33074), .Z(n33218) );
  XNOR U33611 ( .A(n33221), .B(n33220), .Z(n33279) );
  XOR U33612 ( .A(n33278), .B(n33279), .Z(n33281) );
  NANDN U33613 ( .A(n33077), .B(n33076), .Z(n33081) );
  OR U33614 ( .A(n33079), .B(n33078), .Z(n33080) );
  NAND U33615 ( .A(n33081), .B(n33080), .Z(n33280) );
  XOR U33616 ( .A(n33281), .B(n33280), .Z(n33298) );
  OR U33617 ( .A(n33083), .B(n33082), .Z(n33087) );
  NANDN U33618 ( .A(n33085), .B(n33084), .Z(n33086) );
  NAND U33619 ( .A(n33087), .B(n33086), .Z(n33297) );
  NANDN U33620 ( .A(n33089), .B(n33088), .Z(n33093) );
  NANDN U33621 ( .A(n33091), .B(n33090), .Z(n33092) );
  NAND U33622 ( .A(n33093), .B(n33092), .Z(n33286) );
  NANDN U33623 ( .A(n33095), .B(n33094), .Z(n33099) );
  NAND U33624 ( .A(n33097), .B(n33096), .Z(n33098) );
  NAND U33625 ( .A(n33099), .B(n33098), .Z(n33285) );
  NANDN U33626 ( .A(n33101), .B(n33100), .Z(n33105) );
  NAND U33627 ( .A(n33103), .B(n33102), .Z(n33104) );
  NAND U33628 ( .A(n33105), .B(n33104), .Z(n33224) );
  NANDN U33629 ( .A(n33107), .B(n33106), .Z(n33111) );
  NAND U33630 ( .A(n33109), .B(n33108), .Z(n33110) );
  AND U33631 ( .A(n33111), .B(n33110), .Z(n33225) );
  XNOR U33632 ( .A(n33224), .B(n33225), .Z(n33226) );
  XOR U33633 ( .A(b[9]), .B(n36592), .Z(n33248) );
  NANDN U33634 ( .A(n33248), .B(n36925), .Z(n33114) );
  NANDN U33635 ( .A(n33112), .B(n36926), .Z(n33113) );
  NAND U33636 ( .A(n33114), .B(n33113), .Z(n33190) );
  XOR U33637 ( .A(b[15]), .B(n35381), .Z(n33251) );
  OR U33638 ( .A(n33251), .B(n37665), .Z(n33117) );
  NANDN U33639 ( .A(n33115), .B(n37604), .Z(n33116) );
  AND U33640 ( .A(n33117), .B(n33116), .Z(n33188) );
  XNOR U33641 ( .A(b[21]), .B(a[216]), .Z(n33254) );
  NANDN U33642 ( .A(n33254), .B(n38101), .Z(n33120) );
  NANDN U33643 ( .A(n33118), .B(n38102), .Z(n33119) );
  AND U33644 ( .A(n33120), .B(n33119), .Z(n33189) );
  XOR U33645 ( .A(n33190), .B(n33191), .Z(n33179) );
  XOR U33646 ( .A(b[11]), .B(n36280), .Z(n33257) );
  OR U33647 ( .A(n33257), .B(n37311), .Z(n33123) );
  NANDN U33648 ( .A(n33121), .B(n37218), .Z(n33122) );
  NAND U33649 ( .A(n33123), .B(n33122), .Z(n33177) );
  XOR U33650 ( .A(n1053), .B(a[224]), .Z(n33260) );
  NANDN U33651 ( .A(n33260), .B(n37424), .Z(n33126) );
  NANDN U33652 ( .A(n33124), .B(n37425), .Z(n33125) );
  NAND U33653 ( .A(n33126), .B(n33125), .Z(n33176) );
  XOR U33654 ( .A(n33179), .B(n33178), .Z(n33173) );
  NANDN U33655 ( .A(n1049), .B(a[236]), .Z(n33127) );
  XNOR U33656 ( .A(b[1]), .B(n33127), .Z(n33129) );
  IV U33657 ( .A(a[235]), .Z(n37420) );
  NANDN U33658 ( .A(n37420), .B(n1049), .Z(n33128) );
  AND U33659 ( .A(n33129), .B(n33128), .Z(n33197) );
  ANDN U33660 ( .B(b[31]), .A(n33130), .Z(n33194) );
  NANDN U33661 ( .A(n33131), .B(n38490), .Z(n33133) );
  XNOR U33662 ( .A(n1058), .B(a[208]), .Z(n33266) );
  NANDN U33663 ( .A(n1048), .B(n33266), .Z(n33132) );
  NAND U33664 ( .A(n33133), .B(n33132), .Z(n33195) );
  XOR U33665 ( .A(n33194), .B(n33195), .Z(n33196) );
  XNOR U33666 ( .A(n33197), .B(n33196), .Z(n33170) );
  NANDN U33667 ( .A(n33134), .B(n38205), .Z(n33136) );
  XNOR U33668 ( .A(b[23]), .B(a[214]), .Z(n33269) );
  OR U33669 ( .A(n33269), .B(n38268), .Z(n33135) );
  NAND U33670 ( .A(n33136), .B(n33135), .Z(n33239) );
  XNOR U33671 ( .A(b[7]), .B(a[230]), .Z(n33272) );
  NANDN U33672 ( .A(n33272), .B(n36701), .Z(n33139) );
  NAND U33673 ( .A(n33137), .B(n36702), .Z(n33138) );
  NAND U33674 ( .A(n33139), .B(n33138), .Z(n33236) );
  XOR U33675 ( .A(b[25]), .B(a[212]), .Z(n33275) );
  NAND U33676 ( .A(n33275), .B(n38325), .Z(n33142) );
  NAND U33677 ( .A(n33140), .B(n38326), .Z(n33141) );
  AND U33678 ( .A(n33142), .B(n33141), .Z(n33237) );
  XNOR U33679 ( .A(n33236), .B(n33237), .Z(n33238) );
  XNOR U33680 ( .A(n33239), .B(n33238), .Z(n33171) );
  XOR U33681 ( .A(n33173), .B(n33172), .Z(n33227) );
  XNOR U33682 ( .A(n33226), .B(n33227), .Z(n33284) );
  XNOR U33683 ( .A(n33285), .B(n33284), .Z(n33287) );
  XNOR U33684 ( .A(n33286), .B(n33287), .Z(n33296) );
  XOR U33685 ( .A(n33297), .B(n33296), .Z(n33299) );
  NAND U33686 ( .A(n33148), .B(n33147), .Z(n33152) );
  NANDN U33687 ( .A(n33150), .B(n33149), .Z(n33151) );
  AND U33688 ( .A(n33152), .B(n33151), .Z(n33290) );
  XNOR U33689 ( .A(n33291), .B(n33290), .Z(n33292) );
  XOR U33690 ( .A(n33293), .B(n33292), .Z(n33167) );
  XOR U33691 ( .A(n33166), .B(n33167), .Z(n33158) );
  XOR U33692 ( .A(n33159), .B(n33158), .Z(n33160) );
  XNOR U33693 ( .A(n33161), .B(n33160), .Z(n33302) );
  XNOR U33694 ( .A(n33302), .B(sreg[460]), .Z(n33304) );
  NAND U33695 ( .A(n33153), .B(sreg[459]), .Z(n33157) );
  OR U33696 ( .A(n33155), .B(n33154), .Z(n33156) );
  AND U33697 ( .A(n33157), .B(n33156), .Z(n33303) );
  XOR U33698 ( .A(n33304), .B(n33303), .Z(c[460]) );
  NAND U33699 ( .A(n33159), .B(n33158), .Z(n33163) );
  NAND U33700 ( .A(n33161), .B(n33160), .Z(n33162) );
  NAND U33701 ( .A(n33163), .B(n33162), .Z(n33310) );
  NANDN U33702 ( .A(n33165), .B(n33164), .Z(n33169) );
  NAND U33703 ( .A(n33167), .B(n33166), .Z(n33168) );
  NAND U33704 ( .A(n33169), .B(n33168), .Z(n33308) );
  OR U33705 ( .A(n33171), .B(n33170), .Z(n33175) );
  NANDN U33706 ( .A(n33173), .B(n33172), .Z(n33174) );
  NAND U33707 ( .A(n33175), .B(n33174), .Z(n33440) );
  OR U33708 ( .A(n33177), .B(n33176), .Z(n33181) );
  NAND U33709 ( .A(n33179), .B(n33178), .Z(n33180) );
  NAND U33710 ( .A(n33181), .B(n33180), .Z(n33379) );
  OR U33711 ( .A(n33183), .B(n33182), .Z(n33187) );
  NANDN U33712 ( .A(n33185), .B(n33184), .Z(n33186) );
  NAND U33713 ( .A(n33187), .B(n33186), .Z(n33378) );
  OR U33714 ( .A(n33189), .B(n33188), .Z(n33193) );
  NANDN U33715 ( .A(n33191), .B(n33190), .Z(n33192) );
  NAND U33716 ( .A(n33193), .B(n33192), .Z(n33377) );
  XOR U33717 ( .A(n33379), .B(n33380), .Z(n33438) );
  OR U33718 ( .A(n33195), .B(n33194), .Z(n33199) );
  NANDN U33719 ( .A(n33197), .B(n33196), .Z(n33198) );
  NAND U33720 ( .A(n33199), .B(n33198), .Z(n33391) );
  XNOR U33721 ( .A(b[19]), .B(a[219]), .Z(n33335) );
  NANDN U33722 ( .A(n33335), .B(n37934), .Z(n33202) );
  NANDN U33723 ( .A(n33200), .B(n37935), .Z(n33201) );
  NAND U33724 ( .A(n33202), .B(n33201), .Z(n33404) );
  XOR U33725 ( .A(b[27]), .B(a[211]), .Z(n33338) );
  NAND U33726 ( .A(n38423), .B(n33338), .Z(n33205) );
  NAND U33727 ( .A(n33203), .B(n38424), .Z(n33204) );
  NAND U33728 ( .A(n33205), .B(n33204), .Z(n33401) );
  XOR U33729 ( .A(a[233]), .B(n1051), .Z(n33341) );
  NANDN U33730 ( .A(n33341), .B(n36587), .Z(n33208) );
  NANDN U33731 ( .A(n33206), .B(n36588), .Z(n33207) );
  AND U33732 ( .A(n33208), .B(n33207), .Z(n33402) );
  XNOR U33733 ( .A(n33401), .B(n33402), .Z(n33403) );
  XNOR U33734 ( .A(n33404), .B(n33403), .Z(n33390) );
  NAND U33735 ( .A(n33209), .B(n37762), .Z(n33211) );
  XOR U33736 ( .A(b[17]), .B(a[221]), .Z(n33344) );
  NAND U33737 ( .A(n33344), .B(n37764), .Z(n33210) );
  NAND U33738 ( .A(n33211), .B(n33210), .Z(n33362) );
  XNOR U33739 ( .A(b[31]), .B(a[207]), .Z(n33347) );
  NANDN U33740 ( .A(n33347), .B(n38552), .Z(n33214) );
  NANDN U33741 ( .A(n33212), .B(n38553), .Z(n33213) );
  NAND U33742 ( .A(n33214), .B(n33213), .Z(n33359) );
  OR U33743 ( .A(n33215), .B(n36105), .Z(n33217) );
  XOR U33744 ( .A(a[235]), .B(n1050), .Z(n33350) );
  NANDN U33745 ( .A(n33350), .B(n36107), .Z(n33216) );
  AND U33746 ( .A(n33217), .B(n33216), .Z(n33360) );
  XNOR U33747 ( .A(n33359), .B(n33360), .Z(n33361) );
  XOR U33748 ( .A(n33362), .B(n33361), .Z(n33389) );
  XOR U33749 ( .A(n33390), .B(n33389), .Z(n33392) );
  XOR U33750 ( .A(n33391), .B(n33392), .Z(n33437) );
  XOR U33751 ( .A(n33438), .B(n33437), .Z(n33439) );
  XNOR U33752 ( .A(n33440), .B(n33439), .Z(n33326) );
  OR U33753 ( .A(n33219), .B(n33218), .Z(n33223) );
  NAND U33754 ( .A(n33221), .B(n33220), .Z(n33222) );
  NAND U33755 ( .A(n33223), .B(n33222), .Z(n33324) );
  NANDN U33756 ( .A(n33225), .B(n33224), .Z(n33229) );
  NANDN U33757 ( .A(n33227), .B(n33226), .Z(n33228) );
  NAND U33758 ( .A(n33229), .B(n33228), .Z(n33445) );
  OR U33759 ( .A(n33231), .B(n33230), .Z(n33235) );
  NAND U33760 ( .A(n33233), .B(n33232), .Z(n33234) );
  NAND U33761 ( .A(n33235), .B(n33234), .Z(n33444) );
  NANDN U33762 ( .A(n33237), .B(n33236), .Z(n33241) );
  NAND U33763 ( .A(n33239), .B(n33238), .Z(n33240) );
  NAND U33764 ( .A(n33241), .B(n33240), .Z(n33383) );
  NANDN U33765 ( .A(n33243), .B(n33242), .Z(n33247) );
  NAND U33766 ( .A(n33245), .B(n33244), .Z(n33246) );
  AND U33767 ( .A(n33247), .B(n33246), .Z(n33384) );
  XNOR U33768 ( .A(n33383), .B(n33384), .Z(n33385) );
  XNOR U33769 ( .A(n1052), .B(a[229]), .Z(n33413) );
  NAND U33770 ( .A(n36925), .B(n33413), .Z(n33250) );
  NANDN U33771 ( .A(n33248), .B(n36926), .Z(n33249) );
  NAND U33772 ( .A(n33250), .B(n33249), .Z(n33367) );
  XNOR U33773 ( .A(b[15]), .B(a[223]), .Z(n33410) );
  OR U33774 ( .A(n33410), .B(n37665), .Z(n33253) );
  NANDN U33775 ( .A(n33251), .B(n37604), .Z(n33252) );
  AND U33776 ( .A(n33253), .B(n33252), .Z(n33365) );
  XOR U33777 ( .A(n1056), .B(n34670), .Z(n33407) );
  NAND U33778 ( .A(n33407), .B(n38101), .Z(n33256) );
  NANDN U33779 ( .A(n33254), .B(n38102), .Z(n33255) );
  AND U33780 ( .A(n33256), .B(n33255), .Z(n33366) );
  XOR U33781 ( .A(n33367), .B(n33368), .Z(n33356) );
  XNOR U33782 ( .A(b[11]), .B(a[227]), .Z(n33416) );
  OR U33783 ( .A(n33416), .B(n37311), .Z(n33259) );
  NANDN U33784 ( .A(n33257), .B(n37218), .Z(n33258) );
  NAND U33785 ( .A(n33259), .B(n33258), .Z(n33354) );
  XOR U33786 ( .A(n1053), .B(a[225]), .Z(n33419) );
  NANDN U33787 ( .A(n33419), .B(n37424), .Z(n33262) );
  NANDN U33788 ( .A(n33260), .B(n37425), .Z(n33261) );
  AND U33789 ( .A(n33262), .B(n33261), .Z(n33353) );
  XNOR U33790 ( .A(n33354), .B(n33353), .Z(n33355) );
  XOR U33791 ( .A(n33356), .B(n33355), .Z(n33373) );
  NANDN U33792 ( .A(n1049), .B(a[237]), .Z(n33263) );
  XNOR U33793 ( .A(b[1]), .B(n33263), .Z(n33265) );
  IV U33794 ( .A(a[236]), .Z(n37106) );
  NANDN U33795 ( .A(n37106), .B(n1049), .Z(n33264) );
  AND U33796 ( .A(n33265), .B(n33264), .Z(n33331) );
  NAND U33797 ( .A(n33266), .B(n38490), .Z(n33268) );
  XNOR U33798 ( .A(n1058), .B(a[209]), .Z(n33425) );
  NANDN U33799 ( .A(n1048), .B(n33425), .Z(n33267) );
  NAND U33800 ( .A(n33268), .B(n33267), .Z(n33329) );
  NANDN U33801 ( .A(n1059), .B(a[205]), .Z(n33330) );
  XNOR U33802 ( .A(n33329), .B(n33330), .Z(n33332) );
  XOR U33803 ( .A(n33331), .B(n33332), .Z(n33371) );
  NANDN U33804 ( .A(n33269), .B(n38205), .Z(n33271) );
  XOR U33805 ( .A(b[23]), .B(n34725), .Z(n33428) );
  OR U33806 ( .A(n33428), .B(n38268), .Z(n33270) );
  NAND U33807 ( .A(n33271), .B(n33270), .Z(n33398) );
  XNOR U33808 ( .A(b[7]), .B(a[231]), .Z(n33431) );
  NANDN U33809 ( .A(n33431), .B(n36701), .Z(n33274) );
  NANDN U33810 ( .A(n33272), .B(n36702), .Z(n33273) );
  NAND U33811 ( .A(n33274), .B(n33273), .Z(n33395) );
  XOR U33812 ( .A(b[25]), .B(a[213]), .Z(n33434) );
  NAND U33813 ( .A(n33434), .B(n38325), .Z(n33277) );
  NAND U33814 ( .A(n33275), .B(n38326), .Z(n33276) );
  AND U33815 ( .A(n33277), .B(n33276), .Z(n33396) );
  XNOR U33816 ( .A(n33395), .B(n33396), .Z(n33397) );
  XNOR U33817 ( .A(n33398), .B(n33397), .Z(n33372) );
  XOR U33818 ( .A(n33371), .B(n33372), .Z(n33374) );
  XNOR U33819 ( .A(n33373), .B(n33374), .Z(n33386) );
  XNOR U33820 ( .A(n33385), .B(n33386), .Z(n33443) );
  XNOR U33821 ( .A(n33444), .B(n33443), .Z(n33446) );
  XNOR U33822 ( .A(n33445), .B(n33446), .Z(n33323) );
  XNOR U33823 ( .A(n33324), .B(n33323), .Z(n33325) );
  XOR U33824 ( .A(n33326), .B(n33325), .Z(n33320) );
  NANDN U33825 ( .A(n33279), .B(n33278), .Z(n33283) );
  OR U33826 ( .A(n33281), .B(n33280), .Z(n33282) );
  NAND U33827 ( .A(n33283), .B(n33282), .Z(n33317) );
  NAND U33828 ( .A(n33285), .B(n33284), .Z(n33289) );
  NANDN U33829 ( .A(n33287), .B(n33286), .Z(n33288) );
  NAND U33830 ( .A(n33289), .B(n33288), .Z(n33318) );
  XNOR U33831 ( .A(n33317), .B(n33318), .Z(n33319) );
  XNOR U33832 ( .A(n33320), .B(n33319), .Z(n33314) );
  NANDN U33833 ( .A(n33291), .B(n33290), .Z(n33295) );
  NAND U33834 ( .A(n33293), .B(n33292), .Z(n33294) );
  NAND U33835 ( .A(n33295), .B(n33294), .Z(n33311) );
  NANDN U33836 ( .A(n33297), .B(n33296), .Z(n33301) );
  OR U33837 ( .A(n33299), .B(n33298), .Z(n33300) );
  NAND U33838 ( .A(n33301), .B(n33300), .Z(n33312) );
  XNOR U33839 ( .A(n33311), .B(n33312), .Z(n33313) );
  XNOR U33840 ( .A(n33314), .B(n33313), .Z(n33307) );
  XOR U33841 ( .A(n33308), .B(n33307), .Z(n33309) );
  XNOR U33842 ( .A(n33310), .B(n33309), .Z(n33449) );
  XNOR U33843 ( .A(n33449), .B(sreg[461]), .Z(n33451) );
  NAND U33844 ( .A(n33302), .B(sreg[460]), .Z(n33306) );
  OR U33845 ( .A(n33304), .B(n33303), .Z(n33305) );
  AND U33846 ( .A(n33306), .B(n33305), .Z(n33450) );
  XOR U33847 ( .A(n33451), .B(n33450), .Z(c[461]) );
  NANDN U33848 ( .A(n33312), .B(n33311), .Z(n33316) );
  NANDN U33849 ( .A(n33314), .B(n33313), .Z(n33315) );
  NAND U33850 ( .A(n33316), .B(n33315), .Z(n33455) );
  NANDN U33851 ( .A(n33318), .B(n33317), .Z(n33322) );
  NAND U33852 ( .A(n33320), .B(n33319), .Z(n33321) );
  NAND U33853 ( .A(n33322), .B(n33321), .Z(n33460) );
  NANDN U33854 ( .A(n33324), .B(n33323), .Z(n33328) );
  NANDN U33855 ( .A(n33326), .B(n33325), .Z(n33327) );
  NAND U33856 ( .A(n33328), .B(n33327), .Z(n33461) );
  XNOR U33857 ( .A(n33460), .B(n33461), .Z(n33462) );
  NANDN U33858 ( .A(n33330), .B(n33329), .Z(n33334) );
  NAND U33859 ( .A(n33332), .B(n33331), .Z(n33333) );
  NAND U33860 ( .A(n33334), .B(n33333), .Z(n33527) );
  XNOR U33861 ( .A(b[19]), .B(a[220]), .Z(n33472) );
  NANDN U33862 ( .A(n33472), .B(n37934), .Z(n33337) );
  NANDN U33863 ( .A(n33335), .B(n37935), .Z(n33336) );
  NAND U33864 ( .A(n33337), .B(n33336), .Z(n33537) );
  XOR U33865 ( .A(b[27]), .B(a[212]), .Z(n33475) );
  NAND U33866 ( .A(n38423), .B(n33475), .Z(n33340) );
  NAND U33867 ( .A(n33338), .B(n38424), .Z(n33339) );
  NAND U33868 ( .A(n33340), .B(n33339), .Z(n33534) );
  XOR U33869 ( .A(a[234]), .B(n1051), .Z(n33478) );
  NANDN U33870 ( .A(n33478), .B(n36587), .Z(n33343) );
  NANDN U33871 ( .A(n33341), .B(n36588), .Z(n33342) );
  AND U33872 ( .A(n33343), .B(n33342), .Z(n33535) );
  XNOR U33873 ( .A(n33534), .B(n33535), .Z(n33536) );
  XNOR U33874 ( .A(n33537), .B(n33536), .Z(n33525) );
  NAND U33875 ( .A(n33344), .B(n37762), .Z(n33346) );
  XNOR U33876 ( .A(b[17]), .B(a[222]), .Z(n33481) );
  NANDN U33877 ( .A(n33481), .B(n37764), .Z(n33345) );
  NAND U33878 ( .A(n33346), .B(n33345), .Z(n33499) );
  XNOR U33879 ( .A(b[31]), .B(a[208]), .Z(n33484) );
  NANDN U33880 ( .A(n33484), .B(n38552), .Z(n33349) );
  NANDN U33881 ( .A(n33347), .B(n38553), .Z(n33348) );
  NAND U33882 ( .A(n33349), .B(n33348), .Z(n33496) );
  OR U33883 ( .A(n33350), .B(n36105), .Z(n33352) );
  XOR U33884 ( .A(a[236]), .B(n1050), .Z(n33487) );
  NANDN U33885 ( .A(n33487), .B(n36107), .Z(n33351) );
  AND U33886 ( .A(n33352), .B(n33351), .Z(n33497) );
  XNOR U33887 ( .A(n33496), .B(n33497), .Z(n33498) );
  XOR U33888 ( .A(n33499), .B(n33498), .Z(n33524) );
  XNOR U33889 ( .A(n33525), .B(n33524), .Z(n33526) );
  XNOR U33890 ( .A(n33527), .B(n33526), .Z(n33570) );
  NANDN U33891 ( .A(n33354), .B(n33353), .Z(n33358) );
  NAND U33892 ( .A(n33356), .B(n33355), .Z(n33357) );
  NAND U33893 ( .A(n33358), .B(n33357), .Z(n33515) );
  NANDN U33894 ( .A(n33360), .B(n33359), .Z(n33364) );
  NAND U33895 ( .A(n33362), .B(n33361), .Z(n33363) );
  NAND U33896 ( .A(n33364), .B(n33363), .Z(n33513) );
  OR U33897 ( .A(n33366), .B(n33365), .Z(n33370) );
  NANDN U33898 ( .A(n33368), .B(n33367), .Z(n33369) );
  NAND U33899 ( .A(n33370), .B(n33369), .Z(n33512) );
  XNOR U33900 ( .A(n33515), .B(n33514), .Z(n33571) );
  XOR U33901 ( .A(n33570), .B(n33571), .Z(n33573) );
  NANDN U33902 ( .A(n33372), .B(n33371), .Z(n33376) );
  OR U33903 ( .A(n33374), .B(n33373), .Z(n33375) );
  NAND U33904 ( .A(n33376), .B(n33375), .Z(n33572) );
  XOR U33905 ( .A(n33573), .B(n33572), .Z(n33590) );
  OR U33906 ( .A(n33378), .B(n33377), .Z(n33382) );
  NANDN U33907 ( .A(n33380), .B(n33379), .Z(n33381) );
  NAND U33908 ( .A(n33382), .B(n33381), .Z(n33589) );
  NANDN U33909 ( .A(n33384), .B(n33383), .Z(n33388) );
  NANDN U33910 ( .A(n33386), .B(n33385), .Z(n33387) );
  NAND U33911 ( .A(n33388), .B(n33387), .Z(n33578) );
  NANDN U33912 ( .A(n33390), .B(n33389), .Z(n33394) );
  OR U33913 ( .A(n33392), .B(n33391), .Z(n33393) );
  NAND U33914 ( .A(n33394), .B(n33393), .Z(n33577) );
  NANDN U33915 ( .A(n33396), .B(n33395), .Z(n33400) );
  NAND U33916 ( .A(n33398), .B(n33397), .Z(n33399) );
  NAND U33917 ( .A(n33400), .B(n33399), .Z(n33518) );
  NANDN U33918 ( .A(n33402), .B(n33401), .Z(n33406) );
  NAND U33919 ( .A(n33404), .B(n33403), .Z(n33405) );
  AND U33920 ( .A(n33406), .B(n33405), .Z(n33519) );
  XNOR U33921 ( .A(n33518), .B(n33519), .Z(n33520) );
  XOR U33922 ( .A(n1056), .B(a[218]), .Z(n33546) );
  NANDN U33923 ( .A(n33546), .B(n38101), .Z(n33409) );
  NAND U33924 ( .A(n38102), .B(n33407), .Z(n33408) );
  NAND U33925 ( .A(n33409), .B(n33408), .Z(n33508) );
  XNOR U33926 ( .A(b[15]), .B(a[224]), .Z(n33543) );
  OR U33927 ( .A(n33543), .B(n37665), .Z(n33412) );
  NANDN U33928 ( .A(n33410), .B(n37604), .Z(n33411) );
  AND U33929 ( .A(n33412), .B(n33411), .Z(n33509) );
  XNOR U33930 ( .A(n33508), .B(n33509), .Z(n33511) );
  XOR U33931 ( .A(n1052), .B(a[230]), .Z(n33540) );
  NANDN U33932 ( .A(n33540), .B(n36925), .Z(n33415) );
  NAND U33933 ( .A(n36926), .B(n33413), .Z(n33414) );
  NAND U33934 ( .A(n33415), .B(n33414), .Z(n33510) );
  XNOR U33935 ( .A(n33511), .B(n33510), .Z(n33504) );
  XOR U33936 ( .A(b[11]), .B(n36592), .Z(n33549) );
  OR U33937 ( .A(n33549), .B(n37311), .Z(n33418) );
  NANDN U33938 ( .A(n33416), .B(n37218), .Z(n33417) );
  NAND U33939 ( .A(n33418), .B(n33417), .Z(n33503) );
  XOR U33940 ( .A(n1053), .B(a[226]), .Z(n33552) );
  NANDN U33941 ( .A(n33552), .B(n37424), .Z(n33421) );
  NANDN U33942 ( .A(n33419), .B(n37425), .Z(n33420) );
  NAND U33943 ( .A(n33421), .B(n33420), .Z(n33502) );
  XNOR U33944 ( .A(n33503), .B(n33502), .Z(n33505) );
  XNOR U33945 ( .A(n33504), .B(n33505), .Z(n33493) );
  NANDN U33946 ( .A(n1049), .B(a[238]), .Z(n33422) );
  XNOR U33947 ( .A(b[1]), .B(n33422), .Z(n33424) );
  NANDN U33948 ( .A(b[0]), .B(a[237]), .Z(n33423) );
  AND U33949 ( .A(n33424), .B(n33423), .Z(n33468) );
  NAND U33950 ( .A(n38490), .B(n33425), .Z(n33427) );
  XNOR U33951 ( .A(n1058), .B(a[210]), .Z(n33555) );
  NANDN U33952 ( .A(n1048), .B(n33555), .Z(n33426) );
  NAND U33953 ( .A(n33427), .B(n33426), .Z(n33466) );
  NANDN U33954 ( .A(n1059), .B(a[206]), .Z(n33467) );
  XNOR U33955 ( .A(n33466), .B(n33467), .Z(n33469) );
  XNOR U33956 ( .A(n33468), .B(n33469), .Z(n33491) );
  NANDN U33957 ( .A(n33428), .B(n38205), .Z(n33430) );
  XNOR U33958 ( .A(b[23]), .B(a[216]), .Z(n33561) );
  OR U33959 ( .A(n33561), .B(n38268), .Z(n33429) );
  NAND U33960 ( .A(n33430), .B(n33429), .Z(n33531) );
  XNOR U33961 ( .A(a[232]), .B(b[7]), .Z(n33564) );
  NANDN U33962 ( .A(n33564), .B(n36701), .Z(n33433) );
  NANDN U33963 ( .A(n33431), .B(n36702), .Z(n33432) );
  NAND U33964 ( .A(n33433), .B(n33432), .Z(n33528) );
  XOR U33965 ( .A(b[25]), .B(a[214]), .Z(n33567) );
  NAND U33966 ( .A(n33567), .B(n38325), .Z(n33436) );
  NAND U33967 ( .A(n33434), .B(n38326), .Z(n33435) );
  AND U33968 ( .A(n33436), .B(n33435), .Z(n33529) );
  XNOR U33969 ( .A(n33528), .B(n33529), .Z(n33530) );
  XOR U33970 ( .A(n33531), .B(n33530), .Z(n33490) );
  XOR U33971 ( .A(n33493), .B(n33492), .Z(n33521) );
  XNOR U33972 ( .A(n33520), .B(n33521), .Z(n33576) );
  XNOR U33973 ( .A(n33577), .B(n33576), .Z(n33579) );
  XNOR U33974 ( .A(n33578), .B(n33579), .Z(n33588) );
  XOR U33975 ( .A(n33589), .B(n33588), .Z(n33591) );
  NAND U33976 ( .A(n33438), .B(n33437), .Z(n33442) );
  NAND U33977 ( .A(n33440), .B(n33439), .Z(n33441) );
  NAND U33978 ( .A(n33442), .B(n33441), .Z(n33583) );
  NAND U33979 ( .A(n33444), .B(n33443), .Z(n33448) );
  NANDN U33980 ( .A(n33446), .B(n33445), .Z(n33447) );
  AND U33981 ( .A(n33448), .B(n33447), .Z(n33582) );
  XNOR U33982 ( .A(n33583), .B(n33582), .Z(n33584) );
  XOR U33983 ( .A(n33585), .B(n33584), .Z(n33463) );
  XOR U33984 ( .A(n33462), .B(n33463), .Z(n33454) );
  XOR U33985 ( .A(n33455), .B(n33454), .Z(n33456) );
  XNOR U33986 ( .A(n33457), .B(n33456), .Z(n33594) );
  XNOR U33987 ( .A(n33594), .B(sreg[462]), .Z(n33596) );
  NAND U33988 ( .A(n33449), .B(sreg[461]), .Z(n33453) );
  OR U33989 ( .A(n33451), .B(n33450), .Z(n33452) );
  AND U33990 ( .A(n33453), .B(n33452), .Z(n33595) );
  XOR U33991 ( .A(n33596), .B(n33595), .Z(c[462]) );
  NAND U33992 ( .A(n33455), .B(n33454), .Z(n33459) );
  NAND U33993 ( .A(n33457), .B(n33456), .Z(n33458) );
  NAND U33994 ( .A(n33459), .B(n33458), .Z(n33602) );
  NANDN U33995 ( .A(n33461), .B(n33460), .Z(n33465) );
  NAND U33996 ( .A(n33463), .B(n33462), .Z(n33464) );
  NAND U33997 ( .A(n33465), .B(n33464), .Z(n33600) );
  NANDN U33998 ( .A(n33467), .B(n33466), .Z(n33471) );
  NAND U33999 ( .A(n33469), .B(n33468), .Z(n33470) );
  NAND U34000 ( .A(n33471), .B(n33470), .Z(n33670) );
  XNOR U34001 ( .A(b[19]), .B(a[221]), .Z(n33617) );
  NANDN U34002 ( .A(n33617), .B(n37934), .Z(n33474) );
  NANDN U34003 ( .A(n33472), .B(n37935), .Z(n33473) );
  NAND U34004 ( .A(n33474), .B(n33473), .Z(n33680) );
  XOR U34005 ( .A(b[27]), .B(a[213]), .Z(n33620) );
  NAND U34006 ( .A(n38423), .B(n33620), .Z(n33477) );
  NAND U34007 ( .A(n33475), .B(n38424), .Z(n33476) );
  NAND U34008 ( .A(n33477), .B(n33476), .Z(n33677) );
  XOR U34009 ( .A(a[235]), .B(n1051), .Z(n33623) );
  NANDN U34010 ( .A(n33623), .B(n36587), .Z(n33480) );
  NANDN U34011 ( .A(n33478), .B(n36588), .Z(n33479) );
  AND U34012 ( .A(n33480), .B(n33479), .Z(n33678) );
  XNOR U34013 ( .A(n33677), .B(n33678), .Z(n33679) );
  XNOR U34014 ( .A(n33680), .B(n33679), .Z(n33668) );
  NANDN U34015 ( .A(n33481), .B(n37762), .Z(n33483) );
  XOR U34016 ( .A(b[17]), .B(a[223]), .Z(n33626) );
  NAND U34017 ( .A(n33626), .B(n37764), .Z(n33482) );
  NAND U34018 ( .A(n33483), .B(n33482), .Z(n33644) );
  XNOR U34019 ( .A(b[31]), .B(a[209]), .Z(n33629) );
  NANDN U34020 ( .A(n33629), .B(n38552), .Z(n33486) );
  NANDN U34021 ( .A(n33484), .B(n38553), .Z(n33485) );
  NAND U34022 ( .A(n33486), .B(n33485), .Z(n33641) );
  OR U34023 ( .A(n33487), .B(n36105), .Z(n33489) );
  XNOR U34024 ( .A(a[237]), .B(b[3]), .Z(n33632) );
  NANDN U34025 ( .A(n33632), .B(n36107), .Z(n33488) );
  AND U34026 ( .A(n33489), .B(n33488), .Z(n33642) );
  XNOR U34027 ( .A(n33641), .B(n33642), .Z(n33643) );
  XOR U34028 ( .A(n33644), .B(n33643), .Z(n33667) );
  XNOR U34029 ( .A(n33668), .B(n33667), .Z(n33669) );
  XNOR U34030 ( .A(n33670), .B(n33669), .Z(n33719) );
  NANDN U34031 ( .A(n33491), .B(n33490), .Z(n33495) );
  NANDN U34032 ( .A(n33493), .B(n33492), .Z(n33494) );
  NAND U34033 ( .A(n33495), .B(n33494), .Z(n33720) );
  XNOR U34034 ( .A(n33719), .B(n33720), .Z(n33721) );
  NANDN U34035 ( .A(n33497), .B(n33496), .Z(n33501) );
  NAND U34036 ( .A(n33499), .B(n33498), .Z(n33500) );
  NAND U34037 ( .A(n33501), .B(n33500), .Z(n33660) );
  OR U34038 ( .A(n33503), .B(n33502), .Z(n33507) );
  NANDN U34039 ( .A(n33505), .B(n33504), .Z(n33506) );
  NAND U34040 ( .A(n33507), .B(n33506), .Z(n33658) );
  XNOR U34041 ( .A(n33658), .B(n33657), .Z(n33659) );
  XOR U34042 ( .A(n33660), .B(n33659), .Z(n33722) );
  XOR U34043 ( .A(n33721), .B(n33722), .Z(n33732) );
  OR U34044 ( .A(n33513), .B(n33512), .Z(n33517) );
  NAND U34045 ( .A(n33515), .B(n33514), .Z(n33516) );
  NAND U34046 ( .A(n33517), .B(n33516), .Z(n33730) );
  NANDN U34047 ( .A(n33519), .B(n33518), .Z(n33523) );
  NANDN U34048 ( .A(n33521), .B(n33520), .Z(n33522) );
  NAND U34049 ( .A(n33523), .B(n33522), .Z(n33715) );
  NANDN U34050 ( .A(n33529), .B(n33528), .Z(n33533) );
  NAND U34051 ( .A(n33531), .B(n33530), .Z(n33532) );
  NAND U34052 ( .A(n33533), .B(n33532), .Z(n33661) );
  NANDN U34053 ( .A(n33535), .B(n33534), .Z(n33539) );
  NAND U34054 ( .A(n33537), .B(n33536), .Z(n33538) );
  AND U34055 ( .A(n33539), .B(n33538), .Z(n33662) );
  XNOR U34056 ( .A(n33661), .B(n33662), .Z(n33663) );
  XOR U34057 ( .A(n1052), .B(a[231]), .Z(n33689) );
  NANDN U34058 ( .A(n33689), .B(n36925), .Z(n33542) );
  NANDN U34059 ( .A(n33540), .B(n36926), .Z(n33541) );
  NAND U34060 ( .A(n33542), .B(n33541), .Z(n33649) );
  XNOR U34061 ( .A(n1054), .B(a[225]), .Z(n33686) );
  NANDN U34062 ( .A(n37665), .B(n33686), .Z(n33545) );
  NANDN U34063 ( .A(n33543), .B(n37604), .Z(n33544) );
  NAND U34064 ( .A(n33545), .B(n33544), .Z(n33647) );
  XOR U34065 ( .A(n1056), .B(a[219]), .Z(n33683) );
  NANDN U34066 ( .A(n33683), .B(n38101), .Z(n33548) );
  NANDN U34067 ( .A(n33546), .B(n38102), .Z(n33547) );
  NAND U34068 ( .A(n33548), .B(n33547), .Z(n33648) );
  XNOR U34069 ( .A(n33647), .B(n33648), .Z(n33650) );
  XOR U34070 ( .A(n33649), .B(n33650), .Z(n33638) );
  XNOR U34071 ( .A(b[11]), .B(a[229]), .Z(n33692) );
  OR U34072 ( .A(n33692), .B(n37311), .Z(n33551) );
  NANDN U34073 ( .A(n33549), .B(n37218), .Z(n33550) );
  NAND U34074 ( .A(n33551), .B(n33550), .Z(n33636) );
  XOR U34075 ( .A(n1053), .B(a[227]), .Z(n33695) );
  NANDN U34076 ( .A(n33695), .B(n37424), .Z(n33554) );
  NANDN U34077 ( .A(n33552), .B(n37425), .Z(n33553) );
  AND U34078 ( .A(n33554), .B(n33553), .Z(n33635) );
  XNOR U34079 ( .A(n33636), .B(n33635), .Z(n33637) );
  XNOR U34080 ( .A(n33638), .B(n33637), .Z(n33654) );
  NAND U34081 ( .A(n38490), .B(n33555), .Z(n33557) );
  XNOR U34082 ( .A(n1058), .B(a[211]), .Z(n33701) );
  NANDN U34083 ( .A(n1048), .B(n33701), .Z(n33556) );
  NAND U34084 ( .A(n33557), .B(n33556), .Z(n33611) );
  NANDN U34085 ( .A(n1059), .B(a[207]), .Z(n33612) );
  XNOR U34086 ( .A(n33611), .B(n33612), .Z(n33614) );
  NANDN U34087 ( .A(n1049), .B(a[239]), .Z(n33558) );
  XNOR U34088 ( .A(b[1]), .B(n33558), .Z(n33560) );
  IV U34089 ( .A(a[238]), .Z(n37467) );
  NANDN U34090 ( .A(n37467), .B(n1049), .Z(n33559) );
  AND U34091 ( .A(n33560), .B(n33559), .Z(n33613) );
  XNOR U34092 ( .A(n33614), .B(n33613), .Z(n33652) );
  NANDN U34093 ( .A(n33561), .B(n38205), .Z(n33563) );
  XOR U34094 ( .A(b[23]), .B(n34670), .Z(n33704) );
  OR U34095 ( .A(n33704), .B(n38268), .Z(n33562) );
  NAND U34096 ( .A(n33563), .B(n33562), .Z(n33674) );
  XNOR U34097 ( .A(b[7]), .B(a[233]), .Z(n33707) );
  NANDN U34098 ( .A(n33707), .B(n36701), .Z(n33566) );
  NANDN U34099 ( .A(n33564), .B(n36702), .Z(n33565) );
  NAND U34100 ( .A(n33566), .B(n33565), .Z(n33671) );
  XNOR U34101 ( .A(b[25]), .B(a[215]), .Z(n33710) );
  NANDN U34102 ( .A(n33710), .B(n38325), .Z(n33569) );
  NAND U34103 ( .A(n33567), .B(n38326), .Z(n33568) );
  AND U34104 ( .A(n33569), .B(n33568), .Z(n33672) );
  XNOR U34105 ( .A(n33671), .B(n33672), .Z(n33673) );
  XOR U34106 ( .A(n33674), .B(n33673), .Z(n33651) );
  XOR U34107 ( .A(n33654), .B(n33653), .Z(n33664) );
  XOR U34108 ( .A(n33663), .B(n33664), .Z(n33713) );
  XNOR U34109 ( .A(n33714), .B(n33713), .Z(n33716) );
  XNOR U34110 ( .A(n33715), .B(n33716), .Z(n33729) );
  XOR U34111 ( .A(n33730), .B(n33729), .Z(n33731) );
  XNOR U34112 ( .A(n33732), .B(n33731), .Z(n33726) );
  NANDN U34113 ( .A(n33571), .B(n33570), .Z(n33575) );
  OR U34114 ( .A(n33573), .B(n33572), .Z(n33574) );
  NAND U34115 ( .A(n33575), .B(n33574), .Z(n33723) );
  NAND U34116 ( .A(n33577), .B(n33576), .Z(n33581) );
  NANDN U34117 ( .A(n33579), .B(n33578), .Z(n33580) );
  NAND U34118 ( .A(n33581), .B(n33580), .Z(n33724) );
  XNOR U34119 ( .A(n33723), .B(n33724), .Z(n33725) );
  XOR U34120 ( .A(n33726), .B(n33725), .Z(n33607) );
  NANDN U34121 ( .A(n33583), .B(n33582), .Z(n33587) );
  NAND U34122 ( .A(n33585), .B(n33584), .Z(n33586) );
  NAND U34123 ( .A(n33587), .B(n33586), .Z(n33605) );
  NANDN U34124 ( .A(n33589), .B(n33588), .Z(n33593) );
  OR U34125 ( .A(n33591), .B(n33590), .Z(n33592) );
  NAND U34126 ( .A(n33593), .B(n33592), .Z(n33606) );
  XNOR U34127 ( .A(n33605), .B(n33606), .Z(n33608) );
  XOR U34128 ( .A(n33607), .B(n33608), .Z(n33599) );
  XOR U34129 ( .A(n33600), .B(n33599), .Z(n33601) );
  XNOR U34130 ( .A(n33602), .B(n33601), .Z(n33735) );
  XNOR U34131 ( .A(n33735), .B(sreg[463]), .Z(n33737) );
  NAND U34132 ( .A(n33594), .B(sreg[462]), .Z(n33598) );
  OR U34133 ( .A(n33596), .B(n33595), .Z(n33597) );
  AND U34134 ( .A(n33598), .B(n33597), .Z(n33736) );
  XOR U34135 ( .A(n33737), .B(n33736), .Z(c[463]) );
  NAND U34136 ( .A(n33600), .B(n33599), .Z(n33604) );
  NAND U34137 ( .A(n33602), .B(n33601), .Z(n33603) );
  NAND U34138 ( .A(n33604), .B(n33603), .Z(n33743) );
  NANDN U34139 ( .A(n33606), .B(n33605), .Z(n33610) );
  NAND U34140 ( .A(n33608), .B(n33607), .Z(n33609) );
  NAND U34141 ( .A(n33610), .B(n33609), .Z(n33741) );
  NANDN U34142 ( .A(n33612), .B(n33611), .Z(n33616) );
  NAND U34143 ( .A(n33614), .B(n33613), .Z(n33615) );
  NAND U34144 ( .A(n33616), .B(n33615), .Z(n33819) );
  XOR U34145 ( .A(b[19]), .B(n35381), .Z(n33766) );
  NANDN U34146 ( .A(n33766), .B(n37934), .Z(n33619) );
  NANDN U34147 ( .A(n33617), .B(n37935), .Z(n33618) );
  NAND U34148 ( .A(n33619), .B(n33618), .Z(n33829) );
  XOR U34149 ( .A(b[27]), .B(a[214]), .Z(n33769) );
  NAND U34150 ( .A(n38423), .B(n33769), .Z(n33622) );
  NAND U34151 ( .A(n33620), .B(n38424), .Z(n33621) );
  NAND U34152 ( .A(n33622), .B(n33621), .Z(n33826) );
  XOR U34153 ( .A(a[236]), .B(n1051), .Z(n33772) );
  NANDN U34154 ( .A(n33772), .B(n36587), .Z(n33625) );
  NANDN U34155 ( .A(n33623), .B(n36588), .Z(n33624) );
  AND U34156 ( .A(n33625), .B(n33624), .Z(n33827) );
  XNOR U34157 ( .A(n33826), .B(n33827), .Z(n33828) );
  XNOR U34158 ( .A(n33829), .B(n33828), .Z(n33817) );
  NAND U34159 ( .A(n33626), .B(n37762), .Z(n33628) );
  XOR U34160 ( .A(b[17]), .B(a[224]), .Z(n33775) );
  NAND U34161 ( .A(n33775), .B(n37764), .Z(n33627) );
  NAND U34162 ( .A(n33628), .B(n33627), .Z(n33793) );
  XNOR U34163 ( .A(b[31]), .B(a[210]), .Z(n33778) );
  NANDN U34164 ( .A(n33778), .B(n38552), .Z(n33631) );
  NANDN U34165 ( .A(n33629), .B(n38553), .Z(n33630) );
  NAND U34166 ( .A(n33631), .B(n33630), .Z(n33790) );
  OR U34167 ( .A(n33632), .B(n36105), .Z(n33634) );
  XOR U34168 ( .A(a[238]), .B(n1050), .Z(n33781) );
  NANDN U34169 ( .A(n33781), .B(n36107), .Z(n33633) );
  AND U34170 ( .A(n33634), .B(n33633), .Z(n33791) );
  XNOR U34171 ( .A(n33790), .B(n33791), .Z(n33792) );
  XOR U34172 ( .A(n33793), .B(n33792), .Z(n33816) );
  XNOR U34173 ( .A(n33817), .B(n33816), .Z(n33818) );
  XNOR U34174 ( .A(n33819), .B(n33818), .Z(n33757) );
  NANDN U34175 ( .A(n33636), .B(n33635), .Z(n33640) );
  NAND U34176 ( .A(n33638), .B(n33637), .Z(n33639) );
  NAND U34177 ( .A(n33640), .B(n33639), .Z(n33808) );
  NANDN U34178 ( .A(n33642), .B(n33641), .Z(n33646) );
  NAND U34179 ( .A(n33644), .B(n33643), .Z(n33645) );
  NAND U34180 ( .A(n33646), .B(n33645), .Z(n33807) );
  XNOR U34181 ( .A(n33807), .B(n33806), .Z(n33809) );
  XOR U34182 ( .A(n33808), .B(n33809), .Z(n33756) );
  XOR U34183 ( .A(n33757), .B(n33756), .Z(n33758) );
  NANDN U34184 ( .A(n33652), .B(n33651), .Z(n33656) );
  NAND U34185 ( .A(n33654), .B(n33653), .Z(n33655) );
  AND U34186 ( .A(n33656), .B(n33655), .Z(n33759) );
  XNOR U34187 ( .A(n33758), .B(n33759), .Z(n33865) );
  NANDN U34188 ( .A(n33662), .B(n33661), .Z(n33666) );
  NAND U34189 ( .A(n33664), .B(n33663), .Z(n33665) );
  NAND U34190 ( .A(n33666), .B(n33665), .Z(n33753) );
  NANDN U34191 ( .A(n33672), .B(n33671), .Z(n33676) );
  NAND U34192 ( .A(n33674), .B(n33673), .Z(n33675) );
  NAND U34193 ( .A(n33676), .B(n33675), .Z(n33810) );
  NANDN U34194 ( .A(n33678), .B(n33677), .Z(n33682) );
  NAND U34195 ( .A(n33680), .B(n33679), .Z(n33681) );
  AND U34196 ( .A(n33682), .B(n33681), .Z(n33811) );
  XNOR U34197 ( .A(n33810), .B(n33811), .Z(n33812) );
  XNOR U34198 ( .A(b[21]), .B(a[220]), .Z(n33838) );
  NANDN U34199 ( .A(n33838), .B(n38101), .Z(n33685) );
  NANDN U34200 ( .A(n33683), .B(n38102), .Z(n33684) );
  NAND U34201 ( .A(n33685), .B(n33684), .Z(n33802) );
  XOR U34202 ( .A(b[15]), .B(n36280), .Z(n33835) );
  OR U34203 ( .A(n33835), .B(n37665), .Z(n33688) );
  NAND U34204 ( .A(n33686), .B(n37604), .Z(n33687) );
  AND U34205 ( .A(n33688), .B(n33687), .Z(n33803) );
  XNOR U34206 ( .A(n33802), .B(n33803), .Z(n33805) );
  XOR U34207 ( .A(b[9]), .B(n37079), .Z(n33832) );
  NANDN U34208 ( .A(n33832), .B(n36925), .Z(n33691) );
  NANDN U34209 ( .A(n33689), .B(n36926), .Z(n33690) );
  NAND U34210 ( .A(n33691), .B(n33690), .Z(n33804) );
  XNOR U34211 ( .A(n33805), .B(n33804), .Z(n33798) );
  XOR U34212 ( .A(b[11]), .B(n36333), .Z(n33841) );
  OR U34213 ( .A(n33841), .B(n37311), .Z(n33694) );
  NANDN U34214 ( .A(n33692), .B(n37218), .Z(n33693) );
  NAND U34215 ( .A(n33694), .B(n33693), .Z(n33797) );
  XOR U34216 ( .A(n1053), .B(a[228]), .Z(n33844) );
  NANDN U34217 ( .A(n33844), .B(n37424), .Z(n33697) );
  NANDN U34218 ( .A(n33695), .B(n37425), .Z(n33696) );
  NAND U34219 ( .A(n33697), .B(n33696), .Z(n33796) );
  XNOR U34220 ( .A(n33797), .B(n33796), .Z(n33799) );
  XNOR U34221 ( .A(n33798), .B(n33799), .Z(n33787) );
  NANDN U34222 ( .A(n1049), .B(a[240]), .Z(n33698) );
  XNOR U34223 ( .A(b[1]), .B(n33698), .Z(n33700) );
  NANDN U34224 ( .A(b[0]), .B(a[239]), .Z(n33699) );
  AND U34225 ( .A(n33700), .B(n33699), .Z(n33762) );
  NAND U34226 ( .A(n38490), .B(n33701), .Z(n33703) );
  XNOR U34227 ( .A(n1058), .B(a[212]), .Z(n33847) );
  NANDN U34228 ( .A(n1048), .B(n33847), .Z(n33702) );
  NAND U34229 ( .A(n33703), .B(n33702), .Z(n33760) );
  NANDN U34230 ( .A(n1059), .B(a[208]), .Z(n33761) );
  XNOR U34231 ( .A(n33760), .B(n33761), .Z(n33763) );
  XNOR U34232 ( .A(n33762), .B(n33763), .Z(n33785) );
  NANDN U34233 ( .A(n33704), .B(n38205), .Z(n33706) );
  XNOR U34234 ( .A(b[23]), .B(a[218]), .Z(n33853) );
  OR U34235 ( .A(n33853), .B(n38268), .Z(n33705) );
  NAND U34236 ( .A(n33706), .B(n33705), .Z(n33823) );
  XNOR U34237 ( .A(a[234]), .B(b[7]), .Z(n33856) );
  NANDN U34238 ( .A(n33856), .B(n36701), .Z(n33709) );
  NANDN U34239 ( .A(n33707), .B(n36702), .Z(n33708) );
  NAND U34240 ( .A(n33709), .B(n33708), .Z(n33820) );
  XOR U34241 ( .A(b[25]), .B(a[216]), .Z(n33859) );
  NAND U34242 ( .A(n33859), .B(n38325), .Z(n33712) );
  NANDN U34243 ( .A(n33710), .B(n38326), .Z(n33711) );
  AND U34244 ( .A(n33712), .B(n33711), .Z(n33821) );
  XNOR U34245 ( .A(n33820), .B(n33821), .Z(n33822) );
  XOR U34246 ( .A(n33823), .B(n33822), .Z(n33784) );
  XOR U34247 ( .A(n33787), .B(n33786), .Z(n33813) );
  XNOR U34248 ( .A(n33812), .B(n33813), .Z(n33750) );
  XOR U34249 ( .A(n33751), .B(n33750), .Z(n33752) );
  XOR U34250 ( .A(n33753), .B(n33752), .Z(n33863) );
  XNOR U34251 ( .A(n33862), .B(n33863), .Z(n33864) );
  XNOR U34252 ( .A(n33865), .B(n33864), .Z(n33869) );
  NAND U34253 ( .A(n33714), .B(n33713), .Z(n33718) );
  NANDN U34254 ( .A(n33716), .B(n33715), .Z(n33717) );
  NAND U34255 ( .A(n33718), .B(n33717), .Z(n33866) );
  XNOR U34256 ( .A(n33866), .B(n33867), .Z(n33868) );
  XNOR U34257 ( .A(n33869), .B(n33868), .Z(n33747) );
  NANDN U34258 ( .A(n33724), .B(n33723), .Z(n33728) );
  NAND U34259 ( .A(n33726), .B(n33725), .Z(n33727) );
  NAND U34260 ( .A(n33728), .B(n33727), .Z(n33744) );
  NANDN U34261 ( .A(n33730), .B(n33729), .Z(n33734) );
  OR U34262 ( .A(n33732), .B(n33731), .Z(n33733) );
  NAND U34263 ( .A(n33734), .B(n33733), .Z(n33745) );
  XNOR U34264 ( .A(n33744), .B(n33745), .Z(n33746) );
  XNOR U34265 ( .A(n33747), .B(n33746), .Z(n33740) );
  XOR U34266 ( .A(n33741), .B(n33740), .Z(n33742) );
  XNOR U34267 ( .A(n33743), .B(n33742), .Z(n33872) );
  XNOR U34268 ( .A(n33872), .B(sreg[464]), .Z(n33874) );
  NAND U34269 ( .A(n33735), .B(sreg[463]), .Z(n33739) );
  OR U34270 ( .A(n33737), .B(n33736), .Z(n33738) );
  AND U34271 ( .A(n33739), .B(n33738), .Z(n33873) );
  XOR U34272 ( .A(n33874), .B(n33873), .Z(c[464]) );
  NANDN U34273 ( .A(n33745), .B(n33744), .Z(n33749) );
  NANDN U34274 ( .A(n33747), .B(n33746), .Z(n33748) );
  NAND U34275 ( .A(n33749), .B(n33748), .Z(n33877) );
  NAND U34276 ( .A(n33751), .B(n33750), .Z(n33755) );
  NAND U34277 ( .A(n33753), .B(n33752), .Z(n33754) );
  NAND U34278 ( .A(n33755), .B(n33754), .Z(n34005) );
  XNOR U34279 ( .A(n34005), .B(n34006), .Z(n34007) );
  NANDN U34280 ( .A(n33761), .B(n33760), .Z(n33765) );
  NAND U34281 ( .A(n33763), .B(n33762), .Z(n33764) );
  NAND U34282 ( .A(n33765), .B(n33764), .Z(n33950) );
  XNOR U34283 ( .A(b[19]), .B(a[223]), .Z(n33895) );
  NANDN U34284 ( .A(n33895), .B(n37934), .Z(n33768) );
  NANDN U34285 ( .A(n33766), .B(n37935), .Z(n33767) );
  NAND U34286 ( .A(n33768), .B(n33767), .Z(n33960) );
  XNOR U34287 ( .A(b[27]), .B(a[215]), .Z(n33898) );
  NANDN U34288 ( .A(n33898), .B(n38423), .Z(n33771) );
  NAND U34289 ( .A(n33769), .B(n38424), .Z(n33770) );
  NAND U34290 ( .A(n33771), .B(n33770), .Z(n33957) );
  XNOR U34291 ( .A(a[237]), .B(b[5]), .Z(n33901) );
  NANDN U34292 ( .A(n33901), .B(n36587), .Z(n33774) );
  NANDN U34293 ( .A(n33772), .B(n36588), .Z(n33773) );
  AND U34294 ( .A(n33774), .B(n33773), .Z(n33958) );
  XNOR U34295 ( .A(n33957), .B(n33958), .Z(n33959) );
  XNOR U34296 ( .A(n33960), .B(n33959), .Z(n33948) );
  NAND U34297 ( .A(n33775), .B(n37762), .Z(n33777) );
  XNOR U34298 ( .A(b[17]), .B(a[225]), .Z(n33904) );
  NANDN U34299 ( .A(n33904), .B(n37764), .Z(n33776) );
  NAND U34300 ( .A(n33777), .B(n33776), .Z(n33922) );
  XNOR U34301 ( .A(b[31]), .B(a[211]), .Z(n33907) );
  NANDN U34302 ( .A(n33907), .B(n38552), .Z(n33780) );
  NANDN U34303 ( .A(n33778), .B(n38553), .Z(n33779) );
  NAND U34304 ( .A(n33780), .B(n33779), .Z(n33919) );
  OR U34305 ( .A(n33781), .B(n36105), .Z(n33783) );
  XNOR U34306 ( .A(a[239]), .B(b[3]), .Z(n33910) );
  NANDN U34307 ( .A(n33910), .B(n36107), .Z(n33782) );
  AND U34308 ( .A(n33783), .B(n33782), .Z(n33920) );
  XNOR U34309 ( .A(n33919), .B(n33920), .Z(n33921) );
  XOR U34310 ( .A(n33922), .B(n33921), .Z(n33947) );
  XNOR U34311 ( .A(n33948), .B(n33947), .Z(n33949) );
  XNOR U34312 ( .A(n33950), .B(n33949), .Z(n33999) );
  NANDN U34313 ( .A(n33785), .B(n33784), .Z(n33789) );
  NANDN U34314 ( .A(n33787), .B(n33786), .Z(n33788) );
  NAND U34315 ( .A(n33789), .B(n33788), .Z(n34000) );
  XNOR U34316 ( .A(n33999), .B(n34000), .Z(n34001) );
  NANDN U34317 ( .A(n33791), .B(n33790), .Z(n33795) );
  NAND U34318 ( .A(n33793), .B(n33792), .Z(n33794) );
  NAND U34319 ( .A(n33795), .B(n33794), .Z(n33940) );
  OR U34320 ( .A(n33797), .B(n33796), .Z(n33801) );
  NANDN U34321 ( .A(n33799), .B(n33798), .Z(n33800) );
  NAND U34322 ( .A(n33801), .B(n33800), .Z(n33938) );
  XNOR U34323 ( .A(n33938), .B(n33937), .Z(n33939) );
  XOR U34324 ( .A(n33940), .B(n33939), .Z(n34002) );
  XOR U34325 ( .A(n34001), .B(n34002), .Z(n34013) );
  NANDN U34326 ( .A(n33811), .B(n33810), .Z(n33815) );
  NANDN U34327 ( .A(n33813), .B(n33812), .Z(n33814) );
  NAND U34328 ( .A(n33815), .B(n33814), .Z(n33996) );
  NANDN U34329 ( .A(n33821), .B(n33820), .Z(n33825) );
  NAND U34330 ( .A(n33823), .B(n33822), .Z(n33824) );
  NAND U34331 ( .A(n33825), .B(n33824), .Z(n33941) );
  NANDN U34332 ( .A(n33827), .B(n33826), .Z(n33831) );
  NAND U34333 ( .A(n33829), .B(n33828), .Z(n33830) );
  AND U34334 ( .A(n33831), .B(n33830), .Z(n33942) );
  XNOR U34335 ( .A(n33941), .B(n33942), .Z(n33943) );
  XOR U34336 ( .A(b[9]), .B(n37184), .Z(n33963) );
  NANDN U34337 ( .A(n33963), .B(n36925), .Z(n33834) );
  NANDN U34338 ( .A(n33832), .B(n36926), .Z(n33833) );
  NAND U34339 ( .A(n33834), .B(n33833), .Z(n33927) );
  XNOR U34340 ( .A(b[15]), .B(a[227]), .Z(n33966) );
  OR U34341 ( .A(n33966), .B(n37665), .Z(n33837) );
  NANDN U34342 ( .A(n33835), .B(n37604), .Z(n33836) );
  AND U34343 ( .A(n33837), .B(n33836), .Z(n33925) );
  XNOR U34344 ( .A(b[21]), .B(a[221]), .Z(n33969) );
  NANDN U34345 ( .A(n33969), .B(n38101), .Z(n33840) );
  NANDN U34346 ( .A(n33838), .B(n38102), .Z(n33839) );
  AND U34347 ( .A(n33840), .B(n33839), .Z(n33926) );
  XOR U34348 ( .A(n33927), .B(n33928), .Z(n33916) );
  XOR U34349 ( .A(b[11]), .B(n36934), .Z(n33972) );
  OR U34350 ( .A(n33972), .B(n37311), .Z(n33843) );
  NANDN U34351 ( .A(n33841), .B(n37218), .Z(n33842) );
  NAND U34352 ( .A(n33843), .B(n33842), .Z(n33914) );
  XOR U34353 ( .A(n1053), .B(a[229]), .Z(n33975) );
  NANDN U34354 ( .A(n33975), .B(n37424), .Z(n33846) );
  NANDN U34355 ( .A(n33844), .B(n37425), .Z(n33845) );
  AND U34356 ( .A(n33846), .B(n33845), .Z(n33913) );
  XNOR U34357 ( .A(n33914), .B(n33913), .Z(n33915) );
  XOR U34358 ( .A(n33916), .B(n33915), .Z(n33933) );
  NAND U34359 ( .A(n38490), .B(n33847), .Z(n33849) );
  XNOR U34360 ( .A(n1058), .B(a[213]), .Z(n33981) );
  NANDN U34361 ( .A(n1048), .B(n33981), .Z(n33848) );
  NAND U34362 ( .A(n33849), .B(n33848), .Z(n33889) );
  NANDN U34363 ( .A(n1059), .B(a[209]), .Z(n33890) );
  XNOR U34364 ( .A(n33889), .B(n33890), .Z(n33892) );
  NANDN U34365 ( .A(n1049), .B(a[241]), .Z(n33850) );
  XNOR U34366 ( .A(b[1]), .B(n33850), .Z(n33852) );
  IV U34367 ( .A(a[240]), .Z(n37668) );
  NANDN U34368 ( .A(n37668), .B(n1049), .Z(n33851) );
  AND U34369 ( .A(n33852), .B(n33851), .Z(n33891) );
  XOR U34370 ( .A(n33892), .B(n33891), .Z(n33931) );
  NANDN U34371 ( .A(n33853), .B(n38205), .Z(n33855) );
  XNOR U34372 ( .A(b[23]), .B(a[219]), .Z(n33984) );
  OR U34373 ( .A(n33984), .B(n38268), .Z(n33854) );
  NAND U34374 ( .A(n33855), .B(n33854), .Z(n33954) );
  XNOR U34375 ( .A(a[235]), .B(b[7]), .Z(n33987) );
  NANDN U34376 ( .A(n33987), .B(n36701), .Z(n33858) );
  NANDN U34377 ( .A(n33856), .B(n36702), .Z(n33857) );
  NAND U34378 ( .A(n33858), .B(n33857), .Z(n33951) );
  XNOR U34379 ( .A(b[25]), .B(a[217]), .Z(n33990) );
  NANDN U34380 ( .A(n33990), .B(n38325), .Z(n33861) );
  NAND U34381 ( .A(n33859), .B(n38326), .Z(n33860) );
  AND U34382 ( .A(n33861), .B(n33860), .Z(n33952) );
  XNOR U34383 ( .A(n33951), .B(n33952), .Z(n33953) );
  XNOR U34384 ( .A(n33954), .B(n33953), .Z(n33932) );
  XOR U34385 ( .A(n33931), .B(n33932), .Z(n33934) );
  XNOR U34386 ( .A(n33933), .B(n33934), .Z(n33944) );
  XOR U34387 ( .A(n33943), .B(n33944), .Z(n33994) );
  XNOR U34388 ( .A(n33993), .B(n33994), .Z(n33995) );
  XNOR U34389 ( .A(n33996), .B(n33995), .Z(n34011) );
  XNOR U34390 ( .A(n34012), .B(n34011), .Z(n34014) );
  XNOR U34391 ( .A(n34013), .B(n34014), .Z(n34008) );
  XOR U34392 ( .A(n34007), .B(n34008), .Z(n33886) );
  NANDN U34393 ( .A(n33867), .B(n33866), .Z(n33871) );
  NANDN U34394 ( .A(n33869), .B(n33868), .Z(n33870) );
  NAND U34395 ( .A(n33871), .B(n33870), .Z(n33884) );
  XNOR U34396 ( .A(n33883), .B(n33884), .Z(n33885) );
  XNOR U34397 ( .A(n33886), .B(n33885), .Z(n33878) );
  XNOR U34398 ( .A(n33877), .B(n33878), .Z(n33879) );
  XNOR U34399 ( .A(n33880), .B(n33879), .Z(n34017) );
  XNOR U34400 ( .A(n34017), .B(sreg[465]), .Z(n34019) );
  NAND U34401 ( .A(n33872), .B(sreg[464]), .Z(n33876) );
  OR U34402 ( .A(n33874), .B(n33873), .Z(n33875) );
  AND U34403 ( .A(n33876), .B(n33875), .Z(n34018) );
  XOR U34404 ( .A(n34019), .B(n34018), .Z(c[465]) );
  NANDN U34405 ( .A(n33878), .B(n33877), .Z(n33882) );
  NAND U34406 ( .A(n33880), .B(n33879), .Z(n33881) );
  NAND U34407 ( .A(n33882), .B(n33881), .Z(n34025) );
  NANDN U34408 ( .A(n33884), .B(n33883), .Z(n33888) );
  NAND U34409 ( .A(n33886), .B(n33885), .Z(n33887) );
  NAND U34410 ( .A(n33888), .B(n33887), .Z(n34023) );
  NANDN U34411 ( .A(n33890), .B(n33889), .Z(n33894) );
  NAND U34412 ( .A(n33892), .B(n33891), .Z(n33893) );
  NAND U34413 ( .A(n33894), .B(n33893), .Z(n34105) );
  XNOR U34414 ( .A(b[19]), .B(a[224]), .Z(n34048) );
  NANDN U34415 ( .A(n34048), .B(n37934), .Z(n33897) );
  NANDN U34416 ( .A(n33895), .B(n37935), .Z(n33896) );
  NAND U34417 ( .A(n33897), .B(n33896), .Z(n34115) );
  XOR U34418 ( .A(b[27]), .B(a[216]), .Z(n34051) );
  NAND U34419 ( .A(n38423), .B(n34051), .Z(n33900) );
  NANDN U34420 ( .A(n33898), .B(n38424), .Z(n33899) );
  NAND U34421 ( .A(n33900), .B(n33899), .Z(n34112) );
  XOR U34422 ( .A(a[238]), .B(n1051), .Z(n34054) );
  NANDN U34423 ( .A(n34054), .B(n36587), .Z(n33903) );
  NANDN U34424 ( .A(n33901), .B(n36588), .Z(n33902) );
  AND U34425 ( .A(n33903), .B(n33902), .Z(n34113) );
  XNOR U34426 ( .A(n34112), .B(n34113), .Z(n34114) );
  XNOR U34427 ( .A(n34115), .B(n34114), .Z(n34103) );
  NANDN U34428 ( .A(n33904), .B(n37762), .Z(n33906) );
  XNOR U34429 ( .A(b[17]), .B(a[226]), .Z(n34057) );
  NANDN U34430 ( .A(n34057), .B(n37764), .Z(n33905) );
  NAND U34431 ( .A(n33906), .B(n33905), .Z(n34075) );
  XNOR U34432 ( .A(b[31]), .B(a[212]), .Z(n34060) );
  NANDN U34433 ( .A(n34060), .B(n38552), .Z(n33909) );
  NANDN U34434 ( .A(n33907), .B(n38553), .Z(n33908) );
  NAND U34435 ( .A(n33909), .B(n33908), .Z(n34072) );
  OR U34436 ( .A(n33910), .B(n36105), .Z(n33912) );
  XOR U34437 ( .A(a[240]), .B(n1050), .Z(n34063) );
  NANDN U34438 ( .A(n34063), .B(n36107), .Z(n33911) );
  AND U34439 ( .A(n33912), .B(n33911), .Z(n34073) );
  XNOR U34440 ( .A(n34072), .B(n34073), .Z(n34074) );
  XOR U34441 ( .A(n34075), .B(n34074), .Z(n34102) );
  XNOR U34442 ( .A(n34103), .B(n34102), .Z(n34104) );
  XNOR U34443 ( .A(n34105), .B(n34104), .Z(n34148) );
  NANDN U34444 ( .A(n33914), .B(n33913), .Z(n33918) );
  NAND U34445 ( .A(n33916), .B(n33915), .Z(n33917) );
  NAND U34446 ( .A(n33918), .B(n33917), .Z(n34093) );
  NANDN U34447 ( .A(n33920), .B(n33919), .Z(n33924) );
  NAND U34448 ( .A(n33922), .B(n33921), .Z(n33923) );
  NAND U34449 ( .A(n33924), .B(n33923), .Z(n34091) );
  OR U34450 ( .A(n33926), .B(n33925), .Z(n33930) );
  NANDN U34451 ( .A(n33928), .B(n33927), .Z(n33929) );
  NAND U34452 ( .A(n33930), .B(n33929), .Z(n34090) );
  XNOR U34453 ( .A(n34093), .B(n34092), .Z(n34149) );
  XNOR U34454 ( .A(n34148), .B(n34149), .Z(n34150) );
  NANDN U34455 ( .A(n33932), .B(n33931), .Z(n33936) );
  OR U34456 ( .A(n33934), .B(n33933), .Z(n33935) );
  AND U34457 ( .A(n33936), .B(n33935), .Z(n34151) );
  XNOR U34458 ( .A(n34150), .B(n34151), .Z(n34035) );
  NANDN U34459 ( .A(n33942), .B(n33941), .Z(n33946) );
  NANDN U34460 ( .A(n33944), .B(n33943), .Z(n33945) );
  NAND U34461 ( .A(n33946), .B(n33945), .Z(n34157) );
  NANDN U34462 ( .A(n33952), .B(n33951), .Z(n33956) );
  NAND U34463 ( .A(n33954), .B(n33953), .Z(n33955) );
  NAND U34464 ( .A(n33956), .B(n33955), .Z(n34096) );
  NANDN U34465 ( .A(n33958), .B(n33957), .Z(n33962) );
  NAND U34466 ( .A(n33960), .B(n33959), .Z(n33961) );
  AND U34467 ( .A(n33962), .B(n33961), .Z(n34097) );
  XNOR U34468 ( .A(n34096), .B(n34097), .Z(n34098) );
  XOR U34469 ( .A(b[9]), .B(n37080), .Z(n34118) );
  NANDN U34470 ( .A(n34118), .B(n36925), .Z(n33965) );
  NANDN U34471 ( .A(n33963), .B(n36926), .Z(n33964) );
  NAND U34472 ( .A(n33965), .B(n33964), .Z(n34080) );
  XOR U34473 ( .A(b[15]), .B(n36592), .Z(n34121) );
  OR U34474 ( .A(n34121), .B(n37665), .Z(n33968) );
  NANDN U34475 ( .A(n33966), .B(n37604), .Z(n33967) );
  AND U34476 ( .A(n33968), .B(n33967), .Z(n34078) );
  XOR U34477 ( .A(b[21]), .B(n35381), .Z(n34124) );
  NANDN U34478 ( .A(n34124), .B(n38101), .Z(n33971) );
  NANDN U34479 ( .A(n33969), .B(n38102), .Z(n33970) );
  AND U34480 ( .A(n33971), .B(n33970), .Z(n34079) );
  XOR U34481 ( .A(n34080), .B(n34081), .Z(n34069) );
  XOR U34482 ( .A(b[11]), .B(n37079), .Z(n34127) );
  OR U34483 ( .A(n34127), .B(n37311), .Z(n33974) );
  NANDN U34484 ( .A(n33972), .B(n37218), .Z(n33973) );
  NAND U34485 ( .A(n33974), .B(n33973), .Z(n34067) );
  XOR U34486 ( .A(n1053), .B(a[230]), .Z(n34130) );
  NANDN U34487 ( .A(n34130), .B(n37424), .Z(n33977) );
  NANDN U34488 ( .A(n33975), .B(n37425), .Z(n33976) );
  AND U34489 ( .A(n33977), .B(n33976), .Z(n34066) );
  XNOR U34490 ( .A(n34067), .B(n34066), .Z(n34068) );
  XOR U34491 ( .A(n34069), .B(n34068), .Z(n34086) );
  NANDN U34492 ( .A(n1049), .B(a[242]), .Z(n33978) );
  XNOR U34493 ( .A(b[1]), .B(n33978), .Z(n33980) );
  NANDN U34494 ( .A(b[0]), .B(a[241]), .Z(n33979) );
  AND U34495 ( .A(n33980), .B(n33979), .Z(n34044) );
  NAND U34496 ( .A(n38490), .B(n33981), .Z(n33983) );
  XNOR U34497 ( .A(n1058), .B(a[214]), .Z(n34136) );
  NANDN U34498 ( .A(n1048), .B(n34136), .Z(n33982) );
  NAND U34499 ( .A(n33983), .B(n33982), .Z(n34042) );
  NANDN U34500 ( .A(n1059), .B(a[210]), .Z(n34043) );
  XNOR U34501 ( .A(n34042), .B(n34043), .Z(n34045) );
  XOR U34502 ( .A(n34044), .B(n34045), .Z(n34084) );
  NANDN U34503 ( .A(n33984), .B(n38205), .Z(n33986) );
  XNOR U34504 ( .A(b[23]), .B(a[220]), .Z(n34139) );
  OR U34505 ( .A(n34139), .B(n38268), .Z(n33985) );
  NAND U34506 ( .A(n33986), .B(n33985), .Z(n34109) );
  XNOR U34507 ( .A(a[236]), .B(b[7]), .Z(n34142) );
  NANDN U34508 ( .A(n34142), .B(n36701), .Z(n33989) );
  NANDN U34509 ( .A(n33987), .B(n36702), .Z(n33988) );
  NAND U34510 ( .A(n33989), .B(n33988), .Z(n34106) );
  XOR U34511 ( .A(b[25]), .B(a[218]), .Z(n34145) );
  NAND U34512 ( .A(n34145), .B(n38325), .Z(n33992) );
  NANDN U34513 ( .A(n33990), .B(n38326), .Z(n33991) );
  AND U34514 ( .A(n33992), .B(n33991), .Z(n34107) );
  XNOR U34515 ( .A(n34106), .B(n34107), .Z(n34108) );
  XNOR U34516 ( .A(n34109), .B(n34108), .Z(n34085) );
  XOR U34517 ( .A(n34084), .B(n34085), .Z(n34087) );
  XNOR U34518 ( .A(n34086), .B(n34087), .Z(n34099) );
  XOR U34519 ( .A(n34098), .B(n34099), .Z(n34155) );
  XNOR U34520 ( .A(n34154), .B(n34155), .Z(n34156) );
  XOR U34521 ( .A(n34157), .B(n34156), .Z(n34033) );
  XNOR U34522 ( .A(n34032), .B(n34033), .Z(n34034) );
  XNOR U34523 ( .A(n34035), .B(n34034), .Z(n34039) );
  NANDN U34524 ( .A(n33994), .B(n33993), .Z(n33998) );
  NAND U34525 ( .A(n33996), .B(n33995), .Z(n33997) );
  NAND U34526 ( .A(n33998), .B(n33997), .Z(n34036) );
  NANDN U34527 ( .A(n34000), .B(n33999), .Z(n34004) );
  NAND U34528 ( .A(n34002), .B(n34001), .Z(n34003) );
  NAND U34529 ( .A(n34004), .B(n34003), .Z(n34037) );
  XNOR U34530 ( .A(n34036), .B(n34037), .Z(n34038) );
  XNOR U34531 ( .A(n34039), .B(n34038), .Z(n34029) );
  NANDN U34532 ( .A(n34006), .B(n34005), .Z(n34010) );
  NANDN U34533 ( .A(n34008), .B(n34007), .Z(n34009) );
  NAND U34534 ( .A(n34010), .B(n34009), .Z(n34027) );
  OR U34535 ( .A(n34012), .B(n34011), .Z(n34016) );
  OR U34536 ( .A(n34014), .B(n34013), .Z(n34015) );
  AND U34537 ( .A(n34016), .B(n34015), .Z(n34026) );
  XNOR U34538 ( .A(n34027), .B(n34026), .Z(n34028) );
  XNOR U34539 ( .A(n34029), .B(n34028), .Z(n34022) );
  XOR U34540 ( .A(n34023), .B(n34022), .Z(n34024) );
  XNOR U34541 ( .A(n34025), .B(n34024), .Z(n34160) );
  XNOR U34542 ( .A(n34160), .B(sreg[466]), .Z(n34162) );
  NAND U34543 ( .A(n34017), .B(sreg[465]), .Z(n34021) );
  OR U34544 ( .A(n34019), .B(n34018), .Z(n34020) );
  AND U34545 ( .A(n34021), .B(n34020), .Z(n34161) );
  XOR U34546 ( .A(n34162), .B(n34161), .Z(c[466]) );
  NANDN U34547 ( .A(n34027), .B(n34026), .Z(n34031) );
  NANDN U34548 ( .A(n34029), .B(n34028), .Z(n34030) );
  NAND U34549 ( .A(n34031), .B(n34030), .Z(n34166) );
  NANDN U34550 ( .A(n34037), .B(n34036), .Z(n34041) );
  NANDN U34551 ( .A(n34039), .B(n34038), .Z(n34040) );
  NAND U34552 ( .A(n34041), .B(n34040), .Z(n34172) );
  XNOR U34553 ( .A(n34171), .B(n34172), .Z(n34173) );
  NANDN U34554 ( .A(n34043), .B(n34042), .Z(n34047) );
  NAND U34555 ( .A(n34045), .B(n34044), .Z(n34046) );
  NAND U34556 ( .A(n34047), .B(n34046), .Z(n34240) );
  XOR U34557 ( .A(b[19]), .B(n36167), .Z(n34183) );
  NANDN U34558 ( .A(n34183), .B(n37934), .Z(n34050) );
  NANDN U34559 ( .A(n34048), .B(n37935), .Z(n34049) );
  NAND U34560 ( .A(n34050), .B(n34049), .Z(n34250) );
  XNOR U34561 ( .A(b[27]), .B(a[217]), .Z(n34186) );
  NANDN U34562 ( .A(n34186), .B(n38423), .Z(n34053) );
  NAND U34563 ( .A(n34051), .B(n38424), .Z(n34052) );
  NAND U34564 ( .A(n34053), .B(n34052), .Z(n34247) );
  XNOR U34565 ( .A(a[239]), .B(b[5]), .Z(n34189) );
  NANDN U34566 ( .A(n34189), .B(n36587), .Z(n34056) );
  NANDN U34567 ( .A(n34054), .B(n36588), .Z(n34055) );
  AND U34568 ( .A(n34056), .B(n34055), .Z(n34248) );
  XNOR U34569 ( .A(n34247), .B(n34248), .Z(n34249) );
  XNOR U34570 ( .A(n34250), .B(n34249), .Z(n34238) );
  NANDN U34571 ( .A(n34057), .B(n37762), .Z(n34059) );
  XOR U34572 ( .A(b[17]), .B(a[227]), .Z(n34192) );
  NAND U34573 ( .A(n34192), .B(n37764), .Z(n34058) );
  NAND U34574 ( .A(n34059), .B(n34058), .Z(n34210) );
  XNOR U34575 ( .A(b[31]), .B(a[213]), .Z(n34195) );
  NANDN U34576 ( .A(n34195), .B(n38552), .Z(n34062) );
  NANDN U34577 ( .A(n34060), .B(n38553), .Z(n34061) );
  NAND U34578 ( .A(n34062), .B(n34061), .Z(n34207) );
  OR U34579 ( .A(n34063), .B(n36105), .Z(n34065) );
  XNOR U34580 ( .A(a[241]), .B(b[3]), .Z(n34198) );
  NANDN U34581 ( .A(n34198), .B(n36107), .Z(n34064) );
  AND U34582 ( .A(n34065), .B(n34064), .Z(n34208) );
  XNOR U34583 ( .A(n34207), .B(n34208), .Z(n34209) );
  XOR U34584 ( .A(n34210), .B(n34209), .Z(n34237) );
  XNOR U34585 ( .A(n34238), .B(n34237), .Z(n34239) );
  XNOR U34586 ( .A(n34240), .B(n34239), .Z(n34283) );
  NANDN U34587 ( .A(n34067), .B(n34066), .Z(n34071) );
  NAND U34588 ( .A(n34069), .B(n34068), .Z(n34070) );
  NAND U34589 ( .A(n34071), .B(n34070), .Z(n34228) );
  NANDN U34590 ( .A(n34073), .B(n34072), .Z(n34077) );
  NAND U34591 ( .A(n34075), .B(n34074), .Z(n34076) );
  NAND U34592 ( .A(n34077), .B(n34076), .Z(n34226) );
  OR U34593 ( .A(n34079), .B(n34078), .Z(n34083) );
  NANDN U34594 ( .A(n34081), .B(n34080), .Z(n34082) );
  NAND U34595 ( .A(n34083), .B(n34082), .Z(n34225) );
  XNOR U34596 ( .A(n34228), .B(n34227), .Z(n34284) );
  XOR U34597 ( .A(n34283), .B(n34284), .Z(n34286) );
  NANDN U34598 ( .A(n34085), .B(n34084), .Z(n34089) );
  OR U34599 ( .A(n34087), .B(n34086), .Z(n34088) );
  NAND U34600 ( .A(n34089), .B(n34088), .Z(n34285) );
  XOR U34601 ( .A(n34286), .B(n34285), .Z(n34303) );
  OR U34602 ( .A(n34091), .B(n34090), .Z(n34095) );
  NAND U34603 ( .A(n34093), .B(n34092), .Z(n34094) );
  NAND U34604 ( .A(n34095), .B(n34094), .Z(n34302) );
  NANDN U34605 ( .A(n34097), .B(n34096), .Z(n34101) );
  NANDN U34606 ( .A(n34099), .B(n34098), .Z(n34100) );
  NAND U34607 ( .A(n34101), .B(n34100), .Z(n34291) );
  NANDN U34608 ( .A(n34107), .B(n34106), .Z(n34111) );
  NAND U34609 ( .A(n34109), .B(n34108), .Z(n34110) );
  NAND U34610 ( .A(n34111), .B(n34110), .Z(n34231) );
  NANDN U34611 ( .A(n34113), .B(n34112), .Z(n34117) );
  NAND U34612 ( .A(n34115), .B(n34114), .Z(n34116) );
  AND U34613 ( .A(n34117), .B(n34116), .Z(n34232) );
  XNOR U34614 ( .A(n34231), .B(n34232), .Z(n34233) );
  XOR U34615 ( .A(b[9]), .B(n37420), .Z(n34253) );
  NANDN U34616 ( .A(n34253), .B(n36925), .Z(n34120) );
  NANDN U34617 ( .A(n34118), .B(n36926), .Z(n34119) );
  NAND U34618 ( .A(n34120), .B(n34119), .Z(n34215) );
  XNOR U34619 ( .A(b[15]), .B(a[229]), .Z(n34256) );
  OR U34620 ( .A(n34256), .B(n37665), .Z(n34123) );
  NANDN U34621 ( .A(n34121), .B(n37604), .Z(n34122) );
  AND U34622 ( .A(n34123), .B(n34122), .Z(n34213) );
  XNOR U34623 ( .A(b[21]), .B(a[223]), .Z(n34259) );
  NANDN U34624 ( .A(n34259), .B(n38101), .Z(n34126) );
  NANDN U34625 ( .A(n34124), .B(n38102), .Z(n34125) );
  AND U34626 ( .A(n34126), .B(n34125), .Z(n34214) );
  XOR U34627 ( .A(n34215), .B(n34216), .Z(n34204) );
  XOR U34628 ( .A(b[11]), .B(n37184), .Z(n34262) );
  OR U34629 ( .A(n34262), .B(n37311), .Z(n34129) );
  NANDN U34630 ( .A(n34127), .B(n37218), .Z(n34128) );
  NAND U34631 ( .A(n34129), .B(n34128), .Z(n34202) );
  XOR U34632 ( .A(n1053), .B(a[231]), .Z(n34265) );
  NANDN U34633 ( .A(n34265), .B(n37424), .Z(n34132) );
  NANDN U34634 ( .A(n34130), .B(n37425), .Z(n34131) );
  AND U34635 ( .A(n34132), .B(n34131), .Z(n34201) );
  XNOR U34636 ( .A(n34202), .B(n34201), .Z(n34203) );
  XOR U34637 ( .A(n34204), .B(n34203), .Z(n34221) );
  NANDN U34638 ( .A(n1049), .B(a[243]), .Z(n34133) );
  XNOR U34639 ( .A(b[1]), .B(n34133), .Z(n34135) );
  IV U34640 ( .A(a[242]), .Z(n37676) );
  NANDN U34641 ( .A(n37676), .B(n1049), .Z(n34134) );
  AND U34642 ( .A(n34135), .B(n34134), .Z(n34179) );
  NAND U34643 ( .A(n38490), .B(n34136), .Z(n34138) );
  XOR U34644 ( .A(n1058), .B(n34725), .Z(n34271) );
  NANDN U34645 ( .A(n1048), .B(n34271), .Z(n34137) );
  NAND U34646 ( .A(n34138), .B(n34137), .Z(n34177) );
  NANDN U34647 ( .A(n1059), .B(a[211]), .Z(n34178) );
  XNOR U34648 ( .A(n34177), .B(n34178), .Z(n34180) );
  XOR U34649 ( .A(n34179), .B(n34180), .Z(n34219) );
  NANDN U34650 ( .A(n34139), .B(n38205), .Z(n34141) );
  XNOR U34651 ( .A(b[23]), .B(a[221]), .Z(n34274) );
  OR U34652 ( .A(n34274), .B(n38268), .Z(n34140) );
  NAND U34653 ( .A(n34141), .B(n34140), .Z(n34244) );
  XOR U34654 ( .A(a[237]), .B(b[7]), .Z(n34277) );
  NAND U34655 ( .A(n34277), .B(n36701), .Z(n34144) );
  NANDN U34656 ( .A(n34142), .B(n36702), .Z(n34143) );
  NAND U34657 ( .A(n34144), .B(n34143), .Z(n34241) );
  XOR U34658 ( .A(b[25]), .B(a[219]), .Z(n34280) );
  NAND U34659 ( .A(n34280), .B(n38325), .Z(n34147) );
  NAND U34660 ( .A(n34145), .B(n38326), .Z(n34146) );
  AND U34661 ( .A(n34147), .B(n34146), .Z(n34242) );
  XNOR U34662 ( .A(n34241), .B(n34242), .Z(n34243) );
  XNOR U34663 ( .A(n34244), .B(n34243), .Z(n34220) );
  XOR U34664 ( .A(n34219), .B(n34220), .Z(n34222) );
  XNOR U34665 ( .A(n34221), .B(n34222), .Z(n34234) );
  XNOR U34666 ( .A(n34233), .B(n34234), .Z(n34289) );
  XNOR U34667 ( .A(n34290), .B(n34289), .Z(n34292) );
  XNOR U34668 ( .A(n34291), .B(n34292), .Z(n34301) );
  XOR U34669 ( .A(n34302), .B(n34301), .Z(n34304) );
  NANDN U34670 ( .A(n34149), .B(n34148), .Z(n34153) );
  NAND U34671 ( .A(n34151), .B(n34150), .Z(n34152) );
  NAND U34672 ( .A(n34153), .B(n34152), .Z(n34295) );
  NANDN U34673 ( .A(n34155), .B(n34154), .Z(n34159) );
  NAND U34674 ( .A(n34157), .B(n34156), .Z(n34158) );
  NAND U34675 ( .A(n34159), .B(n34158), .Z(n34296) );
  XNOR U34676 ( .A(n34295), .B(n34296), .Z(n34297) );
  XOR U34677 ( .A(n34298), .B(n34297), .Z(n34174) );
  XOR U34678 ( .A(n34173), .B(n34174), .Z(n34165) );
  XOR U34679 ( .A(n34166), .B(n34165), .Z(n34167) );
  XNOR U34680 ( .A(n34168), .B(n34167), .Z(n34307) );
  XNOR U34681 ( .A(n34307), .B(sreg[467]), .Z(n34309) );
  NAND U34682 ( .A(n34160), .B(sreg[466]), .Z(n34164) );
  OR U34683 ( .A(n34162), .B(n34161), .Z(n34163) );
  AND U34684 ( .A(n34164), .B(n34163), .Z(n34308) );
  XOR U34685 ( .A(n34309), .B(n34308), .Z(c[467]) );
  NAND U34686 ( .A(n34166), .B(n34165), .Z(n34170) );
  NAND U34687 ( .A(n34168), .B(n34167), .Z(n34169) );
  NAND U34688 ( .A(n34170), .B(n34169), .Z(n34315) );
  NANDN U34689 ( .A(n34172), .B(n34171), .Z(n34176) );
  NAND U34690 ( .A(n34174), .B(n34173), .Z(n34175) );
  NAND U34691 ( .A(n34176), .B(n34175), .Z(n34313) );
  NANDN U34692 ( .A(n34178), .B(n34177), .Z(n34182) );
  NAND U34693 ( .A(n34180), .B(n34179), .Z(n34181) );
  NAND U34694 ( .A(n34182), .B(n34181), .Z(n34399) );
  XOR U34695 ( .A(b[19]), .B(n36280), .Z(n34366) );
  NANDN U34696 ( .A(n34366), .B(n37934), .Z(n34185) );
  NANDN U34697 ( .A(n34183), .B(n37935), .Z(n34184) );
  NAND U34698 ( .A(n34185), .B(n34184), .Z(n34411) );
  XOR U34699 ( .A(b[27]), .B(a[218]), .Z(n34369) );
  NAND U34700 ( .A(n38423), .B(n34369), .Z(n34188) );
  NANDN U34701 ( .A(n34186), .B(n38424), .Z(n34187) );
  NAND U34702 ( .A(n34188), .B(n34187), .Z(n34408) );
  XOR U34703 ( .A(a[240]), .B(n1051), .Z(n34372) );
  NANDN U34704 ( .A(n34372), .B(n36587), .Z(n34191) );
  NANDN U34705 ( .A(n34189), .B(n36588), .Z(n34190) );
  AND U34706 ( .A(n34191), .B(n34190), .Z(n34409) );
  XNOR U34707 ( .A(n34408), .B(n34409), .Z(n34410) );
  XNOR U34708 ( .A(n34411), .B(n34410), .Z(n34396) );
  NAND U34709 ( .A(n34192), .B(n37762), .Z(n34194) );
  XNOR U34710 ( .A(b[17]), .B(a[228]), .Z(n34375) );
  NANDN U34711 ( .A(n34375), .B(n37764), .Z(n34193) );
  NAND U34712 ( .A(n34194), .B(n34193), .Z(n34350) );
  XNOR U34713 ( .A(b[31]), .B(a[214]), .Z(n34378) );
  NANDN U34714 ( .A(n34378), .B(n38552), .Z(n34197) );
  NANDN U34715 ( .A(n34195), .B(n38553), .Z(n34196) );
  AND U34716 ( .A(n34197), .B(n34196), .Z(n34348) );
  OR U34717 ( .A(n34198), .B(n36105), .Z(n34200) );
  XOR U34718 ( .A(a[242]), .B(n1050), .Z(n34381) );
  NANDN U34719 ( .A(n34381), .B(n36107), .Z(n34199) );
  AND U34720 ( .A(n34200), .B(n34199), .Z(n34349) );
  XOR U34721 ( .A(n34350), .B(n34351), .Z(n34397) );
  XOR U34722 ( .A(n34396), .B(n34397), .Z(n34398) );
  XNOR U34723 ( .A(n34399), .B(n34398), .Z(n34444) );
  NANDN U34724 ( .A(n34202), .B(n34201), .Z(n34206) );
  NAND U34725 ( .A(n34204), .B(n34203), .Z(n34205) );
  NAND U34726 ( .A(n34206), .B(n34205), .Z(n34387) );
  NANDN U34727 ( .A(n34208), .B(n34207), .Z(n34212) );
  NAND U34728 ( .A(n34210), .B(n34209), .Z(n34211) );
  NAND U34729 ( .A(n34212), .B(n34211), .Z(n34385) );
  OR U34730 ( .A(n34214), .B(n34213), .Z(n34218) );
  NANDN U34731 ( .A(n34216), .B(n34215), .Z(n34217) );
  NAND U34732 ( .A(n34218), .B(n34217), .Z(n34384) );
  XNOR U34733 ( .A(n34387), .B(n34386), .Z(n34445) );
  XOR U34734 ( .A(n34444), .B(n34445), .Z(n34447) );
  NANDN U34735 ( .A(n34220), .B(n34219), .Z(n34224) );
  OR U34736 ( .A(n34222), .B(n34221), .Z(n34223) );
  NAND U34737 ( .A(n34224), .B(n34223), .Z(n34446) );
  XOR U34738 ( .A(n34447), .B(n34446), .Z(n34332) );
  OR U34739 ( .A(n34226), .B(n34225), .Z(n34230) );
  NAND U34740 ( .A(n34228), .B(n34227), .Z(n34229) );
  NAND U34741 ( .A(n34230), .B(n34229), .Z(n34331) );
  NANDN U34742 ( .A(n34232), .B(n34231), .Z(n34236) );
  NANDN U34743 ( .A(n34234), .B(n34233), .Z(n34235) );
  NAND U34744 ( .A(n34236), .B(n34235), .Z(n34452) );
  NANDN U34745 ( .A(n34242), .B(n34241), .Z(n34246) );
  NAND U34746 ( .A(n34244), .B(n34243), .Z(n34245) );
  NAND U34747 ( .A(n34246), .B(n34245), .Z(n34390) );
  NANDN U34748 ( .A(n34248), .B(n34247), .Z(n34252) );
  NAND U34749 ( .A(n34250), .B(n34249), .Z(n34251) );
  AND U34750 ( .A(n34252), .B(n34251), .Z(n34391) );
  XNOR U34751 ( .A(n34390), .B(n34391), .Z(n34392) );
  XOR U34752 ( .A(a[236]), .B(n1052), .Z(n34414) );
  NANDN U34753 ( .A(n34414), .B(n36925), .Z(n34255) );
  NANDN U34754 ( .A(n34253), .B(n36926), .Z(n34254) );
  NAND U34755 ( .A(n34255), .B(n34254), .Z(n34356) );
  XOR U34756 ( .A(b[15]), .B(n36333), .Z(n34417) );
  OR U34757 ( .A(n34417), .B(n37665), .Z(n34258) );
  NANDN U34758 ( .A(n34256), .B(n37604), .Z(n34257) );
  AND U34759 ( .A(n34258), .B(n34257), .Z(n34354) );
  XNOR U34760 ( .A(b[21]), .B(a[224]), .Z(n34420) );
  NANDN U34761 ( .A(n34420), .B(n38101), .Z(n34261) );
  NANDN U34762 ( .A(n34259), .B(n38102), .Z(n34260) );
  AND U34763 ( .A(n34261), .B(n34260), .Z(n34355) );
  XOR U34764 ( .A(n34356), .B(n34357), .Z(n34345) );
  XOR U34765 ( .A(b[11]), .B(n37080), .Z(n34423) );
  OR U34766 ( .A(n34423), .B(n37311), .Z(n34264) );
  NANDN U34767 ( .A(n34262), .B(n37218), .Z(n34263) );
  NAND U34768 ( .A(n34264), .B(n34263), .Z(n34343) );
  XOR U34769 ( .A(n1053), .B(a[232]), .Z(n34426) );
  NANDN U34770 ( .A(n34426), .B(n37424), .Z(n34267) );
  NANDN U34771 ( .A(n34265), .B(n37425), .Z(n34266) );
  NAND U34772 ( .A(n34267), .B(n34266), .Z(n34342) );
  XOR U34773 ( .A(n34345), .B(n34344), .Z(n34339) );
  NANDN U34774 ( .A(n1049), .B(a[244]), .Z(n34268) );
  XNOR U34775 ( .A(b[1]), .B(n34268), .Z(n34270) );
  IV U34776 ( .A(a[243]), .Z(n38110) );
  NANDN U34777 ( .A(n38110), .B(n1049), .Z(n34269) );
  AND U34778 ( .A(n34270), .B(n34269), .Z(n34362) );
  NAND U34779 ( .A(n38490), .B(n34271), .Z(n34273) );
  XNOR U34780 ( .A(n1058), .B(a[216]), .Z(n34432) );
  NANDN U34781 ( .A(n1048), .B(n34432), .Z(n34272) );
  NAND U34782 ( .A(n34273), .B(n34272), .Z(n34360) );
  NANDN U34783 ( .A(n1059), .B(a[212]), .Z(n34361) );
  XNOR U34784 ( .A(n34360), .B(n34361), .Z(n34363) );
  XNOR U34785 ( .A(n34362), .B(n34363), .Z(n34337) );
  NANDN U34786 ( .A(n34274), .B(n38205), .Z(n34276) );
  XOR U34787 ( .A(b[23]), .B(n35381), .Z(n34435) );
  OR U34788 ( .A(n34435), .B(n38268), .Z(n34275) );
  NAND U34789 ( .A(n34276), .B(n34275), .Z(n34405) );
  XNOR U34790 ( .A(a[238]), .B(b[7]), .Z(n34438) );
  NANDN U34791 ( .A(n34438), .B(n36701), .Z(n34279) );
  NAND U34792 ( .A(n34277), .B(n36702), .Z(n34278) );
  NAND U34793 ( .A(n34279), .B(n34278), .Z(n34402) );
  XOR U34794 ( .A(b[25]), .B(a[220]), .Z(n34441) );
  NAND U34795 ( .A(n34441), .B(n38325), .Z(n34282) );
  NAND U34796 ( .A(n34280), .B(n38326), .Z(n34281) );
  AND U34797 ( .A(n34282), .B(n34281), .Z(n34403) );
  XNOR U34798 ( .A(n34402), .B(n34403), .Z(n34404) );
  XOR U34799 ( .A(n34405), .B(n34404), .Z(n34336) );
  XOR U34800 ( .A(n34339), .B(n34338), .Z(n34393) );
  XNOR U34801 ( .A(n34392), .B(n34393), .Z(n34450) );
  XNOR U34802 ( .A(n34451), .B(n34450), .Z(n34453) );
  XNOR U34803 ( .A(n34452), .B(n34453), .Z(n34330) );
  XOR U34804 ( .A(n34331), .B(n34330), .Z(n34333) );
  NANDN U34805 ( .A(n34284), .B(n34283), .Z(n34288) );
  OR U34806 ( .A(n34286), .B(n34285), .Z(n34287) );
  NAND U34807 ( .A(n34288), .B(n34287), .Z(n34324) );
  NAND U34808 ( .A(n34290), .B(n34289), .Z(n34294) );
  NANDN U34809 ( .A(n34292), .B(n34291), .Z(n34293) );
  NAND U34810 ( .A(n34294), .B(n34293), .Z(n34325) );
  XNOR U34811 ( .A(n34324), .B(n34325), .Z(n34326) );
  XOR U34812 ( .A(n34327), .B(n34326), .Z(n34320) );
  NANDN U34813 ( .A(n34296), .B(n34295), .Z(n34300) );
  NAND U34814 ( .A(n34298), .B(n34297), .Z(n34299) );
  NAND U34815 ( .A(n34300), .B(n34299), .Z(n34318) );
  NANDN U34816 ( .A(n34302), .B(n34301), .Z(n34306) );
  OR U34817 ( .A(n34304), .B(n34303), .Z(n34305) );
  NAND U34818 ( .A(n34306), .B(n34305), .Z(n34319) );
  XNOR U34819 ( .A(n34318), .B(n34319), .Z(n34321) );
  XOR U34820 ( .A(n34320), .B(n34321), .Z(n34312) );
  XOR U34821 ( .A(n34313), .B(n34312), .Z(n34314) );
  XNOR U34822 ( .A(n34315), .B(n34314), .Z(n34456) );
  XNOR U34823 ( .A(n34456), .B(sreg[468]), .Z(n34458) );
  NAND U34824 ( .A(n34307), .B(sreg[467]), .Z(n34311) );
  OR U34825 ( .A(n34309), .B(n34308), .Z(n34310) );
  AND U34826 ( .A(n34311), .B(n34310), .Z(n34457) );
  XOR U34827 ( .A(n34458), .B(n34457), .Z(c[468]) );
  NAND U34828 ( .A(n34313), .B(n34312), .Z(n34317) );
  NAND U34829 ( .A(n34315), .B(n34314), .Z(n34316) );
  NAND U34830 ( .A(n34317), .B(n34316), .Z(n34464) );
  NANDN U34831 ( .A(n34319), .B(n34318), .Z(n34323) );
  NAND U34832 ( .A(n34321), .B(n34320), .Z(n34322) );
  NAND U34833 ( .A(n34323), .B(n34322), .Z(n34462) );
  NANDN U34834 ( .A(n34325), .B(n34324), .Z(n34329) );
  NAND U34835 ( .A(n34327), .B(n34326), .Z(n34328) );
  NAND U34836 ( .A(n34329), .B(n34328), .Z(n34467) );
  NANDN U34837 ( .A(n34331), .B(n34330), .Z(n34335) );
  OR U34838 ( .A(n34333), .B(n34332), .Z(n34334) );
  NAND U34839 ( .A(n34335), .B(n34334), .Z(n34468) );
  XNOR U34840 ( .A(n34467), .B(n34468), .Z(n34469) );
  NANDN U34841 ( .A(n34337), .B(n34336), .Z(n34341) );
  NANDN U34842 ( .A(n34339), .B(n34338), .Z(n34340) );
  NAND U34843 ( .A(n34341), .B(n34340), .Z(n34584) );
  OR U34844 ( .A(n34343), .B(n34342), .Z(n34347) );
  NAND U34845 ( .A(n34345), .B(n34344), .Z(n34346) );
  NAND U34846 ( .A(n34347), .B(n34346), .Z(n34523) );
  OR U34847 ( .A(n34349), .B(n34348), .Z(n34353) );
  NANDN U34848 ( .A(n34351), .B(n34350), .Z(n34352) );
  NAND U34849 ( .A(n34353), .B(n34352), .Z(n34522) );
  OR U34850 ( .A(n34355), .B(n34354), .Z(n34359) );
  NANDN U34851 ( .A(n34357), .B(n34356), .Z(n34358) );
  NAND U34852 ( .A(n34359), .B(n34358), .Z(n34521) );
  XOR U34853 ( .A(n34523), .B(n34524), .Z(n34581) );
  NANDN U34854 ( .A(n34361), .B(n34360), .Z(n34365) );
  NAND U34855 ( .A(n34363), .B(n34362), .Z(n34364) );
  NAND U34856 ( .A(n34365), .B(n34364), .Z(n34536) );
  XNOR U34857 ( .A(b[19]), .B(a[227]), .Z(n34479) );
  NANDN U34858 ( .A(n34479), .B(n37934), .Z(n34368) );
  NANDN U34859 ( .A(n34366), .B(n37935), .Z(n34367) );
  NAND U34860 ( .A(n34368), .B(n34367), .Z(n34548) );
  XOR U34861 ( .A(b[27]), .B(a[219]), .Z(n34482) );
  NAND U34862 ( .A(n38423), .B(n34482), .Z(n34371) );
  NAND U34863 ( .A(n34369), .B(n38424), .Z(n34370) );
  NAND U34864 ( .A(n34371), .B(n34370), .Z(n34545) );
  XNOR U34865 ( .A(a[241]), .B(b[5]), .Z(n34485) );
  NANDN U34866 ( .A(n34485), .B(n36587), .Z(n34374) );
  NANDN U34867 ( .A(n34372), .B(n36588), .Z(n34373) );
  AND U34868 ( .A(n34374), .B(n34373), .Z(n34546) );
  XNOR U34869 ( .A(n34545), .B(n34546), .Z(n34547) );
  XNOR U34870 ( .A(n34548), .B(n34547), .Z(n34534) );
  NANDN U34871 ( .A(n34375), .B(n37762), .Z(n34377) );
  XOR U34872 ( .A(b[17]), .B(a[229]), .Z(n34488) );
  NAND U34873 ( .A(n34488), .B(n37764), .Z(n34376) );
  NAND U34874 ( .A(n34377), .B(n34376), .Z(n34506) );
  XOR U34875 ( .A(n1059), .B(n34725), .Z(n34491) );
  NAND U34876 ( .A(n34491), .B(n38552), .Z(n34380) );
  NANDN U34877 ( .A(n34378), .B(n38553), .Z(n34379) );
  NAND U34878 ( .A(n34380), .B(n34379), .Z(n34503) );
  OR U34879 ( .A(n34381), .B(n36105), .Z(n34383) );
  XOR U34880 ( .A(a[243]), .B(n1050), .Z(n34494) );
  NANDN U34881 ( .A(n34494), .B(n36107), .Z(n34382) );
  AND U34882 ( .A(n34383), .B(n34382), .Z(n34504) );
  XNOR U34883 ( .A(n34503), .B(n34504), .Z(n34505) );
  XOR U34884 ( .A(n34506), .B(n34505), .Z(n34533) );
  XNOR U34885 ( .A(n34534), .B(n34533), .Z(n34535) );
  XNOR U34886 ( .A(n34536), .B(n34535), .Z(n34582) );
  XNOR U34887 ( .A(n34581), .B(n34582), .Z(n34583) );
  XNOR U34888 ( .A(n34584), .B(n34583), .Z(n34602) );
  OR U34889 ( .A(n34385), .B(n34384), .Z(n34389) );
  NAND U34890 ( .A(n34387), .B(n34386), .Z(n34388) );
  NAND U34891 ( .A(n34389), .B(n34388), .Z(n34600) );
  NANDN U34892 ( .A(n34391), .B(n34390), .Z(n34395) );
  NANDN U34893 ( .A(n34393), .B(n34392), .Z(n34394) );
  NAND U34894 ( .A(n34395), .B(n34394), .Z(n34589) );
  OR U34895 ( .A(n34397), .B(n34396), .Z(n34401) );
  NAND U34896 ( .A(n34399), .B(n34398), .Z(n34400) );
  NAND U34897 ( .A(n34401), .B(n34400), .Z(n34588) );
  NANDN U34898 ( .A(n34403), .B(n34402), .Z(n34407) );
  NAND U34899 ( .A(n34405), .B(n34404), .Z(n34406) );
  NAND U34900 ( .A(n34407), .B(n34406), .Z(n34527) );
  NANDN U34901 ( .A(n34409), .B(n34408), .Z(n34413) );
  NAND U34902 ( .A(n34411), .B(n34410), .Z(n34412) );
  AND U34903 ( .A(n34413), .B(n34412), .Z(n34528) );
  XNOR U34904 ( .A(n34527), .B(n34528), .Z(n34529) );
  XNOR U34905 ( .A(a[237]), .B(n1052), .Z(n34551) );
  NAND U34906 ( .A(n36925), .B(n34551), .Z(n34416) );
  NANDN U34907 ( .A(n34414), .B(n36926), .Z(n34415) );
  NAND U34908 ( .A(n34416), .B(n34415), .Z(n34511) );
  XOR U34909 ( .A(b[15]), .B(n36934), .Z(n34554) );
  OR U34910 ( .A(n34554), .B(n37665), .Z(n34419) );
  NANDN U34911 ( .A(n34417), .B(n37604), .Z(n34418) );
  AND U34912 ( .A(n34419), .B(n34418), .Z(n34509) );
  XOR U34913 ( .A(b[21]), .B(n36167), .Z(n34557) );
  NANDN U34914 ( .A(n34557), .B(n38101), .Z(n34422) );
  NANDN U34915 ( .A(n34420), .B(n38102), .Z(n34421) );
  AND U34916 ( .A(n34422), .B(n34421), .Z(n34510) );
  XOR U34917 ( .A(n34511), .B(n34512), .Z(n34500) );
  XOR U34918 ( .A(b[11]), .B(n37420), .Z(n34560) );
  OR U34919 ( .A(n34560), .B(n37311), .Z(n34425) );
  NANDN U34920 ( .A(n34423), .B(n37218), .Z(n34424) );
  NAND U34921 ( .A(n34425), .B(n34424), .Z(n34498) );
  XOR U34922 ( .A(b[13]), .B(n37184), .Z(n34563) );
  NANDN U34923 ( .A(n34563), .B(n37424), .Z(n34428) );
  NANDN U34924 ( .A(n34426), .B(n37425), .Z(n34427) );
  AND U34925 ( .A(n34428), .B(n34427), .Z(n34497) );
  XNOR U34926 ( .A(n34498), .B(n34497), .Z(n34499) );
  XOR U34927 ( .A(n34500), .B(n34499), .Z(n34517) );
  NANDN U34928 ( .A(n1049), .B(a[245]), .Z(n34429) );
  XNOR U34929 ( .A(b[1]), .B(n34429), .Z(n34431) );
  IV U34930 ( .A(a[244]), .Z(n38034) );
  NANDN U34931 ( .A(n38034), .B(n1049), .Z(n34430) );
  AND U34932 ( .A(n34431), .B(n34430), .Z(n34475) );
  NAND U34933 ( .A(n38490), .B(n34432), .Z(n34434) );
  XOR U34934 ( .A(n1058), .B(n34670), .Z(n34569) );
  NANDN U34935 ( .A(n1048), .B(n34569), .Z(n34433) );
  NAND U34936 ( .A(n34434), .B(n34433), .Z(n34473) );
  NANDN U34937 ( .A(n1059), .B(a[213]), .Z(n34474) );
  XNOR U34938 ( .A(n34473), .B(n34474), .Z(n34476) );
  XOR U34939 ( .A(n34475), .B(n34476), .Z(n34515) );
  NANDN U34940 ( .A(n34435), .B(n38205), .Z(n34437) );
  XNOR U34941 ( .A(b[23]), .B(a[223]), .Z(n34572) );
  OR U34942 ( .A(n34572), .B(n38268), .Z(n34436) );
  NAND U34943 ( .A(n34437), .B(n34436), .Z(n34542) );
  XOR U34944 ( .A(a[239]), .B(b[7]), .Z(n34575) );
  NAND U34945 ( .A(n34575), .B(n36701), .Z(n34440) );
  NANDN U34946 ( .A(n34438), .B(n36702), .Z(n34439) );
  NAND U34947 ( .A(n34440), .B(n34439), .Z(n34539) );
  XOR U34948 ( .A(b[25]), .B(a[221]), .Z(n34578) );
  NAND U34949 ( .A(n34578), .B(n38325), .Z(n34443) );
  NAND U34950 ( .A(n34441), .B(n38326), .Z(n34442) );
  AND U34951 ( .A(n34443), .B(n34442), .Z(n34540) );
  XNOR U34952 ( .A(n34539), .B(n34540), .Z(n34541) );
  XNOR U34953 ( .A(n34542), .B(n34541), .Z(n34516) );
  XOR U34954 ( .A(n34515), .B(n34516), .Z(n34518) );
  XNOR U34955 ( .A(n34517), .B(n34518), .Z(n34530) );
  XNOR U34956 ( .A(n34529), .B(n34530), .Z(n34587) );
  XNOR U34957 ( .A(n34588), .B(n34587), .Z(n34590) );
  XNOR U34958 ( .A(n34589), .B(n34590), .Z(n34599) );
  XNOR U34959 ( .A(n34600), .B(n34599), .Z(n34601) );
  XOR U34960 ( .A(n34602), .B(n34601), .Z(n34596) );
  NANDN U34961 ( .A(n34445), .B(n34444), .Z(n34449) );
  OR U34962 ( .A(n34447), .B(n34446), .Z(n34448) );
  NAND U34963 ( .A(n34449), .B(n34448), .Z(n34593) );
  NAND U34964 ( .A(n34451), .B(n34450), .Z(n34455) );
  NANDN U34965 ( .A(n34453), .B(n34452), .Z(n34454) );
  NAND U34966 ( .A(n34455), .B(n34454), .Z(n34594) );
  XNOR U34967 ( .A(n34593), .B(n34594), .Z(n34595) );
  XOR U34968 ( .A(n34596), .B(n34595), .Z(n34470) );
  XOR U34969 ( .A(n34469), .B(n34470), .Z(n34461) );
  XOR U34970 ( .A(n34462), .B(n34461), .Z(n34463) );
  XNOR U34971 ( .A(n34464), .B(n34463), .Z(n34605) );
  XNOR U34972 ( .A(n34605), .B(sreg[469]), .Z(n34607) );
  NAND U34973 ( .A(n34456), .B(sreg[468]), .Z(n34460) );
  OR U34974 ( .A(n34458), .B(n34457), .Z(n34459) );
  AND U34975 ( .A(n34460), .B(n34459), .Z(n34606) );
  XOR U34976 ( .A(n34607), .B(n34606), .Z(c[469]) );
  NAND U34977 ( .A(n34462), .B(n34461), .Z(n34466) );
  NAND U34978 ( .A(n34464), .B(n34463), .Z(n34465) );
  NAND U34979 ( .A(n34466), .B(n34465), .Z(n34613) );
  NANDN U34980 ( .A(n34468), .B(n34467), .Z(n34472) );
  NAND U34981 ( .A(n34470), .B(n34469), .Z(n34471) );
  NAND U34982 ( .A(n34472), .B(n34471), .Z(n34611) );
  NANDN U34983 ( .A(n34474), .B(n34473), .Z(n34478) );
  NAND U34984 ( .A(n34476), .B(n34475), .Z(n34477) );
  NAND U34985 ( .A(n34478), .B(n34477), .Z(n34692) );
  XOR U34986 ( .A(b[19]), .B(n36592), .Z(n34658) );
  NANDN U34987 ( .A(n34658), .B(n37934), .Z(n34481) );
  NANDN U34988 ( .A(n34479), .B(n37935), .Z(n34480) );
  NAND U34989 ( .A(n34481), .B(n34480), .Z(n34704) );
  XOR U34990 ( .A(b[27]), .B(a[220]), .Z(n34661) );
  NAND U34991 ( .A(n38423), .B(n34661), .Z(n34484) );
  NAND U34992 ( .A(n34482), .B(n38424), .Z(n34483) );
  NAND U34993 ( .A(n34484), .B(n34483), .Z(n34701) );
  XOR U34994 ( .A(a[242]), .B(n1051), .Z(n34664) );
  NANDN U34995 ( .A(n34664), .B(n36587), .Z(n34487) );
  NANDN U34996 ( .A(n34485), .B(n36588), .Z(n34486) );
  AND U34997 ( .A(n34487), .B(n34486), .Z(n34702) );
  XNOR U34998 ( .A(n34701), .B(n34702), .Z(n34703) );
  XNOR U34999 ( .A(n34704), .B(n34703), .Z(n34689) );
  XNOR U35000 ( .A(b[17]), .B(a[230]), .Z(n34667) );
  NANDN U35001 ( .A(n34667), .B(n37764), .Z(n34490) );
  NAND U35002 ( .A(n34488), .B(n37762), .Z(n34489) );
  NAND U35003 ( .A(n34490), .B(n34489), .Z(n34646) );
  XOR U35004 ( .A(n1059), .B(a[216]), .Z(n34671) );
  NANDN U35005 ( .A(n34671), .B(n38552), .Z(n34493) );
  NAND U35006 ( .A(n38553), .B(n34491), .Z(n34492) );
  NAND U35007 ( .A(n34493), .B(n34492), .Z(n34644) );
  OR U35008 ( .A(n34494), .B(n36105), .Z(n34496) );
  XOR U35009 ( .A(a[244]), .B(n1050), .Z(n34674) );
  NANDN U35010 ( .A(n34674), .B(n36107), .Z(n34495) );
  AND U35011 ( .A(n34496), .B(n34495), .Z(n34645) );
  XNOR U35012 ( .A(n34644), .B(n34645), .Z(n34647) );
  XNOR U35013 ( .A(n34646), .B(n34647), .Z(n34690) );
  XOR U35014 ( .A(n34689), .B(n34690), .Z(n34691) );
  XNOR U35015 ( .A(n34692), .B(n34691), .Z(n34738) );
  NANDN U35016 ( .A(n34498), .B(n34497), .Z(n34502) );
  NAND U35017 ( .A(n34500), .B(n34499), .Z(n34501) );
  NAND U35018 ( .A(n34502), .B(n34501), .Z(n34680) );
  NANDN U35019 ( .A(n34504), .B(n34503), .Z(n34508) );
  NAND U35020 ( .A(n34506), .B(n34505), .Z(n34507) );
  NAND U35021 ( .A(n34508), .B(n34507), .Z(n34678) );
  OR U35022 ( .A(n34510), .B(n34509), .Z(n34514) );
  NANDN U35023 ( .A(n34512), .B(n34511), .Z(n34513) );
  NAND U35024 ( .A(n34514), .B(n34513), .Z(n34677) );
  XNOR U35025 ( .A(n34680), .B(n34679), .Z(n34739) );
  XOR U35026 ( .A(n34738), .B(n34739), .Z(n34741) );
  NANDN U35027 ( .A(n34516), .B(n34515), .Z(n34520) );
  OR U35028 ( .A(n34518), .B(n34517), .Z(n34519) );
  NAND U35029 ( .A(n34520), .B(n34519), .Z(n34740) );
  XOR U35030 ( .A(n34741), .B(n34740), .Z(n34630) );
  OR U35031 ( .A(n34522), .B(n34521), .Z(n34526) );
  NANDN U35032 ( .A(n34524), .B(n34523), .Z(n34525) );
  NAND U35033 ( .A(n34526), .B(n34525), .Z(n34629) );
  NANDN U35034 ( .A(n34528), .B(n34527), .Z(n34532) );
  NANDN U35035 ( .A(n34530), .B(n34529), .Z(n34531) );
  NAND U35036 ( .A(n34532), .B(n34531), .Z(n34746) );
  NANDN U35037 ( .A(n34534), .B(n34533), .Z(n34538) );
  NAND U35038 ( .A(n34536), .B(n34535), .Z(n34537) );
  NAND U35039 ( .A(n34538), .B(n34537), .Z(n34745) );
  NANDN U35040 ( .A(n34540), .B(n34539), .Z(n34544) );
  NAND U35041 ( .A(n34542), .B(n34541), .Z(n34543) );
  NAND U35042 ( .A(n34544), .B(n34543), .Z(n34683) );
  NANDN U35043 ( .A(n34546), .B(n34545), .Z(n34550) );
  NAND U35044 ( .A(n34548), .B(n34547), .Z(n34549) );
  AND U35045 ( .A(n34550), .B(n34549), .Z(n34684) );
  XNOR U35046 ( .A(n34683), .B(n34684), .Z(n34685) );
  XOR U35047 ( .A(n37467), .B(b[9]), .Z(n34713) );
  NANDN U35048 ( .A(n34713), .B(n36925), .Z(n34553) );
  NAND U35049 ( .A(n36926), .B(n34551), .Z(n34552) );
  NAND U35050 ( .A(n34553), .B(n34552), .Z(n34650) );
  XNOR U35051 ( .A(n1054), .B(a[232]), .Z(n34710) );
  NANDN U35052 ( .A(n37665), .B(n34710), .Z(n34556) );
  NANDN U35053 ( .A(n34554), .B(n37604), .Z(n34555) );
  NAND U35054 ( .A(n34556), .B(n34555), .Z(n34648) );
  XOR U35055 ( .A(n1056), .B(n36280), .Z(n34707) );
  NAND U35056 ( .A(n34707), .B(n38101), .Z(n34559) );
  NANDN U35057 ( .A(n34557), .B(n38102), .Z(n34558) );
  AND U35058 ( .A(n34559), .B(n34558), .Z(n34649) );
  XNOR U35059 ( .A(n34648), .B(n34649), .Z(n34651) );
  XOR U35060 ( .A(n34650), .B(n34651), .Z(n34643) );
  XOR U35061 ( .A(b[11]), .B(n37106), .Z(n34716) );
  OR U35062 ( .A(n34716), .B(n37311), .Z(n34562) );
  NANDN U35063 ( .A(n34560), .B(n37218), .Z(n34561) );
  NAND U35064 ( .A(n34562), .B(n34561), .Z(n34641) );
  XOR U35065 ( .A(b[13]), .B(n37080), .Z(n34719) );
  NANDN U35066 ( .A(n34719), .B(n37424), .Z(n34565) );
  NANDN U35067 ( .A(n34563), .B(n37425), .Z(n34564) );
  AND U35068 ( .A(n34565), .B(n34564), .Z(n34640) );
  XNOR U35069 ( .A(n34641), .B(n34640), .Z(n34642) );
  XNOR U35070 ( .A(n34643), .B(n34642), .Z(n34636) );
  NANDN U35071 ( .A(n1049), .B(a[246]), .Z(n34566) );
  XNOR U35072 ( .A(b[1]), .B(n34566), .Z(n34568) );
  IV U35073 ( .A(a[245]), .Z(n38213) );
  NANDN U35074 ( .A(n38213), .B(n1049), .Z(n34567) );
  AND U35075 ( .A(n34568), .B(n34567), .Z(n34654) );
  NAND U35076 ( .A(n38490), .B(n34569), .Z(n34571) );
  XNOR U35077 ( .A(b[29]), .B(a[218]), .Z(n34726) );
  OR U35078 ( .A(n34726), .B(n1048), .Z(n34570) );
  NAND U35079 ( .A(n34571), .B(n34570), .Z(n34652) );
  NANDN U35080 ( .A(n1059), .B(a[214]), .Z(n34653) );
  XNOR U35081 ( .A(n34652), .B(n34653), .Z(n34655) );
  XOR U35082 ( .A(n34654), .B(n34655), .Z(n34634) );
  NANDN U35083 ( .A(n34572), .B(n38205), .Z(n34574) );
  XNOR U35084 ( .A(b[23]), .B(a[224]), .Z(n34729) );
  OR U35085 ( .A(n34729), .B(n38268), .Z(n34573) );
  NAND U35086 ( .A(n34574), .B(n34573), .Z(n34698) );
  XNOR U35087 ( .A(a[240]), .B(b[7]), .Z(n34732) );
  NANDN U35088 ( .A(n34732), .B(n36701), .Z(n34577) );
  NAND U35089 ( .A(n34575), .B(n36702), .Z(n34576) );
  NAND U35090 ( .A(n34577), .B(n34576), .Z(n34695) );
  XNOR U35091 ( .A(b[25]), .B(a[222]), .Z(n34735) );
  NANDN U35092 ( .A(n34735), .B(n38325), .Z(n34580) );
  NAND U35093 ( .A(n34578), .B(n38326), .Z(n34579) );
  AND U35094 ( .A(n34580), .B(n34579), .Z(n34696) );
  XNOR U35095 ( .A(n34695), .B(n34696), .Z(n34697) );
  XNOR U35096 ( .A(n34698), .B(n34697), .Z(n34635) );
  XOR U35097 ( .A(n34634), .B(n34635), .Z(n34637) );
  XOR U35098 ( .A(n34685), .B(n34686), .Z(n34744) );
  XNOR U35099 ( .A(n34745), .B(n34744), .Z(n34747) );
  XNOR U35100 ( .A(n34746), .B(n34747), .Z(n34628) );
  XOR U35101 ( .A(n34629), .B(n34628), .Z(n34631) );
  NANDN U35102 ( .A(n34582), .B(n34581), .Z(n34586) );
  NAND U35103 ( .A(n34584), .B(n34583), .Z(n34585) );
  NAND U35104 ( .A(n34586), .B(n34585), .Z(n34623) );
  NAND U35105 ( .A(n34588), .B(n34587), .Z(n34592) );
  NANDN U35106 ( .A(n34590), .B(n34589), .Z(n34591) );
  AND U35107 ( .A(n34592), .B(n34591), .Z(n34622) );
  XNOR U35108 ( .A(n34623), .B(n34622), .Z(n34624) );
  XOR U35109 ( .A(n34625), .B(n34624), .Z(n34618) );
  NANDN U35110 ( .A(n34594), .B(n34593), .Z(n34598) );
  NAND U35111 ( .A(n34596), .B(n34595), .Z(n34597) );
  NAND U35112 ( .A(n34598), .B(n34597), .Z(n34616) );
  NANDN U35113 ( .A(n34600), .B(n34599), .Z(n34604) );
  NANDN U35114 ( .A(n34602), .B(n34601), .Z(n34603) );
  NAND U35115 ( .A(n34604), .B(n34603), .Z(n34617) );
  XNOR U35116 ( .A(n34616), .B(n34617), .Z(n34619) );
  XOR U35117 ( .A(n34618), .B(n34619), .Z(n34610) );
  XOR U35118 ( .A(n34611), .B(n34610), .Z(n34612) );
  XNOR U35119 ( .A(n34613), .B(n34612), .Z(n34750) );
  XNOR U35120 ( .A(n34750), .B(sreg[470]), .Z(n34752) );
  NAND U35121 ( .A(n34605), .B(sreg[469]), .Z(n34609) );
  OR U35122 ( .A(n34607), .B(n34606), .Z(n34608) );
  AND U35123 ( .A(n34609), .B(n34608), .Z(n34751) );
  XOR U35124 ( .A(n34752), .B(n34751), .Z(c[470]) );
  NAND U35125 ( .A(n34611), .B(n34610), .Z(n34615) );
  NAND U35126 ( .A(n34613), .B(n34612), .Z(n34614) );
  NAND U35127 ( .A(n34615), .B(n34614), .Z(n34758) );
  NANDN U35128 ( .A(n34617), .B(n34616), .Z(n34621) );
  NAND U35129 ( .A(n34619), .B(n34618), .Z(n34620) );
  NAND U35130 ( .A(n34621), .B(n34620), .Z(n34756) );
  NANDN U35131 ( .A(n34623), .B(n34622), .Z(n34627) );
  NAND U35132 ( .A(n34625), .B(n34624), .Z(n34626) );
  NAND U35133 ( .A(n34627), .B(n34626), .Z(n34761) );
  NANDN U35134 ( .A(n34629), .B(n34628), .Z(n34633) );
  OR U35135 ( .A(n34631), .B(n34630), .Z(n34632) );
  NAND U35136 ( .A(n34633), .B(n34632), .Z(n34762) );
  XNOR U35137 ( .A(n34761), .B(n34762), .Z(n34763) );
  NANDN U35138 ( .A(n34635), .B(n34634), .Z(n34639) );
  OR U35139 ( .A(n34637), .B(n34636), .Z(n34638) );
  NAND U35140 ( .A(n34639), .B(n34638), .Z(n34776) );
  XNOR U35141 ( .A(n34824), .B(n34823), .Z(n34826) );
  XNOR U35142 ( .A(n34825), .B(n34826), .Z(n34774) );
  NANDN U35143 ( .A(n34653), .B(n34652), .Z(n34657) );
  NAND U35144 ( .A(n34655), .B(n34654), .Z(n34656) );
  NAND U35145 ( .A(n34657), .B(n34656), .Z(n34836) );
  XNOR U35146 ( .A(b[19]), .B(a[229]), .Z(n34785) );
  NANDN U35147 ( .A(n34785), .B(n37934), .Z(n34660) );
  NANDN U35148 ( .A(n34658), .B(n37935), .Z(n34659) );
  NAND U35149 ( .A(n34660), .B(n34659), .Z(n34848) );
  XOR U35150 ( .A(b[27]), .B(a[221]), .Z(n34788) );
  NAND U35151 ( .A(n38423), .B(n34788), .Z(n34663) );
  NAND U35152 ( .A(n34661), .B(n38424), .Z(n34662) );
  NAND U35153 ( .A(n34663), .B(n34662), .Z(n34845) );
  XOR U35154 ( .A(a[243]), .B(n1051), .Z(n34791) );
  NANDN U35155 ( .A(n34791), .B(n36587), .Z(n34666) );
  NANDN U35156 ( .A(n34664), .B(n36588), .Z(n34665) );
  AND U35157 ( .A(n34666), .B(n34665), .Z(n34846) );
  XNOR U35158 ( .A(n34845), .B(n34846), .Z(n34847) );
  XNOR U35159 ( .A(n34848), .B(n34847), .Z(n34833) );
  XNOR U35160 ( .A(b[17]), .B(a[231]), .Z(n34794) );
  NANDN U35161 ( .A(n34794), .B(n37764), .Z(n34669) );
  NANDN U35162 ( .A(n34667), .B(n37762), .Z(n34668) );
  NAND U35163 ( .A(n34669), .B(n34668), .Z(n34809) );
  XOR U35164 ( .A(b[31]), .B(n34670), .Z(n34797) );
  NANDN U35165 ( .A(n34797), .B(n38552), .Z(n34673) );
  NANDN U35166 ( .A(n34671), .B(n38553), .Z(n34672) );
  NAND U35167 ( .A(n34673), .B(n34672), .Z(n34807) );
  OR U35168 ( .A(n34674), .B(n36105), .Z(n34676) );
  XOR U35169 ( .A(a[245]), .B(n1050), .Z(n34800) );
  NANDN U35170 ( .A(n34800), .B(n36107), .Z(n34675) );
  AND U35171 ( .A(n34676), .B(n34675), .Z(n34808) );
  XNOR U35172 ( .A(n34807), .B(n34808), .Z(n34810) );
  XNOR U35173 ( .A(n34809), .B(n34810), .Z(n34834) );
  XOR U35174 ( .A(n34833), .B(n34834), .Z(n34835) );
  XNOR U35175 ( .A(n34836), .B(n34835), .Z(n34773) );
  XOR U35176 ( .A(n34774), .B(n34773), .Z(n34775) );
  XNOR U35177 ( .A(n34776), .B(n34775), .Z(n34890) );
  OR U35178 ( .A(n34678), .B(n34677), .Z(n34682) );
  NAND U35179 ( .A(n34680), .B(n34679), .Z(n34681) );
  NAND U35180 ( .A(n34682), .B(n34681), .Z(n34888) );
  NANDN U35181 ( .A(n34684), .B(n34683), .Z(n34688) );
  NAND U35182 ( .A(n34686), .B(n34685), .Z(n34687) );
  NAND U35183 ( .A(n34688), .B(n34687), .Z(n34769) );
  OR U35184 ( .A(n34690), .B(n34689), .Z(n34694) );
  NAND U35185 ( .A(n34692), .B(n34691), .Z(n34693) );
  NAND U35186 ( .A(n34694), .B(n34693), .Z(n34768) );
  NANDN U35187 ( .A(n34696), .B(n34695), .Z(n34700) );
  NAND U35188 ( .A(n34698), .B(n34697), .Z(n34699) );
  NAND U35189 ( .A(n34700), .B(n34699), .Z(n34827) );
  NANDN U35190 ( .A(n34702), .B(n34701), .Z(n34706) );
  NAND U35191 ( .A(n34704), .B(n34703), .Z(n34705) );
  AND U35192 ( .A(n34706), .B(n34705), .Z(n34828) );
  XNOR U35193 ( .A(n34827), .B(n34828), .Z(n34829) );
  XNOR U35194 ( .A(b[21]), .B(a[227]), .Z(n34857) );
  NANDN U35195 ( .A(n34857), .B(n38101), .Z(n34709) );
  NAND U35196 ( .A(n38102), .B(n34707), .Z(n34708) );
  AND U35197 ( .A(n34709), .B(n34708), .Z(n34817) );
  XOR U35198 ( .A(b[15]), .B(n37184), .Z(n34854) );
  OR U35199 ( .A(n34854), .B(n37665), .Z(n34712) );
  NAND U35200 ( .A(n34710), .B(n37604), .Z(n34711) );
  AND U35201 ( .A(n34712), .B(n34711), .Z(n34818) );
  XOR U35202 ( .A(n34817), .B(n34818), .Z(n34819) );
  XNOR U35203 ( .A(a[239]), .B(b[9]), .Z(n34851) );
  NANDN U35204 ( .A(n34851), .B(n36925), .Z(n34715) );
  NANDN U35205 ( .A(n34713), .B(n36926), .Z(n34714) );
  AND U35206 ( .A(n34715), .B(n34714), .Z(n34820) );
  XNOR U35207 ( .A(n34819), .B(n34820), .Z(n34814) );
  XNOR U35208 ( .A(b[11]), .B(a[237]), .Z(n34860) );
  OR U35209 ( .A(n34860), .B(n37311), .Z(n34718) );
  NANDN U35210 ( .A(n34716), .B(n37218), .Z(n34717) );
  NAND U35211 ( .A(n34718), .B(n34717), .Z(n34812) );
  XOR U35212 ( .A(n1053), .B(n37420), .Z(n34863) );
  NAND U35213 ( .A(n34863), .B(n37424), .Z(n34721) );
  NANDN U35214 ( .A(n34719), .B(n37425), .Z(n34720) );
  NAND U35215 ( .A(n34721), .B(n34720), .Z(n34811) );
  XNOR U35216 ( .A(n34812), .B(n34811), .Z(n34813) );
  NANDN U35217 ( .A(n1049), .B(a[247]), .Z(n34722) );
  XNOR U35218 ( .A(b[1]), .B(n34722), .Z(n34724) );
  IV U35219 ( .A(a[246]), .Z(n38146) );
  NANDN U35220 ( .A(n38146), .B(n1049), .Z(n34723) );
  AND U35221 ( .A(n34724), .B(n34723), .Z(n34782) );
  ANDN U35222 ( .B(b[31]), .A(n34725), .Z(n34779) );
  NANDN U35223 ( .A(n34726), .B(n38490), .Z(n34728) );
  XNOR U35224 ( .A(n1058), .B(a[219]), .Z(n34869) );
  NANDN U35225 ( .A(n1048), .B(n34869), .Z(n34727) );
  NAND U35226 ( .A(n34728), .B(n34727), .Z(n34780) );
  XOR U35227 ( .A(n34779), .B(n34780), .Z(n34781) );
  XNOR U35228 ( .A(n34782), .B(n34781), .Z(n34803) );
  NANDN U35229 ( .A(n34729), .B(n38205), .Z(n34731) );
  XOR U35230 ( .A(b[23]), .B(n36167), .Z(n34872) );
  OR U35231 ( .A(n34872), .B(n38268), .Z(n34730) );
  NAND U35232 ( .A(n34731), .B(n34730), .Z(n34842) );
  XOR U35233 ( .A(a[241]), .B(b[7]), .Z(n34875) );
  NAND U35234 ( .A(n34875), .B(n36701), .Z(n34734) );
  NANDN U35235 ( .A(n34732), .B(n36702), .Z(n34733) );
  NAND U35236 ( .A(n34734), .B(n34733), .Z(n34839) );
  XOR U35237 ( .A(b[25]), .B(a[223]), .Z(n34878) );
  NAND U35238 ( .A(n34878), .B(n38325), .Z(n34737) );
  NANDN U35239 ( .A(n34735), .B(n38326), .Z(n34736) );
  AND U35240 ( .A(n34737), .B(n34736), .Z(n34840) );
  XNOR U35241 ( .A(n34839), .B(n34840), .Z(n34841) );
  XNOR U35242 ( .A(n34842), .B(n34841), .Z(n34804) );
  XNOR U35243 ( .A(n34803), .B(n34804), .Z(n34806) );
  XNOR U35244 ( .A(n34805), .B(n34806), .Z(n34830) );
  XOR U35245 ( .A(n34829), .B(n34830), .Z(n34767) );
  XNOR U35246 ( .A(n34768), .B(n34767), .Z(n34770) );
  XNOR U35247 ( .A(n34769), .B(n34770), .Z(n34887) );
  XNOR U35248 ( .A(n34888), .B(n34887), .Z(n34889) );
  XOR U35249 ( .A(n34890), .B(n34889), .Z(n34884) );
  NANDN U35250 ( .A(n34739), .B(n34738), .Z(n34743) );
  OR U35251 ( .A(n34741), .B(n34740), .Z(n34742) );
  NAND U35252 ( .A(n34743), .B(n34742), .Z(n34881) );
  NAND U35253 ( .A(n34745), .B(n34744), .Z(n34749) );
  NANDN U35254 ( .A(n34747), .B(n34746), .Z(n34748) );
  NAND U35255 ( .A(n34749), .B(n34748), .Z(n34882) );
  XNOR U35256 ( .A(n34881), .B(n34882), .Z(n34883) );
  XOR U35257 ( .A(n34884), .B(n34883), .Z(n34764) );
  XOR U35258 ( .A(n34763), .B(n34764), .Z(n34755) );
  XOR U35259 ( .A(n34756), .B(n34755), .Z(n34757) );
  XNOR U35260 ( .A(n34758), .B(n34757), .Z(n34893) );
  XNOR U35261 ( .A(n34893), .B(sreg[471]), .Z(n34895) );
  NAND U35262 ( .A(n34750), .B(sreg[470]), .Z(n34754) );
  OR U35263 ( .A(n34752), .B(n34751), .Z(n34753) );
  AND U35264 ( .A(n34754), .B(n34753), .Z(n34894) );
  XOR U35265 ( .A(n34895), .B(n34894), .Z(c[471]) );
  NAND U35266 ( .A(n34756), .B(n34755), .Z(n34760) );
  NAND U35267 ( .A(n34758), .B(n34757), .Z(n34759) );
  NAND U35268 ( .A(n34760), .B(n34759), .Z(n34901) );
  NANDN U35269 ( .A(n34762), .B(n34761), .Z(n34766) );
  NAND U35270 ( .A(n34764), .B(n34763), .Z(n34765) );
  NAND U35271 ( .A(n34766), .B(n34765), .Z(n34898) );
  NAND U35272 ( .A(n34768), .B(n34767), .Z(n34772) );
  NANDN U35273 ( .A(n34770), .B(n34769), .Z(n34771) );
  NAND U35274 ( .A(n34772), .B(n34771), .Z(n34910) );
  OR U35275 ( .A(n34774), .B(n34773), .Z(n34778) );
  NAND U35276 ( .A(n34776), .B(n34775), .Z(n34777) );
  AND U35277 ( .A(n34778), .B(n34777), .Z(n34911) );
  XNOR U35278 ( .A(n34910), .B(n34911), .Z(n34912) );
  OR U35279 ( .A(n34780), .B(n34779), .Z(n34784) );
  NANDN U35280 ( .A(n34782), .B(n34781), .Z(n34783) );
  NAND U35281 ( .A(n34784), .B(n34783), .Z(n34978) );
  XOR U35282 ( .A(b[19]), .B(n36333), .Z(n34928) );
  NANDN U35283 ( .A(n34928), .B(n37934), .Z(n34787) );
  NANDN U35284 ( .A(n34785), .B(n37935), .Z(n34786) );
  NAND U35285 ( .A(n34787), .B(n34786), .Z(n35015) );
  XNOR U35286 ( .A(b[27]), .B(a[222]), .Z(n34931) );
  NANDN U35287 ( .A(n34931), .B(n38423), .Z(n34790) );
  NAND U35288 ( .A(n34788), .B(n38424), .Z(n34789) );
  NAND U35289 ( .A(n34790), .B(n34789), .Z(n35012) );
  XOR U35290 ( .A(a[244]), .B(n1051), .Z(n34934) );
  NANDN U35291 ( .A(n34934), .B(n36587), .Z(n34793) );
  NANDN U35292 ( .A(n34791), .B(n36588), .Z(n34792) );
  AND U35293 ( .A(n34793), .B(n34792), .Z(n35013) );
  XNOR U35294 ( .A(n35012), .B(n35013), .Z(n35014) );
  XNOR U35295 ( .A(n35015), .B(n35014), .Z(n34977) );
  NANDN U35296 ( .A(n34794), .B(n37762), .Z(n34796) );
  XNOR U35297 ( .A(b[17]), .B(a[232]), .Z(n34937) );
  NANDN U35298 ( .A(n34937), .B(n37764), .Z(n34795) );
  NAND U35299 ( .A(n34796), .B(n34795), .Z(n34955) );
  XNOR U35300 ( .A(b[31]), .B(a[218]), .Z(n34940) );
  NANDN U35301 ( .A(n34940), .B(n38552), .Z(n34799) );
  NANDN U35302 ( .A(n34797), .B(n38553), .Z(n34798) );
  NAND U35303 ( .A(n34799), .B(n34798), .Z(n34952) );
  OR U35304 ( .A(n34800), .B(n36105), .Z(n34802) );
  XOR U35305 ( .A(a[246]), .B(n1050), .Z(n34943) );
  NANDN U35306 ( .A(n34943), .B(n36107), .Z(n34801) );
  AND U35307 ( .A(n34802), .B(n34801), .Z(n34953) );
  XNOR U35308 ( .A(n34952), .B(n34953), .Z(n34954) );
  XOR U35309 ( .A(n34955), .B(n34954), .Z(n34976) );
  XOR U35310 ( .A(n34977), .B(n34976), .Z(n34979) );
  XNOR U35311 ( .A(n34978), .B(n34979), .Z(n35030) );
  XNOR U35312 ( .A(n35030), .B(n35031), .Z(n35032) );
  OR U35313 ( .A(n34812), .B(n34811), .Z(n34816) );
  OR U35314 ( .A(n34814), .B(n34813), .Z(n34815) );
  AND U35315 ( .A(n34816), .B(n34815), .Z(n35024) );
  OR U35316 ( .A(n34818), .B(n34817), .Z(n34822) );
  NANDN U35317 ( .A(n34820), .B(n34819), .Z(n34821) );
  NAND U35318 ( .A(n34822), .B(n34821), .Z(n35025) );
  XNOR U35319 ( .A(n35024), .B(n35025), .Z(n35026) );
  XOR U35320 ( .A(n35027), .B(n35026), .Z(n35033) );
  XOR U35321 ( .A(n35032), .B(n35033), .Z(n34918) );
  NANDN U35322 ( .A(n34828), .B(n34827), .Z(n34832) );
  NAND U35323 ( .A(n34830), .B(n34829), .Z(n34831) );
  NAND U35324 ( .A(n34832), .B(n34831), .Z(n35039) );
  OR U35325 ( .A(n34834), .B(n34833), .Z(n34838) );
  NAND U35326 ( .A(n34836), .B(n34835), .Z(n34837) );
  NAND U35327 ( .A(n34838), .B(n34837), .Z(n35036) );
  NANDN U35328 ( .A(n34840), .B(n34839), .Z(n34844) );
  NAND U35329 ( .A(n34842), .B(n34841), .Z(n34843) );
  NAND U35330 ( .A(n34844), .B(n34843), .Z(n34970) );
  NANDN U35331 ( .A(n34846), .B(n34845), .Z(n34850) );
  NAND U35332 ( .A(n34848), .B(n34847), .Z(n34849) );
  AND U35333 ( .A(n34850), .B(n34849), .Z(n34971) );
  XNOR U35334 ( .A(n34970), .B(n34971), .Z(n34972) );
  XOR U35335 ( .A(a[240]), .B(n1052), .Z(n34982) );
  NANDN U35336 ( .A(n34982), .B(n36925), .Z(n34853) );
  NANDN U35337 ( .A(n34851), .B(n36926), .Z(n34852) );
  NAND U35338 ( .A(n34853), .B(n34852), .Z(n34960) );
  XOR U35339 ( .A(b[15]), .B(n37080), .Z(n34985) );
  OR U35340 ( .A(n34985), .B(n37665), .Z(n34856) );
  NANDN U35341 ( .A(n34854), .B(n37604), .Z(n34855) );
  AND U35342 ( .A(n34856), .B(n34855), .Z(n34958) );
  XOR U35343 ( .A(b[21]), .B(n36592), .Z(n34988) );
  NANDN U35344 ( .A(n34988), .B(n38101), .Z(n34859) );
  NANDN U35345 ( .A(n34857), .B(n38102), .Z(n34858) );
  AND U35346 ( .A(n34859), .B(n34858), .Z(n34959) );
  XOR U35347 ( .A(n34960), .B(n34961), .Z(n34949) );
  XOR U35348 ( .A(n37467), .B(b[11]), .Z(n34991) );
  OR U35349 ( .A(n34991), .B(n37311), .Z(n34862) );
  NANDN U35350 ( .A(n34860), .B(n37218), .Z(n34861) );
  NAND U35351 ( .A(n34862), .B(n34861), .Z(n34947) );
  XOR U35352 ( .A(n1053), .B(a[236]), .Z(n34994) );
  NANDN U35353 ( .A(n34994), .B(n37424), .Z(n34865) );
  NAND U35354 ( .A(n37425), .B(n34863), .Z(n34864) );
  AND U35355 ( .A(n34865), .B(n34864), .Z(n34946) );
  XNOR U35356 ( .A(n34947), .B(n34946), .Z(n34948) );
  XOR U35357 ( .A(n34949), .B(n34948), .Z(n34966) );
  NANDN U35358 ( .A(n1049), .B(a[248]), .Z(n34866) );
  XNOR U35359 ( .A(b[1]), .B(n34866), .Z(n34868) );
  NANDN U35360 ( .A(b[0]), .B(a[247]), .Z(n34867) );
  AND U35361 ( .A(n34868), .B(n34867), .Z(n34924) );
  NAND U35362 ( .A(n34869), .B(n38490), .Z(n34871) );
  XNOR U35363 ( .A(n1058), .B(a[220]), .Z(n35000) );
  NANDN U35364 ( .A(n1048), .B(n35000), .Z(n34870) );
  NAND U35365 ( .A(n34871), .B(n34870), .Z(n34922) );
  NANDN U35366 ( .A(n1059), .B(a[216]), .Z(n34923) );
  XNOR U35367 ( .A(n34922), .B(n34923), .Z(n34925) );
  XOR U35368 ( .A(n34924), .B(n34925), .Z(n34964) );
  NANDN U35369 ( .A(n34872), .B(n38205), .Z(n34874) );
  XOR U35370 ( .A(b[23]), .B(n36280), .Z(n35003) );
  OR U35371 ( .A(n35003), .B(n38268), .Z(n34873) );
  NAND U35372 ( .A(n34874), .B(n34873), .Z(n35021) );
  XNOR U35373 ( .A(a[242]), .B(b[7]), .Z(n35006) );
  NANDN U35374 ( .A(n35006), .B(n36701), .Z(n34877) );
  NAND U35375 ( .A(n34875), .B(n36702), .Z(n34876) );
  NAND U35376 ( .A(n34877), .B(n34876), .Z(n35018) );
  XOR U35377 ( .A(b[25]), .B(a[224]), .Z(n35009) );
  NAND U35378 ( .A(n35009), .B(n38325), .Z(n34880) );
  NAND U35379 ( .A(n34878), .B(n38326), .Z(n34879) );
  AND U35380 ( .A(n34880), .B(n34879), .Z(n35019) );
  XNOR U35381 ( .A(n35018), .B(n35019), .Z(n35020) );
  XNOR U35382 ( .A(n35021), .B(n35020), .Z(n34965) );
  XOR U35383 ( .A(n34964), .B(n34965), .Z(n34967) );
  XNOR U35384 ( .A(n34966), .B(n34967), .Z(n34973) );
  XOR U35385 ( .A(n34972), .B(n34973), .Z(n35037) );
  XNOR U35386 ( .A(n35036), .B(n35037), .Z(n35038) );
  XNOR U35387 ( .A(n35039), .B(n35038), .Z(n34916) );
  XNOR U35388 ( .A(n34917), .B(n34916), .Z(n34919) );
  XNOR U35389 ( .A(n34918), .B(n34919), .Z(n34913) );
  XOR U35390 ( .A(n34912), .B(n34913), .Z(n34907) );
  NANDN U35391 ( .A(n34882), .B(n34881), .Z(n34886) );
  NAND U35392 ( .A(n34884), .B(n34883), .Z(n34885) );
  NAND U35393 ( .A(n34886), .B(n34885), .Z(n34904) );
  NANDN U35394 ( .A(n34888), .B(n34887), .Z(n34892) );
  NANDN U35395 ( .A(n34890), .B(n34889), .Z(n34891) );
  NAND U35396 ( .A(n34892), .B(n34891), .Z(n34905) );
  XNOR U35397 ( .A(n34904), .B(n34905), .Z(n34906) );
  XNOR U35398 ( .A(n34907), .B(n34906), .Z(n34899) );
  XNOR U35399 ( .A(n34898), .B(n34899), .Z(n34900) );
  XNOR U35400 ( .A(n34901), .B(n34900), .Z(n35042) );
  XNOR U35401 ( .A(n35042), .B(sreg[472]), .Z(n35044) );
  NAND U35402 ( .A(n34893), .B(sreg[471]), .Z(n34897) );
  OR U35403 ( .A(n34895), .B(n34894), .Z(n34896) );
  AND U35404 ( .A(n34897), .B(n34896), .Z(n35043) );
  XOR U35405 ( .A(n35044), .B(n35043), .Z(c[472]) );
  NANDN U35406 ( .A(n34899), .B(n34898), .Z(n34903) );
  NAND U35407 ( .A(n34901), .B(n34900), .Z(n34902) );
  NAND U35408 ( .A(n34903), .B(n34902), .Z(n35050) );
  NANDN U35409 ( .A(n34905), .B(n34904), .Z(n34909) );
  NAND U35410 ( .A(n34907), .B(n34906), .Z(n34908) );
  NAND U35411 ( .A(n34909), .B(n34908), .Z(n35048) );
  NANDN U35412 ( .A(n34911), .B(n34910), .Z(n34915) );
  NANDN U35413 ( .A(n34913), .B(n34912), .Z(n34914) );
  NAND U35414 ( .A(n34915), .B(n34914), .Z(n35054) );
  OR U35415 ( .A(n34917), .B(n34916), .Z(n34921) );
  OR U35416 ( .A(n34919), .B(n34918), .Z(n34920) );
  AND U35417 ( .A(n34921), .B(n34920), .Z(n35053) );
  XNOR U35418 ( .A(n35054), .B(n35053), .Z(n35055) );
  NANDN U35419 ( .A(n34923), .B(n34922), .Z(n34927) );
  NAND U35420 ( .A(n34925), .B(n34924), .Z(n34926) );
  NAND U35421 ( .A(n34927), .B(n34926), .Z(n35122) );
  XOR U35422 ( .A(b[19]), .B(n36934), .Z(n35089) );
  NANDN U35423 ( .A(n35089), .B(n37934), .Z(n34930) );
  NANDN U35424 ( .A(n34928), .B(n37935), .Z(n34929) );
  NAND U35425 ( .A(n34930), .B(n34929), .Z(n35158) );
  XOR U35426 ( .A(b[27]), .B(a[223]), .Z(n35092) );
  NAND U35427 ( .A(n38423), .B(n35092), .Z(n34933) );
  NANDN U35428 ( .A(n34931), .B(n38424), .Z(n34932) );
  NAND U35429 ( .A(n34933), .B(n34932), .Z(n35155) );
  XOR U35430 ( .A(a[245]), .B(n1051), .Z(n35095) );
  NANDN U35431 ( .A(n35095), .B(n36587), .Z(n34936) );
  NANDN U35432 ( .A(n34934), .B(n36588), .Z(n34935) );
  AND U35433 ( .A(n34936), .B(n34935), .Z(n35156) );
  XNOR U35434 ( .A(n35155), .B(n35156), .Z(n35157) );
  XNOR U35435 ( .A(n35158), .B(n35157), .Z(n35119) );
  NANDN U35436 ( .A(n34937), .B(n37762), .Z(n34939) );
  XNOR U35437 ( .A(b[17]), .B(a[233]), .Z(n35098) );
  NANDN U35438 ( .A(n35098), .B(n37764), .Z(n34938) );
  NAND U35439 ( .A(n34939), .B(n34938), .Z(n35073) );
  XNOR U35440 ( .A(b[31]), .B(a[219]), .Z(n35101) );
  NANDN U35441 ( .A(n35101), .B(n38552), .Z(n34942) );
  NANDN U35442 ( .A(n34940), .B(n38553), .Z(n34941) );
  AND U35443 ( .A(n34942), .B(n34941), .Z(n35071) );
  OR U35444 ( .A(n34943), .B(n36105), .Z(n34945) );
  XNOR U35445 ( .A(a[247]), .B(b[3]), .Z(n35104) );
  NANDN U35446 ( .A(n35104), .B(n36107), .Z(n34944) );
  AND U35447 ( .A(n34945), .B(n34944), .Z(n35072) );
  XOR U35448 ( .A(n35073), .B(n35074), .Z(n35120) );
  XOR U35449 ( .A(n35119), .B(n35120), .Z(n35121) );
  XNOR U35450 ( .A(n35122), .B(n35121), .Z(n35167) );
  NANDN U35451 ( .A(n34947), .B(n34946), .Z(n34951) );
  NAND U35452 ( .A(n34949), .B(n34948), .Z(n34950) );
  NAND U35453 ( .A(n34951), .B(n34950), .Z(n35110) );
  NANDN U35454 ( .A(n34953), .B(n34952), .Z(n34957) );
  NAND U35455 ( .A(n34955), .B(n34954), .Z(n34956) );
  NAND U35456 ( .A(n34957), .B(n34956), .Z(n35108) );
  OR U35457 ( .A(n34959), .B(n34958), .Z(n34963) );
  NANDN U35458 ( .A(n34961), .B(n34960), .Z(n34962) );
  NAND U35459 ( .A(n34963), .B(n34962), .Z(n35107) );
  XNOR U35460 ( .A(n35110), .B(n35109), .Z(n35168) );
  XNOR U35461 ( .A(n35167), .B(n35168), .Z(n35169) );
  NANDN U35462 ( .A(n34965), .B(n34964), .Z(n34969) );
  OR U35463 ( .A(n34967), .B(n34966), .Z(n34968) );
  AND U35464 ( .A(n34969), .B(n34968), .Z(n35170) );
  XNOR U35465 ( .A(n35169), .B(n35170), .Z(n35188) );
  NANDN U35466 ( .A(n34971), .B(n34970), .Z(n34975) );
  NANDN U35467 ( .A(n34973), .B(n34972), .Z(n34974) );
  NAND U35468 ( .A(n34975), .B(n34974), .Z(n35176) );
  NANDN U35469 ( .A(n34977), .B(n34976), .Z(n34981) );
  OR U35470 ( .A(n34979), .B(n34978), .Z(n34980) );
  NAND U35471 ( .A(n34981), .B(n34980), .Z(n35173) );
  XNOR U35472 ( .A(a[241]), .B(n1052), .Z(n35125) );
  NAND U35473 ( .A(n36925), .B(n35125), .Z(n34984) );
  NANDN U35474 ( .A(n34982), .B(n36926), .Z(n34983) );
  NAND U35475 ( .A(n34984), .B(n34983), .Z(n35079) );
  XOR U35476 ( .A(b[15]), .B(n37420), .Z(n35128) );
  OR U35477 ( .A(n35128), .B(n37665), .Z(n34987) );
  NANDN U35478 ( .A(n34985), .B(n37604), .Z(n34986) );
  AND U35479 ( .A(n34987), .B(n34986), .Z(n35077) );
  XNOR U35480 ( .A(n1056), .B(a[229]), .Z(n35131) );
  NAND U35481 ( .A(n35131), .B(n38101), .Z(n34990) );
  NANDN U35482 ( .A(n34988), .B(n38102), .Z(n34989) );
  AND U35483 ( .A(n34990), .B(n34989), .Z(n35078) );
  XOR U35484 ( .A(n35079), .B(n35080), .Z(n35068) );
  XNOR U35485 ( .A(a[239]), .B(b[11]), .Z(n35134) );
  OR U35486 ( .A(n35134), .B(n37311), .Z(n34993) );
  NANDN U35487 ( .A(n34991), .B(n37218), .Z(n34992) );
  NAND U35488 ( .A(n34993), .B(n34992), .Z(n35066) );
  XOR U35489 ( .A(n1053), .B(a[237]), .Z(n35137) );
  NANDN U35490 ( .A(n35137), .B(n37424), .Z(n34996) );
  NANDN U35491 ( .A(n34994), .B(n37425), .Z(n34995) );
  NAND U35492 ( .A(n34996), .B(n34995), .Z(n35065) );
  XOR U35493 ( .A(n35068), .B(n35067), .Z(n35062) );
  NANDN U35494 ( .A(n1049), .B(a[249]), .Z(n34997) );
  XNOR U35495 ( .A(b[1]), .B(n34997), .Z(n34999) );
  IV U35496 ( .A(a[248]), .Z(n38272) );
  NANDN U35497 ( .A(n38272), .B(n1049), .Z(n34998) );
  AND U35498 ( .A(n34999), .B(n34998), .Z(n35085) );
  NAND U35499 ( .A(n38490), .B(n35000), .Z(n35002) );
  XNOR U35500 ( .A(n1058), .B(a[221]), .Z(n35143) );
  NANDN U35501 ( .A(n1048), .B(n35143), .Z(n35001) );
  NAND U35502 ( .A(n35002), .B(n35001), .Z(n35083) );
  NANDN U35503 ( .A(n1059), .B(a[217]), .Z(n35084) );
  XNOR U35504 ( .A(n35083), .B(n35084), .Z(n35086) );
  XNOR U35505 ( .A(n35085), .B(n35086), .Z(n35060) );
  NANDN U35506 ( .A(n35003), .B(n38205), .Z(n35005) );
  XNOR U35507 ( .A(b[23]), .B(a[227]), .Z(n35146) );
  OR U35508 ( .A(n35146), .B(n38268), .Z(n35004) );
  NAND U35509 ( .A(n35005), .B(n35004), .Z(n35164) );
  XNOR U35510 ( .A(a[243]), .B(b[7]), .Z(n35149) );
  NANDN U35511 ( .A(n35149), .B(n36701), .Z(n35008) );
  NANDN U35512 ( .A(n35006), .B(n36702), .Z(n35007) );
  NAND U35513 ( .A(n35008), .B(n35007), .Z(n35161) );
  XNOR U35514 ( .A(b[25]), .B(a[225]), .Z(n35152) );
  NANDN U35515 ( .A(n35152), .B(n38325), .Z(n35011) );
  NAND U35516 ( .A(n35009), .B(n38326), .Z(n35010) );
  AND U35517 ( .A(n35011), .B(n35010), .Z(n35162) );
  XNOR U35518 ( .A(n35161), .B(n35162), .Z(n35163) );
  XOR U35519 ( .A(n35164), .B(n35163), .Z(n35059) );
  XNOR U35520 ( .A(n35062), .B(n35061), .Z(n35116) );
  NANDN U35521 ( .A(n35013), .B(n35012), .Z(n35017) );
  NAND U35522 ( .A(n35015), .B(n35014), .Z(n35016) );
  NAND U35523 ( .A(n35017), .B(n35016), .Z(n35114) );
  NANDN U35524 ( .A(n35019), .B(n35018), .Z(n35023) );
  NAND U35525 ( .A(n35021), .B(n35020), .Z(n35022) );
  AND U35526 ( .A(n35023), .B(n35022), .Z(n35113) );
  XNOR U35527 ( .A(n35114), .B(n35113), .Z(n35115) );
  XNOR U35528 ( .A(n35116), .B(n35115), .Z(n35174) );
  XNOR U35529 ( .A(n35173), .B(n35174), .Z(n35175) );
  XOR U35530 ( .A(n35176), .B(n35175), .Z(n35186) );
  OR U35531 ( .A(n35025), .B(n35024), .Z(n35029) );
  OR U35532 ( .A(n35027), .B(n35026), .Z(n35028) );
  AND U35533 ( .A(n35029), .B(n35028), .Z(n35185) );
  XNOR U35534 ( .A(n35186), .B(n35185), .Z(n35187) );
  XNOR U35535 ( .A(n35188), .B(n35187), .Z(n35182) );
  NANDN U35536 ( .A(n35031), .B(n35030), .Z(n35035) );
  NAND U35537 ( .A(n35033), .B(n35032), .Z(n35034) );
  NAND U35538 ( .A(n35035), .B(n35034), .Z(n35179) );
  NANDN U35539 ( .A(n35037), .B(n35036), .Z(n35041) );
  NAND U35540 ( .A(n35039), .B(n35038), .Z(n35040) );
  NAND U35541 ( .A(n35041), .B(n35040), .Z(n35180) );
  XNOR U35542 ( .A(n35179), .B(n35180), .Z(n35181) );
  XOR U35543 ( .A(n35182), .B(n35181), .Z(n35056) );
  XNOR U35544 ( .A(n35055), .B(n35056), .Z(n35047) );
  XOR U35545 ( .A(n35048), .B(n35047), .Z(n35049) );
  XNOR U35546 ( .A(n35050), .B(n35049), .Z(n35191) );
  XNOR U35547 ( .A(n35191), .B(sreg[473]), .Z(n35193) );
  NAND U35548 ( .A(n35042), .B(sreg[472]), .Z(n35046) );
  OR U35549 ( .A(n35044), .B(n35043), .Z(n35045) );
  AND U35550 ( .A(n35046), .B(n35045), .Z(n35192) );
  XOR U35551 ( .A(n35193), .B(n35192), .Z(c[473]) );
  NAND U35552 ( .A(n35048), .B(n35047), .Z(n35052) );
  NAND U35553 ( .A(n35050), .B(n35049), .Z(n35051) );
  NAND U35554 ( .A(n35052), .B(n35051), .Z(n35199) );
  NANDN U35555 ( .A(n35054), .B(n35053), .Z(n35058) );
  NANDN U35556 ( .A(n35056), .B(n35055), .Z(n35057) );
  NAND U35557 ( .A(n35058), .B(n35057), .Z(n35197) );
  NANDN U35558 ( .A(n35060), .B(n35059), .Z(n35064) );
  NANDN U35559 ( .A(n35062), .B(n35061), .Z(n35063) );
  NAND U35560 ( .A(n35064), .B(n35063), .Z(n35327) );
  OR U35561 ( .A(n35066), .B(n35065), .Z(n35070) );
  NAND U35562 ( .A(n35068), .B(n35067), .Z(n35069) );
  NAND U35563 ( .A(n35070), .B(n35069), .Z(n35266) );
  OR U35564 ( .A(n35072), .B(n35071), .Z(n35076) );
  NANDN U35565 ( .A(n35074), .B(n35073), .Z(n35075) );
  NAND U35566 ( .A(n35076), .B(n35075), .Z(n35265) );
  OR U35567 ( .A(n35078), .B(n35077), .Z(n35082) );
  NANDN U35568 ( .A(n35080), .B(n35079), .Z(n35081) );
  NAND U35569 ( .A(n35082), .B(n35081), .Z(n35264) );
  XOR U35570 ( .A(n35266), .B(n35267), .Z(n35324) );
  NANDN U35571 ( .A(n35084), .B(n35083), .Z(n35088) );
  NAND U35572 ( .A(n35086), .B(n35085), .Z(n35087) );
  NAND U35573 ( .A(n35088), .B(n35087), .Z(n35279) );
  XOR U35574 ( .A(b[19]), .B(n37079), .Z(n35224) );
  NANDN U35575 ( .A(n35224), .B(n37934), .Z(n35091) );
  NANDN U35576 ( .A(n35089), .B(n37935), .Z(n35090) );
  NAND U35577 ( .A(n35091), .B(n35090), .Z(n35291) );
  XOR U35578 ( .A(b[27]), .B(a[224]), .Z(n35227) );
  NAND U35579 ( .A(n38423), .B(n35227), .Z(n35094) );
  NAND U35580 ( .A(n35092), .B(n38424), .Z(n35093) );
  NAND U35581 ( .A(n35094), .B(n35093), .Z(n35288) );
  XOR U35582 ( .A(a[246]), .B(n1051), .Z(n35230) );
  NANDN U35583 ( .A(n35230), .B(n36587), .Z(n35097) );
  NANDN U35584 ( .A(n35095), .B(n36588), .Z(n35096) );
  AND U35585 ( .A(n35097), .B(n35096), .Z(n35289) );
  XNOR U35586 ( .A(n35288), .B(n35289), .Z(n35290) );
  XNOR U35587 ( .A(n35291), .B(n35290), .Z(n35277) );
  NANDN U35588 ( .A(n35098), .B(n37762), .Z(n35100) );
  XNOR U35589 ( .A(b[17]), .B(a[234]), .Z(n35233) );
  NANDN U35590 ( .A(n35233), .B(n37764), .Z(n35099) );
  NAND U35591 ( .A(n35100), .B(n35099), .Z(n35251) );
  XNOR U35592 ( .A(b[31]), .B(a[220]), .Z(n35236) );
  NANDN U35593 ( .A(n35236), .B(n38552), .Z(n35103) );
  NANDN U35594 ( .A(n35101), .B(n38553), .Z(n35102) );
  NAND U35595 ( .A(n35103), .B(n35102), .Z(n35248) );
  OR U35596 ( .A(n35104), .B(n36105), .Z(n35106) );
  XOR U35597 ( .A(a[248]), .B(n1050), .Z(n35239) );
  NANDN U35598 ( .A(n35239), .B(n36107), .Z(n35105) );
  AND U35599 ( .A(n35106), .B(n35105), .Z(n35249) );
  XNOR U35600 ( .A(n35248), .B(n35249), .Z(n35250) );
  XOR U35601 ( .A(n35251), .B(n35250), .Z(n35276) );
  XNOR U35602 ( .A(n35277), .B(n35276), .Z(n35278) );
  XNOR U35603 ( .A(n35279), .B(n35278), .Z(n35325) );
  XNOR U35604 ( .A(n35324), .B(n35325), .Z(n35326) );
  XNOR U35605 ( .A(n35327), .B(n35326), .Z(n35215) );
  OR U35606 ( .A(n35108), .B(n35107), .Z(n35112) );
  NAND U35607 ( .A(n35110), .B(n35109), .Z(n35111) );
  NAND U35608 ( .A(n35112), .B(n35111), .Z(n35213) );
  NANDN U35609 ( .A(n35114), .B(n35113), .Z(n35118) );
  NANDN U35610 ( .A(n35116), .B(n35115), .Z(n35117) );
  NAND U35611 ( .A(n35118), .B(n35117), .Z(n35333) );
  OR U35612 ( .A(n35120), .B(n35119), .Z(n35124) );
  NAND U35613 ( .A(n35122), .B(n35121), .Z(n35123) );
  NAND U35614 ( .A(n35124), .B(n35123), .Z(n35330) );
  XOR U35615 ( .A(n37676), .B(b[9]), .Z(n35294) );
  NANDN U35616 ( .A(n35294), .B(n36925), .Z(n35127) );
  NAND U35617 ( .A(n36926), .B(n35125), .Z(n35126) );
  NAND U35618 ( .A(n35127), .B(n35126), .Z(n35256) );
  XOR U35619 ( .A(b[15]), .B(n37106), .Z(n35297) );
  OR U35620 ( .A(n35297), .B(n37665), .Z(n35130) );
  NANDN U35621 ( .A(n35128), .B(n37604), .Z(n35129) );
  NAND U35622 ( .A(n35130), .B(n35129), .Z(n35254) );
  XOR U35623 ( .A(n1056), .B(a[230]), .Z(n35300) );
  NANDN U35624 ( .A(n35300), .B(n38101), .Z(n35133) );
  NAND U35625 ( .A(n38102), .B(n35131), .Z(n35132) );
  NAND U35626 ( .A(n35133), .B(n35132), .Z(n35255) );
  XNOR U35627 ( .A(n35254), .B(n35255), .Z(n35257) );
  XOR U35628 ( .A(n35256), .B(n35257), .Z(n35245) );
  XOR U35629 ( .A(n37668), .B(b[11]), .Z(n35303) );
  OR U35630 ( .A(n35303), .B(n37311), .Z(n35136) );
  NANDN U35631 ( .A(n35134), .B(n37218), .Z(n35135) );
  NAND U35632 ( .A(n35136), .B(n35135), .Z(n35243) );
  XOR U35633 ( .A(n1053), .B(a[238]), .Z(n35306) );
  NANDN U35634 ( .A(n35306), .B(n37424), .Z(n35139) );
  NANDN U35635 ( .A(n35137), .B(n37425), .Z(n35138) );
  AND U35636 ( .A(n35139), .B(n35138), .Z(n35242) );
  XNOR U35637 ( .A(n35243), .B(n35242), .Z(n35244) );
  XNOR U35638 ( .A(n35245), .B(n35244), .Z(n35261) );
  NANDN U35639 ( .A(n1049), .B(a[250]), .Z(n35140) );
  XNOR U35640 ( .A(b[1]), .B(n35140), .Z(n35142) );
  NANDN U35641 ( .A(b[0]), .B(a[249]), .Z(n35141) );
  AND U35642 ( .A(n35142), .B(n35141), .Z(n35220) );
  NAND U35643 ( .A(n38490), .B(n35143), .Z(n35145) );
  XOR U35644 ( .A(n1058), .B(n35381), .Z(n35309) );
  NANDN U35645 ( .A(n1048), .B(n35309), .Z(n35144) );
  NAND U35646 ( .A(n35145), .B(n35144), .Z(n35218) );
  NANDN U35647 ( .A(n1059), .B(a[218]), .Z(n35219) );
  XNOR U35648 ( .A(n35218), .B(n35219), .Z(n35221) );
  XNOR U35649 ( .A(n35220), .B(n35221), .Z(n35259) );
  NANDN U35650 ( .A(n35146), .B(n38205), .Z(n35148) );
  XOR U35651 ( .A(b[23]), .B(n36592), .Z(n35315) );
  OR U35652 ( .A(n35315), .B(n38268), .Z(n35147) );
  NAND U35653 ( .A(n35148), .B(n35147), .Z(n35285) );
  XNOR U35654 ( .A(a[244]), .B(b[7]), .Z(n35318) );
  NANDN U35655 ( .A(n35318), .B(n36701), .Z(n35151) );
  NANDN U35656 ( .A(n35149), .B(n36702), .Z(n35150) );
  NAND U35657 ( .A(n35151), .B(n35150), .Z(n35282) );
  XNOR U35658 ( .A(b[25]), .B(a[226]), .Z(n35321) );
  NANDN U35659 ( .A(n35321), .B(n38325), .Z(n35154) );
  NANDN U35660 ( .A(n35152), .B(n38326), .Z(n35153) );
  AND U35661 ( .A(n35154), .B(n35153), .Z(n35283) );
  XNOR U35662 ( .A(n35282), .B(n35283), .Z(n35284) );
  XOR U35663 ( .A(n35285), .B(n35284), .Z(n35258) );
  XOR U35664 ( .A(n35261), .B(n35260), .Z(n35273) );
  NANDN U35665 ( .A(n35156), .B(n35155), .Z(n35160) );
  NAND U35666 ( .A(n35158), .B(n35157), .Z(n35159) );
  NAND U35667 ( .A(n35160), .B(n35159), .Z(n35271) );
  NANDN U35668 ( .A(n35162), .B(n35161), .Z(n35166) );
  NAND U35669 ( .A(n35164), .B(n35163), .Z(n35165) );
  AND U35670 ( .A(n35166), .B(n35165), .Z(n35270) );
  XNOR U35671 ( .A(n35271), .B(n35270), .Z(n35272) );
  XNOR U35672 ( .A(n35273), .B(n35272), .Z(n35331) );
  XNOR U35673 ( .A(n35330), .B(n35331), .Z(n35332) );
  XNOR U35674 ( .A(n35333), .B(n35332), .Z(n35212) );
  XNOR U35675 ( .A(n35213), .B(n35212), .Z(n35214) );
  XOR U35676 ( .A(n35215), .B(n35214), .Z(n35209) );
  NANDN U35677 ( .A(n35168), .B(n35167), .Z(n35172) );
  NAND U35678 ( .A(n35170), .B(n35169), .Z(n35171) );
  NAND U35679 ( .A(n35172), .B(n35171), .Z(n35206) );
  NANDN U35680 ( .A(n35174), .B(n35173), .Z(n35178) );
  NAND U35681 ( .A(n35176), .B(n35175), .Z(n35177) );
  NAND U35682 ( .A(n35178), .B(n35177), .Z(n35207) );
  XNOR U35683 ( .A(n35206), .B(n35207), .Z(n35208) );
  XNOR U35684 ( .A(n35209), .B(n35208), .Z(n35203) );
  NANDN U35685 ( .A(n35180), .B(n35179), .Z(n35184) );
  NANDN U35686 ( .A(n35182), .B(n35181), .Z(n35183) );
  NAND U35687 ( .A(n35184), .B(n35183), .Z(n35200) );
  OR U35688 ( .A(n35186), .B(n35185), .Z(n35190) );
  OR U35689 ( .A(n35188), .B(n35187), .Z(n35189) );
  AND U35690 ( .A(n35190), .B(n35189), .Z(n35201) );
  XNOR U35691 ( .A(n35200), .B(n35201), .Z(n35202) );
  XNOR U35692 ( .A(n35203), .B(n35202), .Z(n35196) );
  XOR U35693 ( .A(n35197), .B(n35196), .Z(n35198) );
  XNOR U35694 ( .A(n35199), .B(n35198), .Z(n35336) );
  XNOR U35695 ( .A(n35336), .B(sreg[474]), .Z(n35338) );
  NAND U35696 ( .A(n35191), .B(sreg[473]), .Z(n35195) );
  OR U35697 ( .A(n35193), .B(n35192), .Z(n35194) );
  AND U35698 ( .A(n35195), .B(n35194), .Z(n35337) );
  XOR U35699 ( .A(n35338), .B(n35337), .Z(c[474]) );
  NANDN U35700 ( .A(n35201), .B(n35200), .Z(n35205) );
  NANDN U35701 ( .A(n35203), .B(n35202), .Z(n35204) );
  NAND U35702 ( .A(n35205), .B(n35204), .Z(n35342) );
  NANDN U35703 ( .A(n35207), .B(n35206), .Z(n35211) );
  NAND U35704 ( .A(n35209), .B(n35208), .Z(n35210) );
  NAND U35705 ( .A(n35211), .B(n35210), .Z(n35347) );
  NANDN U35706 ( .A(n35213), .B(n35212), .Z(n35217) );
  NANDN U35707 ( .A(n35215), .B(n35214), .Z(n35216) );
  NAND U35708 ( .A(n35217), .B(n35216), .Z(n35348) );
  XNOR U35709 ( .A(n35347), .B(n35348), .Z(n35349) );
  NANDN U35710 ( .A(n35219), .B(n35218), .Z(n35223) );
  NAND U35711 ( .A(n35221), .B(n35220), .Z(n35222) );
  NAND U35712 ( .A(n35223), .B(n35222), .Z(n35423) );
  XOR U35713 ( .A(b[19]), .B(n37184), .Z(n35375) );
  NANDN U35714 ( .A(n35375), .B(n37934), .Z(n35226) );
  NANDN U35715 ( .A(n35224), .B(n37935), .Z(n35225) );
  NAND U35716 ( .A(n35226), .B(n35225), .Z(n35463) );
  XNOR U35717 ( .A(b[27]), .B(a[225]), .Z(n35369) );
  NANDN U35718 ( .A(n35369), .B(n38423), .Z(n35229) );
  NAND U35719 ( .A(n35227), .B(n38424), .Z(n35228) );
  NAND U35720 ( .A(n35229), .B(n35228), .Z(n35460) );
  XNOR U35721 ( .A(a[247]), .B(b[5]), .Z(n35372) );
  NANDN U35722 ( .A(n35372), .B(n36587), .Z(n35232) );
  NANDN U35723 ( .A(n35230), .B(n36588), .Z(n35231) );
  AND U35724 ( .A(n35232), .B(n35231), .Z(n35461) );
  XNOR U35725 ( .A(n35460), .B(n35461), .Z(n35462) );
  XNOR U35726 ( .A(n35463), .B(n35462), .Z(n35421) );
  NANDN U35727 ( .A(n35233), .B(n37762), .Z(n35235) );
  XNOR U35728 ( .A(b[17]), .B(a[235]), .Z(n35378) );
  NANDN U35729 ( .A(n35378), .B(n37764), .Z(n35234) );
  NAND U35730 ( .A(n35235), .B(n35234), .Z(n35397) );
  XNOR U35731 ( .A(b[31]), .B(a[221]), .Z(n35382) );
  NANDN U35732 ( .A(n35382), .B(n38552), .Z(n35238) );
  NANDN U35733 ( .A(n35236), .B(n38553), .Z(n35237) );
  NAND U35734 ( .A(n35238), .B(n35237), .Z(n35394) );
  OR U35735 ( .A(n35239), .B(n36105), .Z(n35241) );
  XNOR U35736 ( .A(a[249]), .B(b[3]), .Z(n35385) );
  NANDN U35737 ( .A(n35385), .B(n36107), .Z(n35240) );
  AND U35738 ( .A(n35241), .B(n35240), .Z(n35395) );
  XNOR U35739 ( .A(n35394), .B(n35395), .Z(n35396) );
  XOR U35740 ( .A(n35397), .B(n35396), .Z(n35420) );
  XNOR U35741 ( .A(n35421), .B(n35420), .Z(n35422) );
  XNOR U35742 ( .A(n35423), .B(n35422), .Z(n35360) );
  NANDN U35743 ( .A(n35243), .B(n35242), .Z(n35247) );
  NAND U35744 ( .A(n35245), .B(n35244), .Z(n35246) );
  NAND U35745 ( .A(n35247), .B(n35246), .Z(n35412) );
  NANDN U35746 ( .A(n35249), .B(n35248), .Z(n35253) );
  NAND U35747 ( .A(n35251), .B(n35250), .Z(n35252) );
  NAND U35748 ( .A(n35253), .B(n35252), .Z(n35411) );
  XNOR U35749 ( .A(n35411), .B(n35410), .Z(n35413) );
  XOR U35750 ( .A(n35412), .B(n35413), .Z(n35359) );
  XOR U35751 ( .A(n35360), .B(n35359), .Z(n35361) );
  NANDN U35752 ( .A(n35259), .B(n35258), .Z(n35263) );
  NAND U35753 ( .A(n35261), .B(n35260), .Z(n35262) );
  NAND U35754 ( .A(n35263), .B(n35262), .Z(n35362) );
  XNOR U35755 ( .A(n35361), .B(n35362), .Z(n35474) );
  OR U35756 ( .A(n35265), .B(n35264), .Z(n35269) );
  NANDN U35757 ( .A(n35267), .B(n35266), .Z(n35268) );
  NAND U35758 ( .A(n35269), .B(n35268), .Z(n35473) );
  NANDN U35759 ( .A(n35271), .B(n35270), .Z(n35275) );
  NANDN U35760 ( .A(n35273), .B(n35272), .Z(n35274) );
  NAND U35761 ( .A(n35275), .B(n35274), .Z(n35356) );
  NANDN U35762 ( .A(n35277), .B(n35276), .Z(n35281) );
  NAND U35763 ( .A(n35279), .B(n35278), .Z(n35280) );
  NAND U35764 ( .A(n35281), .B(n35280), .Z(n35354) );
  NANDN U35765 ( .A(n35283), .B(n35282), .Z(n35287) );
  NAND U35766 ( .A(n35285), .B(n35284), .Z(n35286) );
  NAND U35767 ( .A(n35287), .B(n35286), .Z(n35414) );
  NANDN U35768 ( .A(n35289), .B(n35288), .Z(n35293) );
  NAND U35769 ( .A(n35291), .B(n35290), .Z(n35292) );
  AND U35770 ( .A(n35293), .B(n35292), .Z(n35415) );
  XNOR U35771 ( .A(n35414), .B(n35415), .Z(n35416) );
  XOR U35772 ( .A(a[243]), .B(n1052), .Z(n35424) );
  NANDN U35773 ( .A(n35424), .B(n36925), .Z(n35296) );
  NANDN U35774 ( .A(n35294), .B(n36926), .Z(n35295) );
  NAND U35775 ( .A(n35296), .B(n35295), .Z(n35402) );
  XNOR U35776 ( .A(n1054), .B(a[237]), .Z(n35427) );
  NANDN U35777 ( .A(n37665), .B(n35427), .Z(n35299) );
  NANDN U35778 ( .A(n35297), .B(n37604), .Z(n35298) );
  NAND U35779 ( .A(n35299), .B(n35298), .Z(n35400) );
  XOR U35780 ( .A(b[21]), .B(n36934), .Z(n35430) );
  NANDN U35781 ( .A(n35430), .B(n38101), .Z(n35302) );
  NANDN U35782 ( .A(n35300), .B(n38102), .Z(n35301) );
  NAND U35783 ( .A(n35302), .B(n35301), .Z(n35401) );
  XNOR U35784 ( .A(n35400), .B(n35401), .Z(n35403) );
  XOR U35785 ( .A(n35402), .B(n35403), .Z(n35391) );
  XNOR U35786 ( .A(a[241]), .B(b[11]), .Z(n35433) );
  OR U35787 ( .A(n35433), .B(n37311), .Z(n35305) );
  NANDN U35788 ( .A(n35303), .B(n37218), .Z(n35304) );
  NAND U35789 ( .A(n35305), .B(n35304), .Z(n35389) );
  XOR U35790 ( .A(n1053), .B(a[239]), .Z(n35436) );
  NANDN U35791 ( .A(n35436), .B(n37424), .Z(n35308) );
  NANDN U35792 ( .A(n35306), .B(n37425), .Z(n35307) );
  AND U35793 ( .A(n35308), .B(n35307), .Z(n35388) );
  XNOR U35794 ( .A(n35389), .B(n35388), .Z(n35390) );
  XNOR U35795 ( .A(n35391), .B(n35390), .Z(n35407) );
  NAND U35796 ( .A(n38490), .B(n35309), .Z(n35311) );
  XNOR U35797 ( .A(n1058), .B(a[223]), .Z(n35451) );
  NANDN U35798 ( .A(n1048), .B(n35451), .Z(n35310) );
  NAND U35799 ( .A(n35311), .B(n35310), .Z(n35363) );
  NANDN U35800 ( .A(n1059), .B(a[219]), .Z(n35364) );
  XNOR U35801 ( .A(n35363), .B(n35364), .Z(n35366) );
  NANDN U35802 ( .A(n1049), .B(a[251]), .Z(n35312) );
  XNOR U35803 ( .A(b[1]), .B(n35312), .Z(n35314) );
  IV U35804 ( .A(a[250]), .Z(n38356) );
  NANDN U35805 ( .A(n38356), .B(n1049), .Z(n35313) );
  AND U35806 ( .A(n35314), .B(n35313), .Z(n35365) );
  XNOR U35807 ( .A(n35366), .B(n35365), .Z(n35405) );
  NANDN U35808 ( .A(n35315), .B(n38205), .Z(n35317) );
  XNOR U35809 ( .A(b[23]), .B(a[229]), .Z(n35442) );
  OR U35810 ( .A(n35442), .B(n38268), .Z(n35316) );
  NAND U35811 ( .A(n35317), .B(n35316), .Z(n35457) );
  XNOR U35812 ( .A(a[245]), .B(b[7]), .Z(n35445) );
  NANDN U35813 ( .A(n35445), .B(n36701), .Z(n35320) );
  NANDN U35814 ( .A(n35318), .B(n36702), .Z(n35319) );
  NAND U35815 ( .A(n35320), .B(n35319), .Z(n35454) );
  XOR U35816 ( .A(b[25]), .B(a[227]), .Z(n35439) );
  NAND U35817 ( .A(n35439), .B(n38325), .Z(n35323) );
  NANDN U35818 ( .A(n35321), .B(n38326), .Z(n35322) );
  AND U35819 ( .A(n35323), .B(n35322), .Z(n35455) );
  XNOR U35820 ( .A(n35454), .B(n35455), .Z(n35456) );
  XOR U35821 ( .A(n35457), .B(n35456), .Z(n35404) );
  XOR U35822 ( .A(n35407), .B(n35406), .Z(n35417) );
  XOR U35823 ( .A(n35416), .B(n35417), .Z(n35353) );
  XOR U35824 ( .A(n35354), .B(n35353), .Z(n35355) );
  XNOR U35825 ( .A(n35356), .B(n35355), .Z(n35472) );
  XOR U35826 ( .A(n35473), .B(n35472), .Z(n35475) );
  NANDN U35827 ( .A(n35325), .B(n35324), .Z(n35329) );
  NAND U35828 ( .A(n35327), .B(n35326), .Z(n35328) );
  NAND U35829 ( .A(n35329), .B(n35328), .Z(n35467) );
  NANDN U35830 ( .A(n35331), .B(n35330), .Z(n35335) );
  NANDN U35831 ( .A(n35333), .B(n35332), .Z(n35334) );
  AND U35832 ( .A(n35335), .B(n35334), .Z(n35466) );
  XNOR U35833 ( .A(n35467), .B(n35466), .Z(n35468) );
  XOR U35834 ( .A(n35469), .B(n35468), .Z(n35350) );
  XOR U35835 ( .A(n35349), .B(n35350), .Z(n35341) );
  XOR U35836 ( .A(n35342), .B(n35341), .Z(n35343) );
  XNOR U35837 ( .A(n35344), .B(n35343), .Z(n35478) );
  XNOR U35838 ( .A(n35478), .B(sreg[475]), .Z(n35480) );
  NAND U35839 ( .A(n35336), .B(sreg[474]), .Z(n35340) );
  OR U35840 ( .A(n35338), .B(n35337), .Z(n35339) );
  AND U35841 ( .A(n35340), .B(n35339), .Z(n35479) );
  XOR U35842 ( .A(n35480), .B(n35479), .Z(c[475]) );
  NAND U35843 ( .A(n35342), .B(n35341), .Z(n35346) );
  NAND U35844 ( .A(n35344), .B(n35343), .Z(n35345) );
  NAND U35845 ( .A(n35346), .B(n35345), .Z(n35486) );
  NANDN U35846 ( .A(n35348), .B(n35347), .Z(n35352) );
  NAND U35847 ( .A(n35350), .B(n35349), .Z(n35351) );
  NAND U35848 ( .A(n35352), .B(n35351), .Z(n35483) );
  NAND U35849 ( .A(n35354), .B(n35353), .Z(n35358) );
  NANDN U35850 ( .A(n35356), .B(n35355), .Z(n35357) );
  NAND U35851 ( .A(n35358), .B(n35357), .Z(n35609) );
  XNOR U35852 ( .A(n35609), .B(n35610), .Z(n35611) );
  NANDN U35853 ( .A(n35364), .B(n35363), .Z(n35368) );
  NAND U35854 ( .A(n35366), .B(n35365), .Z(n35367) );
  NAND U35855 ( .A(n35368), .B(n35367), .Z(n35566) );
  XNOR U35856 ( .A(b[27]), .B(a[226]), .Z(n35520) );
  NANDN U35857 ( .A(n35520), .B(n38423), .Z(n35371) );
  NANDN U35858 ( .A(n35369), .B(n38424), .Z(n35370) );
  NAND U35859 ( .A(n35371), .B(n35370), .Z(n35570) );
  XOR U35860 ( .A(a[248]), .B(n1051), .Z(n35523) );
  NANDN U35861 ( .A(n35523), .B(n36587), .Z(n35374) );
  NANDN U35862 ( .A(n35372), .B(n36588), .Z(n35373) );
  NAND U35863 ( .A(n35374), .B(n35373), .Z(n35567) );
  XOR U35864 ( .A(b[19]), .B(n37080), .Z(n35526) );
  NANDN U35865 ( .A(n35526), .B(n37934), .Z(n35377) );
  NANDN U35866 ( .A(n35375), .B(n37935), .Z(n35376) );
  AND U35867 ( .A(n35377), .B(n35376), .Z(n35568) );
  XNOR U35868 ( .A(n35567), .B(n35568), .Z(n35569) );
  XNOR U35869 ( .A(n35570), .B(n35569), .Z(n35564) );
  NANDN U35870 ( .A(n35378), .B(n37762), .Z(n35380) );
  XNOR U35871 ( .A(b[17]), .B(a[236]), .Z(n35511) );
  NANDN U35872 ( .A(n35511), .B(n37764), .Z(n35379) );
  NAND U35873 ( .A(n35380), .B(n35379), .Z(n35544) );
  XOR U35874 ( .A(b[31]), .B(n35381), .Z(n35514) );
  NANDN U35875 ( .A(n35514), .B(n38552), .Z(n35384) );
  NANDN U35876 ( .A(n35382), .B(n38553), .Z(n35383) );
  NAND U35877 ( .A(n35384), .B(n35383), .Z(n35541) );
  OR U35878 ( .A(n35385), .B(n36105), .Z(n35387) );
  XOR U35879 ( .A(a[250]), .B(n1050), .Z(n35517) );
  NANDN U35880 ( .A(n35517), .B(n36107), .Z(n35386) );
  AND U35881 ( .A(n35387), .B(n35386), .Z(n35542) );
  XNOR U35882 ( .A(n35541), .B(n35542), .Z(n35543) );
  XOR U35883 ( .A(n35544), .B(n35543), .Z(n35563) );
  XNOR U35884 ( .A(n35564), .B(n35563), .Z(n35565) );
  XNOR U35885 ( .A(n35566), .B(n35565), .Z(n35502) );
  NANDN U35886 ( .A(n35389), .B(n35388), .Z(n35393) );
  NAND U35887 ( .A(n35391), .B(n35390), .Z(n35392) );
  NAND U35888 ( .A(n35393), .B(n35392), .Z(n35555) );
  NANDN U35889 ( .A(n35395), .B(n35394), .Z(n35399) );
  NAND U35890 ( .A(n35397), .B(n35396), .Z(n35398) );
  NAND U35891 ( .A(n35399), .B(n35398), .Z(n35554) );
  XNOR U35892 ( .A(n35554), .B(n35553), .Z(n35556) );
  XOR U35893 ( .A(n35555), .B(n35556), .Z(n35501) );
  XOR U35894 ( .A(n35502), .B(n35501), .Z(n35503) );
  NANDN U35895 ( .A(n35405), .B(n35404), .Z(n35409) );
  NAND U35896 ( .A(n35407), .B(n35406), .Z(n35408) );
  AND U35897 ( .A(n35409), .B(n35408), .Z(n35504) );
  XOR U35898 ( .A(n35503), .B(n35504), .Z(n35617) );
  NANDN U35899 ( .A(n35415), .B(n35414), .Z(n35419) );
  NAND U35900 ( .A(n35417), .B(n35416), .Z(n35418) );
  NAND U35901 ( .A(n35419), .B(n35418), .Z(n35498) );
  XOR U35902 ( .A(a[244]), .B(n1052), .Z(n35594) );
  NANDN U35903 ( .A(n35594), .B(n36925), .Z(n35426) );
  NANDN U35904 ( .A(n35424), .B(n36926), .Z(n35425) );
  NAND U35905 ( .A(n35426), .B(n35425), .Z(n35550) );
  XOR U35906 ( .A(b[15]), .B(n37467), .Z(n35597) );
  OR U35907 ( .A(n35597), .B(n37665), .Z(n35429) );
  NAND U35908 ( .A(n35427), .B(n37604), .Z(n35428) );
  NAND U35909 ( .A(n35429), .B(n35428), .Z(n35547) );
  XOR U35910 ( .A(b[21]), .B(n37079), .Z(n35600) );
  NANDN U35911 ( .A(n35600), .B(n38101), .Z(n35432) );
  NANDN U35912 ( .A(n35430), .B(n38102), .Z(n35431) );
  AND U35913 ( .A(n35432), .B(n35431), .Z(n35548) );
  XNOR U35914 ( .A(n35547), .B(n35548), .Z(n35549) );
  XNOR U35915 ( .A(n35550), .B(n35549), .Z(n35538) );
  XOR U35916 ( .A(n37676), .B(b[11]), .Z(n35606) );
  OR U35917 ( .A(n35606), .B(n37311), .Z(n35435) );
  NANDN U35918 ( .A(n35433), .B(n37218), .Z(n35434) );
  NAND U35919 ( .A(n35435), .B(n35434), .Z(n35536) );
  XOR U35920 ( .A(n37668), .B(b[13]), .Z(n35603) );
  NANDN U35921 ( .A(n35603), .B(n37424), .Z(n35438) );
  NANDN U35922 ( .A(n35436), .B(n37425), .Z(n35437) );
  AND U35923 ( .A(n35438), .B(n35437), .Z(n35535) );
  XNOR U35924 ( .A(n35536), .B(n35535), .Z(n35537) );
  XNOR U35925 ( .A(n35538), .B(n35537), .Z(n35508) );
  XNOR U35926 ( .A(b[25]), .B(a[228]), .Z(n35591) );
  NANDN U35927 ( .A(n35591), .B(n38325), .Z(n35441) );
  NAND U35928 ( .A(n35439), .B(n38326), .Z(n35440) );
  NAND U35929 ( .A(n35441), .B(n35440), .Z(n35576) );
  NANDN U35930 ( .A(n35442), .B(n38205), .Z(n35444) );
  XOR U35931 ( .A(b[23]), .B(n36333), .Z(n35585) );
  OR U35932 ( .A(n35585), .B(n38268), .Z(n35443) );
  NAND U35933 ( .A(n35444), .B(n35443), .Z(n35573) );
  XNOR U35934 ( .A(a[246]), .B(b[7]), .Z(n35588) );
  NANDN U35935 ( .A(n35588), .B(n36701), .Z(n35447) );
  NANDN U35936 ( .A(n35445), .B(n36702), .Z(n35446) );
  AND U35937 ( .A(n35447), .B(n35446), .Z(n35574) );
  XNOR U35938 ( .A(n35573), .B(n35574), .Z(n35575) );
  XNOR U35939 ( .A(n35576), .B(n35575), .Z(n35505) );
  NANDN U35940 ( .A(n1049), .B(a[252]), .Z(n35448) );
  XNOR U35941 ( .A(b[1]), .B(n35448), .Z(n35450) );
  NANDN U35942 ( .A(b[0]), .B(a[251]), .Z(n35449) );
  AND U35943 ( .A(n35450), .B(n35449), .Z(n35531) );
  NAND U35944 ( .A(n38490), .B(n35451), .Z(n35453) );
  XNOR U35945 ( .A(n1058), .B(a[224]), .Z(n35582) );
  NANDN U35946 ( .A(n1048), .B(n35582), .Z(n35452) );
  NAND U35947 ( .A(n35453), .B(n35452), .Z(n35529) );
  NANDN U35948 ( .A(n1059), .B(a[220]), .Z(n35530) );
  XNOR U35949 ( .A(n35529), .B(n35530), .Z(n35532) );
  XOR U35950 ( .A(n35531), .B(n35532), .Z(n35506) );
  XNOR U35951 ( .A(n35505), .B(n35506), .Z(n35507) );
  XOR U35952 ( .A(n35508), .B(n35507), .Z(n35560) );
  NANDN U35953 ( .A(n35455), .B(n35454), .Z(n35459) );
  NAND U35954 ( .A(n35457), .B(n35456), .Z(n35458) );
  NAND U35955 ( .A(n35459), .B(n35458), .Z(n35557) );
  NANDN U35956 ( .A(n35461), .B(n35460), .Z(n35465) );
  NAND U35957 ( .A(n35463), .B(n35462), .Z(n35464) );
  AND U35958 ( .A(n35465), .B(n35464), .Z(n35558) );
  XNOR U35959 ( .A(n35557), .B(n35558), .Z(n35559) );
  XNOR U35960 ( .A(n35560), .B(n35559), .Z(n35496) );
  XNOR U35961 ( .A(n35495), .B(n35496), .Z(n35497) );
  XNOR U35962 ( .A(n35498), .B(n35497), .Z(n35615) );
  XNOR U35963 ( .A(n35616), .B(n35615), .Z(n35618) );
  XNOR U35964 ( .A(n35617), .B(n35618), .Z(n35612) );
  XOR U35965 ( .A(n35611), .B(n35612), .Z(n35492) );
  NANDN U35966 ( .A(n35467), .B(n35466), .Z(n35471) );
  NAND U35967 ( .A(n35469), .B(n35468), .Z(n35470) );
  NAND U35968 ( .A(n35471), .B(n35470), .Z(n35489) );
  NANDN U35969 ( .A(n35473), .B(n35472), .Z(n35477) );
  OR U35970 ( .A(n35475), .B(n35474), .Z(n35476) );
  NAND U35971 ( .A(n35477), .B(n35476), .Z(n35490) );
  XNOR U35972 ( .A(n35489), .B(n35490), .Z(n35491) );
  XNOR U35973 ( .A(n35492), .B(n35491), .Z(n35484) );
  XNOR U35974 ( .A(n35483), .B(n35484), .Z(n35485) );
  XNOR U35975 ( .A(n35486), .B(n35485), .Z(n35621) );
  XNOR U35976 ( .A(n35621), .B(sreg[476]), .Z(n35623) );
  NAND U35977 ( .A(n35478), .B(sreg[475]), .Z(n35482) );
  OR U35978 ( .A(n35480), .B(n35479), .Z(n35481) );
  AND U35979 ( .A(n35482), .B(n35481), .Z(n35622) );
  XOR U35980 ( .A(n35623), .B(n35622), .Z(c[476]) );
  NANDN U35981 ( .A(n35484), .B(n35483), .Z(n35488) );
  NAND U35982 ( .A(n35486), .B(n35485), .Z(n35487) );
  NAND U35983 ( .A(n35488), .B(n35487), .Z(n35629) );
  NANDN U35984 ( .A(n35490), .B(n35489), .Z(n35494) );
  NAND U35985 ( .A(n35492), .B(n35491), .Z(n35493) );
  NAND U35986 ( .A(n35494), .B(n35493), .Z(n35626) );
  NANDN U35987 ( .A(n35496), .B(n35495), .Z(n35500) );
  NAND U35988 ( .A(n35498), .B(n35497), .Z(n35499) );
  NAND U35989 ( .A(n35500), .B(n35499), .Z(n35758) );
  XNOR U35990 ( .A(n35758), .B(n35759), .Z(n35760) );
  NANDN U35991 ( .A(n35506), .B(n35505), .Z(n35510) );
  NANDN U35992 ( .A(n35508), .B(n35507), .Z(n35509) );
  NAND U35993 ( .A(n35510), .B(n35509), .Z(n35647) );
  NANDN U35994 ( .A(n35511), .B(n37762), .Z(n35513) );
  XOR U35995 ( .A(b[17]), .B(a[237]), .Z(n35656) );
  NAND U35996 ( .A(n35656), .B(n37764), .Z(n35512) );
  NAND U35997 ( .A(n35513), .B(n35512), .Z(n35689) );
  XNOR U35998 ( .A(b[31]), .B(a[223]), .Z(n35659) );
  NANDN U35999 ( .A(n35659), .B(n38552), .Z(n35516) );
  NANDN U36000 ( .A(n35514), .B(n38553), .Z(n35515) );
  NAND U36001 ( .A(n35516), .B(n35515), .Z(n35686) );
  OR U36002 ( .A(n35517), .B(n36105), .Z(n35519) );
  XNOR U36003 ( .A(a[251]), .B(b[3]), .Z(n35662) );
  NANDN U36004 ( .A(n35662), .B(n36107), .Z(n35518) );
  AND U36005 ( .A(n35519), .B(n35518), .Z(n35687) );
  XNOR U36006 ( .A(n35686), .B(n35687), .Z(n35688) );
  XNOR U36007 ( .A(n35689), .B(n35688), .Z(n35710) );
  XOR U36008 ( .A(b[27]), .B(a[227]), .Z(n35665) );
  NAND U36009 ( .A(n38423), .B(n35665), .Z(n35522) );
  NANDN U36010 ( .A(n35520), .B(n38424), .Z(n35521) );
  NAND U36011 ( .A(n35522), .B(n35521), .Z(n35755) );
  XNOR U36012 ( .A(a[249]), .B(b[5]), .Z(n35668) );
  NANDN U36013 ( .A(n35668), .B(n36587), .Z(n35525) );
  NANDN U36014 ( .A(n35523), .B(n36588), .Z(n35524) );
  NAND U36015 ( .A(n35525), .B(n35524), .Z(n35752) );
  XOR U36016 ( .A(b[19]), .B(n37420), .Z(n35671) );
  NANDN U36017 ( .A(n35671), .B(n37934), .Z(n35528) );
  NANDN U36018 ( .A(n35526), .B(n37935), .Z(n35527) );
  AND U36019 ( .A(n35528), .B(n35527), .Z(n35753) );
  XNOR U36020 ( .A(n35752), .B(n35753), .Z(n35754) );
  XOR U36021 ( .A(n35755), .B(n35754), .Z(n35711) );
  XNOR U36022 ( .A(n35710), .B(n35711), .Z(n35712) );
  NANDN U36023 ( .A(n35530), .B(n35529), .Z(n35534) );
  NAND U36024 ( .A(n35532), .B(n35531), .Z(n35533) );
  AND U36025 ( .A(n35534), .B(n35533), .Z(n35713) );
  XNOR U36026 ( .A(n35712), .B(n35713), .Z(n35645) );
  NANDN U36027 ( .A(n35536), .B(n35535), .Z(n35540) );
  NAND U36028 ( .A(n35538), .B(n35537), .Z(n35539) );
  NAND U36029 ( .A(n35540), .B(n35539), .Z(n35701) );
  NANDN U36030 ( .A(n35542), .B(n35541), .Z(n35546) );
  NAND U36031 ( .A(n35544), .B(n35543), .Z(n35545) );
  NAND U36032 ( .A(n35546), .B(n35545), .Z(n35699) );
  NANDN U36033 ( .A(n35548), .B(n35547), .Z(n35552) );
  NAND U36034 ( .A(n35550), .B(n35549), .Z(n35551) );
  AND U36035 ( .A(n35552), .B(n35551), .Z(n35698) );
  XNOR U36036 ( .A(n35699), .B(n35698), .Z(n35700) );
  XOR U36037 ( .A(n35701), .B(n35700), .Z(n35644) );
  XNOR U36038 ( .A(n35645), .B(n35644), .Z(n35646) );
  XOR U36039 ( .A(n35647), .B(n35646), .Z(n35766) );
  NANDN U36040 ( .A(n35558), .B(n35557), .Z(n35562) );
  NAND U36041 ( .A(n35560), .B(n35559), .Z(n35561) );
  NAND U36042 ( .A(n35562), .B(n35561), .Z(n35641) );
  NANDN U36043 ( .A(n35568), .B(n35567), .Z(n35572) );
  NAND U36044 ( .A(n35570), .B(n35569), .Z(n35571) );
  NAND U36045 ( .A(n35572), .B(n35571), .Z(n35705) );
  NANDN U36046 ( .A(n35574), .B(n35573), .Z(n35578) );
  NAND U36047 ( .A(n35576), .B(n35575), .Z(n35577) );
  AND U36048 ( .A(n35578), .B(n35577), .Z(n35704) );
  XNOR U36049 ( .A(n35705), .B(n35704), .Z(n35706) );
  NANDN U36050 ( .A(n1049), .B(a[253]), .Z(n35579) );
  XNOR U36051 ( .A(b[1]), .B(n35579), .Z(n35581) );
  IV U36052 ( .A(a[252]), .Z(n38531) );
  NANDN U36053 ( .A(n38531), .B(n1049), .Z(n35580) );
  AND U36054 ( .A(n35581), .B(n35580), .Z(n35676) );
  NAND U36055 ( .A(n38490), .B(n35582), .Z(n35584) );
  XOR U36056 ( .A(b[29]), .B(n36167), .Z(n35743) );
  OR U36057 ( .A(n35743), .B(n1048), .Z(n35583) );
  NAND U36058 ( .A(n35584), .B(n35583), .Z(n35674) );
  NANDN U36059 ( .A(n1059), .B(a[221]), .Z(n35675) );
  XNOR U36060 ( .A(n35674), .B(n35675), .Z(n35677) );
  XOR U36061 ( .A(n35676), .B(n35677), .Z(n35653) );
  NANDN U36062 ( .A(n35585), .B(n38205), .Z(n35587) );
  XOR U36063 ( .A(b[23]), .B(n36934), .Z(n35734) );
  OR U36064 ( .A(n35734), .B(n38268), .Z(n35586) );
  NAND U36065 ( .A(n35587), .B(n35586), .Z(n35749) );
  XOR U36066 ( .A(a[247]), .B(b[7]), .Z(n35737) );
  NAND U36067 ( .A(n35737), .B(n36701), .Z(n35590) );
  NANDN U36068 ( .A(n35588), .B(n36702), .Z(n35589) );
  NAND U36069 ( .A(n35590), .B(n35589), .Z(n35746) );
  XOR U36070 ( .A(b[25]), .B(a[229]), .Z(n35731) );
  NAND U36071 ( .A(n35731), .B(n38325), .Z(n35593) );
  NANDN U36072 ( .A(n35591), .B(n38326), .Z(n35592) );
  AND U36073 ( .A(n35593), .B(n35592), .Z(n35747) );
  XNOR U36074 ( .A(n35746), .B(n35747), .Z(n35748) );
  XNOR U36075 ( .A(n35749), .B(n35748), .Z(n35650) );
  XOR U36076 ( .A(a[245]), .B(n1052), .Z(n35728) );
  NANDN U36077 ( .A(n35728), .B(n36925), .Z(n35596) );
  NANDN U36078 ( .A(n35594), .B(n36926), .Z(n35595) );
  NAND U36079 ( .A(n35596), .B(n35595), .Z(n35695) );
  XNOR U36080 ( .A(b[15]), .B(a[239]), .Z(n35722) );
  OR U36081 ( .A(n35722), .B(n37665), .Z(n35599) );
  NANDN U36082 ( .A(n35597), .B(n37604), .Z(n35598) );
  NAND U36083 ( .A(n35599), .B(n35598), .Z(n35692) );
  XOR U36084 ( .A(b[21]), .B(n37184), .Z(n35725) );
  NANDN U36085 ( .A(n35725), .B(n38101), .Z(n35602) );
  NANDN U36086 ( .A(n35600), .B(n38102), .Z(n35601) );
  AND U36087 ( .A(n35602), .B(n35601), .Z(n35693) );
  XNOR U36088 ( .A(n35692), .B(n35693), .Z(n35694) );
  XNOR U36089 ( .A(n35695), .B(n35694), .Z(n35683) );
  XNOR U36090 ( .A(a[241]), .B(b[13]), .Z(n35719) );
  NANDN U36091 ( .A(n35719), .B(n37424), .Z(n35605) );
  NANDN U36092 ( .A(n35603), .B(n37425), .Z(n35604) );
  NAND U36093 ( .A(n35605), .B(n35604), .Z(n35681) );
  XNOR U36094 ( .A(a[243]), .B(b[11]), .Z(n35716) );
  OR U36095 ( .A(n35716), .B(n37311), .Z(n35608) );
  NANDN U36096 ( .A(n35606), .B(n37218), .Z(n35607) );
  AND U36097 ( .A(n35608), .B(n35607), .Z(n35680) );
  XNOR U36098 ( .A(n35681), .B(n35680), .Z(n35682) );
  XNOR U36099 ( .A(n35683), .B(n35682), .Z(n35651) );
  XOR U36100 ( .A(n35653), .B(n35652), .Z(n35707) );
  XNOR U36101 ( .A(n35706), .B(n35707), .Z(n35639) );
  XNOR U36102 ( .A(n35638), .B(n35639), .Z(n35640) );
  XNOR U36103 ( .A(n35641), .B(n35640), .Z(n35764) );
  XNOR U36104 ( .A(n35765), .B(n35764), .Z(n35767) );
  XNOR U36105 ( .A(n35766), .B(n35767), .Z(n35761) );
  XOR U36106 ( .A(n35760), .B(n35761), .Z(n35635) );
  NANDN U36107 ( .A(n35610), .B(n35609), .Z(n35614) );
  NANDN U36108 ( .A(n35612), .B(n35611), .Z(n35613) );
  NAND U36109 ( .A(n35614), .B(n35613), .Z(n35633) );
  OR U36110 ( .A(n35616), .B(n35615), .Z(n35620) );
  OR U36111 ( .A(n35618), .B(n35617), .Z(n35619) );
  AND U36112 ( .A(n35620), .B(n35619), .Z(n35632) );
  XNOR U36113 ( .A(n35633), .B(n35632), .Z(n35634) );
  XNOR U36114 ( .A(n35635), .B(n35634), .Z(n35627) );
  XNOR U36115 ( .A(n35626), .B(n35627), .Z(n35628) );
  XNOR U36116 ( .A(n35629), .B(n35628), .Z(n35770) );
  XNOR U36117 ( .A(n35770), .B(sreg[477]), .Z(n35772) );
  NAND U36118 ( .A(n35621), .B(sreg[476]), .Z(n35625) );
  OR U36119 ( .A(n35623), .B(n35622), .Z(n35624) );
  AND U36120 ( .A(n35625), .B(n35624), .Z(n35771) );
  XOR U36121 ( .A(n35772), .B(n35771), .Z(c[477]) );
  NANDN U36122 ( .A(n35627), .B(n35626), .Z(n35631) );
  NAND U36123 ( .A(n35629), .B(n35628), .Z(n35630) );
  NAND U36124 ( .A(n35631), .B(n35630), .Z(n35778) );
  NANDN U36125 ( .A(n35633), .B(n35632), .Z(n35637) );
  NAND U36126 ( .A(n35635), .B(n35634), .Z(n35636) );
  NAND U36127 ( .A(n35637), .B(n35636), .Z(n35775) );
  NANDN U36128 ( .A(n35639), .B(n35638), .Z(n35643) );
  NAND U36129 ( .A(n35641), .B(n35640), .Z(n35642) );
  NAND U36130 ( .A(n35643), .B(n35642), .Z(n35791) );
  NANDN U36131 ( .A(n35645), .B(n35644), .Z(n35649) );
  NAND U36132 ( .A(n35647), .B(n35646), .Z(n35648) );
  NAND U36133 ( .A(n35649), .B(n35648), .Z(n35792) );
  XNOR U36134 ( .A(n35791), .B(n35792), .Z(n35793) );
  NANDN U36135 ( .A(n35651), .B(n35650), .Z(n35655) );
  NANDN U36136 ( .A(n35653), .B(n35652), .Z(n35654) );
  NAND U36137 ( .A(n35655), .B(n35654), .Z(n35914) );
  NAND U36138 ( .A(n35656), .B(n37762), .Z(n35658) );
  XNOR U36139 ( .A(b[17]), .B(a[238]), .Z(n35872) );
  NANDN U36140 ( .A(n35872), .B(n37764), .Z(n35657) );
  NAND U36141 ( .A(n35658), .B(n35657), .Z(n35896) );
  XNOR U36142 ( .A(b[31]), .B(a[224]), .Z(n35875) );
  NANDN U36143 ( .A(n35875), .B(n38552), .Z(n35661) );
  NANDN U36144 ( .A(n35659), .B(n38553), .Z(n35660) );
  NAND U36145 ( .A(n35661), .B(n35660), .Z(n35893) );
  OR U36146 ( .A(n35662), .B(n36105), .Z(n35664) );
  XOR U36147 ( .A(a[252]), .B(n1050), .Z(n35878) );
  NANDN U36148 ( .A(n35878), .B(n36107), .Z(n35663) );
  AND U36149 ( .A(n35664), .B(n35663), .Z(n35894) );
  XNOR U36150 ( .A(n35893), .B(n35894), .Z(n35895) );
  XNOR U36151 ( .A(n35896), .B(n35895), .Z(n35803) );
  XNOR U36152 ( .A(b[27]), .B(a[228]), .Z(n35863) );
  NANDN U36153 ( .A(n35863), .B(n38423), .Z(n35667) );
  NAND U36154 ( .A(n35665), .B(n38424), .Z(n35666) );
  NAND U36155 ( .A(n35667), .B(n35666), .Z(n35848) );
  XOR U36156 ( .A(a[250]), .B(n1051), .Z(n35866) );
  NANDN U36157 ( .A(n35866), .B(n36587), .Z(n35670) );
  NANDN U36158 ( .A(n35668), .B(n36588), .Z(n35669) );
  NAND U36159 ( .A(n35670), .B(n35669), .Z(n35845) );
  XOR U36160 ( .A(b[19]), .B(n37106), .Z(n35869) );
  NANDN U36161 ( .A(n35869), .B(n37934), .Z(n35673) );
  NANDN U36162 ( .A(n35671), .B(n37935), .Z(n35672) );
  AND U36163 ( .A(n35673), .B(n35672), .Z(n35846) );
  XNOR U36164 ( .A(n35845), .B(n35846), .Z(n35847) );
  XOR U36165 ( .A(n35848), .B(n35847), .Z(n35804) );
  XNOR U36166 ( .A(n35803), .B(n35804), .Z(n35805) );
  NANDN U36167 ( .A(n35675), .B(n35674), .Z(n35679) );
  NAND U36168 ( .A(n35677), .B(n35676), .Z(n35678) );
  AND U36169 ( .A(n35679), .B(n35678), .Z(n35806) );
  XNOR U36170 ( .A(n35805), .B(n35806), .Z(n35912) );
  NANDN U36171 ( .A(n35681), .B(n35680), .Z(n35685) );
  NAND U36172 ( .A(n35683), .B(n35682), .Z(n35684) );
  NAND U36173 ( .A(n35685), .B(n35684), .Z(n35854) );
  NANDN U36174 ( .A(n35687), .B(n35686), .Z(n35691) );
  NAND U36175 ( .A(n35689), .B(n35688), .Z(n35690) );
  NAND U36176 ( .A(n35691), .B(n35690), .Z(n35852) );
  NANDN U36177 ( .A(n35693), .B(n35692), .Z(n35697) );
  NAND U36178 ( .A(n35695), .B(n35694), .Z(n35696) );
  AND U36179 ( .A(n35697), .B(n35696), .Z(n35851) );
  XNOR U36180 ( .A(n35852), .B(n35851), .Z(n35853) );
  XOR U36181 ( .A(n35854), .B(n35853), .Z(n35911) );
  XNOR U36182 ( .A(n35912), .B(n35911), .Z(n35913) );
  XNOR U36183 ( .A(n35914), .B(n35913), .Z(n35790) );
  NANDN U36184 ( .A(n35699), .B(n35698), .Z(n35703) );
  NAND U36185 ( .A(n35701), .B(n35700), .Z(n35702) );
  NAND U36186 ( .A(n35703), .B(n35702), .Z(n35788) );
  NANDN U36187 ( .A(n35705), .B(n35704), .Z(n35709) );
  NANDN U36188 ( .A(n35707), .B(n35706), .Z(n35708) );
  NAND U36189 ( .A(n35709), .B(n35708), .Z(n35906) );
  NANDN U36190 ( .A(n35711), .B(n35710), .Z(n35715) );
  NAND U36191 ( .A(n35713), .B(n35712), .Z(n35714) );
  AND U36192 ( .A(n35715), .B(n35714), .Z(n35905) );
  XNOR U36193 ( .A(n35906), .B(n35905), .Z(n35907) );
  XNOR U36194 ( .A(n38034), .B(b[11]), .Z(n35836) );
  NANDN U36195 ( .A(n37311), .B(n35836), .Z(n35718) );
  NANDN U36196 ( .A(n35716), .B(n37218), .Z(n35717) );
  NAND U36197 ( .A(n35718), .B(n35717), .Z(n35902) );
  XOR U36198 ( .A(n37676), .B(n1053), .Z(n35833) );
  NAND U36199 ( .A(n35833), .B(n37424), .Z(n35721) );
  NANDN U36200 ( .A(n35719), .B(n37425), .Z(n35720) );
  NAND U36201 ( .A(n35721), .B(n35720), .Z(n35899) );
  XOR U36202 ( .A(b[15]), .B(n37668), .Z(n35824) );
  OR U36203 ( .A(n35824), .B(n37665), .Z(n35724) );
  NANDN U36204 ( .A(n35722), .B(n37604), .Z(n35723) );
  NAND U36205 ( .A(n35724), .B(n35723), .Z(n35890) );
  XOR U36206 ( .A(b[21]), .B(n37080), .Z(n35827) );
  NANDN U36207 ( .A(n35827), .B(n38101), .Z(n35727) );
  NANDN U36208 ( .A(n35725), .B(n38102), .Z(n35726) );
  NAND U36209 ( .A(n35727), .B(n35726), .Z(n35887) );
  XOR U36210 ( .A(a[246]), .B(n1052), .Z(n35830) );
  NANDN U36211 ( .A(n35830), .B(n36925), .Z(n35730) );
  NANDN U36212 ( .A(n35728), .B(n36926), .Z(n35729) );
  AND U36213 ( .A(n35730), .B(n35729), .Z(n35888) );
  XNOR U36214 ( .A(n35887), .B(n35888), .Z(n35889) );
  XNOR U36215 ( .A(n35890), .B(n35889), .Z(n35900) );
  XNOR U36216 ( .A(n35899), .B(n35900), .Z(n35901) );
  XNOR U36217 ( .A(n35902), .B(n35901), .Z(n35859) );
  XNOR U36218 ( .A(b[25]), .B(a[230]), .Z(n35809) );
  NANDN U36219 ( .A(n35809), .B(n38325), .Z(n35733) );
  NAND U36220 ( .A(n35731), .B(n38326), .Z(n35732) );
  NAND U36221 ( .A(n35733), .B(n35732), .Z(n35842) );
  NANDN U36222 ( .A(n35734), .B(n38205), .Z(n35736) );
  XOR U36223 ( .A(b[23]), .B(n37079), .Z(n35812) );
  OR U36224 ( .A(n35812), .B(n38268), .Z(n35735) );
  NAND U36225 ( .A(n35736), .B(n35735), .Z(n35839) );
  XNOR U36226 ( .A(a[248]), .B(b[7]), .Z(n35815) );
  NANDN U36227 ( .A(n35815), .B(n36701), .Z(n35739) );
  NAND U36228 ( .A(n35737), .B(n36702), .Z(n35738) );
  AND U36229 ( .A(n35739), .B(n35738), .Z(n35840) );
  XNOR U36230 ( .A(n35839), .B(n35840), .Z(n35841) );
  XNOR U36231 ( .A(n35842), .B(n35841), .Z(n35857) );
  NAND U36232 ( .A(a[222]), .B(b[31]), .Z(n35884) );
  NANDN U36233 ( .A(n1049), .B(a[254]), .Z(n35740) );
  XNOR U36234 ( .A(b[1]), .B(n35740), .Z(n35742) );
  NANDN U36235 ( .A(b[0]), .B(a[253]), .Z(n35741) );
  AND U36236 ( .A(n35742), .B(n35741), .Z(n35882) );
  NANDN U36237 ( .A(n35743), .B(n38490), .Z(n35745) );
  XNOR U36238 ( .A(n1058), .B(a[226]), .Z(n35821) );
  NANDN U36239 ( .A(n1048), .B(n35821), .Z(n35744) );
  AND U36240 ( .A(n35745), .B(n35744), .Z(n35881) );
  XNOR U36241 ( .A(n35882), .B(n35881), .Z(n35883) );
  XNOR U36242 ( .A(n35884), .B(n35883), .Z(n35858) );
  XOR U36243 ( .A(n35857), .B(n35858), .Z(n35860) );
  XNOR U36244 ( .A(n35859), .B(n35860), .Z(n35800) );
  NANDN U36245 ( .A(n35747), .B(n35746), .Z(n35751) );
  NAND U36246 ( .A(n35749), .B(n35748), .Z(n35750) );
  NAND U36247 ( .A(n35751), .B(n35750), .Z(n35797) );
  NANDN U36248 ( .A(n35753), .B(n35752), .Z(n35757) );
  NAND U36249 ( .A(n35755), .B(n35754), .Z(n35756) );
  AND U36250 ( .A(n35757), .B(n35756), .Z(n35798) );
  XNOR U36251 ( .A(n35797), .B(n35798), .Z(n35799) );
  XOR U36252 ( .A(n35800), .B(n35799), .Z(n35908) );
  XNOR U36253 ( .A(n35907), .B(n35908), .Z(n35787) );
  XNOR U36254 ( .A(n35788), .B(n35787), .Z(n35789) );
  XOR U36255 ( .A(n35790), .B(n35789), .Z(n35794) );
  XNOR U36256 ( .A(n35793), .B(n35794), .Z(n35784) );
  NANDN U36257 ( .A(n35759), .B(n35758), .Z(n35763) );
  NANDN U36258 ( .A(n35761), .B(n35760), .Z(n35762) );
  NAND U36259 ( .A(n35763), .B(n35762), .Z(n35782) );
  OR U36260 ( .A(n35765), .B(n35764), .Z(n35769) );
  OR U36261 ( .A(n35767), .B(n35766), .Z(n35768) );
  AND U36262 ( .A(n35769), .B(n35768), .Z(n35781) );
  XNOR U36263 ( .A(n35782), .B(n35781), .Z(n35783) );
  XNOR U36264 ( .A(n35784), .B(n35783), .Z(n35776) );
  XNOR U36265 ( .A(n35775), .B(n35776), .Z(n35777) );
  XNOR U36266 ( .A(n35778), .B(n35777), .Z(n35915) );
  XNOR U36267 ( .A(n35915), .B(sreg[478]), .Z(n35917) );
  NAND U36268 ( .A(n35770), .B(sreg[477]), .Z(n35774) );
  OR U36269 ( .A(n35772), .B(n35771), .Z(n35773) );
  AND U36270 ( .A(n35774), .B(n35773), .Z(n35916) );
  XOR U36271 ( .A(n35917), .B(n35916), .Z(c[478]) );
  NANDN U36272 ( .A(n35776), .B(n35775), .Z(n35780) );
  NAND U36273 ( .A(n35778), .B(n35777), .Z(n35779) );
  NAND U36274 ( .A(n35780), .B(n35779), .Z(n35923) );
  NANDN U36275 ( .A(n35782), .B(n35781), .Z(n35786) );
  NAND U36276 ( .A(n35784), .B(n35783), .Z(n35785) );
  NAND U36277 ( .A(n35786), .B(n35785), .Z(n35920) );
  NANDN U36278 ( .A(n35792), .B(n35791), .Z(n35796) );
  NAND U36279 ( .A(n35794), .B(n35793), .Z(n35795) );
  AND U36280 ( .A(n35796), .B(n35795), .Z(n36056) );
  XNOR U36281 ( .A(n36055), .B(n36056), .Z(n36057) );
  NANDN U36282 ( .A(n35798), .B(n35797), .Z(n35802) );
  NANDN U36283 ( .A(n35800), .B(n35799), .Z(n35801) );
  NAND U36284 ( .A(n35802), .B(n35801), .Z(n36040) );
  NANDN U36285 ( .A(n35804), .B(n35803), .Z(n35808) );
  NAND U36286 ( .A(n35806), .B(n35805), .Z(n35807) );
  NAND U36287 ( .A(n35808), .B(n35807), .Z(n36037) );
  XNOR U36288 ( .A(b[25]), .B(n36934), .Z(n35953) );
  NAND U36289 ( .A(n35953), .B(n38325), .Z(n35811) );
  NANDN U36290 ( .A(n35809), .B(n38326), .Z(n35810) );
  NAND U36291 ( .A(n35811), .B(n35810), .Z(n35947) );
  NANDN U36292 ( .A(n35812), .B(n38205), .Z(n35814) );
  XOR U36293 ( .A(n1057), .B(n37184), .Z(n35959) );
  NANDN U36294 ( .A(n38268), .B(n35959), .Z(n35813) );
  NAND U36295 ( .A(n35814), .B(n35813), .Z(n35944) );
  XOR U36296 ( .A(a[249]), .B(b[7]), .Z(n35956) );
  NAND U36297 ( .A(n35956), .B(n36701), .Z(n35817) );
  NANDN U36298 ( .A(n35815), .B(n36702), .Z(n35816) );
  AND U36299 ( .A(n35817), .B(n35816), .Z(n35945) );
  XNOR U36300 ( .A(n35944), .B(n35945), .Z(n35946) );
  XOR U36301 ( .A(n35947), .B(n35946), .Z(n35989) );
  NANDN U36302 ( .A(n1049), .B(a[255]), .Z(n35818) );
  XNOR U36303 ( .A(b[1]), .B(n35818), .Z(n35820) );
  IV U36304 ( .A(a[254]), .Z(n38532) );
  NANDN U36305 ( .A(n38532), .B(n1049), .Z(n35819) );
  AND U36306 ( .A(n35820), .B(n35819), .Z(n36015) );
  NAND U36307 ( .A(n35821), .B(n38490), .Z(n35823) );
  XNOR U36308 ( .A(n1058), .B(a[227]), .Z(n35950) );
  NANDN U36309 ( .A(n1048), .B(n35950), .Z(n35822) );
  NAND U36310 ( .A(n35823), .B(n35822), .Z(n36013) );
  NANDN U36311 ( .A(n1059), .B(a[223]), .Z(n36014) );
  XNOR U36312 ( .A(n36013), .B(n36014), .Z(n36016) );
  XOR U36313 ( .A(n36015), .B(n36016), .Z(n35990) );
  XNOR U36314 ( .A(n35989), .B(n35990), .Z(n35992) );
  XNOR U36315 ( .A(b[15]), .B(a[241]), .Z(n35962) );
  OR U36316 ( .A(n35962), .B(n37665), .Z(n35826) );
  NANDN U36317 ( .A(n35824), .B(n37604), .Z(n35825) );
  NAND U36318 ( .A(n35826), .B(n35825), .Z(n36034) );
  XOR U36319 ( .A(b[21]), .B(n37420), .Z(n35965) );
  NANDN U36320 ( .A(n35965), .B(n38101), .Z(n35829) );
  NANDN U36321 ( .A(n35827), .B(n38102), .Z(n35828) );
  NAND U36322 ( .A(n35829), .B(n35828), .Z(n36031) );
  XNOR U36323 ( .A(a[247]), .B(b[9]), .Z(n35968) );
  NANDN U36324 ( .A(n35968), .B(n36925), .Z(n35832) );
  NANDN U36325 ( .A(n35830), .B(n36926), .Z(n35831) );
  AND U36326 ( .A(n35832), .B(n35831), .Z(n36032) );
  XNOR U36327 ( .A(n36031), .B(n36032), .Z(n36033) );
  XNOR U36328 ( .A(n36034), .B(n36033), .Z(n36022) );
  XOR U36329 ( .A(n38110), .B(b[13]), .Z(n35971) );
  NANDN U36330 ( .A(n35971), .B(n37424), .Z(n35835) );
  NAND U36331 ( .A(n37425), .B(n35833), .Z(n35834) );
  NAND U36332 ( .A(n35835), .B(n35834), .Z(n36020) );
  XOR U36333 ( .A(n38213), .B(b[11]), .Z(n35974) );
  OR U36334 ( .A(n35974), .B(n37311), .Z(n35838) );
  NAND U36335 ( .A(n37218), .B(n35836), .Z(n35837) );
  AND U36336 ( .A(n35838), .B(n35837), .Z(n36019) );
  XNOR U36337 ( .A(n36020), .B(n36019), .Z(n36021) );
  XOR U36338 ( .A(n36022), .B(n36021), .Z(n35991) );
  XNOR U36339 ( .A(n35992), .B(n35991), .Z(n35935) );
  NANDN U36340 ( .A(n35840), .B(n35839), .Z(n35844) );
  NAND U36341 ( .A(n35842), .B(n35841), .Z(n35843) );
  NAND U36342 ( .A(n35844), .B(n35843), .Z(n35932) );
  NANDN U36343 ( .A(n35846), .B(n35845), .Z(n35850) );
  NAND U36344 ( .A(n35848), .B(n35847), .Z(n35849) );
  AND U36345 ( .A(n35850), .B(n35849), .Z(n35933) );
  XNOR U36346 ( .A(n35932), .B(n35933), .Z(n35934) );
  XOR U36347 ( .A(n35935), .B(n35934), .Z(n36038) );
  XOR U36348 ( .A(n36037), .B(n36038), .Z(n36039) );
  XNOR U36349 ( .A(n36040), .B(n36039), .Z(n36052) );
  NANDN U36350 ( .A(n35852), .B(n35851), .Z(n35856) );
  NAND U36351 ( .A(n35854), .B(n35853), .Z(n35855) );
  NAND U36352 ( .A(n35856), .B(n35855), .Z(n36049) );
  NANDN U36353 ( .A(n35858), .B(n35857), .Z(n35862) );
  NANDN U36354 ( .A(n35860), .B(n35859), .Z(n35861) );
  NAND U36355 ( .A(n35862), .B(n35861), .Z(n36046) );
  XOR U36356 ( .A(b[27]), .B(a[229]), .Z(n36007) );
  NAND U36357 ( .A(n38423), .B(n36007), .Z(n35865) );
  NANDN U36358 ( .A(n35863), .B(n38424), .Z(n35864) );
  NAND U36359 ( .A(n35865), .B(n35864), .Z(n35941) );
  XNOR U36360 ( .A(a[251]), .B(b[5]), .Z(n36010) );
  NANDN U36361 ( .A(n36010), .B(n36587), .Z(n35868) );
  NANDN U36362 ( .A(n35866), .B(n36588), .Z(n35867) );
  NAND U36363 ( .A(n35868), .B(n35867), .Z(n35938) );
  XNOR U36364 ( .A(b[19]), .B(a[237]), .Z(n36004) );
  NANDN U36365 ( .A(n36004), .B(n37934), .Z(n35871) );
  NANDN U36366 ( .A(n35869), .B(n37935), .Z(n35870) );
  AND U36367 ( .A(n35871), .B(n35870), .Z(n35939) );
  XNOR U36368 ( .A(n35938), .B(n35939), .Z(n35940) );
  XNOR U36369 ( .A(n35941), .B(n35940), .Z(n35978) );
  NANDN U36370 ( .A(n35872), .B(n37762), .Z(n35874) );
  XOR U36371 ( .A(b[17]), .B(a[239]), .Z(n35995) );
  NAND U36372 ( .A(n35995), .B(n37764), .Z(n35873) );
  NAND U36373 ( .A(n35874), .B(n35873), .Z(n36028) );
  XOR U36374 ( .A(b[31]), .B(n36167), .Z(n35998) );
  NANDN U36375 ( .A(n35998), .B(n38552), .Z(n35877) );
  NANDN U36376 ( .A(n35875), .B(n38553), .Z(n35876) );
  NAND U36377 ( .A(n35877), .B(n35876), .Z(n36025) );
  OR U36378 ( .A(n35878), .B(n36105), .Z(n35880) );
  XNOR U36379 ( .A(a[253]), .B(b[3]), .Z(n36001) );
  NANDN U36380 ( .A(n36001), .B(n36107), .Z(n35879) );
  AND U36381 ( .A(n35880), .B(n35879), .Z(n36026) );
  XNOR U36382 ( .A(n36025), .B(n36026), .Z(n36027) );
  XOR U36383 ( .A(n36028), .B(n36027), .Z(n35977) );
  XOR U36384 ( .A(n35978), .B(n35977), .Z(n35980) );
  NANDN U36385 ( .A(n35882), .B(n35881), .Z(n35886) );
  NAND U36386 ( .A(n35884), .B(n35883), .Z(n35885) );
  NAND U36387 ( .A(n35886), .B(n35885), .Z(n35979) );
  XNOR U36388 ( .A(n35980), .B(n35979), .Z(n36043) );
  NANDN U36389 ( .A(n35888), .B(n35887), .Z(n35892) );
  NAND U36390 ( .A(n35890), .B(n35889), .Z(n35891) );
  NAND U36391 ( .A(n35892), .B(n35891), .Z(n35984) );
  NANDN U36392 ( .A(n35894), .B(n35893), .Z(n35898) );
  NAND U36393 ( .A(n35896), .B(n35895), .Z(n35897) );
  AND U36394 ( .A(n35898), .B(n35897), .Z(n35983) );
  XNOR U36395 ( .A(n35984), .B(n35983), .Z(n35985) );
  NANDN U36396 ( .A(n35900), .B(n35899), .Z(n35904) );
  NAND U36397 ( .A(n35902), .B(n35901), .Z(n35903) );
  AND U36398 ( .A(n35904), .B(n35903), .Z(n35986) );
  XNOR U36399 ( .A(n35985), .B(n35986), .Z(n36044) );
  XNOR U36400 ( .A(n36043), .B(n36044), .Z(n36045) );
  XNOR U36401 ( .A(n36046), .B(n36045), .Z(n36050) );
  XNOR U36402 ( .A(n36049), .B(n36050), .Z(n36051) );
  XOR U36403 ( .A(n36052), .B(n36051), .Z(n35929) );
  NANDN U36404 ( .A(n35906), .B(n35905), .Z(n35910) );
  NANDN U36405 ( .A(n35908), .B(n35907), .Z(n35909) );
  NAND U36406 ( .A(n35910), .B(n35909), .Z(n35926) );
  XNOR U36407 ( .A(n35926), .B(n35927), .Z(n35928) );
  XOR U36408 ( .A(n35929), .B(n35928), .Z(n36058) );
  XNOR U36409 ( .A(n36057), .B(n36058), .Z(n35921) );
  XNOR U36410 ( .A(n35920), .B(n35921), .Z(n35922) );
  XNOR U36411 ( .A(n35923), .B(n35922), .Z(n36061) );
  XNOR U36412 ( .A(n36061), .B(sreg[479]), .Z(n36063) );
  NAND U36413 ( .A(n35915), .B(sreg[478]), .Z(n35919) );
  OR U36414 ( .A(n35917), .B(n35916), .Z(n35918) );
  AND U36415 ( .A(n35919), .B(n35918), .Z(n36062) );
  XOR U36416 ( .A(n36063), .B(n36062), .Z(c[479]) );
  NANDN U36417 ( .A(n35921), .B(n35920), .Z(n35925) );
  NAND U36418 ( .A(n35923), .B(n35922), .Z(n35924) );
  NAND U36419 ( .A(n35925), .B(n35924), .Z(n36071) );
  NANDN U36420 ( .A(n35927), .B(n35926), .Z(n35931) );
  NANDN U36421 ( .A(n35929), .B(n35928), .Z(n35930) );
  NAND U36422 ( .A(n35931), .B(n35930), .Z(n36207) );
  NANDN U36423 ( .A(n35933), .B(n35932), .Z(n35937) );
  NANDN U36424 ( .A(n35935), .B(n35934), .Z(n35936) );
  NAND U36425 ( .A(n35937), .B(n35936), .Z(n36089) );
  NANDN U36426 ( .A(n35939), .B(n35938), .Z(n35943) );
  NAND U36427 ( .A(n35941), .B(n35940), .Z(n35942) );
  NAND U36428 ( .A(n35943), .B(n35942), .Z(n36187) );
  NANDN U36429 ( .A(n35945), .B(n35944), .Z(n35949) );
  NAND U36430 ( .A(n35947), .B(n35946), .Z(n35948) );
  AND U36431 ( .A(n35949), .B(n35948), .Z(n36186) );
  XNOR U36432 ( .A(n36187), .B(n36186), .Z(n36188) );
  NAND U36433 ( .A(n38490), .B(n35950), .Z(n35952) );
  XOR U36434 ( .A(b[29]), .B(n36592), .Z(n36168) );
  OR U36435 ( .A(n36168), .B(n1048), .Z(n35951) );
  NAND U36436 ( .A(n35952), .B(n35951), .Z(n36119) );
  NANDN U36437 ( .A(n1059), .B(a[224]), .Z(n36120) );
  XNOR U36438 ( .A(n36119), .B(n36120), .Z(n36121) );
  XNOR U36439 ( .A(n36122), .B(n36121), .Z(n36096) );
  XNOR U36440 ( .A(b[25]), .B(a[232]), .Z(n36102) );
  NANDN U36441 ( .A(n36102), .B(n38325), .Z(n35955) );
  NAND U36442 ( .A(n38326), .B(n35953), .Z(n35954) );
  NAND U36443 ( .A(n35955), .B(n35954), .Z(n36181) );
  XNOR U36444 ( .A(a[250]), .B(b[7]), .Z(n36149) );
  NANDN U36445 ( .A(n36149), .B(n36701), .Z(n35958) );
  NAND U36446 ( .A(n36702), .B(n35956), .Z(n35957) );
  AND U36447 ( .A(n35958), .B(n35957), .Z(n36180) );
  XNOR U36448 ( .A(n36181), .B(n36180), .Z(n36182) );
  XOR U36449 ( .A(b[23]), .B(n37080), .Z(n36158) );
  OR U36450 ( .A(n36158), .B(n38268), .Z(n35961) );
  NAND U36451 ( .A(n38205), .B(n35959), .Z(n35960) );
  AND U36452 ( .A(n35961), .B(n35960), .Z(n36183) );
  XNOR U36453 ( .A(n36182), .B(n36183), .Z(n36097) );
  XOR U36454 ( .A(n36096), .B(n36097), .Z(n36099) );
  XOR U36455 ( .A(a[242]), .B(n1054), .Z(n36113) );
  OR U36456 ( .A(n36113), .B(n37665), .Z(n35964) );
  NANDN U36457 ( .A(n35962), .B(n37604), .Z(n35963) );
  NAND U36458 ( .A(n35964), .B(n35963), .Z(n36140) );
  XOR U36459 ( .A(b[21]), .B(n37106), .Z(n36161) );
  NANDN U36460 ( .A(n36161), .B(n38101), .Z(n35967) );
  NANDN U36461 ( .A(n35965), .B(n38102), .Z(n35966) );
  NAND U36462 ( .A(n35967), .B(n35966), .Z(n36137) );
  XOR U36463 ( .A(a[248]), .B(n1052), .Z(n36143) );
  NANDN U36464 ( .A(n36143), .B(n36925), .Z(n35970) );
  NANDN U36465 ( .A(n35968), .B(n36926), .Z(n35969) );
  AND U36466 ( .A(n35970), .B(n35969), .Z(n36138) );
  XNOR U36467 ( .A(n36137), .B(n36138), .Z(n36139) );
  XNOR U36468 ( .A(n36140), .B(n36139), .Z(n36128) );
  XOR U36469 ( .A(a[244]), .B(n1053), .Z(n36152) );
  NANDN U36470 ( .A(n36152), .B(n37424), .Z(n35973) );
  NANDN U36471 ( .A(n35971), .B(n37425), .Z(n35972) );
  NAND U36472 ( .A(n35973), .B(n35972), .Z(n36126) );
  XNOR U36473 ( .A(a[246]), .B(b[11]), .Z(n36146) );
  OR U36474 ( .A(n36146), .B(n37311), .Z(n35976) );
  NANDN U36475 ( .A(n35974), .B(n37218), .Z(n35975) );
  AND U36476 ( .A(n35976), .B(n35975), .Z(n36125) );
  XNOR U36477 ( .A(n36126), .B(n36125), .Z(n36127) );
  XOR U36478 ( .A(n36128), .B(n36127), .Z(n36098) );
  XNOR U36479 ( .A(n36099), .B(n36098), .Z(n36189) );
  XNOR U36480 ( .A(n36188), .B(n36189), .Z(n36086) );
  NANDN U36481 ( .A(n35978), .B(n35977), .Z(n35982) );
  OR U36482 ( .A(n35980), .B(n35979), .Z(n35981) );
  AND U36483 ( .A(n35982), .B(n35981), .Z(n36087) );
  XNOR U36484 ( .A(n36086), .B(n36087), .Z(n36088) );
  XNOR U36485 ( .A(n36089), .B(n36088), .Z(n36198) );
  NANDN U36486 ( .A(n35984), .B(n35983), .Z(n35988) );
  NAND U36487 ( .A(n35986), .B(n35985), .Z(n35987) );
  AND U36488 ( .A(n35988), .B(n35987), .Z(n36199) );
  XOR U36489 ( .A(n36198), .B(n36199), .Z(n36201) );
  OR U36490 ( .A(n35990), .B(n35989), .Z(n35994) );
  NANDN U36491 ( .A(n35992), .B(n35991), .Z(n35993) );
  NAND U36492 ( .A(n35994), .B(n35993), .Z(n36080) );
  NAND U36493 ( .A(n35995), .B(n37762), .Z(n35997) );
  XNOR U36494 ( .A(b[17]), .B(a[240]), .Z(n36110) );
  NANDN U36495 ( .A(n36110), .B(n37764), .Z(n35996) );
  NAND U36496 ( .A(n35997), .B(n35996), .Z(n36134) );
  XOR U36497 ( .A(n1059), .B(n36280), .Z(n36171) );
  NAND U36498 ( .A(n36171), .B(n38552), .Z(n36000) );
  NANDN U36499 ( .A(n35998), .B(n38553), .Z(n35999) );
  NAND U36500 ( .A(n36000), .B(n35999), .Z(n36131) );
  OR U36501 ( .A(n36001), .B(n36105), .Z(n36003) );
  XOR U36502 ( .A(a[254]), .B(n1050), .Z(n36106) );
  NANDN U36503 ( .A(n36106), .B(n36107), .Z(n36002) );
  AND U36504 ( .A(n36003), .B(n36002), .Z(n36132) );
  XNOR U36505 ( .A(n36131), .B(n36132), .Z(n36133) );
  XNOR U36506 ( .A(n36134), .B(n36133), .Z(n36192) );
  XOR U36507 ( .A(b[19]), .B(n37467), .Z(n36155) );
  NANDN U36508 ( .A(n36155), .B(n37934), .Z(n36006) );
  NANDN U36509 ( .A(n36004), .B(n37935), .Z(n36005) );
  NAND U36510 ( .A(n36006), .B(n36005), .Z(n36177) );
  XNOR U36511 ( .A(b[27]), .B(n36333), .Z(n36116) );
  NAND U36512 ( .A(n38423), .B(n36116), .Z(n36009) );
  NAND U36513 ( .A(n36007), .B(n38424), .Z(n36008) );
  NAND U36514 ( .A(n36009), .B(n36008), .Z(n36174) );
  XOR U36515 ( .A(a[252]), .B(n1051), .Z(n36164) );
  NANDN U36516 ( .A(n36164), .B(n36587), .Z(n36012) );
  NANDN U36517 ( .A(n36010), .B(n36588), .Z(n36011) );
  AND U36518 ( .A(n36012), .B(n36011), .Z(n36175) );
  XNOR U36519 ( .A(n36174), .B(n36175), .Z(n36176) );
  XOR U36520 ( .A(n36177), .B(n36176), .Z(n36193) );
  XNOR U36521 ( .A(n36192), .B(n36193), .Z(n36194) );
  NANDN U36522 ( .A(n36014), .B(n36013), .Z(n36018) );
  NAND U36523 ( .A(n36016), .B(n36015), .Z(n36017) );
  AND U36524 ( .A(n36018), .B(n36017), .Z(n36195) );
  XNOR U36525 ( .A(n36194), .B(n36195), .Z(n36081) );
  XNOR U36526 ( .A(n36080), .B(n36081), .Z(n36082) );
  NANDN U36527 ( .A(n36020), .B(n36019), .Z(n36024) );
  NAND U36528 ( .A(n36022), .B(n36021), .Z(n36023) );
  NAND U36529 ( .A(n36024), .B(n36023), .Z(n36093) );
  NANDN U36530 ( .A(n36026), .B(n36025), .Z(n36030) );
  NAND U36531 ( .A(n36028), .B(n36027), .Z(n36029) );
  NAND U36532 ( .A(n36030), .B(n36029), .Z(n36091) );
  NANDN U36533 ( .A(n36032), .B(n36031), .Z(n36036) );
  NAND U36534 ( .A(n36034), .B(n36033), .Z(n36035) );
  AND U36535 ( .A(n36036), .B(n36035), .Z(n36090) );
  XNOR U36536 ( .A(n36091), .B(n36090), .Z(n36092) );
  XOR U36537 ( .A(n36093), .B(n36092), .Z(n36083) );
  XOR U36538 ( .A(n36082), .B(n36083), .Z(n36200) );
  XOR U36539 ( .A(n36201), .B(n36200), .Z(n36077) );
  OR U36540 ( .A(n36038), .B(n36037), .Z(n36042) );
  NAND U36541 ( .A(n36040), .B(n36039), .Z(n36041) );
  NAND U36542 ( .A(n36042), .B(n36041), .Z(n36074) );
  NANDN U36543 ( .A(n36044), .B(n36043), .Z(n36048) );
  NAND U36544 ( .A(n36046), .B(n36045), .Z(n36047) );
  NAND U36545 ( .A(n36048), .B(n36047), .Z(n36075) );
  XNOR U36546 ( .A(n36074), .B(n36075), .Z(n36076) );
  XNOR U36547 ( .A(n36077), .B(n36076), .Z(n36205) );
  NANDN U36548 ( .A(n36050), .B(n36049), .Z(n36054) );
  NAND U36549 ( .A(n36052), .B(n36051), .Z(n36053) );
  AND U36550 ( .A(n36054), .B(n36053), .Z(n36204) );
  XNOR U36551 ( .A(n36205), .B(n36204), .Z(n36206) );
  XNOR U36552 ( .A(n36207), .B(n36206), .Z(n36068) );
  NANDN U36553 ( .A(n36056), .B(n36055), .Z(n36060) );
  NANDN U36554 ( .A(n36058), .B(n36057), .Z(n36059) );
  NAND U36555 ( .A(n36060), .B(n36059), .Z(n36069) );
  XNOR U36556 ( .A(n36068), .B(n36069), .Z(n36070) );
  XOR U36557 ( .A(n36071), .B(n36070), .Z(n36067) );
  NAND U36558 ( .A(n36061), .B(sreg[479]), .Z(n36065) );
  OR U36559 ( .A(n36063), .B(n36062), .Z(n36064) );
  AND U36560 ( .A(n36065), .B(n36064), .Z(n36066) );
  XOR U36561 ( .A(n36067), .B(n36066), .Z(c[480]) );
  OR U36562 ( .A(n36067), .B(n36066), .Z(n36351) );
  NANDN U36563 ( .A(n36069), .B(n36068), .Z(n36073) );
  NAND U36564 ( .A(n36071), .B(n36070), .Z(n36072) );
  NAND U36565 ( .A(n36073), .B(n36072), .Z(n36213) );
  NANDN U36566 ( .A(n36075), .B(n36074), .Z(n36079) );
  NAND U36567 ( .A(n36077), .B(n36076), .Z(n36078) );
  NAND U36568 ( .A(n36079), .B(n36078), .Z(n36219) );
  NANDN U36569 ( .A(n36081), .B(n36080), .Z(n36085) );
  NAND U36570 ( .A(n36083), .B(n36082), .Z(n36084) );
  NAND U36571 ( .A(n36085), .B(n36084), .Z(n36220) );
  XNOR U36572 ( .A(n36220), .B(n36221), .Z(n36222) );
  NANDN U36573 ( .A(n36091), .B(n36090), .Z(n36095) );
  NAND U36574 ( .A(n36093), .B(n36092), .Z(n36094) );
  NAND U36575 ( .A(n36095), .B(n36094), .Z(n36345) );
  NANDN U36576 ( .A(n36097), .B(n36096), .Z(n36101) );
  NANDN U36577 ( .A(n36099), .B(n36098), .Z(n36100) );
  NAND U36578 ( .A(n36101), .B(n36100), .Z(n36299) );
  XNOR U36579 ( .A(b[25]), .B(a[233]), .Z(n36259) );
  NANDN U36580 ( .A(n36259), .B(n38325), .Z(n36104) );
  NANDN U36581 ( .A(n36102), .B(n38326), .Z(n36103) );
  NAND U36582 ( .A(n36104), .B(n36103), .Z(n36235) );
  OR U36583 ( .A(n36106), .B(n36105), .Z(n36109) );
  IV U36584 ( .A(a[255]), .Z(n38595) );
  XNOR U36585 ( .A(n38595), .B(b[3]), .Z(n36277) );
  NAND U36586 ( .A(n36277), .B(n36107), .Z(n36108) );
  NAND U36587 ( .A(n36109), .B(n36108), .Z(n36232) );
  NANDN U36588 ( .A(n36110), .B(n37762), .Z(n36112) );
  XOR U36589 ( .A(b[17]), .B(a[241]), .Z(n36273) );
  NAND U36590 ( .A(n36273), .B(n37764), .Z(n36111) );
  AND U36591 ( .A(n36112), .B(n36111), .Z(n36233) );
  XNOR U36592 ( .A(n36232), .B(n36233), .Z(n36234) );
  XNOR U36593 ( .A(n36235), .B(n36234), .Z(n36294) );
  XNOR U36594 ( .A(n38110), .B(b[15]), .Z(n36329) );
  NANDN U36595 ( .A(n37665), .B(n36329), .Z(n36115) );
  NANDN U36596 ( .A(n36113), .B(n37604), .Z(n36114) );
  AND U36597 ( .A(n36115), .B(n36114), .Z(n36262) );
  XNOR U36598 ( .A(b[1]), .B(n36262), .Z(n36264) );
  XNOR U36599 ( .A(b[27]), .B(a[231]), .Z(n36270) );
  NANDN U36600 ( .A(n36270), .B(n38423), .Z(n36118) );
  NAND U36601 ( .A(n38424), .B(n36116), .Z(n36117) );
  AND U36602 ( .A(n36118), .B(n36117), .Z(n36263) );
  XNOR U36603 ( .A(n36264), .B(n36263), .Z(n36293) );
  XOR U36604 ( .A(n36294), .B(n36293), .Z(n36295) );
  NANDN U36605 ( .A(n36120), .B(n36119), .Z(n36124) );
  NAND U36606 ( .A(n36122), .B(n36121), .Z(n36123) );
  AND U36607 ( .A(n36124), .B(n36123), .Z(n36296) );
  XNOR U36608 ( .A(n36295), .B(n36296), .Z(n36300) );
  XNOR U36609 ( .A(n36299), .B(n36300), .Z(n36301) );
  NANDN U36610 ( .A(n36126), .B(n36125), .Z(n36130) );
  NAND U36611 ( .A(n36128), .B(n36127), .Z(n36129) );
  NAND U36612 ( .A(n36130), .B(n36129), .Z(n36320) );
  NANDN U36613 ( .A(n36132), .B(n36131), .Z(n36136) );
  NAND U36614 ( .A(n36134), .B(n36133), .Z(n36135) );
  NAND U36615 ( .A(n36136), .B(n36135), .Z(n36318) );
  NANDN U36616 ( .A(n36138), .B(n36137), .Z(n36142) );
  NAND U36617 ( .A(n36140), .B(n36139), .Z(n36141) );
  AND U36618 ( .A(n36142), .B(n36141), .Z(n36317) );
  XNOR U36619 ( .A(n36318), .B(n36317), .Z(n36319) );
  XOR U36620 ( .A(n36320), .B(n36319), .Z(n36302) );
  XOR U36621 ( .A(n36301), .B(n36302), .Z(n36344) );
  XNOR U36622 ( .A(n36345), .B(n36344), .Z(n36346) );
  XNOR U36623 ( .A(a[249]), .B(b[9]), .Z(n36244) );
  NANDN U36624 ( .A(n36244), .B(n36925), .Z(n36145) );
  NANDN U36625 ( .A(n36143), .B(n36926), .Z(n36144) );
  NAND U36626 ( .A(n36145), .B(n36144), .Z(n36229) );
  XOR U36627 ( .A(a[247]), .B(b[11]), .Z(n36256) );
  NANDN U36628 ( .A(n37311), .B(n36256), .Z(n36148) );
  NANDN U36629 ( .A(n36146), .B(n37218), .Z(n36147) );
  NAND U36630 ( .A(n36148), .B(n36147), .Z(n36226) );
  XOR U36631 ( .A(a[251]), .B(b[7]), .Z(n36247) );
  NAND U36632 ( .A(n36247), .B(n36701), .Z(n36151) );
  NANDN U36633 ( .A(n36149), .B(n36702), .Z(n36150) );
  NAND U36634 ( .A(n36151), .B(n36150), .Z(n36241) );
  XOR U36635 ( .A(a[245]), .B(n1053), .Z(n36253) );
  NANDN U36636 ( .A(n36253), .B(n37424), .Z(n36154) );
  NANDN U36637 ( .A(n36152), .B(n37425), .Z(n36153) );
  NAND U36638 ( .A(n36154), .B(n36153), .Z(n36238) );
  XNOR U36639 ( .A(n1055), .B(a[239]), .Z(n36281) );
  NAND U36640 ( .A(n36281), .B(n37934), .Z(n36157) );
  NANDN U36641 ( .A(n36155), .B(n37935), .Z(n36156) );
  AND U36642 ( .A(n36157), .B(n36156), .Z(n36239) );
  XNOR U36643 ( .A(n36238), .B(n36239), .Z(n36240) );
  XNOR U36644 ( .A(n36241), .B(n36240), .Z(n36227) );
  XNOR U36645 ( .A(n36226), .B(n36227), .Z(n36228) );
  XOR U36646 ( .A(n36229), .B(n36228), .Z(n36290) );
  NANDN U36647 ( .A(n36158), .B(n38205), .Z(n36160) );
  XOR U36648 ( .A(b[23]), .B(n37420), .Z(n36267) );
  OR U36649 ( .A(n36267), .B(n38268), .Z(n36159) );
  NAND U36650 ( .A(n36160), .B(n36159), .Z(n36326) );
  XNOR U36651 ( .A(b[21]), .B(a[237]), .Z(n36250) );
  NANDN U36652 ( .A(n36250), .B(n38101), .Z(n36163) );
  NANDN U36653 ( .A(n36161), .B(n38102), .Z(n36162) );
  NAND U36654 ( .A(n36163), .B(n36162), .Z(n36323) );
  XNOR U36655 ( .A(a[253]), .B(n1051), .Z(n36284) );
  NAND U36656 ( .A(n36284), .B(n36587), .Z(n36166) );
  NANDN U36657 ( .A(n36164), .B(n36588), .Z(n36165) );
  AND U36658 ( .A(n36166), .B(n36165), .Z(n36324) );
  XNOR U36659 ( .A(n36323), .B(n36324), .Z(n36325) );
  XOR U36660 ( .A(n36326), .B(n36325), .Z(n36288) );
  ANDN U36661 ( .B(b[31]), .A(n36167), .Z(n36396) );
  IV U36662 ( .A(n36396), .Z(n36551) );
  NANDN U36663 ( .A(n36168), .B(n38490), .Z(n36170) );
  XNOR U36664 ( .A(n1058), .B(a[229]), .Z(n36332) );
  NANDN U36665 ( .A(n1048), .B(n36332), .Z(n36169) );
  AND U36666 ( .A(n36170), .B(n36169), .Z(n36339) );
  XOR U36667 ( .A(n36551), .B(n36339), .Z(n36341) );
  XNOR U36668 ( .A(b[31]), .B(a[227]), .Z(n36336) );
  NANDN U36669 ( .A(n36336), .B(n38552), .Z(n36173) );
  NAND U36670 ( .A(n38553), .B(n36171), .Z(n36172) );
  NAND U36671 ( .A(n36173), .B(n36172), .Z(n36340) );
  XOR U36672 ( .A(n36341), .B(n36340), .Z(n36287) );
  XOR U36673 ( .A(n36288), .B(n36287), .Z(n36289) );
  XOR U36674 ( .A(n36290), .B(n36289), .Z(n36314) );
  NANDN U36675 ( .A(n36175), .B(n36174), .Z(n36179) );
  NAND U36676 ( .A(n36177), .B(n36176), .Z(n36178) );
  NAND U36677 ( .A(n36179), .B(n36178), .Z(n36311) );
  NANDN U36678 ( .A(n36181), .B(n36180), .Z(n36185) );
  NAND U36679 ( .A(n36183), .B(n36182), .Z(n36184) );
  NAND U36680 ( .A(n36185), .B(n36184), .Z(n36312) );
  XNOR U36681 ( .A(n36311), .B(n36312), .Z(n36313) );
  XNOR U36682 ( .A(n36314), .B(n36313), .Z(n36308) );
  NANDN U36683 ( .A(n36187), .B(n36186), .Z(n36191) );
  NAND U36684 ( .A(n36189), .B(n36188), .Z(n36190) );
  NAND U36685 ( .A(n36191), .B(n36190), .Z(n36305) );
  NANDN U36686 ( .A(n36193), .B(n36192), .Z(n36197) );
  NAND U36687 ( .A(n36195), .B(n36194), .Z(n36196) );
  AND U36688 ( .A(n36197), .B(n36196), .Z(n36306) );
  XNOR U36689 ( .A(n36305), .B(n36306), .Z(n36307) );
  XOR U36690 ( .A(n36308), .B(n36307), .Z(n36347) );
  XOR U36691 ( .A(n36346), .B(n36347), .Z(n36223) );
  XNOR U36692 ( .A(n36222), .B(n36223), .Z(n36216) );
  NANDN U36693 ( .A(n36199), .B(n36198), .Z(n36203) );
  NANDN U36694 ( .A(n36201), .B(n36200), .Z(n36202) );
  NAND U36695 ( .A(n36203), .B(n36202), .Z(n36217) );
  XNOR U36696 ( .A(n36216), .B(n36217), .Z(n36218) );
  XNOR U36697 ( .A(n36219), .B(n36218), .Z(n36210) );
  NANDN U36698 ( .A(n36205), .B(n36204), .Z(n36209) );
  NAND U36699 ( .A(n36207), .B(n36206), .Z(n36208) );
  NAND U36700 ( .A(n36209), .B(n36208), .Z(n36211) );
  XNOR U36701 ( .A(n36210), .B(n36211), .Z(n36212) );
  XOR U36702 ( .A(n36213), .B(n36212), .Z(n36350) );
  XOR U36703 ( .A(n36351), .B(n36350), .Z(c[481]) );
  NANDN U36704 ( .A(n36211), .B(n36210), .Z(n36215) );
  NAND U36705 ( .A(n36213), .B(n36212), .Z(n36214) );
  AND U36706 ( .A(n36215), .B(n36214), .Z(n36357) );
  NANDN U36707 ( .A(n36221), .B(n36220), .Z(n36225) );
  NAND U36708 ( .A(n36223), .B(n36222), .Z(n36224) );
  NAND U36709 ( .A(n36225), .B(n36224), .Z(n36485) );
  NANDN U36710 ( .A(n36227), .B(n36226), .Z(n36231) );
  NAND U36711 ( .A(n36229), .B(n36228), .Z(n36230) );
  NAND U36712 ( .A(n36231), .B(n36230), .Z(n36469) );
  NANDN U36713 ( .A(n36233), .B(n36232), .Z(n36237) );
  NAND U36714 ( .A(n36235), .B(n36234), .Z(n36236) );
  NAND U36715 ( .A(n36237), .B(n36236), .Z(n36468) );
  NANDN U36716 ( .A(n36239), .B(n36238), .Z(n36243) );
  NAND U36717 ( .A(n36241), .B(n36240), .Z(n36242) );
  NAND U36718 ( .A(n36243), .B(n36242), .Z(n36380) );
  XOR U36719 ( .A(a[250]), .B(n1052), .Z(n36457) );
  NANDN U36720 ( .A(n36457), .B(n36925), .Z(n36246) );
  NANDN U36721 ( .A(n36244), .B(n36926), .Z(n36245) );
  NAND U36722 ( .A(n36246), .B(n36245), .Z(n36414) );
  XNOR U36723 ( .A(a[252]), .B(b[7]), .Z(n36430) );
  NANDN U36724 ( .A(n36430), .B(n36701), .Z(n36249) );
  NAND U36725 ( .A(n36247), .B(n36702), .Z(n36248) );
  NAND U36726 ( .A(n36249), .B(n36248), .Z(n36411) );
  XOR U36727 ( .A(b[21]), .B(n37467), .Z(n36436) );
  NANDN U36728 ( .A(n36436), .B(n38101), .Z(n36252) );
  NANDN U36729 ( .A(n36250), .B(n38102), .Z(n36251) );
  AND U36730 ( .A(n36252), .B(n36251), .Z(n36412) );
  XNOR U36731 ( .A(n36411), .B(n36412), .Z(n36413) );
  XNOR U36732 ( .A(n36414), .B(n36413), .Z(n36378) );
  XOR U36733 ( .A(a[246]), .B(n1053), .Z(n36384) );
  NANDN U36734 ( .A(n36384), .B(n37424), .Z(n36255) );
  NANDN U36735 ( .A(n36253), .B(n37425), .Z(n36254) );
  NAND U36736 ( .A(n36255), .B(n36254), .Z(n36448) );
  XNOR U36737 ( .A(a[248]), .B(b[11]), .Z(n36421) );
  OR U36738 ( .A(n36421), .B(n37311), .Z(n36258) );
  NAND U36739 ( .A(n36256), .B(n37218), .Z(n36257) );
  NAND U36740 ( .A(n36258), .B(n36257), .Z(n36445) );
  XNOR U36741 ( .A(b[25]), .B(a[234]), .Z(n36424) );
  NANDN U36742 ( .A(n36424), .B(n38325), .Z(n36261) );
  NANDN U36743 ( .A(n36259), .B(n38326), .Z(n36260) );
  AND U36744 ( .A(n36261), .B(n36260), .Z(n36446) );
  XNOR U36745 ( .A(n36445), .B(n36446), .Z(n36447) );
  XOR U36746 ( .A(n36448), .B(n36447), .Z(n36379) );
  XOR U36747 ( .A(n36378), .B(n36379), .Z(n36381) );
  XOR U36748 ( .A(n36380), .B(n36381), .Z(n36467) );
  XOR U36749 ( .A(n36468), .B(n36467), .Z(n36470) );
  XNOR U36750 ( .A(n36469), .B(n36470), .Z(n36478) );
  NAND U36751 ( .A(b[1]), .B(n36262), .Z(n36266) );
  NANDN U36752 ( .A(n36264), .B(n36263), .Z(n36265) );
  NAND U36753 ( .A(n36266), .B(n36265), .Z(n36420) );
  NANDN U36754 ( .A(n36267), .B(n38205), .Z(n36269) );
  XOR U36755 ( .A(b[23]), .B(n37106), .Z(n36451) );
  OR U36756 ( .A(n36451), .B(n38268), .Z(n36268) );
  NAND U36757 ( .A(n36269), .B(n36268), .Z(n36402) );
  XNOR U36758 ( .A(b[27]), .B(a[232]), .Z(n36427) );
  NANDN U36759 ( .A(n36427), .B(n38423), .Z(n36272) );
  NANDN U36760 ( .A(n36270), .B(n38424), .Z(n36271) );
  NAND U36761 ( .A(n36272), .B(n36271), .Z(n36399) );
  NAND U36762 ( .A(n36273), .B(n37762), .Z(n36275) );
  XNOR U36763 ( .A(b[17]), .B(a[242]), .Z(n36390) );
  NANDN U36764 ( .A(n36390), .B(n37764), .Z(n36274) );
  AND U36765 ( .A(n36275), .B(n36274), .Z(n36400) );
  XNOR U36766 ( .A(n36399), .B(n36400), .Z(n36401) );
  XNOR U36767 ( .A(n36402), .B(n36401), .Z(n36418) );
  NAND U36768 ( .A(b[1]), .B(b[2]), .Z(n36460) );
  XOR U36769 ( .A(n1050), .B(n36460), .Z(n36279) );
  XNOR U36770 ( .A(b[2]), .B(b[1]), .Z(n36276) );
  NANDN U36771 ( .A(n36277), .B(n36276), .Z(n36278) );
  AND U36772 ( .A(n36279), .B(n36278), .Z(n36393) );
  NANDN U36773 ( .A(n36280), .B(b[31]), .Z(n36394) );
  XNOR U36774 ( .A(n36393), .B(n36394), .Z(n36395) );
  XOR U36775 ( .A(n36551), .B(n36395), .Z(n36408) );
  XOR U36776 ( .A(n1055), .B(a[240]), .Z(n36464) );
  NANDN U36777 ( .A(n36464), .B(n37934), .Z(n36283) );
  NAND U36778 ( .A(n37935), .B(n36281), .Z(n36282) );
  NAND U36779 ( .A(n36283), .B(n36282), .Z(n36406) );
  XOR U36780 ( .A(n38532), .B(b[5]), .Z(n36461) );
  NANDN U36781 ( .A(n36461), .B(n36587), .Z(n36286) );
  NAND U36782 ( .A(n36588), .B(n36284), .Z(n36285) );
  AND U36783 ( .A(n36286), .B(n36285), .Z(n36405) );
  XNOR U36784 ( .A(n36406), .B(n36405), .Z(n36407) );
  XNOR U36785 ( .A(n36408), .B(n36407), .Z(n36417) );
  XOR U36786 ( .A(n36418), .B(n36417), .Z(n36419) );
  XNOR U36787 ( .A(n36420), .B(n36419), .Z(n36363) );
  NANDN U36788 ( .A(n36288), .B(n36287), .Z(n36292) );
  OR U36789 ( .A(n36290), .B(n36289), .Z(n36291) );
  NAND U36790 ( .A(n36292), .B(n36291), .Z(n36361) );
  NAND U36791 ( .A(n36294), .B(n36293), .Z(n36298) );
  NAND U36792 ( .A(n36296), .B(n36295), .Z(n36297) );
  AND U36793 ( .A(n36298), .B(n36297), .Z(n36360) );
  XNOR U36794 ( .A(n36361), .B(n36360), .Z(n36362) );
  XOR U36795 ( .A(n36363), .B(n36362), .Z(n36477) );
  XNOR U36796 ( .A(n36478), .B(n36477), .Z(n36480) );
  NANDN U36797 ( .A(n36300), .B(n36299), .Z(n36304) );
  NAND U36798 ( .A(n36302), .B(n36301), .Z(n36303) );
  NAND U36799 ( .A(n36304), .B(n36303), .Z(n36479) );
  XNOR U36800 ( .A(n36480), .B(n36479), .Z(n36476) );
  NANDN U36801 ( .A(n36306), .B(n36305), .Z(n36310) );
  NANDN U36802 ( .A(n36308), .B(n36307), .Z(n36309) );
  NAND U36803 ( .A(n36310), .B(n36309), .Z(n36474) );
  NANDN U36804 ( .A(n36312), .B(n36311), .Z(n36316) );
  NANDN U36805 ( .A(n36314), .B(n36313), .Z(n36315) );
  NAND U36806 ( .A(n36316), .B(n36315), .Z(n36369) );
  NANDN U36807 ( .A(n36318), .B(n36317), .Z(n36322) );
  NAND U36808 ( .A(n36320), .B(n36319), .Z(n36321) );
  NAND U36809 ( .A(n36322), .B(n36321), .Z(n36367) );
  NANDN U36810 ( .A(n36324), .B(n36323), .Z(n36328) );
  NAND U36811 ( .A(n36326), .B(n36325), .Z(n36327) );
  NAND U36812 ( .A(n36328), .B(n36327), .Z(n36374) );
  XOR U36813 ( .A(a[244]), .B(n1054), .Z(n36387) );
  OR U36814 ( .A(n36387), .B(n37665), .Z(n36331) );
  NAND U36815 ( .A(n36329), .B(n37604), .Z(n36330) );
  NAND U36816 ( .A(n36331), .B(n36330), .Z(n36442) );
  NAND U36817 ( .A(n36332), .B(n38490), .Z(n36335) );
  XOR U36818 ( .A(n1058), .B(n36333), .Z(n36454) );
  NANDN U36819 ( .A(n1048), .B(n36454), .Z(n36334) );
  NAND U36820 ( .A(n36335), .B(n36334), .Z(n36439) );
  XOR U36821 ( .A(b[31]), .B(n36592), .Z(n36433) );
  NANDN U36822 ( .A(n36433), .B(n38552), .Z(n36338) );
  NANDN U36823 ( .A(n36336), .B(n38553), .Z(n36337) );
  AND U36824 ( .A(n36338), .B(n36337), .Z(n36440) );
  XNOR U36825 ( .A(n36439), .B(n36440), .Z(n36441) );
  XNOR U36826 ( .A(n36442), .B(n36441), .Z(n36372) );
  NANDN U36827 ( .A(n36551), .B(n36339), .Z(n36343) );
  OR U36828 ( .A(n36341), .B(n36340), .Z(n36342) );
  AND U36829 ( .A(n36343), .B(n36342), .Z(n36373) );
  XOR U36830 ( .A(n36372), .B(n36373), .Z(n36375) );
  XOR U36831 ( .A(n36374), .B(n36375), .Z(n36366) );
  XOR U36832 ( .A(n36367), .B(n36366), .Z(n36368) );
  XNOR U36833 ( .A(n36369), .B(n36368), .Z(n36473) );
  XOR U36834 ( .A(n36474), .B(n36473), .Z(n36475) );
  XNOR U36835 ( .A(n36476), .B(n36475), .Z(n36483) );
  NAND U36836 ( .A(n36345), .B(n36344), .Z(n36349) );
  OR U36837 ( .A(n36347), .B(n36346), .Z(n36348) );
  NAND U36838 ( .A(n36349), .B(n36348), .Z(n36484) );
  XOR U36839 ( .A(n36483), .B(n36484), .Z(n36486) );
  XOR U36840 ( .A(n36485), .B(n36486), .Z(n36354) );
  XOR U36841 ( .A(n36355), .B(n36354), .Z(n36356) );
  XNOR U36842 ( .A(n36357), .B(n36356), .Z(n36353) );
  OR U36843 ( .A(n36351), .B(n36350), .Z(n36352) );
  XOR U36844 ( .A(n36353), .B(n36352), .Z(c[482]) );
  OR U36845 ( .A(n36353), .B(n36352), .Z(n36490) );
  OR U36846 ( .A(n36355), .B(n36354), .Z(n36359) );
  NANDN U36847 ( .A(n36357), .B(n36356), .Z(n36358) );
  AND U36848 ( .A(n36359), .B(n36358), .Z(n36494) );
  NANDN U36849 ( .A(n36361), .B(n36360), .Z(n36365) );
  NAND U36850 ( .A(n36363), .B(n36362), .Z(n36364) );
  NAND U36851 ( .A(n36365), .B(n36364), .Z(n36503) );
  NAND U36852 ( .A(n36367), .B(n36366), .Z(n36371) );
  NANDN U36853 ( .A(n36369), .B(n36368), .Z(n36370) );
  NAND U36854 ( .A(n36371), .B(n36370), .Z(n36504) );
  XNOR U36855 ( .A(n36503), .B(n36504), .Z(n36505) );
  NANDN U36856 ( .A(n36373), .B(n36372), .Z(n36377) );
  OR U36857 ( .A(n36375), .B(n36374), .Z(n36376) );
  NAND U36858 ( .A(n36377), .B(n36376), .Z(n36516) );
  NANDN U36859 ( .A(n36379), .B(n36378), .Z(n36383) );
  OR U36860 ( .A(n36381), .B(n36380), .Z(n36382) );
  NAND U36861 ( .A(n36383), .B(n36382), .Z(n36514) );
  XNOR U36862 ( .A(a[247]), .B(b[13]), .Z(n36563) );
  NANDN U36863 ( .A(n36563), .B(n37424), .Z(n36386) );
  NANDN U36864 ( .A(n36384), .B(n37425), .Z(n36385) );
  NAND U36865 ( .A(n36386), .B(n36385), .Z(n36569) );
  XOR U36866 ( .A(a[245]), .B(n1054), .Z(n36557) );
  OR U36867 ( .A(n36557), .B(n37665), .Z(n36389) );
  NANDN U36868 ( .A(n36387), .B(n37604), .Z(n36388) );
  NAND U36869 ( .A(n36389), .B(n36388), .Z(n36566) );
  NANDN U36870 ( .A(n36390), .B(n37762), .Z(n36392) );
  XNOR U36871 ( .A(b[17]), .B(a[243]), .Z(n36560) );
  NANDN U36872 ( .A(n36560), .B(n37764), .Z(n36391) );
  AND U36873 ( .A(n36392), .B(n36391), .Z(n36567) );
  XNOR U36874 ( .A(n36566), .B(n36567), .Z(n36568) );
  XNOR U36875 ( .A(n36569), .B(n36568), .Z(n36623) );
  NANDN U36876 ( .A(n36394), .B(n36393), .Z(n36398) );
  NANDN U36877 ( .A(n36396), .B(n36395), .Z(n36397) );
  NAND U36878 ( .A(n36398), .B(n36397), .Z(n36621) );
  NANDN U36879 ( .A(n36400), .B(n36399), .Z(n36404) );
  NAND U36880 ( .A(n36402), .B(n36401), .Z(n36403) );
  AND U36881 ( .A(n36404), .B(n36403), .Z(n36620) );
  XNOR U36882 ( .A(n36621), .B(n36620), .Z(n36622) );
  XNOR U36883 ( .A(n36623), .B(n36622), .Z(n36520) );
  NANDN U36884 ( .A(n36406), .B(n36405), .Z(n36410) );
  NANDN U36885 ( .A(n36408), .B(n36407), .Z(n36409) );
  NAND U36886 ( .A(n36410), .B(n36409), .Z(n36517) );
  NANDN U36887 ( .A(n36412), .B(n36411), .Z(n36416) );
  NAND U36888 ( .A(n36414), .B(n36413), .Z(n36415) );
  NAND U36889 ( .A(n36416), .B(n36415), .Z(n36518) );
  XNOR U36890 ( .A(n36517), .B(n36518), .Z(n36519) );
  XNOR U36891 ( .A(n36520), .B(n36519), .Z(n36513) );
  XOR U36892 ( .A(n36514), .B(n36513), .Z(n36515) );
  XNOR U36893 ( .A(n36516), .B(n36515), .Z(n36512) );
  XOR U36894 ( .A(a[249]), .B(b[11]), .Z(n36608) );
  NANDN U36895 ( .A(n37311), .B(n36608), .Z(n36423) );
  NANDN U36896 ( .A(n36421), .B(n37218), .Z(n36422) );
  NAND U36897 ( .A(n36423), .B(n36422), .Z(n36599) );
  XNOR U36898 ( .A(b[25]), .B(a[235]), .Z(n36605) );
  NANDN U36899 ( .A(n36605), .B(n38325), .Z(n36426) );
  NANDN U36900 ( .A(n36424), .B(n38326), .Z(n36425) );
  NAND U36901 ( .A(n36426), .B(n36425), .Z(n36596) );
  XNOR U36902 ( .A(b[27]), .B(a[233]), .Z(n36581) );
  NANDN U36903 ( .A(n36581), .B(n38423), .Z(n36429) );
  NANDN U36904 ( .A(n36427), .B(n38424), .Z(n36428) );
  AND U36905 ( .A(n36429), .B(n36428), .Z(n36597) );
  XNOR U36906 ( .A(n36596), .B(n36597), .Z(n36598) );
  XNOR U36907 ( .A(n36599), .B(n36598), .Z(n36529) );
  XOR U36908 ( .A(a[253]), .B(b[7]), .Z(n36611) );
  NAND U36909 ( .A(n36611), .B(n36701), .Z(n36432) );
  NANDN U36910 ( .A(n36430), .B(n36702), .Z(n36431) );
  NAND U36911 ( .A(n36432), .B(n36431), .Z(n36542) );
  XNOR U36912 ( .A(n1059), .B(a[229]), .Z(n36593) );
  NAND U36913 ( .A(n36593), .B(n38552), .Z(n36435) );
  NANDN U36914 ( .A(n36433), .B(n38553), .Z(n36434) );
  NAND U36915 ( .A(n36435), .B(n36434), .Z(n36539) );
  XNOR U36916 ( .A(b[21]), .B(a[239]), .Z(n36578) );
  NANDN U36917 ( .A(n36578), .B(n38101), .Z(n36438) );
  NANDN U36918 ( .A(n36436), .B(n38102), .Z(n36437) );
  AND U36919 ( .A(n36438), .B(n36437), .Z(n36540) );
  XNOR U36920 ( .A(n36539), .B(n36540), .Z(n36541) );
  XOR U36921 ( .A(n36542), .B(n36541), .Z(n36530) );
  XNOR U36922 ( .A(n36529), .B(n36530), .Z(n36531) );
  NANDN U36923 ( .A(n36440), .B(n36439), .Z(n36444) );
  NAND U36924 ( .A(n36442), .B(n36441), .Z(n36443) );
  AND U36925 ( .A(n36444), .B(n36443), .Z(n36532) );
  XNOR U36926 ( .A(n36531), .B(n36532), .Z(n36536) );
  NANDN U36927 ( .A(n36446), .B(n36445), .Z(n36450) );
  NAND U36928 ( .A(n36448), .B(n36447), .Z(n36449) );
  NAND U36929 ( .A(n36450), .B(n36449), .Z(n36525) );
  NANDN U36930 ( .A(n36451), .B(n38205), .Z(n36453) );
  XNOR U36931 ( .A(b[23]), .B(a[237]), .Z(n36602) );
  OR U36932 ( .A(n36602), .B(n38268), .Z(n36452) );
  NAND U36933 ( .A(n36453), .B(n36452), .Z(n36575) );
  NAND U36934 ( .A(n38490), .B(n36454), .Z(n36456) );
  XOR U36935 ( .A(n1058), .B(n36934), .Z(n36614) );
  NANDN U36936 ( .A(n1048), .B(n36614), .Z(n36455) );
  NAND U36937 ( .A(n36456), .B(n36455), .Z(n36572) );
  XNOR U36938 ( .A(a[251]), .B(b[9]), .Z(n36584) );
  NANDN U36939 ( .A(n36584), .B(n36925), .Z(n36459) );
  NANDN U36940 ( .A(n36457), .B(n36926), .Z(n36458) );
  AND U36941 ( .A(n36459), .B(n36458), .Z(n36573) );
  XNOR U36942 ( .A(n36572), .B(n36573), .Z(n36574) );
  XNOR U36943 ( .A(n36575), .B(n36574), .Z(n36523) );
  ANDN U36944 ( .B(n36460), .A(n1050), .Z(n36552) );
  XNOR U36945 ( .A(n36552), .B(n36551), .Z(n36554) );
  NANDN U36946 ( .A(n1059), .B(a[227]), .Z(n36553) );
  XNOR U36947 ( .A(n36554), .B(n36553), .Z(n36545) );
  XOR U36948 ( .A(n38595), .B(b[5]), .Z(n36589) );
  NANDN U36949 ( .A(n36589), .B(n36587), .Z(n36463) );
  NANDN U36950 ( .A(n36461), .B(n36588), .Z(n36462) );
  NAND U36951 ( .A(n36463), .B(n36462), .Z(n36546) );
  XNOR U36952 ( .A(n36545), .B(n36546), .Z(n36547) );
  XNOR U36953 ( .A(b[19]), .B(a[241]), .Z(n36617) );
  NANDN U36954 ( .A(n36617), .B(n37934), .Z(n36466) );
  NANDN U36955 ( .A(n36464), .B(n37935), .Z(n36465) );
  AND U36956 ( .A(n36466), .B(n36465), .Z(n36548) );
  XNOR U36957 ( .A(n36547), .B(n36548), .Z(n36524) );
  XOR U36958 ( .A(n36523), .B(n36524), .Z(n36526) );
  XOR U36959 ( .A(n36525), .B(n36526), .Z(n36535) );
  XNOR U36960 ( .A(n36536), .B(n36535), .Z(n36537) );
  XNOR U36961 ( .A(n36538), .B(n36537), .Z(n36509) );
  NANDN U36962 ( .A(n36468), .B(n36467), .Z(n36472) );
  OR U36963 ( .A(n36470), .B(n36469), .Z(n36471) );
  NAND U36964 ( .A(n36472), .B(n36471), .Z(n36510) );
  XNOR U36965 ( .A(n36509), .B(n36510), .Z(n36511) );
  XOR U36966 ( .A(n36512), .B(n36511), .Z(n36506) );
  XNOR U36967 ( .A(n36505), .B(n36506), .Z(n36500) );
  NAND U36968 ( .A(n36478), .B(n36477), .Z(n36482) );
  OR U36969 ( .A(n36480), .B(n36479), .Z(n36481) );
  NAND U36970 ( .A(n36482), .B(n36481), .Z(n36498) );
  XNOR U36971 ( .A(n36497), .B(n36498), .Z(n36499) );
  XNOR U36972 ( .A(n36500), .B(n36499), .Z(n36492) );
  NANDN U36973 ( .A(n36484), .B(n36483), .Z(n36488) );
  OR U36974 ( .A(n36486), .B(n36485), .Z(n36487) );
  AND U36975 ( .A(n36488), .B(n36487), .Z(n36491) );
  XNOR U36976 ( .A(n36492), .B(n36491), .Z(n36493) );
  XNOR U36977 ( .A(n36494), .B(n36493), .Z(n36489) );
  XOR U36978 ( .A(n36490), .B(n36489), .Z(c[483]) );
  OR U36979 ( .A(n36490), .B(n36489), .Z(n36758) );
  NANDN U36980 ( .A(n36492), .B(n36491), .Z(n36496) );
  NANDN U36981 ( .A(n36494), .B(n36493), .Z(n36495) );
  NAND U36982 ( .A(n36496), .B(n36495), .Z(n36629) );
  NANDN U36983 ( .A(n36498), .B(n36497), .Z(n36502) );
  NAND U36984 ( .A(n36500), .B(n36499), .Z(n36501) );
  NAND U36985 ( .A(n36502), .B(n36501), .Z(n36626) );
  NANDN U36986 ( .A(n36504), .B(n36503), .Z(n36508) );
  NAND U36987 ( .A(n36506), .B(n36505), .Z(n36507) );
  NAND U36988 ( .A(n36508), .B(n36507), .Z(n36754) );
  NANDN U36989 ( .A(n36518), .B(n36517), .Z(n36522) );
  NANDN U36990 ( .A(n36520), .B(n36519), .Z(n36521) );
  NAND U36991 ( .A(n36522), .B(n36521), .Z(n36742) );
  NANDN U36992 ( .A(n36524), .B(n36523), .Z(n36528) );
  OR U36993 ( .A(n36526), .B(n36525), .Z(n36527) );
  NAND U36994 ( .A(n36528), .B(n36527), .Z(n36739) );
  NANDN U36995 ( .A(n36530), .B(n36529), .Z(n36534) );
  NAND U36996 ( .A(n36532), .B(n36531), .Z(n36533) );
  AND U36997 ( .A(n36534), .B(n36533), .Z(n36740) );
  XNOR U36998 ( .A(n36739), .B(n36740), .Z(n36741) );
  XNOR U36999 ( .A(n36742), .B(n36741), .Z(n36633) );
  XNOR U37000 ( .A(n36632), .B(n36633), .Z(n36634) );
  NANDN U37001 ( .A(n36540), .B(n36539), .Z(n36544) );
  NAND U37002 ( .A(n36542), .B(n36541), .Z(n36543) );
  NAND U37003 ( .A(n36544), .B(n36543), .Z(n36733) );
  NANDN U37004 ( .A(n36546), .B(n36545), .Z(n36550) );
  NAND U37005 ( .A(n36548), .B(n36547), .Z(n36549) );
  NAND U37006 ( .A(n36550), .B(n36549), .Z(n36734) );
  XNOR U37007 ( .A(n36733), .B(n36734), .Z(n36735) );
  OR U37008 ( .A(n36552), .B(n36551), .Z(n36556) );
  OR U37009 ( .A(n36554), .B(n36553), .Z(n36555) );
  AND U37010 ( .A(n36556), .B(n36555), .Z(n36715) );
  XOR U37011 ( .A(a[246]), .B(n1054), .Z(n36683) );
  OR U37012 ( .A(n36683), .B(n37665), .Z(n36559) );
  NANDN U37013 ( .A(n36557), .B(n37604), .Z(n36558) );
  NAND U37014 ( .A(n36559), .B(n36558), .Z(n36668) );
  NANDN U37015 ( .A(n36560), .B(n37762), .Z(n36562) );
  XNOR U37016 ( .A(a[244]), .B(b[17]), .Z(n36689) );
  NANDN U37017 ( .A(n36689), .B(n37764), .Z(n36561) );
  NAND U37018 ( .A(n36562), .B(n36561), .Z(n36665) );
  XOR U37019 ( .A(a[248]), .B(n1053), .Z(n36686) );
  NANDN U37020 ( .A(n36686), .B(n37424), .Z(n36565) );
  NANDN U37021 ( .A(n36563), .B(n37425), .Z(n36564) );
  AND U37022 ( .A(n36565), .B(n36564), .Z(n36666) );
  XNOR U37023 ( .A(n36665), .B(n36666), .Z(n36667) );
  XNOR U37024 ( .A(n36668), .B(n36667), .Z(n36716) );
  XNOR U37025 ( .A(n36715), .B(n36716), .Z(n36717) );
  NANDN U37026 ( .A(n36567), .B(n36566), .Z(n36571) );
  NAND U37027 ( .A(n36569), .B(n36568), .Z(n36570) );
  AND U37028 ( .A(n36571), .B(n36570), .Z(n36718) );
  XOR U37029 ( .A(n36735), .B(n36736), .Z(n36745) );
  NANDN U37030 ( .A(n36573), .B(n36572), .Z(n36577) );
  NAND U37031 ( .A(n36575), .B(n36574), .Z(n36576) );
  NAND U37032 ( .A(n36577), .B(n36576), .Z(n36729) );
  XOR U37033 ( .A(b[21]), .B(n37668), .Z(n36706) );
  NANDN U37034 ( .A(n36706), .B(n38101), .Z(n36580) );
  NANDN U37035 ( .A(n36578), .B(n38102), .Z(n36579) );
  NAND U37036 ( .A(n36580), .B(n36579), .Z(n36674) );
  XNOR U37037 ( .A(b[27]), .B(a[234]), .Z(n36655) );
  NANDN U37038 ( .A(n36655), .B(n38423), .Z(n36583) );
  NANDN U37039 ( .A(n36581), .B(n38424), .Z(n36582) );
  NAND U37040 ( .A(n36583), .B(n36582), .Z(n36671) );
  XOR U37041 ( .A(a[252]), .B(n1052), .Z(n36652) );
  NANDN U37042 ( .A(n36652), .B(n36925), .Z(n36586) );
  NANDN U37043 ( .A(n36584), .B(n36926), .Z(n36585) );
  AND U37044 ( .A(n36586), .B(n36585), .Z(n36672) );
  XNOR U37045 ( .A(n36671), .B(n36672), .Z(n36673) );
  XNOR U37046 ( .A(n36674), .B(n36673), .Z(n36727) );
  NANDN U37047 ( .A(n1051), .B(n36587), .Z(n36591) );
  NANDN U37048 ( .A(n36589), .B(n36588), .Z(n36590) );
  NAND U37049 ( .A(n36591), .B(n36590), .Z(n36644) );
  ANDN U37050 ( .B(b[31]), .A(n36592), .Z(n36658) );
  XNOR U37051 ( .A(n36644), .B(n36658), .Z(n36645) );
  XOR U37052 ( .A(n1059), .B(a[230]), .Z(n36659) );
  NANDN U37053 ( .A(n36659), .B(n38552), .Z(n36595) );
  NAND U37054 ( .A(n38553), .B(n36593), .Z(n36594) );
  AND U37055 ( .A(n36595), .B(n36594), .Z(n36646) );
  XNOR U37056 ( .A(n36645), .B(n36646), .Z(n36728) );
  XOR U37057 ( .A(n36727), .B(n36728), .Z(n36730) );
  XNOR U37058 ( .A(n36729), .B(n36730), .Z(n36638) );
  NANDN U37059 ( .A(n36597), .B(n36596), .Z(n36601) );
  NAND U37060 ( .A(n36599), .B(n36598), .Z(n36600) );
  NAND U37061 ( .A(n36601), .B(n36600), .Z(n36723) );
  NANDN U37062 ( .A(n36602), .B(n38205), .Z(n36604) );
  XOR U37063 ( .A(b[23]), .B(n37467), .Z(n36649) );
  OR U37064 ( .A(n36649), .B(n38268), .Z(n36603) );
  NAND U37065 ( .A(n36604), .B(n36603), .Z(n36680) );
  XNOR U37066 ( .A(b[25]), .B(a[236]), .Z(n36692) );
  NANDN U37067 ( .A(n36692), .B(n38325), .Z(n36607) );
  NANDN U37068 ( .A(n36605), .B(n38326), .Z(n36606) );
  NAND U37069 ( .A(n36607), .B(n36606), .Z(n36677) );
  XNOR U37070 ( .A(a[250]), .B(b[11]), .Z(n36695) );
  OR U37071 ( .A(n36695), .B(n37311), .Z(n36610) );
  NAND U37072 ( .A(n36608), .B(n37218), .Z(n36609) );
  AND U37073 ( .A(n36610), .B(n36609), .Z(n36678) );
  XNOR U37074 ( .A(n36677), .B(n36678), .Z(n36679) );
  XNOR U37075 ( .A(n36680), .B(n36679), .Z(n36721) );
  XNOR U37076 ( .A(a[254]), .B(b[7]), .Z(n36703) );
  NANDN U37077 ( .A(n36703), .B(n36701), .Z(n36613) );
  NAND U37078 ( .A(n36611), .B(n36702), .Z(n36612) );
  NAND U37079 ( .A(n36613), .B(n36612), .Z(n36712) );
  NAND U37080 ( .A(n38490), .B(n36614), .Z(n36616) );
  XOR U37081 ( .A(n1058), .B(n37079), .Z(n36698) );
  NANDN U37082 ( .A(n1048), .B(n36698), .Z(n36615) );
  NAND U37083 ( .A(n36616), .B(n36615), .Z(n36709) );
  XOR U37084 ( .A(n1055), .B(n37676), .Z(n36662) );
  NAND U37085 ( .A(n36662), .B(n37934), .Z(n36619) );
  NANDN U37086 ( .A(n36617), .B(n37935), .Z(n36618) );
  AND U37087 ( .A(n36619), .B(n36618), .Z(n36710) );
  XNOR U37088 ( .A(n36709), .B(n36710), .Z(n36711) );
  XOR U37089 ( .A(n36712), .B(n36711), .Z(n36722) );
  XOR U37090 ( .A(n36721), .B(n36722), .Z(n36724) );
  XOR U37091 ( .A(n36723), .B(n36724), .Z(n36639) );
  XNOR U37092 ( .A(n36638), .B(n36639), .Z(n36640) );
  NANDN U37093 ( .A(n36621), .B(n36620), .Z(n36625) );
  NAND U37094 ( .A(n36623), .B(n36622), .Z(n36624) );
  NAND U37095 ( .A(n36625), .B(n36624), .Z(n36641) );
  XNOR U37096 ( .A(n36640), .B(n36641), .Z(n36746) );
  XNOR U37097 ( .A(n36745), .B(n36746), .Z(n36747) );
  XNOR U37098 ( .A(n36748), .B(n36747), .Z(n36635) );
  XNOR U37099 ( .A(n36634), .B(n36635), .Z(n36752) );
  XNOR U37100 ( .A(n36751), .B(n36752), .Z(n36753) );
  XOR U37101 ( .A(n36754), .B(n36753), .Z(n36627) );
  XNOR U37102 ( .A(n36626), .B(n36627), .Z(n36628) );
  XOR U37103 ( .A(n36629), .B(n36628), .Z(n36757) );
  XOR U37104 ( .A(n36758), .B(n36757), .Z(c[484]) );
  NANDN U37105 ( .A(n36627), .B(n36626), .Z(n36631) );
  NAND U37106 ( .A(n36629), .B(n36628), .Z(n36630) );
  NAND U37107 ( .A(n36631), .B(n36630), .Z(n36763) );
  NANDN U37108 ( .A(n36633), .B(n36632), .Z(n36637) );
  NANDN U37109 ( .A(n36635), .B(n36634), .Z(n36636) );
  NAND U37110 ( .A(n36637), .B(n36636), .Z(n36882) );
  NANDN U37111 ( .A(n36639), .B(n36638), .Z(n36643) );
  NANDN U37112 ( .A(n36641), .B(n36640), .Z(n36642) );
  NAND U37113 ( .A(n36643), .B(n36642), .Z(n36878) );
  IV U37114 ( .A(n36658), .Z(n36863) );
  OR U37115 ( .A(n36644), .B(n36863), .Z(n36648) );
  NAND U37116 ( .A(n36646), .B(n36645), .Z(n36647) );
  NAND U37117 ( .A(n36648), .B(n36647), .Z(n36790) );
  NANDN U37118 ( .A(n36649), .B(n38205), .Z(n36651) );
  XNOR U37119 ( .A(n1057), .B(a[239]), .Z(n36817) );
  NANDN U37120 ( .A(n38268), .B(n36817), .Z(n36650) );
  NAND U37121 ( .A(n36651), .B(n36650), .Z(n36857) );
  XNOR U37122 ( .A(a[253]), .B(b[9]), .Z(n36826) );
  NANDN U37123 ( .A(n36826), .B(n36925), .Z(n36654) );
  NANDN U37124 ( .A(n36652), .B(n36926), .Z(n36653) );
  NAND U37125 ( .A(n36654), .B(n36653), .Z(n36854) );
  XNOR U37126 ( .A(b[27]), .B(a[235]), .Z(n36805) );
  NANDN U37127 ( .A(n36805), .B(n38423), .Z(n36657) );
  NANDN U37128 ( .A(n36655), .B(n38424), .Z(n36656) );
  AND U37129 ( .A(n36657), .B(n36656), .Z(n36855) );
  XNOR U37130 ( .A(n36854), .B(n36855), .Z(n36856) );
  XNOR U37131 ( .A(n36857), .B(n36856), .Z(n36787) );
  NANDN U37132 ( .A(n1059), .B(a[229]), .Z(n36860) );
  XOR U37133 ( .A(n36861), .B(n36860), .Z(n36862) );
  XOR U37134 ( .A(n36658), .B(n36862), .Z(n36794) );
  XOR U37135 ( .A(n1059), .B(a[231]), .Z(n36833) );
  NANDN U37136 ( .A(n36833), .B(n38552), .Z(n36661) );
  NANDN U37137 ( .A(n36659), .B(n38553), .Z(n36660) );
  NAND U37138 ( .A(n36661), .B(n36660), .Z(n36793) );
  XOR U37139 ( .A(n36794), .B(n36793), .Z(n36795) );
  XOR U37140 ( .A(n1055), .B(a[243]), .Z(n36814) );
  NANDN U37141 ( .A(n36814), .B(n37934), .Z(n36664) );
  NAND U37142 ( .A(n37935), .B(n36662), .Z(n36663) );
  AND U37143 ( .A(n36664), .B(n36663), .Z(n36796) );
  XNOR U37144 ( .A(n36795), .B(n36796), .Z(n36788) );
  XNOR U37145 ( .A(n36787), .B(n36788), .Z(n36789) );
  XNOR U37146 ( .A(n36790), .B(n36789), .Z(n36839) );
  NANDN U37147 ( .A(n36666), .B(n36665), .Z(n36670) );
  NAND U37148 ( .A(n36668), .B(n36667), .Z(n36669) );
  NAND U37149 ( .A(n36670), .B(n36669), .Z(n36837) );
  NANDN U37150 ( .A(n36672), .B(n36671), .Z(n36676) );
  NAND U37151 ( .A(n36674), .B(n36673), .Z(n36675) );
  AND U37152 ( .A(n36676), .B(n36675), .Z(n36836) );
  XNOR U37153 ( .A(n36837), .B(n36836), .Z(n36838) );
  XNOR U37154 ( .A(n36839), .B(n36838), .Z(n36781) );
  NANDN U37155 ( .A(n36678), .B(n36677), .Z(n36682) );
  NAND U37156 ( .A(n36680), .B(n36679), .Z(n36681) );
  NAND U37157 ( .A(n36682), .B(n36681), .Z(n36780) );
  XNOR U37158 ( .A(a[247]), .B(b[15]), .Z(n36866) );
  OR U37159 ( .A(n36866), .B(n37665), .Z(n36685) );
  NANDN U37160 ( .A(n36683), .B(n37604), .Z(n36684) );
  NAND U37161 ( .A(n36685), .B(n36684), .Z(n36845) );
  XNOR U37162 ( .A(a[249]), .B(b[13]), .Z(n36869) );
  NANDN U37163 ( .A(n36869), .B(n37424), .Z(n36688) );
  NANDN U37164 ( .A(n36686), .B(n37425), .Z(n36687) );
  NAND U37165 ( .A(n36688), .B(n36687), .Z(n36842) );
  NANDN U37166 ( .A(n36689), .B(n37762), .Z(n36691) );
  XNOR U37167 ( .A(a[245]), .B(b[17]), .Z(n36811) );
  NANDN U37168 ( .A(n36811), .B(n37764), .Z(n36690) );
  NAND U37169 ( .A(n36691), .B(n36690), .Z(n36802) );
  XOR U37170 ( .A(b[25]), .B(a[237]), .Z(n36872) );
  NAND U37171 ( .A(n36872), .B(n38325), .Z(n36694) );
  NANDN U37172 ( .A(n36692), .B(n38326), .Z(n36693) );
  NAND U37173 ( .A(n36694), .B(n36693), .Z(n36799) );
  XOR U37174 ( .A(a[251]), .B(b[11]), .Z(n36823) );
  NANDN U37175 ( .A(n37311), .B(n36823), .Z(n36697) );
  NANDN U37176 ( .A(n36695), .B(n37218), .Z(n36696) );
  AND U37177 ( .A(n36697), .B(n36696), .Z(n36800) );
  XNOR U37178 ( .A(n36799), .B(n36800), .Z(n36801) );
  XNOR U37179 ( .A(n36802), .B(n36801), .Z(n36843) );
  XNOR U37180 ( .A(n36842), .B(n36843), .Z(n36844) );
  XNOR U37181 ( .A(n36845), .B(n36844), .Z(n36786) );
  NAND U37182 ( .A(n38490), .B(n36698), .Z(n36700) );
  XOR U37183 ( .A(n1058), .B(n37184), .Z(n36808) );
  NANDN U37184 ( .A(n1048), .B(n36808), .Z(n36699) );
  NAND U37185 ( .A(n36700), .B(n36699), .Z(n36851) );
  XNOR U37186 ( .A(n38595), .B(b[7]), .Z(n36830) );
  NAND U37187 ( .A(n36830), .B(n36701), .Z(n36705) );
  NANDN U37188 ( .A(n36703), .B(n36702), .Z(n36704) );
  NAND U37189 ( .A(n36705), .B(n36704), .Z(n36848) );
  XNOR U37190 ( .A(b[21]), .B(a[241]), .Z(n36820) );
  NANDN U37191 ( .A(n36820), .B(n38101), .Z(n36708) );
  NANDN U37192 ( .A(n36706), .B(n38102), .Z(n36707) );
  AND U37193 ( .A(n36708), .B(n36707), .Z(n36849) );
  XNOR U37194 ( .A(n36848), .B(n36849), .Z(n36850) );
  XNOR U37195 ( .A(n36851), .B(n36850), .Z(n36783) );
  NANDN U37196 ( .A(n36710), .B(n36709), .Z(n36714) );
  NAND U37197 ( .A(n36712), .B(n36711), .Z(n36713) );
  NAND U37198 ( .A(n36714), .B(n36713), .Z(n36784) );
  XNOR U37199 ( .A(n36783), .B(n36784), .Z(n36785) );
  XOR U37200 ( .A(n36786), .B(n36785), .Z(n36779) );
  XOR U37201 ( .A(n36780), .B(n36779), .Z(n36782) );
  XOR U37202 ( .A(n36781), .B(n36782), .Z(n36875) );
  OR U37203 ( .A(n36716), .B(n36715), .Z(n36720) );
  OR U37204 ( .A(n36718), .B(n36717), .Z(n36719) );
  AND U37205 ( .A(n36720), .B(n36719), .Z(n36876) );
  XNOR U37206 ( .A(n36875), .B(n36876), .Z(n36877) );
  XNOR U37207 ( .A(n36878), .B(n36877), .Z(n36879) );
  NANDN U37208 ( .A(n36722), .B(n36721), .Z(n36726) );
  OR U37209 ( .A(n36724), .B(n36723), .Z(n36725) );
  NAND U37210 ( .A(n36726), .B(n36725), .Z(n36773) );
  NANDN U37211 ( .A(n36728), .B(n36727), .Z(n36732) );
  OR U37212 ( .A(n36730), .B(n36729), .Z(n36731) );
  AND U37213 ( .A(n36732), .B(n36731), .Z(n36774) );
  XNOR U37214 ( .A(n36773), .B(n36774), .Z(n36775) );
  NANDN U37215 ( .A(n36734), .B(n36733), .Z(n36738) );
  NANDN U37216 ( .A(n36736), .B(n36735), .Z(n36737) );
  NAND U37217 ( .A(n36738), .B(n36737), .Z(n36776) );
  XOR U37218 ( .A(n36775), .B(n36776), .Z(n36767) );
  NANDN U37219 ( .A(n36740), .B(n36739), .Z(n36744) );
  NAND U37220 ( .A(n36742), .B(n36741), .Z(n36743) );
  NAND U37221 ( .A(n36744), .B(n36743), .Z(n36768) );
  XNOR U37222 ( .A(n36767), .B(n36768), .Z(n36769) );
  NANDN U37223 ( .A(n36746), .B(n36745), .Z(n36750) );
  NAND U37224 ( .A(n36748), .B(n36747), .Z(n36749) );
  NAND U37225 ( .A(n36750), .B(n36749), .Z(n36770) );
  XNOR U37226 ( .A(n36769), .B(n36770), .Z(n36880) );
  XNOR U37227 ( .A(n36879), .B(n36880), .Z(n36881) );
  XNOR U37228 ( .A(n36882), .B(n36881), .Z(n36761) );
  NANDN U37229 ( .A(n36752), .B(n36751), .Z(n36756) );
  NAND U37230 ( .A(n36754), .B(n36753), .Z(n36755) );
  AND U37231 ( .A(n36756), .B(n36755), .Z(n36762) );
  XOR U37232 ( .A(n36761), .B(n36762), .Z(n36764) );
  XOR U37233 ( .A(n36763), .B(n36764), .Z(n36759) );
  OR U37234 ( .A(n36758), .B(n36757), .Z(n36760) );
  XNOR U37235 ( .A(n36759), .B(n36760), .Z(c[485]) );
  NANDN U37236 ( .A(n36760), .B(n36759), .Z(n36885) );
  NANDN U37237 ( .A(n36762), .B(n36761), .Z(n36766) );
  OR U37238 ( .A(n36764), .B(n36763), .Z(n36765) );
  NAND U37239 ( .A(n36766), .B(n36765), .Z(n37003) );
  NANDN U37240 ( .A(n36768), .B(n36767), .Z(n36772) );
  NANDN U37241 ( .A(n36770), .B(n36769), .Z(n36771) );
  NAND U37242 ( .A(n36772), .B(n36771), .Z(n36889) );
  NANDN U37243 ( .A(n36774), .B(n36773), .Z(n36778) );
  NANDN U37244 ( .A(n36776), .B(n36775), .Z(n36777) );
  NAND U37245 ( .A(n36778), .B(n36777), .Z(n36894) );
  NANDN U37246 ( .A(n36788), .B(n36787), .Z(n36792) );
  NAND U37247 ( .A(n36790), .B(n36789), .Z(n36791) );
  NAND U37248 ( .A(n36792), .B(n36791), .Z(n36978) );
  OR U37249 ( .A(n36794), .B(n36793), .Z(n36798) );
  NAND U37250 ( .A(n36796), .B(n36795), .Z(n36797) );
  NAND U37251 ( .A(n36798), .B(n36797), .Z(n36983) );
  NANDN U37252 ( .A(n36800), .B(n36799), .Z(n36804) );
  NAND U37253 ( .A(n36802), .B(n36801), .Z(n36803) );
  NAND U37254 ( .A(n36804), .B(n36803), .Z(n36984) );
  XNOR U37255 ( .A(n36983), .B(n36984), .Z(n36985) );
  XNOR U37256 ( .A(b[27]), .B(a[236]), .Z(n36953) );
  NANDN U37257 ( .A(n36953), .B(n38423), .Z(n36807) );
  NANDN U37258 ( .A(n36805), .B(n38424), .Z(n36806) );
  NAND U37259 ( .A(n36807), .B(n36806), .Z(n36911) );
  NAND U37260 ( .A(n38490), .B(n36808), .Z(n36810) );
  XOR U37261 ( .A(n1058), .B(n37080), .Z(n36935) );
  NANDN U37262 ( .A(n1048), .B(n36935), .Z(n36809) );
  NAND U37263 ( .A(n36810), .B(n36809), .Z(n36908) );
  NANDN U37264 ( .A(n36811), .B(n37762), .Z(n36813) );
  XNOR U37265 ( .A(a[246]), .B(b[17]), .Z(n36965) );
  NANDN U37266 ( .A(n36965), .B(n37764), .Z(n36812) );
  AND U37267 ( .A(n36813), .B(n36812), .Z(n36909) );
  XNOR U37268 ( .A(n36908), .B(n36909), .Z(n36910) );
  XNOR U37269 ( .A(n36911), .B(n36910), .Z(n36974) );
  XOR U37270 ( .A(n38034), .B(b[19]), .Z(n36962) );
  NANDN U37271 ( .A(n36962), .B(n37934), .Z(n36816) );
  NANDN U37272 ( .A(n36814), .B(n37935), .Z(n36815) );
  NAND U37273 ( .A(n36816), .B(n36815), .Z(n36972) );
  XOR U37274 ( .A(b[23]), .B(n37668), .Z(n36941) );
  OR U37275 ( .A(n36941), .B(n38268), .Z(n36819) );
  NAND U37276 ( .A(n38205), .B(n36817), .Z(n36818) );
  AND U37277 ( .A(n36819), .B(n36818), .Z(n36971) );
  XNOR U37278 ( .A(n36972), .B(n36971), .Z(n36973) );
  XOR U37279 ( .A(n36974), .B(n36973), .Z(n36997) );
  XOR U37280 ( .A(b[21]), .B(n37676), .Z(n36930) );
  NANDN U37281 ( .A(n36930), .B(n38101), .Z(n36822) );
  NANDN U37282 ( .A(n36820), .B(n38102), .Z(n36821) );
  NAND U37283 ( .A(n36822), .B(n36821), .Z(n36917) );
  XNOR U37284 ( .A(a[252]), .B(b[11]), .Z(n36956) );
  OR U37285 ( .A(n36956), .B(n37311), .Z(n36825) );
  NAND U37286 ( .A(n36823), .B(n37218), .Z(n36824) );
  NAND U37287 ( .A(n36825), .B(n36824), .Z(n36914) );
  XOR U37288 ( .A(a[254]), .B(n1052), .Z(n36927) );
  NANDN U37289 ( .A(n36927), .B(n36925), .Z(n36828) );
  NANDN U37290 ( .A(n36826), .B(n36926), .Z(n36827) );
  AND U37291 ( .A(n36828), .B(n36827), .Z(n36915) );
  XNOR U37292 ( .A(n36914), .B(n36915), .Z(n36916) );
  XNOR U37293 ( .A(n36917), .B(n36916), .Z(n36995) );
  NANDN U37294 ( .A(n1051), .B(b[6]), .Z(n36933) );
  XNOR U37295 ( .A(b[7]), .B(n36933), .Z(n36832) );
  XOR U37296 ( .A(b[6]), .B(n1051), .Z(n36829) );
  NANDN U37297 ( .A(n36830), .B(n36829), .Z(n36831) );
  AND U37298 ( .A(n36832), .B(n36831), .Z(n36920) );
  AND U37299 ( .A(a[230]), .B(b[31]), .Z(n37086) );
  XNOR U37300 ( .A(n36920), .B(n37086), .Z(n36921) );
  XOR U37301 ( .A(b[31]), .B(n37079), .Z(n36938) );
  NANDN U37302 ( .A(n36938), .B(n38552), .Z(n36835) );
  NANDN U37303 ( .A(n36833), .B(n38553), .Z(n36834) );
  AND U37304 ( .A(n36835), .B(n36834), .Z(n36922) );
  XNOR U37305 ( .A(n36921), .B(n36922), .Z(n36996) );
  XOR U37306 ( .A(n36995), .B(n36996), .Z(n36998) );
  XNOR U37307 ( .A(n36997), .B(n36998), .Z(n36986) );
  XOR U37308 ( .A(n36985), .B(n36986), .Z(n36977) );
  XOR U37309 ( .A(n36978), .B(n36977), .Z(n36979) );
  XNOR U37310 ( .A(n36980), .B(n36979), .Z(n36901) );
  NANDN U37311 ( .A(n36837), .B(n36836), .Z(n36841) );
  NANDN U37312 ( .A(n36839), .B(n36838), .Z(n36840) );
  NAND U37313 ( .A(n36841), .B(n36840), .Z(n36899) );
  NANDN U37314 ( .A(n36843), .B(n36842), .Z(n36847) );
  NAND U37315 ( .A(n36845), .B(n36844), .Z(n36846) );
  NAND U37316 ( .A(n36847), .B(n36846), .Z(n36904) );
  NANDN U37317 ( .A(n36849), .B(n36848), .Z(n36853) );
  NAND U37318 ( .A(n36851), .B(n36850), .Z(n36852) );
  NAND U37319 ( .A(n36853), .B(n36852), .Z(n36903) );
  NANDN U37320 ( .A(n36855), .B(n36854), .Z(n36859) );
  NAND U37321 ( .A(n36857), .B(n36856), .Z(n36858) );
  NAND U37322 ( .A(n36859), .B(n36858), .Z(n36989) );
  OR U37323 ( .A(n36861), .B(n36860), .Z(n36865) );
  NANDN U37324 ( .A(n36863), .B(n36862), .Z(n36864) );
  AND U37325 ( .A(n36865), .B(n36864), .Z(n36990) );
  XNOR U37326 ( .A(n36989), .B(n36990), .Z(n36991) );
  XOR U37327 ( .A(a[248]), .B(n1054), .Z(n36968) );
  OR U37328 ( .A(n36968), .B(n37665), .Z(n36868) );
  NANDN U37329 ( .A(n36866), .B(n37604), .Z(n36867) );
  NAND U37330 ( .A(n36868), .B(n36867), .Z(n36947) );
  XOR U37331 ( .A(n38356), .B(n1053), .Z(n36959) );
  NAND U37332 ( .A(n36959), .B(n37424), .Z(n36871) );
  NANDN U37333 ( .A(n36869), .B(n37425), .Z(n36870) );
  NAND U37334 ( .A(n36871), .B(n36870), .Z(n36944) );
  XNOR U37335 ( .A(b[25]), .B(a[238]), .Z(n36950) );
  NANDN U37336 ( .A(n36950), .B(n38325), .Z(n36874) );
  NAND U37337 ( .A(n36872), .B(n38326), .Z(n36873) );
  AND U37338 ( .A(n36874), .B(n36873), .Z(n36945) );
  XNOR U37339 ( .A(n36944), .B(n36945), .Z(n36946) );
  XOR U37340 ( .A(n36947), .B(n36946), .Z(n36992) );
  XOR U37341 ( .A(n36991), .B(n36992), .Z(n36902) );
  XNOR U37342 ( .A(n36903), .B(n36902), .Z(n36905) );
  XNOR U37343 ( .A(n36904), .B(n36905), .Z(n36898) );
  XNOR U37344 ( .A(n36899), .B(n36898), .Z(n36900) );
  XOR U37345 ( .A(n36901), .B(n36900), .Z(n36892) );
  XOR U37346 ( .A(n36893), .B(n36892), .Z(n36895) );
  XNOR U37347 ( .A(n36894), .B(n36895), .Z(n36887) );
  XOR U37348 ( .A(n36887), .B(n36886), .Z(n36888) );
  XOR U37349 ( .A(n36889), .B(n36888), .Z(n37001) );
  XOR U37350 ( .A(n37001), .B(n37002), .Z(n36883) );
  XOR U37351 ( .A(n37003), .B(n36883), .Z(n36884) );
  XNOR U37352 ( .A(n36885), .B(n36884), .Z(c[486]) );
  NANDN U37353 ( .A(n36885), .B(n36884), .Z(n37125) );
  NAND U37354 ( .A(n36887), .B(n36886), .Z(n36891) );
  NANDN U37355 ( .A(n36889), .B(n36888), .Z(n36890) );
  NAND U37356 ( .A(n36891), .B(n36890), .Z(n37006) );
  NANDN U37357 ( .A(n36893), .B(n36892), .Z(n36897) );
  OR U37358 ( .A(n36895), .B(n36894), .Z(n36896) );
  NAND U37359 ( .A(n36897), .B(n36896), .Z(n37011) );
  NAND U37360 ( .A(n36903), .B(n36902), .Z(n36907) );
  NANDN U37361 ( .A(n36905), .B(n36904), .Z(n36906) );
  NAND U37362 ( .A(n36907), .B(n36906), .Z(n37121) );
  NANDN U37363 ( .A(n36909), .B(n36908), .Z(n36913) );
  NAND U37364 ( .A(n36911), .B(n36910), .Z(n36912) );
  NAND U37365 ( .A(n36913), .B(n36912), .Z(n37026) );
  NANDN U37366 ( .A(n36915), .B(n36914), .Z(n36919) );
  NAND U37367 ( .A(n36917), .B(n36916), .Z(n36918) );
  AND U37368 ( .A(n36919), .B(n36918), .Z(n37027) );
  XNOR U37369 ( .A(n37026), .B(n37027), .Z(n37028) );
  NANDN U37370 ( .A(n36920), .B(n37086), .Z(n36924) );
  NAND U37371 ( .A(n36922), .B(n36921), .Z(n36923) );
  NAND U37372 ( .A(n36924), .B(n36923), .Z(n37035) );
  XNOR U37373 ( .A(n38595), .B(b[9]), .Z(n37076) );
  NAND U37374 ( .A(n36925), .B(n37076), .Z(n36929) );
  NANDN U37375 ( .A(n36927), .B(n36926), .Z(n36928) );
  NAND U37376 ( .A(n36929), .B(n36928), .Z(n37112) );
  XOR U37377 ( .A(n1056), .B(n38110), .Z(n37109) );
  NAND U37378 ( .A(n37109), .B(n38101), .Z(n36932) );
  NANDN U37379 ( .A(n36930), .B(n38102), .Z(n36931) );
  AND U37380 ( .A(n36932), .B(n36931), .Z(n37113) );
  XNOR U37381 ( .A(n37112), .B(n37113), .Z(n37114) );
  AND U37382 ( .A(n36933), .B(b[7]), .Z(n37085) );
  NANDN U37383 ( .A(n36934), .B(b[31]), .Z(n37084) );
  XOR U37384 ( .A(n37085), .B(n37084), .Z(n37087) );
  XNOR U37385 ( .A(n37086), .B(n37087), .Z(n37115) );
  XNOR U37386 ( .A(n37114), .B(n37115), .Z(n37032) );
  NAND U37387 ( .A(n38490), .B(n36935), .Z(n36937) );
  XOR U37388 ( .A(b[29]), .B(n37420), .Z(n37105) );
  OR U37389 ( .A(n37105), .B(n1048), .Z(n36936) );
  NAND U37390 ( .A(n36937), .B(n36936), .Z(n37093) );
  XOR U37391 ( .A(b[31]), .B(n37184), .Z(n37081) );
  NANDN U37392 ( .A(n37081), .B(n38552), .Z(n36940) );
  NANDN U37393 ( .A(n36938), .B(n38553), .Z(n36939) );
  NAND U37394 ( .A(n36940), .B(n36939), .Z(n37090) );
  NANDN U37395 ( .A(n36941), .B(n38205), .Z(n36943) );
  XNOR U37396 ( .A(n1057), .B(a[241]), .Z(n37048) );
  NANDN U37397 ( .A(n38268), .B(n37048), .Z(n36942) );
  AND U37398 ( .A(n36943), .B(n36942), .Z(n37091) );
  XNOR U37399 ( .A(n37090), .B(n37091), .Z(n37092) );
  XOR U37400 ( .A(n37093), .B(n37092), .Z(n37033) );
  XOR U37401 ( .A(n37032), .B(n37033), .Z(n37034) );
  XOR U37402 ( .A(n37035), .B(n37034), .Z(n37029) );
  XOR U37403 ( .A(n37028), .B(n37029), .Z(n37119) );
  NANDN U37404 ( .A(n36945), .B(n36944), .Z(n36949) );
  NAND U37405 ( .A(n36947), .B(n36946), .Z(n36948) );
  NAND U37406 ( .A(n36949), .B(n36948), .Z(n37042) );
  XOR U37407 ( .A(b[25]), .B(a[239]), .Z(n37054) );
  NAND U37408 ( .A(n37054), .B(n38325), .Z(n36952) );
  NANDN U37409 ( .A(n36950), .B(n38326), .Z(n36951) );
  NAND U37410 ( .A(n36952), .B(n36951), .Z(n37072) );
  XOR U37411 ( .A(b[27]), .B(a[237]), .Z(n37051) );
  NAND U37412 ( .A(n38423), .B(n37051), .Z(n36955) );
  NANDN U37413 ( .A(n36953), .B(n38424), .Z(n36954) );
  NAND U37414 ( .A(n36955), .B(n36954), .Z(n37069) );
  XOR U37415 ( .A(a[253]), .B(b[11]), .Z(n37102) );
  NANDN U37416 ( .A(n37311), .B(n37102), .Z(n36958) );
  NANDN U37417 ( .A(n36956), .B(n37218), .Z(n36957) );
  AND U37418 ( .A(n36958), .B(n36957), .Z(n37070) );
  XNOR U37419 ( .A(n37069), .B(n37070), .Z(n37071) );
  XNOR U37420 ( .A(n37072), .B(n37071), .Z(n37039) );
  XOR U37421 ( .A(a[251]), .B(n1053), .Z(n37060) );
  NANDN U37422 ( .A(n37060), .B(n37424), .Z(n36961) );
  NAND U37423 ( .A(n37425), .B(n36959), .Z(n36960) );
  NAND U37424 ( .A(n36961), .B(n36960), .Z(n37097) );
  XOR U37425 ( .A(b[19]), .B(n38213), .Z(n37063) );
  NANDN U37426 ( .A(n37063), .B(n37934), .Z(n36964) );
  NANDN U37427 ( .A(n36962), .B(n37935), .Z(n36963) );
  AND U37428 ( .A(n36964), .B(n36963), .Z(n37096) );
  XNOR U37429 ( .A(n37097), .B(n37096), .Z(n37098) );
  XOR U37430 ( .A(a[247]), .B(b[17]), .Z(n37057) );
  NAND U37431 ( .A(n37764), .B(n37057), .Z(n36967) );
  NANDN U37432 ( .A(n36965), .B(n37762), .Z(n36966) );
  AND U37433 ( .A(n36967), .B(n36966), .Z(n37099) );
  XNOR U37434 ( .A(n37098), .B(n37099), .Z(n37037) );
  XNOR U37435 ( .A(a[249]), .B(b[15]), .Z(n37066) );
  OR U37436 ( .A(n37066), .B(n37665), .Z(n36970) );
  NANDN U37437 ( .A(n36968), .B(n37604), .Z(n36969) );
  AND U37438 ( .A(n36970), .B(n36969), .Z(n37036) );
  XNOR U37439 ( .A(n37037), .B(n37036), .Z(n37038) );
  XOR U37440 ( .A(n37039), .B(n37038), .Z(n37043) );
  XNOR U37441 ( .A(n37042), .B(n37043), .Z(n37044) );
  NANDN U37442 ( .A(n36972), .B(n36971), .Z(n36976) );
  NAND U37443 ( .A(n36974), .B(n36973), .Z(n36975) );
  AND U37444 ( .A(n36976), .B(n36975), .Z(n37045) );
  XNOR U37445 ( .A(n37044), .B(n37045), .Z(n37118) );
  XOR U37446 ( .A(n37119), .B(n37118), .Z(n37120) );
  XOR U37447 ( .A(n37121), .B(n37120), .Z(n37017) );
  NAND U37448 ( .A(n36978), .B(n36977), .Z(n36982) );
  NAND U37449 ( .A(n36980), .B(n36979), .Z(n36981) );
  NAND U37450 ( .A(n36982), .B(n36981), .Z(n37014) );
  NANDN U37451 ( .A(n36984), .B(n36983), .Z(n36988) );
  NAND U37452 ( .A(n36986), .B(n36985), .Z(n36987) );
  NAND U37453 ( .A(n36988), .B(n36987), .Z(n37023) );
  NANDN U37454 ( .A(n36990), .B(n36989), .Z(n36994) );
  NAND U37455 ( .A(n36992), .B(n36991), .Z(n36993) );
  NAND U37456 ( .A(n36994), .B(n36993), .Z(n37020) );
  NANDN U37457 ( .A(n36996), .B(n36995), .Z(n37000) );
  NANDN U37458 ( .A(n36998), .B(n36997), .Z(n36999) );
  NAND U37459 ( .A(n37000), .B(n36999), .Z(n37021) );
  XNOR U37460 ( .A(n37020), .B(n37021), .Z(n37022) );
  XOR U37461 ( .A(n37023), .B(n37022), .Z(n37015) );
  XOR U37462 ( .A(n37014), .B(n37015), .Z(n37016) );
  XNOR U37463 ( .A(n37017), .B(n37016), .Z(n37009) );
  XNOR U37464 ( .A(n37008), .B(n37009), .Z(n37010) );
  XNOR U37465 ( .A(n37011), .B(n37010), .Z(n37005) );
  XNOR U37466 ( .A(n37005), .B(n37007), .Z(n37004) );
  XNOR U37467 ( .A(n37006), .B(n37004), .Z(n37124) );
  XNOR U37468 ( .A(n37125), .B(n37124), .Z(c[487]) );
  NANDN U37469 ( .A(n37009), .B(n37008), .Z(n37013) );
  NAND U37470 ( .A(n37011), .B(n37010), .Z(n37012) );
  NAND U37471 ( .A(n37013), .B(n37012), .Z(n37128) );
  OR U37472 ( .A(n37015), .B(n37014), .Z(n37019) );
  NAND U37473 ( .A(n37017), .B(n37016), .Z(n37018) );
  NAND U37474 ( .A(n37019), .B(n37018), .Z(n37234) );
  NANDN U37475 ( .A(n37021), .B(n37020), .Z(n37025) );
  NANDN U37476 ( .A(n37023), .B(n37022), .Z(n37024) );
  NAND U37477 ( .A(n37025), .B(n37024), .Z(n37134) );
  NANDN U37478 ( .A(n37027), .B(n37026), .Z(n37031) );
  NANDN U37479 ( .A(n37029), .B(n37028), .Z(n37030) );
  NAND U37480 ( .A(n37031), .B(n37030), .Z(n37228) );
  NANDN U37481 ( .A(n37037), .B(n37036), .Z(n37041) );
  NAND U37482 ( .A(n37039), .B(n37038), .Z(n37040) );
  NAND U37483 ( .A(n37041), .B(n37040), .Z(n37226) );
  XNOR U37484 ( .A(n37225), .B(n37226), .Z(n37227) );
  XNOR U37485 ( .A(n37228), .B(n37227), .Z(n37135) );
  XNOR U37486 ( .A(n37134), .B(n37135), .Z(n37136) );
  NANDN U37487 ( .A(n37043), .B(n37042), .Z(n37047) );
  NAND U37488 ( .A(n37045), .B(n37044), .Z(n37046) );
  NAND U37489 ( .A(n37047), .B(n37046), .Z(n37143) );
  XOR U37490 ( .A(n1057), .B(a[242]), .Z(n37222) );
  OR U37491 ( .A(n37222), .B(n38268), .Z(n37050) );
  NAND U37492 ( .A(n38205), .B(n37048), .Z(n37049) );
  NAND U37493 ( .A(n37050), .B(n37049), .Z(n37192) );
  XNOR U37494 ( .A(b[27]), .B(n37467), .Z(n37177) );
  NAND U37495 ( .A(n38423), .B(n37177), .Z(n37053) );
  NAND U37496 ( .A(n37051), .B(n38424), .Z(n37052) );
  AND U37497 ( .A(n37053), .B(n37052), .Z(n37191) );
  XOR U37498 ( .A(n37192), .B(n37191), .Z(n37194) );
  XOR U37499 ( .A(b[25]), .B(n37668), .Z(n37174) );
  NANDN U37500 ( .A(n37174), .B(n38325), .Z(n37056) );
  NAND U37501 ( .A(n38326), .B(n37054), .Z(n37055) );
  NAND U37502 ( .A(n37056), .B(n37055), .Z(n37193) );
  XNOR U37503 ( .A(n37194), .B(n37193), .Z(n37161) );
  NAND U37504 ( .A(n37057), .B(n37762), .Z(n37059) );
  XNOR U37505 ( .A(a[248]), .B(b[17]), .Z(n37209) );
  NANDN U37506 ( .A(n37209), .B(n37764), .Z(n37058) );
  NAND U37507 ( .A(n37059), .B(n37058), .Z(n37158) );
  XOR U37508 ( .A(n38531), .B(b[13]), .Z(n37215) );
  NANDN U37509 ( .A(n37215), .B(n37424), .Z(n37062) );
  NANDN U37510 ( .A(n37060), .B(n37425), .Z(n37061) );
  NAND U37511 ( .A(n37062), .B(n37061), .Z(n37201) );
  XOR U37512 ( .A(a[246]), .B(n1055), .Z(n37180) );
  NANDN U37513 ( .A(n37180), .B(n37934), .Z(n37065) );
  NANDN U37514 ( .A(n37063), .B(n37935), .Z(n37064) );
  AND U37515 ( .A(n37065), .B(n37064), .Z(n37200) );
  XOR U37516 ( .A(n37201), .B(n37200), .Z(n37203) );
  XNOR U37517 ( .A(n38356), .B(b[15]), .Z(n37212) );
  NANDN U37518 ( .A(n37665), .B(n37212), .Z(n37068) );
  NANDN U37519 ( .A(n37066), .B(n37604), .Z(n37067) );
  NAND U37520 ( .A(n37068), .B(n37067), .Z(n37202) );
  XOR U37521 ( .A(n37203), .B(n37202), .Z(n37159) );
  XNOR U37522 ( .A(n37158), .B(n37159), .Z(n37160) );
  XNOR U37523 ( .A(n37161), .B(n37160), .Z(n37149) );
  NANDN U37524 ( .A(n37070), .B(n37069), .Z(n37074) );
  NAND U37525 ( .A(n37072), .B(n37071), .Z(n37073) );
  NAND U37526 ( .A(n37074), .B(n37073), .Z(n37167) );
  XOR U37527 ( .A(n1052), .B(n37183), .Z(n37078) );
  XNOR U37528 ( .A(b[8]), .B(b[7]), .Z(n37075) );
  NANDN U37529 ( .A(n37076), .B(n37075), .Z(n37077) );
  AND U37530 ( .A(n37078), .B(n37077), .Z(n37197) );
  ANDN U37531 ( .B(b[31]), .A(n37079), .Z(n37269) );
  XNOR U37532 ( .A(n37197), .B(n37269), .Z(n37198) );
  XOR U37533 ( .A(n1059), .B(n37080), .Z(n37185) );
  NAND U37534 ( .A(n37185), .B(n38552), .Z(n37083) );
  NANDN U37535 ( .A(n37081), .B(n38553), .Z(n37082) );
  AND U37536 ( .A(n37083), .B(n37082), .Z(n37199) );
  XOR U37537 ( .A(n37198), .B(n37199), .Z(n37165) );
  OR U37538 ( .A(n37085), .B(n37084), .Z(n37089) );
  NAND U37539 ( .A(n37087), .B(n37086), .Z(n37088) );
  NAND U37540 ( .A(n37089), .B(n37088), .Z(n37164) );
  XNOR U37541 ( .A(n37165), .B(n37164), .Z(n37166) );
  XNOR U37542 ( .A(n37167), .B(n37166), .Z(n37146) );
  NANDN U37543 ( .A(n37091), .B(n37090), .Z(n37095) );
  NAND U37544 ( .A(n37093), .B(n37092), .Z(n37094) );
  NAND U37545 ( .A(n37095), .B(n37094), .Z(n37147) );
  XNOR U37546 ( .A(n37146), .B(n37147), .Z(n37148) );
  XOR U37547 ( .A(n37149), .B(n37148), .Z(n37141) );
  NANDN U37548 ( .A(n37097), .B(n37096), .Z(n37101) );
  NAND U37549 ( .A(n37099), .B(n37098), .Z(n37100) );
  NAND U37550 ( .A(n37101), .B(n37100), .Z(n37155) );
  XOR U37551 ( .A(n38532), .B(b[11]), .Z(n37219) );
  OR U37552 ( .A(n37219), .B(n37311), .Z(n37104) );
  NAND U37553 ( .A(n37218), .B(n37102), .Z(n37103) );
  NAND U37554 ( .A(n37104), .B(n37103), .Z(n37170) );
  NANDN U37555 ( .A(n37105), .B(n38490), .Z(n37108) );
  XOR U37556 ( .A(n1058), .B(n37106), .Z(n37206) );
  NANDN U37557 ( .A(n1048), .B(n37206), .Z(n37107) );
  NAND U37558 ( .A(n37108), .B(n37107), .Z(n37168) );
  XOR U37559 ( .A(n1056), .B(a[244]), .Z(n37188) );
  NANDN U37560 ( .A(n37188), .B(n38101), .Z(n37111) );
  NAND U37561 ( .A(n38102), .B(n37109), .Z(n37110) );
  NAND U37562 ( .A(n37111), .B(n37110), .Z(n37169) );
  XOR U37563 ( .A(n37168), .B(n37169), .Z(n37171) );
  XNOR U37564 ( .A(n37170), .B(n37171), .Z(n37152) );
  NANDN U37565 ( .A(n37113), .B(n37112), .Z(n37117) );
  NANDN U37566 ( .A(n37115), .B(n37114), .Z(n37116) );
  NAND U37567 ( .A(n37117), .B(n37116), .Z(n37153) );
  XNOR U37568 ( .A(n37152), .B(n37153), .Z(n37154) );
  XOR U37569 ( .A(n37155), .B(n37154), .Z(n37140) );
  XOR U37570 ( .A(n37141), .B(n37140), .Z(n37142) );
  XOR U37571 ( .A(n37143), .B(n37142), .Z(n37137) );
  XNOR U37572 ( .A(n37136), .B(n37137), .Z(n37231) );
  NAND U37573 ( .A(n37119), .B(n37118), .Z(n37123) );
  NANDN U37574 ( .A(n37121), .B(n37120), .Z(n37122) );
  AND U37575 ( .A(n37123), .B(n37122), .Z(n37232) );
  XNOR U37576 ( .A(n37231), .B(n37232), .Z(n37233) );
  XNOR U37577 ( .A(n37234), .B(n37233), .Z(n37129) );
  XNOR U37578 ( .A(n37128), .B(n37129), .Z(n37130) );
  XNOR U37579 ( .A(n37131), .B(n37130), .Z(n37126) );
  NANDN U37580 ( .A(n37125), .B(n37124), .Z(n37127) );
  XNOR U37581 ( .A(n37126), .B(n37127), .Z(c[488]) );
  NANDN U37582 ( .A(n37127), .B(n37126), .Z(n37340) );
  NANDN U37583 ( .A(n37129), .B(n37128), .Z(n37133) );
  NANDN U37584 ( .A(n37131), .B(n37130), .Z(n37132) );
  NAND U37585 ( .A(n37133), .B(n37132), .Z(n37238) );
  NANDN U37586 ( .A(n37135), .B(n37134), .Z(n37139) );
  NAND U37587 ( .A(n37137), .B(n37136), .Z(n37138) );
  NAND U37588 ( .A(n37139), .B(n37138), .Z(n37242) );
  OR U37589 ( .A(n37141), .B(n37140), .Z(n37145) );
  NAND U37590 ( .A(n37143), .B(n37142), .Z(n37144) );
  NAND U37591 ( .A(n37145), .B(n37144), .Z(n37240) );
  NANDN U37592 ( .A(n37147), .B(n37146), .Z(n37151) );
  NAND U37593 ( .A(n37149), .B(n37148), .Z(n37150) );
  NAND U37594 ( .A(n37151), .B(n37150), .Z(n37254) );
  NANDN U37595 ( .A(n37153), .B(n37152), .Z(n37157) );
  NAND U37596 ( .A(n37155), .B(n37154), .Z(n37156) );
  NAND U37597 ( .A(n37157), .B(n37156), .Z(n37251) );
  NANDN U37598 ( .A(n37159), .B(n37158), .Z(n37163) );
  NAND U37599 ( .A(n37161), .B(n37160), .Z(n37162) );
  NAND U37600 ( .A(n37163), .B(n37162), .Z(n37252) );
  XNOR U37601 ( .A(n37251), .B(n37252), .Z(n37253) );
  XNOR U37602 ( .A(n37254), .B(n37253), .Z(n37248) );
  NAND U37603 ( .A(n37169), .B(n37168), .Z(n37173) );
  NAND U37604 ( .A(n37171), .B(n37170), .Z(n37172) );
  NAND U37605 ( .A(n37173), .B(n37172), .Z(n37292) );
  XNOR U37606 ( .A(b[25]), .B(a[241]), .Z(n37301) );
  NANDN U37607 ( .A(n37301), .B(n38325), .Z(n37176) );
  NANDN U37608 ( .A(n37174), .B(n38326), .Z(n37175) );
  NAND U37609 ( .A(n37176), .B(n37175), .Z(n37338) );
  XNOR U37610 ( .A(b[27]), .B(a[239]), .Z(n37317) );
  NANDN U37611 ( .A(n37317), .B(n38423), .Z(n37179) );
  NAND U37612 ( .A(n38424), .B(n37177), .Z(n37178) );
  NAND U37613 ( .A(n37179), .B(n37178), .Z(n37335) );
  XNOR U37614 ( .A(a[247]), .B(n1055), .Z(n37307) );
  NAND U37615 ( .A(n37307), .B(n37934), .Z(n37182) );
  NANDN U37616 ( .A(n37180), .B(n37935), .Z(n37181) );
  AND U37617 ( .A(n37182), .B(n37181), .Z(n37336) );
  XNOR U37618 ( .A(n37335), .B(n37336), .Z(n37337) );
  XOR U37619 ( .A(n37338), .B(n37337), .Z(n37290) );
  NANDN U37620 ( .A(n1052), .B(n37183), .Z(n37268) );
  ANDN U37621 ( .B(b[31]), .A(n37184), .Z(n37267) );
  XOR U37622 ( .A(n37268), .B(n37267), .Z(n37270) );
  XOR U37623 ( .A(n37269), .B(n37270), .Z(n37295) );
  XOR U37624 ( .A(n1059), .B(a[235]), .Z(n37314) );
  NANDN U37625 ( .A(n37314), .B(n38552), .Z(n37187) );
  NAND U37626 ( .A(n38553), .B(n37185), .Z(n37186) );
  NAND U37627 ( .A(n37187), .B(n37186), .Z(n37296) );
  XOR U37628 ( .A(n37295), .B(n37296), .Z(n37297) );
  XOR U37629 ( .A(n1056), .B(a[245]), .Z(n37304) );
  NANDN U37630 ( .A(n37304), .B(n38101), .Z(n37190) );
  NANDN U37631 ( .A(n37188), .B(n38102), .Z(n37189) );
  NAND U37632 ( .A(n37190), .B(n37189), .Z(n37298) );
  XNOR U37633 ( .A(n37297), .B(n37298), .Z(n37289) );
  XOR U37634 ( .A(n37290), .B(n37289), .Z(n37291) );
  XNOR U37635 ( .A(n37292), .B(n37291), .Z(n37265) );
  NANDN U37636 ( .A(n37192), .B(n37191), .Z(n37196) );
  OR U37637 ( .A(n37194), .B(n37193), .Z(n37195) );
  NAND U37638 ( .A(n37196), .B(n37195), .Z(n37264) );
  XOR U37639 ( .A(n37264), .B(n37263), .Z(n37266) );
  XNOR U37640 ( .A(n37265), .B(n37266), .Z(n37258) );
  NANDN U37641 ( .A(n37201), .B(n37200), .Z(n37205) );
  OR U37642 ( .A(n37203), .B(n37202), .Z(n37204) );
  NAND U37643 ( .A(n37205), .B(n37204), .Z(n37286) );
  NAND U37644 ( .A(n37206), .B(n38490), .Z(n37208) );
  XNOR U37645 ( .A(b[29]), .B(a[237]), .Z(n37320) );
  OR U37646 ( .A(n37320), .B(n1048), .Z(n37207) );
  NAND U37647 ( .A(n37208), .B(n37207), .Z(n37282) );
  XNOR U37648 ( .A(a[249]), .B(b[17]), .Z(n37323) );
  NANDN U37649 ( .A(n37323), .B(n37764), .Z(n37211) );
  NANDN U37650 ( .A(n37209), .B(n37762), .Z(n37210) );
  NAND U37651 ( .A(n37211), .B(n37210), .Z(n37279) );
  XNOR U37652 ( .A(a[251]), .B(b[15]), .Z(n37329) );
  OR U37653 ( .A(n37329), .B(n37665), .Z(n37214) );
  NAND U37654 ( .A(n37212), .B(n37604), .Z(n37213) );
  AND U37655 ( .A(n37214), .B(n37213), .Z(n37280) );
  XNOR U37656 ( .A(n37279), .B(n37280), .Z(n37281) );
  XOR U37657 ( .A(n37282), .B(n37281), .Z(n37283) );
  XOR U37658 ( .A(a[253]), .B(n1053), .Z(n37332) );
  NANDN U37659 ( .A(n37332), .B(n37424), .Z(n37217) );
  NANDN U37660 ( .A(n37215), .B(n37425), .Z(n37216) );
  NAND U37661 ( .A(n37217), .B(n37216), .Z(n37275) );
  XNOR U37662 ( .A(a[255]), .B(b[11]), .Z(n37310) );
  OR U37663 ( .A(n37310), .B(n37311), .Z(n37221) );
  NANDN U37664 ( .A(n37219), .B(n37218), .Z(n37220) );
  NAND U37665 ( .A(n37221), .B(n37220), .Z(n37273) );
  XOR U37666 ( .A(n1057), .B(a[243]), .Z(n37326) );
  OR U37667 ( .A(n37326), .B(n38268), .Z(n37224) );
  NANDN U37668 ( .A(n37222), .B(n38205), .Z(n37223) );
  NAND U37669 ( .A(n37224), .B(n37223), .Z(n37274) );
  XOR U37670 ( .A(n37273), .B(n37274), .Z(n37276) );
  XOR U37671 ( .A(n37275), .B(n37276), .Z(n37284) );
  XOR U37672 ( .A(n37283), .B(n37284), .Z(n37285) );
  XOR U37673 ( .A(n37286), .B(n37285), .Z(n37257) );
  XOR U37674 ( .A(n37258), .B(n37257), .Z(n37259) );
  XOR U37675 ( .A(n37260), .B(n37259), .Z(n37245) );
  NANDN U37676 ( .A(n37226), .B(n37225), .Z(n37230) );
  NAND U37677 ( .A(n37228), .B(n37227), .Z(n37229) );
  AND U37678 ( .A(n37230), .B(n37229), .Z(n37246) );
  XNOR U37679 ( .A(n37245), .B(n37246), .Z(n37247) );
  XOR U37680 ( .A(n37248), .B(n37247), .Z(n37239) );
  XOR U37681 ( .A(n37240), .B(n37239), .Z(n37241) );
  XOR U37682 ( .A(n37242), .B(n37241), .Z(n37236) );
  XNOR U37683 ( .A(n37236), .B(n37237), .Z(n37235) );
  XOR U37684 ( .A(n37238), .B(n37235), .Z(n37339) );
  XNOR U37685 ( .A(n37340), .B(n37339), .Z(c[489]) );
  NAND U37686 ( .A(n37240), .B(n37239), .Z(n37244) );
  NAND U37687 ( .A(n37242), .B(n37241), .Z(n37243) );
  NAND U37688 ( .A(n37244), .B(n37243), .Z(n37343) );
  NANDN U37689 ( .A(n37246), .B(n37245), .Z(n37250) );
  NAND U37690 ( .A(n37248), .B(n37247), .Z(n37249) );
  NAND U37691 ( .A(n37250), .B(n37249), .Z(n37352) );
  NANDN U37692 ( .A(n37252), .B(n37251), .Z(n37256) );
  NAND U37693 ( .A(n37254), .B(n37253), .Z(n37255) );
  NAND U37694 ( .A(n37256), .B(n37255), .Z(n37350) );
  NAND U37695 ( .A(n37258), .B(n37257), .Z(n37262) );
  NANDN U37696 ( .A(n37260), .B(n37259), .Z(n37261) );
  NAND U37697 ( .A(n37262), .B(n37261), .Z(n37441) );
  NAND U37698 ( .A(n37268), .B(n37267), .Z(n37272) );
  NAND U37699 ( .A(n37270), .B(n37269), .Z(n37271) );
  NAND U37700 ( .A(n37272), .B(n37271), .Z(n37364) );
  NAND U37701 ( .A(n37274), .B(n37273), .Z(n37278) );
  NAND U37702 ( .A(n37276), .B(n37275), .Z(n37277) );
  NAND U37703 ( .A(n37278), .B(n37277), .Z(n37362) );
  XOR U37704 ( .A(n37362), .B(n37361), .Z(n37363) );
  XOR U37705 ( .A(n37364), .B(n37363), .Z(n37432) );
  OR U37706 ( .A(n37284), .B(n37283), .Z(n37288) );
  NAND U37707 ( .A(n37286), .B(n37285), .Z(n37287) );
  NAND U37708 ( .A(n37288), .B(n37287), .Z(n37433) );
  XNOR U37709 ( .A(n37432), .B(n37433), .Z(n37434) );
  NANDN U37710 ( .A(n37290), .B(n37289), .Z(n37294) );
  OR U37711 ( .A(n37292), .B(n37291), .Z(n37293) );
  NAND U37712 ( .A(n37294), .B(n37293), .Z(n37358) );
  OR U37713 ( .A(n37296), .B(n37295), .Z(n37300) );
  NANDN U37714 ( .A(n37298), .B(n37297), .Z(n37299) );
  NAND U37715 ( .A(n37300), .B(n37299), .Z(n37373) );
  XOR U37716 ( .A(b[25]), .B(n37676), .Z(n37399) );
  NANDN U37717 ( .A(n37399), .B(n38325), .Z(n37303) );
  NANDN U37718 ( .A(n37301), .B(n38326), .Z(n37302) );
  NAND U37719 ( .A(n37303), .B(n37302), .Z(n37383) );
  XOR U37720 ( .A(n1056), .B(a[246]), .Z(n37429) );
  NANDN U37721 ( .A(n37429), .B(n38101), .Z(n37306) );
  NANDN U37722 ( .A(n37304), .B(n38102), .Z(n37305) );
  NAND U37723 ( .A(n37306), .B(n37305), .Z(n37381) );
  XOR U37724 ( .A(a[248]), .B(n1055), .Z(n37405) );
  NANDN U37725 ( .A(n37405), .B(n37934), .Z(n37309) );
  NAND U37726 ( .A(n37935), .B(n37307), .Z(n37308) );
  NAND U37727 ( .A(n37309), .B(n37308), .Z(n37382) );
  XOR U37728 ( .A(n37381), .B(n37382), .Z(n37384) );
  XOR U37729 ( .A(n37383), .B(n37384), .Z(n37374) );
  XNOR U37730 ( .A(n37373), .B(n37374), .Z(n37375) );
  NANDN U37731 ( .A(n1052), .B(b[10]), .Z(n37419) );
  XNOR U37732 ( .A(b[11]), .B(n37419), .Z(n37313) );
  NAND U37733 ( .A(n37311), .B(n37310), .Z(n37312) );
  AND U37734 ( .A(n37313), .B(n37312), .Z(n37408) );
  AND U37735 ( .A(a[234]), .B(b[31]), .Z(n37513) );
  XOR U37736 ( .A(n37408), .B(n37513), .Z(n37410) );
  XOR U37737 ( .A(n1059), .B(a[236]), .Z(n37416) );
  NANDN U37738 ( .A(n37416), .B(n38552), .Z(n37316) );
  NANDN U37739 ( .A(n37314), .B(n38553), .Z(n37315) );
  NAND U37740 ( .A(n37316), .B(n37315), .Z(n37409) );
  XOR U37741 ( .A(n37410), .B(n37409), .Z(n37376) );
  XOR U37742 ( .A(n37375), .B(n37376), .Z(n37356) );
  XOR U37743 ( .A(b[27]), .B(n37668), .Z(n37402) );
  NANDN U37744 ( .A(n37402), .B(n38423), .Z(n37319) );
  NANDN U37745 ( .A(n37317), .B(n38424), .Z(n37318) );
  NAND U37746 ( .A(n37319), .B(n37318), .Z(n37380) );
  NANDN U37747 ( .A(n37320), .B(n38490), .Z(n37322) );
  XOR U37748 ( .A(b[29]), .B(n37467), .Z(n37421) );
  OR U37749 ( .A(n37421), .B(n1048), .Z(n37321) );
  NAND U37750 ( .A(n37322), .B(n37321), .Z(n37377) );
  NANDN U37751 ( .A(n37323), .B(n37762), .Z(n37325) );
  XNOR U37752 ( .A(a[250]), .B(b[17]), .Z(n37393) );
  NANDN U37753 ( .A(n37393), .B(n37764), .Z(n37324) );
  AND U37754 ( .A(n37325), .B(n37324), .Z(n37378) );
  XNOR U37755 ( .A(n37377), .B(n37378), .Z(n37379) );
  XOR U37756 ( .A(n37380), .B(n37379), .Z(n37367) );
  XOR U37757 ( .A(n1057), .B(a[244]), .Z(n37413) );
  OR U37758 ( .A(n37413), .B(n38268), .Z(n37328) );
  NANDN U37759 ( .A(n37326), .B(n38205), .Z(n37327) );
  NAND U37760 ( .A(n37328), .B(n37327), .Z(n37389) );
  XOR U37761 ( .A(a[252]), .B(n1054), .Z(n37396) );
  OR U37762 ( .A(n37396), .B(n37665), .Z(n37331) );
  NANDN U37763 ( .A(n37329), .B(n37604), .Z(n37330) );
  NAND U37764 ( .A(n37331), .B(n37330), .Z(n37387) );
  XOR U37765 ( .A(n38532), .B(b[13]), .Z(n37426) );
  NANDN U37766 ( .A(n37426), .B(n37424), .Z(n37334) );
  NANDN U37767 ( .A(n37332), .B(n37425), .Z(n37333) );
  NAND U37768 ( .A(n37334), .B(n37333), .Z(n37388) );
  XOR U37769 ( .A(n37387), .B(n37388), .Z(n37390) );
  XOR U37770 ( .A(n37389), .B(n37390), .Z(n37368) );
  XOR U37771 ( .A(n37367), .B(n37368), .Z(n37369) );
  XNOR U37772 ( .A(n37369), .B(n37370), .Z(n37355) );
  XOR U37773 ( .A(n37356), .B(n37355), .Z(n37357) );
  XOR U37774 ( .A(n37358), .B(n37357), .Z(n37435) );
  XOR U37775 ( .A(n37434), .B(n37435), .Z(n37438) );
  XOR U37776 ( .A(n37439), .B(n37438), .Z(n37440) );
  XNOR U37777 ( .A(n37441), .B(n37440), .Z(n37349) );
  XNOR U37778 ( .A(n37350), .B(n37349), .Z(n37351) );
  XNOR U37779 ( .A(n37352), .B(n37351), .Z(n37344) );
  XNOR U37780 ( .A(n37343), .B(n37344), .Z(n37346) );
  XOR U37781 ( .A(n37345), .B(n37346), .Z(n37341) );
  NANDN U37782 ( .A(n37340), .B(n37339), .Z(n37342) );
  XNOR U37783 ( .A(n37341), .B(n37342), .Z(c[490]) );
  NANDN U37784 ( .A(n37342), .B(n37341), .Z(n37542) );
  NANDN U37785 ( .A(n37344), .B(n37343), .Z(n37348) );
  NAND U37786 ( .A(n37346), .B(n37345), .Z(n37347) );
  AND U37787 ( .A(n37348), .B(n37347), .Z(n37536) );
  NANDN U37788 ( .A(n37350), .B(n37349), .Z(n37354) );
  NAND U37789 ( .A(n37352), .B(n37351), .Z(n37353) );
  AND U37790 ( .A(n37354), .B(n37353), .Z(n37534) );
  NANDN U37791 ( .A(n37356), .B(n37355), .Z(n37360) );
  OR U37792 ( .A(n37358), .B(n37357), .Z(n37359) );
  NAND U37793 ( .A(n37360), .B(n37359), .Z(n37451) );
  OR U37794 ( .A(n37362), .B(n37361), .Z(n37366) );
  NANDN U37795 ( .A(n37364), .B(n37363), .Z(n37365) );
  NAND U37796 ( .A(n37366), .B(n37365), .Z(n37452) );
  XNOR U37797 ( .A(n37451), .B(n37452), .Z(n37453) );
  OR U37798 ( .A(n37368), .B(n37367), .Z(n37372) );
  NAND U37799 ( .A(n37370), .B(n37369), .Z(n37371) );
  NAND U37800 ( .A(n37372), .B(n37371), .Z(n37530) );
  XNOR U37801 ( .A(n37530), .B(n37529), .Z(n37531) );
  NAND U37802 ( .A(n37382), .B(n37381), .Z(n37386) );
  NAND U37803 ( .A(n37384), .B(n37383), .Z(n37385) );
  NAND U37804 ( .A(n37386), .B(n37385), .Z(n37524) );
  NAND U37805 ( .A(n37388), .B(n37387), .Z(n37392) );
  NAND U37806 ( .A(n37390), .B(n37389), .Z(n37391) );
  NAND U37807 ( .A(n37392), .B(n37391), .Z(n37518) );
  XNOR U37808 ( .A(a[251]), .B(b[17]), .Z(n37502) );
  NANDN U37809 ( .A(n37502), .B(n37764), .Z(n37395) );
  NANDN U37810 ( .A(n37393), .B(n37762), .Z(n37394) );
  NAND U37811 ( .A(n37395), .B(n37394), .Z(n37480) );
  XNOR U37812 ( .A(a[253]), .B(n1054), .Z(n37505) );
  NANDN U37813 ( .A(n37665), .B(n37505), .Z(n37398) );
  NANDN U37814 ( .A(n37396), .B(n37604), .Z(n37397) );
  NAND U37815 ( .A(n37398), .B(n37397), .Z(n37478) );
  XNOR U37816 ( .A(b[25]), .B(a[243]), .Z(n37508) );
  NANDN U37817 ( .A(n37508), .B(n38325), .Z(n37401) );
  NANDN U37818 ( .A(n37399), .B(n38326), .Z(n37400) );
  NAND U37819 ( .A(n37401), .B(n37400), .Z(n37457) );
  XOR U37820 ( .A(b[27]), .B(a[241]), .Z(n37493) );
  NAND U37821 ( .A(n38423), .B(n37493), .Z(n37404) );
  NANDN U37822 ( .A(n37402), .B(n38424), .Z(n37403) );
  NAND U37823 ( .A(n37404), .B(n37403), .Z(n37455) );
  XNOR U37824 ( .A(a[249]), .B(b[19]), .Z(n37487) );
  NANDN U37825 ( .A(n37487), .B(n37934), .Z(n37407) );
  NANDN U37826 ( .A(n37405), .B(n37935), .Z(n37406) );
  AND U37827 ( .A(n37407), .B(n37406), .Z(n37456) );
  XNOR U37828 ( .A(n37455), .B(n37456), .Z(n37458) );
  XOR U37829 ( .A(n37457), .B(n37458), .Z(n37477) );
  XOR U37830 ( .A(n37478), .B(n37477), .Z(n37479) );
  XOR U37831 ( .A(n37480), .B(n37479), .Z(n37517) );
  XOR U37832 ( .A(n37518), .B(n37517), .Z(n37519) );
  NANDN U37833 ( .A(n37408), .B(n37513), .Z(n37412) );
  OR U37834 ( .A(n37410), .B(n37409), .Z(n37411) );
  NAND U37835 ( .A(n37412), .B(n37411), .Z(n37474) );
  XOR U37836 ( .A(b[23]), .B(n38213), .Z(n37499) );
  OR U37837 ( .A(n37499), .B(n38268), .Z(n37415) );
  NANDN U37838 ( .A(n37413), .B(n38205), .Z(n37414) );
  NAND U37839 ( .A(n37415), .B(n37414), .Z(n37462) );
  XNOR U37840 ( .A(b[31]), .B(a[237]), .Z(n37468) );
  NANDN U37841 ( .A(n37468), .B(n38552), .Z(n37418) );
  NANDN U37842 ( .A(n37416), .B(n38553), .Z(n37417) );
  NAND U37843 ( .A(n37418), .B(n37417), .Z(n37459) );
  AND U37844 ( .A(n37419), .B(b[11]), .Z(n37512) );
  NANDN U37845 ( .A(n37420), .B(b[31]), .Z(n37511) );
  XOR U37846 ( .A(n37512), .B(n37511), .Z(n37514) );
  XNOR U37847 ( .A(n37513), .B(n37514), .Z(n37460) );
  XNOR U37848 ( .A(n37459), .B(n37460), .Z(n37461) );
  XOR U37849 ( .A(n37462), .B(n37461), .Z(n37471) );
  NANDN U37850 ( .A(n37421), .B(n38490), .Z(n37423) );
  XNOR U37851 ( .A(n1058), .B(a[239]), .Z(n37496) );
  NANDN U37852 ( .A(n1048), .B(n37496), .Z(n37422) );
  NAND U37853 ( .A(n37423), .B(n37422), .Z(n37483) );
  XOR U37854 ( .A(a[255]), .B(n1053), .Z(n37463) );
  NANDN U37855 ( .A(n37463), .B(n37424), .Z(n37428) );
  NANDN U37856 ( .A(n37426), .B(n37425), .Z(n37427) );
  NAND U37857 ( .A(n37428), .B(n37427), .Z(n37481) );
  XNOR U37858 ( .A(b[21]), .B(a[247]), .Z(n37490) );
  NANDN U37859 ( .A(n37490), .B(n38101), .Z(n37431) );
  NANDN U37860 ( .A(n37429), .B(n38102), .Z(n37430) );
  NAND U37861 ( .A(n37431), .B(n37430), .Z(n37482) );
  XOR U37862 ( .A(n37481), .B(n37482), .Z(n37484) );
  XOR U37863 ( .A(n37483), .B(n37484), .Z(n37472) );
  XNOR U37864 ( .A(n37471), .B(n37472), .Z(n37473) );
  XOR U37865 ( .A(n37474), .B(n37473), .Z(n37520) );
  XOR U37866 ( .A(n37519), .B(n37520), .Z(n37523) );
  XOR U37867 ( .A(n37524), .B(n37523), .Z(n37525) );
  XOR U37868 ( .A(n37526), .B(n37525), .Z(n37532) );
  XOR U37869 ( .A(n37531), .B(n37532), .Z(n37454) );
  XOR U37870 ( .A(n37453), .B(n37454), .Z(n37445) );
  NANDN U37871 ( .A(n37433), .B(n37432), .Z(n37437) );
  NAND U37872 ( .A(n37435), .B(n37434), .Z(n37436) );
  NAND U37873 ( .A(n37437), .B(n37436), .Z(n37446) );
  XOR U37874 ( .A(n37445), .B(n37446), .Z(n37447) );
  NAND U37875 ( .A(n37439), .B(n37438), .Z(n37443) );
  NANDN U37876 ( .A(n37441), .B(n37440), .Z(n37442) );
  NAND U37877 ( .A(n37443), .B(n37442), .Z(n37448) );
  XNOR U37878 ( .A(n37447), .B(n37448), .Z(n37535) );
  IV U37879 ( .A(n37535), .Z(n37533) );
  XOR U37880 ( .A(n37534), .B(n37533), .Z(n37444) );
  XOR U37881 ( .A(n37536), .B(n37444), .Z(n37541) );
  XNOR U37882 ( .A(n37542), .B(n37541), .Z(c[491]) );
  OR U37883 ( .A(n37446), .B(n37445), .Z(n37450) );
  NANDN U37884 ( .A(n37448), .B(n37447), .Z(n37449) );
  NAND U37885 ( .A(n37450), .B(n37449), .Z(n37545) );
  XNOR U37886 ( .A(n37554), .B(n37555), .Z(n37556) );
  NAND U37887 ( .A(b[11]), .B(b[12]), .Z(n37603) );
  XOR U37888 ( .A(n1053), .B(n37603), .Z(n37466) );
  XNOR U37889 ( .A(b[12]), .B(b[11]), .Z(n37464) );
  NAND U37890 ( .A(n37464), .B(n37463), .Z(n37465) );
  AND U37891 ( .A(n37466), .B(n37465), .Z(n37612) );
  AND U37892 ( .A(a[236]), .B(b[31]), .Z(n37653) );
  XOR U37893 ( .A(b[31]), .B(n37467), .Z(n37576) );
  NANDN U37894 ( .A(n37576), .B(n38552), .Z(n37470) );
  NANDN U37895 ( .A(n37468), .B(n38553), .Z(n37469) );
  AND U37896 ( .A(n37470), .B(n37469), .Z(n37611) );
  XOR U37897 ( .A(n37653), .B(n37611), .Z(n37613) );
  XOR U37898 ( .A(n37612), .B(n37613), .Z(n37557) );
  XNOR U37899 ( .A(n37556), .B(n37557), .Z(n37622) );
  NAND U37900 ( .A(n37472), .B(n37471), .Z(n37476) );
  OR U37901 ( .A(n37474), .B(n37473), .Z(n37475) );
  NAND U37902 ( .A(n37476), .B(n37475), .Z(n37623) );
  XNOR U37903 ( .A(n37622), .B(n37623), .Z(n37624) );
  NAND U37904 ( .A(n37482), .B(n37481), .Z(n37486) );
  NAND U37905 ( .A(n37484), .B(n37483), .Z(n37485) );
  NAND U37906 ( .A(n37486), .B(n37485), .Z(n37559) );
  XOR U37907 ( .A(a[250]), .B(n1055), .Z(n37585) );
  NANDN U37908 ( .A(n37585), .B(n37934), .Z(n37489) );
  NANDN U37909 ( .A(n37487), .B(n37935), .Z(n37488) );
  NAND U37910 ( .A(n37489), .B(n37488), .Z(n37594) );
  XOR U37911 ( .A(n38272), .B(n1056), .Z(n37588) );
  NAND U37912 ( .A(n37588), .B(n38101), .Z(n37492) );
  NANDN U37913 ( .A(n37490), .B(n38102), .Z(n37491) );
  NAND U37914 ( .A(n37492), .B(n37491), .Z(n37591) );
  XNOR U37915 ( .A(b[27]), .B(a[242]), .Z(n37579) );
  NANDN U37916 ( .A(n37579), .B(n38423), .Z(n37495) );
  NAND U37917 ( .A(n37493), .B(n38424), .Z(n37494) );
  NAND U37918 ( .A(n37495), .B(n37494), .Z(n37600) );
  NAND U37919 ( .A(n37496), .B(n38490), .Z(n37498) );
  XOR U37920 ( .A(n1058), .B(n37668), .Z(n37582) );
  NANDN U37921 ( .A(n1048), .B(n37582), .Z(n37497) );
  AND U37922 ( .A(n37498), .B(n37497), .Z(n37597) );
  NANDN U37923 ( .A(n37499), .B(n38205), .Z(n37501) );
  XOR U37924 ( .A(b[23]), .B(n38146), .Z(n37570) );
  OR U37925 ( .A(n37570), .B(n38268), .Z(n37500) );
  AND U37926 ( .A(n37501), .B(n37500), .Z(n37598) );
  XNOR U37927 ( .A(n37600), .B(n37599), .Z(n37592) );
  XNOR U37928 ( .A(n37591), .B(n37592), .Z(n37593) );
  XNOR U37929 ( .A(n37594), .B(n37593), .Z(n37618) );
  NANDN U37930 ( .A(n37502), .B(n37762), .Z(n37504) );
  XNOR U37931 ( .A(a[252]), .B(b[17]), .Z(n37573) );
  NANDN U37932 ( .A(n37573), .B(n37764), .Z(n37503) );
  NAND U37933 ( .A(n37504), .B(n37503), .Z(n37567) );
  XOR U37934 ( .A(a[254]), .B(n1054), .Z(n37605) );
  OR U37935 ( .A(n37605), .B(n37665), .Z(n37507) );
  NAND U37936 ( .A(n37505), .B(n37604), .Z(n37506) );
  NAND U37937 ( .A(n37507), .B(n37506), .Z(n37564) );
  XNOR U37938 ( .A(b[25]), .B(n38034), .Z(n37608) );
  NAND U37939 ( .A(n37608), .B(n38325), .Z(n37510) );
  NANDN U37940 ( .A(n37508), .B(n38326), .Z(n37509) );
  AND U37941 ( .A(n37510), .B(n37509), .Z(n37565) );
  XNOR U37942 ( .A(n37564), .B(n37565), .Z(n37566) );
  XNOR U37943 ( .A(n37567), .B(n37566), .Z(n37617) );
  OR U37944 ( .A(n37512), .B(n37511), .Z(n37516) );
  NAND U37945 ( .A(n37514), .B(n37513), .Z(n37515) );
  AND U37946 ( .A(n37516), .B(n37515), .Z(n37616) );
  XOR U37947 ( .A(n37617), .B(n37616), .Z(n37619) );
  XOR U37948 ( .A(n37618), .B(n37619), .Z(n37558) );
  XNOR U37949 ( .A(n37559), .B(n37558), .Z(n37560) );
  XOR U37950 ( .A(n37561), .B(n37560), .Z(n37625) );
  XOR U37951 ( .A(n37624), .B(n37625), .Z(n37631) );
  NAND U37952 ( .A(n37518), .B(n37517), .Z(n37522) );
  NAND U37953 ( .A(n37520), .B(n37519), .Z(n37521) );
  NAND U37954 ( .A(n37522), .B(n37521), .Z(n37628) );
  NAND U37955 ( .A(n37524), .B(n37523), .Z(n37528) );
  NAND U37956 ( .A(n37526), .B(n37525), .Z(n37527) );
  AND U37957 ( .A(n37528), .B(n37527), .Z(n37629) );
  XNOR U37958 ( .A(n37628), .B(n37629), .Z(n37630) );
  XNOR U37959 ( .A(n37631), .B(n37630), .Z(n37549) );
  XOR U37960 ( .A(n37549), .B(n37548), .Z(n37550) );
  XOR U37961 ( .A(n37551), .B(n37550), .Z(n37546) );
  NANDN U37962 ( .A(n37533), .B(n37534), .Z(n37539) );
  NOR U37963 ( .A(n37535), .B(n37534), .Z(n37537) );
  NANDN U37964 ( .A(n37537), .B(n37536), .Z(n37538) );
  NAND U37965 ( .A(n37539), .B(n37538), .Z(n37547) );
  XNOR U37966 ( .A(n37546), .B(n37547), .Z(n37540) );
  XNOR U37967 ( .A(n37545), .B(n37540), .Z(n37543) );
  NANDN U37968 ( .A(n37542), .B(n37541), .Z(n37544) );
  XNOR U37969 ( .A(n37543), .B(n37544), .Z(c[492]) );
  NANDN U37970 ( .A(n37544), .B(n37543), .Z(n37721) );
  NAND U37971 ( .A(n37549), .B(n37548), .Z(n37553) );
  NANDN U37972 ( .A(n37551), .B(n37550), .Z(n37552) );
  AND U37973 ( .A(n37553), .B(n37552), .Z(n37717) );
  NANDN U37974 ( .A(n37559), .B(n37558), .Z(n37563) );
  NANDN U37975 ( .A(n37561), .B(n37560), .Z(n37562) );
  NAND U37976 ( .A(n37563), .B(n37562), .Z(n37713) );
  XNOR U37977 ( .A(n37712), .B(n37713), .Z(n37714) );
  NANDN U37978 ( .A(n37565), .B(n37564), .Z(n37569) );
  NAND U37979 ( .A(n37567), .B(n37566), .Z(n37568) );
  NAND U37980 ( .A(n37569), .B(n37568), .Z(n37644) );
  NANDN U37981 ( .A(n37570), .B(n38205), .Z(n37572) );
  XNOR U37982 ( .A(b[23]), .B(a[247]), .Z(n37685) );
  OR U37983 ( .A(n37685), .B(n38268), .Z(n37571) );
  NAND U37984 ( .A(n37572), .B(n37571), .Z(n37697) );
  NANDN U37985 ( .A(n37573), .B(n37762), .Z(n37575) );
  XOR U37986 ( .A(a[253]), .B(b[17]), .Z(n37688) );
  NAND U37987 ( .A(n37688), .B(n37764), .Z(n37574) );
  NAND U37988 ( .A(n37575), .B(n37574), .Z(n37694) );
  XNOR U37989 ( .A(b[31]), .B(a[239]), .Z(n37669) );
  NANDN U37990 ( .A(n37669), .B(n38552), .Z(n37578) );
  NANDN U37991 ( .A(n37576), .B(n38553), .Z(n37577) );
  AND U37992 ( .A(n37578), .B(n37577), .Z(n37695) );
  XNOR U37993 ( .A(n37694), .B(n37695), .Z(n37696) );
  XNOR U37994 ( .A(n37697), .B(n37696), .Z(n37650) );
  XNOR U37995 ( .A(b[27]), .B(a[243]), .Z(n37672) );
  NANDN U37996 ( .A(n37672), .B(n38423), .Z(n37581) );
  NANDN U37997 ( .A(n37579), .B(n38424), .Z(n37580) );
  NAND U37998 ( .A(n37581), .B(n37580), .Z(n37703) );
  NAND U37999 ( .A(n38490), .B(n37582), .Z(n37584) );
  XNOR U38000 ( .A(n1058), .B(a[241]), .Z(n37675) );
  NANDN U38001 ( .A(n1048), .B(n37675), .Z(n37583) );
  NAND U38002 ( .A(n37584), .B(n37583), .Z(n37700) );
  XNOR U38003 ( .A(a[251]), .B(n1055), .Z(n37691) );
  NAND U38004 ( .A(n37691), .B(n37934), .Z(n37587) );
  NANDN U38005 ( .A(n37585), .B(n37935), .Z(n37586) );
  AND U38006 ( .A(n37587), .B(n37586), .Z(n37701) );
  XNOR U38007 ( .A(n37700), .B(n37701), .Z(n37702) );
  XNOR U38008 ( .A(n37703), .B(n37702), .Z(n37647) );
  XNOR U38009 ( .A(a[249]), .B(b[21]), .Z(n37682) );
  NANDN U38010 ( .A(n37682), .B(n38101), .Z(n37590) );
  NAND U38011 ( .A(n38102), .B(n37588), .Z(n37589) );
  NAND U38012 ( .A(n37590), .B(n37589), .Z(n37648) );
  XNOR U38013 ( .A(n37647), .B(n37648), .Z(n37649) );
  XOR U38014 ( .A(n37650), .B(n37649), .Z(n37643) );
  XNOR U38015 ( .A(n37644), .B(n37643), .Z(n37645) );
  NANDN U38016 ( .A(n37592), .B(n37591), .Z(n37596) );
  NAND U38017 ( .A(n37594), .B(n37593), .Z(n37595) );
  AND U38018 ( .A(n37596), .B(n37595), .Z(n37646) );
  XNOR U38019 ( .A(n37645), .B(n37646), .Z(n37708) );
  OR U38020 ( .A(n37598), .B(n37597), .Z(n37602) );
  NAND U38021 ( .A(n37600), .B(n37599), .Z(n37601) );
  NAND U38022 ( .A(n37602), .B(n37601), .Z(n37640) );
  NAND U38023 ( .A(b[13]), .B(n37603), .Z(n37651) );
  NANDN U38024 ( .A(n1059), .B(a[237]), .Z(n37652) );
  XOR U38025 ( .A(n37651), .B(n37652), .Z(n37654) );
  XNOR U38026 ( .A(n37653), .B(n37654), .Z(n37657) );
  NANDN U38027 ( .A(n37605), .B(n37604), .Z(n37607) );
  XOR U38028 ( .A(a[255]), .B(n1054), .Z(n37664) );
  OR U38029 ( .A(n37664), .B(n37665), .Z(n37606) );
  NAND U38030 ( .A(n37607), .B(n37606), .Z(n37658) );
  XOR U38031 ( .A(n37657), .B(n37658), .Z(n37659) );
  XNOR U38032 ( .A(b[25]), .B(a[245]), .Z(n37679) );
  NANDN U38033 ( .A(n37679), .B(n38325), .Z(n37610) );
  NAND U38034 ( .A(n38326), .B(n37608), .Z(n37609) );
  AND U38035 ( .A(n37610), .B(n37609), .Z(n37660) );
  XOR U38036 ( .A(n37659), .B(n37660), .Z(n37639) );
  XNOR U38037 ( .A(n37640), .B(n37639), .Z(n37641) );
  OR U38038 ( .A(n37653), .B(n37611), .Z(n37615) );
  NAND U38039 ( .A(n37613), .B(n37612), .Z(n37614) );
  AND U38040 ( .A(n37615), .B(n37614), .Z(n37642) );
  XNOR U38041 ( .A(n37641), .B(n37642), .Z(n37707) );
  NAND U38042 ( .A(n37617), .B(n37616), .Z(n37621) );
  NAND U38043 ( .A(n37619), .B(n37618), .Z(n37620) );
  AND U38044 ( .A(n37621), .B(n37620), .Z(n37706) );
  XOR U38045 ( .A(n37707), .B(n37706), .Z(n37709) );
  XOR U38046 ( .A(n37708), .B(n37709), .Z(n37715) );
  XNOR U38047 ( .A(n37714), .B(n37715), .Z(n37633) );
  NANDN U38048 ( .A(n37623), .B(n37622), .Z(n37627) );
  NANDN U38049 ( .A(n37625), .B(n37624), .Z(n37626) );
  AND U38050 ( .A(n37627), .B(n37626), .Z(n37634) );
  XNOR U38051 ( .A(n37633), .B(n37634), .Z(n37635) );
  XNOR U38052 ( .A(n37635), .B(n37636), .Z(n37716) );
  XNOR U38053 ( .A(n37717), .B(n37716), .Z(n37632) );
  XNOR U38054 ( .A(n37718), .B(n37632), .Z(n37720) );
  XOR U38055 ( .A(n37721), .B(n37720), .Z(c[493]) );
  NANDN U38056 ( .A(n37634), .B(n37633), .Z(n37638) );
  NANDN U38057 ( .A(n37636), .B(n37635), .Z(n37637) );
  NAND U38058 ( .A(n37638), .B(n37637), .Z(n37801) );
  XNOR U38059 ( .A(n37729), .B(n37728), .Z(n37730) );
  NANDN U38060 ( .A(n37652), .B(n37651), .Z(n37656) );
  NANDN U38061 ( .A(n37654), .B(n37653), .Z(n37655) );
  NAND U38062 ( .A(n37656), .B(n37655), .Z(n37738) );
  OR U38063 ( .A(n37658), .B(n37657), .Z(n37662) );
  NAND U38064 ( .A(n37660), .B(n37659), .Z(n37661) );
  NAND U38065 ( .A(n37662), .B(n37661), .Z(n37739) );
  XNOR U38066 ( .A(n37738), .B(n37739), .Z(n37740) );
  XOR U38067 ( .A(n1054), .B(n37663), .Z(n37667) );
  NAND U38068 ( .A(n37665), .B(n37664), .Z(n37666) );
  AND U38069 ( .A(n37667), .B(n37666), .Z(n37789) );
  AND U38070 ( .A(a[238]), .B(b[31]), .Z(n37853) );
  XOR U38071 ( .A(b[31]), .B(n37668), .Z(n37773) );
  NANDN U38072 ( .A(n37773), .B(n38552), .Z(n37671) );
  NANDN U38073 ( .A(n37669), .B(n38553), .Z(n37670) );
  AND U38074 ( .A(n37671), .B(n37670), .Z(n37788) );
  XOR U38075 ( .A(n37853), .B(n37788), .Z(n37790) );
  XOR U38076 ( .A(n37789), .B(n37790), .Z(n37741) );
  XOR U38077 ( .A(n37740), .B(n37741), .Z(n37734) );
  XNOR U38078 ( .A(n37735), .B(n37734), .Z(n37736) );
  XNOR U38079 ( .A(b[27]), .B(a[244]), .Z(n37779) );
  NANDN U38080 ( .A(n37779), .B(n38423), .Z(n37674) );
  NANDN U38081 ( .A(n37672), .B(n38424), .Z(n37673) );
  NAND U38082 ( .A(n37674), .B(n37673), .Z(n37770) );
  NAND U38083 ( .A(n38490), .B(n37675), .Z(n37678) );
  XOR U38084 ( .A(n1058), .B(n37676), .Z(n37782) );
  NANDN U38085 ( .A(n1048), .B(n37782), .Z(n37677) );
  NAND U38086 ( .A(n37678), .B(n37677), .Z(n37767) );
  XNOR U38087 ( .A(b[25]), .B(a[246]), .Z(n37776) );
  NANDN U38088 ( .A(n37776), .B(n38325), .Z(n37681) );
  NANDN U38089 ( .A(n37679), .B(n38326), .Z(n37680) );
  AND U38090 ( .A(n37681), .B(n37680), .Z(n37768) );
  XNOR U38091 ( .A(n37767), .B(n37768), .Z(n37769) );
  XNOR U38092 ( .A(n37770), .B(n37769), .Z(n37796) );
  XOR U38093 ( .A(a[250]), .B(n1056), .Z(n37785) );
  NANDN U38094 ( .A(n37785), .B(n38101), .Z(n37684) );
  NANDN U38095 ( .A(n37682), .B(n38102), .Z(n37683) );
  NAND U38096 ( .A(n37684), .B(n37683), .Z(n37753) );
  NANDN U38097 ( .A(n37685), .B(n38205), .Z(n37687) );
  XOR U38098 ( .A(b[23]), .B(n38272), .Z(n37756) );
  OR U38099 ( .A(n37756), .B(n38268), .Z(n37686) );
  NAND U38100 ( .A(n37687), .B(n37686), .Z(n37750) );
  NAND U38101 ( .A(n37688), .B(n37762), .Z(n37690) );
  XNOR U38102 ( .A(a[254]), .B(b[17]), .Z(n37763) );
  NANDN U38103 ( .A(n37763), .B(n37764), .Z(n37689) );
  AND U38104 ( .A(n37690), .B(n37689), .Z(n37751) );
  XNOR U38105 ( .A(n37750), .B(n37751), .Z(n37752) );
  XNOR U38106 ( .A(n37753), .B(n37752), .Z(n37793) );
  XOR U38107 ( .A(a[252]), .B(n1055), .Z(n37759) );
  NANDN U38108 ( .A(n37759), .B(n37934), .Z(n37693) );
  NAND U38109 ( .A(n37935), .B(n37691), .Z(n37692) );
  NAND U38110 ( .A(n37693), .B(n37692), .Z(n37794) );
  XNOR U38111 ( .A(n37793), .B(n37794), .Z(n37795) );
  XOR U38112 ( .A(n37796), .B(n37795), .Z(n37747) );
  NANDN U38113 ( .A(n37695), .B(n37694), .Z(n37699) );
  NAND U38114 ( .A(n37697), .B(n37696), .Z(n37698) );
  NAND U38115 ( .A(n37699), .B(n37698), .Z(n37744) );
  NANDN U38116 ( .A(n37701), .B(n37700), .Z(n37705) );
  NAND U38117 ( .A(n37703), .B(n37702), .Z(n37704) );
  AND U38118 ( .A(n37705), .B(n37704), .Z(n37745) );
  XNOR U38119 ( .A(n37744), .B(n37745), .Z(n37746) );
  XOR U38120 ( .A(n37747), .B(n37746), .Z(n37737) );
  XNOR U38121 ( .A(n37736), .B(n37737), .Z(n37731) );
  XNOR U38122 ( .A(n37730), .B(n37731), .Z(n37724) );
  NAND U38123 ( .A(n37707), .B(n37706), .Z(n37711) );
  NAND U38124 ( .A(n37709), .B(n37708), .Z(n37710) );
  NAND U38125 ( .A(n37711), .B(n37710), .Z(n37725) );
  XNOR U38126 ( .A(n37724), .B(n37725), .Z(n37726) );
  XNOR U38127 ( .A(n37726), .B(n37727), .Z(n37800) );
  IV U38128 ( .A(n37800), .Z(n37799) );
  XOR U38129 ( .A(n37799), .B(n37802), .Z(n37719) );
  XNOR U38130 ( .A(n37801), .B(n37719), .Z(n37722) );
  OR U38131 ( .A(n37721), .B(n37720), .Z(n37723) );
  XNOR U38132 ( .A(n37722), .B(n37723), .Z(c[494]) );
  NANDN U38133 ( .A(n37723), .B(n37722), .Z(n37884) );
  NANDN U38134 ( .A(n37729), .B(n37728), .Z(n37733) );
  NAND U38135 ( .A(n37731), .B(n37730), .Z(n37732) );
  NAND U38136 ( .A(n37733), .B(n37732), .Z(n37879) );
  NANDN U38137 ( .A(n37739), .B(n37738), .Z(n37743) );
  NAND U38138 ( .A(n37741), .B(n37740), .Z(n37742) );
  NAND U38139 ( .A(n37743), .B(n37742), .Z(n37871) );
  NANDN U38140 ( .A(n37745), .B(n37744), .Z(n37749) );
  NANDN U38141 ( .A(n37747), .B(n37746), .Z(n37748) );
  AND U38142 ( .A(n37749), .B(n37748), .Z(n37872) );
  XNOR U38143 ( .A(n37871), .B(n37872), .Z(n37873) );
  NANDN U38144 ( .A(n37751), .B(n37750), .Z(n37755) );
  NAND U38145 ( .A(n37753), .B(n37752), .Z(n37754) );
  NAND U38146 ( .A(n37755), .B(n37754), .Z(n37863) );
  NANDN U38147 ( .A(n37756), .B(n38205), .Z(n37758) );
  XNOR U38148 ( .A(n1057), .B(a[249]), .Z(n37842) );
  NANDN U38149 ( .A(n38268), .B(n37842), .Z(n37757) );
  NAND U38150 ( .A(n37758), .B(n37757), .Z(n37810) );
  XNOR U38151 ( .A(a[253]), .B(n1055), .Z(n37816) );
  NAND U38152 ( .A(n37816), .B(n37934), .Z(n37761) );
  NANDN U38153 ( .A(n37759), .B(n37935), .Z(n37760) );
  NAND U38154 ( .A(n37761), .B(n37760), .Z(n37807) );
  NANDN U38155 ( .A(n37763), .B(n37762), .Z(n37766) );
  XNOR U38156 ( .A(n38595), .B(b[17]), .Z(n37824) );
  NAND U38157 ( .A(n37824), .B(n37764), .Z(n37765) );
  AND U38158 ( .A(n37766), .B(n37765), .Z(n37808) );
  XNOR U38159 ( .A(n37807), .B(n37808), .Z(n37809) );
  XNOR U38160 ( .A(n37810), .B(n37809), .Z(n37861) );
  NANDN U38161 ( .A(n37768), .B(n37767), .Z(n37772) );
  NAND U38162 ( .A(n37770), .B(n37769), .Z(n37771) );
  NAND U38163 ( .A(n37772), .B(n37771), .Z(n37862) );
  XOR U38164 ( .A(n37861), .B(n37862), .Z(n37864) );
  XNOR U38165 ( .A(n37863), .B(n37864), .Z(n37870) );
  XNOR U38166 ( .A(n1059), .B(a[241]), .Z(n37827) );
  NAND U38167 ( .A(n37827), .B(n38552), .Z(n37775) );
  NANDN U38168 ( .A(n37773), .B(n38553), .Z(n37774) );
  NAND U38169 ( .A(n37775), .B(n37774), .Z(n37830) );
  XOR U38170 ( .A(b[25]), .B(a[247]), .Z(n37848) );
  NAND U38171 ( .A(n37848), .B(n38325), .Z(n37778) );
  NANDN U38172 ( .A(n37776), .B(n38326), .Z(n37777) );
  AND U38173 ( .A(n37778), .B(n37777), .Z(n37831) );
  XNOR U38174 ( .A(n37830), .B(n37831), .Z(n37832) );
  NANDN U38175 ( .A(n1059), .B(a[239]), .Z(n37852) );
  XNOR U38176 ( .A(n37851), .B(n37852), .Z(n37854) );
  XOR U38177 ( .A(n37853), .B(n37854), .Z(n37833) );
  XOR U38178 ( .A(n37832), .B(n37833), .Z(n37860) );
  XNOR U38179 ( .A(b[27]), .B(n38213), .Z(n37819) );
  NAND U38180 ( .A(n38423), .B(n37819), .Z(n37781) );
  NANDN U38181 ( .A(n37779), .B(n38424), .Z(n37780) );
  NAND U38182 ( .A(n37781), .B(n37780), .Z(n37839) );
  NAND U38183 ( .A(n38490), .B(n37782), .Z(n37784) );
  XOR U38184 ( .A(b[29]), .B(n38110), .Z(n37845) );
  OR U38185 ( .A(n37845), .B(n1048), .Z(n37783) );
  NAND U38186 ( .A(n37784), .B(n37783), .Z(n37836) );
  XNOR U38187 ( .A(a[251]), .B(n1056), .Z(n37813) );
  NAND U38188 ( .A(n37813), .B(n38101), .Z(n37787) );
  NANDN U38189 ( .A(n37785), .B(n38102), .Z(n37786) );
  AND U38190 ( .A(n37787), .B(n37786), .Z(n37837) );
  XNOR U38191 ( .A(n37836), .B(n37837), .Z(n37838) );
  XNOR U38192 ( .A(n37839), .B(n37838), .Z(n37857) );
  OR U38193 ( .A(n37853), .B(n37788), .Z(n37792) );
  NAND U38194 ( .A(n37790), .B(n37789), .Z(n37791) );
  NAND U38195 ( .A(n37792), .B(n37791), .Z(n37858) );
  XNOR U38196 ( .A(n37857), .B(n37858), .Z(n37859) );
  XNOR U38197 ( .A(n37860), .B(n37859), .Z(n37867) );
  NANDN U38198 ( .A(n37794), .B(n37793), .Z(n37798) );
  NAND U38199 ( .A(n37796), .B(n37795), .Z(n37797) );
  NAND U38200 ( .A(n37798), .B(n37797), .Z(n37868) );
  XNOR U38201 ( .A(n37867), .B(n37868), .Z(n37869) );
  XNOR U38202 ( .A(n37870), .B(n37869), .Z(n37874) );
  XNOR U38203 ( .A(n37873), .B(n37874), .Z(n37877) );
  XNOR U38204 ( .A(n37878), .B(n37877), .Z(n37880) );
  XOR U38205 ( .A(n37879), .B(n37880), .Z(n37804) );
  XNOR U38206 ( .A(n37804), .B(n37806), .Z(n37803) );
  XNOR U38207 ( .A(n37805), .B(n37803), .Z(n37883) );
  XNOR U38208 ( .A(n37884), .B(n37883), .Z(c[495]) );
  NANDN U38209 ( .A(n37808), .B(n37807), .Z(n37812) );
  NAND U38210 ( .A(n37810), .B(n37809), .Z(n37811) );
  NAND U38211 ( .A(n37812), .B(n37811), .Z(n37924) );
  XOR U38212 ( .A(n38531), .B(b[21]), .Z(n37954) );
  NANDN U38213 ( .A(n37954), .B(n38101), .Z(n37815) );
  NAND U38214 ( .A(n38102), .B(n37813), .Z(n37814) );
  NAND U38215 ( .A(n37815), .B(n37814), .Z(n37913) );
  XOR U38216 ( .A(a[254]), .B(n1055), .Z(n37936) );
  NANDN U38217 ( .A(n37936), .B(n37934), .Z(n37818) );
  NAND U38218 ( .A(n37935), .B(n37816), .Z(n37817) );
  NAND U38219 ( .A(n37818), .B(n37817), .Z(n37911) );
  XNOR U38220 ( .A(b[27]), .B(a[246]), .Z(n37939) );
  NANDN U38221 ( .A(n37939), .B(n38423), .Z(n37821) );
  NAND U38222 ( .A(n38424), .B(n37819), .Z(n37820) );
  NAND U38223 ( .A(n37821), .B(n37820), .Z(n37912) );
  XOR U38224 ( .A(n37911), .B(n37912), .Z(n37914) );
  XNOR U38225 ( .A(n37913), .B(n37914), .Z(n37922) );
  XNOR U38226 ( .A(b[17]), .B(n37822), .Z(n37826) );
  XOR U38227 ( .A(b[16]), .B(n1054), .Z(n37823) );
  NANDN U38228 ( .A(n37824), .B(n37823), .Z(n37825) );
  AND U38229 ( .A(n37826), .B(n37825), .Z(n37918) );
  AND U38230 ( .A(a[240]), .B(b[31]), .Z(n38026) );
  XOR U38231 ( .A(n1059), .B(a[242]), .Z(n37951) );
  NANDN U38232 ( .A(n37951), .B(n38552), .Z(n37829) );
  NAND U38233 ( .A(n38553), .B(n37827), .Z(n37828) );
  NAND U38234 ( .A(n37829), .B(n37828), .Z(n37917) );
  XNOR U38235 ( .A(n38026), .B(n37917), .Z(n37919) );
  XOR U38236 ( .A(n37918), .B(n37919), .Z(n37923) );
  XOR U38237 ( .A(n37922), .B(n37923), .Z(n37925) );
  XNOR U38238 ( .A(n37924), .B(n37925), .Z(n37899) );
  NANDN U38239 ( .A(n37831), .B(n37830), .Z(n37835) );
  NANDN U38240 ( .A(n37833), .B(n37832), .Z(n37834) );
  AND U38241 ( .A(n37835), .B(n37834), .Z(n37900) );
  XNOR U38242 ( .A(n37899), .B(n37900), .Z(n37901) );
  NANDN U38243 ( .A(n37837), .B(n37836), .Z(n37841) );
  NAND U38244 ( .A(n37839), .B(n37838), .Z(n37840) );
  NAND U38245 ( .A(n37841), .B(n37840), .Z(n37908) );
  XOR U38246 ( .A(a[250]), .B(n1057), .Z(n37945) );
  OR U38247 ( .A(n37945), .B(n38268), .Z(n37844) );
  NAND U38248 ( .A(n38205), .B(n37842), .Z(n37843) );
  NAND U38249 ( .A(n37844), .B(n37843), .Z(n37929) );
  NANDN U38250 ( .A(n37845), .B(n38490), .Z(n37847) );
  XNOR U38251 ( .A(n1058), .B(a[244]), .Z(n37942) );
  NANDN U38252 ( .A(n1048), .B(n37942), .Z(n37846) );
  AND U38253 ( .A(n37847), .B(n37846), .Z(n37928) );
  XNOR U38254 ( .A(n37929), .B(n37928), .Z(n37930) );
  XOR U38255 ( .A(b[25]), .B(n38272), .Z(n37948) );
  NANDN U38256 ( .A(n37948), .B(n38325), .Z(n37850) );
  NAND U38257 ( .A(n38326), .B(n37848), .Z(n37849) );
  NAND U38258 ( .A(n37850), .B(n37849), .Z(n37931) );
  XOR U38259 ( .A(n37930), .B(n37931), .Z(n37905) );
  OR U38260 ( .A(n37852), .B(n37851), .Z(n37856) );
  NANDN U38261 ( .A(n37854), .B(n37853), .Z(n37855) );
  AND U38262 ( .A(n37856), .B(n37855), .Z(n37906) );
  XNOR U38263 ( .A(n37905), .B(n37906), .Z(n37907) );
  XNOR U38264 ( .A(n37908), .B(n37907), .Z(n37902) );
  XOR U38265 ( .A(n37901), .B(n37902), .Z(n37896) );
  NANDN U38266 ( .A(n37862), .B(n37861), .Z(n37866) );
  OR U38267 ( .A(n37864), .B(n37863), .Z(n37865) );
  AND U38268 ( .A(n37866), .B(n37865), .Z(n37894) );
  XNOR U38269 ( .A(n37893), .B(n37894), .Z(n37895) );
  XNOR U38270 ( .A(n37896), .B(n37895), .Z(n37958) );
  XNOR U38271 ( .A(n37958), .B(n37957), .Z(n37959) );
  NANDN U38272 ( .A(n37872), .B(n37871), .Z(n37876) );
  NANDN U38273 ( .A(n37874), .B(n37873), .Z(n37875) );
  NAND U38274 ( .A(n37876), .B(n37875), .Z(n37960) );
  XOR U38275 ( .A(n37959), .B(n37960), .Z(n37887) );
  NAND U38276 ( .A(n37878), .B(n37877), .Z(n37882) );
  NANDN U38277 ( .A(n37880), .B(n37879), .Z(n37881) );
  AND U38278 ( .A(n37882), .B(n37881), .Z(n37888) );
  XNOR U38279 ( .A(n37887), .B(n37888), .Z(n37889) );
  XNOR U38280 ( .A(n37890), .B(n37889), .Z(n37885) );
  NANDN U38281 ( .A(n37884), .B(n37883), .Z(n37886) );
  XNOR U38282 ( .A(n37885), .B(n37886), .Z(c[496]) );
  NANDN U38283 ( .A(n37886), .B(n37885), .Z(n38039) );
  NANDN U38284 ( .A(n37888), .B(n37887), .Z(n37892) );
  NANDN U38285 ( .A(n37890), .B(n37889), .Z(n37891) );
  AND U38286 ( .A(n37892), .B(n37891), .Z(n37966) );
  NANDN U38287 ( .A(n37894), .B(n37893), .Z(n37898) );
  NAND U38288 ( .A(n37896), .B(n37895), .Z(n37897) );
  NAND U38289 ( .A(n37898), .B(n37897), .Z(n37970) );
  NANDN U38290 ( .A(n37900), .B(n37899), .Z(n37904) );
  NANDN U38291 ( .A(n37902), .B(n37901), .Z(n37903) );
  NAND U38292 ( .A(n37904), .B(n37903), .Z(n37967) );
  NANDN U38293 ( .A(n37906), .B(n37905), .Z(n37910) );
  NAND U38294 ( .A(n37908), .B(n37907), .Z(n37909) );
  NAND U38295 ( .A(n37910), .B(n37909), .Z(n37981) );
  NAND U38296 ( .A(n37912), .B(n37911), .Z(n37916) );
  NAND U38297 ( .A(n37914), .B(n37913), .Z(n37915) );
  NAND U38298 ( .A(n37916), .B(n37915), .Z(n37979) );
  NANDN U38299 ( .A(n38026), .B(n37917), .Z(n37921) );
  NAND U38300 ( .A(n37919), .B(n37918), .Z(n37920) );
  NAND U38301 ( .A(n37921), .B(n37920), .Z(n37980) );
  XOR U38302 ( .A(n37979), .B(n37980), .Z(n37982) );
  XNOR U38303 ( .A(n37981), .B(n37982), .Z(n37976) );
  NANDN U38304 ( .A(n37923), .B(n37922), .Z(n37927) );
  OR U38305 ( .A(n37925), .B(n37924), .Z(n37926) );
  NAND U38306 ( .A(n37927), .B(n37926), .Z(n37973) );
  NANDN U38307 ( .A(n37929), .B(n37928), .Z(n37933) );
  NANDN U38308 ( .A(n37931), .B(n37930), .Z(n37932) );
  NAND U38309 ( .A(n37933), .B(n37932), .Z(n37988) );
  XNOR U38310 ( .A(n38595), .B(b[19]), .Z(n38031) );
  NAND U38311 ( .A(n38031), .B(n37934), .Z(n37938) );
  NANDN U38312 ( .A(n37936), .B(n37935), .Z(n37937) );
  NAND U38313 ( .A(n37938), .B(n37937), .Z(n38018) );
  XOR U38314 ( .A(b[27]), .B(a[247]), .Z(n38009) );
  NAND U38315 ( .A(n38423), .B(n38009), .Z(n37941) );
  NANDN U38316 ( .A(n37939), .B(n38424), .Z(n37940) );
  AND U38317 ( .A(n37941), .B(n37940), .Z(n38019) );
  XNOR U38318 ( .A(n38018), .B(n38019), .Z(n38020) );
  NANDN U38319 ( .A(n1059), .B(a[241]), .Z(n38024) );
  XOR U38320 ( .A(n38025), .B(n38024), .Z(n38027) );
  XNOR U38321 ( .A(n38026), .B(n38027), .Z(n38021) );
  XOR U38322 ( .A(n38020), .B(n38021), .Z(n37985) );
  NAND U38323 ( .A(n37942), .B(n38490), .Z(n37944) );
  XOR U38324 ( .A(n1058), .B(n38213), .Z(n38006) );
  NANDN U38325 ( .A(n1048), .B(n38006), .Z(n37943) );
  NAND U38326 ( .A(n37944), .B(n37943), .Z(n37994) );
  NANDN U38327 ( .A(n37945), .B(n38205), .Z(n37947) );
  XNOR U38328 ( .A(a[251]), .B(b[23]), .Z(n38015) );
  OR U38329 ( .A(n38015), .B(n38268), .Z(n37946) );
  NAND U38330 ( .A(n37947), .B(n37946), .Z(n37991) );
  XOR U38331 ( .A(b[25]), .B(a[249]), .Z(n38003) );
  NAND U38332 ( .A(n38325), .B(n38003), .Z(n37950) );
  NANDN U38333 ( .A(n37948), .B(n38326), .Z(n37949) );
  NAND U38334 ( .A(n37950), .B(n37949), .Z(n37998) );
  XOR U38335 ( .A(b[31]), .B(n38110), .Z(n38035) );
  NANDN U38336 ( .A(n38035), .B(n38552), .Z(n37953) );
  NANDN U38337 ( .A(n37951), .B(n38553), .Z(n37952) );
  AND U38338 ( .A(n37953), .B(n37952), .Z(n37997) );
  XNOR U38339 ( .A(n37998), .B(n37997), .Z(n37999) );
  XNOR U38340 ( .A(a[253]), .B(b[21]), .Z(n38012) );
  NANDN U38341 ( .A(n38012), .B(n38101), .Z(n37956) );
  NANDN U38342 ( .A(n37954), .B(n38102), .Z(n37955) );
  NAND U38343 ( .A(n37956), .B(n37955), .Z(n38000) );
  XNOR U38344 ( .A(n37999), .B(n38000), .Z(n37992) );
  XNOR U38345 ( .A(n37991), .B(n37992), .Z(n37993) );
  XOR U38346 ( .A(n37994), .B(n37993), .Z(n37986) );
  XNOR U38347 ( .A(n37985), .B(n37986), .Z(n37987) );
  XNOR U38348 ( .A(n37988), .B(n37987), .Z(n37974) );
  XNOR U38349 ( .A(n37973), .B(n37974), .Z(n37975) );
  XOR U38350 ( .A(n37976), .B(n37975), .Z(n37968) );
  XNOR U38351 ( .A(n37967), .B(n37968), .Z(n37969) );
  XOR U38352 ( .A(n37970), .B(n37969), .Z(n37964) );
  NANDN U38353 ( .A(n37958), .B(n37957), .Z(n37962) );
  NANDN U38354 ( .A(n37960), .B(n37959), .Z(n37961) );
  AND U38355 ( .A(n37962), .B(n37961), .Z(n37965) );
  XOR U38356 ( .A(n37964), .B(n37965), .Z(n37963) );
  XOR U38357 ( .A(n37966), .B(n37963), .Z(n38038) );
  XNOR U38358 ( .A(n38039), .B(n38038), .Z(c[497]) );
  NANDN U38359 ( .A(n37968), .B(n37967), .Z(n37972) );
  NANDN U38360 ( .A(n37970), .B(n37969), .Z(n37971) );
  NAND U38361 ( .A(n37972), .B(n37971), .Z(n38043) );
  NANDN U38362 ( .A(n37974), .B(n37973), .Z(n37978) );
  NAND U38363 ( .A(n37976), .B(n37975), .Z(n37977) );
  NAND U38364 ( .A(n37978), .B(n37977), .Z(n38051) );
  NAND U38365 ( .A(n37980), .B(n37979), .Z(n37984) );
  NAND U38366 ( .A(n37982), .B(n37981), .Z(n37983) );
  NAND U38367 ( .A(n37984), .B(n37983), .Z(n38049) );
  NANDN U38368 ( .A(n37986), .B(n37985), .Z(n37990) );
  NAND U38369 ( .A(n37988), .B(n37987), .Z(n37989) );
  NAND U38370 ( .A(n37990), .B(n37989), .Z(n38057) );
  NANDN U38371 ( .A(n37992), .B(n37991), .Z(n37996) );
  NAND U38372 ( .A(n37994), .B(n37993), .Z(n37995) );
  NAND U38373 ( .A(n37996), .B(n37995), .Z(n38055) );
  NANDN U38374 ( .A(n37998), .B(n37997), .Z(n38002) );
  NANDN U38375 ( .A(n38000), .B(n37999), .Z(n38001) );
  NAND U38376 ( .A(n38002), .B(n38001), .Z(n38060) );
  XNOR U38377 ( .A(b[25]), .B(n38356), .Z(n38098) );
  NAND U38378 ( .A(n38098), .B(n38325), .Z(n38005) );
  NAND U38379 ( .A(n38003), .B(n38326), .Z(n38004) );
  NAND U38380 ( .A(n38005), .B(n38004), .Z(n38086) );
  NAND U38381 ( .A(n38490), .B(n38006), .Z(n38008) );
  XOR U38382 ( .A(n1058), .B(n38146), .Z(n38089) );
  NANDN U38383 ( .A(n1048), .B(n38089), .Z(n38007) );
  NAND U38384 ( .A(n38008), .B(n38007), .Z(n38083) );
  XNOR U38385 ( .A(b[27]), .B(a[248]), .Z(n38106) );
  NANDN U38386 ( .A(n38106), .B(n38423), .Z(n38011) );
  NAND U38387 ( .A(n38009), .B(n38424), .Z(n38010) );
  AND U38388 ( .A(n38011), .B(n38010), .Z(n38084) );
  XNOR U38389 ( .A(n38083), .B(n38084), .Z(n38085) );
  XNOR U38390 ( .A(n38086), .B(n38085), .Z(n38069) );
  XOR U38391 ( .A(a[254]), .B(n1056), .Z(n38103) );
  NANDN U38392 ( .A(n38103), .B(n38101), .Z(n38014) );
  NANDN U38393 ( .A(n38012), .B(n38102), .Z(n38013) );
  NAND U38394 ( .A(n38014), .B(n38013), .Z(n38066) );
  NANDN U38395 ( .A(n38015), .B(n38205), .Z(n38017) );
  XOR U38396 ( .A(n38531), .B(n1057), .Z(n38095) );
  NANDN U38397 ( .A(n38268), .B(n38095), .Z(n38016) );
  AND U38398 ( .A(n38017), .B(n38016), .Z(n38067) );
  XNOR U38399 ( .A(n38066), .B(n38067), .Z(n38068) );
  XOR U38400 ( .A(n38069), .B(n38068), .Z(n38061) );
  XOR U38401 ( .A(n38060), .B(n38061), .Z(n38062) );
  NANDN U38402 ( .A(n38019), .B(n38018), .Z(n38023) );
  NANDN U38403 ( .A(n38021), .B(n38020), .Z(n38022) );
  NAND U38404 ( .A(n38023), .B(n38022), .Z(n38074) );
  OR U38405 ( .A(n38025), .B(n38024), .Z(n38029) );
  NAND U38406 ( .A(n38027), .B(n38026), .Z(n38028) );
  NAND U38407 ( .A(n38029), .B(n38028), .Z(n38073) );
  NAND U38408 ( .A(b[18]), .B(b[17]), .Z(n38109) );
  XOR U38409 ( .A(n1055), .B(n38109), .Z(n38033) );
  XNOR U38410 ( .A(b[18]), .B(b[17]), .Z(n38030) );
  NANDN U38411 ( .A(n38031), .B(n38030), .Z(n38032) );
  AND U38412 ( .A(n38033), .B(n38032), .Z(n38079) );
  AND U38413 ( .A(a[242]), .B(b[31]), .Z(n38162) );
  XOR U38414 ( .A(n1059), .B(n38034), .Z(n38092) );
  NAND U38415 ( .A(n38092), .B(n38552), .Z(n38037) );
  NANDN U38416 ( .A(n38035), .B(n38553), .Z(n38036) );
  AND U38417 ( .A(n38037), .B(n38036), .Z(n38078) );
  XOR U38418 ( .A(n38162), .B(n38078), .Z(n38080) );
  XOR U38419 ( .A(n38079), .B(n38080), .Z(n38072) );
  XNOR U38420 ( .A(n38073), .B(n38072), .Z(n38075) );
  XNOR U38421 ( .A(n38074), .B(n38075), .Z(n38063) );
  XOR U38422 ( .A(n38062), .B(n38063), .Z(n38054) );
  XNOR U38423 ( .A(n38055), .B(n38054), .Z(n38056) );
  XOR U38424 ( .A(n38057), .B(n38056), .Z(n38048) );
  XOR U38425 ( .A(n38049), .B(n38048), .Z(n38050) );
  XNOR U38426 ( .A(n38051), .B(n38050), .Z(n38042) );
  XOR U38427 ( .A(n38043), .B(n38042), .Z(n38044) );
  XNOR U38428 ( .A(n38045), .B(n38044), .Z(n38040) );
  NANDN U38429 ( .A(n38039), .B(n38038), .Z(n38041) );
  XNOR U38430 ( .A(n38040), .B(n38041), .Z(c[498]) );
  NANDN U38431 ( .A(n38041), .B(n38040), .Z(n38113) );
  NAND U38432 ( .A(n38043), .B(n38042), .Z(n38047) );
  NANDN U38433 ( .A(n38045), .B(n38044), .Z(n38046) );
  NAND U38434 ( .A(n38047), .B(n38046), .Z(n38116) );
  NAND U38435 ( .A(n38049), .B(n38048), .Z(n38053) );
  NANDN U38436 ( .A(n38051), .B(n38050), .Z(n38052) );
  AND U38437 ( .A(n38053), .B(n38052), .Z(n38115) );
  NAND U38438 ( .A(n38055), .B(n38054), .Z(n38059) );
  OR U38439 ( .A(n38057), .B(n38056), .Z(n38058) );
  NAND U38440 ( .A(n38059), .B(n38058), .Z(n38120) );
  OR U38441 ( .A(n38061), .B(n38060), .Z(n38065) );
  NAND U38442 ( .A(n38063), .B(n38062), .Z(n38064) );
  NAND U38443 ( .A(n38065), .B(n38064), .Z(n38118) );
  NANDN U38444 ( .A(n38067), .B(n38066), .Z(n38071) );
  NANDN U38445 ( .A(n38069), .B(n38068), .Z(n38070) );
  NAND U38446 ( .A(n38071), .B(n38070), .Z(n38123) );
  NAND U38447 ( .A(n38073), .B(n38072), .Z(n38077) );
  NANDN U38448 ( .A(n38075), .B(n38074), .Z(n38076) );
  AND U38449 ( .A(n38077), .B(n38076), .Z(n38124) );
  XNOR U38450 ( .A(n38123), .B(n38124), .Z(n38125) );
  OR U38451 ( .A(n38162), .B(n38078), .Z(n38082) );
  NAND U38452 ( .A(n38080), .B(n38079), .Z(n38081) );
  NAND U38453 ( .A(n38082), .B(n38081), .Z(n38174) );
  NANDN U38454 ( .A(n38084), .B(n38083), .Z(n38088) );
  NAND U38455 ( .A(n38086), .B(n38085), .Z(n38087) );
  AND U38456 ( .A(n38088), .B(n38087), .Z(n38175) );
  XNOR U38457 ( .A(n38174), .B(n38175), .Z(n38176) );
  NAND U38458 ( .A(n38490), .B(n38089), .Z(n38091) );
  XNOR U38459 ( .A(b[29]), .B(a[247]), .Z(n38138) );
  OR U38460 ( .A(n38138), .B(n1048), .Z(n38090) );
  NAND U38461 ( .A(n38091), .B(n38090), .Z(n38150) );
  XOR U38462 ( .A(n1059), .B(a[245]), .Z(n38147) );
  NANDN U38463 ( .A(n38147), .B(n38552), .Z(n38094) );
  NAND U38464 ( .A(n38553), .B(n38092), .Z(n38093) );
  NAND U38465 ( .A(n38094), .B(n38093), .Z(n38157) );
  XNOR U38466 ( .A(a[253]), .B(b[23]), .Z(n38132) );
  OR U38467 ( .A(n38132), .B(n38268), .Z(n38097) );
  NAND U38468 ( .A(n38205), .B(n38095), .Z(n38096) );
  AND U38469 ( .A(n38097), .B(n38096), .Z(n38156) );
  XNOR U38470 ( .A(n38157), .B(n38156), .Z(n38158) );
  XOR U38471 ( .A(b[25]), .B(a[251]), .Z(n38129) );
  NAND U38472 ( .A(n38325), .B(n38129), .Z(n38100) );
  NAND U38473 ( .A(n38326), .B(n38098), .Z(n38099) );
  NAND U38474 ( .A(n38100), .B(n38099), .Z(n38159) );
  XNOR U38475 ( .A(n38158), .B(n38159), .Z(n38151) );
  XNOR U38476 ( .A(n38150), .B(n38151), .Z(n38152) );
  XNOR U38477 ( .A(n38595), .B(b[21]), .Z(n38143) );
  NAND U38478 ( .A(n38143), .B(n38101), .Z(n38105) );
  NANDN U38479 ( .A(n38103), .B(n38102), .Z(n38104) );
  NAND U38480 ( .A(n38105), .B(n38104), .Z(n38168) );
  XOR U38481 ( .A(b[27]), .B(a[249]), .Z(n38135) );
  NAND U38482 ( .A(n38423), .B(n38135), .Z(n38108) );
  NANDN U38483 ( .A(n38106), .B(n38424), .Z(n38107) );
  AND U38484 ( .A(n38108), .B(n38107), .Z(n38169) );
  XNOR U38485 ( .A(n38168), .B(n38169), .Z(n38170) );
  ANDN U38486 ( .B(n38109), .A(n1055), .Z(n38163) );
  XOR U38487 ( .A(n38163), .B(n38162), .Z(n38165) );
  NANDN U38488 ( .A(n38110), .B(b[31]), .Z(n38164) );
  XOR U38489 ( .A(n38165), .B(n38164), .Z(n38171) );
  XOR U38490 ( .A(n38170), .B(n38171), .Z(n38153) );
  XOR U38491 ( .A(n38152), .B(n38153), .Z(n38177) );
  XOR U38492 ( .A(n38176), .B(n38177), .Z(n38126) );
  XOR U38493 ( .A(n38125), .B(n38126), .Z(n38117) );
  XOR U38494 ( .A(n38118), .B(n38117), .Z(n38119) );
  XOR U38495 ( .A(n38120), .B(n38119), .Z(n38114) );
  XNOR U38496 ( .A(n38115), .B(n38114), .Z(n38111) );
  XOR U38497 ( .A(n38116), .B(n38111), .Z(n38112) );
  XNOR U38498 ( .A(n38113), .B(n38112), .Z(c[499]) );
  NANDN U38499 ( .A(n38113), .B(n38112), .Z(n38234) );
  NAND U38500 ( .A(n38118), .B(n38117), .Z(n38122) );
  NAND U38501 ( .A(n38120), .B(n38119), .Z(n38121) );
  AND U38502 ( .A(n38122), .B(n38121), .Z(n38182) );
  NANDN U38503 ( .A(n38124), .B(n38123), .Z(n38128) );
  NAND U38504 ( .A(n38126), .B(n38125), .Z(n38127) );
  NAND U38505 ( .A(n38128), .B(n38127), .Z(n38187) );
  XNOR U38506 ( .A(a[252]), .B(b[25]), .Z(n38214) );
  NANDN U38507 ( .A(n38214), .B(n38325), .Z(n38131) );
  NAND U38508 ( .A(n38129), .B(n38326), .Z(n38130) );
  NAND U38509 ( .A(n38131), .B(n38130), .Z(n38202) );
  NANDN U38510 ( .A(n38132), .B(n38205), .Z(n38134) );
  XOR U38511 ( .A(a[254]), .B(n1057), .Z(n38206) );
  OR U38512 ( .A(n38206), .B(n38268), .Z(n38133) );
  NAND U38513 ( .A(n38134), .B(n38133), .Z(n38199) );
  XNOR U38514 ( .A(b[27]), .B(a[250]), .Z(n38209) );
  NANDN U38515 ( .A(n38209), .B(n38423), .Z(n38137) );
  NAND U38516 ( .A(n38135), .B(n38424), .Z(n38136) );
  AND U38517 ( .A(n38137), .B(n38136), .Z(n38200) );
  XNOR U38518 ( .A(n38199), .B(n38200), .Z(n38201) );
  XNOR U38519 ( .A(n38202), .B(n38201), .Z(n38223) );
  NANDN U38520 ( .A(n38138), .B(n38490), .Z(n38140) );
  XNOR U38521 ( .A(n1058), .B(a[248]), .Z(n38217) );
  NANDN U38522 ( .A(n1048), .B(n38217), .Z(n38139) );
  NAND U38523 ( .A(n38140), .B(n38139), .Z(n38224) );
  XNOR U38524 ( .A(n38223), .B(n38224), .Z(n38225) );
  XOR U38525 ( .A(n1056), .B(n38212), .Z(n38145) );
  XOR U38526 ( .A(n38141), .B(b[19]), .Z(n38142) );
  NANDN U38527 ( .A(n38143), .B(n38142), .Z(n38144) );
  AND U38528 ( .A(n38145), .B(n38144), .Z(n38196) );
  AND U38529 ( .A(a[244]), .B(b[31]), .Z(n38290) );
  XNOR U38530 ( .A(n38196), .B(n38290), .Z(n38197) );
  XOR U38531 ( .A(b[31]), .B(n38146), .Z(n38220) );
  NANDN U38532 ( .A(n38220), .B(n38552), .Z(n38149) );
  NANDN U38533 ( .A(n38147), .B(n38553), .Z(n38148) );
  AND U38534 ( .A(n38149), .B(n38148), .Z(n38198) );
  XNOR U38535 ( .A(n38197), .B(n38198), .Z(n38226) );
  XNOR U38536 ( .A(n38225), .B(n38226), .Z(n38190) );
  NANDN U38537 ( .A(n38151), .B(n38150), .Z(n38155) );
  NAND U38538 ( .A(n38153), .B(n38152), .Z(n38154) );
  AND U38539 ( .A(n38155), .B(n38154), .Z(n38191) );
  XNOR U38540 ( .A(n38190), .B(n38191), .Z(n38193) );
  NANDN U38541 ( .A(n38157), .B(n38156), .Z(n38161) );
  NANDN U38542 ( .A(n38159), .B(n38158), .Z(n38160) );
  NAND U38543 ( .A(n38161), .B(n38160), .Z(n38230) );
  NANDN U38544 ( .A(n38163), .B(n38162), .Z(n38167) );
  OR U38545 ( .A(n38165), .B(n38164), .Z(n38166) );
  NAND U38546 ( .A(n38167), .B(n38166), .Z(n38228) );
  NANDN U38547 ( .A(n38169), .B(n38168), .Z(n38173) );
  NAND U38548 ( .A(n38171), .B(n38170), .Z(n38172) );
  AND U38549 ( .A(n38173), .B(n38172), .Z(n38227) );
  XNOR U38550 ( .A(n38228), .B(n38227), .Z(n38229) );
  XNOR U38551 ( .A(n38230), .B(n38229), .Z(n38192) );
  XNOR U38552 ( .A(n38193), .B(n38192), .Z(n38184) );
  NANDN U38553 ( .A(n38175), .B(n38174), .Z(n38179) );
  NAND U38554 ( .A(n38177), .B(n38176), .Z(n38178) );
  AND U38555 ( .A(n38179), .B(n38178), .Z(n38185) );
  XNOR U38556 ( .A(n38184), .B(n38185), .Z(n38186) );
  XOR U38557 ( .A(n38187), .B(n38186), .Z(n38181) );
  XNOR U38558 ( .A(n38182), .B(n38181), .Z(n38180) );
  XOR U38559 ( .A(n38183), .B(n38180), .Z(n38233) );
  XNOR U38560 ( .A(n38234), .B(n38233), .Z(c[500]) );
  NANDN U38561 ( .A(n38185), .B(n38184), .Z(n38189) );
  NAND U38562 ( .A(n38187), .B(n38186), .Z(n38188) );
  NAND U38563 ( .A(n38189), .B(n38188), .Z(n38236) );
  NAND U38564 ( .A(n38191), .B(n38190), .Z(n38195) );
  OR U38565 ( .A(n38193), .B(n38192), .Z(n38194) );
  NAND U38566 ( .A(n38195), .B(n38194), .Z(n38244) );
  NANDN U38567 ( .A(n38200), .B(n38199), .Z(n38204) );
  NAND U38568 ( .A(n38202), .B(n38201), .Z(n38203) );
  NAND U38569 ( .A(n38204), .B(n38203), .Z(n38255) );
  NANDN U38570 ( .A(n38206), .B(n38205), .Z(n38208) );
  XNOR U38571 ( .A(n38595), .B(b[23]), .Z(n38269) );
  NANDN U38572 ( .A(n38268), .B(n38269), .Z(n38207) );
  NAND U38573 ( .A(n38208), .B(n38207), .Z(n38282) );
  XOR U38574 ( .A(b[27]), .B(a[251]), .Z(n38259) );
  NAND U38575 ( .A(n38423), .B(n38259), .Z(n38211) );
  NANDN U38576 ( .A(n38209), .B(n38424), .Z(n38210) );
  AND U38577 ( .A(n38211), .B(n38210), .Z(n38283) );
  XNOR U38578 ( .A(n38282), .B(n38283), .Z(n38284) );
  NANDN U38579 ( .A(n1056), .B(n38212), .Z(n38289) );
  ANDN U38580 ( .B(b[31]), .A(n38213), .Z(n38288) );
  XNOR U38581 ( .A(n38289), .B(n38288), .Z(n38291) );
  XOR U38582 ( .A(n38290), .B(n38291), .Z(n38285) );
  XNOR U38583 ( .A(n38284), .B(n38285), .Z(n38253) );
  XOR U38584 ( .A(a[253]), .B(b[25]), .Z(n38262) );
  NAND U38585 ( .A(n38262), .B(n38325), .Z(n38216) );
  NANDN U38586 ( .A(n38214), .B(n38326), .Z(n38215) );
  NAND U38587 ( .A(n38216), .B(n38215), .Z(n38279) );
  NAND U38588 ( .A(n38217), .B(n38490), .Z(n38219) );
  XNOR U38589 ( .A(n1058), .B(a[249]), .Z(n38265) );
  NANDN U38590 ( .A(n1048), .B(n38265), .Z(n38218) );
  NAND U38591 ( .A(n38219), .B(n38218), .Z(n38276) );
  XNOR U38592 ( .A(n1059), .B(a[247]), .Z(n38273) );
  NAND U38593 ( .A(n38273), .B(n38552), .Z(n38222) );
  NANDN U38594 ( .A(n38220), .B(n38553), .Z(n38221) );
  AND U38595 ( .A(n38222), .B(n38221), .Z(n38277) );
  XNOR U38596 ( .A(n38276), .B(n38277), .Z(n38278) );
  XOR U38597 ( .A(n38279), .B(n38278), .Z(n38254) );
  XNOR U38598 ( .A(n38253), .B(n38254), .Z(n38256) );
  XOR U38599 ( .A(n38255), .B(n38256), .Z(n38248) );
  XOR U38600 ( .A(n38247), .B(n38248), .Z(n38249) );
  XNOR U38601 ( .A(n38249), .B(n38250), .Z(n38242) );
  NANDN U38602 ( .A(n38228), .B(n38227), .Z(n38232) );
  NAND U38603 ( .A(n38230), .B(n38229), .Z(n38231) );
  AND U38604 ( .A(n38232), .B(n38231), .Z(n38241) );
  XNOR U38605 ( .A(n38242), .B(n38241), .Z(n38243) );
  XNOR U38606 ( .A(n38244), .B(n38243), .Z(n38235) );
  XNOR U38607 ( .A(n38236), .B(n38235), .Z(n38238) );
  XNOR U38608 ( .A(n38237), .B(n38238), .Z(n38294) );
  NANDN U38609 ( .A(n38234), .B(n38233), .Z(n38295) );
  XNOR U38610 ( .A(n38294), .B(n38295), .Z(c[501]) );
  NAND U38611 ( .A(n38236), .B(n38235), .Z(n38240) );
  NANDN U38612 ( .A(n38238), .B(n38237), .Z(n38239) );
  NAND U38613 ( .A(n38240), .B(n38239), .Z(n38300) );
  NANDN U38614 ( .A(n38242), .B(n38241), .Z(n38246) );
  NANDN U38615 ( .A(n38244), .B(n38243), .Z(n38245) );
  NAND U38616 ( .A(n38246), .B(n38245), .Z(n38299) );
  OR U38617 ( .A(n38248), .B(n38247), .Z(n38252) );
  NAND U38618 ( .A(n38250), .B(n38249), .Z(n38251) );
  NAND U38619 ( .A(n38252), .B(n38251), .Z(n38307) );
  NAND U38620 ( .A(n38254), .B(n38253), .Z(n38258) );
  NANDN U38621 ( .A(n38256), .B(n38255), .Z(n38257) );
  NAND U38622 ( .A(n38258), .B(n38257), .Z(n38304) );
  XNOR U38623 ( .A(b[27]), .B(a[252]), .Z(n38322) );
  NANDN U38624 ( .A(n38322), .B(n38423), .Z(n38261) );
  NAND U38625 ( .A(n38259), .B(n38424), .Z(n38260) );
  NAND U38626 ( .A(n38261), .B(n38260), .Z(n38311) );
  XNOR U38627 ( .A(a[254]), .B(b[25]), .Z(n38327) );
  NANDN U38628 ( .A(n38327), .B(n38325), .Z(n38264) );
  NAND U38629 ( .A(n38262), .B(n38326), .Z(n38263) );
  NAND U38630 ( .A(n38264), .B(n38263), .Z(n38308) );
  NAND U38631 ( .A(n38490), .B(n38265), .Z(n38267) );
  XOR U38632 ( .A(n1058), .B(n38356), .Z(n38330) );
  NANDN U38633 ( .A(n1048), .B(n38330), .Z(n38266) );
  AND U38634 ( .A(n38267), .B(n38266), .Z(n38309) );
  XNOR U38635 ( .A(n38308), .B(n38309), .Z(n38310) );
  XNOR U38636 ( .A(n38311), .B(n38310), .Z(n38334) );
  NANDN U38637 ( .A(n1056), .B(b[22]), .Z(n38333) );
  XOR U38638 ( .A(n1057), .B(n38333), .Z(n38271) );
  NANDN U38639 ( .A(n38269), .B(n38268), .Z(n38270) );
  AND U38640 ( .A(n38271), .B(n38270), .Z(n38314) );
  AND U38641 ( .A(a[246]), .B(b[31]), .Z(n38368) );
  XNOR U38642 ( .A(n38314), .B(n38368), .Z(n38315) );
  XOR U38643 ( .A(b[31]), .B(n38272), .Z(n38319) );
  NANDN U38644 ( .A(n38319), .B(n38552), .Z(n38275) );
  NAND U38645 ( .A(n38553), .B(n38273), .Z(n38274) );
  AND U38646 ( .A(n38275), .B(n38274), .Z(n38316) );
  XNOR U38647 ( .A(n38315), .B(n38316), .Z(n38335) );
  XOR U38648 ( .A(n38334), .B(n38335), .Z(n38337) );
  NANDN U38649 ( .A(n38277), .B(n38276), .Z(n38281) );
  NAND U38650 ( .A(n38279), .B(n38278), .Z(n38280) );
  NAND U38651 ( .A(n38281), .B(n38280), .Z(n38336) );
  XNOR U38652 ( .A(n38337), .B(n38336), .Z(n38343) );
  NANDN U38653 ( .A(n38283), .B(n38282), .Z(n38287) );
  NANDN U38654 ( .A(n38285), .B(n38284), .Z(n38286) );
  NAND U38655 ( .A(n38287), .B(n38286), .Z(n38340) );
  NAND U38656 ( .A(n38289), .B(n38288), .Z(n38293) );
  NANDN U38657 ( .A(n38291), .B(n38290), .Z(n38292) );
  AND U38658 ( .A(n38293), .B(n38292), .Z(n38341) );
  XNOR U38659 ( .A(n38340), .B(n38341), .Z(n38342) );
  XNOR U38660 ( .A(n38343), .B(n38342), .Z(n38305) );
  XNOR U38661 ( .A(n38304), .B(n38305), .Z(n38306) );
  XOR U38662 ( .A(n38307), .B(n38306), .Z(n38298) );
  XNOR U38663 ( .A(n38299), .B(n38298), .Z(n38301) );
  XNOR U38664 ( .A(n38300), .B(n38301), .Z(n38296) );
  NANDN U38665 ( .A(n38295), .B(n38294), .Z(n38297) );
  XNOR U38666 ( .A(n38296), .B(n38297), .Z(c[502]) );
  NANDN U38667 ( .A(n38297), .B(n38296), .Z(n38393) );
  NAND U38668 ( .A(n38299), .B(n38298), .Z(n38303) );
  NANDN U38669 ( .A(n38301), .B(n38300), .Z(n38302) );
  AND U38670 ( .A(n38303), .B(n38302), .Z(n38349) );
  NANDN U38671 ( .A(n38309), .B(n38308), .Z(n38313) );
  NAND U38672 ( .A(n38311), .B(n38310), .Z(n38312) );
  NAND U38673 ( .A(n38313), .B(n38312), .Z(n38387) );
  NANDN U38674 ( .A(n38314), .B(n38368), .Z(n38318) );
  NAND U38675 ( .A(n38316), .B(n38315), .Z(n38317) );
  NAND U38676 ( .A(n38318), .B(n38317), .Z(n38385) );
  XNOR U38677 ( .A(n1059), .B(a[249]), .Z(n38357) );
  NAND U38678 ( .A(n38357), .B(n38552), .Z(n38321) );
  NANDN U38679 ( .A(n38319), .B(n38553), .Z(n38320) );
  NAND U38680 ( .A(n38321), .B(n38320), .Z(n38380) );
  XOR U38681 ( .A(b[27]), .B(a[253]), .Z(n38375) );
  NAND U38682 ( .A(n38423), .B(n38375), .Z(n38324) );
  NANDN U38683 ( .A(n38322), .B(n38424), .Z(n38323) );
  NAND U38684 ( .A(n38324), .B(n38323), .Z(n38379) );
  XNOR U38685 ( .A(n38595), .B(b[25]), .Z(n38353) );
  NAND U38686 ( .A(n38353), .B(n38325), .Z(n38329) );
  NANDN U38687 ( .A(n38327), .B(n38326), .Z(n38328) );
  NAND U38688 ( .A(n38329), .B(n38328), .Z(n38360) );
  NAND U38689 ( .A(n38490), .B(n38330), .Z(n38332) );
  XNOR U38690 ( .A(n1058), .B(a[251]), .Z(n38372) );
  NANDN U38691 ( .A(n1048), .B(n38372), .Z(n38331) );
  AND U38692 ( .A(n38332), .B(n38331), .Z(n38361) );
  XNOR U38693 ( .A(n38360), .B(n38361), .Z(n38362) );
  ANDN U38694 ( .B(n38333), .A(n1057), .Z(n38367) );
  NANDN U38695 ( .A(n1059), .B(a[247]), .Z(n38366) );
  XOR U38696 ( .A(n38367), .B(n38366), .Z(n38369) );
  XNOR U38697 ( .A(n38368), .B(n38369), .Z(n38363) );
  XNOR U38698 ( .A(n38362), .B(n38363), .Z(n38378) );
  XNOR U38699 ( .A(n38379), .B(n38378), .Z(n38381) );
  XNOR U38700 ( .A(n38380), .B(n38381), .Z(n38384) );
  XNOR U38701 ( .A(n38385), .B(n38384), .Z(n38386) );
  XNOR U38702 ( .A(n38387), .B(n38386), .Z(n38388) );
  NANDN U38703 ( .A(n38335), .B(n38334), .Z(n38339) );
  OR U38704 ( .A(n38337), .B(n38336), .Z(n38338) );
  AND U38705 ( .A(n38339), .B(n38338), .Z(n38389) );
  XNOR U38706 ( .A(n38388), .B(n38389), .Z(n38390) );
  NANDN U38707 ( .A(n38341), .B(n38340), .Z(n38345) );
  NAND U38708 ( .A(n38343), .B(n38342), .Z(n38344) );
  AND U38709 ( .A(n38345), .B(n38344), .Z(n38391) );
  XOR U38710 ( .A(n38390), .B(n38391), .Z(n38348) );
  XOR U38711 ( .A(n38347), .B(n38348), .Z(n38346) );
  XNOR U38712 ( .A(n38349), .B(n38346), .Z(n38392) );
  XOR U38713 ( .A(n38393), .B(n38392), .Z(c[503]) );
  XNOR U38714 ( .A(b[25]), .B(n38350), .Z(n38355) );
  XOR U38715 ( .A(n38351), .B(b[23]), .Z(n38352) );
  NANDN U38716 ( .A(n38353), .B(n38352), .Z(n38354) );
  AND U38717 ( .A(n38355), .B(n38354), .Z(n38418) );
  AND U38718 ( .A(a[248]), .B(b[31]), .Z(n38457) );
  XOR U38719 ( .A(n38418), .B(n38457), .Z(n38420) );
  XOR U38720 ( .A(b[31]), .B(n38356), .Z(n38431) );
  NANDN U38721 ( .A(n38431), .B(n38552), .Z(n38359) );
  NAND U38722 ( .A(n38553), .B(n38357), .Z(n38358) );
  NAND U38723 ( .A(n38359), .B(n38358), .Z(n38419) );
  XNOR U38724 ( .A(n38420), .B(n38419), .Z(n38406) );
  NANDN U38725 ( .A(n38361), .B(n38360), .Z(n38365) );
  NANDN U38726 ( .A(n38363), .B(n38362), .Z(n38364) );
  AND U38727 ( .A(n38365), .B(n38364), .Z(n38407) );
  XNOR U38728 ( .A(n38406), .B(n38407), .Z(n38408) );
  OR U38729 ( .A(n38367), .B(n38366), .Z(n38371) );
  NAND U38730 ( .A(n38369), .B(n38368), .Z(n38370) );
  NAND U38731 ( .A(n38371), .B(n38370), .Z(n38415) );
  NAND U38732 ( .A(n38490), .B(n38372), .Z(n38374) );
  XOR U38733 ( .A(n1058), .B(n38531), .Z(n38428) );
  NANDN U38734 ( .A(n1048), .B(n38428), .Z(n38373) );
  NAND U38735 ( .A(n38374), .B(n38373), .Z(n38412) );
  XNOR U38736 ( .A(b[27]), .B(a[254]), .Z(n38425) );
  NANDN U38737 ( .A(n38425), .B(n38423), .Z(n38377) );
  NAND U38738 ( .A(n38375), .B(n38424), .Z(n38376) );
  AND U38739 ( .A(n38377), .B(n38376), .Z(n38413) );
  XNOR U38740 ( .A(n38412), .B(n38413), .Z(n38414) );
  XNOR U38741 ( .A(n38415), .B(n38414), .Z(n38409) );
  XOR U38742 ( .A(n38408), .B(n38409), .Z(n38400) );
  NAND U38743 ( .A(n38379), .B(n38378), .Z(n38383) );
  NANDN U38744 ( .A(n38381), .B(n38380), .Z(n38382) );
  NAND U38745 ( .A(n38383), .B(n38382), .Z(n38401) );
  XNOR U38746 ( .A(n38400), .B(n38401), .Z(n38402) );
  XOR U38747 ( .A(n38402), .B(n38403), .Z(n38394) );
  XNOR U38748 ( .A(n38394), .B(n38395), .Z(n38397) );
  XOR U38749 ( .A(n38396), .B(n38397), .Z(n38434) );
  OR U38750 ( .A(n38393), .B(n38392), .Z(n38435) );
  XNOR U38751 ( .A(n38434), .B(n38435), .Z(c[504]) );
  NANDN U38752 ( .A(n38395), .B(n38394), .Z(n38399) );
  NAND U38753 ( .A(n38397), .B(n38396), .Z(n38398) );
  NAND U38754 ( .A(n38399), .B(n38398), .Z(n38441) );
  NANDN U38755 ( .A(n38401), .B(n38400), .Z(n38405) );
  NANDN U38756 ( .A(n38403), .B(n38402), .Z(n38404) );
  NAND U38757 ( .A(n38405), .B(n38404), .Z(n38439) );
  NANDN U38758 ( .A(n38407), .B(n38406), .Z(n38411) );
  NANDN U38759 ( .A(n38409), .B(n38408), .Z(n38410) );
  NAND U38760 ( .A(n38411), .B(n38410), .Z(n38473) );
  NANDN U38761 ( .A(n38413), .B(n38412), .Z(n38417) );
  NAND U38762 ( .A(n38415), .B(n38414), .Z(n38416) );
  NAND U38763 ( .A(n38417), .B(n38416), .Z(n38472) );
  NANDN U38764 ( .A(n38418), .B(n38457), .Z(n38422) );
  OR U38765 ( .A(n38420), .B(n38419), .Z(n38421) );
  NAND U38766 ( .A(n38422), .B(n38421), .Z(n38469) );
  XNOR U38767 ( .A(b[27]), .B(n38595), .Z(n38446) );
  NAND U38768 ( .A(n38423), .B(n38446), .Z(n38427) );
  NANDN U38769 ( .A(n38425), .B(n38424), .Z(n38426) );
  NAND U38770 ( .A(n38427), .B(n38426), .Z(n38468) );
  NAND U38771 ( .A(n38490), .B(n38428), .Z(n38430) );
  XNOR U38772 ( .A(n1058), .B(a[253]), .Z(n38452) );
  NANDN U38773 ( .A(n1048), .B(n38452), .Z(n38429) );
  NAND U38774 ( .A(n38430), .B(n38429), .Z(n38461) );
  XNOR U38775 ( .A(n1059), .B(a[251]), .Z(n38449) );
  NAND U38776 ( .A(n38449), .B(n38552), .Z(n38433) );
  NANDN U38777 ( .A(n38431), .B(n38553), .Z(n38432) );
  AND U38778 ( .A(n38433), .B(n38432), .Z(n38462) );
  XNOR U38779 ( .A(n38461), .B(n38462), .Z(n38463) );
  NANDN U38780 ( .A(n1059), .B(a[249]), .Z(n38455) );
  XOR U38781 ( .A(n38456), .B(n38455), .Z(n38458) );
  XNOR U38782 ( .A(n38457), .B(n38458), .Z(n38464) );
  XNOR U38783 ( .A(n38463), .B(n38464), .Z(n38467) );
  XNOR U38784 ( .A(n38468), .B(n38467), .Z(n38470) );
  XOR U38785 ( .A(n38469), .B(n38470), .Z(n38471) );
  XNOR U38786 ( .A(n38472), .B(n38471), .Z(n38474) );
  XNOR U38787 ( .A(n38473), .B(n38474), .Z(n38438) );
  XNOR U38788 ( .A(n38439), .B(n38438), .Z(n38440) );
  XNOR U38789 ( .A(n38441), .B(n38440), .Z(n38437) );
  NANDN U38790 ( .A(n38435), .B(n38434), .Z(n38436) );
  XOR U38791 ( .A(n38437), .B(n38436), .Z(c[505]) );
  OR U38792 ( .A(n38437), .B(n38436), .Z(n38506) );
  NANDN U38793 ( .A(n38439), .B(n38438), .Z(n38443) );
  NAND U38794 ( .A(n38441), .B(n38440), .Z(n38442) );
  AND U38795 ( .A(n38443), .B(n38442), .Z(n38480) );
  XNOR U38796 ( .A(b[27]), .B(n38444), .Z(n38448) );
  XNOR U38797 ( .A(b[26]), .B(b[25]), .Z(n38445) );
  NANDN U38798 ( .A(n38446), .B(n38445), .Z(n38447) );
  AND U38799 ( .A(n38448), .B(n38447), .Z(n38494) );
  AND U38800 ( .A(a[250]), .B(b[31]), .Z(n38523) );
  XOR U38801 ( .A(n38494), .B(n38523), .Z(n38496) );
  XOR U38802 ( .A(b[31]), .B(n38531), .Z(n38487) );
  NANDN U38803 ( .A(n38487), .B(n38552), .Z(n38451) );
  NAND U38804 ( .A(n38553), .B(n38449), .Z(n38450) );
  NAND U38805 ( .A(n38451), .B(n38450), .Z(n38495) );
  XNOR U38806 ( .A(n38496), .B(n38495), .Z(n38484) );
  NAND U38807 ( .A(n38490), .B(n38452), .Z(n38454) );
  XOR U38808 ( .A(b[29]), .B(n38532), .Z(n38491) );
  OR U38809 ( .A(n38491), .B(n1048), .Z(n38453) );
  NAND U38810 ( .A(n38454), .B(n38453), .Z(n38481) );
  OR U38811 ( .A(n38456), .B(n38455), .Z(n38460) );
  NAND U38812 ( .A(n38458), .B(n38457), .Z(n38459) );
  AND U38813 ( .A(n38460), .B(n38459), .Z(n38482) );
  XNOR U38814 ( .A(n38481), .B(n38482), .Z(n38483) );
  XNOR U38815 ( .A(n38484), .B(n38483), .Z(n38499) );
  NANDN U38816 ( .A(n38462), .B(n38461), .Z(n38466) );
  NANDN U38817 ( .A(n38464), .B(n38463), .Z(n38465) );
  NAND U38818 ( .A(n38466), .B(n38465), .Z(n38500) );
  XOR U38819 ( .A(n38499), .B(n38500), .Z(n38502) );
  XOR U38820 ( .A(n38502), .B(n38501), .Z(n38479) );
  NAND U38821 ( .A(n38472), .B(n38471), .Z(n38476) );
  NANDN U38822 ( .A(n38474), .B(n38473), .Z(n38475) );
  AND U38823 ( .A(n38476), .B(n38475), .Z(n38478) );
  XNOR U38824 ( .A(n38479), .B(n38478), .Z(n38477) );
  XOR U38825 ( .A(n38480), .B(n38477), .Z(n38505) );
  XNOR U38826 ( .A(n38506), .B(n38505), .Z(c[506]) );
  NANDN U38827 ( .A(n38482), .B(n38481), .Z(n38486) );
  NAND U38828 ( .A(n38484), .B(n38483), .Z(n38485) );
  NAND U38829 ( .A(n38486), .B(n38485), .Z(n38539) );
  XNOR U38830 ( .A(b[31]), .B(a[253]), .Z(n38533) );
  NANDN U38831 ( .A(n38533), .B(n38552), .Z(n38489) );
  NANDN U38832 ( .A(n38487), .B(n38553), .Z(n38488) );
  NAND U38833 ( .A(n38489), .B(n38488), .Z(n38515) );
  NANDN U38834 ( .A(n38491), .B(n38490), .Z(n38493) );
  XNOR U38835 ( .A(n1058), .B(a[255]), .Z(n38528) );
  NANDN U38836 ( .A(n1048), .B(n38528), .Z(n38492) );
  AND U38837 ( .A(n38493), .B(n38492), .Z(n38516) );
  XNOR U38838 ( .A(n38515), .B(n38516), .Z(n38517) );
  NANDN U38839 ( .A(n1059), .B(a[251]), .Z(n38521) );
  XOR U38840 ( .A(n38522), .B(n38521), .Z(n38524) );
  XNOR U38841 ( .A(n38523), .B(n38524), .Z(n38518) );
  XOR U38842 ( .A(n38517), .B(n38518), .Z(n38536) );
  NANDN U38843 ( .A(n38494), .B(n38523), .Z(n38498) );
  OR U38844 ( .A(n38496), .B(n38495), .Z(n38497) );
  AND U38845 ( .A(n38498), .B(n38497), .Z(n38537) );
  XNOR U38846 ( .A(n38536), .B(n38537), .Z(n38538) );
  XOR U38847 ( .A(n38539), .B(n38538), .Z(n38509) );
  NANDN U38848 ( .A(n38500), .B(n38499), .Z(n38504) );
  OR U38849 ( .A(n38502), .B(n38501), .Z(n38503) );
  NAND U38850 ( .A(n38504), .B(n38503), .Z(n38510) );
  XNOR U38851 ( .A(n38509), .B(n38510), .Z(n38511) );
  XNOR U38852 ( .A(n38512), .B(n38511), .Z(n38507) );
  NANDN U38853 ( .A(n38506), .B(n38505), .Z(n38508) );
  XNOR U38854 ( .A(n38507), .B(n38508), .Z(c[507]) );
  NANDN U38855 ( .A(n38508), .B(n38507), .Z(n38564) );
  NANDN U38856 ( .A(n38510), .B(n38509), .Z(n38514) );
  NANDN U38857 ( .A(n38512), .B(n38511), .Z(n38513) );
  AND U38858 ( .A(n38514), .B(n38513), .Z(n38545) );
  NANDN U38859 ( .A(n38516), .B(n38515), .Z(n38520) );
  NANDN U38860 ( .A(n38518), .B(n38517), .Z(n38519) );
  NAND U38861 ( .A(n38520), .B(n38519), .Z(n38548) );
  OR U38862 ( .A(n38522), .B(n38521), .Z(n38526) );
  NAND U38863 ( .A(n38524), .B(n38523), .Z(n38525) );
  NAND U38864 ( .A(n38526), .B(n38525), .Z(n38547) );
  XOR U38865 ( .A(n1058), .B(n38527), .Z(n38530) );
  NANDN U38866 ( .A(n38528), .B(n1048), .Z(n38529) );
  NAND U38867 ( .A(n38530), .B(n38529), .Z(n38560) );
  ANDN U38868 ( .B(b[31]), .A(n38531), .Z(n38557) );
  IV U38869 ( .A(n38557), .Z(n38569) );
  XOR U38870 ( .A(b[31]), .B(n38532), .Z(n38554) );
  NANDN U38871 ( .A(n38554), .B(n38552), .Z(n38535) );
  NANDN U38872 ( .A(n38533), .B(n38553), .Z(n38534) );
  AND U38873 ( .A(n38535), .B(n38534), .Z(n38558) );
  XNOR U38874 ( .A(n38569), .B(n38558), .Z(n38559) );
  XNOR U38875 ( .A(n38547), .B(n38546), .Z(n38549) );
  XOR U38876 ( .A(n38548), .B(n38549), .Z(n38543) );
  NANDN U38877 ( .A(n38537), .B(n38536), .Z(n38541) );
  NANDN U38878 ( .A(n38539), .B(n38538), .Z(n38540) );
  AND U38879 ( .A(n38541), .B(n38540), .Z(n38544) );
  XOR U38880 ( .A(n38543), .B(n38544), .Z(n38542) );
  XOR U38881 ( .A(n38545), .B(n38542), .Z(n38563) );
  XNOR U38882 ( .A(n38564), .B(n38563), .Z(c[508]) );
  NAND U38883 ( .A(n38547), .B(n38546), .Z(n38551) );
  NANDN U38884 ( .A(n38549), .B(n38548), .Z(n38550) );
  NAND U38885 ( .A(n38551), .B(n38550), .Z(n38578) );
  XOR U38886 ( .A(b[31]), .B(n38595), .Z(n38573) );
  NANDN U38887 ( .A(n38573), .B(n38552), .Z(n38556) );
  NANDN U38888 ( .A(n38554), .B(n38553), .Z(n38555) );
  AND U38889 ( .A(n38556), .B(n38555), .Z(n38584) );
  OR U38890 ( .A(n38558), .B(n38557), .Z(n38562) );
  NANDN U38891 ( .A(n38560), .B(n38559), .Z(n38561) );
  AND U38892 ( .A(n38562), .B(n38561), .Z(n38585) );
  XOR U38893 ( .A(n38584), .B(n38585), .Z(n38586) );
  NANDN U38894 ( .A(n1059), .B(a[253]), .Z(n38568) );
  XNOR U38895 ( .A(n38567), .B(n38568), .Z(n38570) );
  XNOR U38896 ( .A(n38569), .B(n38570), .Z(n38587) );
  XOR U38897 ( .A(n38586), .B(n38587), .Z(n38579) );
  XNOR U38898 ( .A(n38578), .B(n38579), .Z(n38580) );
  XNOR U38899 ( .A(n38581), .B(n38580), .Z(n38565) );
  NANDN U38900 ( .A(n38564), .B(n38563), .Z(n38566) );
  XNOR U38901 ( .A(n38565), .B(n38566), .Z(c[509]) );
  NANDN U38902 ( .A(n38566), .B(n38565), .Z(n38604) );
  AND U38903 ( .A(a[254]), .B(b[31]), .Z(n38591) );
  OR U38904 ( .A(n38568), .B(n38567), .Z(n38572) );
  OR U38905 ( .A(n38570), .B(n38569), .Z(n38571) );
  NAND U38906 ( .A(n38572), .B(n38571), .Z(n38590) );
  ANDN U38907 ( .B(b[30]), .A(n1058), .Z(n38594) );
  XOR U38908 ( .A(b[31]), .B(n38594), .Z(n38576) );
  NAND U38909 ( .A(n38574), .B(n38573), .Z(n38575) );
  AND U38910 ( .A(n38576), .B(n38575), .Z(n38577) );
  XNOR U38911 ( .A(n38590), .B(n38577), .Z(n38592) );
  XNOR U38912 ( .A(n38591), .B(n38592), .Z(n38600) );
  NANDN U38913 ( .A(n38579), .B(n38578), .Z(n38583) );
  NANDN U38914 ( .A(n38581), .B(n38580), .Z(n38582) );
  NAND U38915 ( .A(n38583), .B(n38582), .Z(n38598) );
  OR U38916 ( .A(n38585), .B(n38584), .Z(n38589) );
  NANDN U38917 ( .A(n38587), .B(n38586), .Z(n38588) );
  NAND U38918 ( .A(n38589), .B(n38588), .Z(n38597) );
  XOR U38919 ( .A(n38598), .B(n38597), .Z(n38599) );
  XOR U38920 ( .A(n38600), .B(n38599), .Z(n38603) );
  XOR U38921 ( .A(n38604), .B(n38603), .Z(c[510]) );
  XNOR U38922 ( .A(n38591), .B(n38590), .Z(n38593) );
  NAND U38923 ( .A(n38593), .B(n38592), .Z(n38610) );
  XOR U38924 ( .A(n38595), .B(n38594), .Z(n38596) );
  ANDN U38925 ( .B(n38596), .A(n1059), .Z(n38608) );
  NOR U38926 ( .A(n38598), .B(n38597), .Z(n38602) );
  AND U38927 ( .A(n38600), .B(n38599), .Z(n38601) );
  OR U38928 ( .A(n38602), .B(n38601), .Z(n38606) );
  OR U38929 ( .A(n38604), .B(n38603), .Z(n38605) );
  NAND U38930 ( .A(n38606), .B(n38605), .Z(n38607) );
  XNOR U38931 ( .A(n38608), .B(n38607), .Z(n38609) );
  XOR U38932 ( .A(n38610), .B(n38609), .Z(c[511]) );
endmodule

