
module mult_N128_CC128 ( clk, rst, a, b, c );
  input [127:0] a;
  input [0:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614;
  wire   [127:1] swire;
  wire   [255:128] sreg;

  DFF \sreg_reg[128]  ( .D(swire[1]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[129]  ( .D(swire[2]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[130]  ( .D(swire[3]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[131]  ( .D(swire[4]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[132]  ( .D(swire[5]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[133]  ( .D(swire[6]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[134]  ( .D(swire[7]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[135]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[136]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[137]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[138]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[139]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[140]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[141]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[142]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[143]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[144]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[145]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[146]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[147]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[148]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[149]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[150]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[151]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[152]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[153]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[154]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[155]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[156]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[157]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[158]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[159]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[160]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[161]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[162]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[163]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[164]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[165]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[166]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[167]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[168]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[169]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[170]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[171]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[172]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[173]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[174]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[175]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[176]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[177]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[178]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[179]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[180]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[181]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[182]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[183]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[184]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[185]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[186]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[187]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[188]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[189]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[190]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[191]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[192]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[193]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[194]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[195]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[196]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[197]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[198]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[199]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[200]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[201]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[202]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[203]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[204]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[205]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[206]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[207]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[208]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[209]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[210]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[211]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[212]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[213]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[214]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[215]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[216]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[217]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[218]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[219]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[220]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[221]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[222]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[223]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[224]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[225]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[226]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[227]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[228]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[229]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[230]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[231]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[232]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[233]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[234]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[235]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[236]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[237]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[238]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[239]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[240]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[241]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[242]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[243]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[244]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[245]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[246]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[247]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[248]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[249]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[250]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[251]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[252]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[253]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[254]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[3]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[2]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[1]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U4 ( .A(n224), .B(n221), .Z(n222) );
  XNOR U5 ( .A(n239), .B(n236), .Z(n237) );
  XNOR U6 ( .A(n254), .B(n251), .Z(n252) );
  XNOR U7 ( .A(n271), .B(n266), .Z(n267) );
  XNOR U8 ( .A(n286), .B(n283), .Z(n284) );
  XNOR U9 ( .A(n301), .B(n298), .Z(n299) );
  XNOR U10 ( .A(n316), .B(n313), .Z(n314) );
  XNOR U11 ( .A(n325), .B(n324), .Z(n7) );
  XNOR U12 ( .A(n334), .B(n333), .Z(n13) );
  XNOR U13 ( .A(n343), .B(n342), .Z(n19) );
  XNOR U14 ( .A(n352), .B(n351), .Z(n27) );
  XNOR U15 ( .A(n361), .B(n360), .Z(n33) );
  XNOR U16 ( .A(n370), .B(n369), .Z(n39) );
  XNOR U17 ( .A(n379), .B(n378), .Z(n47) );
  XNOR U18 ( .A(n388), .B(n387), .Z(n53) );
  XNOR U19 ( .A(n397), .B(n396), .Z(n59) );
  XNOR U20 ( .A(n406), .B(n405), .Z(n65) );
  XNOR U21 ( .A(n415), .B(n414), .Z(n73) );
  XNOR U22 ( .A(n424), .B(n423), .Z(n79) );
  XNOR U23 ( .A(n433), .B(n432), .Z(n85) );
  XNOR U24 ( .A(n442), .B(n441), .Z(n93) );
  XNOR U25 ( .A(n451), .B(n450), .Z(n99) );
  XNOR U26 ( .A(n460), .B(n459), .Z(n105) );
  XNOR U27 ( .A(n469), .B(n468), .Z(n113) );
  XNOR U28 ( .A(n478), .B(n477), .Z(n119) );
  XNOR U29 ( .A(n487), .B(n486), .Z(n125) );
  XNOR U30 ( .A(n496), .B(n495), .Z(n131) );
  XNOR U31 ( .A(n505), .B(n504), .Z(n139) );
  XNOR U32 ( .A(n514), .B(n513), .Z(n145) );
  XNOR U33 ( .A(n523), .B(n522), .Z(n151) );
  XNOR U34 ( .A(n532), .B(n531), .Z(n159) );
  XNOR U35 ( .A(n541), .B(n540), .Z(n165) );
  XNOR U36 ( .A(n550), .B(n549), .Z(n171) );
  XNOR U37 ( .A(n559), .B(n558), .Z(n179) );
  XNOR U38 ( .A(n568), .B(n567), .Z(n185) );
  XNOR U39 ( .A(n577), .B(n576), .Z(n191) );
  XNOR U40 ( .A(n586), .B(n585), .Z(n269) );
  XNOR U41 ( .A(n595), .B(n594), .Z(n45) );
  XNOR U42 ( .A(n604), .B(n603), .Z(n111) );
  XNOR U43 ( .A(n212), .B(n209), .Z(n210) );
  XNOR U44 ( .A(n229), .B(n226), .Z(n227) );
  XNOR U45 ( .A(n244), .B(n241), .Z(n242) );
  XNOR U46 ( .A(n259), .B(n256), .Z(n257) );
  XNOR U47 ( .A(n276), .B(n273), .Z(n274) );
  XNOR U48 ( .A(n291), .B(n288), .Z(n289) );
  XNOR U49 ( .A(n306), .B(n303), .Z(n304) );
  XNOR U50 ( .A(n319), .B(n318), .Z(n4) );
  XNOR U51 ( .A(n328), .B(n327), .Z(n9) );
  XNOR U52 ( .A(n337), .B(n336), .Z(n15) );
  XNOR U53 ( .A(n346), .B(n345), .Z(n21) );
  XNOR U54 ( .A(n355), .B(n354), .Z(n29) );
  XNOR U55 ( .A(n364), .B(n363), .Z(n35) );
  XNOR U56 ( .A(n373), .B(n372), .Z(n41) );
  XNOR U57 ( .A(n382), .B(n381), .Z(n49) );
  XNOR U58 ( .A(n391), .B(n390), .Z(n55) );
  XNOR U59 ( .A(n400), .B(n399), .Z(n61) );
  XNOR U60 ( .A(n409), .B(n408), .Z(n69) );
  XNOR U61 ( .A(n418), .B(n417), .Z(n75) );
  XNOR U62 ( .A(n427), .B(n426), .Z(n81) );
  XNOR U63 ( .A(n436), .B(n435), .Z(n87) );
  XNOR U64 ( .A(n445), .B(n444), .Z(n95) );
  XNOR U65 ( .A(n454), .B(n453), .Z(n101) );
  XNOR U66 ( .A(n463), .B(n462), .Z(n107) );
  XNOR U67 ( .A(n472), .B(n471), .Z(n115) );
  XNOR U68 ( .A(n481), .B(n480), .Z(n121) );
  XNOR U69 ( .A(n490), .B(n489), .Z(n127) );
  XNOR U70 ( .A(n499), .B(n498), .Z(n135) );
  XNOR U71 ( .A(n508), .B(n507), .Z(n141) );
  XNOR U72 ( .A(n517), .B(n516), .Z(n147) );
  XNOR U73 ( .A(n526), .B(n525), .Z(n153) );
  XNOR U74 ( .A(n535), .B(n534), .Z(n161) );
  XNOR U75 ( .A(n544), .B(n543), .Z(n167) );
  XNOR U76 ( .A(n553), .B(n552), .Z(n173) );
  XNOR U77 ( .A(n562), .B(n561), .Z(n181) );
  XNOR U78 ( .A(n571), .B(n570), .Z(n187) );
  XNOR U79 ( .A(n580), .B(n579), .Z(n193) );
  XNOR U80 ( .A(n589), .B(n588), .Z(n2) );
  XNOR U81 ( .A(n598), .B(n597), .Z(n67) );
  XNOR U82 ( .A(n607), .B(n606), .Z(n133) );
  XNOR U83 ( .A(n219), .B(n214), .Z(n215) );
  XNOR U84 ( .A(n234), .B(n231), .Z(n232) );
  XNOR U85 ( .A(n249), .B(n246), .Z(n247) );
  XNOR U86 ( .A(n264), .B(n261), .Z(n262) );
  XNOR U87 ( .A(n281), .B(n278), .Z(n279) );
  XNOR U88 ( .A(n296), .B(n293), .Z(n294) );
  XNOR U89 ( .A(n311), .B(n308), .Z(n309) );
  XNOR U90 ( .A(n322), .B(n321), .Z(n5) );
  XNOR U91 ( .A(n331), .B(n330), .Z(n11) );
  XNOR U92 ( .A(n340), .B(n339), .Z(n17) );
  XNOR U93 ( .A(n349), .B(n348), .Z(n25) );
  XNOR U94 ( .A(n358), .B(n357), .Z(n31) );
  XNOR U95 ( .A(n367), .B(n366), .Z(n37) );
  XNOR U96 ( .A(n376), .B(n375), .Z(n43) );
  XNOR U97 ( .A(n385), .B(n384), .Z(n51) );
  XNOR U98 ( .A(n394), .B(n393), .Z(n57) );
  XNOR U99 ( .A(n403), .B(n402), .Z(n63) );
  XNOR U100 ( .A(n412), .B(n411), .Z(n71) );
  XNOR U101 ( .A(n421), .B(n420), .Z(n77) );
  XNOR U102 ( .A(n430), .B(n429), .Z(n83) );
  XNOR U103 ( .A(n439), .B(n438), .Z(n91) );
  XNOR U104 ( .A(n448), .B(n447), .Z(n97) );
  XNOR U105 ( .A(n457), .B(n456), .Z(n103) );
  XNOR U106 ( .A(n466), .B(n465), .Z(n109) );
  XNOR U107 ( .A(n475), .B(n474), .Z(n117) );
  XNOR U108 ( .A(n484), .B(n483), .Z(n123) );
  XNOR U109 ( .A(n493), .B(n492), .Z(n129) );
  XNOR U110 ( .A(n502), .B(n501), .Z(n137) );
  XNOR U111 ( .A(n511), .B(n510), .Z(n143) );
  XNOR U112 ( .A(n520), .B(n519), .Z(n149) );
  XNOR U113 ( .A(n529), .B(n528), .Z(n157) );
  XNOR U114 ( .A(n538), .B(n537), .Z(n163) );
  XNOR U115 ( .A(n547), .B(n546), .Z(n169) );
  XNOR U116 ( .A(n556), .B(n555), .Z(n175) );
  XNOR U117 ( .A(n565), .B(n564), .Z(n183) );
  XNOR U118 ( .A(n574), .B(n573), .Z(n189) );
  XNOR U119 ( .A(n583), .B(n582), .Z(n217) );
  XNOR U120 ( .A(n592), .B(n591), .Z(n23) );
  XNOR U121 ( .A(n601), .B(n600), .Z(n89) );
  XOR U122 ( .A(n610), .B(n609), .Z(n155) );
  XNOR U123 ( .A(n1), .B(n2), .Z(swire[9]) );
  XNOR U124 ( .A(n3), .B(n4), .Z(swire[99]) );
  XNOR U125 ( .A(n5), .B(n6), .Z(swire[98]) );
  XNOR U126 ( .A(n7), .B(n8), .Z(swire[97]) );
  XNOR U127 ( .A(n9), .B(n10), .Z(swire[96]) );
  XNOR U128 ( .A(n11), .B(n12), .Z(swire[95]) );
  XNOR U129 ( .A(n13), .B(n14), .Z(swire[94]) );
  XNOR U130 ( .A(n15), .B(n16), .Z(swire[93]) );
  XNOR U131 ( .A(n17), .B(n18), .Z(swire[92]) );
  XNOR U132 ( .A(n19), .B(n20), .Z(swire[91]) );
  XNOR U133 ( .A(n21), .B(n22), .Z(swire[90]) );
  XNOR U134 ( .A(n23), .B(n24), .Z(swire[8]) );
  XNOR U135 ( .A(n25), .B(n26), .Z(swire[89]) );
  XNOR U136 ( .A(n27), .B(n28), .Z(swire[88]) );
  XNOR U137 ( .A(n29), .B(n30), .Z(swire[87]) );
  XNOR U138 ( .A(n31), .B(n32), .Z(swire[86]) );
  XNOR U139 ( .A(n33), .B(n34), .Z(swire[85]) );
  XNOR U140 ( .A(n35), .B(n36), .Z(swire[84]) );
  XNOR U141 ( .A(n37), .B(n38), .Z(swire[83]) );
  XNOR U142 ( .A(n39), .B(n40), .Z(swire[82]) );
  XNOR U143 ( .A(n41), .B(n42), .Z(swire[81]) );
  XNOR U144 ( .A(n43), .B(n44), .Z(swire[80]) );
  XNOR U145 ( .A(n45), .B(n46), .Z(swire[7]) );
  XNOR U146 ( .A(n47), .B(n48), .Z(swire[79]) );
  XNOR U147 ( .A(n49), .B(n50), .Z(swire[78]) );
  XNOR U148 ( .A(n51), .B(n52), .Z(swire[77]) );
  XNOR U149 ( .A(n53), .B(n54), .Z(swire[76]) );
  XNOR U150 ( .A(n55), .B(n56), .Z(swire[75]) );
  XNOR U151 ( .A(n57), .B(n58), .Z(swire[74]) );
  XNOR U152 ( .A(n59), .B(n60), .Z(swire[73]) );
  XNOR U153 ( .A(n61), .B(n62), .Z(swire[72]) );
  XNOR U154 ( .A(n63), .B(n64), .Z(swire[71]) );
  XNOR U155 ( .A(n65), .B(n66), .Z(swire[70]) );
  XNOR U156 ( .A(n67), .B(n68), .Z(swire[6]) );
  XNOR U157 ( .A(n69), .B(n70), .Z(swire[69]) );
  XNOR U158 ( .A(n71), .B(n72), .Z(swire[68]) );
  XNOR U159 ( .A(n73), .B(n74), .Z(swire[67]) );
  XNOR U160 ( .A(n75), .B(n76), .Z(swire[66]) );
  XNOR U161 ( .A(n77), .B(n78), .Z(swire[65]) );
  XNOR U162 ( .A(n79), .B(n80), .Z(swire[64]) );
  XNOR U163 ( .A(n81), .B(n82), .Z(swire[63]) );
  XNOR U164 ( .A(n83), .B(n84), .Z(swire[62]) );
  XNOR U165 ( .A(n85), .B(n86), .Z(swire[61]) );
  XNOR U166 ( .A(n87), .B(n88), .Z(swire[60]) );
  XNOR U167 ( .A(n89), .B(n90), .Z(swire[5]) );
  XNOR U168 ( .A(n91), .B(n92), .Z(swire[59]) );
  XNOR U169 ( .A(n93), .B(n94), .Z(swire[58]) );
  XNOR U170 ( .A(n95), .B(n96), .Z(swire[57]) );
  XNOR U171 ( .A(n97), .B(n98), .Z(swire[56]) );
  XNOR U172 ( .A(n99), .B(n100), .Z(swire[55]) );
  XNOR U173 ( .A(n101), .B(n102), .Z(swire[54]) );
  XNOR U174 ( .A(n103), .B(n104), .Z(swire[53]) );
  XNOR U175 ( .A(n105), .B(n106), .Z(swire[52]) );
  XNOR U176 ( .A(n107), .B(n108), .Z(swire[51]) );
  XNOR U177 ( .A(n109), .B(n110), .Z(swire[50]) );
  XNOR U178 ( .A(n111), .B(n112), .Z(swire[4]) );
  XNOR U179 ( .A(n113), .B(n114), .Z(swire[49]) );
  XNOR U180 ( .A(n115), .B(n116), .Z(swire[48]) );
  XNOR U181 ( .A(n117), .B(n118), .Z(swire[47]) );
  XNOR U182 ( .A(n119), .B(n120), .Z(swire[46]) );
  XNOR U183 ( .A(n121), .B(n122), .Z(swire[45]) );
  XNOR U184 ( .A(n123), .B(n124), .Z(swire[44]) );
  XNOR U185 ( .A(n125), .B(n126), .Z(swire[43]) );
  XNOR U186 ( .A(n127), .B(n128), .Z(swire[42]) );
  XNOR U187 ( .A(n129), .B(n130), .Z(swire[41]) );
  XNOR U188 ( .A(n131), .B(n132), .Z(swire[40]) );
  XNOR U189 ( .A(n133), .B(n134), .Z(swire[3]) );
  XNOR U190 ( .A(n135), .B(n136), .Z(swire[39]) );
  XNOR U191 ( .A(n137), .B(n138), .Z(swire[38]) );
  XNOR U192 ( .A(n139), .B(n140), .Z(swire[37]) );
  XNOR U193 ( .A(n141), .B(n142), .Z(swire[36]) );
  XNOR U194 ( .A(n143), .B(n144), .Z(swire[35]) );
  XNOR U195 ( .A(n145), .B(n146), .Z(swire[34]) );
  XNOR U196 ( .A(n147), .B(n148), .Z(swire[33]) );
  XNOR U197 ( .A(n149), .B(n150), .Z(swire[32]) );
  XNOR U198 ( .A(n151), .B(n152), .Z(swire[31]) );
  XNOR U199 ( .A(n153), .B(n154), .Z(swire[30]) );
  XOR U200 ( .A(n155), .B(n156), .Z(swire[2]) );
  XNOR U201 ( .A(n157), .B(n158), .Z(swire[29]) );
  XNOR U202 ( .A(n159), .B(n160), .Z(swire[28]) );
  XNOR U203 ( .A(n161), .B(n162), .Z(swire[27]) );
  XNOR U204 ( .A(n163), .B(n164), .Z(swire[26]) );
  XNOR U205 ( .A(n165), .B(n166), .Z(swire[25]) );
  XNOR U206 ( .A(n167), .B(n168), .Z(swire[24]) );
  XNOR U207 ( .A(n169), .B(n170), .Z(swire[23]) );
  XNOR U208 ( .A(n171), .B(n172), .Z(swire[22]) );
  XNOR U209 ( .A(n173), .B(n174), .Z(swire[21]) );
  XNOR U210 ( .A(n175), .B(n176), .Z(swire[20]) );
  XOR U211 ( .A(n177), .B(n178), .Z(swire[1]) );
  XNOR U212 ( .A(n179), .B(n180), .Z(swire[19]) );
  XNOR U213 ( .A(n181), .B(n182), .Z(swire[18]) );
  XNOR U214 ( .A(n183), .B(n184), .Z(swire[17]) );
  XNOR U215 ( .A(n185), .B(n186), .Z(swire[16]) );
  XNOR U216 ( .A(n187), .B(n188), .Z(swire[15]) );
  XNOR U217 ( .A(n189), .B(n190), .Z(swire[14]) );
  XNOR U218 ( .A(n191), .B(n192), .Z(swire[13]) );
  XNOR U219 ( .A(n193), .B(n194), .Z(swire[12]) );
  AND U220 ( .A(a[127]), .B(b[0]), .Z(swire[127]) );
  XOR U221 ( .A(sreg[254]), .B(n195), .Z(swire[126]) );
  AND U222 ( .A(a[126]), .B(b[0]), .Z(n195) );
  XOR U223 ( .A(sreg[253]), .B(n196), .Z(swire[125]) );
  AND U224 ( .A(a[125]), .B(b[0]), .Z(n196) );
  XOR U225 ( .A(sreg[252]), .B(n197), .Z(swire[124]) );
  AND U226 ( .A(a[124]), .B(b[0]), .Z(n197) );
  XOR U227 ( .A(sreg[251]), .B(n198), .Z(swire[123]) );
  AND U228 ( .A(a[123]), .B(b[0]), .Z(n198) );
  XOR U229 ( .A(n199), .B(n200), .Z(swire[122]) );
  XNOR U230 ( .A(sreg[250]), .B(n201), .Z(n200) );
  XNOR U231 ( .A(n202), .B(n201), .Z(n199) );
  XNOR U232 ( .A(n203), .B(n204), .Z(n201) );
  ANDN U233 ( .B(n205), .A(n206), .Z(n203) );
  AND U234 ( .A(a[122]), .B(b[0]), .Z(n202) );
  XNOR U235 ( .A(n205), .B(n206), .Z(swire[121]) );
  XNOR U236 ( .A(sreg[249]), .B(n204), .Z(n206) );
  XOR U237 ( .A(n207), .B(n204), .Z(n205) );
  XNOR U238 ( .A(n208), .B(n209), .Z(n204) );
  ANDN U239 ( .B(n210), .A(n211), .Z(n208) );
  AND U240 ( .A(a[121]), .B(b[0]), .Z(n207) );
  XNOR U241 ( .A(n210), .B(n211), .Z(swire[120]) );
  XOR U242 ( .A(sreg[248]), .B(n209), .Z(n211) );
  XOR U243 ( .A(n213), .B(n214), .Z(n209) );
  ANDN U244 ( .B(n215), .A(n216), .Z(n213) );
  AND U245 ( .A(a[120]), .B(b[0]), .Z(n212) );
  XNOR U246 ( .A(n217), .B(n218), .Z(swire[11]) );
  XNOR U247 ( .A(n215), .B(n216), .Z(swire[119]) );
  XOR U248 ( .A(sreg[247]), .B(n214), .Z(n216) );
  XOR U249 ( .A(n220), .B(n221), .Z(n214) );
  ANDN U250 ( .B(n222), .A(n223), .Z(n220) );
  AND U251 ( .A(a[119]), .B(b[0]), .Z(n219) );
  XNOR U252 ( .A(n222), .B(n223), .Z(swire[118]) );
  XOR U253 ( .A(sreg[246]), .B(n221), .Z(n223) );
  XOR U254 ( .A(n225), .B(n226), .Z(n221) );
  ANDN U255 ( .B(n227), .A(n228), .Z(n225) );
  AND U256 ( .A(a[118]), .B(b[0]), .Z(n224) );
  XNOR U257 ( .A(n227), .B(n228), .Z(swire[117]) );
  XOR U258 ( .A(sreg[245]), .B(n226), .Z(n228) );
  XOR U259 ( .A(n230), .B(n231), .Z(n226) );
  ANDN U260 ( .B(n232), .A(n233), .Z(n230) );
  AND U261 ( .A(a[117]), .B(b[0]), .Z(n229) );
  XNOR U262 ( .A(n232), .B(n233), .Z(swire[116]) );
  XOR U263 ( .A(sreg[244]), .B(n231), .Z(n233) );
  XOR U264 ( .A(n235), .B(n236), .Z(n231) );
  ANDN U265 ( .B(n237), .A(n238), .Z(n235) );
  AND U266 ( .A(a[116]), .B(b[0]), .Z(n234) );
  XNOR U267 ( .A(n237), .B(n238), .Z(swire[115]) );
  XOR U268 ( .A(sreg[243]), .B(n236), .Z(n238) );
  XOR U269 ( .A(n240), .B(n241), .Z(n236) );
  ANDN U270 ( .B(n242), .A(n243), .Z(n240) );
  AND U271 ( .A(a[115]), .B(b[0]), .Z(n239) );
  XNOR U272 ( .A(n242), .B(n243), .Z(swire[114]) );
  XOR U273 ( .A(sreg[242]), .B(n241), .Z(n243) );
  XOR U274 ( .A(n245), .B(n246), .Z(n241) );
  ANDN U275 ( .B(n247), .A(n248), .Z(n245) );
  AND U276 ( .A(a[114]), .B(b[0]), .Z(n244) );
  XNOR U277 ( .A(n247), .B(n248), .Z(swire[113]) );
  XOR U278 ( .A(sreg[241]), .B(n246), .Z(n248) );
  XOR U279 ( .A(n250), .B(n251), .Z(n246) );
  ANDN U280 ( .B(n252), .A(n253), .Z(n250) );
  AND U281 ( .A(a[113]), .B(b[0]), .Z(n249) );
  XNOR U282 ( .A(n252), .B(n253), .Z(swire[112]) );
  XOR U283 ( .A(sreg[240]), .B(n251), .Z(n253) );
  XOR U284 ( .A(n255), .B(n256), .Z(n251) );
  ANDN U285 ( .B(n257), .A(n258), .Z(n255) );
  AND U286 ( .A(a[112]), .B(b[0]), .Z(n254) );
  XNOR U287 ( .A(n257), .B(n258), .Z(swire[111]) );
  XOR U288 ( .A(sreg[239]), .B(n256), .Z(n258) );
  XOR U289 ( .A(n260), .B(n261), .Z(n256) );
  ANDN U290 ( .B(n262), .A(n263), .Z(n260) );
  AND U291 ( .A(a[111]), .B(b[0]), .Z(n259) );
  XNOR U292 ( .A(n262), .B(n263), .Z(swire[110]) );
  XOR U293 ( .A(sreg[238]), .B(n261), .Z(n263) );
  XOR U294 ( .A(n265), .B(n266), .Z(n261) );
  ANDN U295 ( .B(n267), .A(n268), .Z(n265) );
  AND U296 ( .A(a[110]), .B(b[0]), .Z(n264) );
  XNOR U297 ( .A(n269), .B(n270), .Z(swire[10]) );
  XNOR U298 ( .A(n267), .B(n268), .Z(swire[109]) );
  XOR U299 ( .A(sreg[237]), .B(n266), .Z(n268) );
  XOR U300 ( .A(n272), .B(n273), .Z(n266) );
  ANDN U301 ( .B(n274), .A(n275), .Z(n272) );
  AND U302 ( .A(a[109]), .B(b[0]), .Z(n271) );
  XNOR U303 ( .A(n274), .B(n275), .Z(swire[108]) );
  XOR U304 ( .A(sreg[236]), .B(n273), .Z(n275) );
  XOR U305 ( .A(n277), .B(n278), .Z(n273) );
  ANDN U306 ( .B(n279), .A(n280), .Z(n277) );
  AND U307 ( .A(a[108]), .B(b[0]), .Z(n276) );
  XNOR U308 ( .A(n279), .B(n280), .Z(swire[107]) );
  XOR U309 ( .A(sreg[235]), .B(n278), .Z(n280) );
  XOR U310 ( .A(n282), .B(n283), .Z(n278) );
  ANDN U311 ( .B(n284), .A(n285), .Z(n282) );
  AND U312 ( .A(a[107]), .B(b[0]), .Z(n281) );
  XNOR U313 ( .A(n284), .B(n285), .Z(swire[106]) );
  XOR U314 ( .A(sreg[234]), .B(n283), .Z(n285) );
  XOR U315 ( .A(n287), .B(n288), .Z(n283) );
  ANDN U316 ( .B(n289), .A(n290), .Z(n287) );
  AND U317 ( .A(a[106]), .B(b[0]), .Z(n286) );
  XNOR U318 ( .A(n289), .B(n290), .Z(swire[105]) );
  XOR U319 ( .A(sreg[233]), .B(n288), .Z(n290) );
  XOR U320 ( .A(n292), .B(n293), .Z(n288) );
  ANDN U321 ( .B(n294), .A(n295), .Z(n292) );
  AND U322 ( .A(a[105]), .B(b[0]), .Z(n291) );
  XNOR U323 ( .A(n294), .B(n295), .Z(swire[104]) );
  XOR U324 ( .A(sreg[232]), .B(n293), .Z(n295) );
  XOR U325 ( .A(n297), .B(n298), .Z(n293) );
  ANDN U326 ( .B(n299), .A(n300), .Z(n297) );
  AND U327 ( .A(a[104]), .B(b[0]), .Z(n296) );
  XNOR U328 ( .A(n299), .B(n300), .Z(swire[103]) );
  XOR U329 ( .A(sreg[231]), .B(n298), .Z(n300) );
  XOR U330 ( .A(n302), .B(n303), .Z(n298) );
  ANDN U331 ( .B(n304), .A(n305), .Z(n302) );
  AND U332 ( .A(a[103]), .B(b[0]), .Z(n301) );
  XNOR U333 ( .A(n304), .B(n305), .Z(swire[102]) );
  XOR U334 ( .A(sreg[230]), .B(n303), .Z(n305) );
  XOR U335 ( .A(n307), .B(n308), .Z(n303) );
  ANDN U336 ( .B(n309), .A(n310), .Z(n307) );
  AND U337 ( .A(a[102]), .B(b[0]), .Z(n306) );
  XNOR U338 ( .A(n309), .B(n310), .Z(swire[101]) );
  XOR U339 ( .A(sreg[229]), .B(n308), .Z(n310) );
  XOR U340 ( .A(n312), .B(n313), .Z(n308) );
  ANDN U341 ( .B(n314), .A(n315), .Z(n312) );
  AND U342 ( .A(a[101]), .B(b[0]), .Z(n311) );
  XNOR U343 ( .A(n314), .B(n315), .Z(swire[100]) );
  XOR U344 ( .A(sreg[228]), .B(n313), .Z(n315) );
  XOR U345 ( .A(n317), .B(n318), .Z(n313) );
  ANDN U346 ( .B(n4), .A(n3), .Z(n317) );
  XOR U347 ( .A(sreg[227]), .B(n318), .Z(n3) );
  XOR U348 ( .A(n320), .B(n321), .Z(n318) );
  ANDN U349 ( .B(n5), .A(n6), .Z(n320) );
  XOR U350 ( .A(sreg[226]), .B(n321), .Z(n6) );
  XOR U351 ( .A(n323), .B(n324), .Z(n321) );
  ANDN U352 ( .B(n7), .A(n8), .Z(n323) );
  XOR U353 ( .A(sreg[225]), .B(n324), .Z(n8) );
  XOR U354 ( .A(n326), .B(n327), .Z(n324) );
  ANDN U355 ( .B(n9), .A(n10), .Z(n326) );
  XOR U356 ( .A(sreg[224]), .B(n327), .Z(n10) );
  XOR U357 ( .A(n329), .B(n330), .Z(n327) );
  ANDN U358 ( .B(n11), .A(n12), .Z(n329) );
  XOR U359 ( .A(sreg[223]), .B(n330), .Z(n12) );
  XOR U360 ( .A(n332), .B(n333), .Z(n330) );
  ANDN U361 ( .B(n13), .A(n14), .Z(n332) );
  XOR U362 ( .A(sreg[222]), .B(n333), .Z(n14) );
  XOR U363 ( .A(n335), .B(n336), .Z(n333) );
  ANDN U364 ( .B(n15), .A(n16), .Z(n335) );
  XOR U365 ( .A(sreg[221]), .B(n336), .Z(n16) );
  XOR U366 ( .A(n338), .B(n339), .Z(n336) );
  ANDN U367 ( .B(n17), .A(n18), .Z(n338) );
  XOR U368 ( .A(sreg[220]), .B(n339), .Z(n18) );
  XOR U369 ( .A(n341), .B(n342), .Z(n339) );
  ANDN U370 ( .B(n19), .A(n20), .Z(n341) );
  XOR U371 ( .A(sreg[219]), .B(n342), .Z(n20) );
  XOR U372 ( .A(n344), .B(n345), .Z(n342) );
  ANDN U373 ( .B(n21), .A(n22), .Z(n344) );
  XOR U374 ( .A(sreg[218]), .B(n345), .Z(n22) );
  XOR U375 ( .A(n347), .B(n348), .Z(n345) );
  ANDN U376 ( .B(n25), .A(n26), .Z(n347) );
  XOR U377 ( .A(sreg[217]), .B(n348), .Z(n26) );
  XOR U378 ( .A(n350), .B(n351), .Z(n348) );
  ANDN U379 ( .B(n27), .A(n28), .Z(n350) );
  XOR U380 ( .A(sreg[216]), .B(n351), .Z(n28) );
  XOR U381 ( .A(n353), .B(n354), .Z(n351) );
  ANDN U382 ( .B(n29), .A(n30), .Z(n353) );
  XOR U383 ( .A(sreg[215]), .B(n354), .Z(n30) );
  XOR U384 ( .A(n356), .B(n357), .Z(n354) );
  ANDN U385 ( .B(n31), .A(n32), .Z(n356) );
  XOR U386 ( .A(sreg[214]), .B(n357), .Z(n32) );
  XOR U387 ( .A(n359), .B(n360), .Z(n357) );
  ANDN U388 ( .B(n33), .A(n34), .Z(n359) );
  XOR U389 ( .A(sreg[213]), .B(n360), .Z(n34) );
  XOR U390 ( .A(n362), .B(n363), .Z(n360) );
  ANDN U391 ( .B(n35), .A(n36), .Z(n362) );
  XOR U392 ( .A(sreg[212]), .B(n363), .Z(n36) );
  XOR U393 ( .A(n365), .B(n366), .Z(n363) );
  ANDN U394 ( .B(n37), .A(n38), .Z(n365) );
  XOR U395 ( .A(sreg[211]), .B(n366), .Z(n38) );
  XOR U396 ( .A(n368), .B(n369), .Z(n366) );
  ANDN U397 ( .B(n39), .A(n40), .Z(n368) );
  XOR U398 ( .A(sreg[210]), .B(n369), .Z(n40) );
  XOR U399 ( .A(n371), .B(n372), .Z(n369) );
  ANDN U400 ( .B(n41), .A(n42), .Z(n371) );
  XOR U401 ( .A(sreg[209]), .B(n372), .Z(n42) );
  XOR U402 ( .A(n374), .B(n375), .Z(n372) );
  ANDN U403 ( .B(n43), .A(n44), .Z(n374) );
  XOR U404 ( .A(sreg[208]), .B(n375), .Z(n44) );
  XOR U405 ( .A(n377), .B(n378), .Z(n375) );
  ANDN U406 ( .B(n47), .A(n48), .Z(n377) );
  XOR U407 ( .A(sreg[207]), .B(n378), .Z(n48) );
  XOR U408 ( .A(n380), .B(n381), .Z(n378) );
  ANDN U409 ( .B(n49), .A(n50), .Z(n380) );
  XOR U410 ( .A(sreg[206]), .B(n381), .Z(n50) );
  XOR U411 ( .A(n383), .B(n384), .Z(n381) );
  ANDN U412 ( .B(n51), .A(n52), .Z(n383) );
  XOR U413 ( .A(sreg[205]), .B(n384), .Z(n52) );
  XOR U414 ( .A(n386), .B(n387), .Z(n384) );
  ANDN U415 ( .B(n53), .A(n54), .Z(n386) );
  XOR U416 ( .A(sreg[204]), .B(n387), .Z(n54) );
  XOR U417 ( .A(n389), .B(n390), .Z(n387) );
  ANDN U418 ( .B(n55), .A(n56), .Z(n389) );
  XOR U419 ( .A(sreg[203]), .B(n390), .Z(n56) );
  XOR U420 ( .A(n392), .B(n393), .Z(n390) );
  ANDN U421 ( .B(n57), .A(n58), .Z(n392) );
  XOR U422 ( .A(sreg[202]), .B(n393), .Z(n58) );
  XOR U423 ( .A(n395), .B(n396), .Z(n393) );
  ANDN U424 ( .B(n59), .A(n60), .Z(n395) );
  XOR U425 ( .A(sreg[201]), .B(n396), .Z(n60) );
  XOR U426 ( .A(n398), .B(n399), .Z(n396) );
  ANDN U427 ( .B(n61), .A(n62), .Z(n398) );
  XOR U428 ( .A(sreg[200]), .B(n399), .Z(n62) );
  XOR U429 ( .A(n401), .B(n402), .Z(n399) );
  ANDN U430 ( .B(n63), .A(n64), .Z(n401) );
  XOR U431 ( .A(sreg[199]), .B(n402), .Z(n64) );
  XOR U432 ( .A(n404), .B(n405), .Z(n402) );
  ANDN U433 ( .B(n65), .A(n66), .Z(n404) );
  XOR U434 ( .A(sreg[198]), .B(n405), .Z(n66) );
  XOR U435 ( .A(n407), .B(n408), .Z(n405) );
  ANDN U436 ( .B(n69), .A(n70), .Z(n407) );
  XOR U437 ( .A(sreg[197]), .B(n408), .Z(n70) );
  XOR U438 ( .A(n410), .B(n411), .Z(n408) );
  ANDN U439 ( .B(n71), .A(n72), .Z(n410) );
  XOR U440 ( .A(sreg[196]), .B(n411), .Z(n72) );
  XOR U441 ( .A(n413), .B(n414), .Z(n411) );
  ANDN U442 ( .B(n73), .A(n74), .Z(n413) );
  XOR U443 ( .A(sreg[195]), .B(n414), .Z(n74) );
  XOR U444 ( .A(n416), .B(n417), .Z(n414) );
  ANDN U445 ( .B(n75), .A(n76), .Z(n416) );
  XOR U446 ( .A(sreg[194]), .B(n417), .Z(n76) );
  XOR U447 ( .A(n419), .B(n420), .Z(n417) );
  ANDN U448 ( .B(n77), .A(n78), .Z(n419) );
  XOR U449 ( .A(sreg[193]), .B(n420), .Z(n78) );
  XOR U450 ( .A(n422), .B(n423), .Z(n420) );
  ANDN U451 ( .B(n79), .A(n80), .Z(n422) );
  XOR U452 ( .A(sreg[192]), .B(n423), .Z(n80) );
  XOR U453 ( .A(n425), .B(n426), .Z(n423) );
  ANDN U454 ( .B(n81), .A(n82), .Z(n425) );
  XOR U455 ( .A(sreg[191]), .B(n426), .Z(n82) );
  XOR U456 ( .A(n428), .B(n429), .Z(n426) );
  ANDN U457 ( .B(n83), .A(n84), .Z(n428) );
  XOR U458 ( .A(sreg[190]), .B(n429), .Z(n84) );
  XOR U459 ( .A(n431), .B(n432), .Z(n429) );
  ANDN U460 ( .B(n85), .A(n86), .Z(n431) );
  XOR U461 ( .A(sreg[189]), .B(n432), .Z(n86) );
  XOR U462 ( .A(n434), .B(n435), .Z(n432) );
  ANDN U463 ( .B(n87), .A(n88), .Z(n434) );
  XOR U464 ( .A(sreg[188]), .B(n435), .Z(n88) );
  XOR U465 ( .A(n437), .B(n438), .Z(n435) );
  ANDN U466 ( .B(n91), .A(n92), .Z(n437) );
  XOR U467 ( .A(sreg[187]), .B(n438), .Z(n92) );
  XOR U468 ( .A(n440), .B(n441), .Z(n438) );
  ANDN U469 ( .B(n93), .A(n94), .Z(n440) );
  XOR U470 ( .A(sreg[186]), .B(n441), .Z(n94) );
  XOR U471 ( .A(n443), .B(n444), .Z(n441) );
  ANDN U472 ( .B(n95), .A(n96), .Z(n443) );
  XOR U473 ( .A(sreg[185]), .B(n444), .Z(n96) );
  XOR U474 ( .A(n446), .B(n447), .Z(n444) );
  ANDN U475 ( .B(n97), .A(n98), .Z(n446) );
  XOR U476 ( .A(sreg[184]), .B(n447), .Z(n98) );
  XOR U477 ( .A(n449), .B(n450), .Z(n447) );
  ANDN U478 ( .B(n99), .A(n100), .Z(n449) );
  XOR U479 ( .A(sreg[183]), .B(n450), .Z(n100) );
  XOR U480 ( .A(n452), .B(n453), .Z(n450) );
  ANDN U481 ( .B(n101), .A(n102), .Z(n452) );
  XOR U482 ( .A(sreg[182]), .B(n453), .Z(n102) );
  XOR U483 ( .A(n455), .B(n456), .Z(n453) );
  ANDN U484 ( .B(n103), .A(n104), .Z(n455) );
  XOR U485 ( .A(sreg[181]), .B(n456), .Z(n104) );
  XOR U486 ( .A(n458), .B(n459), .Z(n456) );
  ANDN U487 ( .B(n105), .A(n106), .Z(n458) );
  XOR U488 ( .A(sreg[180]), .B(n459), .Z(n106) );
  XOR U489 ( .A(n461), .B(n462), .Z(n459) );
  ANDN U490 ( .B(n107), .A(n108), .Z(n461) );
  XOR U491 ( .A(sreg[179]), .B(n462), .Z(n108) );
  XOR U492 ( .A(n464), .B(n465), .Z(n462) );
  ANDN U493 ( .B(n109), .A(n110), .Z(n464) );
  XOR U494 ( .A(sreg[178]), .B(n465), .Z(n110) );
  XOR U495 ( .A(n467), .B(n468), .Z(n465) );
  ANDN U496 ( .B(n113), .A(n114), .Z(n467) );
  XOR U497 ( .A(sreg[177]), .B(n468), .Z(n114) );
  XOR U498 ( .A(n470), .B(n471), .Z(n468) );
  ANDN U499 ( .B(n115), .A(n116), .Z(n470) );
  XOR U500 ( .A(sreg[176]), .B(n471), .Z(n116) );
  XOR U501 ( .A(n473), .B(n474), .Z(n471) );
  ANDN U502 ( .B(n117), .A(n118), .Z(n473) );
  XOR U503 ( .A(sreg[175]), .B(n474), .Z(n118) );
  XOR U504 ( .A(n476), .B(n477), .Z(n474) );
  ANDN U505 ( .B(n119), .A(n120), .Z(n476) );
  XOR U506 ( .A(sreg[174]), .B(n477), .Z(n120) );
  XOR U507 ( .A(n479), .B(n480), .Z(n477) );
  ANDN U508 ( .B(n121), .A(n122), .Z(n479) );
  XOR U509 ( .A(sreg[173]), .B(n480), .Z(n122) );
  XOR U510 ( .A(n482), .B(n483), .Z(n480) );
  ANDN U511 ( .B(n123), .A(n124), .Z(n482) );
  XOR U512 ( .A(sreg[172]), .B(n483), .Z(n124) );
  XOR U513 ( .A(n485), .B(n486), .Z(n483) );
  ANDN U514 ( .B(n125), .A(n126), .Z(n485) );
  XOR U515 ( .A(sreg[171]), .B(n486), .Z(n126) );
  XOR U516 ( .A(n488), .B(n489), .Z(n486) );
  ANDN U517 ( .B(n127), .A(n128), .Z(n488) );
  XOR U518 ( .A(sreg[170]), .B(n489), .Z(n128) );
  XOR U519 ( .A(n491), .B(n492), .Z(n489) );
  ANDN U520 ( .B(n129), .A(n130), .Z(n491) );
  XOR U521 ( .A(sreg[169]), .B(n492), .Z(n130) );
  XOR U522 ( .A(n494), .B(n495), .Z(n492) );
  ANDN U523 ( .B(n131), .A(n132), .Z(n494) );
  XOR U524 ( .A(sreg[168]), .B(n495), .Z(n132) );
  XOR U525 ( .A(n497), .B(n498), .Z(n495) );
  ANDN U526 ( .B(n135), .A(n136), .Z(n497) );
  XOR U527 ( .A(sreg[167]), .B(n498), .Z(n136) );
  XOR U528 ( .A(n500), .B(n501), .Z(n498) );
  ANDN U529 ( .B(n137), .A(n138), .Z(n500) );
  XOR U530 ( .A(sreg[166]), .B(n501), .Z(n138) );
  XOR U531 ( .A(n503), .B(n504), .Z(n501) );
  ANDN U532 ( .B(n139), .A(n140), .Z(n503) );
  XOR U533 ( .A(sreg[165]), .B(n504), .Z(n140) );
  XOR U534 ( .A(n506), .B(n507), .Z(n504) );
  ANDN U535 ( .B(n141), .A(n142), .Z(n506) );
  XOR U536 ( .A(sreg[164]), .B(n507), .Z(n142) );
  XOR U537 ( .A(n509), .B(n510), .Z(n507) );
  ANDN U538 ( .B(n143), .A(n144), .Z(n509) );
  XOR U539 ( .A(sreg[163]), .B(n510), .Z(n144) );
  XOR U540 ( .A(n512), .B(n513), .Z(n510) );
  ANDN U541 ( .B(n145), .A(n146), .Z(n512) );
  XOR U542 ( .A(sreg[162]), .B(n513), .Z(n146) );
  XOR U543 ( .A(n515), .B(n516), .Z(n513) );
  ANDN U544 ( .B(n147), .A(n148), .Z(n515) );
  XOR U545 ( .A(sreg[161]), .B(n516), .Z(n148) );
  XOR U546 ( .A(n518), .B(n519), .Z(n516) );
  ANDN U547 ( .B(n149), .A(n150), .Z(n518) );
  XOR U548 ( .A(sreg[160]), .B(n519), .Z(n150) );
  XOR U549 ( .A(n521), .B(n522), .Z(n519) );
  ANDN U550 ( .B(n151), .A(n152), .Z(n521) );
  XOR U551 ( .A(sreg[159]), .B(n522), .Z(n152) );
  XOR U552 ( .A(n524), .B(n525), .Z(n522) );
  ANDN U553 ( .B(n153), .A(n154), .Z(n524) );
  XOR U554 ( .A(sreg[158]), .B(n525), .Z(n154) );
  XOR U555 ( .A(n527), .B(n528), .Z(n525) );
  ANDN U556 ( .B(n157), .A(n158), .Z(n527) );
  XOR U557 ( .A(sreg[157]), .B(n528), .Z(n158) );
  XOR U558 ( .A(n530), .B(n531), .Z(n528) );
  ANDN U559 ( .B(n159), .A(n160), .Z(n530) );
  XOR U560 ( .A(sreg[156]), .B(n531), .Z(n160) );
  XOR U561 ( .A(n533), .B(n534), .Z(n531) );
  ANDN U562 ( .B(n161), .A(n162), .Z(n533) );
  XOR U563 ( .A(sreg[155]), .B(n534), .Z(n162) );
  XOR U564 ( .A(n536), .B(n537), .Z(n534) );
  ANDN U565 ( .B(n163), .A(n164), .Z(n536) );
  XOR U566 ( .A(sreg[154]), .B(n537), .Z(n164) );
  XOR U567 ( .A(n539), .B(n540), .Z(n537) );
  ANDN U568 ( .B(n165), .A(n166), .Z(n539) );
  XOR U569 ( .A(sreg[153]), .B(n540), .Z(n166) );
  XOR U570 ( .A(n542), .B(n543), .Z(n540) );
  ANDN U571 ( .B(n167), .A(n168), .Z(n542) );
  XOR U572 ( .A(sreg[152]), .B(n543), .Z(n168) );
  XOR U573 ( .A(n545), .B(n546), .Z(n543) );
  ANDN U574 ( .B(n169), .A(n170), .Z(n545) );
  XOR U575 ( .A(sreg[151]), .B(n546), .Z(n170) );
  XOR U576 ( .A(n548), .B(n549), .Z(n546) );
  ANDN U577 ( .B(n171), .A(n172), .Z(n548) );
  XOR U578 ( .A(sreg[150]), .B(n549), .Z(n172) );
  XOR U579 ( .A(n551), .B(n552), .Z(n549) );
  ANDN U580 ( .B(n173), .A(n174), .Z(n551) );
  XOR U581 ( .A(sreg[149]), .B(n552), .Z(n174) );
  XOR U582 ( .A(n554), .B(n555), .Z(n552) );
  ANDN U583 ( .B(n175), .A(n176), .Z(n554) );
  XOR U584 ( .A(sreg[148]), .B(n555), .Z(n176) );
  XOR U585 ( .A(n557), .B(n558), .Z(n555) );
  ANDN U586 ( .B(n179), .A(n180), .Z(n557) );
  XOR U587 ( .A(sreg[147]), .B(n558), .Z(n180) );
  XOR U588 ( .A(n560), .B(n561), .Z(n558) );
  ANDN U589 ( .B(n181), .A(n182), .Z(n560) );
  XOR U590 ( .A(sreg[146]), .B(n561), .Z(n182) );
  XOR U591 ( .A(n563), .B(n564), .Z(n561) );
  ANDN U592 ( .B(n183), .A(n184), .Z(n563) );
  XOR U593 ( .A(sreg[145]), .B(n564), .Z(n184) );
  XOR U594 ( .A(n566), .B(n567), .Z(n564) );
  ANDN U595 ( .B(n185), .A(n186), .Z(n566) );
  XOR U596 ( .A(sreg[144]), .B(n567), .Z(n186) );
  XOR U597 ( .A(n569), .B(n570), .Z(n567) );
  ANDN U598 ( .B(n187), .A(n188), .Z(n569) );
  XOR U599 ( .A(sreg[143]), .B(n570), .Z(n188) );
  XOR U600 ( .A(n572), .B(n573), .Z(n570) );
  ANDN U601 ( .B(n189), .A(n190), .Z(n572) );
  XOR U602 ( .A(sreg[142]), .B(n573), .Z(n190) );
  XOR U603 ( .A(n575), .B(n576), .Z(n573) );
  ANDN U604 ( .B(n191), .A(n192), .Z(n575) );
  XOR U605 ( .A(sreg[141]), .B(n576), .Z(n192) );
  XOR U606 ( .A(n578), .B(n579), .Z(n576) );
  ANDN U607 ( .B(n193), .A(n194), .Z(n578) );
  XOR U608 ( .A(sreg[140]), .B(n579), .Z(n194) );
  XOR U609 ( .A(n581), .B(n582), .Z(n579) );
  ANDN U610 ( .B(n217), .A(n218), .Z(n581) );
  XOR U611 ( .A(sreg[139]), .B(n582), .Z(n218) );
  XOR U612 ( .A(n584), .B(n585), .Z(n582) );
  ANDN U613 ( .B(n269), .A(n270), .Z(n584) );
  XOR U614 ( .A(sreg[138]), .B(n585), .Z(n270) );
  XOR U615 ( .A(n587), .B(n588), .Z(n585) );
  ANDN U616 ( .B(n2), .A(n1), .Z(n587) );
  XOR U617 ( .A(sreg[137]), .B(n588), .Z(n1) );
  XOR U618 ( .A(n590), .B(n591), .Z(n588) );
  ANDN U619 ( .B(n23), .A(n24), .Z(n590) );
  XOR U620 ( .A(sreg[136]), .B(n591), .Z(n24) );
  XOR U621 ( .A(n593), .B(n594), .Z(n591) );
  ANDN U622 ( .B(n45), .A(n46), .Z(n593) );
  XOR U623 ( .A(sreg[135]), .B(n594), .Z(n46) );
  XOR U624 ( .A(n596), .B(n597), .Z(n594) );
  ANDN U625 ( .B(n67), .A(n68), .Z(n596) );
  XOR U626 ( .A(sreg[134]), .B(n597), .Z(n68) );
  XOR U627 ( .A(n599), .B(n600), .Z(n597) );
  ANDN U628 ( .B(n89), .A(n90), .Z(n599) );
  XOR U629 ( .A(sreg[133]), .B(n600), .Z(n90) );
  XOR U630 ( .A(n602), .B(n603), .Z(n600) );
  ANDN U631 ( .B(n111), .A(n112), .Z(n602) );
  XOR U632 ( .A(sreg[132]), .B(n603), .Z(n112) );
  XOR U633 ( .A(n605), .B(n606), .Z(n603) );
  ANDN U634 ( .B(n133), .A(n134), .Z(n605) );
  XOR U635 ( .A(sreg[131]), .B(n606), .Z(n134) );
  XOR U636 ( .A(n608), .B(n609), .Z(n606) );
  NOR U637 ( .A(n156), .B(n155), .Z(n608) );
  AND U638 ( .A(a[2]), .B(b[0]), .Z(n610) );
  XOR U639 ( .A(sreg[130]), .B(n609), .Z(n156) );
  XOR U640 ( .A(n611), .B(n612), .Z(n609) );
  NAND U641 ( .A(n177), .B(n178), .Z(n612) );
  XOR U642 ( .A(sreg[129]), .B(n611), .Z(n178) );
  XNOR U643 ( .A(n611), .B(n613), .Z(n177) );
  NAND U644 ( .A(b[0]), .B(a[1]), .Z(n613) );
  ANDN U645 ( .B(sreg[128]), .A(n614), .Z(n611) );
  AND U646 ( .A(a[3]), .B(b[0]), .Z(n607) );
  AND U647 ( .A(a[4]), .B(b[0]), .Z(n604) );
  AND U648 ( .A(a[5]), .B(b[0]), .Z(n601) );
  AND U649 ( .A(a[6]), .B(b[0]), .Z(n598) );
  AND U650 ( .A(a[7]), .B(b[0]), .Z(n595) );
  AND U651 ( .A(a[8]), .B(b[0]), .Z(n592) );
  AND U652 ( .A(a[9]), .B(b[0]), .Z(n589) );
  AND U653 ( .A(a[10]), .B(b[0]), .Z(n586) );
  AND U654 ( .A(a[11]), .B(b[0]), .Z(n583) );
  AND U655 ( .A(a[12]), .B(b[0]), .Z(n580) );
  AND U656 ( .A(a[13]), .B(b[0]), .Z(n577) );
  AND U657 ( .A(a[14]), .B(b[0]), .Z(n574) );
  AND U658 ( .A(a[15]), .B(b[0]), .Z(n571) );
  AND U659 ( .A(a[16]), .B(b[0]), .Z(n568) );
  AND U660 ( .A(a[17]), .B(b[0]), .Z(n565) );
  AND U661 ( .A(a[18]), .B(b[0]), .Z(n562) );
  AND U662 ( .A(a[19]), .B(b[0]), .Z(n559) );
  AND U663 ( .A(a[20]), .B(b[0]), .Z(n556) );
  AND U664 ( .A(a[21]), .B(b[0]), .Z(n553) );
  AND U665 ( .A(a[22]), .B(b[0]), .Z(n550) );
  AND U666 ( .A(a[23]), .B(b[0]), .Z(n547) );
  AND U667 ( .A(a[24]), .B(b[0]), .Z(n544) );
  AND U668 ( .A(a[25]), .B(b[0]), .Z(n541) );
  AND U669 ( .A(a[26]), .B(b[0]), .Z(n538) );
  AND U670 ( .A(a[27]), .B(b[0]), .Z(n535) );
  AND U671 ( .A(a[28]), .B(b[0]), .Z(n532) );
  AND U672 ( .A(a[29]), .B(b[0]), .Z(n529) );
  AND U673 ( .A(a[30]), .B(b[0]), .Z(n526) );
  AND U674 ( .A(a[31]), .B(b[0]), .Z(n523) );
  AND U675 ( .A(a[32]), .B(b[0]), .Z(n520) );
  AND U676 ( .A(a[33]), .B(b[0]), .Z(n517) );
  AND U677 ( .A(a[34]), .B(b[0]), .Z(n514) );
  AND U678 ( .A(a[35]), .B(b[0]), .Z(n511) );
  AND U679 ( .A(a[36]), .B(b[0]), .Z(n508) );
  AND U680 ( .A(a[37]), .B(b[0]), .Z(n505) );
  AND U681 ( .A(a[38]), .B(b[0]), .Z(n502) );
  AND U682 ( .A(a[39]), .B(b[0]), .Z(n499) );
  AND U683 ( .A(a[40]), .B(b[0]), .Z(n496) );
  AND U684 ( .A(a[41]), .B(b[0]), .Z(n493) );
  AND U685 ( .A(a[42]), .B(b[0]), .Z(n490) );
  AND U686 ( .A(a[43]), .B(b[0]), .Z(n487) );
  AND U687 ( .A(a[44]), .B(b[0]), .Z(n484) );
  AND U688 ( .A(a[45]), .B(b[0]), .Z(n481) );
  AND U689 ( .A(a[46]), .B(b[0]), .Z(n478) );
  AND U690 ( .A(a[47]), .B(b[0]), .Z(n475) );
  AND U691 ( .A(a[48]), .B(b[0]), .Z(n472) );
  AND U692 ( .A(a[49]), .B(b[0]), .Z(n469) );
  AND U693 ( .A(a[50]), .B(b[0]), .Z(n466) );
  AND U694 ( .A(a[51]), .B(b[0]), .Z(n463) );
  AND U695 ( .A(a[52]), .B(b[0]), .Z(n460) );
  AND U696 ( .A(a[53]), .B(b[0]), .Z(n457) );
  AND U697 ( .A(a[54]), .B(b[0]), .Z(n454) );
  AND U698 ( .A(a[55]), .B(b[0]), .Z(n451) );
  AND U699 ( .A(a[56]), .B(b[0]), .Z(n448) );
  AND U700 ( .A(a[57]), .B(b[0]), .Z(n445) );
  AND U701 ( .A(a[58]), .B(b[0]), .Z(n442) );
  AND U702 ( .A(a[59]), .B(b[0]), .Z(n439) );
  AND U703 ( .A(a[60]), .B(b[0]), .Z(n436) );
  AND U704 ( .A(a[61]), .B(b[0]), .Z(n433) );
  AND U705 ( .A(a[62]), .B(b[0]), .Z(n430) );
  AND U706 ( .A(a[63]), .B(b[0]), .Z(n427) );
  AND U707 ( .A(a[64]), .B(b[0]), .Z(n424) );
  AND U708 ( .A(a[65]), .B(b[0]), .Z(n421) );
  AND U709 ( .A(a[66]), .B(b[0]), .Z(n418) );
  AND U710 ( .A(a[67]), .B(b[0]), .Z(n415) );
  AND U711 ( .A(a[68]), .B(b[0]), .Z(n412) );
  AND U712 ( .A(a[69]), .B(b[0]), .Z(n409) );
  AND U713 ( .A(a[70]), .B(b[0]), .Z(n406) );
  AND U714 ( .A(a[71]), .B(b[0]), .Z(n403) );
  AND U715 ( .A(a[72]), .B(b[0]), .Z(n400) );
  AND U716 ( .A(a[73]), .B(b[0]), .Z(n397) );
  AND U717 ( .A(a[74]), .B(b[0]), .Z(n394) );
  AND U718 ( .A(a[75]), .B(b[0]), .Z(n391) );
  AND U719 ( .A(a[76]), .B(b[0]), .Z(n388) );
  AND U720 ( .A(a[77]), .B(b[0]), .Z(n385) );
  AND U721 ( .A(a[78]), .B(b[0]), .Z(n382) );
  AND U722 ( .A(a[79]), .B(b[0]), .Z(n379) );
  AND U723 ( .A(a[80]), .B(b[0]), .Z(n376) );
  AND U724 ( .A(a[81]), .B(b[0]), .Z(n373) );
  AND U725 ( .A(a[82]), .B(b[0]), .Z(n370) );
  AND U726 ( .A(a[83]), .B(b[0]), .Z(n367) );
  AND U727 ( .A(a[84]), .B(b[0]), .Z(n364) );
  AND U728 ( .A(a[85]), .B(b[0]), .Z(n361) );
  AND U729 ( .A(a[86]), .B(b[0]), .Z(n358) );
  AND U730 ( .A(a[87]), .B(b[0]), .Z(n355) );
  AND U731 ( .A(a[88]), .B(b[0]), .Z(n352) );
  AND U732 ( .A(a[89]), .B(b[0]), .Z(n349) );
  AND U733 ( .A(a[90]), .B(b[0]), .Z(n346) );
  AND U734 ( .A(a[91]), .B(b[0]), .Z(n343) );
  AND U735 ( .A(a[92]), .B(b[0]), .Z(n340) );
  AND U736 ( .A(a[93]), .B(b[0]), .Z(n337) );
  AND U737 ( .A(a[94]), .B(b[0]), .Z(n334) );
  AND U738 ( .A(a[95]), .B(b[0]), .Z(n331) );
  AND U739 ( .A(a[96]), .B(b[0]), .Z(n328) );
  AND U740 ( .A(a[97]), .B(b[0]), .Z(n325) );
  AND U741 ( .A(a[98]), .B(b[0]), .Z(n322) );
  AND U742 ( .A(a[99]), .B(b[0]), .Z(n319) );
  AND U743 ( .A(a[100]), .B(b[0]), .Z(n316) );
  XNOR U744 ( .A(sreg[128]), .B(n614), .Z(c[127]) );
  NAND U745 ( .A(a[0]), .B(b[0]), .Z(n614) );
endmodule

